//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 0 0 0 1 1 1 1 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 0 0 0 1 1 0 1 1 0 0 0 0 0 0 1 1 0 1 1 1 0 1 0 1 0 0 1 0 0 0 1 1 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:26:59 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n694, new_n695, new_n696,
    new_n697, new_n698, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n710, new_n711, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n719, new_n720, new_n721,
    new_n722, new_n723, new_n724, new_n725, new_n727, new_n728, new_n729,
    new_n730, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n758, new_n759,
    new_n760, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n789,
    new_n790, new_n791, new_n792, new_n793, new_n794, new_n795, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n912, new_n913, new_n914, new_n915, new_n916, new_n917,
    new_n918, new_n919, new_n920, new_n921, new_n922, new_n923, new_n924,
    new_n925, new_n926, new_n927, new_n928, new_n929, new_n930, new_n931,
    new_n932, new_n933, new_n934, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n948, new_n949, new_n950, new_n952, new_n953, new_n954, new_n955,
    new_n956, new_n957, new_n958, new_n959, new_n960, new_n961, new_n962,
    new_n963, new_n964, new_n965, new_n966, new_n967, new_n968, new_n970,
    new_n971, new_n972, new_n973, new_n974, new_n975, new_n976, new_n977,
    new_n978, new_n979, new_n980, new_n981, new_n982, new_n983, new_n984,
    new_n985, new_n986, new_n987, new_n989, new_n990, new_n991, new_n992,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1017, new_n1018,
    new_n1019, new_n1021, new_n1022, new_n1023, new_n1024, new_n1025,
    new_n1026, new_n1027, new_n1028, new_n1029, new_n1030, new_n1031,
    new_n1032, new_n1033;
  INV_X1    g000(.A(G221), .ZN(new_n187));
  XNOR2_X1  g001(.A(KEYINPUT9), .B(G234), .ZN(new_n188));
  INV_X1    g002(.A(new_n188), .ZN(new_n189));
  INV_X1    g003(.A(G902), .ZN(new_n190));
  AOI21_X1  g004(.A(new_n187), .B1(new_n189), .B2(new_n190), .ZN(new_n191));
  INV_X1    g005(.A(new_n191), .ZN(new_n192));
  INV_X1    g006(.A(KEYINPUT76), .ZN(new_n193));
  INV_X1    g007(.A(G107), .ZN(new_n194));
  OAI21_X1  g008(.A(new_n193), .B1(new_n194), .B2(G104), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n194), .A2(G104), .ZN(new_n196));
  INV_X1    g010(.A(G104), .ZN(new_n197));
  NAND3_X1  g011(.A1(new_n197), .A2(KEYINPUT76), .A3(G107), .ZN(new_n198));
  NAND3_X1  g012(.A1(new_n195), .A2(new_n196), .A3(new_n198), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n199), .A2(G101), .ZN(new_n200));
  INV_X1    g014(.A(G101), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n197), .A2(G107), .ZN(new_n202));
  AND3_X1   g016(.A1(new_n194), .A2(KEYINPUT3), .A3(G104), .ZN(new_n203));
  AOI21_X1  g017(.A(KEYINPUT3), .B1(new_n194), .B2(G104), .ZN(new_n204));
  OAI211_X1 g018(.A(new_n201), .B(new_n202), .C1(new_n203), .C2(new_n204), .ZN(new_n205));
  NAND3_X1  g019(.A1(new_n200), .A2(new_n205), .A3(KEYINPUT77), .ZN(new_n206));
  INV_X1    g020(.A(KEYINPUT77), .ZN(new_n207));
  NAND3_X1  g021(.A1(new_n199), .A2(new_n207), .A3(G101), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n206), .A2(new_n208), .ZN(new_n209));
  INV_X1    g023(.A(G119), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n210), .A2(G116), .ZN(new_n211));
  OR2_X1    g025(.A1(new_n211), .A2(KEYINPUT5), .ZN(new_n212));
  AND2_X1   g026(.A1(new_n212), .A2(G113), .ZN(new_n213));
  XNOR2_X1  g027(.A(G116), .B(G119), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n214), .A2(KEYINPUT5), .ZN(new_n215));
  XOR2_X1   g029(.A(KEYINPUT2), .B(G113), .Z(new_n216));
  AOI22_X1  g030(.A1(new_n213), .A2(new_n215), .B1(new_n214), .B2(new_n216), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n209), .A2(new_n217), .ZN(new_n218));
  INV_X1    g032(.A(KEYINPUT3), .ZN(new_n219));
  OAI21_X1  g033(.A(new_n219), .B1(new_n197), .B2(G107), .ZN(new_n220));
  NAND3_X1  g034(.A1(new_n194), .A2(KEYINPUT3), .A3(G104), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n220), .A2(new_n221), .ZN(new_n222));
  AOI21_X1  g036(.A(new_n201), .B1(new_n222), .B2(new_n202), .ZN(new_n223));
  INV_X1    g037(.A(KEYINPUT4), .ZN(new_n224));
  NAND2_X1  g038(.A1(new_n216), .A2(new_n214), .ZN(new_n225));
  INV_X1    g039(.A(G116), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n226), .A2(G119), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n211), .A2(new_n227), .ZN(new_n228));
  XNOR2_X1  g042(.A(KEYINPUT2), .B(G113), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n228), .A2(new_n229), .ZN(new_n230));
  AOI22_X1  g044(.A1(new_n223), .A2(new_n224), .B1(new_n225), .B2(new_n230), .ZN(new_n231));
  OAI21_X1  g045(.A(new_n202), .B1(new_n203), .B2(new_n204), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n232), .A2(G101), .ZN(new_n233));
  NAND3_X1  g047(.A1(new_n233), .A2(KEYINPUT4), .A3(new_n205), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n231), .A2(new_n234), .ZN(new_n235));
  XNOR2_X1  g049(.A(G110), .B(G122), .ZN(new_n236));
  NAND3_X1  g050(.A1(new_n218), .A2(new_n235), .A3(new_n236), .ZN(new_n237));
  AOI22_X1  g051(.A1(new_n209), .A2(new_n217), .B1(new_n231), .B2(new_n234), .ZN(new_n238));
  XOR2_X1   g052(.A(new_n236), .B(KEYINPUT83), .Z(new_n239));
  OAI211_X1 g053(.A(new_n237), .B(KEYINPUT6), .C1(new_n238), .C2(new_n239), .ZN(new_n240));
  INV_X1    g054(.A(G146), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n241), .A2(G143), .ZN(new_n242));
  INV_X1    g056(.A(G143), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n243), .A2(G146), .ZN(new_n244));
  NAND4_X1  g058(.A1(new_n242), .A2(new_n244), .A3(KEYINPUT0), .A4(G128), .ZN(new_n245));
  XNOR2_X1  g059(.A(G143), .B(G146), .ZN(new_n246));
  XNOR2_X1  g060(.A(KEYINPUT0), .B(G128), .ZN(new_n247));
  OAI21_X1  g061(.A(new_n245), .B1(new_n246), .B2(new_n247), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n248), .A2(G125), .ZN(new_n249));
  OAI21_X1  g063(.A(KEYINPUT1), .B1(new_n243), .B2(G146), .ZN(new_n250));
  NOR2_X1   g064(.A1(new_n243), .A2(G146), .ZN(new_n251));
  NOR2_X1   g065(.A1(new_n241), .A2(G143), .ZN(new_n252));
  OAI211_X1 g066(.A(G128), .B(new_n250), .C1(new_n251), .C2(new_n252), .ZN(new_n253));
  INV_X1    g067(.A(G128), .ZN(new_n254));
  OAI211_X1 g068(.A(new_n242), .B(new_n244), .C1(KEYINPUT1), .C2(new_n254), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n253), .A2(new_n255), .ZN(new_n256));
  INV_X1    g070(.A(new_n256), .ZN(new_n257));
  OAI21_X1  g071(.A(new_n249), .B1(new_n257), .B2(G125), .ZN(new_n258));
  INV_X1    g072(.A(G224), .ZN(new_n259));
  NOR2_X1   g073(.A1(new_n259), .A2(G953), .ZN(new_n260));
  XNOR2_X1  g074(.A(new_n258), .B(new_n260), .ZN(new_n261));
  INV_X1    g075(.A(KEYINPUT84), .ZN(new_n262));
  AOI21_X1  g076(.A(new_n239), .B1(new_n218), .B2(new_n235), .ZN(new_n263));
  INV_X1    g077(.A(KEYINPUT6), .ZN(new_n264));
  AOI21_X1  g078(.A(new_n262), .B1(new_n263), .B2(new_n264), .ZN(new_n265));
  NOR4_X1   g079(.A1(new_n238), .A2(KEYINPUT84), .A3(KEYINPUT6), .A4(new_n239), .ZN(new_n266));
  OAI211_X1 g080(.A(new_n240), .B(new_n261), .C1(new_n265), .C2(new_n266), .ZN(new_n267));
  OAI21_X1  g081(.A(KEYINPUT7), .B1(new_n259), .B2(G953), .ZN(new_n268));
  OR2_X1    g082(.A1(new_n258), .A2(new_n268), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n258), .A2(new_n268), .ZN(new_n270));
  AND3_X1   g084(.A1(new_n237), .A2(new_n269), .A3(new_n270), .ZN(new_n271));
  XNOR2_X1  g085(.A(new_n209), .B(new_n217), .ZN(new_n272));
  XNOR2_X1  g086(.A(new_n236), .B(KEYINPUT8), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n272), .A2(new_n273), .ZN(new_n274));
  AOI21_X1  g088(.A(G902), .B1(new_n271), .B2(new_n274), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n267), .A2(new_n275), .ZN(new_n276));
  OAI21_X1  g090(.A(G210), .B1(G237), .B2(G902), .ZN(new_n277));
  INV_X1    g091(.A(new_n277), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n276), .A2(new_n278), .ZN(new_n279));
  NAND3_X1  g093(.A1(new_n267), .A2(new_n275), .A3(new_n277), .ZN(new_n280));
  NAND3_X1  g094(.A1(new_n279), .A2(KEYINPUT85), .A3(new_n280), .ZN(new_n281));
  NOR2_X1   g095(.A1(new_n280), .A2(KEYINPUT85), .ZN(new_n282));
  INV_X1    g096(.A(new_n282), .ZN(new_n283));
  NAND2_X1  g097(.A1(G234), .A2(G237), .ZN(new_n284));
  INV_X1    g098(.A(G953), .ZN(new_n285));
  NAND3_X1  g099(.A1(new_n284), .A2(G952), .A3(new_n285), .ZN(new_n286));
  INV_X1    g100(.A(new_n286), .ZN(new_n287));
  NAND3_X1  g101(.A1(new_n284), .A2(G902), .A3(G953), .ZN(new_n288));
  INV_X1    g102(.A(new_n288), .ZN(new_n289));
  XNOR2_X1  g103(.A(KEYINPUT21), .B(G898), .ZN(new_n290));
  AOI21_X1  g104(.A(new_n287), .B1(new_n289), .B2(new_n290), .ZN(new_n291));
  OAI21_X1  g105(.A(G214), .B1(G237), .B2(G902), .ZN(new_n292));
  INV_X1    g106(.A(new_n292), .ZN(new_n293));
  NOR2_X1   g107(.A1(new_n291), .A2(new_n293), .ZN(new_n294));
  NAND3_X1  g108(.A1(new_n281), .A2(new_n283), .A3(new_n294), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n254), .A2(G143), .ZN(new_n296));
  OAI21_X1  g110(.A(KEYINPUT91), .B1(new_n254), .B2(G143), .ZN(new_n297));
  INV_X1    g111(.A(KEYINPUT91), .ZN(new_n298));
  NAND3_X1  g112(.A1(new_n298), .A2(new_n243), .A3(G128), .ZN(new_n299));
  AND2_X1   g113(.A1(new_n297), .A2(new_n299), .ZN(new_n300));
  OAI21_X1  g114(.A(new_n296), .B1(new_n300), .B2(KEYINPUT13), .ZN(new_n301));
  AND3_X1   g115(.A1(new_n297), .A2(new_n299), .A3(KEYINPUT13), .ZN(new_n302));
  OAI21_X1  g116(.A(G134), .B1(new_n301), .B2(new_n302), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n297), .A2(new_n299), .ZN(new_n304));
  INV_X1    g118(.A(G134), .ZN(new_n305));
  NAND3_X1  g119(.A1(new_n304), .A2(new_n305), .A3(new_n296), .ZN(new_n306));
  XNOR2_X1  g120(.A(G116), .B(G122), .ZN(new_n307));
  XNOR2_X1  g121(.A(new_n307), .B(new_n194), .ZN(new_n308));
  NAND3_X1  g122(.A1(new_n303), .A2(new_n306), .A3(new_n308), .ZN(new_n309));
  INV_X1    g123(.A(KEYINPUT14), .ZN(new_n310));
  NAND3_X1  g124(.A1(new_n310), .A2(new_n226), .A3(G122), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n311), .A2(KEYINPUT92), .ZN(new_n312));
  INV_X1    g126(.A(G122), .ZN(new_n313));
  OAI21_X1  g127(.A(KEYINPUT14), .B1(new_n313), .B2(G116), .ZN(new_n314));
  OAI211_X1 g128(.A(new_n312), .B(new_n314), .C1(new_n226), .C2(G122), .ZN(new_n315));
  NOR2_X1   g129(.A1(new_n311), .A2(KEYINPUT92), .ZN(new_n316));
  OAI21_X1  g130(.A(G107), .B1(new_n315), .B2(new_n316), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n307), .A2(new_n194), .ZN(new_n318));
  INV_X1    g132(.A(new_n306), .ZN(new_n319));
  AOI21_X1  g133(.A(new_n305), .B1(new_n304), .B2(new_n296), .ZN(new_n320));
  OAI211_X1 g134(.A(new_n317), .B(new_n318), .C1(new_n319), .C2(new_n320), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n309), .A2(new_n321), .ZN(new_n322));
  INV_X1    g136(.A(G217), .ZN(new_n323));
  NOR3_X1   g137(.A1(new_n188), .A2(new_n323), .A3(G953), .ZN(new_n324));
  INV_X1    g138(.A(new_n324), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n322), .A2(new_n325), .ZN(new_n326));
  NAND3_X1  g140(.A1(new_n309), .A2(new_n321), .A3(new_n324), .ZN(new_n327));
  AOI21_X1  g141(.A(G902), .B1(new_n326), .B2(new_n327), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n328), .A2(KEYINPUT93), .ZN(new_n329));
  INV_X1    g143(.A(G478), .ZN(new_n330));
  NOR2_X1   g144(.A1(new_n330), .A2(KEYINPUT15), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n329), .A2(new_n331), .ZN(new_n332));
  OAI211_X1 g146(.A(new_n328), .B(KEYINPUT93), .C1(KEYINPUT15), .C2(new_n330), .ZN(new_n333));
  AND2_X1   g147(.A1(new_n332), .A2(new_n333), .ZN(new_n334));
  INV_X1    g148(.A(KEYINPUT20), .ZN(new_n335));
  XNOR2_X1  g149(.A(G113), .B(G122), .ZN(new_n336));
  XNOR2_X1  g150(.A(new_n336), .B(new_n197), .ZN(new_n337));
  INV_X1    g151(.A(G237), .ZN(new_n338));
  NAND3_X1  g152(.A1(new_n338), .A2(new_n285), .A3(G214), .ZN(new_n339));
  NOR2_X1   g153(.A1(KEYINPUT86), .A2(G143), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n339), .A2(new_n340), .ZN(new_n341));
  NOR2_X1   g155(.A1(G237), .A2(G953), .ZN(new_n342));
  OAI211_X1 g156(.A(new_n342), .B(G214), .C1(KEYINPUT86), .C2(G143), .ZN(new_n343));
  NAND2_X1  g157(.A1(KEYINPUT18), .A2(G131), .ZN(new_n344));
  NAND3_X1  g158(.A1(new_n341), .A2(new_n343), .A3(new_n344), .ZN(new_n345));
  INV_X1    g159(.A(G140), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n346), .A2(G125), .ZN(new_n347));
  INV_X1    g161(.A(G125), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n348), .A2(G140), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n347), .A2(new_n349), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n350), .A2(G146), .ZN(new_n351));
  XNOR2_X1  g165(.A(G125), .B(G140), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n352), .A2(new_n241), .ZN(new_n353));
  NAND2_X1  g167(.A1(new_n351), .A2(new_n353), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n341), .A2(new_n343), .ZN(new_n355));
  INV_X1    g169(.A(new_n344), .ZN(new_n356));
  AOI21_X1  g170(.A(KEYINPUT87), .B1(new_n355), .B2(new_n356), .ZN(new_n357));
  INV_X1    g171(.A(KEYINPUT87), .ZN(new_n358));
  AOI211_X1 g172(.A(new_n358), .B(new_n344), .C1(new_n341), .C2(new_n343), .ZN(new_n359));
  OAI211_X1 g173(.A(new_n345), .B(new_n354), .C1(new_n357), .C2(new_n359), .ZN(new_n360));
  NAND3_X1  g174(.A1(new_n347), .A2(new_n349), .A3(KEYINPUT16), .ZN(new_n361));
  OR3_X1    g175(.A1(new_n348), .A2(KEYINPUT16), .A3(G140), .ZN(new_n362));
  NAND3_X1  g176(.A1(new_n361), .A2(new_n362), .A3(G146), .ZN(new_n363));
  INV_X1    g177(.A(KEYINPUT71), .ZN(new_n364));
  NAND2_X1  g178(.A1(new_n363), .A2(new_n364), .ZN(new_n365));
  AOI21_X1  g179(.A(G146), .B1(new_n361), .B2(new_n362), .ZN(new_n366));
  NOR2_X1   g180(.A1(new_n365), .A2(new_n366), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n361), .A2(new_n362), .ZN(new_n368));
  NAND3_X1  g182(.A1(new_n368), .A2(KEYINPUT71), .A3(new_n241), .ZN(new_n369));
  INV_X1    g183(.A(new_n369), .ZN(new_n370));
  INV_X1    g184(.A(KEYINPUT17), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n355), .A2(G131), .ZN(new_n372));
  OAI22_X1  g186(.A1(new_n367), .A2(new_n370), .B1(new_n371), .B2(new_n372), .ZN(new_n373));
  INV_X1    g187(.A(G131), .ZN(new_n374));
  NAND3_X1  g188(.A1(new_n341), .A2(new_n343), .A3(new_n374), .ZN(new_n375));
  INV_X1    g189(.A(KEYINPUT88), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n375), .A2(new_n376), .ZN(new_n377));
  NAND4_X1  g191(.A1(new_n341), .A2(new_n343), .A3(KEYINPUT88), .A4(new_n374), .ZN(new_n378));
  NAND3_X1  g192(.A1(new_n377), .A2(new_n378), .A3(new_n372), .ZN(new_n379));
  NOR2_X1   g193(.A1(new_n379), .A2(KEYINPUT17), .ZN(new_n380));
  OAI211_X1 g194(.A(new_n337), .B(new_n360), .C1(new_n373), .C2(new_n380), .ZN(new_n381));
  INV_X1    g195(.A(new_n337), .ZN(new_n382));
  XOR2_X1   g196(.A(KEYINPUT89), .B(KEYINPUT19), .Z(new_n383));
  NAND2_X1  g197(.A1(new_n383), .A2(new_n352), .ZN(new_n384));
  INV_X1    g198(.A(KEYINPUT89), .ZN(new_n385));
  OAI21_X1  g199(.A(new_n350), .B1(new_n385), .B2(KEYINPUT19), .ZN(new_n386));
  NAND3_X1  g200(.A1(new_n384), .A2(new_n386), .A3(new_n241), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n387), .A2(new_n363), .ZN(new_n388));
  AOI21_X1  g202(.A(new_n374), .B1(new_n341), .B2(new_n343), .ZN(new_n389));
  AOI21_X1  g203(.A(new_n389), .B1(new_n376), .B2(new_n375), .ZN(new_n390));
  AOI21_X1  g204(.A(new_n388), .B1(new_n390), .B2(new_n378), .ZN(new_n391));
  NAND2_X1  g205(.A1(new_n354), .A2(new_n345), .ZN(new_n392));
  INV_X1    g206(.A(new_n357), .ZN(new_n393));
  NAND3_X1  g207(.A1(new_n355), .A2(KEYINPUT87), .A3(new_n356), .ZN(new_n394));
  AOI21_X1  g208(.A(new_n392), .B1(new_n393), .B2(new_n394), .ZN(new_n395));
  OAI21_X1  g209(.A(new_n382), .B1(new_n391), .B2(new_n395), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n381), .A2(new_n396), .ZN(new_n397));
  NOR2_X1   g211(.A1(G475), .A2(G902), .ZN(new_n398));
  AOI21_X1  g212(.A(new_n335), .B1(new_n397), .B2(new_n398), .ZN(new_n399));
  INV_X1    g213(.A(new_n398), .ZN(new_n400));
  AOI211_X1 g214(.A(KEYINPUT20), .B(new_n400), .C1(new_n381), .C2(new_n396), .ZN(new_n401));
  OAI21_X1  g215(.A(new_n360), .B1(new_n373), .B2(new_n380), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n402), .A2(new_n382), .ZN(new_n403));
  AOI21_X1  g217(.A(G902), .B1(new_n403), .B2(new_n381), .ZN(new_n404));
  INV_X1    g218(.A(G475), .ZN(new_n405));
  OAI22_X1  g219(.A1(new_n399), .A2(new_n401), .B1(new_n404), .B2(new_n405), .ZN(new_n406));
  NOR2_X1   g220(.A1(new_n406), .A2(KEYINPUT90), .ZN(new_n407));
  INV_X1    g221(.A(KEYINPUT90), .ZN(new_n408));
  NAND3_X1  g222(.A1(new_n379), .A2(new_n363), .A3(new_n387), .ZN(new_n409));
  AOI21_X1  g223(.A(new_n337), .B1(new_n409), .B2(new_n360), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n368), .A2(new_n241), .ZN(new_n411));
  NAND3_X1  g225(.A1(new_n411), .A2(new_n364), .A3(new_n363), .ZN(new_n412));
  AOI22_X1  g226(.A1(new_n412), .A2(new_n369), .B1(KEYINPUT17), .B2(new_n389), .ZN(new_n413));
  NAND3_X1  g227(.A1(new_n390), .A2(new_n371), .A3(new_n378), .ZN(new_n414));
  AOI21_X1  g228(.A(new_n395), .B1(new_n413), .B2(new_n414), .ZN(new_n415));
  AOI21_X1  g229(.A(new_n410), .B1(new_n415), .B2(new_n337), .ZN(new_n416));
  OAI21_X1  g230(.A(KEYINPUT20), .B1(new_n416), .B2(new_n400), .ZN(new_n417));
  NAND3_X1  g231(.A1(new_n397), .A2(new_n335), .A3(new_n398), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n417), .A2(new_n418), .ZN(new_n419));
  NOR2_X1   g233(.A1(new_n415), .A2(new_n337), .ZN(new_n420));
  INV_X1    g234(.A(new_n381), .ZN(new_n421));
  OAI21_X1  g235(.A(new_n190), .B1(new_n420), .B2(new_n421), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n422), .A2(G475), .ZN(new_n423));
  AOI21_X1  g237(.A(new_n408), .B1(new_n419), .B2(new_n423), .ZN(new_n424));
  OAI21_X1  g238(.A(new_n334), .B1(new_n407), .B2(new_n424), .ZN(new_n425));
  NOR2_X1   g239(.A1(new_n295), .A2(new_n425), .ZN(new_n426));
  XNOR2_X1  g240(.A(G110), .B(G140), .ZN(new_n427));
  AND2_X1   g241(.A1(new_n285), .A2(G227), .ZN(new_n428));
  XNOR2_X1  g242(.A(new_n427), .B(new_n428), .ZN(new_n429));
  INV_X1    g243(.A(KEYINPUT78), .ZN(new_n430));
  AND3_X1   g244(.A1(new_n199), .A2(new_n207), .A3(G101), .ZN(new_n431));
  AOI21_X1  g245(.A(new_n207), .B1(new_n199), .B2(G101), .ZN(new_n432));
  AOI21_X1  g246(.A(new_n431), .B1(new_n205), .B2(new_n432), .ZN(new_n433));
  OAI21_X1  g247(.A(new_n430), .B1(new_n433), .B2(new_n256), .ZN(new_n434));
  AOI21_X1  g248(.A(new_n256), .B1(new_n206), .B2(new_n208), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n435), .A2(KEYINPUT78), .ZN(new_n436));
  NAND2_X1  g250(.A1(new_n433), .A2(new_n256), .ZN(new_n437));
  NAND3_X1  g251(.A1(new_n434), .A2(new_n436), .A3(new_n437), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n305), .A2(G137), .ZN(new_n439));
  INV_X1    g253(.A(G137), .ZN(new_n440));
  AOI21_X1  g254(.A(KEYINPUT64), .B1(new_n440), .B2(G134), .ZN(new_n441));
  INV_X1    g255(.A(KEYINPUT11), .ZN(new_n442));
  OAI21_X1  g256(.A(new_n439), .B1(new_n441), .B2(new_n442), .ZN(new_n443));
  AOI211_X1 g257(.A(KEYINPUT64), .B(KEYINPUT11), .C1(new_n440), .C2(G134), .ZN(new_n444));
  NOR3_X1   g258(.A1(new_n443), .A2(G131), .A3(new_n444), .ZN(new_n445));
  NOR2_X1   g259(.A1(new_n440), .A2(G134), .ZN(new_n446));
  INV_X1    g260(.A(KEYINPUT64), .ZN(new_n447));
  OAI21_X1  g261(.A(new_n447), .B1(new_n305), .B2(G137), .ZN(new_n448));
  AOI21_X1  g262(.A(new_n446), .B1(new_n448), .B2(KEYINPUT11), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n441), .A2(new_n442), .ZN(new_n450));
  AOI21_X1  g264(.A(new_n374), .B1(new_n449), .B2(new_n450), .ZN(new_n451));
  NOR2_X1   g265(.A1(new_n445), .A2(new_n451), .ZN(new_n452));
  INV_X1    g266(.A(new_n452), .ZN(new_n453));
  AND3_X1   g267(.A1(new_n438), .A2(KEYINPUT12), .A3(new_n453), .ZN(new_n454));
  AOI21_X1  g268(.A(KEYINPUT12), .B1(new_n438), .B2(new_n453), .ZN(new_n455));
  NOR2_X1   g269(.A1(new_n454), .A2(new_n455), .ZN(new_n456));
  INV_X1    g270(.A(KEYINPUT10), .ZN(new_n457));
  NAND3_X1  g271(.A1(new_n434), .A2(new_n457), .A3(new_n436), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n435), .A2(KEYINPUT10), .ZN(new_n459));
  INV_X1    g273(.A(new_n248), .ZN(new_n460));
  OAI211_X1 g274(.A(new_n234), .B(new_n460), .C1(KEYINPUT4), .C2(new_n233), .ZN(new_n461));
  AND2_X1   g275(.A1(new_n459), .A2(new_n461), .ZN(new_n462));
  NAND3_X1  g276(.A1(new_n458), .A2(new_n462), .A3(new_n452), .ZN(new_n463));
  INV_X1    g277(.A(new_n463), .ZN(new_n464));
  OAI21_X1  g278(.A(new_n429), .B1(new_n456), .B2(new_n464), .ZN(new_n465));
  INV_X1    g279(.A(KEYINPUT80), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n458), .A2(new_n462), .ZN(new_n467));
  AOI21_X1  g281(.A(new_n466), .B1(new_n467), .B2(new_n453), .ZN(new_n468));
  AOI211_X1 g282(.A(KEYINPUT80), .B(new_n452), .C1(new_n458), .C2(new_n462), .ZN(new_n469));
  INV_X1    g283(.A(new_n429), .ZN(new_n470));
  NAND2_X1  g284(.A1(new_n463), .A2(new_n470), .ZN(new_n471));
  OAI22_X1  g285(.A1(new_n468), .A2(new_n469), .B1(new_n471), .B2(KEYINPUT79), .ZN(new_n472));
  AND2_X1   g286(.A1(new_n471), .A2(KEYINPUT79), .ZN(new_n473));
  OAI21_X1  g287(.A(new_n465), .B1(new_n472), .B2(new_n473), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n474), .A2(KEYINPUT81), .ZN(new_n475));
  INV_X1    g289(.A(KEYINPUT81), .ZN(new_n476));
  OAI211_X1 g290(.A(new_n465), .B(new_n476), .C1(new_n472), .C2(new_n473), .ZN(new_n477));
  AND3_X1   g291(.A1(new_n475), .A2(G469), .A3(new_n477), .ZN(new_n478));
  INV_X1    g292(.A(G469), .ZN(new_n479));
  OAI21_X1  g293(.A(KEYINPUT82), .B1(new_n456), .B2(new_n471), .ZN(new_n480));
  NAND2_X1  g294(.A1(new_n459), .A2(new_n461), .ZN(new_n481));
  AOI21_X1  g295(.A(KEYINPUT78), .B1(new_n209), .B2(new_n257), .ZN(new_n482));
  AOI211_X1 g296(.A(new_n430), .B(new_n256), .C1(new_n206), .C2(new_n208), .ZN(new_n483));
  NOR2_X1   g297(.A1(new_n482), .A2(new_n483), .ZN(new_n484));
  AOI21_X1  g298(.A(new_n481), .B1(new_n484), .B2(new_n457), .ZN(new_n485));
  AOI21_X1  g299(.A(new_n429), .B1(new_n485), .B2(new_n452), .ZN(new_n486));
  INV_X1    g300(.A(KEYINPUT82), .ZN(new_n487));
  OAI211_X1 g301(.A(new_n486), .B(new_n487), .C1(new_n454), .C2(new_n455), .ZN(new_n488));
  NAND2_X1  g302(.A1(new_n480), .A2(new_n488), .ZN(new_n489));
  OAI21_X1  g303(.A(KEYINPUT80), .B1(new_n485), .B2(new_n452), .ZN(new_n490));
  NAND3_X1  g304(.A1(new_n467), .A2(new_n466), .A3(new_n453), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  AOI21_X1  g306(.A(new_n470), .B1(new_n492), .B2(new_n463), .ZN(new_n493));
  OAI211_X1 g307(.A(new_n479), .B(new_n190), .C1(new_n489), .C2(new_n493), .ZN(new_n494));
  NOR2_X1   g308(.A1(new_n479), .A2(new_n190), .ZN(new_n495));
  INV_X1    g309(.A(new_n495), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n494), .A2(new_n496), .ZN(new_n497));
  OAI211_X1 g311(.A(new_n192), .B(new_n426), .C1(new_n478), .C2(new_n497), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n254), .A2(G119), .ZN(new_n499));
  NAND2_X1  g313(.A1(new_n210), .A2(G128), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  XNOR2_X1  g315(.A(KEYINPUT24), .B(G110), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  INV_X1    g317(.A(KEYINPUT23), .ZN(new_n504));
  OAI21_X1  g318(.A(new_n504), .B1(new_n210), .B2(G128), .ZN(new_n505));
  NAND3_X1  g319(.A1(new_n254), .A2(KEYINPUT23), .A3(G119), .ZN(new_n506));
  NAND3_X1  g320(.A1(new_n505), .A2(new_n500), .A3(new_n506), .ZN(new_n507));
  OAI21_X1  g321(.A(new_n503), .B1(G110), .B2(new_n507), .ZN(new_n508));
  NAND3_X1  g322(.A1(new_n508), .A2(new_n363), .A3(new_n353), .ZN(new_n509));
  INV_X1    g323(.A(new_n509), .ZN(new_n510));
  NOR2_X1   g324(.A1(new_n501), .A2(new_n502), .ZN(new_n511));
  INV_X1    g325(.A(G110), .ZN(new_n512));
  INV_X1    g326(.A(KEYINPUT70), .ZN(new_n513));
  AOI21_X1  g327(.A(new_n512), .B1(new_n507), .B2(new_n513), .ZN(new_n514));
  NAND4_X1  g328(.A1(new_n505), .A2(new_n506), .A3(KEYINPUT70), .A4(new_n500), .ZN(new_n515));
  AOI21_X1  g329(.A(new_n511), .B1(new_n514), .B2(new_n515), .ZN(new_n516));
  NAND3_X1  g330(.A1(new_n516), .A2(new_n412), .A3(new_n369), .ZN(new_n517));
  INV_X1    g331(.A(KEYINPUT72), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  NAND4_X1  g333(.A1(new_n516), .A2(new_n412), .A3(KEYINPUT72), .A4(new_n369), .ZN(new_n520));
  AOI21_X1  g334(.A(new_n510), .B1(new_n519), .B2(new_n520), .ZN(new_n521));
  XNOR2_X1  g335(.A(KEYINPUT22), .B(G137), .ZN(new_n522));
  AND3_X1   g336(.A1(new_n285), .A2(G221), .A3(G234), .ZN(new_n523));
  XOR2_X1   g337(.A(new_n522), .B(new_n523), .Z(new_n524));
  AOI21_X1  g338(.A(G902), .B1(new_n521), .B2(new_n524), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n519), .A2(new_n520), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n526), .A2(new_n509), .ZN(new_n527));
  INV_X1    g341(.A(new_n524), .ZN(new_n528));
  AOI21_X1  g342(.A(KEYINPUT73), .B1(new_n527), .B2(new_n528), .ZN(new_n529));
  INV_X1    g343(.A(KEYINPUT73), .ZN(new_n530));
  NOR3_X1   g344(.A1(new_n521), .A2(new_n530), .A3(new_n524), .ZN(new_n531));
  OAI21_X1  g345(.A(new_n525), .B1(new_n529), .B2(new_n531), .ZN(new_n532));
  NOR2_X1   g346(.A1(KEYINPUT74), .A2(KEYINPUT25), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  INV_X1    g348(.A(new_n533), .ZN(new_n535));
  OAI211_X1 g349(.A(new_n525), .B(new_n535), .C1(new_n529), .C2(new_n531), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n534), .A2(new_n536), .ZN(new_n537));
  AOI21_X1  g351(.A(new_n323), .B1(G234), .B2(new_n190), .ZN(new_n538));
  AOI21_X1  g352(.A(KEYINPUT75), .B1(new_n537), .B2(new_n538), .ZN(new_n539));
  INV_X1    g353(.A(KEYINPUT75), .ZN(new_n540));
  INV_X1    g354(.A(new_n538), .ZN(new_n541));
  AOI211_X1 g355(.A(new_n540), .B(new_n541), .C1(new_n534), .C2(new_n536), .ZN(new_n542));
  NOR2_X1   g356(.A1(new_n539), .A2(new_n542), .ZN(new_n543));
  XNOR2_X1  g357(.A(KEYINPUT68), .B(KEYINPUT32), .ZN(new_n544));
  NAND2_X1  g358(.A1(new_n342), .A2(G210), .ZN(new_n545));
  XNOR2_X1  g359(.A(new_n545), .B(KEYINPUT27), .ZN(new_n546));
  XNOR2_X1  g360(.A(KEYINPUT26), .B(G101), .ZN(new_n547));
  XNOR2_X1  g361(.A(new_n546), .B(new_n547), .ZN(new_n548));
  XNOR2_X1  g362(.A(new_n548), .B(KEYINPUT65), .ZN(new_n549));
  INV_X1    g363(.A(KEYINPUT28), .ZN(new_n550));
  NAND2_X1  g364(.A1(new_n225), .A2(new_n230), .ZN(new_n551));
  OAI21_X1  g365(.A(G131), .B1(new_n443), .B2(new_n444), .ZN(new_n552));
  NAND3_X1  g366(.A1(new_n449), .A2(new_n374), .A3(new_n450), .ZN(new_n553));
  AOI21_X1  g367(.A(new_n248), .B1(new_n552), .B2(new_n553), .ZN(new_n554));
  NOR2_X1   g368(.A1(new_n305), .A2(G137), .ZN(new_n555));
  OAI21_X1  g369(.A(G131), .B1(new_n555), .B2(new_n446), .ZN(new_n556));
  NAND3_X1  g370(.A1(new_n253), .A2(new_n255), .A3(new_n556), .ZN(new_n557));
  NOR2_X1   g371(.A1(new_n445), .A2(new_n557), .ZN(new_n558));
  OAI21_X1  g372(.A(new_n551), .B1(new_n554), .B2(new_n558), .ZN(new_n559));
  OAI21_X1  g373(.A(new_n460), .B1(new_n445), .B2(new_n451), .ZN(new_n560));
  INV_X1    g374(.A(new_n551), .ZN(new_n561));
  NAND4_X1  g375(.A1(new_n553), .A2(new_n255), .A3(new_n253), .A4(new_n556), .ZN(new_n562));
  NAND3_X1  g376(.A1(new_n560), .A2(new_n561), .A3(new_n562), .ZN(new_n563));
  AOI21_X1  g377(.A(new_n550), .B1(new_n559), .B2(new_n563), .ZN(new_n564));
  INV_X1    g378(.A(KEYINPUT66), .ZN(new_n565));
  AOI21_X1  g379(.A(new_n565), .B1(new_n563), .B2(new_n550), .ZN(new_n566));
  NOR2_X1   g380(.A1(new_n564), .A2(new_n566), .ZN(new_n567));
  AOI211_X1 g381(.A(new_n565), .B(new_n550), .C1(new_n559), .C2(new_n563), .ZN(new_n568));
  OAI21_X1  g382(.A(new_n549), .B1(new_n567), .B2(new_n568), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n569), .A2(KEYINPUT67), .ZN(new_n570));
  NOR3_X1   g384(.A1(new_n554), .A2(new_n558), .A3(KEYINPUT30), .ZN(new_n571));
  INV_X1    g385(.A(KEYINPUT30), .ZN(new_n572));
  AOI21_X1  g386(.A(new_n572), .B1(new_n560), .B2(new_n562), .ZN(new_n573));
  OAI21_X1  g387(.A(new_n551), .B1(new_n571), .B2(new_n573), .ZN(new_n574));
  NAND3_X1  g388(.A1(new_n574), .A2(new_n548), .A3(new_n563), .ZN(new_n575));
  INV_X1    g389(.A(KEYINPUT31), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n575), .A2(new_n576), .ZN(new_n577));
  INV_X1    g391(.A(new_n563), .ZN(new_n578));
  OAI21_X1  g392(.A(KEYINPUT30), .B1(new_n554), .B2(new_n558), .ZN(new_n579));
  NAND3_X1  g393(.A1(new_n560), .A2(new_n572), .A3(new_n562), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  AOI21_X1  g395(.A(new_n578), .B1(new_n581), .B2(new_n551), .ZN(new_n582));
  NAND3_X1  g396(.A1(new_n582), .A2(KEYINPUT31), .A3(new_n548), .ZN(new_n583));
  NAND2_X1  g397(.A1(new_n577), .A2(new_n583), .ZN(new_n584));
  INV_X1    g398(.A(KEYINPUT67), .ZN(new_n585));
  OAI211_X1 g399(.A(new_n585), .B(new_n549), .C1(new_n567), .C2(new_n568), .ZN(new_n586));
  NAND3_X1  g400(.A1(new_n570), .A2(new_n584), .A3(new_n586), .ZN(new_n587));
  NOR2_X1   g401(.A1(G472), .A2(G902), .ZN(new_n588));
  AOI21_X1  g402(.A(new_n544), .B1(new_n587), .B2(new_n588), .ZN(new_n589));
  INV_X1    g403(.A(new_n589), .ZN(new_n590));
  NAND3_X1  g404(.A1(new_n587), .A2(KEYINPUT32), .A3(new_n588), .ZN(new_n591));
  INV_X1    g405(.A(KEYINPUT69), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n564), .A2(new_n592), .ZN(new_n593));
  OAI21_X1  g407(.A(KEYINPUT69), .B1(new_n578), .B2(KEYINPUT28), .ZN(new_n594));
  OAI21_X1  g408(.A(new_n593), .B1(new_n564), .B2(new_n594), .ZN(new_n595));
  INV_X1    g409(.A(new_n548), .ZN(new_n596));
  INV_X1    g410(.A(KEYINPUT29), .ZN(new_n597));
  NOR2_X1   g411(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n595), .A2(new_n598), .ZN(new_n599));
  NOR3_X1   g413(.A1(new_n567), .A2(new_n568), .A3(new_n549), .ZN(new_n600));
  OAI21_X1  g414(.A(new_n597), .B1(new_n582), .B2(new_n548), .ZN(new_n601));
  OAI211_X1 g415(.A(new_n599), .B(new_n190), .C1(new_n600), .C2(new_n601), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n602), .A2(G472), .ZN(new_n603));
  NAND3_X1  g417(.A1(new_n590), .A2(new_n591), .A3(new_n603), .ZN(new_n604));
  NAND3_X1  g418(.A1(new_n527), .A2(KEYINPUT73), .A3(new_n528), .ZN(new_n605));
  OAI21_X1  g419(.A(new_n530), .B1(new_n521), .B2(new_n524), .ZN(new_n606));
  AOI22_X1  g420(.A1(new_n605), .A2(new_n606), .B1(new_n521), .B2(new_n524), .ZN(new_n607));
  NOR2_X1   g421(.A1(new_n538), .A2(G902), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  NAND3_X1  g423(.A1(new_n543), .A2(new_n604), .A3(new_n609), .ZN(new_n610));
  NOR2_X1   g424(.A1(new_n498), .A2(new_n610), .ZN(new_n611));
  XNOR2_X1  g425(.A(new_n611), .B(new_n201), .ZN(G3));
  OAI21_X1  g426(.A(new_n192), .B1(new_n478), .B2(new_n497), .ZN(new_n613));
  NAND2_X1  g427(.A1(new_n406), .A2(KEYINPUT90), .ZN(new_n614));
  NAND3_X1  g428(.A1(new_n419), .A2(new_n408), .A3(new_n423), .ZN(new_n615));
  NAND2_X1  g429(.A1(new_n326), .A2(new_n327), .ZN(new_n616));
  NAND2_X1  g430(.A1(new_n616), .A2(KEYINPUT33), .ZN(new_n617));
  INV_X1    g431(.A(KEYINPUT33), .ZN(new_n618));
  NAND3_X1  g432(.A1(new_n326), .A2(new_n618), .A3(new_n327), .ZN(new_n619));
  NAND3_X1  g433(.A1(new_n617), .A2(G478), .A3(new_n619), .ZN(new_n620));
  NOR2_X1   g434(.A1(new_n330), .A2(new_n190), .ZN(new_n621));
  AOI21_X1  g435(.A(new_n621), .B1(new_n328), .B2(new_n330), .ZN(new_n622));
  AND2_X1   g436(.A1(new_n620), .A2(new_n622), .ZN(new_n623));
  NAND3_X1  g437(.A1(new_n614), .A2(new_n615), .A3(new_n623), .ZN(new_n624));
  NAND2_X1  g438(.A1(new_n587), .A2(new_n190), .ZN(new_n625));
  AOI22_X1  g439(.A1(new_n625), .A2(G472), .B1(new_n588), .B2(new_n587), .ZN(new_n626));
  INV_X1    g440(.A(new_n536), .ZN(new_n627));
  NAND2_X1  g441(.A1(new_n605), .A2(new_n606), .ZN(new_n628));
  AOI21_X1  g442(.A(new_n535), .B1(new_n628), .B2(new_n525), .ZN(new_n629));
  OAI21_X1  g443(.A(new_n538), .B1(new_n627), .B2(new_n629), .ZN(new_n630));
  NAND2_X1  g444(.A1(new_n630), .A2(new_n540), .ZN(new_n631));
  NAND3_X1  g445(.A1(new_n537), .A2(KEYINPUT75), .A3(new_n538), .ZN(new_n632));
  NAND4_X1  g446(.A1(new_n626), .A2(new_n631), .A3(new_n632), .A4(new_n609), .ZN(new_n633));
  NOR3_X1   g447(.A1(new_n613), .A2(new_n624), .A3(new_n633), .ZN(new_n634));
  INV_X1    g448(.A(new_n291), .ZN(new_n635));
  NAND2_X1  g449(.A1(new_n279), .A2(new_n280), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n636), .A2(new_n292), .ZN(new_n637));
  INV_X1    g451(.A(new_n637), .ZN(new_n638));
  NAND3_X1  g452(.A1(new_n634), .A2(new_n635), .A3(new_n638), .ZN(new_n639));
  XOR2_X1   g453(.A(KEYINPUT34), .B(G104), .Z(new_n640));
  XNOR2_X1  g454(.A(new_n639), .B(new_n640), .ZN(new_n641));
  XNOR2_X1  g455(.A(KEYINPUT94), .B(KEYINPUT95), .ZN(new_n642));
  XNOR2_X1  g456(.A(new_n641), .B(new_n642), .ZN(G6));
  AND2_X1   g457(.A1(new_n494), .A2(new_n496), .ZN(new_n644));
  NAND3_X1  g458(.A1(new_n475), .A2(G469), .A3(new_n477), .ZN(new_n645));
  AOI21_X1  g459(.A(new_n191), .B1(new_n644), .B2(new_n645), .ZN(new_n646));
  INV_X1    g460(.A(new_n633), .ZN(new_n647));
  NAND3_X1  g461(.A1(new_n636), .A2(new_n635), .A3(new_n292), .ZN(new_n648));
  INV_X1    g462(.A(new_n406), .ZN(new_n649));
  NAND2_X1  g463(.A1(new_n332), .A2(new_n333), .ZN(new_n650));
  NAND2_X1  g464(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  NOR2_X1   g465(.A1(new_n648), .A2(new_n651), .ZN(new_n652));
  NAND3_X1  g466(.A1(new_n646), .A2(new_n647), .A3(new_n652), .ZN(new_n653));
  XOR2_X1   g467(.A(KEYINPUT35), .B(G107), .Z(new_n654));
  XNOR2_X1  g468(.A(new_n653), .B(new_n654), .ZN(G9));
  NOR2_X1   g469(.A1(new_n528), .A2(KEYINPUT36), .ZN(new_n656));
  XNOR2_X1  g470(.A(new_n527), .B(new_n656), .ZN(new_n657));
  NAND2_X1  g471(.A1(new_n657), .A2(new_n608), .ZN(new_n658));
  NAND3_X1  g472(.A1(new_n631), .A2(new_n632), .A3(new_n658), .ZN(new_n659));
  NAND2_X1  g473(.A1(new_n659), .A2(new_n626), .ZN(new_n660));
  NOR2_X1   g474(.A1(new_n498), .A2(new_n660), .ZN(new_n661));
  XNOR2_X1  g475(.A(KEYINPUT37), .B(G110), .ZN(new_n662));
  XNOR2_X1  g476(.A(new_n661), .B(new_n662), .ZN(G12));
  AND2_X1   g477(.A1(new_n591), .A2(new_n603), .ZN(new_n664));
  AOI21_X1  g478(.A(new_n637), .B1(new_n664), .B2(new_n590), .ZN(new_n665));
  XOR2_X1   g479(.A(new_n286), .B(KEYINPUT96), .Z(new_n666));
  INV_X1    g480(.A(new_n666), .ZN(new_n667));
  INV_X1    g481(.A(G900), .ZN(new_n668));
  AOI21_X1  g482(.A(new_n667), .B1(new_n668), .B2(new_n289), .ZN(new_n669));
  NOR2_X1   g483(.A1(new_n651), .A2(new_n669), .ZN(new_n670));
  NAND4_X1  g484(.A1(new_n646), .A2(new_n659), .A3(new_n665), .A4(new_n670), .ZN(new_n671));
  XNOR2_X1  g485(.A(new_n671), .B(G128), .ZN(G30));
  XOR2_X1   g486(.A(new_n669), .B(KEYINPUT39), .Z(new_n673));
  NAND2_X1  g487(.A1(new_n646), .A2(new_n673), .ZN(new_n674));
  AND2_X1   g488(.A1(new_n674), .A2(KEYINPUT40), .ZN(new_n675));
  NOR2_X1   g489(.A1(new_n674), .A2(KEYINPUT40), .ZN(new_n676));
  NAND2_X1  g490(.A1(new_n559), .A2(new_n563), .ZN(new_n677));
  AOI22_X1  g491(.A1(new_n582), .A2(new_n548), .B1(new_n677), .B2(new_n549), .ZN(new_n678));
  OAI21_X1  g492(.A(G472), .B1(new_n678), .B2(G902), .ZN(new_n679));
  NAND2_X1  g493(.A1(new_n591), .A2(new_n679), .ZN(new_n680));
  NOR2_X1   g494(.A1(new_n680), .A2(new_n589), .ZN(new_n681));
  NOR2_X1   g495(.A1(new_n659), .A2(new_n681), .ZN(new_n682));
  AND3_X1   g496(.A1(new_n267), .A2(new_n275), .A3(new_n277), .ZN(new_n683));
  AOI21_X1  g497(.A(new_n277), .B1(new_n267), .B2(new_n275), .ZN(new_n684));
  NOR2_X1   g498(.A1(new_n683), .A2(new_n684), .ZN(new_n685));
  AOI21_X1  g499(.A(new_n282), .B1(new_n685), .B2(KEYINPUT85), .ZN(new_n686));
  XNOR2_X1  g500(.A(new_n686), .B(KEYINPUT38), .ZN(new_n687));
  AOI21_X1  g501(.A(new_n293), .B1(new_n332), .B2(new_n333), .ZN(new_n688));
  NAND3_X1  g502(.A1(new_n614), .A2(new_n688), .A3(new_n615), .ZN(new_n689));
  INV_X1    g503(.A(new_n689), .ZN(new_n690));
  NAND3_X1  g504(.A1(new_n682), .A2(new_n687), .A3(new_n690), .ZN(new_n691));
  NOR3_X1   g505(.A1(new_n675), .A2(new_n676), .A3(new_n691), .ZN(new_n692));
  XNOR2_X1  g506(.A(new_n692), .B(new_n243), .ZN(G45));
  INV_X1    g507(.A(new_n624), .ZN(new_n694));
  INV_X1    g508(.A(new_n669), .ZN(new_n695));
  NAND2_X1  g509(.A1(new_n694), .A2(new_n695), .ZN(new_n696));
  AOI21_X1  g510(.A(new_n696), .B1(new_n543), .B2(new_n658), .ZN(new_n697));
  NAND3_X1  g511(.A1(new_n646), .A2(new_n697), .A3(new_n665), .ZN(new_n698));
  XNOR2_X1  g512(.A(new_n698), .B(G146), .ZN(G48));
  NOR2_X1   g513(.A1(new_n648), .A2(new_n624), .ZN(new_n700));
  NAND4_X1  g514(.A1(new_n543), .A2(new_n604), .A3(new_n609), .A4(new_n700), .ZN(new_n701));
  AOI21_X1  g515(.A(new_n464), .B1(new_n490), .B2(new_n491), .ZN(new_n702));
  OAI211_X1 g516(.A(new_n480), .B(new_n488), .C1(new_n470), .C2(new_n702), .ZN(new_n703));
  NAND2_X1  g517(.A1(new_n703), .A2(new_n190), .ZN(new_n704));
  NAND2_X1  g518(.A1(new_n704), .A2(G469), .ZN(new_n705));
  NAND3_X1  g519(.A1(new_n705), .A2(new_n192), .A3(new_n494), .ZN(new_n706));
  NOR2_X1   g520(.A1(new_n701), .A2(new_n706), .ZN(new_n707));
  XOR2_X1   g521(.A(KEYINPUT41), .B(G113), .Z(new_n708));
  XNOR2_X1  g522(.A(new_n707), .B(new_n708), .ZN(G15));
  NAND4_X1  g523(.A1(new_n543), .A2(new_n604), .A3(new_n609), .A4(new_n652), .ZN(new_n710));
  NOR2_X1   g524(.A1(new_n710), .A2(new_n706), .ZN(new_n711));
  XNOR2_X1  g525(.A(new_n711), .B(new_n226), .ZN(G18));
  INV_X1    g526(.A(new_n494), .ZN(new_n713));
  AOI21_X1  g527(.A(new_n479), .B1(new_n703), .B2(new_n190), .ZN(new_n714));
  NOR3_X1   g528(.A1(new_n713), .A2(new_n714), .A3(new_n191), .ZN(new_n715));
  NOR2_X1   g529(.A1(new_n425), .A2(new_n291), .ZN(new_n716));
  NAND4_X1  g530(.A1(new_n715), .A2(new_n659), .A3(new_n665), .A4(new_n716), .ZN(new_n717));
  XNOR2_X1  g531(.A(new_n717), .B(G119), .ZN(G21));
  OAI211_X1 g532(.A(new_n593), .B(new_n549), .C1(new_n564), .C2(new_n594), .ZN(new_n719));
  NAND2_X1  g533(.A1(new_n584), .A2(new_n719), .ZN(new_n720));
  AOI22_X1  g534(.A1(new_n625), .A2(G472), .B1(new_n588), .B2(new_n720), .ZN(new_n721));
  NAND4_X1  g535(.A1(new_n721), .A2(new_n631), .A3(new_n632), .A4(new_n609), .ZN(new_n722));
  INV_X1    g536(.A(new_n722), .ZN(new_n723));
  NOR3_X1   g537(.A1(new_n689), .A2(new_n685), .A3(new_n291), .ZN(new_n724));
  NAND3_X1  g538(.A1(new_n723), .A2(new_n715), .A3(new_n724), .ZN(new_n725));
  XNOR2_X1  g539(.A(new_n725), .B(G122), .ZN(G24));
  NOR2_X1   g540(.A1(new_n624), .A2(new_n669), .ZN(new_n727));
  AND3_X1   g541(.A1(new_n659), .A2(new_n727), .A3(new_n721), .ZN(new_n728));
  NOR4_X1   g542(.A1(new_n713), .A2(new_n714), .A3(new_n191), .A4(new_n637), .ZN(new_n729));
  NAND2_X1  g543(.A1(new_n728), .A2(new_n729), .ZN(new_n730));
  XNOR2_X1  g544(.A(new_n730), .B(G125), .ZN(G27));
  OAI21_X1  g545(.A(KEYINPUT97), .B1(new_n686), .B2(new_n293), .ZN(new_n732));
  OAI211_X1 g546(.A(new_n465), .B(G469), .C1(new_n472), .C2(new_n473), .ZN(new_n733));
  NAND3_X1  g547(.A1(new_n494), .A2(new_n496), .A3(new_n733), .ZN(new_n734));
  NAND2_X1  g548(.A1(new_n281), .A2(new_n283), .ZN(new_n735));
  INV_X1    g549(.A(KEYINPUT97), .ZN(new_n736));
  NAND3_X1  g550(.A1(new_n735), .A2(new_n736), .A3(new_n292), .ZN(new_n737));
  NAND4_X1  g551(.A1(new_n732), .A2(new_n192), .A3(new_n734), .A4(new_n737), .ZN(new_n738));
  NOR2_X1   g552(.A1(new_n738), .A2(new_n696), .ZN(new_n739));
  NAND3_X1  g553(.A1(new_n631), .A2(new_n632), .A3(new_n609), .ZN(new_n740));
  NAND2_X1  g554(.A1(new_n591), .A2(new_n603), .ZN(new_n741));
  AOI21_X1  g555(.A(KEYINPUT32), .B1(new_n587), .B2(new_n588), .ZN(new_n742));
  NOR2_X1   g556(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  NOR2_X1   g557(.A1(new_n740), .A2(new_n743), .ZN(new_n744));
  NAND3_X1  g558(.A1(new_n739), .A2(KEYINPUT42), .A3(new_n744), .ZN(new_n745));
  INV_X1    g559(.A(new_n745), .ZN(new_n746));
  XOR2_X1   g560(.A(KEYINPUT99), .B(KEYINPUT42), .Z(new_n747));
  NOR3_X1   g561(.A1(new_n738), .A2(new_n610), .A3(new_n696), .ZN(new_n748));
  AOI21_X1  g562(.A(new_n747), .B1(new_n748), .B2(KEYINPUT98), .ZN(new_n749));
  INV_X1    g563(.A(new_n738), .ZN(new_n750));
  NOR2_X1   g564(.A1(new_n741), .A2(new_n589), .ZN(new_n751));
  NOR2_X1   g565(.A1(new_n740), .A2(new_n751), .ZN(new_n752));
  NAND3_X1  g566(.A1(new_n750), .A2(new_n752), .A3(new_n727), .ZN(new_n753));
  INV_X1    g567(.A(KEYINPUT98), .ZN(new_n754));
  NAND2_X1  g568(.A1(new_n753), .A2(new_n754), .ZN(new_n755));
  AOI21_X1  g569(.A(new_n746), .B1(new_n749), .B2(new_n755), .ZN(new_n756));
  XNOR2_X1  g570(.A(new_n756), .B(new_n374), .ZN(G33));
  NAND4_X1  g571(.A1(new_n543), .A2(new_n604), .A3(new_n609), .A4(new_n670), .ZN(new_n758));
  NOR2_X1   g572(.A1(new_n738), .A2(new_n758), .ZN(new_n759));
  XOR2_X1   g573(.A(KEYINPUT100), .B(G134), .Z(new_n760));
  XNOR2_X1  g574(.A(new_n759), .B(new_n760), .ZN(G36));
  NAND2_X1  g575(.A1(new_n475), .A2(new_n477), .ZN(new_n762));
  INV_X1    g576(.A(KEYINPUT45), .ZN(new_n763));
  NAND2_X1  g577(.A1(new_n762), .A2(new_n763), .ZN(new_n764));
  OAI211_X1 g578(.A(new_n764), .B(G469), .C1(new_n763), .C2(new_n474), .ZN(new_n765));
  XNOR2_X1  g579(.A(new_n765), .B(KEYINPUT101), .ZN(new_n766));
  NAND2_X1  g580(.A1(new_n766), .A2(new_n496), .ZN(new_n767));
  INV_X1    g581(.A(KEYINPUT46), .ZN(new_n768));
  OAI21_X1  g582(.A(new_n494), .B1(new_n767), .B2(new_n768), .ZN(new_n769));
  INV_X1    g583(.A(KEYINPUT102), .ZN(new_n770));
  AND2_X1   g584(.A1(new_n769), .A2(new_n770), .ZN(new_n771));
  NAND2_X1  g585(.A1(new_n767), .A2(new_n768), .ZN(new_n772));
  OAI21_X1  g586(.A(new_n772), .B1(new_n769), .B2(new_n770), .ZN(new_n773));
  NOR2_X1   g587(.A1(new_n771), .A2(new_n773), .ZN(new_n774));
  NOR2_X1   g588(.A1(new_n774), .A2(new_n191), .ZN(new_n775));
  NAND2_X1  g589(.A1(new_n732), .A2(new_n737), .ZN(new_n776));
  NOR2_X1   g590(.A1(new_n407), .A2(new_n424), .ZN(new_n777));
  INV_X1    g591(.A(new_n777), .ZN(new_n778));
  NAND2_X1  g592(.A1(new_n778), .A2(new_n623), .ZN(new_n779));
  XOR2_X1   g593(.A(new_n779), .B(KEYINPUT43), .Z(new_n780));
  INV_X1    g594(.A(new_n626), .ZN(new_n781));
  NAND3_X1  g595(.A1(new_n780), .A2(new_n781), .A3(new_n659), .ZN(new_n782));
  INV_X1    g596(.A(KEYINPUT44), .ZN(new_n783));
  AOI21_X1  g597(.A(new_n776), .B1(new_n782), .B2(new_n783), .ZN(new_n784));
  OAI21_X1  g598(.A(new_n784), .B1(new_n783), .B2(new_n782), .ZN(new_n785));
  INV_X1    g599(.A(new_n785), .ZN(new_n786));
  NAND3_X1  g600(.A1(new_n775), .A2(new_n673), .A3(new_n786), .ZN(new_n787));
  XNOR2_X1  g601(.A(new_n787), .B(G137), .ZN(G39));
  INV_X1    g602(.A(KEYINPUT47), .ZN(new_n789));
  OAI21_X1  g603(.A(new_n789), .B1(new_n774), .B2(new_n191), .ZN(new_n790));
  OAI211_X1 g604(.A(KEYINPUT47), .B(new_n192), .C1(new_n771), .C2(new_n773), .ZN(new_n791));
  AND2_X1   g605(.A1(new_n790), .A2(new_n791), .ZN(new_n792));
  INV_X1    g606(.A(new_n776), .ZN(new_n793));
  NAND4_X1  g607(.A1(new_n793), .A2(new_n751), .A3(new_n740), .A4(new_n727), .ZN(new_n794));
  NOR2_X1   g608(.A1(new_n792), .A2(new_n794), .ZN(new_n795));
  XNOR2_X1  g609(.A(new_n795), .B(new_n346), .ZN(G42));
  NOR4_X1   g610(.A1(new_n687), .A2(new_n191), .A3(new_n293), .A4(new_n779), .ZN(new_n797));
  NOR3_X1   g611(.A1(new_n740), .A2(new_n589), .A3(new_n680), .ZN(new_n798));
  NOR2_X1   g612(.A1(new_n713), .A2(new_n714), .ZN(new_n799));
  INV_X1    g613(.A(new_n799), .ZN(new_n800));
  OR2_X1    g614(.A1(new_n800), .A2(KEYINPUT49), .ZN(new_n801));
  NAND2_X1  g615(.A1(new_n800), .A2(KEYINPUT49), .ZN(new_n802));
  NAND4_X1  g616(.A1(new_n797), .A2(new_n798), .A3(new_n801), .A4(new_n802), .ZN(new_n803));
  AND2_X1   g617(.A1(new_n734), .A2(new_n192), .ZN(new_n804));
  NAND4_X1  g618(.A1(new_n777), .A2(new_n636), .A3(new_n695), .A4(new_n688), .ZN(new_n805));
  INV_X1    g619(.A(new_n805), .ZN(new_n806));
  NAND3_X1  g620(.A1(new_n804), .A2(new_n682), .A3(new_n806), .ZN(new_n807));
  NAND4_X1  g621(.A1(new_n671), .A2(new_n698), .A3(new_n730), .A4(new_n807), .ZN(new_n808));
  NAND2_X1  g622(.A1(new_n808), .A2(KEYINPUT52), .ZN(new_n809));
  OAI211_X1 g623(.A(new_n752), .B(new_n715), .C1(new_n652), .C2(new_n700), .ZN(new_n810));
  NAND3_X1  g624(.A1(new_n810), .A2(new_n717), .A3(new_n725), .ZN(new_n811));
  NAND3_X1  g625(.A1(new_n645), .A2(new_n496), .A3(new_n494), .ZN(new_n812));
  NOR3_X1   g626(.A1(new_n650), .A2(new_n406), .A3(new_n669), .ZN(new_n813));
  INV_X1    g627(.A(new_n813), .ZN(new_n814));
  AOI21_X1  g628(.A(new_n814), .B1(new_n664), .B2(new_n590), .ZN(new_n815));
  NAND4_X1  g629(.A1(new_n812), .A2(new_n815), .A3(new_n192), .A4(new_n659), .ZN(new_n816));
  OAI22_X1  g630(.A1(new_n816), .A2(new_n776), .B1(new_n738), .B2(new_n758), .ZN(new_n817));
  NOR2_X1   g631(.A1(new_n811), .A2(new_n817), .ZN(new_n818));
  NOR3_X1   g632(.A1(new_n659), .A2(new_n681), .A3(new_n805), .ZN(new_n819));
  AOI21_X1  g633(.A(KEYINPUT52), .B1(new_n819), .B2(new_n804), .ZN(new_n820));
  NAND4_X1  g634(.A1(new_n820), .A2(new_n671), .A3(new_n698), .A4(new_n730), .ZN(new_n821));
  AND2_X1   g635(.A1(new_n659), .A2(new_n721), .ZN(new_n822));
  NAND2_X1  g636(.A1(new_n739), .A2(new_n822), .ZN(new_n823));
  NAND4_X1  g637(.A1(new_n809), .A2(new_n818), .A3(new_n821), .A4(new_n823), .ZN(new_n824));
  NAND2_X1  g638(.A1(new_n646), .A2(new_n647), .ZN(new_n825));
  INV_X1    g639(.A(KEYINPUT103), .ZN(new_n826));
  OAI21_X1  g640(.A(new_n650), .B1(new_n407), .B2(new_n424), .ZN(new_n827));
  OAI21_X1  g641(.A(new_n826), .B1(new_n295), .B2(new_n827), .ZN(new_n828));
  AOI21_X1  g642(.A(new_n334), .B1(new_n614), .B2(new_n615), .ZN(new_n829));
  NAND4_X1  g643(.A1(new_n686), .A2(new_n829), .A3(KEYINPUT103), .A4(new_n294), .ZN(new_n830));
  NAND2_X1  g644(.A1(new_n828), .A2(new_n830), .ZN(new_n831));
  OAI221_X1 g645(.A(KEYINPUT104), .B1(new_n498), .B2(new_n660), .C1(new_n825), .C2(new_n831), .ZN(new_n832));
  INV_X1    g646(.A(KEYINPUT104), .ZN(new_n833));
  NOR3_X1   g647(.A1(new_n613), .A2(new_n831), .A3(new_n633), .ZN(new_n834));
  OAI21_X1  g648(.A(new_n833), .B1(new_n834), .B2(new_n661), .ZN(new_n835));
  INV_X1    g649(.A(new_n295), .ZN(new_n836));
  AOI21_X1  g650(.A(new_n611), .B1(new_n634), .B2(new_n836), .ZN(new_n837));
  NAND3_X1  g651(.A1(new_n832), .A2(new_n835), .A3(new_n837), .ZN(new_n838));
  NOR3_X1   g652(.A1(new_n824), .A2(new_n756), .A3(new_n838), .ZN(new_n839));
  NOR2_X1   g653(.A1(new_n839), .A2(KEYINPUT53), .ZN(new_n840));
  AOI21_X1  g654(.A(new_n706), .B1(new_n701), .B2(new_n710), .ZN(new_n841));
  NAND4_X1  g655(.A1(new_n659), .A2(new_n604), .A3(new_n716), .A4(new_n638), .ZN(new_n842));
  NAND4_X1  g656(.A1(new_n724), .A2(new_n705), .A3(new_n192), .A4(new_n494), .ZN(new_n843));
  OAI22_X1  g657(.A1(new_n842), .A2(new_n706), .B1(new_n843), .B2(new_n722), .ZN(new_n844));
  NOR2_X1   g658(.A1(new_n841), .A2(new_n844), .ZN(new_n845));
  NAND3_X1  g659(.A1(new_n659), .A2(new_n604), .A3(new_n813), .ZN(new_n846));
  NOR2_X1   g660(.A1(new_n613), .A2(new_n846), .ZN(new_n847));
  INV_X1    g661(.A(new_n758), .ZN(new_n848));
  AOI22_X1  g662(.A1(new_n847), .A2(new_n793), .B1(new_n750), .B2(new_n848), .ZN(new_n849));
  AND4_X1   g663(.A1(new_n821), .A2(new_n823), .A3(new_n845), .A4(new_n849), .ZN(new_n850));
  AND3_X1   g664(.A1(new_n832), .A2(new_n835), .A3(new_n837), .ZN(new_n851));
  INV_X1    g665(.A(new_n747), .ZN(new_n852));
  OAI21_X1  g666(.A(new_n852), .B1(new_n753), .B2(new_n754), .ZN(new_n853));
  NOR2_X1   g667(.A1(new_n748), .A2(KEYINPUT98), .ZN(new_n854));
  OAI21_X1  g668(.A(new_n745), .B1(new_n853), .B2(new_n854), .ZN(new_n855));
  NAND4_X1  g669(.A1(new_n850), .A2(new_n851), .A3(new_n855), .A4(new_n809), .ZN(new_n856));
  INV_X1    g670(.A(KEYINPUT53), .ZN(new_n857));
  NOR2_X1   g671(.A1(new_n856), .A2(new_n857), .ZN(new_n858));
  OAI21_X1  g672(.A(KEYINPUT54), .B1(new_n840), .B2(new_n858), .ZN(new_n859));
  INV_X1    g673(.A(KEYINPUT105), .ZN(new_n860));
  NAND2_X1  g674(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  OAI211_X1 g675(.A(KEYINPUT105), .B(KEYINPUT54), .C1(new_n840), .C2(new_n858), .ZN(new_n862));
  NAND2_X1  g676(.A1(new_n861), .A2(new_n862), .ZN(new_n863));
  INV_X1    g677(.A(KEYINPUT107), .ZN(new_n864));
  OAI21_X1  g678(.A(new_n864), .B1(new_n856), .B2(new_n857), .ZN(new_n865));
  NOR2_X1   g679(.A1(new_n824), .A2(new_n838), .ZN(new_n866));
  NAND4_X1  g680(.A1(new_n866), .A2(KEYINPUT107), .A3(KEYINPUT53), .A4(new_n855), .ZN(new_n867));
  NAND2_X1  g681(.A1(new_n865), .A2(new_n867), .ZN(new_n868));
  INV_X1    g682(.A(KEYINPUT54), .ZN(new_n869));
  OAI21_X1  g683(.A(KEYINPUT106), .B1(new_n839), .B2(KEYINPUT53), .ZN(new_n870));
  INV_X1    g684(.A(KEYINPUT106), .ZN(new_n871));
  NAND3_X1  g685(.A1(new_n856), .A2(new_n871), .A3(new_n857), .ZN(new_n872));
  NAND4_X1  g686(.A1(new_n868), .A2(new_n869), .A3(new_n870), .A4(new_n872), .ZN(new_n873));
  INV_X1    g687(.A(KEYINPUT108), .ZN(new_n874));
  NAND2_X1  g688(.A1(new_n873), .A2(new_n874), .ZN(new_n875));
  AND2_X1   g689(.A1(new_n870), .A2(new_n872), .ZN(new_n876));
  NAND4_X1  g690(.A1(new_n876), .A2(KEYINPUT108), .A3(new_n869), .A4(new_n868), .ZN(new_n877));
  NAND3_X1  g691(.A1(new_n863), .A2(new_n875), .A3(new_n877), .ZN(new_n878));
  INV_X1    g692(.A(G952), .ZN(new_n879));
  AND2_X1   g693(.A1(new_n780), .A2(new_n667), .ZN(new_n880));
  AND2_X1   g694(.A1(new_n880), .A2(new_n723), .ZN(new_n881));
  AOI211_X1 g695(.A(new_n879), .B(G953), .C1(new_n881), .C2(new_n729), .ZN(new_n882));
  NOR2_X1   g696(.A1(new_n776), .A2(new_n706), .ZN(new_n883));
  AND2_X1   g697(.A1(new_n880), .A2(new_n883), .ZN(new_n884));
  NAND4_X1  g698(.A1(new_n884), .A2(KEYINPUT111), .A3(KEYINPUT48), .A4(new_n744), .ZN(new_n885));
  NAND2_X1  g699(.A1(new_n884), .A2(new_n744), .ZN(new_n886));
  XOR2_X1   g700(.A(KEYINPUT111), .B(KEYINPUT48), .Z(new_n887));
  NAND2_X1  g701(.A1(new_n886), .A2(new_n887), .ZN(new_n888));
  AND3_X1   g702(.A1(new_n883), .A2(new_n287), .A3(new_n798), .ZN(new_n889));
  NAND2_X1  g703(.A1(new_n889), .A2(new_n694), .ZN(new_n890));
  NAND4_X1  g704(.A1(new_n882), .A2(new_n885), .A3(new_n888), .A4(new_n890), .ZN(new_n891));
  NAND2_X1  g705(.A1(new_n881), .A2(new_n793), .ZN(new_n892));
  NAND2_X1  g706(.A1(new_n799), .A2(new_n191), .ZN(new_n893));
  AOI21_X1  g707(.A(new_n892), .B1(new_n792), .B2(new_n893), .ZN(new_n894));
  AND2_X1   g708(.A1(new_n884), .A2(new_n822), .ZN(new_n895));
  NOR3_X1   g709(.A1(new_n687), .A2(new_n706), .A3(new_n292), .ZN(new_n896));
  NAND2_X1  g710(.A1(new_n881), .A2(new_n896), .ZN(new_n897));
  XNOR2_X1  g711(.A(new_n897), .B(KEYINPUT50), .ZN(new_n898));
  NOR2_X1   g712(.A1(new_n777), .A2(new_n623), .ZN(new_n899));
  AOI211_X1 g713(.A(new_n895), .B(new_n898), .C1(new_n889), .C2(new_n899), .ZN(new_n900));
  NOR2_X1   g714(.A1(new_n900), .A2(KEYINPUT110), .ZN(new_n901));
  OAI21_X1  g715(.A(KEYINPUT51), .B1(new_n894), .B2(new_n901), .ZN(new_n902));
  XNOR2_X1  g716(.A(new_n893), .B(KEYINPUT109), .ZN(new_n903));
  NAND3_X1  g717(.A1(new_n790), .A2(new_n791), .A3(new_n903), .ZN(new_n904));
  INV_X1    g718(.A(KEYINPUT51), .ZN(new_n905));
  NAND4_X1  g719(.A1(new_n904), .A2(new_n905), .A3(new_n793), .A4(new_n881), .ZN(new_n906));
  OAI211_X1 g720(.A(new_n906), .B(new_n900), .C1(KEYINPUT110), .C2(new_n905), .ZN(new_n907));
  AOI211_X1 g721(.A(new_n878), .B(new_n891), .C1(new_n902), .C2(new_n907), .ZN(new_n908));
  NOR2_X1   g722(.A1(G952), .A2(G953), .ZN(new_n909));
  XNOR2_X1  g723(.A(new_n909), .B(KEYINPUT112), .ZN(new_n910));
  OAI21_X1  g724(.A(new_n803), .B1(new_n908), .B2(new_n910), .ZN(G75));
  NAND2_X1  g725(.A1(new_n876), .A2(new_n868), .ZN(new_n912));
  NAND3_X1  g726(.A1(new_n912), .A2(G210), .A3(G902), .ZN(new_n913));
  INV_X1    g727(.A(KEYINPUT113), .ZN(new_n914));
  OR2_X1    g728(.A1(new_n913), .A2(new_n914), .ZN(new_n915));
  AOI21_X1  g729(.A(KEYINPUT56), .B1(new_n913), .B2(new_n914), .ZN(new_n916));
  NAND2_X1  g730(.A1(new_n915), .A2(new_n916), .ZN(new_n917));
  OAI21_X1  g731(.A(new_n240), .B1(new_n265), .B2(new_n266), .ZN(new_n918));
  XNOR2_X1  g732(.A(new_n918), .B(new_n261), .ZN(new_n919));
  XOR2_X1   g733(.A(new_n919), .B(KEYINPUT55), .Z(new_n920));
  NAND2_X1  g734(.A1(new_n917), .A2(new_n920), .ZN(new_n921));
  NOR2_X1   g735(.A1(new_n285), .A2(G952), .ZN(new_n922));
  INV_X1    g736(.A(new_n922), .ZN(new_n923));
  NAND2_X1  g737(.A1(new_n913), .A2(KEYINPUT114), .ZN(new_n924));
  INV_X1    g738(.A(KEYINPUT114), .ZN(new_n925));
  NAND4_X1  g739(.A1(new_n912), .A2(new_n925), .A3(G210), .A4(G902), .ZN(new_n926));
  NOR2_X1   g740(.A1(new_n920), .A2(KEYINPUT56), .ZN(new_n927));
  NAND3_X1  g741(.A1(new_n924), .A2(new_n926), .A3(new_n927), .ZN(new_n928));
  NAND4_X1  g742(.A1(new_n921), .A2(KEYINPUT115), .A3(new_n923), .A4(new_n928), .ZN(new_n929));
  INV_X1    g743(.A(KEYINPUT115), .ZN(new_n930));
  NAND2_X1  g744(.A1(new_n928), .A2(new_n923), .ZN(new_n931));
  INV_X1    g745(.A(new_n920), .ZN(new_n932));
  AOI21_X1  g746(.A(new_n932), .B1(new_n915), .B2(new_n916), .ZN(new_n933));
  OAI21_X1  g747(.A(new_n930), .B1(new_n931), .B2(new_n933), .ZN(new_n934));
  NAND2_X1  g748(.A1(new_n929), .A2(new_n934), .ZN(G51));
  AND2_X1   g749(.A1(new_n865), .A2(new_n867), .ZN(new_n936));
  NAND2_X1  g750(.A1(new_n870), .A2(new_n872), .ZN(new_n937));
  OAI21_X1  g751(.A(KEYINPUT54), .B1(new_n936), .B2(new_n937), .ZN(new_n938));
  INV_X1    g752(.A(KEYINPUT116), .ZN(new_n939));
  NAND3_X1  g753(.A1(new_n938), .A2(new_n939), .A3(new_n873), .ZN(new_n940));
  NAND3_X1  g754(.A1(new_n912), .A2(KEYINPUT116), .A3(KEYINPUT54), .ZN(new_n941));
  XNOR2_X1  g755(.A(new_n495), .B(KEYINPUT57), .ZN(new_n942));
  NAND3_X1  g756(.A1(new_n940), .A2(new_n941), .A3(new_n942), .ZN(new_n943));
  NAND2_X1  g757(.A1(new_n943), .A2(new_n703), .ZN(new_n944));
  NAND2_X1  g758(.A1(new_n912), .A2(G902), .ZN(new_n945));
  OR2_X1    g759(.A1(new_n945), .A2(new_n766), .ZN(new_n946));
  AOI21_X1  g760(.A(new_n922), .B1(new_n944), .B2(new_n946), .ZN(G54));
  INV_X1    g761(.A(KEYINPUT58), .ZN(new_n948));
  NOR3_X1   g762(.A1(new_n945), .A2(new_n948), .A3(new_n405), .ZN(new_n949));
  OAI21_X1  g763(.A(new_n923), .B1(new_n949), .B2(new_n397), .ZN(new_n950));
  AOI21_X1  g764(.A(new_n950), .B1(new_n397), .B2(new_n949), .ZN(G60));
  NAND2_X1  g765(.A1(new_n617), .A2(new_n619), .ZN(new_n952));
  XOR2_X1   g766(.A(new_n952), .B(KEYINPUT117), .Z(new_n953));
  XNOR2_X1  g767(.A(KEYINPUT118), .B(KEYINPUT59), .ZN(new_n954));
  XOR2_X1   g768(.A(new_n954), .B(new_n621), .Z(new_n955));
  NOR2_X1   g769(.A1(new_n953), .A2(new_n955), .ZN(new_n956));
  NAND3_X1  g770(.A1(new_n940), .A2(new_n941), .A3(new_n956), .ZN(new_n957));
  INV_X1    g771(.A(KEYINPUT119), .ZN(new_n958));
  NAND2_X1  g772(.A1(new_n957), .A2(new_n958), .ZN(new_n959));
  NAND4_X1  g773(.A1(new_n940), .A2(new_n941), .A3(KEYINPUT119), .A4(new_n956), .ZN(new_n960));
  NAND2_X1  g774(.A1(new_n959), .A2(new_n960), .ZN(new_n961));
  INV_X1    g775(.A(new_n955), .ZN(new_n962));
  NAND2_X1  g776(.A1(new_n878), .A2(new_n962), .ZN(new_n963));
  AOI21_X1  g777(.A(new_n922), .B1(new_n963), .B2(new_n953), .ZN(new_n964));
  NAND2_X1  g778(.A1(new_n961), .A2(new_n964), .ZN(new_n965));
  INV_X1    g779(.A(KEYINPUT120), .ZN(new_n966));
  NAND2_X1  g780(.A1(new_n965), .A2(new_n966), .ZN(new_n967));
  NAND3_X1  g781(.A1(new_n961), .A2(new_n964), .A3(KEYINPUT120), .ZN(new_n968));
  NAND2_X1  g782(.A1(new_n967), .A2(new_n968), .ZN(G63));
  INV_X1    g783(.A(KEYINPUT61), .ZN(new_n970));
  NAND2_X1  g784(.A1(G217), .A2(G902), .ZN(new_n971));
  XNOR2_X1  g785(.A(new_n971), .B(KEYINPUT122), .ZN(new_n972));
  XOR2_X1   g786(.A(KEYINPUT121), .B(KEYINPUT60), .Z(new_n973));
  XNOR2_X1  g787(.A(new_n972), .B(new_n973), .ZN(new_n974));
  NAND2_X1  g788(.A1(new_n912), .A2(new_n974), .ZN(new_n975));
  INV_X1    g789(.A(new_n607), .ZN(new_n976));
  NAND2_X1  g790(.A1(new_n975), .A2(new_n976), .ZN(new_n977));
  NAND3_X1  g791(.A1(new_n977), .A2(KEYINPUT123), .A3(new_n923), .ZN(new_n978));
  NAND3_X1  g792(.A1(new_n912), .A2(new_n657), .A3(new_n974), .ZN(new_n979));
  NAND2_X1  g793(.A1(new_n978), .A2(new_n979), .ZN(new_n980));
  AOI21_X1  g794(.A(KEYINPUT123), .B1(new_n977), .B2(new_n923), .ZN(new_n981));
  OAI21_X1  g795(.A(new_n970), .B1(new_n980), .B2(new_n981), .ZN(new_n982));
  INV_X1    g796(.A(KEYINPUT124), .ZN(new_n983));
  NOR2_X1   g797(.A1(new_n977), .A2(new_n983), .ZN(new_n984));
  NAND2_X1  g798(.A1(new_n977), .A2(new_n983), .ZN(new_n985));
  NOR2_X1   g799(.A1(new_n922), .A2(new_n970), .ZN(new_n986));
  NAND3_X1  g800(.A1(new_n985), .A2(new_n979), .A3(new_n986), .ZN(new_n987));
  OAI21_X1  g801(.A(new_n982), .B1(new_n984), .B2(new_n987), .ZN(G66));
  OAI21_X1  g802(.A(G953), .B1(new_n290), .B2(new_n259), .ZN(new_n989));
  NOR2_X1   g803(.A1(new_n838), .A2(new_n811), .ZN(new_n990));
  OAI21_X1  g804(.A(new_n989), .B1(new_n990), .B2(G953), .ZN(new_n991));
  OAI21_X1  g805(.A(new_n918), .B1(G898), .B2(new_n285), .ZN(new_n992));
  XNOR2_X1  g806(.A(new_n991), .B(new_n992), .ZN(G69));
  NAND2_X1  g807(.A1(new_n384), .A2(new_n386), .ZN(new_n994));
  XOR2_X1   g808(.A(new_n994), .B(KEYINPUT125), .Z(new_n995));
  XNOR2_X1  g809(.A(new_n581), .B(new_n995), .ZN(new_n996));
  OR2_X1    g810(.A1(new_n792), .A2(new_n794), .ZN(new_n997));
  NAND3_X1  g811(.A1(new_n671), .A2(new_n698), .A3(new_n730), .ZN(new_n998));
  NOR2_X1   g812(.A1(new_n692), .A2(new_n998), .ZN(new_n999));
  XOR2_X1   g813(.A(new_n999), .B(KEYINPUT62), .Z(new_n1000));
  OAI21_X1  g814(.A(new_n752), .B1(new_n694), .B2(new_n829), .ZN(new_n1001));
  NOR3_X1   g815(.A1(new_n674), .A2(new_n1001), .A3(new_n776), .ZN(new_n1002));
  NOR2_X1   g816(.A1(new_n1000), .A2(new_n1002), .ZN(new_n1003));
  AND2_X1   g817(.A1(new_n787), .A2(new_n1003), .ZN(new_n1004));
  NAND2_X1  g818(.A1(new_n997), .A2(new_n1004), .ZN(new_n1005));
  AOI21_X1  g819(.A(new_n996), .B1(new_n1005), .B2(new_n285), .ZN(new_n1006));
  INV_X1    g820(.A(new_n996), .ZN(new_n1007));
  AOI21_X1  g821(.A(new_n1007), .B1(G900), .B2(G953), .ZN(new_n1008));
  INV_X1    g822(.A(new_n1008), .ZN(new_n1009));
  NOR3_X1   g823(.A1(new_n756), .A2(new_n759), .A3(new_n998), .ZN(new_n1010));
  NAND2_X1  g824(.A1(new_n775), .A2(new_n673), .ZN(new_n1011));
  NOR2_X1   g825(.A1(new_n689), .A2(new_n685), .ZN(new_n1012));
  AOI21_X1  g826(.A(new_n786), .B1(new_n1012), .B2(new_n744), .ZN(new_n1013));
  OAI21_X1  g827(.A(new_n1010), .B1(new_n1011), .B2(new_n1013), .ZN(new_n1014));
  NOR2_X1   g828(.A1(new_n795), .A2(new_n1014), .ZN(new_n1015));
  AOI21_X1  g829(.A(new_n1009), .B1(new_n1015), .B2(new_n285), .ZN(new_n1016));
  AOI21_X1  g830(.A(new_n285), .B1(G227), .B2(G900), .ZN(new_n1017));
  OR3_X1    g831(.A1(new_n1006), .A2(new_n1016), .A3(new_n1017), .ZN(new_n1018));
  OAI21_X1  g832(.A(new_n1017), .B1(new_n1006), .B2(new_n1016), .ZN(new_n1019));
  NAND2_X1  g833(.A1(new_n1018), .A2(new_n1019), .ZN(G72));
  NAND2_X1  g834(.A1(new_n582), .A2(new_n596), .ZN(new_n1021));
  NAND2_X1  g835(.A1(new_n1015), .A2(new_n990), .ZN(new_n1022));
  NAND2_X1  g836(.A1(G472), .A2(G902), .ZN(new_n1023));
  XNOR2_X1  g837(.A(new_n1023), .B(KEYINPUT127), .ZN(new_n1024));
  XOR2_X1   g838(.A(KEYINPUT126), .B(KEYINPUT63), .Z(new_n1025));
  XNOR2_X1  g839(.A(new_n1024), .B(new_n1025), .ZN(new_n1026));
  AOI21_X1  g840(.A(new_n1021), .B1(new_n1022), .B2(new_n1026), .ZN(new_n1027));
  OR2_X1    g841(.A1(new_n582), .A2(new_n596), .ZN(new_n1028));
  NAND3_X1  g842(.A1(new_n997), .A2(new_n990), .A3(new_n1004), .ZN(new_n1029));
  AOI21_X1  g843(.A(new_n1028), .B1(new_n1029), .B2(new_n1026), .ZN(new_n1030));
  NOR2_X1   g844(.A1(new_n840), .A2(new_n858), .ZN(new_n1031));
  NAND3_X1  g845(.A1(new_n1028), .A2(new_n1026), .A3(new_n1021), .ZN(new_n1032));
  OAI21_X1  g846(.A(new_n923), .B1(new_n1031), .B2(new_n1032), .ZN(new_n1033));
  NOR3_X1   g847(.A1(new_n1027), .A2(new_n1030), .A3(new_n1033), .ZN(G57));
endmodule


