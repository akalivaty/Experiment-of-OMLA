//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 1 0 1 1 1 1 1 1 1 1 0 1 0 0 1 0 1 1 0 0 0 0 1 1 0 1 0 1 0 0 1 1 0 0 0 1 1 1 0 0 1 1 1 1 0 1 0 1 1 0 0 0 0 0 0 1 1 0 1 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:19:06 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n677, new_n678,
    new_n679, new_n680, new_n681, new_n682, new_n683, new_n684, new_n685,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n692, new_n693,
    new_n694, new_n696, new_n697, new_n698, new_n699, new_n700, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n728, new_n729, new_n730, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n750, new_n751, new_n752, new_n753, new_n755, new_n756,
    new_n757, new_n758, new_n759, new_n761, new_n762, new_n763, new_n765,
    new_n767, new_n768, new_n769, new_n770, new_n771, new_n772, new_n773,
    new_n774, new_n775, new_n776, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n789,
    new_n790, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n831, new_n832, new_n833, new_n834,
    new_n836, new_n838, new_n839, new_n840, new_n841, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n868, new_n869, new_n871, new_n872, new_n873, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n883, new_n884,
    new_n886, new_n887, new_n888, new_n889, new_n890, new_n891, new_n892,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n909,
    new_n910, new_n911, new_n913, new_n914, new_n915, new_n916, new_n918,
    new_n919, new_n920;
  XOR2_X1   g000(.A(G113gat), .B(G120gat), .Z(new_n202));
  INV_X1    g001(.A(KEYINPUT1), .ZN(new_n203));
  INV_X1    g002(.A(KEYINPUT69), .ZN(new_n204));
  XNOR2_X1  g003(.A(G127gat), .B(G134gat), .ZN(new_n205));
  OAI211_X1 g004(.A(new_n202), .B(new_n203), .C1(new_n204), .C2(new_n205), .ZN(new_n206));
  XOR2_X1   g005(.A(G127gat), .B(G134gat), .Z(new_n207));
  NAND2_X1  g006(.A1(new_n204), .A2(new_n203), .ZN(new_n208));
  XNOR2_X1  g007(.A(G113gat), .B(G120gat), .ZN(new_n209));
  OAI211_X1 g008(.A(new_n207), .B(new_n208), .C1(KEYINPUT1), .C2(new_n209), .ZN(new_n210));
  AND2_X1   g009(.A1(new_n206), .A2(new_n210), .ZN(new_n211));
  AND2_X1   g010(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n212));
  NOR2_X1   g011(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n213));
  OR2_X1    g012(.A1(new_n212), .A2(new_n213), .ZN(new_n214));
  INV_X1    g013(.A(G190gat), .ZN(new_n215));
  OAI21_X1  g014(.A(KEYINPUT68), .B1(KEYINPUT67), .B2(KEYINPUT28), .ZN(new_n216));
  OR2_X1    g015(.A1(KEYINPUT68), .A2(KEYINPUT28), .ZN(new_n217));
  NAND4_X1  g016(.A1(new_n214), .A2(new_n215), .A3(new_n216), .A4(new_n217), .ZN(new_n218));
  OAI21_X1  g017(.A(new_n215), .B1(new_n212), .B2(new_n213), .ZN(new_n219));
  INV_X1    g018(.A(new_n216), .ZN(new_n220));
  AOI22_X1  g019(.A1(new_n219), .A2(new_n220), .B1(G183gat), .B2(G190gat), .ZN(new_n221));
  NAND2_X1  g020(.A1(G169gat), .A2(G176gat), .ZN(new_n222));
  INV_X1    g021(.A(G169gat), .ZN(new_n223));
  INV_X1    g022(.A(G176gat), .ZN(new_n224));
  AND3_X1   g023(.A1(new_n223), .A2(new_n224), .A3(KEYINPUT26), .ZN(new_n225));
  AOI21_X1  g024(.A(KEYINPUT26), .B1(new_n223), .B2(new_n224), .ZN(new_n226));
  OAI21_X1  g025(.A(new_n222), .B1(new_n225), .B2(new_n226), .ZN(new_n227));
  NAND3_X1  g026(.A1(new_n218), .A2(new_n221), .A3(new_n227), .ZN(new_n228));
  NAND3_X1  g027(.A1(new_n223), .A2(new_n224), .A3(KEYINPUT23), .ZN(new_n229));
  INV_X1    g028(.A(KEYINPUT23), .ZN(new_n230));
  OAI21_X1  g029(.A(new_n230), .B1(G169gat), .B2(G176gat), .ZN(new_n231));
  NAND3_X1  g030(.A1(new_n229), .A2(new_n231), .A3(new_n222), .ZN(new_n232));
  INV_X1    g031(.A(KEYINPUT65), .ZN(new_n233));
  NAND2_X1  g032(.A1(new_n232), .A2(new_n233), .ZN(new_n234));
  INV_X1    g033(.A(KEYINPUT64), .ZN(new_n235));
  INV_X1    g034(.A(G183gat), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n236), .A2(new_n215), .ZN(new_n237));
  NAND3_X1  g036(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n238));
  NAND2_X1  g037(.A1(new_n237), .A2(new_n238), .ZN(new_n239));
  AOI21_X1  g038(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n240));
  OAI21_X1  g039(.A(new_n235), .B1(new_n239), .B2(new_n240), .ZN(new_n241));
  OR2_X1    g040(.A1(KEYINPUT65), .A2(KEYINPUT25), .ZN(new_n242));
  NAND4_X1  g041(.A1(new_n229), .A2(new_n231), .A3(new_n222), .A4(new_n242), .ZN(new_n243));
  INV_X1    g042(.A(new_n240), .ZN(new_n244));
  NAND4_X1  g043(.A1(new_n244), .A2(KEYINPUT64), .A3(new_n238), .A4(new_n237), .ZN(new_n245));
  NAND4_X1  g044(.A1(new_n234), .A2(new_n241), .A3(new_n243), .A4(new_n245), .ZN(new_n246));
  NOR2_X1   g045(.A1(new_n239), .A2(new_n240), .ZN(new_n247));
  OAI21_X1  g046(.A(KEYINPUT25), .B1(new_n247), .B2(new_n232), .ZN(new_n248));
  AND3_X1   g047(.A1(new_n246), .A2(KEYINPUT66), .A3(new_n248), .ZN(new_n249));
  AOI21_X1  g048(.A(KEYINPUT66), .B1(new_n246), .B2(new_n248), .ZN(new_n250));
  OAI211_X1 g049(.A(new_n211), .B(new_n228), .C1(new_n249), .C2(new_n250), .ZN(new_n251));
  INV_X1    g050(.A(KEYINPUT70), .ZN(new_n252));
  NAND2_X1  g051(.A1(new_n251), .A2(new_n252), .ZN(new_n253));
  NAND2_X1  g052(.A1(new_n246), .A2(new_n248), .ZN(new_n254));
  INV_X1    g053(.A(KEYINPUT66), .ZN(new_n255));
  NAND2_X1  g054(.A1(new_n254), .A2(new_n255), .ZN(new_n256));
  NAND3_X1  g055(.A1(new_n246), .A2(KEYINPUT66), .A3(new_n248), .ZN(new_n257));
  NAND2_X1  g056(.A1(new_n256), .A2(new_n257), .ZN(new_n258));
  NAND4_X1  g057(.A1(new_n258), .A2(KEYINPUT70), .A3(new_n211), .A4(new_n228), .ZN(new_n259));
  OAI21_X1  g058(.A(new_n228), .B1(new_n249), .B2(new_n250), .ZN(new_n260));
  NAND2_X1  g059(.A1(new_n206), .A2(new_n210), .ZN(new_n261));
  NAND2_X1  g060(.A1(new_n260), .A2(new_n261), .ZN(new_n262));
  NAND3_X1  g061(.A1(new_n253), .A2(new_n259), .A3(new_n262), .ZN(new_n263));
  NAND2_X1  g062(.A1(G227gat), .A2(G233gat), .ZN(new_n264));
  INV_X1    g063(.A(new_n264), .ZN(new_n265));
  AOI21_X1  g064(.A(KEYINPUT33), .B1(new_n263), .B2(new_n265), .ZN(new_n266));
  NOR2_X1   g065(.A1(new_n263), .A2(new_n265), .ZN(new_n267));
  XNOR2_X1  g066(.A(G15gat), .B(G43gat), .ZN(new_n268));
  XNOR2_X1  g067(.A(G71gat), .B(G99gat), .ZN(new_n269));
  XOR2_X1   g068(.A(new_n268), .B(new_n269), .Z(new_n270));
  INV_X1    g069(.A(new_n270), .ZN(new_n271));
  NOR3_X1   g070(.A1(new_n266), .A2(new_n267), .A3(new_n271), .ZN(new_n272));
  AND3_X1   g071(.A1(new_n253), .A2(new_n259), .A3(new_n262), .ZN(new_n273));
  INV_X1    g072(.A(KEYINPUT33), .ZN(new_n274));
  OAI211_X1 g073(.A(new_n273), .B(new_n264), .C1(new_n274), .C2(new_n271), .ZN(new_n275));
  INV_X1    g074(.A(new_n275), .ZN(new_n276));
  INV_X1    g075(.A(KEYINPUT34), .ZN(new_n277));
  NAND2_X1  g076(.A1(new_n263), .A2(new_n265), .ZN(new_n278));
  AOI21_X1  g077(.A(new_n277), .B1(new_n278), .B2(KEYINPUT32), .ZN(new_n279));
  INV_X1    g078(.A(KEYINPUT32), .ZN(new_n280));
  AOI211_X1 g079(.A(new_n280), .B(KEYINPUT34), .C1(new_n263), .C2(new_n265), .ZN(new_n281));
  OAI22_X1  g080(.A1(new_n272), .A2(new_n276), .B1(new_n279), .B2(new_n281), .ZN(new_n282));
  NAND2_X1  g081(.A1(new_n278), .A2(new_n274), .ZN(new_n283));
  NAND2_X1  g082(.A1(new_n273), .A2(new_n264), .ZN(new_n284));
  NAND3_X1  g083(.A1(new_n283), .A2(new_n284), .A3(new_n270), .ZN(new_n285));
  NAND2_X1  g084(.A1(new_n278), .A2(KEYINPUT32), .ZN(new_n286));
  NAND2_X1  g085(.A1(new_n286), .A2(KEYINPUT34), .ZN(new_n287));
  NAND3_X1  g086(.A1(new_n278), .A2(KEYINPUT32), .A3(new_n277), .ZN(new_n288));
  NAND4_X1  g087(.A1(new_n285), .A2(new_n287), .A3(new_n288), .A4(new_n275), .ZN(new_n289));
  XNOR2_X1  g088(.A(G78gat), .B(G106gat), .ZN(new_n290));
  XNOR2_X1  g089(.A(KEYINPUT31), .B(G50gat), .ZN(new_n291));
  XOR2_X1   g090(.A(new_n290), .B(new_n291), .Z(new_n292));
  INV_X1    g091(.A(new_n292), .ZN(new_n293));
  INV_X1    g092(.A(G228gat), .ZN(new_n294));
  INV_X1    g093(.A(G233gat), .ZN(new_n295));
  NOR2_X1   g094(.A1(new_n294), .A2(new_n295), .ZN(new_n296));
  INV_X1    g095(.A(new_n296), .ZN(new_n297));
  XOR2_X1   g096(.A(G211gat), .B(G218gat), .Z(new_n298));
  AOI21_X1  g097(.A(KEYINPUT22), .B1(G211gat), .B2(G218gat), .ZN(new_n299));
  AND2_X1   g098(.A1(G197gat), .A2(G204gat), .ZN(new_n300));
  NOR2_X1   g099(.A1(G197gat), .A2(G204gat), .ZN(new_n301));
  NOR2_X1   g100(.A1(new_n300), .A2(new_n301), .ZN(new_n302));
  OAI21_X1  g101(.A(new_n298), .B1(new_n299), .B2(new_n302), .ZN(new_n303));
  XNOR2_X1  g102(.A(G211gat), .B(G218gat), .ZN(new_n304));
  INV_X1    g103(.A(new_n299), .ZN(new_n305));
  OAI211_X1 g104(.A(new_n304), .B(new_n305), .C1(new_n301), .C2(new_n300), .ZN(new_n306));
  NAND3_X1  g105(.A1(new_n303), .A2(new_n306), .A3(KEYINPUT71), .ZN(new_n307));
  INV_X1    g106(.A(KEYINPUT29), .ZN(new_n308));
  INV_X1    g107(.A(KEYINPUT71), .ZN(new_n309));
  OAI211_X1 g108(.A(new_n298), .B(new_n309), .C1(new_n299), .C2(new_n302), .ZN(new_n310));
  NAND3_X1  g109(.A1(new_n307), .A2(new_n308), .A3(new_n310), .ZN(new_n311));
  INV_X1    g110(.A(KEYINPUT3), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n311), .A2(new_n312), .ZN(new_n313));
  NAND2_X1  g112(.A1(G155gat), .A2(G162gat), .ZN(new_n314));
  NAND2_X1  g113(.A1(new_n314), .A2(KEYINPUT2), .ZN(new_n315));
  NAND2_X1  g114(.A1(new_n315), .A2(KEYINPUT76), .ZN(new_n316));
  XNOR2_X1  g115(.A(G155gat), .B(G162gat), .ZN(new_n317));
  XNOR2_X1  g116(.A(G141gat), .B(G148gat), .ZN(new_n318));
  AND2_X1   g117(.A1(new_n314), .A2(KEYINPUT2), .ZN(new_n319));
  OAI211_X1 g118(.A(new_n316), .B(new_n317), .C1(new_n318), .C2(new_n319), .ZN(new_n320));
  INV_X1    g119(.A(G141gat), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n321), .A2(G148gat), .ZN(new_n322));
  INV_X1    g121(.A(G148gat), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n323), .A2(G141gat), .ZN(new_n324));
  NAND2_X1  g123(.A1(new_n322), .A2(new_n324), .ZN(new_n325));
  AND2_X1   g124(.A1(G155gat), .A2(G162gat), .ZN(new_n326));
  NOR2_X1   g125(.A1(G155gat), .A2(G162gat), .ZN(new_n327));
  NOR2_X1   g126(.A1(new_n326), .A2(new_n327), .ZN(new_n328));
  OAI211_X1 g127(.A(new_n315), .B(new_n325), .C1(new_n328), .C2(KEYINPUT76), .ZN(new_n329));
  AND2_X1   g128(.A1(new_n320), .A2(new_n329), .ZN(new_n330));
  AOI21_X1  g129(.A(new_n297), .B1(new_n313), .B2(new_n330), .ZN(new_n331));
  INV_X1    g130(.A(KEYINPUT77), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n320), .A2(new_n329), .ZN(new_n333));
  AOI21_X1  g132(.A(new_n332), .B1(new_n333), .B2(new_n312), .ZN(new_n334));
  AOI211_X1 g133(.A(KEYINPUT77), .B(KEYINPUT3), .C1(new_n320), .C2(new_n329), .ZN(new_n335));
  OAI21_X1  g134(.A(new_n308), .B1(new_n334), .B2(new_n335), .ZN(new_n336));
  INV_X1    g135(.A(new_n336), .ZN(new_n337));
  NAND2_X1  g136(.A1(new_n307), .A2(new_n310), .ZN(new_n338));
  INV_X1    g137(.A(KEYINPUT72), .ZN(new_n339));
  NAND2_X1  g138(.A1(new_n338), .A2(new_n339), .ZN(new_n340));
  NAND3_X1  g139(.A1(new_n307), .A2(KEYINPUT72), .A3(new_n310), .ZN(new_n341));
  NAND2_X1  g140(.A1(new_n340), .A2(new_n341), .ZN(new_n342));
  OAI21_X1  g141(.A(new_n331), .B1(new_n337), .B2(new_n342), .ZN(new_n343));
  INV_X1    g142(.A(G22gat), .ZN(new_n344));
  NAND2_X1  g143(.A1(new_n303), .A2(new_n306), .ZN(new_n345));
  NAND2_X1  g144(.A1(new_n345), .A2(new_n308), .ZN(new_n346));
  AOI21_X1  g145(.A(new_n333), .B1(new_n346), .B2(new_n312), .ZN(new_n347));
  AOI21_X1  g146(.A(new_n347), .B1(new_n336), .B2(new_n338), .ZN(new_n348));
  OAI211_X1 g147(.A(new_n343), .B(new_n344), .C1(new_n296), .C2(new_n348), .ZN(new_n349));
  INV_X1    g148(.A(new_n349), .ZN(new_n350));
  INV_X1    g149(.A(new_n338), .ZN(new_n351));
  NAND2_X1  g150(.A1(new_n333), .A2(new_n312), .ZN(new_n352));
  NAND2_X1  g151(.A1(new_n352), .A2(KEYINPUT77), .ZN(new_n353));
  NAND3_X1  g152(.A1(new_n333), .A2(new_n332), .A3(new_n312), .ZN(new_n354));
  NAND2_X1  g153(.A1(new_n353), .A2(new_n354), .ZN(new_n355));
  AOI21_X1  g154(.A(new_n351), .B1(new_n355), .B2(new_n308), .ZN(new_n356));
  OAI21_X1  g155(.A(new_n297), .B1(new_n356), .B2(new_n347), .ZN(new_n357));
  AOI21_X1  g156(.A(new_n344), .B1(new_n357), .B2(new_n343), .ZN(new_n358));
  OAI21_X1  g157(.A(KEYINPUT83), .B1(new_n350), .B2(new_n358), .ZN(new_n359));
  NAND2_X1  g158(.A1(new_n357), .A2(new_n343), .ZN(new_n360));
  NAND2_X1  g159(.A1(new_n360), .A2(G22gat), .ZN(new_n361));
  INV_X1    g160(.A(KEYINPUT83), .ZN(new_n362));
  NAND3_X1  g161(.A1(new_n361), .A2(new_n362), .A3(new_n349), .ZN(new_n363));
  AOI21_X1  g162(.A(new_n293), .B1(new_n359), .B2(new_n363), .ZN(new_n364));
  NAND2_X1  g163(.A1(new_n361), .A2(new_n349), .ZN(new_n365));
  AOI21_X1  g164(.A(new_n292), .B1(new_n365), .B2(KEYINPUT83), .ZN(new_n366));
  OAI211_X1 g165(.A(new_n282), .B(new_n289), .C1(new_n364), .C2(new_n366), .ZN(new_n367));
  XOR2_X1   g166(.A(KEYINPUT80), .B(KEYINPUT0), .Z(new_n368));
  XNOR2_X1  g167(.A(G1gat), .B(G29gat), .ZN(new_n369));
  XNOR2_X1  g168(.A(new_n368), .B(new_n369), .ZN(new_n370));
  XNOR2_X1  g169(.A(G57gat), .B(G85gat), .ZN(new_n371));
  XOR2_X1   g170(.A(new_n370), .B(new_n371), .Z(new_n372));
  INV_X1    g171(.A(new_n372), .ZN(new_n373));
  XNOR2_X1  g172(.A(KEYINPUT78), .B(KEYINPUT4), .ZN(new_n374));
  NAND4_X1  g173(.A1(new_n333), .A2(new_n206), .A3(new_n210), .A4(new_n374), .ZN(new_n375));
  NAND3_X1  g174(.A1(new_n333), .A2(new_n206), .A3(new_n210), .ZN(new_n376));
  AOI22_X1  g175(.A1(KEYINPUT81), .A2(new_n375), .B1(new_n376), .B2(KEYINPUT4), .ZN(new_n377));
  INV_X1    g176(.A(KEYINPUT81), .ZN(new_n378));
  NAND4_X1  g177(.A1(new_n211), .A2(new_n378), .A3(new_n333), .A4(new_n374), .ZN(new_n379));
  AOI22_X1  g178(.A1(new_n330), .A2(KEYINPUT3), .B1(new_n206), .B2(new_n210), .ZN(new_n380));
  AOI22_X1  g179(.A1(new_n377), .A2(new_n379), .B1(new_n355), .B2(new_n380), .ZN(new_n381));
  INV_X1    g180(.A(KEYINPUT82), .ZN(new_n382));
  NAND2_X1  g181(.A1(G225gat), .A2(G233gat), .ZN(new_n383));
  INV_X1    g182(.A(new_n383), .ZN(new_n384));
  NOR2_X1   g183(.A1(new_n384), .A2(KEYINPUT5), .ZN(new_n385));
  NAND3_X1  g184(.A1(new_n381), .A2(new_n382), .A3(new_n385), .ZN(new_n386));
  NAND2_X1  g185(.A1(new_n375), .A2(KEYINPUT81), .ZN(new_n387));
  NAND2_X1  g186(.A1(new_n376), .A2(KEYINPUT4), .ZN(new_n388));
  NAND3_X1  g187(.A1(new_n387), .A2(new_n379), .A3(new_n388), .ZN(new_n389));
  OAI21_X1  g188(.A(new_n380), .B1(new_n334), .B2(new_n335), .ZN(new_n390));
  NAND3_X1  g189(.A1(new_n389), .A2(new_n390), .A3(new_n385), .ZN(new_n391));
  NAND2_X1  g190(.A1(new_n391), .A2(KEYINPUT82), .ZN(new_n392));
  NAND2_X1  g191(.A1(new_n386), .A2(new_n392), .ZN(new_n393));
  XNOR2_X1  g192(.A(new_n261), .B(new_n333), .ZN(new_n394));
  OAI21_X1  g193(.A(KEYINPUT5), .B1(new_n394), .B2(new_n383), .ZN(new_n395));
  INV_X1    g194(.A(KEYINPUT79), .ZN(new_n396));
  OR2_X1    g195(.A1(new_n395), .A2(new_n396), .ZN(new_n397));
  NAND2_X1  g196(.A1(new_n376), .A2(new_n374), .ZN(new_n398));
  NAND3_X1  g197(.A1(new_n211), .A2(KEYINPUT4), .A3(new_n333), .ZN(new_n399));
  AND3_X1   g198(.A1(new_n398), .A2(new_n383), .A3(new_n399), .ZN(new_n400));
  AOI22_X1  g199(.A1(new_n395), .A2(new_n396), .B1(new_n400), .B2(new_n390), .ZN(new_n401));
  NAND2_X1  g200(.A1(new_n397), .A2(new_n401), .ZN(new_n402));
  AOI21_X1  g201(.A(new_n373), .B1(new_n393), .B2(new_n402), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n403), .A2(KEYINPUT6), .ZN(new_n404));
  INV_X1    g203(.A(KEYINPUT6), .ZN(new_n405));
  AOI22_X1  g204(.A1(new_n392), .A2(new_n386), .B1(new_n397), .B2(new_n401), .ZN(new_n406));
  OAI21_X1  g205(.A(new_n405), .B1(new_n406), .B2(new_n373), .ZN(new_n407));
  AND3_X1   g206(.A1(new_n393), .A2(new_n402), .A3(new_n373), .ZN(new_n408));
  OAI21_X1  g207(.A(new_n404), .B1(new_n407), .B2(new_n408), .ZN(new_n409));
  NAND3_X1  g208(.A1(new_n228), .A2(new_n246), .A3(new_n248), .ZN(new_n410));
  NAND2_X1  g209(.A1(new_n410), .A2(new_n308), .ZN(new_n411));
  NAND2_X1  g210(.A1(G226gat), .A2(G233gat), .ZN(new_n412));
  XOR2_X1   g211(.A(new_n412), .B(KEYINPUT73), .Z(new_n413));
  INV_X1    g212(.A(new_n413), .ZN(new_n414));
  NAND2_X1  g213(.A1(new_n411), .A2(new_n414), .ZN(new_n415));
  INV_X1    g214(.A(new_n228), .ZN(new_n416));
  AOI21_X1  g215(.A(new_n416), .B1(new_n256), .B2(new_n257), .ZN(new_n417));
  XOR2_X1   g216(.A(new_n413), .B(KEYINPUT74), .Z(new_n418));
  OAI211_X1 g217(.A(new_n415), .B(new_n351), .C1(new_n417), .C2(new_n418), .ZN(new_n419));
  INV_X1    g218(.A(new_n419), .ZN(new_n420));
  INV_X1    g219(.A(new_n342), .ZN(new_n421));
  OAI21_X1  g220(.A(new_n418), .B1(new_n417), .B2(KEYINPUT29), .ZN(new_n422));
  NAND2_X1  g221(.A1(new_n410), .A2(new_n413), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n422), .A2(new_n423), .ZN(new_n424));
  AOI21_X1  g223(.A(new_n420), .B1(new_n421), .B2(new_n424), .ZN(new_n425));
  INV_X1    g224(.A(KEYINPUT30), .ZN(new_n426));
  XNOR2_X1  g225(.A(G8gat), .B(G36gat), .ZN(new_n427));
  XNOR2_X1  g226(.A(G64gat), .B(G92gat), .ZN(new_n428));
  XNOR2_X1  g227(.A(new_n427), .B(new_n428), .ZN(new_n429));
  INV_X1    g228(.A(new_n429), .ZN(new_n430));
  NAND3_X1  g229(.A1(new_n425), .A2(new_n426), .A3(new_n430), .ZN(new_n431));
  NAND2_X1  g230(.A1(new_n424), .A2(new_n421), .ZN(new_n432));
  NAND3_X1  g231(.A1(new_n432), .A2(new_n419), .A3(new_n430), .ZN(new_n433));
  NAND2_X1  g232(.A1(new_n433), .A2(KEYINPUT30), .ZN(new_n434));
  XOR2_X1   g233(.A(new_n429), .B(KEYINPUT75), .Z(new_n435));
  NOR2_X1   g234(.A1(new_n425), .A2(new_n435), .ZN(new_n436));
  OAI21_X1  g235(.A(new_n431), .B1(new_n434), .B2(new_n436), .ZN(new_n437));
  NAND2_X1  g236(.A1(new_n409), .A2(new_n437), .ZN(new_n438));
  OAI21_X1  g237(.A(KEYINPUT35), .B1(new_n367), .B2(new_n438), .ZN(new_n439));
  AND2_X1   g238(.A1(new_n282), .A2(new_n289), .ZN(new_n440));
  NAND2_X1  g239(.A1(new_n359), .A2(new_n293), .ZN(new_n441));
  AND2_X1   g240(.A1(new_n359), .A2(new_n363), .ZN(new_n442));
  OAI21_X1  g241(.A(new_n441), .B1(new_n442), .B2(new_n293), .ZN(new_n443));
  INV_X1    g242(.A(new_n403), .ZN(new_n444));
  NAND2_X1  g243(.A1(new_n406), .A2(new_n373), .ZN(new_n445));
  NAND3_X1  g244(.A1(new_n444), .A2(new_n445), .A3(new_n405), .ZN(new_n446));
  AND3_X1   g245(.A1(new_n403), .A2(KEYINPUT87), .A3(KEYINPUT6), .ZN(new_n447));
  AOI21_X1  g246(.A(KEYINPUT87), .B1(new_n403), .B2(KEYINPUT6), .ZN(new_n448));
  OAI21_X1  g247(.A(new_n446), .B1(new_n447), .B2(new_n448), .ZN(new_n449));
  AOI21_X1  g248(.A(new_n426), .B1(new_n425), .B2(new_n430), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n432), .A2(new_n419), .ZN(new_n451));
  INV_X1    g250(.A(new_n435), .ZN(new_n452));
  NAND2_X1  g251(.A1(new_n451), .A2(new_n452), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n450), .A2(new_n453), .ZN(new_n454));
  AOI21_X1  g253(.A(KEYINPUT35), .B1(new_n454), .B2(new_n431), .ZN(new_n455));
  NAND4_X1  g254(.A1(new_n440), .A2(new_n443), .A3(new_n449), .A4(new_n455), .ZN(new_n456));
  AND2_X1   g255(.A1(new_n439), .A2(new_n456), .ZN(new_n457));
  INV_X1    g256(.A(KEYINPUT39), .ZN(new_n458));
  INV_X1    g257(.A(KEYINPUT84), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n389), .A2(new_n390), .ZN(new_n460));
  AOI21_X1  g259(.A(new_n459), .B1(new_n460), .B2(new_n384), .ZN(new_n461));
  AOI211_X1 g260(.A(KEYINPUT84), .B(new_n383), .C1(new_n389), .C2(new_n390), .ZN(new_n462));
  OAI21_X1  g261(.A(new_n458), .B1(new_n461), .B2(new_n462), .ZN(new_n463));
  OAI21_X1  g262(.A(KEYINPUT84), .B1(new_n381), .B2(new_n383), .ZN(new_n464));
  NAND3_X1  g263(.A1(new_n460), .A2(new_n459), .A3(new_n384), .ZN(new_n465));
  AOI21_X1  g264(.A(new_n458), .B1(new_n394), .B2(new_n383), .ZN(new_n466));
  NAND3_X1  g265(.A1(new_n464), .A2(new_n465), .A3(new_n466), .ZN(new_n467));
  NAND3_X1  g266(.A1(new_n463), .A2(new_n467), .A3(new_n373), .ZN(new_n468));
  INV_X1    g267(.A(KEYINPUT40), .ZN(new_n469));
  NAND2_X1  g268(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  NAND4_X1  g269(.A1(new_n463), .A2(new_n467), .A3(KEYINPUT40), .A4(new_n373), .ZN(new_n471));
  NAND3_X1  g270(.A1(new_n470), .A2(new_n444), .A3(new_n471), .ZN(new_n472));
  OAI21_X1  g271(.A(KEYINPUT85), .B1(new_n472), .B2(new_n437), .ZN(new_n473));
  AND4_X1   g272(.A1(new_n426), .A2(new_n432), .A3(new_n419), .A4(new_n430), .ZN(new_n474));
  AOI21_X1  g273(.A(new_n474), .B1(new_n450), .B2(new_n453), .ZN(new_n475));
  INV_X1    g274(.A(KEYINPUT85), .ZN(new_n476));
  AOI21_X1  g275(.A(new_n403), .B1(new_n468), .B2(new_n469), .ZN(new_n477));
  NAND4_X1  g276(.A1(new_n475), .A2(new_n476), .A3(new_n471), .A4(new_n477), .ZN(new_n478));
  NAND2_X1  g277(.A1(new_n473), .A2(new_n478), .ZN(new_n479));
  INV_X1    g278(.A(KEYINPUT37), .ZN(new_n480));
  NOR2_X1   g279(.A1(new_n425), .A2(new_n480), .ZN(new_n481));
  NAND2_X1  g280(.A1(new_n260), .A2(new_n308), .ZN(new_n482));
  AOI22_X1  g281(.A1(new_n482), .A2(new_n418), .B1(new_n413), .B2(new_n410), .ZN(new_n483));
  OAI211_X1 g282(.A(new_n480), .B(new_n419), .C1(new_n483), .C2(new_n342), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n484), .A2(new_n429), .ZN(new_n485));
  OAI21_X1  g284(.A(KEYINPUT38), .B1(new_n481), .B2(new_n485), .ZN(new_n486));
  NAND2_X1  g285(.A1(new_n483), .A2(new_n342), .ZN(new_n487));
  OAI21_X1  g286(.A(new_n415), .B1(new_n417), .B2(new_n418), .ZN(new_n488));
  NAND2_X1  g287(.A1(new_n488), .A2(new_n338), .ZN(new_n489));
  NAND2_X1  g288(.A1(new_n487), .A2(new_n489), .ZN(new_n490));
  NAND2_X1  g289(.A1(new_n490), .A2(KEYINPUT37), .ZN(new_n491));
  INV_X1    g290(.A(KEYINPUT86), .ZN(new_n492));
  NOR2_X1   g291(.A1(new_n435), .A2(KEYINPUT38), .ZN(new_n493));
  NAND4_X1  g292(.A1(new_n491), .A2(new_n492), .A3(new_n484), .A4(new_n493), .ZN(new_n494));
  NAND2_X1  g293(.A1(new_n484), .A2(new_n493), .ZN(new_n495));
  AOI21_X1  g294(.A(new_n480), .B1(new_n487), .B2(new_n489), .ZN(new_n496));
  OAI21_X1  g295(.A(KEYINPUT86), .B1(new_n495), .B2(new_n496), .ZN(new_n497));
  NAND4_X1  g296(.A1(new_n486), .A2(new_n494), .A3(new_n497), .A4(new_n433), .ZN(new_n498));
  NOR2_X1   g297(.A1(new_n498), .A2(new_n449), .ZN(new_n499));
  OAI21_X1  g298(.A(new_n443), .B1(new_n479), .B2(new_n499), .ZN(new_n500));
  NOR2_X1   g299(.A1(new_n443), .A2(new_n438), .ZN(new_n501));
  INV_X1    g300(.A(new_n501), .ZN(new_n502));
  NAND2_X1  g301(.A1(new_n500), .A2(new_n502), .ZN(new_n503));
  NAND2_X1  g302(.A1(new_n282), .A2(new_n289), .ZN(new_n504));
  INV_X1    g303(.A(KEYINPUT36), .ZN(new_n505));
  NAND2_X1  g304(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  NAND3_X1  g305(.A1(new_n282), .A2(new_n289), .A3(KEYINPUT36), .ZN(new_n507));
  NAND2_X1  g306(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  AOI21_X1  g307(.A(new_n457), .B1(new_n503), .B2(new_n508), .ZN(new_n509));
  NAND2_X1  g308(.A1(KEYINPUT96), .A2(KEYINPUT18), .ZN(new_n510));
  NAND2_X1  g309(.A1(G229gat), .A2(G233gat), .ZN(new_n511));
  INV_X1    g310(.A(G8gat), .ZN(new_n512));
  XNOR2_X1  g311(.A(G15gat), .B(G22gat), .ZN(new_n513));
  AND2_X1   g312(.A1(new_n513), .A2(KEYINPUT93), .ZN(new_n514));
  NOR2_X1   g313(.A1(new_n513), .A2(KEYINPUT93), .ZN(new_n515));
  OR3_X1    g314(.A1(new_n514), .A2(new_n515), .A3(G1gat), .ZN(new_n516));
  AOI21_X1  g315(.A(new_n512), .B1(new_n516), .B2(KEYINPUT94), .ZN(new_n517));
  INV_X1    g316(.A(KEYINPUT16), .ZN(new_n518));
  OAI22_X1  g317(.A1(new_n514), .A2(new_n515), .B1(new_n518), .B2(G1gat), .ZN(new_n519));
  NAND2_X1  g318(.A1(new_n516), .A2(new_n519), .ZN(new_n520));
  OR2_X1    g319(.A1(new_n517), .A2(new_n520), .ZN(new_n521));
  NAND2_X1  g320(.A1(new_n517), .A2(new_n520), .ZN(new_n522));
  NAND2_X1  g321(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  NAND2_X1  g322(.A1(G29gat), .A2(G36gat), .ZN(new_n524));
  XNOR2_X1  g323(.A(new_n524), .B(KEYINPUT91), .ZN(new_n525));
  INV_X1    g324(.A(KEYINPUT14), .ZN(new_n526));
  INV_X1    g325(.A(G29gat), .ZN(new_n527));
  INV_X1    g326(.A(G36gat), .ZN(new_n528));
  NAND4_X1  g327(.A1(new_n526), .A2(new_n527), .A3(new_n528), .A4(KEYINPUT90), .ZN(new_n529));
  NAND3_X1  g328(.A1(new_n526), .A2(new_n527), .A3(new_n528), .ZN(new_n530));
  OAI21_X1  g329(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n531));
  NAND2_X1  g330(.A1(new_n530), .A2(new_n531), .ZN(new_n532));
  OAI211_X1 g331(.A(new_n525), .B(new_n529), .C1(KEYINPUT90), .C2(new_n532), .ZN(new_n533));
  XNOR2_X1  g332(.A(G43gat), .B(G50gat), .ZN(new_n534));
  INV_X1    g333(.A(KEYINPUT89), .ZN(new_n535));
  NAND3_X1  g334(.A1(new_n534), .A2(new_n535), .A3(KEYINPUT15), .ZN(new_n536));
  NAND2_X1  g335(.A1(new_n534), .A2(KEYINPUT15), .ZN(new_n537));
  INV_X1    g336(.A(KEYINPUT15), .ZN(new_n538));
  INV_X1    g337(.A(G43gat), .ZN(new_n539));
  NOR2_X1   g338(.A1(new_n539), .A2(G50gat), .ZN(new_n540));
  INV_X1    g339(.A(G50gat), .ZN(new_n541));
  NOR2_X1   g340(.A1(new_n541), .A2(G43gat), .ZN(new_n542));
  OAI21_X1  g341(.A(new_n538), .B1(new_n540), .B2(new_n542), .ZN(new_n543));
  NAND3_X1  g342(.A1(new_n537), .A2(new_n543), .A3(KEYINPUT89), .ZN(new_n544));
  AOI21_X1  g343(.A(new_n533), .B1(new_n536), .B2(new_n544), .ZN(new_n545));
  AOI21_X1  g344(.A(new_n537), .B1(new_n524), .B2(new_n532), .ZN(new_n546));
  OR2_X1    g345(.A1(new_n545), .A2(new_n546), .ZN(new_n547));
  NAND2_X1  g346(.A1(new_n523), .A2(new_n547), .ZN(new_n548));
  NOR2_X1   g347(.A1(new_n545), .A2(new_n546), .ZN(new_n549));
  OAI21_X1  g348(.A(KEYINPUT92), .B1(new_n549), .B2(KEYINPUT17), .ZN(new_n550));
  INV_X1    g349(.A(KEYINPUT92), .ZN(new_n551));
  INV_X1    g350(.A(KEYINPUT17), .ZN(new_n552));
  NAND3_X1  g351(.A1(new_n547), .A2(new_n551), .A3(new_n552), .ZN(new_n553));
  AND3_X1   g352(.A1(new_n549), .A2(KEYINPUT95), .A3(KEYINPUT17), .ZN(new_n554));
  AOI21_X1  g353(.A(KEYINPUT95), .B1(new_n549), .B2(KEYINPUT17), .ZN(new_n555));
  OAI211_X1 g354(.A(new_n550), .B(new_n553), .C1(new_n554), .C2(new_n555), .ZN(new_n556));
  OAI211_X1 g355(.A(new_n511), .B(new_n548), .C1(new_n556), .C2(new_n523), .ZN(new_n557));
  NOR2_X1   g356(.A1(KEYINPUT96), .A2(KEYINPUT18), .ZN(new_n558));
  OAI21_X1  g357(.A(new_n510), .B1(new_n557), .B2(new_n558), .ZN(new_n559));
  OR2_X1    g358(.A1(new_n556), .A2(new_n523), .ZN(new_n560));
  INV_X1    g359(.A(new_n510), .ZN(new_n561));
  NAND4_X1  g360(.A1(new_n560), .A2(new_n561), .A3(new_n511), .A4(new_n548), .ZN(new_n562));
  XNOR2_X1  g361(.A(new_n523), .B(new_n547), .ZN(new_n563));
  XOR2_X1   g362(.A(new_n511), .B(KEYINPUT13), .Z(new_n564));
  NAND2_X1  g363(.A1(new_n563), .A2(new_n564), .ZN(new_n565));
  NAND3_X1  g364(.A1(new_n559), .A2(new_n562), .A3(new_n565), .ZN(new_n566));
  XNOR2_X1  g365(.A(KEYINPUT88), .B(KEYINPUT11), .ZN(new_n567));
  XNOR2_X1  g366(.A(G113gat), .B(G141gat), .ZN(new_n568));
  XNOR2_X1  g367(.A(new_n567), .B(new_n568), .ZN(new_n569));
  XOR2_X1   g368(.A(G169gat), .B(G197gat), .Z(new_n570));
  XNOR2_X1  g369(.A(new_n569), .B(new_n570), .ZN(new_n571));
  XNOR2_X1  g370(.A(new_n571), .B(KEYINPUT12), .ZN(new_n572));
  INV_X1    g371(.A(new_n572), .ZN(new_n573));
  NAND2_X1  g372(.A1(new_n566), .A2(new_n573), .ZN(new_n574));
  NAND4_X1  g373(.A1(new_n559), .A2(new_n562), .A3(new_n572), .A4(new_n565), .ZN(new_n575));
  NAND2_X1  g374(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  INV_X1    g375(.A(new_n576), .ZN(new_n577));
  NOR2_X1   g376(.A1(new_n509), .A2(new_n577), .ZN(new_n578));
  INV_X1    g377(.A(KEYINPUT7), .ZN(new_n579));
  INV_X1    g378(.A(G85gat), .ZN(new_n580));
  INV_X1    g379(.A(G92gat), .ZN(new_n581));
  OAI21_X1  g380(.A(new_n579), .B1(new_n580), .B2(new_n581), .ZN(new_n582));
  NAND3_X1  g381(.A1(KEYINPUT7), .A2(G85gat), .A3(G92gat), .ZN(new_n583));
  OAI211_X1 g382(.A(new_n582), .B(new_n583), .C1(G85gat), .C2(G92gat), .ZN(new_n584));
  AND3_X1   g383(.A1(KEYINPUT101), .A2(G99gat), .A3(G106gat), .ZN(new_n585));
  AOI21_X1  g384(.A(KEYINPUT101), .B1(G99gat), .B2(G106gat), .ZN(new_n586));
  INV_X1    g385(.A(KEYINPUT8), .ZN(new_n587));
  NOR3_X1   g386(.A1(new_n585), .A2(new_n586), .A3(new_n587), .ZN(new_n588));
  XOR2_X1   g387(.A(G99gat), .B(G106gat), .Z(new_n589));
  OR3_X1    g388(.A1(new_n584), .A2(new_n588), .A3(new_n589), .ZN(new_n590));
  OAI21_X1  g389(.A(new_n589), .B1(new_n584), .B2(new_n588), .ZN(new_n591));
  AND2_X1   g390(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  NAND2_X1  g391(.A1(G232gat), .A2(G233gat), .ZN(new_n593));
  XOR2_X1   g392(.A(new_n593), .B(KEYINPUT100), .Z(new_n594));
  INV_X1    g393(.A(new_n594), .ZN(new_n595));
  AOI22_X1  g394(.A1(new_n547), .A2(new_n592), .B1(KEYINPUT41), .B2(new_n595), .ZN(new_n596));
  OAI21_X1  g395(.A(new_n596), .B1(new_n556), .B2(new_n592), .ZN(new_n597));
  XOR2_X1   g396(.A(G134gat), .B(G162gat), .Z(new_n598));
  NAND2_X1  g397(.A1(new_n597), .A2(new_n598), .ZN(new_n599));
  NOR2_X1   g398(.A1(new_n595), .A2(KEYINPUT41), .ZN(new_n600));
  XNOR2_X1  g399(.A(G190gat), .B(G218gat), .ZN(new_n601));
  XNOR2_X1  g400(.A(new_n600), .B(new_n601), .ZN(new_n602));
  INV_X1    g401(.A(new_n598), .ZN(new_n603));
  OAI211_X1 g402(.A(new_n603), .B(new_n596), .C1(new_n556), .C2(new_n592), .ZN(new_n604));
  AND3_X1   g403(.A1(new_n599), .A2(new_n602), .A3(new_n604), .ZN(new_n605));
  AOI21_X1  g404(.A(new_n602), .B1(new_n599), .B2(new_n604), .ZN(new_n606));
  NOR2_X1   g405(.A1(new_n605), .A2(new_n606), .ZN(new_n607));
  AOI21_X1  g406(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n608));
  OR2_X1    g407(.A1(new_n608), .A2(KEYINPUT97), .ZN(new_n609));
  XOR2_X1   g408(.A(G57gat), .B(G64gat), .Z(new_n610));
  NAND2_X1  g409(.A1(new_n608), .A2(KEYINPUT97), .ZN(new_n611));
  NAND3_X1  g410(.A1(new_n609), .A2(new_n610), .A3(new_n611), .ZN(new_n612));
  XNOR2_X1  g411(.A(G71gat), .B(G78gat), .ZN(new_n613));
  XNOR2_X1  g412(.A(new_n612), .B(new_n613), .ZN(new_n614));
  NAND2_X1  g413(.A1(new_n614), .A2(KEYINPUT21), .ZN(new_n615));
  NAND3_X1  g414(.A1(new_n521), .A2(new_n522), .A3(new_n615), .ZN(new_n616));
  XOR2_X1   g415(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n617));
  INV_X1    g416(.A(new_n617), .ZN(new_n618));
  XNOR2_X1  g417(.A(new_n616), .B(new_n618), .ZN(new_n619));
  XOR2_X1   g418(.A(new_n612), .B(new_n613), .Z(new_n620));
  INV_X1    g419(.A(G127gat), .ZN(new_n621));
  XNOR2_X1  g420(.A(KEYINPUT98), .B(KEYINPUT21), .ZN(new_n622));
  NAND3_X1  g421(.A1(new_n620), .A2(new_n621), .A3(new_n622), .ZN(new_n623));
  INV_X1    g422(.A(new_n623), .ZN(new_n624));
  AOI21_X1  g423(.A(new_n621), .B1(new_n620), .B2(new_n622), .ZN(new_n625));
  OAI21_X1  g424(.A(G155gat), .B1(new_n624), .B2(new_n625), .ZN(new_n626));
  INV_X1    g425(.A(new_n625), .ZN(new_n627));
  INV_X1    g426(.A(G155gat), .ZN(new_n628));
  NAND3_X1  g427(.A1(new_n627), .A2(new_n628), .A3(new_n623), .ZN(new_n629));
  NAND2_X1  g428(.A1(new_n626), .A2(new_n629), .ZN(new_n630));
  NAND2_X1  g429(.A1(G231gat), .A2(G233gat), .ZN(new_n631));
  XNOR2_X1  g430(.A(new_n631), .B(KEYINPUT99), .ZN(new_n632));
  XNOR2_X1  g431(.A(new_n632), .B(new_n236), .ZN(new_n633));
  XNOR2_X1  g432(.A(new_n633), .B(G211gat), .ZN(new_n634));
  INV_X1    g433(.A(new_n634), .ZN(new_n635));
  NAND2_X1  g434(.A1(new_n630), .A2(new_n635), .ZN(new_n636));
  NAND3_X1  g435(.A1(new_n626), .A2(new_n629), .A3(new_n634), .ZN(new_n637));
  AND3_X1   g436(.A1(new_n619), .A2(new_n636), .A3(new_n637), .ZN(new_n638));
  AOI21_X1  g437(.A(new_n619), .B1(new_n636), .B2(new_n637), .ZN(new_n639));
  OR2_X1    g438(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  OAI21_X1  g439(.A(KEYINPUT102), .B1(new_n607), .B2(new_n640), .ZN(new_n641));
  NOR2_X1   g440(.A1(new_n638), .A2(new_n639), .ZN(new_n642));
  INV_X1    g441(.A(KEYINPUT102), .ZN(new_n643));
  OAI211_X1 g442(.A(new_n642), .B(new_n643), .C1(new_n605), .C2(new_n606), .ZN(new_n644));
  NAND2_X1  g443(.A1(new_n641), .A2(new_n644), .ZN(new_n645));
  INV_X1    g444(.A(G230gat), .ZN(new_n646));
  NOR2_X1   g445(.A1(new_n646), .A2(new_n295), .ZN(new_n647));
  INV_X1    g446(.A(new_n647), .ZN(new_n648));
  NAND2_X1  g447(.A1(new_n590), .A2(new_n591), .ZN(new_n649));
  NAND2_X1  g448(.A1(new_n620), .A2(new_n649), .ZN(new_n650));
  NAND3_X1  g449(.A1(new_n614), .A2(new_n590), .A3(new_n591), .ZN(new_n651));
  NAND3_X1  g450(.A1(new_n650), .A2(KEYINPUT103), .A3(new_n651), .ZN(new_n652));
  OR3_X1    g451(.A1(new_n592), .A2(KEYINPUT103), .A3(new_n614), .ZN(new_n653));
  AOI21_X1  g452(.A(KEYINPUT10), .B1(new_n652), .B2(new_n653), .ZN(new_n654));
  NAND3_X1  g453(.A1(new_n592), .A2(KEYINPUT10), .A3(new_n614), .ZN(new_n655));
  INV_X1    g454(.A(new_n655), .ZN(new_n656));
  OAI21_X1  g455(.A(new_n648), .B1(new_n654), .B2(new_n656), .ZN(new_n657));
  AND2_X1   g456(.A1(new_n652), .A2(new_n653), .ZN(new_n658));
  NAND2_X1  g457(.A1(new_n658), .A2(new_n647), .ZN(new_n659));
  NAND2_X1  g458(.A1(new_n657), .A2(new_n659), .ZN(new_n660));
  XNOR2_X1  g459(.A(G120gat), .B(G148gat), .ZN(new_n661));
  XNOR2_X1  g460(.A(G176gat), .B(G204gat), .ZN(new_n662));
  XNOR2_X1  g461(.A(new_n661), .B(new_n662), .ZN(new_n663));
  NAND2_X1  g462(.A1(new_n660), .A2(new_n663), .ZN(new_n664));
  INV_X1    g463(.A(new_n663), .ZN(new_n665));
  NAND3_X1  g464(.A1(new_n657), .A2(new_n659), .A3(new_n665), .ZN(new_n666));
  NAND2_X1  g465(.A1(new_n664), .A2(new_n666), .ZN(new_n667));
  INV_X1    g466(.A(KEYINPUT104), .ZN(new_n668));
  NAND2_X1  g467(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  NAND3_X1  g468(.A1(new_n664), .A2(KEYINPUT104), .A3(new_n666), .ZN(new_n670));
  NAND2_X1  g469(.A1(new_n669), .A2(new_n670), .ZN(new_n671));
  NOR2_X1   g470(.A1(new_n645), .A2(new_n671), .ZN(new_n672));
  NAND2_X1  g471(.A1(new_n578), .A2(new_n672), .ZN(new_n673));
  NOR2_X1   g472(.A1(new_n673), .A2(new_n409), .ZN(new_n674));
  XNOR2_X1  g473(.A(KEYINPUT105), .B(G1gat), .ZN(new_n675));
  XNOR2_X1  g474(.A(new_n674), .B(new_n675), .ZN(G1324gat));
  INV_X1    g475(.A(KEYINPUT106), .ZN(new_n677));
  INV_X1    g476(.A(new_n673), .ZN(new_n678));
  NAND2_X1  g477(.A1(new_n678), .A2(new_n475), .ZN(new_n679));
  XNOR2_X1  g478(.A(KEYINPUT16), .B(G8gat), .ZN(new_n680));
  NOR2_X1   g479(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  AOI21_X1  g480(.A(new_n677), .B1(new_n681), .B2(KEYINPUT42), .ZN(new_n682));
  INV_X1    g481(.A(KEYINPUT42), .ZN(new_n683));
  NOR4_X1   g482(.A1(new_n679), .A2(KEYINPUT106), .A3(new_n683), .A4(new_n680), .ZN(new_n684));
  AOI21_X1  g483(.A(new_n683), .B1(new_n679), .B2(G8gat), .ZN(new_n685));
  OAI22_X1  g484(.A1(new_n682), .A2(new_n684), .B1(new_n685), .B2(new_n681), .ZN(G1325gat));
  AND3_X1   g485(.A1(new_n282), .A2(new_n289), .A3(KEYINPUT36), .ZN(new_n687));
  AOI21_X1  g486(.A(KEYINPUT36), .B1(new_n282), .B2(new_n289), .ZN(new_n688));
  OAI21_X1  g487(.A(KEYINPUT107), .B1(new_n687), .B2(new_n688), .ZN(new_n689));
  INV_X1    g488(.A(KEYINPUT107), .ZN(new_n690));
  NAND3_X1  g489(.A1(new_n506), .A2(new_n690), .A3(new_n507), .ZN(new_n691));
  AND2_X1   g490(.A1(new_n689), .A2(new_n691), .ZN(new_n692));
  AND3_X1   g491(.A1(new_n678), .A2(G15gat), .A3(new_n692), .ZN(new_n693));
  AOI21_X1  g492(.A(G15gat), .B1(new_n678), .B2(new_n440), .ZN(new_n694));
  NOR2_X1   g493(.A1(new_n693), .A2(new_n694), .ZN(G1326gat));
  INV_X1    g494(.A(new_n443), .ZN(new_n696));
  NAND3_X1  g495(.A1(new_n678), .A2(new_n344), .A3(new_n696), .ZN(new_n697));
  OAI21_X1  g496(.A(G22gat), .B1(new_n673), .B2(new_n443), .ZN(new_n698));
  NAND2_X1  g497(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  XNOR2_X1  g498(.A(KEYINPUT108), .B(KEYINPUT43), .ZN(new_n700));
  XNOR2_X1  g499(.A(new_n699), .B(new_n700), .ZN(G1327gat));
  INV_X1    g500(.A(new_n671), .ZN(new_n702));
  NAND2_X1  g501(.A1(new_n702), .A2(new_n640), .ZN(new_n703));
  INV_X1    g502(.A(new_n607), .ZN(new_n704));
  NOR2_X1   g503(.A1(new_n703), .A2(new_n704), .ZN(new_n705));
  XNOR2_X1  g504(.A(new_n705), .B(KEYINPUT109), .ZN(new_n706));
  NAND2_X1  g505(.A1(new_n578), .A2(new_n706), .ZN(new_n707));
  NOR3_X1   g506(.A1(new_n707), .A2(G29gat), .A3(new_n409), .ZN(new_n708));
  XOR2_X1   g507(.A(new_n708), .B(KEYINPUT45), .Z(new_n709));
  INV_X1    g508(.A(KEYINPUT112), .ZN(new_n710));
  OAI21_X1  g509(.A(KEYINPUT44), .B1(new_n509), .B2(new_n704), .ZN(new_n711));
  OAI211_X1 g510(.A(new_n473), .B(new_n478), .C1(new_n449), .C2(new_n498), .ZN(new_n712));
  AOI21_X1  g511(.A(new_n501), .B1(new_n712), .B2(new_n443), .ZN(new_n713));
  AND3_X1   g512(.A1(new_n439), .A2(new_n456), .A3(KEYINPUT110), .ZN(new_n714));
  AOI21_X1  g513(.A(KEYINPUT110), .B1(new_n439), .B2(new_n456), .ZN(new_n715));
  OAI22_X1  g514(.A1(new_n713), .A2(new_n692), .B1(new_n714), .B2(new_n715), .ZN(new_n716));
  XOR2_X1   g515(.A(KEYINPUT111), .B(KEYINPUT44), .Z(new_n717));
  NAND3_X1  g516(.A1(new_n716), .A2(new_n607), .A3(new_n717), .ZN(new_n718));
  NAND2_X1  g517(.A1(new_n711), .A2(new_n718), .ZN(new_n719));
  NOR2_X1   g518(.A1(new_n703), .A2(new_n577), .ZN(new_n720));
  AOI21_X1  g519(.A(new_n710), .B1(new_n719), .B2(new_n720), .ZN(new_n721));
  INV_X1    g520(.A(new_n721), .ZN(new_n722));
  INV_X1    g521(.A(new_n720), .ZN(new_n723));
  AOI211_X1 g522(.A(KEYINPUT112), .B(new_n723), .C1(new_n711), .C2(new_n718), .ZN(new_n724));
  INV_X1    g523(.A(new_n724), .ZN(new_n725));
  AOI21_X1  g524(.A(new_n409), .B1(new_n722), .B2(new_n725), .ZN(new_n726));
  OAI21_X1  g525(.A(new_n709), .B1(new_n726), .B2(new_n527), .ZN(G1328gat));
  NOR3_X1   g526(.A1(new_n707), .A2(G36gat), .A3(new_n437), .ZN(new_n728));
  XNOR2_X1  g527(.A(new_n728), .B(KEYINPUT46), .ZN(new_n729));
  AOI21_X1  g528(.A(new_n437), .B1(new_n722), .B2(new_n725), .ZN(new_n730));
  OAI21_X1  g529(.A(new_n729), .B1(new_n730), .B2(new_n528), .ZN(G1329gat));
  NOR3_X1   g530(.A1(new_n707), .A2(G43gat), .A3(new_n504), .ZN(new_n732));
  INV_X1    g531(.A(KEYINPUT47), .ZN(new_n733));
  NOR2_X1   g532(.A1(new_n732), .A2(new_n733), .ZN(new_n734));
  INV_X1    g533(.A(new_n719), .ZN(new_n735));
  INV_X1    g534(.A(new_n692), .ZN(new_n736));
  NOR3_X1   g535(.A1(new_n735), .A2(new_n736), .A3(new_n723), .ZN(new_n737));
  OAI21_X1  g536(.A(new_n734), .B1(new_n737), .B2(new_n539), .ZN(new_n738));
  OAI21_X1  g537(.A(new_n692), .B1(new_n721), .B2(new_n724), .ZN(new_n739));
  AOI21_X1  g538(.A(new_n732), .B1(new_n739), .B2(G43gat), .ZN(new_n740));
  OAI21_X1  g539(.A(new_n738), .B1(new_n740), .B2(KEYINPUT47), .ZN(G1330gat));
  NOR3_X1   g540(.A1(new_n707), .A2(G50gat), .A3(new_n443), .ZN(new_n742));
  INV_X1    g541(.A(KEYINPUT48), .ZN(new_n743));
  NOR2_X1   g542(.A1(new_n742), .A2(new_n743), .ZN(new_n744));
  NOR3_X1   g543(.A1(new_n735), .A2(new_n443), .A3(new_n723), .ZN(new_n745));
  OAI21_X1  g544(.A(new_n744), .B1(new_n745), .B2(new_n541), .ZN(new_n746));
  OAI21_X1  g545(.A(new_n696), .B1(new_n721), .B2(new_n724), .ZN(new_n747));
  AOI21_X1  g546(.A(new_n742), .B1(new_n747), .B2(G50gat), .ZN(new_n748));
  OAI21_X1  g547(.A(new_n746), .B1(new_n748), .B2(KEYINPUT48), .ZN(G1331gat));
  NOR3_X1   g548(.A1(new_n645), .A2(new_n576), .A3(new_n702), .ZN(new_n750));
  AND2_X1   g549(.A1(new_n716), .A2(new_n750), .ZN(new_n751));
  INV_X1    g550(.A(new_n409), .ZN(new_n752));
  NAND2_X1  g551(.A1(new_n751), .A2(new_n752), .ZN(new_n753));
  XNOR2_X1  g552(.A(new_n753), .B(G57gat), .ZN(G1332gat));
  NAND2_X1  g553(.A1(new_n751), .A2(new_n475), .ZN(new_n755));
  OAI21_X1  g554(.A(new_n755), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n756));
  XOR2_X1   g555(.A(KEYINPUT49), .B(G64gat), .Z(new_n757));
  OAI21_X1  g556(.A(new_n756), .B1(new_n755), .B2(new_n757), .ZN(new_n758));
  XNOR2_X1  g557(.A(KEYINPUT113), .B(KEYINPUT114), .ZN(new_n759));
  XNOR2_X1  g558(.A(new_n758), .B(new_n759), .ZN(G1333gat));
  AOI21_X1  g559(.A(G71gat), .B1(new_n751), .B2(new_n440), .ZN(new_n761));
  AND2_X1   g560(.A1(new_n692), .A2(G71gat), .ZN(new_n762));
  AOI21_X1  g561(.A(new_n761), .B1(new_n751), .B2(new_n762), .ZN(new_n763));
  XOR2_X1   g562(.A(new_n763), .B(KEYINPUT50), .Z(G1334gat));
  NAND2_X1  g563(.A1(new_n751), .A2(new_n696), .ZN(new_n765));
  XNOR2_X1  g564(.A(new_n765), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g565(.A1(new_n576), .A2(new_n642), .ZN(new_n767));
  NAND3_X1  g566(.A1(new_n719), .A2(new_n671), .A3(new_n767), .ZN(new_n768));
  OAI21_X1  g567(.A(G85gat), .B1(new_n768), .B2(new_n409), .ZN(new_n769));
  AND2_X1   g568(.A1(new_n716), .A2(new_n607), .ZN(new_n770));
  AOI21_X1  g569(.A(KEYINPUT51), .B1(new_n770), .B2(new_n767), .ZN(new_n771));
  INV_X1    g570(.A(new_n771), .ZN(new_n772));
  NAND3_X1  g571(.A1(new_n770), .A2(KEYINPUT51), .A3(new_n767), .ZN(new_n773));
  NAND2_X1  g572(.A1(new_n772), .A2(new_n773), .ZN(new_n774));
  INV_X1    g573(.A(new_n774), .ZN(new_n775));
  NAND3_X1  g574(.A1(new_n671), .A2(new_n752), .A3(new_n580), .ZN(new_n776));
  OAI21_X1  g575(.A(new_n769), .B1(new_n775), .B2(new_n776), .ZN(G1336gat));
  INV_X1    g576(.A(KEYINPUT115), .ZN(new_n778));
  NOR3_X1   g577(.A1(new_n702), .A2(G92gat), .A3(new_n437), .ZN(new_n779));
  INV_X1    g578(.A(new_n773), .ZN(new_n780));
  OAI211_X1 g579(.A(new_n778), .B(new_n779), .C1(new_n780), .C2(new_n771), .ZN(new_n781));
  OAI21_X1  g580(.A(G92gat), .B1(new_n768), .B2(new_n437), .ZN(new_n782));
  INV_X1    g581(.A(KEYINPUT116), .ZN(new_n783));
  NAND3_X1  g582(.A1(new_n781), .A2(new_n782), .A3(new_n783), .ZN(new_n784));
  INV_X1    g583(.A(KEYINPUT52), .ZN(new_n785));
  AOI21_X1  g584(.A(KEYINPUT115), .B1(new_n783), .B2(KEYINPUT52), .ZN(new_n786));
  AOI21_X1  g585(.A(new_n786), .B1(new_n774), .B2(new_n779), .ZN(new_n787));
  AOI22_X1  g586(.A1(new_n784), .A2(new_n785), .B1(new_n787), .B2(new_n782), .ZN(G1337gat));
  OAI21_X1  g587(.A(G99gat), .B1(new_n768), .B2(new_n736), .ZN(new_n789));
  OR3_X1    g588(.A1(new_n702), .A2(G99gat), .A3(new_n504), .ZN(new_n790));
  OAI21_X1  g589(.A(new_n789), .B1(new_n775), .B2(new_n790), .ZN(G1338gat));
  OAI21_X1  g590(.A(G106gat), .B1(new_n768), .B2(new_n443), .ZN(new_n792));
  INV_X1    g591(.A(new_n792), .ZN(new_n793));
  NOR3_X1   g592(.A1(new_n702), .A2(G106gat), .A3(new_n443), .ZN(new_n794));
  XOR2_X1   g593(.A(new_n794), .B(KEYINPUT117), .Z(new_n795));
  INV_X1    g594(.A(new_n795), .ZN(new_n796));
  AOI21_X1  g595(.A(new_n796), .B1(new_n772), .B2(new_n773), .ZN(new_n797));
  OAI21_X1  g596(.A(KEYINPUT53), .B1(new_n793), .B2(new_n797), .ZN(new_n798));
  INV_X1    g597(.A(KEYINPUT53), .ZN(new_n799));
  OAI211_X1 g598(.A(new_n792), .B(new_n799), .C1(new_n775), .C2(new_n796), .ZN(new_n800));
  NAND2_X1  g599(.A1(new_n798), .A2(new_n800), .ZN(G1339gat));
  OAI211_X1 g600(.A(new_n647), .B(new_n655), .C1(new_n658), .C2(KEYINPUT10), .ZN(new_n802));
  NAND3_X1  g601(.A1(new_n802), .A2(new_n657), .A3(KEYINPUT54), .ZN(new_n803));
  INV_X1    g602(.A(KEYINPUT54), .ZN(new_n804));
  OAI211_X1 g603(.A(new_n804), .B(new_n648), .C1(new_n654), .C2(new_n656), .ZN(new_n805));
  INV_X1    g604(.A(KEYINPUT118), .ZN(new_n806));
  AND3_X1   g605(.A1(new_n805), .A2(new_n806), .A3(new_n663), .ZN(new_n807));
  AOI21_X1  g606(.A(new_n806), .B1(new_n805), .B2(new_n663), .ZN(new_n808));
  OAI21_X1  g607(.A(new_n803), .B1(new_n807), .B2(new_n808), .ZN(new_n809));
  INV_X1    g608(.A(KEYINPUT55), .ZN(new_n810));
  NAND2_X1  g609(.A1(new_n809), .A2(new_n810), .ZN(new_n811));
  OAI211_X1 g610(.A(KEYINPUT55), .B(new_n803), .C1(new_n807), .C2(new_n808), .ZN(new_n812));
  NAND4_X1  g611(.A1(new_n576), .A2(new_n666), .A3(new_n811), .A4(new_n812), .ZN(new_n813));
  AOI21_X1  g612(.A(new_n511), .B1(new_n560), .B2(new_n548), .ZN(new_n814));
  NOR2_X1   g613(.A1(new_n563), .A2(new_n564), .ZN(new_n815));
  OAI21_X1  g614(.A(new_n571), .B1(new_n814), .B2(new_n815), .ZN(new_n816));
  AND2_X1   g615(.A1(new_n575), .A2(new_n816), .ZN(new_n817));
  AOI21_X1  g616(.A(new_n607), .B1(new_n817), .B2(new_n671), .ZN(new_n818));
  NAND2_X1  g617(.A1(new_n813), .A2(new_n818), .ZN(new_n819));
  NAND3_X1  g618(.A1(new_n811), .A2(new_n666), .A3(new_n812), .ZN(new_n820));
  NAND2_X1  g619(.A1(new_n575), .A2(new_n816), .ZN(new_n821));
  OAI21_X1  g620(.A(new_n607), .B1(new_n820), .B2(new_n821), .ZN(new_n822));
  NAND3_X1  g621(.A1(new_n819), .A2(new_n640), .A3(new_n822), .ZN(new_n823));
  AND4_X1   g622(.A1(new_n577), .A2(new_n641), .A3(new_n702), .A4(new_n644), .ZN(new_n824));
  INV_X1    g623(.A(new_n824), .ZN(new_n825));
  NAND2_X1  g624(.A1(new_n823), .A2(new_n825), .ZN(new_n826));
  NOR3_X1   g625(.A1(new_n367), .A2(new_n409), .A3(new_n475), .ZN(new_n827));
  NAND2_X1  g626(.A1(new_n826), .A2(new_n827), .ZN(new_n828));
  NOR2_X1   g627(.A1(new_n828), .A2(new_n577), .ZN(new_n829));
  XOR2_X1   g628(.A(new_n829), .B(G113gat), .Z(G1340gat));
  NOR2_X1   g629(.A1(new_n828), .A2(new_n702), .ZN(new_n831));
  INV_X1    g630(.A(G120gat), .ZN(new_n832));
  OAI21_X1  g631(.A(new_n831), .B1(KEYINPUT119), .B2(new_n832), .ZN(new_n833));
  XNOR2_X1  g632(.A(KEYINPUT119), .B(G120gat), .ZN(new_n834));
  OAI21_X1  g633(.A(new_n833), .B1(new_n831), .B2(new_n834), .ZN(G1341gat));
  NOR2_X1   g634(.A1(new_n828), .A2(new_n640), .ZN(new_n836));
  XNOR2_X1  g635(.A(new_n836), .B(new_n621), .ZN(G1342gat));
  NOR3_X1   g636(.A1(new_n828), .A2(G134gat), .A3(new_n704), .ZN(new_n838));
  XNOR2_X1  g637(.A(new_n838), .B(KEYINPUT120), .ZN(new_n839));
  NAND3_X1  g638(.A1(new_n826), .A2(new_n607), .A3(new_n827), .ZN(new_n840));
  AOI22_X1  g639(.A1(new_n839), .A2(KEYINPUT56), .B1(G134gat), .B2(new_n840), .ZN(new_n841));
  OAI21_X1  g640(.A(new_n841), .B1(KEYINPUT56), .B2(new_n839), .ZN(G1343gat));
  INV_X1    g641(.A(KEYINPUT57), .ZN(new_n843));
  AOI21_X1  g642(.A(new_n642), .B1(new_n813), .B2(new_n818), .ZN(new_n844));
  AOI21_X1  g643(.A(new_n824), .B1(new_n844), .B2(new_n822), .ZN(new_n845));
  OAI21_X1  g644(.A(new_n843), .B1(new_n845), .B2(new_n443), .ZN(new_n846));
  NAND3_X1  g645(.A1(new_n826), .A2(KEYINPUT57), .A3(new_n696), .ZN(new_n847));
  NAND2_X1  g646(.A1(new_n846), .A2(new_n847), .ZN(new_n848));
  AOI211_X1 g647(.A(new_n409), .B(new_n475), .C1(new_n689), .C2(new_n691), .ZN(new_n849));
  XNOR2_X1  g648(.A(new_n849), .B(KEYINPUT121), .ZN(new_n850));
  NAND2_X1  g649(.A1(new_n848), .A2(new_n850), .ZN(new_n851));
  OAI21_X1  g650(.A(G141gat), .B1(new_n851), .B2(new_n577), .ZN(new_n852));
  NOR2_X1   g651(.A1(new_n845), .A2(new_n443), .ZN(new_n853));
  AND2_X1   g652(.A1(new_n853), .A2(new_n849), .ZN(new_n854));
  NAND3_X1  g653(.A1(new_n854), .A2(new_n321), .A3(new_n576), .ZN(new_n855));
  NAND2_X1  g654(.A1(new_n852), .A2(new_n855), .ZN(new_n856));
  XNOR2_X1  g655(.A(new_n856), .B(KEYINPUT58), .ZN(G1344gat));
  NAND3_X1  g656(.A1(new_n854), .A2(new_n323), .A3(new_n671), .ZN(new_n858));
  NAND3_X1  g657(.A1(new_n848), .A2(new_n671), .A3(new_n850), .ZN(new_n859));
  INV_X1    g658(.A(KEYINPUT59), .ZN(new_n860));
  AND3_X1   g659(.A1(new_n859), .A2(new_n860), .A3(G148gat), .ZN(new_n861));
  AOI21_X1  g660(.A(new_n860), .B1(new_n859), .B2(G148gat), .ZN(new_n862));
  OAI21_X1  g661(.A(new_n858), .B1(new_n861), .B2(new_n862), .ZN(new_n863));
  NAND2_X1  g662(.A1(new_n863), .A2(KEYINPUT122), .ZN(new_n864));
  INV_X1    g663(.A(KEYINPUT122), .ZN(new_n865));
  OAI211_X1 g664(.A(new_n865), .B(new_n858), .C1(new_n861), .C2(new_n862), .ZN(new_n866));
  NAND2_X1  g665(.A1(new_n864), .A2(new_n866), .ZN(G1345gat));
  NOR3_X1   g666(.A1(new_n851), .A2(new_n628), .A3(new_n640), .ZN(new_n868));
  AOI21_X1  g667(.A(G155gat), .B1(new_n854), .B2(new_n642), .ZN(new_n869));
  NOR2_X1   g668(.A1(new_n868), .A2(new_n869), .ZN(G1346gat));
  AND2_X1   g669(.A1(new_n854), .A2(new_n607), .ZN(new_n871));
  NAND2_X1  g670(.A1(new_n607), .A2(G162gat), .ZN(new_n872));
  OAI22_X1  g671(.A1(new_n871), .A2(G162gat), .B1(new_n851), .B2(new_n872), .ZN(new_n873));
  XNOR2_X1  g672(.A(new_n873), .B(KEYINPUT123), .ZN(G1347gat));
  NOR2_X1   g673(.A1(new_n845), .A2(new_n752), .ZN(new_n875));
  NOR2_X1   g674(.A1(new_n367), .A2(new_n437), .ZN(new_n876));
  NAND2_X1  g675(.A1(new_n875), .A2(new_n876), .ZN(new_n877));
  OAI21_X1  g676(.A(G169gat), .B1(new_n877), .B2(new_n577), .ZN(new_n878));
  XNOR2_X1  g677(.A(new_n876), .B(KEYINPUT124), .ZN(new_n879));
  NAND2_X1  g678(.A1(new_n875), .A2(new_n879), .ZN(new_n880));
  NAND2_X1  g679(.A1(new_n576), .A2(new_n223), .ZN(new_n881));
  OAI21_X1  g680(.A(new_n878), .B1(new_n880), .B2(new_n881), .ZN(G1348gat));
  NOR3_X1   g681(.A1(new_n877), .A2(new_n224), .A3(new_n702), .ZN(new_n883));
  NAND3_X1  g682(.A1(new_n875), .A2(new_n671), .A3(new_n879), .ZN(new_n884));
  AOI21_X1  g683(.A(new_n883), .B1(new_n224), .B2(new_n884), .ZN(G1349gat));
  NAND4_X1  g684(.A1(new_n875), .A2(new_n214), .A3(new_n642), .A4(new_n879), .ZN(new_n886));
  XOR2_X1   g685(.A(new_n886), .B(KEYINPUT125), .Z(new_n887));
  OAI21_X1  g686(.A(G183gat), .B1(new_n877), .B2(new_n640), .ZN(new_n888));
  NAND2_X1  g687(.A1(new_n887), .A2(new_n888), .ZN(new_n889));
  NAND2_X1  g688(.A1(new_n889), .A2(KEYINPUT60), .ZN(new_n890));
  INV_X1    g689(.A(KEYINPUT60), .ZN(new_n891));
  NAND3_X1  g690(.A1(new_n887), .A2(new_n891), .A3(new_n888), .ZN(new_n892));
  NAND2_X1  g691(.A1(new_n890), .A2(new_n892), .ZN(G1350gat));
  OAI21_X1  g692(.A(G190gat), .B1(new_n877), .B2(new_n704), .ZN(new_n894));
  NAND3_X1  g693(.A1(new_n894), .A2(KEYINPUT126), .A3(KEYINPUT61), .ZN(new_n895));
  OAI21_X1  g694(.A(new_n895), .B1(KEYINPUT61), .B2(new_n894), .ZN(new_n896));
  AOI21_X1  g695(.A(KEYINPUT126), .B1(new_n894), .B2(KEYINPUT61), .ZN(new_n897));
  NAND2_X1  g696(.A1(new_n607), .A2(new_n215), .ZN(new_n898));
  OAI22_X1  g697(.A1(new_n896), .A2(new_n897), .B1(new_n880), .B2(new_n898), .ZN(G1351gat));
  NOR3_X1   g698(.A1(new_n692), .A2(new_n752), .A3(new_n437), .ZN(new_n900));
  NAND2_X1  g699(.A1(new_n853), .A2(new_n900), .ZN(new_n901));
  OR3_X1    g700(.A1(new_n901), .A2(G197gat), .A3(new_n577), .ZN(new_n902));
  NAND2_X1  g701(.A1(new_n848), .A2(new_n900), .ZN(new_n903));
  INV_X1    g702(.A(new_n903), .ZN(new_n904));
  NAND2_X1  g703(.A1(new_n904), .A2(new_n576), .ZN(new_n905));
  AND2_X1   g704(.A1(new_n905), .A2(KEYINPUT127), .ZN(new_n906));
  OAI21_X1  g705(.A(G197gat), .B1(new_n905), .B2(KEYINPUT127), .ZN(new_n907));
  OAI21_X1  g706(.A(new_n902), .B1(new_n906), .B2(new_n907), .ZN(G1352gat));
  NOR3_X1   g707(.A1(new_n901), .A2(G204gat), .A3(new_n702), .ZN(new_n909));
  XNOR2_X1  g708(.A(new_n909), .B(KEYINPUT62), .ZN(new_n910));
  OAI21_X1  g709(.A(G204gat), .B1(new_n903), .B2(new_n702), .ZN(new_n911));
  NAND2_X1  g710(.A1(new_n910), .A2(new_n911), .ZN(G1353gat));
  NAND2_X1  g711(.A1(new_n904), .A2(new_n642), .ZN(new_n913));
  AND3_X1   g712(.A1(new_n913), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n914));
  AOI21_X1  g713(.A(KEYINPUT63), .B1(new_n913), .B2(G211gat), .ZN(new_n915));
  OR2_X1    g714(.A1(new_n640), .A2(G211gat), .ZN(new_n916));
  OAI22_X1  g715(.A1(new_n914), .A2(new_n915), .B1(new_n901), .B2(new_n916), .ZN(G1354gat));
  INV_X1    g716(.A(G218gat), .ZN(new_n918));
  NOR3_X1   g717(.A1(new_n903), .A2(new_n918), .A3(new_n704), .ZN(new_n919));
  NAND3_X1  g718(.A1(new_n853), .A2(new_n607), .A3(new_n900), .ZN(new_n920));
  AOI21_X1  g719(.A(new_n919), .B1(new_n918), .B2(new_n920), .ZN(G1355gat));
endmodule


