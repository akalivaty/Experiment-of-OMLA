//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 1 1 0 0 1 1 1 0 0 0 0 1 0 0 1 1 0 1 1 1 1 0 1 1 0 0 0 1 1 1 1 1 0 1 0 1 0 0 0 1 0 0 0 1 1 0 0 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:27:14 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n614, new_n615,
    new_n616, new_n617, new_n618, new_n619, new_n620, new_n621, new_n622,
    new_n623, new_n625, new_n626, new_n627, new_n628, new_n629, new_n630,
    new_n631, new_n632, new_n633, new_n634, new_n635, new_n636, new_n637,
    new_n638, new_n639, new_n640, new_n641, new_n643, new_n644, new_n645,
    new_n646, new_n647, new_n648, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n671, new_n672, new_n673, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n682, new_n684, new_n685,
    new_n686, new_n687, new_n688, new_n689, new_n690, new_n692, new_n693,
    new_n694, new_n695, new_n696, new_n697, new_n698, new_n699, new_n700,
    new_n701, new_n702, new_n703, new_n704, new_n705, new_n707, new_n708,
    new_n709, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n731,
    new_n732, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n896, new_n897, new_n898,
    new_n900, new_n901, new_n902, new_n903, new_n904, new_n905, new_n906,
    new_n907, new_n908, new_n909, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n922,
    new_n923, new_n924, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n961, new_n962, new_n963, new_n964, new_n965, new_n966,
    new_n967, new_n968, new_n969;
  INV_X1    g000(.A(G146), .ZN(new_n187));
  INV_X1    g001(.A(KEYINPUT16), .ZN(new_n188));
  OR2_X1    g002(.A1(KEYINPUT75), .A2(G125), .ZN(new_n189));
  NAND2_X1  g003(.A1(KEYINPUT75), .A2(G125), .ZN(new_n190));
  NAND3_X1  g004(.A1(new_n189), .A2(G140), .A3(new_n190), .ZN(new_n191));
  NOR2_X1   g005(.A1(G125), .A2(G140), .ZN(new_n192));
  INV_X1    g006(.A(new_n192), .ZN(new_n193));
  AOI21_X1  g007(.A(new_n188), .B1(new_n191), .B2(new_n193), .ZN(new_n194));
  AND2_X1   g008(.A1(KEYINPUT75), .A2(G125), .ZN(new_n195));
  NOR2_X1   g009(.A1(KEYINPUT75), .A2(G125), .ZN(new_n196));
  NOR4_X1   g010(.A1(new_n195), .A2(new_n196), .A3(KEYINPUT16), .A4(G140), .ZN(new_n197));
  OAI21_X1  g011(.A(new_n187), .B1(new_n194), .B2(new_n197), .ZN(new_n198));
  NOR2_X1   g012(.A1(new_n195), .A2(new_n196), .ZN(new_n199));
  INV_X1    g013(.A(G140), .ZN(new_n200));
  NAND3_X1  g014(.A1(new_n199), .A2(new_n188), .A3(new_n200), .ZN(new_n201));
  AOI21_X1  g015(.A(new_n192), .B1(new_n199), .B2(G140), .ZN(new_n202));
  OAI211_X1 g016(.A(G146), .B(new_n201), .C1(new_n202), .C2(new_n188), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n198), .A2(new_n203), .ZN(new_n204));
  INV_X1    g018(.A(new_n204), .ZN(new_n205));
  INV_X1    g019(.A(G237), .ZN(new_n206));
  INV_X1    g020(.A(G953), .ZN(new_n207));
  NAND3_X1  g021(.A1(new_n206), .A2(new_n207), .A3(G214), .ZN(new_n208));
  INV_X1    g022(.A(G143), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  NOR2_X1   g024(.A1(G237), .A2(G953), .ZN(new_n211));
  NAND3_X1  g025(.A1(new_n211), .A2(G143), .A3(G214), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n210), .A2(new_n212), .ZN(new_n213));
  NAND3_X1  g027(.A1(new_n213), .A2(KEYINPUT17), .A3(G131), .ZN(new_n214));
  AND4_X1   g028(.A1(G143), .A2(new_n206), .A3(new_n207), .A4(G214), .ZN(new_n215));
  AOI21_X1  g029(.A(G143), .B1(new_n211), .B2(G214), .ZN(new_n216));
  OAI21_X1  g030(.A(G131), .B1(new_n215), .B2(new_n216), .ZN(new_n217));
  INV_X1    g031(.A(KEYINPUT17), .ZN(new_n218));
  INV_X1    g032(.A(G131), .ZN(new_n219));
  NAND3_X1  g033(.A1(new_n210), .A2(new_n219), .A3(new_n212), .ZN(new_n220));
  NAND3_X1  g034(.A1(new_n217), .A2(new_n218), .A3(new_n220), .ZN(new_n221));
  INV_X1    g035(.A(KEYINPUT89), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  NAND4_X1  g037(.A1(new_n217), .A2(new_n220), .A3(KEYINPUT89), .A4(new_n218), .ZN(new_n224));
  NAND4_X1  g038(.A1(new_n205), .A2(new_n214), .A3(new_n223), .A4(new_n224), .ZN(new_n225));
  INV_X1    g039(.A(KEYINPUT92), .ZN(new_n226));
  NAND2_X1  g040(.A1(KEYINPUT18), .A2(G131), .ZN(new_n227));
  XNOR2_X1  g041(.A(new_n213), .B(new_n227), .ZN(new_n228));
  XNOR2_X1  g042(.A(G125), .B(G140), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n229), .A2(new_n187), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n191), .A2(new_n193), .ZN(new_n231));
  OAI21_X1  g045(.A(new_n230), .B1(new_n231), .B2(new_n187), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n228), .A2(new_n232), .ZN(new_n233));
  NAND3_X1  g047(.A1(new_n225), .A2(new_n226), .A3(new_n233), .ZN(new_n234));
  XNOR2_X1  g048(.A(G113), .B(G122), .ZN(new_n235));
  XNOR2_X1  g049(.A(new_n235), .B(G104), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n223), .A2(new_n224), .ZN(new_n237));
  NAND3_X1  g051(.A1(new_n198), .A2(new_n203), .A3(new_n214), .ZN(new_n238));
  OAI21_X1  g052(.A(new_n233), .B1(new_n237), .B2(new_n238), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n239), .A2(KEYINPUT92), .ZN(new_n240));
  NAND3_X1  g054(.A1(new_n234), .A2(new_n236), .A3(new_n240), .ZN(new_n241));
  INV_X1    g055(.A(KEYINPUT88), .ZN(new_n242));
  XNOR2_X1  g056(.A(new_n236), .B(new_n242), .ZN(new_n243));
  NAND4_X1  g057(.A1(new_n225), .A2(KEYINPUT90), .A3(new_n233), .A4(new_n243), .ZN(new_n244));
  OAI211_X1 g058(.A(new_n233), .B(new_n243), .C1(new_n237), .C2(new_n238), .ZN(new_n245));
  INV_X1    g059(.A(KEYINPUT90), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n245), .A2(new_n246), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n244), .A2(new_n247), .ZN(new_n248));
  AOI21_X1  g062(.A(G902), .B1(new_n241), .B2(new_n248), .ZN(new_n249));
  OR2_X1    g063(.A1(new_n249), .A2(KEYINPUT93), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n249), .A2(KEYINPUT93), .ZN(new_n251));
  NAND3_X1  g065(.A1(new_n250), .A2(G475), .A3(new_n251), .ZN(new_n252));
  INV_X1    g066(.A(KEYINPUT19), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n229), .A2(new_n253), .ZN(new_n254));
  OAI211_X1 g068(.A(new_n187), .B(new_n254), .C1(new_n231), .C2(new_n253), .ZN(new_n255));
  NAND3_X1  g069(.A1(new_n203), .A2(new_n255), .A3(KEYINPUT87), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n217), .A2(new_n220), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n256), .A2(new_n257), .ZN(new_n258));
  AOI21_X1  g072(.A(KEYINPUT87), .B1(new_n203), .B2(new_n255), .ZN(new_n259));
  OAI21_X1  g073(.A(new_n233), .B1(new_n258), .B2(new_n259), .ZN(new_n260));
  AOI22_X1  g074(.A1(new_n244), .A2(new_n247), .B1(new_n260), .B2(new_n236), .ZN(new_n261));
  NOR4_X1   g075(.A1(new_n261), .A2(KEYINPUT20), .A3(G475), .A4(G902), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n260), .A2(new_n236), .ZN(new_n263));
  AND2_X1   g077(.A1(new_n245), .A2(new_n246), .ZN(new_n264));
  NOR2_X1   g078(.A1(new_n245), .A2(new_n246), .ZN(new_n265));
  OAI21_X1  g079(.A(new_n263), .B1(new_n264), .B2(new_n265), .ZN(new_n266));
  INV_X1    g080(.A(G475), .ZN(new_n267));
  INV_X1    g081(.A(G902), .ZN(new_n268));
  NAND3_X1  g082(.A1(new_n266), .A2(new_n267), .A3(new_n268), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n269), .A2(KEYINPUT20), .ZN(new_n270));
  INV_X1    g084(.A(KEYINPUT91), .ZN(new_n271));
  AOI21_X1  g085(.A(new_n262), .B1(new_n270), .B2(new_n271), .ZN(new_n272));
  NOR3_X1   g086(.A1(new_n269), .A2(KEYINPUT91), .A3(KEYINPUT20), .ZN(new_n273));
  OAI21_X1  g087(.A(new_n252), .B1(new_n272), .B2(new_n273), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n274), .A2(KEYINPUT94), .ZN(new_n275));
  INV_X1    g089(.A(KEYINPUT94), .ZN(new_n276));
  OAI211_X1 g090(.A(new_n252), .B(new_n276), .C1(new_n272), .C2(new_n273), .ZN(new_n277));
  XNOR2_X1  g091(.A(G116), .B(G122), .ZN(new_n278));
  INV_X1    g092(.A(G107), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n278), .A2(new_n279), .ZN(new_n280));
  INV_X1    g094(.A(G116), .ZN(new_n281));
  NAND3_X1  g095(.A1(new_n281), .A2(KEYINPUT14), .A3(G122), .ZN(new_n282));
  INV_X1    g096(.A(new_n278), .ZN(new_n283));
  OAI211_X1 g097(.A(G107), .B(new_n282), .C1(new_n283), .C2(KEYINPUT14), .ZN(new_n284));
  XNOR2_X1  g098(.A(G128), .B(G143), .ZN(new_n285));
  XNOR2_X1  g099(.A(new_n285), .B(KEYINPUT96), .ZN(new_n286));
  INV_X1    g100(.A(G134), .ZN(new_n287));
  AND2_X1   g101(.A1(new_n286), .A2(new_n287), .ZN(new_n288));
  NOR2_X1   g102(.A1(new_n286), .A2(new_n287), .ZN(new_n289));
  OAI211_X1 g103(.A(new_n280), .B(new_n284), .C1(new_n288), .C2(new_n289), .ZN(new_n290));
  NAND3_X1  g104(.A1(new_n209), .A2(KEYINPUT13), .A3(G128), .ZN(new_n291));
  XOR2_X1   g105(.A(new_n291), .B(KEYINPUT95), .Z(new_n292));
  INV_X1    g106(.A(G128), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n293), .A2(G143), .ZN(new_n294));
  NOR2_X1   g108(.A1(new_n293), .A2(G143), .ZN(new_n295));
  OAI21_X1  g109(.A(new_n294), .B1(new_n295), .B2(KEYINPUT13), .ZN(new_n296));
  OAI21_X1  g110(.A(G134), .B1(new_n292), .B2(new_n296), .ZN(new_n297));
  XNOR2_X1  g111(.A(new_n278), .B(new_n279), .ZN(new_n298));
  NAND2_X1  g112(.A1(new_n297), .A2(new_n298), .ZN(new_n299));
  OAI21_X1  g113(.A(new_n290), .B1(new_n288), .B2(new_n299), .ZN(new_n300));
  XOR2_X1   g114(.A(KEYINPUT9), .B(G234), .Z(new_n301));
  NAND3_X1  g115(.A1(new_n301), .A2(G217), .A3(new_n207), .ZN(new_n302));
  XNOR2_X1  g116(.A(new_n300), .B(new_n302), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n303), .A2(new_n268), .ZN(new_n304));
  INV_X1    g118(.A(KEYINPUT15), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n305), .A2(G478), .ZN(new_n306));
  XNOR2_X1  g120(.A(new_n304), .B(new_n306), .ZN(new_n307));
  INV_X1    g121(.A(new_n307), .ZN(new_n308));
  AND2_X1   g122(.A1(new_n207), .A2(G952), .ZN(new_n309));
  NAND2_X1  g123(.A1(G234), .A2(G237), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n309), .A2(new_n310), .ZN(new_n311));
  XNOR2_X1  g125(.A(new_n311), .B(KEYINPUT97), .ZN(new_n312));
  XOR2_X1   g126(.A(KEYINPUT21), .B(G898), .Z(new_n313));
  NAND3_X1  g127(.A1(new_n310), .A2(G902), .A3(G953), .ZN(new_n314));
  OAI21_X1  g128(.A(new_n312), .B1(new_n313), .B2(new_n314), .ZN(new_n315));
  INV_X1    g129(.A(new_n315), .ZN(new_n316));
  NOR2_X1   g130(.A1(new_n308), .A2(new_n316), .ZN(new_n317));
  NAND3_X1  g131(.A1(new_n275), .A2(new_n277), .A3(new_n317), .ZN(new_n318));
  OAI21_X1  g132(.A(G214), .B1(G237), .B2(G902), .ZN(new_n319));
  INV_X1    g133(.A(new_n301), .ZN(new_n320));
  OAI21_X1  g134(.A(G221), .B1(new_n320), .B2(G902), .ZN(new_n321));
  INV_X1    g135(.A(new_n321), .ZN(new_n322));
  NOR2_X1   g136(.A1(new_n279), .A2(G104), .ZN(new_n323));
  INV_X1    g137(.A(KEYINPUT3), .ZN(new_n324));
  NAND3_X1  g138(.A1(new_n324), .A2(new_n279), .A3(G104), .ZN(new_n325));
  INV_X1    g139(.A(KEYINPUT79), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n325), .A2(new_n326), .ZN(new_n327));
  NAND4_X1  g141(.A1(new_n324), .A2(new_n279), .A3(KEYINPUT79), .A4(G104), .ZN(new_n328));
  AOI21_X1  g142(.A(new_n323), .B1(new_n327), .B2(new_n328), .ZN(new_n329));
  INV_X1    g143(.A(KEYINPUT78), .ZN(new_n330));
  INV_X1    g144(.A(G104), .ZN(new_n331));
  NOR2_X1   g145(.A1(new_n331), .A2(G107), .ZN(new_n332));
  OAI21_X1  g146(.A(new_n330), .B1(new_n332), .B2(new_n324), .ZN(new_n333));
  OAI211_X1 g147(.A(KEYINPUT78), .B(KEYINPUT3), .C1(new_n331), .C2(G107), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n333), .A2(new_n334), .ZN(new_n335));
  INV_X1    g149(.A(G101), .ZN(new_n336));
  NAND3_X1  g150(.A1(new_n329), .A2(new_n335), .A3(new_n336), .ZN(new_n337));
  NOR2_X1   g151(.A1(new_n293), .A2(KEYINPUT1), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n187), .A2(G143), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n209), .A2(G146), .ZN(new_n340));
  NAND3_X1  g154(.A1(new_n338), .A2(new_n339), .A3(new_n340), .ZN(new_n341));
  OAI211_X1 g155(.A(new_n209), .B(G146), .C1(new_n293), .C2(KEYINPUT1), .ZN(new_n342));
  NAND3_X1  g156(.A1(new_n293), .A2(new_n187), .A3(G143), .ZN(new_n343));
  NAND3_X1  g157(.A1(new_n341), .A2(new_n342), .A3(new_n343), .ZN(new_n344));
  OAI21_X1  g158(.A(G101), .B1(new_n323), .B2(new_n332), .ZN(new_n345));
  NAND4_X1  g159(.A1(new_n337), .A2(KEYINPUT10), .A3(new_n344), .A4(new_n345), .ZN(new_n346));
  INV_X1    g160(.A(KEYINPUT82), .ZN(new_n347));
  XNOR2_X1  g161(.A(new_n346), .B(new_n347), .ZN(new_n348));
  INV_X1    g162(.A(KEYINPUT65), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n339), .A2(new_n340), .ZN(new_n350));
  NAND2_X1  g164(.A1(KEYINPUT0), .A2(G128), .ZN(new_n351));
  OAI21_X1  g165(.A(new_n349), .B1(new_n350), .B2(new_n351), .ZN(new_n352));
  INV_X1    g166(.A(new_n351), .ZN(new_n353));
  NOR2_X1   g167(.A1(KEYINPUT0), .A2(G128), .ZN(new_n354));
  NOR2_X1   g168(.A1(new_n353), .A2(new_n354), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n355), .A2(new_n350), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n352), .A2(new_n356), .ZN(new_n357));
  NAND3_X1  g171(.A1(new_n355), .A2(new_n349), .A3(new_n350), .ZN(new_n358));
  AND2_X1   g172(.A1(new_n357), .A2(new_n358), .ZN(new_n359));
  NAND2_X1  g173(.A1(new_n329), .A2(new_n335), .ZN(new_n360));
  INV_X1    g174(.A(KEYINPUT80), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n360), .A2(new_n361), .ZN(new_n362));
  INV_X1    g176(.A(KEYINPUT4), .ZN(new_n363));
  NAND3_X1  g177(.A1(new_n329), .A2(new_n335), .A3(KEYINPUT80), .ZN(new_n364));
  NAND4_X1  g178(.A1(new_n362), .A2(new_n363), .A3(G101), .A4(new_n364), .ZN(new_n365));
  AND3_X1   g179(.A1(new_n329), .A2(KEYINPUT80), .A3(new_n335), .ZN(new_n366));
  AOI21_X1  g180(.A(KEYINPUT80), .B1(new_n329), .B2(new_n335), .ZN(new_n367));
  NOR3_X1   g181(.A1(new_n366), .A2(new_n367), .A3(new_n336), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n337), .A2(KEYINPUT4), .ZN(new_n369));
  OAI211_X1 g183(.A(new_n359), .B(new_n365), .C1(new_n368), .C2(new_n369), .ZN(new_n370));
  INV_X1    g184(.A(KEYINPUT68), .ZN(new_n371));
  INV_X1    g185(.A(G137), .ZN(new_n372));
  NOR2_X1   g186(.A1(new_n372), .A2(G134), .ZN(new_n373));
  OAI21_X1  g187(.A(KEYINPUT11), .B1(new_n287), .B2(G137), .ZN(new_n374));
  INV_X1    g188(.A(KEYINPUT11), .ZN(new_n375));
  NAND3_X1  g189(.A1(new_n375), .A2(new_n372), .A3(G134), .ZN(new_n376));
  AOI211_X1 g190(.A(G131), .B(new_n373), .C1(new_n374), .C2(new_n376), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n374), .A2(new_n376), .ZN(new_n378));
  INV_X1    g192(.A(new_n373), .ZN(new_n379));
  AOI21_X1  g193(.A(new_n219), .B1(new_n378), .B2(new_n379), .ZN(new_n380));
  OAI21_X1  g194(.A(new_n371), .B1(new_n377), .B2(new_n380), .ZN(new_n381));
  AOI21_X1  g195(.A(new_n375), .B1(G134), .B2(new_n372), .ZN(new_n382));
  NOR3_X1   g196(.A1(new_n287), .A2(KEYINPUT11), .A3(G137), .ZN(new_n383));
  OAI21_X1  g197(.A(new_n379), .B1(new_n382), .B2(new_n383), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n384), .A2(G131), .ZN(new_n385));
  NAND3_X1  g199(.A1(new_n378), .A2(new_n219), .A3(new_n379), .ZN(new_n386));
  NAND3_X1  g200(.A1(new_n385), .A2(new_n386), .A3(KEYINPUT68), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n381), .A2(new_n387), .ZN(new_n388));
  INV_X1    g202(.A(new_n388), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n342), .A2(new_n343), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n390), .A2(KEYINPUT81), .ZN(new_n391));
  INV_X1    g205(.A(KEYINPUT81), .ZN(new_n392));
  NAND3_X1  g206(.A1(new_n342), .A2(new_n392), .A3(new_n343), .ZN(new_n393));
  NAND3_X1  g207(.A1(new_n391), .A2(new_n341), .A3(new_n393), .ZN(new_n394));
  NAND3_X1  g208(.A1(new_n337), .A2(new_n394), .A3(new_n345), .ZN(new_n395));
  INV_X1    g209(.A(new_n395), .ZN(new_n396));
  OR2_X1    g210(.A1(new_n396), .A2(KEYINPUT10), .ZN(new_n397));
  NAND4_X1  g211(.A1(new_n348), .A2(new_n370), .A3(new_n389), .A4(new_n397), .ZN(new_n398));
  XNOR2_X1  g212(.A(G110), .B(G140), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n207), .A2(G227), .ZN(new_n400));
  XNOR2_X1  g214(.A(new_n399), .B(new_n400), .ZN(new_n401));
  AND2_X1   g215(.A1(new_n398), .A2(new_n401), .ZN(new_n402));
  NAND3_X1  g216(.A1(new_n348), .A2(new_n370), .A3(new_n397), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n403), .A2(new_n388), .ZN(new_n404));
  NOR2_X1   g218(.A1(new_n377), .A2(new_n380), .ZN(new_n405));
  INV_X1    g219(.A(new_n405), .ZN(new_n406));
  AOI21_X1  g220(.A(new_n344), .B1(new_n337), .B2(new_n345), .ZN(new_n407));
  OAI211_X1 g221(.A(KEYINPUT12), .B(new_n406), .C1(new_n396), .C2(new_n407), .ZN(new_n408));
  INV_X1    g222(.A(KEYINPUT83), .ZN(new_n409));
  NAND2_X1  g223(.A1(new_n408), .A2(new_n409), .ZN(new_n410));
  AND2_X1   g224(.A1(new_n337), .A2(new_n345), .ZN(new_n411));
  OAI21_X1  g225(.A(new_n395), .B1(new_n411), .B2(new_n344), .ZN(new_n412));
  NAND4_X1  g226(.A1(new_n412), .A2(KEYINPUT83), .A3(KEYINPUT12), .A4(new_n406), .ZN(new_n413));
  OAI21_X1  g227(.A(new_n388), .B1(new_n396), .B2(new_n407), .ZN(new_n414));
  INV_X1    g228(.A(KEYINPUT12), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n414), .A2(new_n415), .ZN(new_n416));
  NAND3_X1  g230(.A1(new_n410), .A2(new_n413), .A3(new_n416), .ZN(new_n417));
  NAND2_X1  g231(.A1(new_n417), .A2(new_n398), .ZN(new_n418));
  XOR2_X1   g232(.A(new_n401), .B(KEYINPUT77), .Z(new_n419));
  AOI22_X1  g233(.A1(new_n402), .A2(new_n404), .B1(new_n418), .B2(new_n419), .ZN(new_n420));
  OAI21_X1  g234(.A(G469), .B1(new_n420), .B2(G902), .ZN(new_n421));
  INV_X1    g235(.A(G469), .ZN(new_n422));
  AOI21_X1  g236(.A(new_n401), .B1(new_n404), .B2(new_n398), .ZN(new_n423));
  AND3_X1   g237(.A1(new_n417), .A2(new_n398), .A3(new_n401), .ZN(new_n424));
  OAI211_X1 g238(.A(new_n422), .B(new_n268), .C1(new_n423), .C2(new_n424), .ZN(new_n425));
  AOI21_X1  g239(.A(new_n322), .B1(new_n421), .B2(new_n425), .ZN(new_n426));
  XOR2_X1   g240(.A(G110), .B(G122), .Z(new_n427));
  INV_X1    g241(.A(new_n427), .ZN(new_n428));
  XNOR2_X1  g242(.A(KEYINPUT67), .B(G119), .ZN(new_n429));
  NOR2_X1   g243(.A1(new_n429), .A2(new_n281), .ZN(new_n430));
  INV_X1    g244(.A(G119), .ZN(new_n431));
  NOR2_X1   g245(.A1(new_n431), .A2(G116), .ZN(new_n432));
  OR2_X1    g246(.A1(new_n430), .A2(new_n432), .ZN(new_n433));
  XNOR2_X1  g247(.A(KEYINPUT2), .B(G113), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n433), .A2(new_n434), .ZN(new_n435));
  OR3_X1    g249(.A1(new_n430), .A2(new_n434), .A3(new_n432), .ZN(new_n436));
  NAND2_X1  g250(.A1(new_n435), .A2(new_n436), .ZN(new_n437));
  OAI211_X1 g251(.A(new_n437), .B(new_n365), .C1(new_n368), .C2(new_n369), .ZN(new_n438));
  INV_X1    g252(.A(KEYINPUT5), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n430), .A2(new_n439), .ZN(new_n440));
  OAI211_X1 g254(.A(G113), .B(new_n440), .C1(new_n433), .C2(new_n439), .ZN(new_n441));
  NAND3_X1  g255(.A1(new_n441), .A2(new_n411), .A3(new_n436), .ZN(new_n442));
  AOI21_X1  g256(.A(new_n428), .B1(new_n438), .B2(new_n442), .ZN(new_n443));
  NOR2_X1   g257(.A1(new_n443), .A2(KEYINPUT6), .ZN(new_n444));
  INV_X1    g258(.A(new_n444), .ZN(new_n445));
  NAND3_X1  g259(.A1(new_n438), .A2(new_n442), .A3(new_n428), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n446), .A2(KEYINPUT84), .ZN(new_n447));
  INV_X1    g261(.A(KEYINPUT84), .ZN(new_n448));
  NAND4_X1  g262(.A1(new_n438), .A2(new_n448), .A3(new_n442), .A4(new_n428), .ZN(new_n449));
  AOI21_X1  g263(.A(new_n443), .B1(new_n447), .B2(new_n449), .ZN(new_n450));
  INV_X1    g264(.A(KEYINPUT6), .ZN(new_n451));
  OAI21_X1  g265(.A(new_n445), .B1(new_n450), .B2(new_n451), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n357), .A2(new_n358), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n453), .A2(new_n199), .ZN(new_n454));
  OAI21_X1  g268(.A(new_n454), .B1(new_n344), .B2(new_n199), .ZN(new_n455));
  INV_X1    g269(.A(G224), .ZN(new_n456));
  NOR2_X1   g270(.A1(new_n456), .A2(G953), .ZN(new_n457));
  XOR2_X1   g271(.A(new_n455), .B(new_n457), .Z(new_n458));
  INV_X1    g272(.A(new_n458), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n452), .A2(new_n459), .ZN(new_n460));
  OAI21_X1  g274(.A(G210), .B1(G237), .B2(G902), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n447), .A2(new_n449), .ZN(new_n462));
  INV_X1    g276(.A(KEYINPUT86), .ZN(new_n463));
  OAI21_X1  g277(.A(KEYINPUT7), .B1(new_n456), .B2(G953), .ZN(new_n464));
  AOI21_X1  g278(.A(new_n455), .B1(new_n463), .B2(new_n464), .ZN(new_n465));
  OR2_X1    g279(.A1(new_n464), .A2(new_n463), .ZN(new_n466));
  XNOR2_X1  g280(.A(new_n465), .B(new_n466), .ZN(new_n467));
  AOI21_X1  g281(.A(new_n411), .B1(new_n436), .B2(new_n441), .ZN(new_n468));
  INV_X1    g282(.A(KEYINPUT85), .ZN(new_n469));
  NOR2_X1   g283(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  XNOR2_X1  g284(.A(new_n470), .B(new_n442), .ZN(new_n471));
  XNOR2_X1  g285(.A(new_n427), .B(KEYINPUT8), .ZN(new_n472));
  OAI211_X1 g286(.A(new_n462), .B(new_n467), .C1(new_n471), .C2(new_n472), .ZN(new_n473));
  AND4_X1   g287(.A1(new_n268), .A2(new_n460), .A3(new_n461), .A4(new_n473), .ZN(new_n474));
  AOI21_X1  g288(.A(G902), .B1(new_n452), .B2(new_n459), .ZN(new_n475));
  AOI21_X1  g289(.A(new_n461), .B1(new_n475), .B2(new_n473), .ZN(new_n476));
  OAI211_X1 g290(.A(new_n319), .B(new_n426), .C1(new_n474), .C2(new_n476), .ZN(new_n477));
  NOR2_X1   g291(.A1(new_n318), .A2(new_n477), .ZN(new_n478));
  INV_X1    g292(.A(KEYINPUT32), .ZN(new_n479));
  INV_X1    g293(.A(KEYINPUT71), .ZN(new_n480));
  INV_X1    g294(.A(KEYINPUT31), .ZN(new_n481));
  AOI21_X1  g295(.A(new_n453), .B1(new_n381), .B2(new_n387), .ZN(new_n482));
  NAND3_X1  g296(.A1(new_n287), .A2(KEYINPUT66), .A3(G137), .ZN(new_n483));
  OAI21_X1  g297(.A(new_n483), .B1(new_n287), .B2(G137), .ZN(new_n484));
  NOR2_X1   g298(.A1(new_n373), .A2(KEYINPUT66), .ZN(new_n485));
  OAI21_X1  g299(.A(G131), .B1(new_n484), .B2(new_n485), .ZN(new_n486));
  NAND3_X1  g300(.A1(new_n486), .A2(new_n386), .A3(new_n344), .ZN(new_n487));
  INV_X1    g301(.A(new_n487), .ZN(new_n488));
  NOR3_X1   g302(.A1(new_n482), .A2(new_n437), .A3(new_n488), .ZN(new_n489));
  XNOR2_X1  g303(.A(KEYINPUT26), .B(KEYINPUT27), .ZN(new_n490));
  XNOR2_X1  g304(.A(new_n490), .B(G101), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n211), .A2(G210), .ZN(new_n492));
  XNOR2_X1  g306(.A(new_n491), .B(new_n492), .ZN(new_n493));
  INV_X1    g307(.A(new_n493), .ZN(new_n494));
  NOR2_X1   g308(.A1(new_n489), .A2(new_n494), .ZN(new_n495));
  AOI21_X1  g309(.A(new_n488), .B1(new_n388), .B2(new_n359), .ZN(new_n496));
  OAI21_X1  g310(.A(new_n487), .B1(new_n453), .B2(new_n405), .ZN(new_n497));
  XNOR2_X1  g311(.A(KEYINPUT64), .B(KEYINPUT30), .ZN(new_n498));
  AOI22_X1  g312(.A1(new_n496), .A2(KEYINPUT30), .B1(new_n497), .B2(new_n498), .ZN(new_n499));
  AOI21_X1  g313(.A(KEYINPUT69), .B1(new_n499), .B2(new_n437), .ZN(new_n500));
  NOR3_X1   g314(.A1(new_n377), .A2(new_n380), .A3(new_n371), .ZN(new_n501));
  AOI21_X1  g315(.A(KEYINPUT68), .B1(new_n385), .B2(new_n386), .ZN(new_n502));
  OAI21_X1  g316(.A(new_n359), .B1(new_n501), .B2(new_n502), .ZN(new_n503));
  NAND3_X1  g317(.A1(new_n503), .A2(KEYINPUT30), .A3(new_n487), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n497), .A2(new_n498), .ZN(new_n505));
  NAND4_X1  g319(.A1(new_n504), .A2(KEYINPUT69), .A3(new_n437), .A4(new_n505), .ZN(new_n506));
  INV_X1    g320(.A(new_n506), .ZN(new_n507));
  OAI211_X1 g321(.A(new_n481), .B(new_n495), .C1(new_n500), .C2(new_n507), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n508), .A2(KEYINPUT70), .ZN(new_n509));
  INV_X1    g323(.A(new_n489), .ZN(new_n510));
  NAND2_X1  g324(.A1(new_n510), .A2(new_n493), .ZN(new_n511));
  NAND3_X1  g325(.A1(new_n504), .A2(new_n437), .A3(new_n505), .ZN(new_n512));
  INV_X1    g326(.A(KEYINPUT69), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  AOI21_X1  g328(.A(new_n511), .B1(new_n514), .B2(new_n506), .ZN(new_n515));
  INV_X1    g329(.A(KEYINPUT70), .ZN(new_n516));
  NAND3_X1  g330(.A1(new_n515), .A2(new_n516), .A3(new_n481), .ZN(new_n517));
  NAND2_X1  g331(.A1(new_n509), .A2(new_n517), .ZN(new_n518));
  OAI21_X1  g332(.A(new_n495), .B1(new_n500), .B2(new_n507), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n497), .A2(new_n437), .ZN(new_n520));
  INV_X1    g334(.A(KEYINPUT28), .ZN(new_n521));
  NOR2_X1   g335(.A1(new_n489), .A2(new_n521), .ZN(new_n522));
  NOR4_X1   g336(.A1(new_n482), .A2(new_n437), .A3(KEYINPUT28), .A4(new_n488), .ZN(new_n523));
  OAI21_X1  g337(.A(new_n520), .B1(new_n522), .B2(new_n523), .ZN(new_n524));
  AOI22_X1  g338(.A1(new_n519), .A2(KEYINPUT31), .B1(new_n494), .B2(new_n524), .ZN(new_n525));
  AOI21_X1  g339(.A(G902), .B1(new_n518), .B2(new_n525), .ZN(new_n526));
  INV_X1    g340(.A(G472), .ZN(new_n527));
  AOI21_X1  g341(.A(new_n480), .B1(new_n526), .B2(new_n527), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n524), .A2(new_n494), .ZN(new_n529));
  OAI21_X1  g343(.A(new_n529), .B1(new_n515), .B2(new_n481), .ZN(new_n530));
  AOI21_X1  g344(.A(new_n530), .B1(new_n517), .B2(new_n509), .ZN(new_n531));
  NOR4_X1   g345(.A1(new_n531), .A2(KEYINPUT71), .A3(G472), .A4(G902), .ZN(new_n532));
  OAI21_X1  g346(.A(new_n479), .B1(new_n528), .B2(new_n532), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n514), .A2(new_n506), .ZN(new_n534));
  NAND3_X1  g348(.A1(new_n534), .A2(new_n510), .A3(new_n494), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n524), .A2(new_n493), .ZN(new_n536));
  AOI21_X1  g350(.A(KEYINPUT29), .B1(new_n535), .B2(new_n536), .ZN(new_n537));
  OR2_X1    g351(.A1(new_n522), .A2(new_n523), .ZN(new_n538));
  OAI21_X1  g352(.A(new_n437), .B1(new_n482), .B2(new_n488), .ZN(new_n539));
  NAND4_X1  g353(.A1(new_n538), .A2(KEYINPUT29), .A3(new_n493), .A4(new_n539), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n540), .A2(new_n268), .ZN(new_n541));
  OAI21_X1  g355(.A(G472), .B1(new_n537), .B2(new_n541), .ZN(new_n542));
  INV_X1    g356(.A(KEYINPUT72), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  NOR2_X1   g358(.A1(new_n508), .A2(KEYINPUT70), .ZN(new_n545));
  AOI21_X1  g359(.A(new_n516), .B1(new_n515), .B2(new_n481), .ZN(new_n546));
  OAI21_X1  g360(.A(new_n525), .B1(new_n545), .B2(new_n546), .ZN(new_n547));
  NAND4_X1  g361(.A1(new_n547), .A2(KEYINPUT32), .A3(new_n527), .A4(new_n268), .ZN(new_n548));
  OAI211_X1 g362(.A(KEYINPUT72), .B(G472), .C1(new_n537), .C2(new_n541), .ZN(new_n549));
  NAND3_X1  g363(.A1(new_n544), .A2(new_n548), .A3(new_n549), .ZN(new_n550));
  INV_X1    g364(.A(new_n550), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n533), .A2(new_n551), .ZN(new_n552));
  NOR2_X1   g366(.A1(new_n431), .A2(G128), .ZN(new_n553));
  XOR2_X1   g367(.A(KEYINPUT67), .B(G119), .Z(new_n554));
  AOI21_X1  g368(.A(new_n553), .B1(new_n554), .B2(G128), .ZN(new_n555));
  XOR2_X1   g369(.A(KEYINPUT24), .B(G110), .Z(new_n556));
  NAND2_X1  g370(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  XOR2_X1   g371(.A(new_n557), .B(KEYINPUT73), .Z(new_n558));
  INV_X1    g372(.A(KEYINPUT23), .ZN(new_n559));
  OAI21_X1  g373(.A(new_n559), .B1(new_n554), .B2(G128), .ZN(new_n560));
  OAI21_X1  g374(.A(new_n560), .B1(new_n555), .B2(new_n559), .ZN(new_n561));
  XNOR2_X1  g375(.A(new_n561), .B(KEYINPUT74), .ZN(new_n562));
  INV_X1    g376(.A(G110), .ZN(new_n563));
  OAI211_X1 g377(.A(new_n558), .B(new_n204), .C1(new_n562), .C2(new_n563), .ZN(new_n564));
  OAI22_X1  g378(.A1(new_n561), .A2(G110), .B1(new_n555), .B2(new_n556), .ZN(new_n565));
  NAND3_X1  g379(.A1(new_n565), .A2(new_n203), .A3(new_n230), .ZN(new_n566));
  NAND3_X1  g380(.A1(new_n207), .A2(G221), .A3(G234), .ZN(new_n567));
  XNOR2_X1  g381(.A(new_n567), .B(KEYINPUT22), .ZN(new_n568));
  XNOR2_X1  g382(.A(new_n568), .B(new_n372), .ZN(new_n569));
  AND3_X1   g383(.A1(new_n564), .A2(new_n566), .A3(new_n569), .ZN(new_n570));
  XOR2_X1   g384(.A(new_n569), .B(KEYINPUT76), .Z(new_n571));
  AOI21_X1  g385(.A(new_n571), .B1(new_n564), .B2(new_n566), .ZN(new_n572));
  NOR2_X1   g386(.A1(new_n570), .A2(new_n572), .ZN(new_n573));
  OAI21_X1  g387(.A(KEYINPUT25), .B1(new_n573), .B2(G902), .ZN(new_n574));
  INV_X1    g388(.A(G217), .ZN(new_n575));
  AOI21_X1  g389(.A(new_n575), .B1(G234), .B2(new_n268), .ZN(new_n576));
  INV_X1    g390(.A(KEYINPUT25), .ZN(new_n577));
  OAI211_X1 g391(.A(new_n577), .B(new_n268), .C1(new_n570), .C2(new_n572), .ZN(new_n578));
  NAND3_X1  g392(.A1(new_n574), .A2(new_n576), .A3(new_n578), .ZN(new_n579));
  INV_X1    g393(.A(new_n573), .ZN(new_n580));
  NOR2_X1   g394(.A1(new_n576), .A2(G902), .ZN(new_n581));
  NAND2_X1  g395(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  NAND2_X1  g396(.A1(new_n579), .A2(new_n582), .ZN(new_n583));
  INV_X1    g397(.A(new_n583), .ZN(new_n584));
  NAND3_X1  g398(.A1(new_n478), .A2(new_n552), .A3(new_n584), .ZN(new_n585));
  XOR2_X1   g399(.A(KEYINPUT98), .B(G101), .Z(new_n586));
  XNOR2_X1  g400(.A(new_n585), .B(new_n586), .ZN(G3));
  XOR2_X1   g401(.A(new_n303), .B(KEYINPUT33), .Z(new_n588));
  NOR2_X1   g402(.A1(new_n588), .A2(G902), .ZN(new_n589));
  XOR2_X1   g403(.A(KEYINPUT99), .B(G478), .Z(new_n590));
  AOI22_X1  g404(.A1(new_n589), .A2(G478), .B1(new_n304), .B2(new_n590), .ZN(new_n591));
  AOI21_X1  g405(.A(new_n591), .B1(new_n275), .B2(new_n277), .ZN(new_n592));
  INV_X1    g406(.A(new_n319), .ZN(new_n593));
  INV_X1    g407(.A(new_n443), .ZN(new_n594));
  NAND2_X1  g408(.A1(new_n462), .A2(new_n594), .ZN(new_n595));
  AOI21_X1  g409(.A(new_n444), .B1(new_n595), .B2(KEYINPUT6), .ZN(new_n596));
  OAI211_X1 g410(.A(new_n268), .B(new_n473), .C1(new_n596), .C2(new_n458), .ZN(new_n597));
  INV_X1    g411(.A(new_n461), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n597), .A2(new_n598), .ZN(new_n599));
  NAND3_X1  g413(.A1(new_n475), .A2(new_n461), .A3(new_n473), .ZN(new_n600));
  AOI21_X1  g414(.A(new_n593), .B1(new_n599), .B2(new_n600), .ZN(new_n601));
  AND3_X1   g415(.A1(new_n592), .A2(new_n601), .A3(new_n315), .ZN(new_n602));
  NAND3_X1  g416(.A1(new_n547), .A2(new_n527), .A3(new_n268), .ZN(new_n603));
  NAND2_X1  g417(.A1(new_n603), .A2(KEYINPUT71), .ZN(new_n604));
  NAND3_X1  g418(.A1(new_n526), .A2(new_n480), .A3(new_n527), .ZN(new_n605));
  NAND2_X1  g419(.A1(new_n547), .A2(new_n268), .ZN(new_n606));
  AOI22_X1  g420(.A1(new_n604), .A2(new_n605), .B1(G472), .B2(new_n606), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n421), .A2(new_n425), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n608), .A2(new_n321), .ZN(new_n609));
  NOR2_X1   g423(.A1(new_n609), .A2(new_n583), .ZN(new_n610));
  NAND3_X1  g424(.A1(new_n602), .A2(new_n607), .A3(new_n610), .ZN(new_n611));
  XOR2_X1   g425(.A(KEYINPUT34), .B(G104), .Z(new_n612));
  XNOR2_X1  g426(.A(new_n611), .B(new_n612), .ZN(G6));
  XNOR2_X1  g427(.A(new_n315), .B(KEYINPUT100), .ZN(new_n614));
  AOI211_X1 g428(.A(new_n593), .B(new_n614), .C1(new_n599), .C2(new_n600), .ZN(new_n615));
  AND3_X1   g429(.A1(new_n615), .A2(new_n607), .A3(new_n610), .ZN(new_n616));
  INV_X1    g430(.A(KEYINPUT20), .ZN(new_n617));
  AOI21_X1  g431(.A(G475), .B1(new_n248), .B2(new_n263), .ZN(new_n618));
  AOI21_X1  g432(.A(new_n617), .B1(new_n618), .B2(new_n268), .ZN(new_n619));
  OAI21_X1  g433(.A(new_n252), .B1(new_n262), .B2(new_n619), .ZN(new_n620));
  NOR2_X1   g434(.A1(new_n620), .A2(new_n307), .ZN(new_n621));
  NAND2_X1  g435(.A1(new_n616), .A2(new_n621), .ZN(new_n622));
  XOR2_X1   g436(.A(KEYINPUT35), .B(G107), .Z(new_n623));
  XNOR2_X1  g437(.A(new_n622), .B(new_n623), .ZN(G9));
  INV_X1    g438(.A(new_n277), .ZN(new_n625));
  NAND3_X1  g439(.A1(new_n618), .A2(new_n617), .A3(new_n268), .ZN(new_n626));
  OAI21_X1  g440(.A(new_n626), .B1(new_n619), .B2(KEYINPUT91), .ZN(new_n627));
  NAND3_X1  g441(.A1(new_n270), .A2(new_n271), .A3(new_n262), .ZN(new_n628));
  NAND2_X1  g442(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  AOI21_X1  g443(.A(new_n276), .B1(new_n629), .B2(new_n252), .ZN(new_n630));
  NOR2_X1   g444(.A1(new_n625), .A2(new_n630), .ZN(new_n631));
  NAND4_X1  g445(.A1(new_n631), .A2(new_n601), .A3(new_n426), .A4(new_n317), .ZN(new_n632));
  INV_X1    g446(.A(new_n607), .ZN(new_n633));
  NOR2_X1   g447(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  NAND2_X1  g448(.A1(new_n564), .A2(new_n566), .ZN(new_n635));
  NOR2_X1   g449(.A1(new_n571), .A2(KEYINPUT36), .ZN(new_n636));
  XNOR2_X1  g450(.A(new_n635), .B(new_n636), .ZN(new_n637));
  NAND2_X1  g451(.A1(new_n637), .A2(new_n581), .ZN(new_n638));
  NAND2_X1  g452(.A1(new_n579), .A2(new_n638), .ZN(new_n639));
  NAND2_X1  g453(.A1(new_n634), .A2(new_n639), .ZN(new_n640));
  XNOR2_X1  g454(.A(new_n640), .B(KEYINPUT37), .ZN(new_n641));
  XNOR2_X1  g455(.A(new_n641), .B(new_n563), .ZN(G12));
  INV_X1    g456(.A(new_n639), .ZN(new_n643));
  AOI21_X1  g457(.A(new_n643), .B1(new_n533), .B2(new_n551), .ZN(new_n644));
  INV_X1    g458(.A(new_n477), .ZN(new_n645));
  XNOR2_X1  g459(.A(KEYINPUT101), .B(G900), .ZN(new_n646));
  OAI21_X1  g460(.A(new_n312), .B1(new_n314), .B2(new_n646), .ZN(new_n647));
  NAND4_X1  g461(.A1(new_n644), .A2(new_n645), .A3(new_n621), .A4(new_n647), .ZN(new_n648));
  XNOR2_X1  g462(.A(new_n648), .B(G128), .ZN(G30));
  NAND2_X1  g463(.A1(new_n599), .A2(new_n600), .ZN(new_n650));
  INV_X1    g464(.A(KEYINPUT102), .ZN(new_n651));
  XNOR2_X1  g465(.A(new_n650), .B(new_n651), .ZN(new_n652));
  XNOR2_X1  g466(.A(new_n652), .B(KEYINPUT38), .ZN(new_n653));
  AOI21_X1  g467(.A(new_n493), .B1(new_n510), .B2(new_n539), .ZN(new_n654));
  XOR2_X1   g468(.A(new_n654), .B(KEYINPUT103), .Z(new_n655));
  NOR3_X1   g469(.A1(new_n655), .A2(KEYINPUT104), .A3(new_n515), .ZN(new_n656));
  NOR2_X1   g470(.A1(new_n656), .A2(G902), .ZN(new_n657));
  OAI21_X1  g471(.A(KEYINPUT104), .B1(new_n655), .B2(new_n515), .ZN(new_n658));
  AND2_X1   g472(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  OAI211_X1 g473(.A(new_n533), .B(new_n548), .C1(new_n527), .C2(new_n659), .ZN(new_n660));
  NOR3_X1   g474(.A1(new_n631), .A2(new_n593), .A3(new_n307), .ZN(new_n661));
  AND2_X1   g475(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  XOR2_X1   g476(.A(new_n647), .B(KEYINPUT105), .Z(new_n663));
  XNOR2_X1  g477(.A(new_n663), .B(KEYINPUT39), .ZN(new_n664));
  OAI21_X1  g478(.A(KEYINPUT40), .B1(new_n609), .B2(new_n664), .ZN(new_n665));
  NOR2_X1   g479(.A1(new_n609), .A2(new_n664), .ZN(new_n666));
  INV_X1    g480(.A(KEYINPUT40), .ZN(new_n667));
  AOI21_X1  g481(.A(new_n639), .B1(new_n666), .B2(new_n667), .ZN(new_n668));
  NAND4_X1  g482(.A1(new_n653), .A2(new_n662), .A3(new_n665), .A4(new_n668), .ZN(new_n669));
  XNOR2_X1  g483(.A(new_n669), .B(G143), .ZN(G45));
  NAND2_X1  g484(.A1(new_n592), .A2(new_n647), .ZN(new_n671));
  INV_X1    g485(.A(new_n671), .ZN(new_n672));
  NAND3_X1  g486(.A1(new_n672), .A2(new_n644), .A3(new_n645), .ZN(new_n673));
  XNOR2_X1  g487(.A(new_n673), .B(G146), .ZN(G48));
  AOI21_X1  g488(.A(new_n583), .B1(new_n533), .B2(new_n551), .ZN(new_n675));
  OAI21_X1  g489(.A(new_n268), .B1(new_n423), .B2(new_n424), .ZN(new_n676));
  NAND2_X1  g490(.A1(new_n676), .A2(G469), .ZN(new_n677));
  AND3_X1   g491(.A1(new_n677), .A2(new_n321), .A3(new_n425), .ZN(new_n678));
  NAND3_X1  g492(.A1(new_n602), .A2(new_n675), .A3(new_n678), .ZN(new_n679));
  XNOR2_X1  g493(.A(new_n679), .B(KEYINPUT41), .ZN(new_n680));
  XNOR2_X1  g494(.A(new_n680), .B(G113), .ZN(G15));
  NAND4_X1  g495(.A1(new_n675), .A2(new_n615), .A3(new_n621), .A4(new_n678), .ZN(new_n682));
  XNOR2_X1  g496(.A(new_n682), .B(G116), .ZN(G18));
  OAI211_X1 g497(.A(new_n319), .B(new_n678), .C1(new_n474), .C2(new_n476), .ZN(new_n684));
  NAND2_X1  g498(.A1(new_n684), .A2(KEYINPUT106), .ZN(new_n685));
  INV_X1    g499(.A(KEYINPUT106), .ZN(new_n686));
  NAND4_X1  g500(.A1(new_n650), .A2(new_n686), .A3(new_n319), .A4(new_n678), .ZN(new_n687));
  NAND2_X1  g501(.A1(new_n685), .A2(new_n687), .ZN(new_n688));
  INV_X1    g502(.A(new_n318), .ZN(new_n689));
  NAND3_X1  g503(.A1(new_n688), .A2(new_n644), .A3(new_n689), .ZN(new_n690));
  XNOR2_X1  g504(.A(new_n690), .B(G119), .ZN(G21));
  NAND2_X1  g505(.A1(new_n606), .A2(G472), .ZN(new_n692));
  NAND2_X1  g506(.A1(new_n519), .A2(KEYINPUT31), .ZN(new_n693));
  AND2_X1   g507(.A1(new_n538), .A2(new_n539), .ZN(new_n694));
  OAI211_X1 g508(.A(new_n518), .B(new_n693), .C1(new_n493), .C2(new_n694), .ZN(new_n695));
  NOR2_X1   g509(.A1(G472), .A2(G902), .ZN(new_n696));
  NAND2_X1  g510(.A1(new_n695), .A2(new_n696), .ZN(new_n697));
  NAND3_X1  g511(.A1(new_n692), .A2(new_n697), .A3(new_n584), .ZN(new_n698));
  NAND2_X1  g512(.A1(new_n698), .A2(KEYINPUT107), .ZN(new_n699));
  INV_X1    g513(.A(KEYINPUT107), .ZN(new_n700));
  NAND4_X1  g514(.A1(new_n692), .A2(new_n697), .A3(new_n584), .A4(new_n700), .ZN(new_n701));
  NAND2_X1  g515(.A1(new_n699), .A2(new_n701), .ZN(new_n702));
  AOI211_X1 g516(.A(new_n307), .B(new_n614), .C1(new_n275), .C2(new_n277), .ZN(new_n703));
  INV_X1    g517(.A(new_n684), .ZN(new_n704));
  NAND3_X1  g518(.A1(new_n702), .A2(new_n703), .A3(new_n704), .ZN(new_n705));
  XNOR2_X1  g519(.A(new_n705), .B(G122), .ZN(G24));
  NAND3_X1  g520(.A1(new_n692), .A2(new_n697), .A3(new_n639), .ZN(new_n707));
  INV_X1    g521(.A(new_n707), .ZN(new_n708));
  NAND3_X1  g522(.A1(new_n672), .A2(new_n688), .A3(new_n708), .ZN(new_n709));
  XNOR2_X1  g523(.A(new_n709), .B(G125), .ZN(G27));
  NAND3_X1  g524(.A1(new_n599), .A2(new_n319), .A3(new_n600), .ZN(new_n711));
  NAND2_X1  g525(.A1(new_n711), .A2(KEYINPUT109), .ZN(new_n712));
  NAND2_X1  g526(.A1(new_n609), .A2(KEYINPUT108), .ZN(new_n713));
  INV_X1    g527(.A(KEYINPUT108), .ZN(new_n714));
  NAND2_X1  g528(.A1(new_n426), .A2(new_n714), .ZN(new_n715));
  NAND2_X1  g529(.A1(new_n713), .A2(new_n715), .ZN(new_n716));
  INV_X1    g530(.A(KEYINPUT109), .ZN(new_n717));
  NAND4_X1  g531(.A1(new_n599), .A2(new_n717), .A3(new_n319), .A4(new_n600), .ZN(new_n718));
  NAND3_X1  g532(.A1(new_n712), .A2(new_n716), .A3(new_n718), .ZN(new_n719));
  INV_X1    g533(.A(new_n719), .ZN(new_n720));
  AND3_X1   g534(.A1(new_n603), .A2(KEYINPUT110), .A3(new_n479), .ZN(new_n721));
  AOI21_X1  g535(.A(KEYINPUT110), .B1(new_n603), .B2(new_n479), .ZN(new_n722));
  NOR2_X1   g536(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  AOI21_X1  g537(.A(new_n583), .B1(new_n723), .B2(new_n551), .ZN(new_n724));
  NAND4_X1  g538(.A1(new_n720), .A2(new_n724), .A3(KEYINPUT42), .A4(new_n672), .ZN(new_n725));
  AOI21_X1  g539(.A(KEYINPUT32), .B1(new_n604), .B2(new_n605), .ZN(new_n726));
  OAI21_X1  g540(.A(new_n584), .B1(new_n726), .B2(new_n550), .ZN(new_n727));
  NOR3_X1   g541(.A1(new_n719), .A2(new_n727), .A3(new_n671), .ZN(new_n728));
  OAI21_X1  g542(.A(new_n725), .B1(new_n728), .B2(KEYINPUT42), .ZN(new_n729));
  XNOR2_X1  g543(.A(new_n729), .B(G131), .ZN(G33));
  NAND2_X1  g544(.A1(new_n621), .A2(new_n647), .ZN(new_n731));
  NOR3_X1   g545(.A1(new_n719), .A2(new_n727), .A3(new_n731), .ZN(new_n732));
  XNOR2_X1  g546(.A(new_n732), .B(new_n287), .ZN(G36));
  NAND2_X1  g547(.A1(new_n631), .A2(KEYINPUT112), .ZN(new_n734));
  INV_X1    g548(.A(KEYINPUT43), .ZN(new_n735));
  NAND2_X1  g549(.A1(new_n734), .A2(new_n735), .ZN(new_n736));
  NAND2_X1  g550(.A1(new_n275), .A2(new_n277), .ZN(new_n737));
  NOR2_X1   g551(.A1(new_n737), .A2(new_n591), .ZN(new_n738));
  NAND2_X1  g552(.A1(new_n736), .A2(new_n738), .ZN(new_n739));
  INV_X1    g553(.A(new_n738), .ZN(new_n740));
  NAND3_X1  g554(.A1(new_n740), .A2(new_n734), .A3(new_n735), .ZN(new_n741));
  NAND2_X1  g555(.A1(new_n739), .A2(new_n741), .ZN(new_n742));
  NAND3_X1  g556(.A1(new_n742), .A2(new_n633), .A3(new_n639), .ZN(new_n743));
  INV_X1    g557(.A(KEYINPUT44), .ZN(new_n744));
  NAND2_X1  g558(.A1(new_n743), .A2(new_n744), .ZN(new_n745));
  NAND2_X1  g559(.A1(new_n712), .A2(new_n718), .ZN(new_n746));
  INV_X1    g560(.A(new_n746), .ZN(new_n747));
  NAND4_X1  g561(.A1(new_n742), .A2(KEYINPUT44), .A3(new_n633), .A4(new_n639), .ZN(new_n748));
  OR2_X1    g562(.A1(new_n420), .A2(KEYINPUT45), .ZN(new_n749));
  NAND2_X1  g563(.A1(new_n420), .A2(KEYINPUT45), .ZN(new_n750));
  NAND3_X1  g564(.A1(new_n749), .A2(G469), .A3(new_n750), .ZN(new_n751));
  NAND2_X1  g565(.A1(G469), .A2(G902), .ZN(new_n752));
  NAND3_X1  g566(.A1(new_n751), .A2(KEYINPUT46), .A3(new_n752), .ZN(new_n753));
  NAND2_X1  g567(.A1(new_n753), .A2(new_n425), .ZN(new_n754));
  INV_X1    g568(.A(KEYINPUT111), .ZN(new_n755));
  NAND2_X1  g569(.A1(new_n754), .A2(new_n755), .ZN(new_n756));
  NAND3_X1  g570(.A1(new_n753), .A2(KEYINPUT111), .A3(new_n425), .ZN(new_n757));
  AND2_X1   g571(.A1(new_n751), .A2(new_n752), .ZN(new_n758));
  OAI211_X1 g572(.A(new_n756), .B(new_n757), .C1(KEYINPUT46), .C2(new_n758), .ZN(new_n759));
  NAND2_X1  g573(.A1(new_n759), .A2(new_n321), .ZN(new_n760));
  NOR2_X1   g574(.A1(new_n760), .A2(new_n664), .ZN(new_n761));
  NAND4_X1  g575(.A1(new_n745), .A2(new_n747), .A3(new_n748), .A4(new_n761), .ZN(new_n762));
  XNOR2_X1  g576(.A(new_n762), .B(G137), .ZN(G39));
  XNOR2_X1  g577(.A(KEYINPUT113), .B(KEYINPUT47), .ZN(new_n764));
  AND3_X1   g578(.A1(new_n759), .A2(new_n321), .A3(new_n764), .ZN(new_n765));
  NOR2_X1   g579(.A1(KEYINPUT113), .A2(KEYINPUT47), .ZN(new_n766));
  AOI21_X1  g580(.A(new_n766), .B1(new_n759), .B2(new_n321), .ZN(new_n767));
  NOR3_X1   g581(.A1(new_n765), .A2(new_n767), .A3(new_n552), .ZN(new_n768));
  NAND4_X1  g582(.A1(new_n768), .A2(new_n583), .A3(new_n672), .A4(new_n747), .ZN(new_n769));
  XNOR2_X1  g583(.A(new_n769), .B(KEYINPUT114), .ZN(new_n770));
  XNOR2_X1  g584(.A(new_n770), .B(G140), .ZN(G42));
  INV_X1    g585(.A(new_n653), .ZN(new_n772));
  AND2_X1   g586(.A1(new_n677), .A2(new_n425), .ZN(new_n773));
  XNOR2_X1  g587(.A(new_n773), .B(KEYINPUT49), .ZN(new_n774));
  NOR4_X1   g588(.A1(new_n660), .A2(new_n740), .A3(new_n583), .A4(new_n322), .ZN(new_n775));
  NAND4_X1  g589(.A1(new_n772), .A2(new_n319), .A3(new_n774), .A4(new_n775), .ZN(new_n776));
  INV_X1    g590(.A(new_n647), .ZN(new_n777));
  NOR3_X1   g591(.A1(new_n609), .A2(new_n639), .A3(new_n777), .ZN(new_n778));
  NAND4_X1  g592(.A1(new_n660), .A2(new_n661), .A3(new_n650), .A4(new_n778), .ZN(new_n779));
  NAND4_X1  g593(.A1(new_n779), .A2(new_n709), .A3(new_n648), .A4(new_n673), .ZN(new_n780));
  XOR2_X1   g594(.A(KEYINPUT118), .B(KEYINPUT52), .Z(new_n781));
  NAND2_X1  g595(.A1(new_n780), .A2(new_n781), .ZN(new_n782));
  AOI21_X1  g596(.A(KEYINPUT117), .B1(new_n709), .B2(new_n648), .ZN(new_n783));
  INV_X1    g597(.A(new_n673), .ZN(new_n784));
  NOR2_X1   g598(.A1(new_n783), .A2(new_n784), .ZN(new_n785));
  NAND3_X1  g599(.A1(new_n709), .A2(new_n648), .A3(KEYINPUT117), .ZN(new_n786));
  NAND3_X1  g600(.A1(new_n785), .A2(new_n779), .A3(new_n786), .ZN(new_n787));
  INV_X1    g601(.A(KEYINPUT52), .ZN(new_n788));
  OAI21_X1  g602(.A(new_n782), .B1(new_n787), .B2(new_n788), .ZN(new_n789));
  AND4_X1   g603(.A1(new_n679), .A2(new_n682), .A3(new_n690), .A4(new_n705), .ZN(new_n790));
  NAND4_X1  g604(.A1(new_n615), .A2(new_n607), .A3(new_n592), .A4(new_n610), .ZN(new_n791));
  OAI21_X1  g605(.A(new_n791), .B1(new_n727), .B2(new_n632), .ZN(new_n792));
  INV_X1    g606(.A(KEYINPUT115), .ZN(new_n793));
  NAND2_X1  g607(.A1(new_n792), .A2(new_n793), .ZN(new_n794));
  OAI211_X1 g608(.A(new_n791), .B(KEYINPUT115), .C1(new_n727), .C2(new_n632), .ZN(new_n795));
  NAND2_X1  g609(.A1(new_n794), .A2(new_n795), .ZN(new_n796));
  NOR2_X1   g610(.A1(new_n737), .A2(new_n307), .ZN(new_n797));
  AOI22_X1  g611(.A1(new_n634), .A2(new_n639), .B1(new_n616), .B2(new_n797), .ZN(new_n798));
  NAND3_X1  g612(.A1(new_n790), .A2(new_n796), .A3(new_n798), .ZN(new_n799));
  NOR3_X1   g613(.A1(new_n719), .A2(new_n671), .A3(new_n707), .ZN(new_n800));
  NOR2_X1   g614(.A1(new_n609), .A2(new_n620), .ZN(new_n801));
  OAI211_X1 g615(.A(new_n639), .B(new_n801), .C1(new_n726), .C2(new_n550), .ZN(new_n802));
  NOR2_X1   g616(.A1(new_n308), .A2(new_n777), .ZN(new_n803));
  NAND3_X1  g617(.A1(new_n712), .A2(new_n718), .A3(new_n803), .ZN(new_n804));
  NOR2_X1   g618(.A1(new_n802), .A2(new_n804), .ZN(new_n805));
  NOR3_X1   g619(.A1(new_n732), .A2(new_n800), .A3(new_n805), .ZN(new_n806));
  NAND2_X1  g620(.A1(new_n806), .A2(new_n729), .ZN(new_n807));
  NOR2_X1   g621(.A1(new_n799), .A2(new_n807), .ZN(new_n808));
  NAND3_X1  g622(.A1(new_n789), .A2(KEYINPUT53), .A3(new_n808), .ZN(new_n809));
  INV_X1    g623(.A(KEYINPUT54), .ZN(new_n810));
  XNOR2_X1  g624(.A(new_n780), .B(KEYINPUT52), .ZN(new_n811));
  INV_X1    g625(.A(new_n795), .ZN(new_n812));
  AOI21_X1  g626(.A(KEYINPUT115), .B1(new_n585), .B2(new_n791), .ZN(new_n813));
  OAI21_X1  g627(.A(new_n798), .B1(new_n812), .B2(new_n813), .ZN(new_n814));
  NAND4_X1  g628(.A1(new_n679), .A2(new_n682), .A3(new_n690), .A4(new_n705), .ZN(new_n815));
  NOR2_X1   g629(.A1(new_n814), .A2(new_n815), .ZN(new_n816));
  AND2_X1   g630(.A1(new_n806), .A2(new_n729), .ZN(new_n817));
  INV_X1    g631(.A(KEYINPUT116), .ZN(new_n818));
  NAND3_X1  g632(.A1(new_n816), .A2(new_n817), .A3(new_n818), .ZN(new_n819));
  OAI21_X1  g633(.A(KEYINPUT116), .B1(new_n799), .B2(new_n807), .ZN(new_n820));
  AOI21_X1  g634(.A(new_n811), .B1(new_n819), .B2(new_n820), .ZN(new_n821));
  XNOR2_X1  g635(.A(KEYINPUT119), .B(KEYINPUT53), .ZN(new_n822));
  OAI211_X1 g636(.A(new_n809), .B(new_n810), .C1(new_n821), .C2(new_n822), .ZN(new_n823));
  INV_X1    g637(.A(new_n823), .ZN(new_n824));
  AOI21_X1  g638(.A(new_n312), .B1(new_n739), .B2(new_n741), .ZN(new_n825));
  AND2_X1   g639(.A1(new_n825), .A2(new_n702), .ZN(new_n826));
  NAND2_X1  g640(.A1(new_n826), .A2(new_n688), .ZN(new_n827));
  NAND2_X1  g641(.A1(new_n747), .A2(new_n678), .ZN(new_n828));
  NOR2_X1   g642(.A1(new_n828), .A2(new_n583), .ZN(new_n829));
  NOR2_X1   g643(.A1(new_n660), .A2(new_n312), .ZN(new_n830));
  NAND3_X1  g644(.A1(new_n829), .A2(new_n592), .A3(new_n830), .ZN(new_n831));
  NAND3_X1  g645(.A1(new_n827), .A2(new_n309), .A3(new_n831), .ZN(new_n832));
  INV_X1    g646(.A(KEYINPUT121), .ZN(new_n833));
  NAND2_X1  g647(.A1(new_n832), .A2(new_n833), .ZN(new_n834));
  NAND4_X1  g648(.A1(new_n827), .A2(KEYINPUT121), .A3(new_n309), .A4(new_n831), .ZN(new_n835));
  AOI211_X1 g649(.A(new_n312), .B(new_n828), .C1(new_n739), .C2(new_n741), .ZN(new_n836));
  NAND2_X1  g650(.A1(new_n836), .A2(new_n724), .ZN(new_n837));
  OR2_X1    g651(.A1(new_n837), .A2(KEYINPUT48), .ZN(new_n838));
  NAND2_X1  g652(.A1(new_n837), .A2(KEYINPUT48), .ZN(new_n839));
  AOI22_X1  g653(.A1(new_n834), .A2(new_n835), .B1(new_n838), .B2(new_n839), .ZN(new_n840));
  INV_X1    g654(.A(KEYINPUT50), .ZN(new_n841));
  NOR2_X1   g655(.A1(new_n653), .A2(new_n319), .ZN(new_n842));
  INV_X1    g656(.A(new_n842), .ZN(new_n843));
  NAND3_X1  g657(.A1(new_n825), .A2(new_n678), .A3(new_n702), .ZN(new_n844));
  OAI21_X1  g658(.A(new_n841), .B1(new_n843), .B2(new_n844), .ZN(new_n845));
  NAND4_X1  g659(.A1(new_n826), .A2(KEYINPUT50), .A3(new_n678), .A4(new_n842), .ZN(new_n846));
  AND2_X1   g660(.A1(new_n845), .A2(new_n846), .ZN(new_n847));
  NAND2_X1  g661(.A1(new_n773), .A2(new_n322), .ZN(new_n848));
  OAI21_X1  g662(.A(new_n848), .B1(new_n765), .B2(new_n767), .ZN(new_n849));
  NAND3_X1  g663(.A1(new_n826), .A2(new_n849), .A3(new_n747), .ZN(new_n850));
  NAND2_X1  g664(.A1(new_n836), .A2(new_n708), .ZN(new_n851));
  NAND4_X1  g665(.A1(new_n829), .A2(new_n631), .A3(new_n591), .A4(new_n830), .ZN(new_n852));
  NAND3_X1  g666(.A1(new_n850), .A2(new_n851), .A3(new_n852), .ZN(new_n853));
  NOR3_X1   g667(.A1(new_n847), .A2(new_n853), .A3(KEYINPUT51), .ZN(new_n854));
  INV_X1    g668(.A(KEYINPUT51), .ZN(new_n855));
  INV_X1    g669(.A(new_n853), .ZN(new_n856));
  NAND2_X1  g670(.A1(new_n845), .A2(new_n846), .ZN(new_n857));
  AOI21_X1  g671(.A(new_n855), .B1(new_n856), .B2(new_n857), .ZN(new_n858));
  OAI21_X1  g672(.A(new_n840), .B1(new_n854), .B2(new_n858), .ZN(new_n859));
  INV_X1    g673(.A(new_n811), .ZN(new_n860));
  AOI21_X1  g674(.A(new_n818), .B1(new_n816), .B2(new_n817), .ZN(new_n861));
  NOR3_X1   g675(.A1(new_n799), .A2(new_n807), .A3(KEYINPUT116), .ZN(new_n862));
  OAI211_X1 g676(.A(new_n822), .B(new_n860), .C1(new_n861), .C2(new_n862), .ZN(new_n863));
  NAND2_X1  g677(.A1(new_n863), .A2(KEYINPUT120), .ZN(new_n864));
  OAI21_X1  g678(.A(new_n789), .B1(new_n861), .B2(new_n862), .ZN(new_n865));
  INV_X1    g679(.A(KEYINPUT53), .ZN(new_n866));
  NAND2_X1  g680(.A1(new_n865), .A2(new_n866), .ZN(new_n867));
  INV_X1    g681(.A(KEYINPUT120), .ZN(new_n868));
  NAND3_X1  g682(.A1(new_n821), .A2(new_n868), .A3(new_n822), .ZN(new_n869));
  NAND3_X1  g683(.A1(new_n864), .A2(new_n867), .A3(new_n869), .ZN(new_n870));
  AOI211_X1 g684(.A(new_n824), .B(new_n859), .C1(KEYINPUT54), .C2(new_n870), .ZN(new_n871));
  NOR2_X1   g685(.A1(G952), .A2(G953), .ZN(new_n872));
  OAI21_X1  g686(.A(new_n776), .B1(new_n871), .B2(new_n872), .ZN(G75));
  NAND2_X1  g687(.A1(new_n596), .A2(new_n458), .ZN(new_n874));
  NAND2_X1  g688(.A1(new_n874), .A2(new_n460), .ZN(new_n875));
  XNOR2_X1  g689(.A(new_n875), .B(KEYINPUT55), .ZN(new_n876));
  INV_X1    g690(.A(new_n876), .ZN(new_n877));
  OAI21_X1  g691(.A(new_n860), .B1(new_n861), .B2(new_n862), .ZN(new_n878));
  INV_X1    g692(.A(new_n822), .ZN(new_n879));
  NAND2_X1  g693(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  AOI21_X1  g694(.A(new_n268), .B1(new_n880), .B2(new_n809), .ZN(new_n881));
  NAND2_X1  g695(.A1(new_n881), .A2(G210), .ZN(new_n882));
  INV_X1    g696(.A(KEYINPUT56), .ZN(new_n883));
  AOI21_X1  g697(.A(new_n877), .B1(new_n882), .B2(new_n883), .ZN(new_n884));
  AOI211_X1 g698(.A(KEYINPUT56), .B(new_n876), .C1(new_n881), .C2(G210), .ZN(new_n885));
  NOR2_X1   g699(.A1(new_n207), .A2(G952), .ZN(new_n886));
  NOR3_X1   g700(.A1(new_n884), .A2(new_n885), .A3(new_n886), .ZN(G51));
  XOR2_X1   g701(.A(new_n752), .B(KEYINPUT57), .Z(new_n888));
  AOI21_X1  g702(.A(new_n810), .B1(new_n880), .B2(new_n809), .ZN(new_n889));
  OAI21_X1  g703(.A(new_n888), .B1(new_n889), .B2(new_n824), .ZN(new_n890));
  NOR2_X1   g704(.A1(new_n423), .A2(new_n424), .ZN(new_n891));
  XOR2_X1   g705(.A(new_n891), .B(KEYINPUT122), .Z(new_n892));
  NAND2_X1  g706(.A1(new_n890), .A2(new_n892), .ZN(new_n893));
  NAND4_X1  g707(.A1(new_n881), .A2(G469), .A3(new_n749), .A4(new_n750), .ZN(new_n894));
  AOI21_X1  g708(.A(new_n886), .B1(new_n893), .B2(new_n894), .ZN(G54));
  NAND3_X1  g709(.A1(new_n881), .A2(KEYINPUT58), .A3(G475), .ZN(new_n896));
  AND2_X1   g710(.A1(new_n896), .A2(new_n261), .ZN(new_n897));
  NOR2_X1   g711(.A1(new_n896), .A2(new_n261), .ZN(new_n898));
  NOR3_X1   g712(.A1(new_n897), .A2(new_n898), .A3(new_n886), .ZN(G60));
  NAND2_X1  g713(.A1(G478), .A2(G902), .ZN(new_n900));
  XOR2_X1   g714(.A(new_n900), .B(KEYINPUT59), .Z(new_n901));
  NOR2_X1   g715(.A1(new_n588), .A2(new_n901), .ZN(new_n902));
  OAI21_X1  g716(.A(new_n902), .B1(new_n889), .B2(new_n824), .ZN(new_n903));
  INV_X1    g717(.A(new_n886), .ZN(new_n904));
  NAND2_X1  g718(.A1(new_n903), .A2(new_n904), .ZN(new_n905));
  NAND2_X1  g719(.A1(new_n870), .A2(KEYINPUT54), .ZN(new_n906));
  NAND2_X1  g720(.A1(new_n906), .A2(new_n823), .ZN(new_n907));
  INV_X1    g721(.A(new_n901), .ZN(new_n908));
  NAND2_X1  g722(.A1(new_n907), .A2(new_n908), .ZN(new_n909));
  AOI21_X1  g723(.A(new_n905), .B1(new_n909), .B2(new_n588), .ZN(G63));
  XNOR2_X1  g724(.A(KEYINPUT123), .B(KEYINPUT60), .ZN(new_n911));
  NOR2_X1   g725(.A1(new_n575), .A2(new_n268), .ZN(new_n912));
  XNOR2_X1  g726(.A(new_n911), .B(new_n912), .ZN(new_n913));
  NOR2_X1   g727(.A1(new_n821), .A2(new_n822), .ZN(new_n914));
  INV_X1    g728(.A(new_n809), .ZN(new_n915));
  OAI211_X1 g729(.A(new_n637), .B(new_n913), .C1(new_n914), .C2(new_n915), .ZN(new_n916));
  INV_X1    g730(.A(new_n913), .ZN(new_n917));
  AOI21_X1  g731(.A(new_n917), .B1(new_n880), .B2(new_n809), .ZN(new_n918));
  OAI211_X1 g732(.A(new_n916), .B(new_n904), .C1(new_n918), .C2(new_n580), .ZN(new_n919));
  INV_X1    g733(.A(KEYINPUT61), .ZN(new_n920));
  XNOR2_X1  g734(.A(new_n919), .B(new_n920), .ZN(G66));
  AOI21_X1  g735(.A(new_n207), .B1(new_n313), .B2(G224), .ZN(new_n922));
  AOI21_X1  g736(.A(new_n922), .B1(new_n799), .B2(new_n207), .ZN(new_n923));
  OAI21_X1  g737(.A(new_n596), .B1(G898), .B2(new_n207), .ZN(new_n924));
  XOR2_X1   g738(.A(new_n923), .B(new_n924), .Z(G69));
  NAND3_X1  g739(.A1(new_n785), .A2(new_n669), .A3(new_n786), .ZN(new_n926));
  INV_X1    g740(.A(KEYINPUT62), .ZN(new_n927));
  XNOR2_X1  g741(.A(new_n926), .B(new_n927), .ZN(new_n928));
  AND2_X1   g742(.A1(new_n762), .A2(new_n769), .ZN(new_n929));
  OR2_X1    g743(.A1(new_n797), .A2(new_n592), .ZN(new_n930));
  NAND4_X1  g744(.A1(new_n930), .A2(new_n675), .A3(new_n666), .A4(new_n747), .ZN(new_n931));
  NAND3_X1  g745(.A1(new_n928), .A2(new_n929), .A3(new_n931), .ZN(new_n932));
  NAND2_X1  g746(.A1(new_n932), .A2(new_n207), .ZN(new_n933));
  XNOR2_X1  g747(.A(new_n499), .B(KEYINPUT124), .ZN(new_n934));
  OAI21_X1  g748(.A(new_n254), .B1(new_n231), .B2(new_n253), .ZN(new_n935));
  XNOR2_X1  g749(.A(new_n934), .B(new_n935), .ZN(new_n936));
  NAND2_X1  g750(.A1(new_n933), .A2(new_n936), .ZN(new_n937));
  NAND2_X1  g751(.A1(new_n937), .A2(KEYINPUT125), .ZN(new_n938));
  INV_X1    g752(.A(KEYINPUT125), .ZN(new_n939));
  NAND3_X1  g753(.A1(new_n933), .A2(new_n939), .A3(new_n936), .ZN(new_n940));
  AOI21_X1  g754(.A(new_n207), .B1(G227), .B2(G900), .ZN(new_n941));
  INV_X1    g755(.A(new_n941), .ZN(new_n942));
  AND2_X1   g756(.A1(new_n761), .A2(new_n724), .ZN(new_n943));
  AND3_X1   g757(.A1(new_n737), .A2(new_n601), .A3(new_n308), .ZN(new_n944));
  AOI21_X1  g758(.A(new_n732), .B1(new_n943), .B2(new_n944), .ZN(new_n945));
  AND3_X1   g759(.A1(new_n945), .A2(new_n769), .A3(new_n729), .ZN(new_n946));
  AND2_X1   g760(.A1(new_n785), .A2(new_n786), .ZN(new_n947));
  INV_X1    g761(.A(KEYINPUT126), .ZN(new_n948));
  AND3_X1   g762(.A1(new_n762), .A2(new_n947), .A3(new_n948), .ZN(new_n949));
  AOI21_X1  g763(.A(new_n948), .B1(new_n762), .B2(new_n947), .ZN(new_n950));
  OAI211_X1 g764(.A(new_n946), .B(new_n207), .C1(new_n949), .C2(new_n950), .ZN(new_n951));
  INV_X1    g765(.A(new_n936), .ZN(new_n952));
  NAND2_X1  g766(.A1(G900), .A2(G953), .ZN(new_n953));
  NAND3_X1  g767(.A1(new_n951), .A2(new_n952), .A3(new_n953), .ZN(new_n954));
  NAND4_X1  g768(.A1(new_n938), .A2(new_n940), .A3(new_n942), .A4(new_n954), .ZN(new_n955));
  INV_X1    g769(.A(KEYINPUT127), .ZN(new_n956));
  NAND2_X1  g770(.A1(new_n954), .A2(new_n956), .ZN(new_n957));
  NAND4_X1  g771(.A1(new_n951), .A2(KEYINPUT127), .A3(new_n952), .A4(new_n953), .ZN(new_n958));
  AND3_X1   g772(.A1(new_n957), .A2(new_n937), .A3(new_n958), .ZN(new_n959));
  OAI21_X1  g773(.A(new_n955), .B1(new_n959), .B2(new_n942), .ZN(G72));
  NAND2_X1  g774(.A1(G472), .A2(G902), .ZN(new_n961));
  XOR2_X1   g775(.A(new_n961), .B(KEYINPUT63), .Z(new_n962));
  INV_X1    g776(.A(new_n534), .ZN(new_n963));
  OAI21_X1  g777(.A(new_n493), .B1(new_n963), .B2(new_n489), .ZN(new_n964));
  AND4_X1   g778(.A1(new_n535), .A2(new_n870), .A3(new_n962), .A4(new_n964), .ZN(new_n965));
  OAI211_X1 g779(.A(new_n946), .B(new_n816), .C1(new_n949), .C2(new_n950), .ZN(new_n966));
  AOI21_X1  g780(.A(new_n535), .B1(new_n966), .B2(new_n962), .ZN(new_n967));
  NAND4_X1  g781(.A1(new_n928), .A2(new_n816), .A3(new_n929), .A4(new_n931), .ZN(new_n968));
  AOI21_X1  g782(.A(new_n964), .B1(new_n968), .B2(new_n962), .ZN(new_n969));
  NOR4_X1   g783(.A1(new_n965), .A2(new_n886), .A3(new_n967), .A4(new_n969), .ZN(G57));
endmodule


