//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 0 1 1 1 1 0 0 0 1 0 0 0 1 0 0 0 1 1 1 0 1 0 1 1 1 0 1 1 1 1 0 1 0 0 0 1 0 1 1 1 0 1 0 0 1 0 1 1 0 1 0 1 1 1 0 0 1 0 0 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:27:30 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n635, new_n636, new_n637,
    new_n638, new_n639, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n653, new_n654, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n690, new_n691, new_n692, new_n693, new_n694, new_n695, new_n696,
    new_n697, new_n698, new_n699, new_n700, new_n701, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n710, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n721,
    new_n722, new_n723, new_n724, new_n725, new_n726, new_n728, new_n729,
    new_n730, new_n731, new_n732, new_n733, new_n734, new_n735, new_n736,
    new_n737, new_n738, new_n739, new_n740, new_n741, new_n742, new_n743,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n760, new_n761, new_n762, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n783, new_n784, new_n785, new_n786, new_n787, new_n788, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n897, new_n898,
    new_n899, new_n900, new_n902, new_n903, new_n904, new_n905, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n916, new_n917, new_n918, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n954, new_n955, new_n956, new_n957, new_n958, new_n959,
    new_n960, new_n961, new_n962, new_n963;
  INV_X1    g000(.A(KEYINPUT11), .ZN(new_n187));
  NOR2_X1   g001(.A1(new_n187), .A2(KEYINPUT64), .ZN(new_n188));
  INV_X1    g002(.A(G134), .ZN(new_n189));
  NOR2_X1   g003(.A1(new_n189), .A2(G137), .ZN(new_n190));
  NAND2_X1  g004(.A1(new_n187), .A2(KEYINPUT64), .ZN(new_n191));
  AOI21_X1  g005(.A(new_n188), .B1(new_n190), .B2(new_n191), .ZN(new_n192));
  INV_X1    g006(.A(KEYINPUT64), .ZN(new_n193));
  INV_X1    g007(.A(G137), .ZN(new_n194));
  NAND4_X1  g008(.A1(new_n193), .A2(new_n194), .A3(KEYINPUT11), .A4(G134), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n189), .A2(G137), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n195), .A2(new_n196), .ZN(new_n197));
  NOR3_X1   g011(.A1(new_n192), .A2(new_n197), .A3(G131), .ZN(new_n198));
  INV_X1    g012(.A(G131), .ZN(new_n199));
  NOR2_X1   g013(.A1(new_n194), .A2(G134), .ZN(new_n200));
  AOI21_X1  g014(.A(new_n200), .B1(new_n188), .B2(new_n190), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n193), .A2(KEYINPUT11), .ZN(new_n202));
  NOR2_X1   g016(.A1(new_n193), .A2(KEYINPUT11), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n194), .A2(G134), .ZN(new_n204));
  OAI21_X1  g018(.A(new_n202), .B1(new_n203), .B2(new_n204), .ZN(new_n205));
  AOI21_X1  g019(.A(new_n199), .B1(new_n201), .B2(new_n205), .ZN(new_n206));
  NOR2_X1   g020(.A1(new_n198), .A2(new_n206), .ZN(new_n207));
  INV_X1    g021(.A(new_n207), .ZN(new_n208));
  INV_X1    g022(.A(KEYINPUT10), .ZN(new_n209));
  INV_X1    g023(.A(G107), .ZN(new_n210));
  NAND3_X1  g024(.A1(new_n210), .A2(KEYINPUT78), .A3(G104), .ZN(new_n211));
  INV_X1    g025(.A(G104), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n212), .A2(G107), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n211), .A2(new_n213), .ZN(new_n214));
  AOI21_X1  g028(.A(KEYINPUT78), .B1(new_n210), .B2(G104), .ZN(new_n215));
  OAI21_X1  g029(.A(G101), .B1(new_n214), .B2(new_n215), .ZN(new_n216));
  OAI21_X1  g030(.A(KEYINPUT3), .B1(new_n212), .B2(G107), .ZN(new_n217));
  INV_X1    g031(.A(KEYINPUT3), .ZN(new_n218));
  NAND3_X1  g032(.A1(new_n218), .A2(new_n210), .A3(G104), .ZN(new_n219));
  INV_X1    g033(.A(G101), .ZN(new_n220));
  NAND4_X1  g034(.A1(new_n217), .A2(new_n219), .A3(new_n220), .A4(new_n213), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n216), .A2(new_n221), .ZN(new_n222));
  INV_X1    g036(.A(KEYINPUT1), .ZN(new_n223));
  INV_X1    g037(.A(G146), .ZN(new_n224));
  NAND2_X1  g038(.A1(new_n224), .A2(G143), .ZN(new_n225));
  INV_X1    g039(.A(G143), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n226), .A2(G146), .ZN(new_n227));
  AND4_X1   g041(.A1(new_n223), .A2(new_n225), .A3(new_n227), .A4(G128), .ZN(new_n228));
  OAI21_X1  g042(.A(KEYINPUT1), .B1(new_n226), .B2(G146), .ZN(new_n229));
  AOI22_X1  g043(.A1(new_n229), .A2(G128), .B1(new_n225), .B2(new_n227), .ZN(new_n230));
  NOR2_X1   g044(.A1(new_n228), .A2(new_n230), .ZN(new_n231));
  OAI21_X1  g045(.A(new_n209), .B1(new_n222), .B2(new_n231), .ZN(new_n232));
  NAND3_X1  g046(.A1(new_n217), .A2(new_n219), .A3(new_n213), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n233), .A2(G101), .ZN(new_n234));
  NAND3_X1  g048(.A1(new_n234), .A2(KEYINPUT4), .A3(new_n221), .ZN(new_n235));
  NOR2_X1   g049(.A1(KEYINPUT0), .A2(G128), .ZN(new_n236));
  XNOR2_X1  g050(.A(G143), .B(G146), .ZN(new_n237));
  NAND2_X1  g051(.A1(KEYINPUT0), .A2(G128), .ZN(new_n238));
  AOI21_X1  g052(.A(new_n236), .B1(new_n237), .B2(new_n238), .ZN(new_n239));
  OAI21_X1  g053(.A(new_n239), .B1(new_n237), .B2(new_n238), .ZN(new_n240));
  INV_X1    g054(.A(KEYINPUT4), .ZN(new_n241));
  NAND3_X1  g055(.A1(new_n233), .A2(new_n241), .A3(G101), .ZN(new_n242));
  NAND3_X1  g056(.A1(new_n235), .A2(new_n240), .A3(new_n242), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n232), .A2(new_n243), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n229), .A2(G128), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n225), .A2(new_n227), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n245), .A2(new_n246), .ZN(new_n247));
  NAND3_X1  g061(.A1(new_n237), .A2(G128), .A3(new_n229), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n247), .A2(new_n248), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n249), .A2(KEYINPUT10), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n222), .A2(KEYINPUT79), .ZN(new_n251));
  INV_X1    g065(.A(KEYINPUT79), .ZN(new_n252));
  NAND3_X1  g066(.A1(new_n216), .A2(new_n252), .A3(new_n221), .ZN(new_n253));
  AOI21_X1  g067(.A(new_n250), .B1(new_n251), .B2(new_n253), .ZN(new_n254));
  OAI21_X1  g068(.A(new_n208), .B1(new_n244), .B2(new_n254), .ZN(new_n255));
  AND3_X1   g069(.A1(new_n216), .A2(new_n252), .A3(new_n221), .ZN(new_n256));
  AOI21_X1  g070(.A(new_n252), .B1(new_n216), .B2(new_n221), .ZN(new_n257));
  OAI211_X1 g071(.A(KEYINPUT10), .B(new_n249), .C1(new_n256), .C2(new_n257), .ZN(new_n258));
  NAND4_X1  g072(.A1(new_n258), .A2(new_n207), .A3(new_n232), .A4(new_n243), .ZN(new_n259));
  INV_X1    g073(.A(KEYINPUT80), .ZN(new_n260));
  NAND3_X1  g074(.A1(new_n255), .A2(new_n259), .A3(new_n260), .ZN(new_n261));
  OAI211_X1 g075(.A(KEYINPUT80), .B(new_n208), .C1(new_n244), .C2(new_n254), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n261), .A2(new_n262), .ZN(new_n263));
  XNOR2_X1  g077(.A(G110), .B(G140), .ZN(new_n264));
  INV_X1    g078(.A(G227), .ZN(new_n265));
  NOR2_X1   g079(.A1(new_n265), .A2(G953), .ZN(new_n266));
  XNOR2_X1  g080(.A(new_n264), .B(new_n266), .ZN(new_n267));
  INV_X1    g081(.A(new_n267), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n263), .A2(new_n268), .ZN(new_n269));
  NOR3_X1   g083(.A1(new_n256), .A2(new_n257), .A3(new_n249), .ZN(new_n270));
  NOR2_X1   g084(.A1(new_n222), .A2(new_n231), .ZN(new_n271));
  OAI21_X1  g085(.A(new_n208), .B1(new_n270), .B2(new_n271), .ZN(new_n272));
  NAND2_X1  g086(.A1(new_n272), .A2(KEYINPUT12), .ZN(new_n273));
  INV_X1    g087(.A(KEYINPUT12), .ZN(new_n274));
  OAI211_X1 g088(.A(new_n274), .B(new_n208), .C1(new_n270), .C2(new_n271), .ZN(new_n275));
  NAND3_X1  g089(.A1(new_n273), .A2(new_n275), .A3(new_n259), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n276), .A2(new_n267), .ZN(new_n277));
  AOI21_X1  g091(.A(G902), .B1(new_n269), .B2(new_n277), .ZN(new_n278));
  INV_X1    g092(.A(new_n278), .ZN(new_n279));
  INV_X1    g093(.A(KEYINPUT81), .ZN(new_n280));
  NAND3_X1  g094(.A1(new_n279), .A2(new_n280), .A3(G469), .ZN(new_n281));
  INV_X1    g095(.A(G469), .ZN(new_n282));
  OAI21_X1  g096(.A(KEYINPUT81), .B1(new_n278), .B2(new_n282), .ZN(new_n283));
  NAND3_X1  g097(.A1(new_n261), .A2(new_n267), .A3(new_n262), .ZN(new_n284));
  NAND4_X1  g098(.A1(new_n273), .A2(new_n275), .A3(new_n259), .A4(new_n268), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n284), .A2(new_n285), .ZN(new_n286));
  INV_X1    g100(.A(G902), .ZN(new_n287));
  NAND3_X1  g101(.A1(new_n286), .A2(new_n282), .A3(new_n287), .ZN(new_n288));
  NAND3_X1  g102(.A1(new_n281), .A2(new_n283), .A3(new_n288), .ZN(new_n289));
  XOR2_X1   g103(.A(KEYINPUT9), .B(G234), .Z(new_n290));
  XNOR2_X1  g104(.A(new_n290), .B(KEYINPUT76), .ZN(new_n291));
  OAI21_X1  g105(.A(G221), .B1(new_n291), .B2(G902), .ZN(new_n292));
  XNOR2_X1  g106(.A(new_n292), .B(KEYINPUT77), .ZN(new_n293));
  INV_X1    g107(.A(new_n293), .ZN(new_n294));
  AND2_X1   g108(.A1(new_n289), .A2(new_n294), .ZN(new_n295));
  INV_X1    g109(.A(KEYINPUT89), .ZN(new_n296));
  INV_X1    g110(.A(G953), .ZN(new_n297));
  INV_X1    g111(.A(KEYINPUT68), .ZN(new_n298));
  NOR2_X1   g112(.A1(new_n298), .A2(G237), .ZN(new_n299));
  INV_X1    g113(.A(G237), .ZN(new_n300));
  NOR2_X1   g114(.A1(new_n300), .A2(KEYINPUT68), .ZN(new_n301));
  OAI211_X1 g115(.A(G214), .B(new_n297), .C1(new_n299), .C2(new_n301), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n302), .A2(new_n226), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n300), .A2(KEYINPUT68), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n298), .A2(G237), .ZN(new_n305));
  AOI21_X1  g119(.A(G953), .B1(new_n304), .B2(new_n305), .ZN(new_n306));
  NAND3_X1  g120(.A1(new_n306), .A2(G143), .A3(G214), .ZN(new_n307));
  NAND2_X1  g121(.A1(KEYINPUT18), .A2(G131), .ZN(new_n308));
  NAND3_X1  g122(.A1(new_n303), .A2(new_n307), .A3(new_n308), .ZN(new_n309));
  INV_X1    g123(.A(KEYINPUT85), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n309), .A2(new_n310), .ZN(new_n311));
  NAND4_X1  g125(.A1(new_n303), .A2(KEYINPUT85), .A3(new_n307), .A4(new_n308), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n311), .A2(new_n312), .ZN(new_n313));
  NAND2_X1  g127(.A1(new_n303), .A2(new_n307), .ZN(new_n314));
  INV_X1    g128(.A(new_n308), .ZN(new_n315));
  INV_X1    g129(.A(G140), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n316), .A2(G125), .ZN(new_n317));
  INV_X1    g131(.A(G125), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n318), .A2(G140), .ZN(new_n319));
  INV_X1    g133(.A(KEYINPUT73), .ZN(new_n320));
  NAND3_X1  g134(.A1(new_n317), .A2(new_n319), .A3(new_n320), .ZN(new_n321));
  NAND3_X1  g135(.A1(new_n318), .A2(KEYINPUT73), .A3(G140), .ZN(new_n322));
  AND2_X1   g136(.A1(new_n321), .A2(new_n322), .ZN(new_n323));
  NAND2_X1  g137(.A1(new_n323), .A2(G146), .ZN(new_n324));
  NAND3_X1  g138(.A1(new_n317), .A2(new_n319), .A3(new_n224), .ZN(new_n325));
  AOI22_X1  g139(.A1(new_n314), .A2(new_n315), .B1(new_n324), .B2(new_n325), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n313), .A2(new_n326), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n304), .A2(new_n305), .ZN(new_n328));
  AND4_X1   g142(.A1(G143), .A2(new_n328), .A3(G214), .A4(new_n297), .ZN(new_n329));
  AOI21_X1  g143(.A(G143), .B1(new_n306), .B2(G214), .ZN(new_n330));
  OAI21_X1  g144(.A(G131), .B1(new_n329), .B2(new_n330), .ZN(new_n331));
  INV_X1    g145(.A(KEYINPUT17), .ZN(new_n332));
  NAND3_X1  g146(.A1(new_n303), .A2(new_n199), .A3(new_n307), .ZN(new_n333));
  NAND3_X1  g147(.A1(new_n331), .A2(new_n332), .A3(new_n333), .ZN(new_n334));
  NAND3_X1  g148(.A1(new_n321), .A2(KEYINPUT16), .A3(new_n322), .ZN(new_n335));
  INV_X1    g149(.A(KEYINPUT16), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n317), .A2(new_n336), .ZN(new_n337));
  AND3_X1   g151(.A1(new_n335), .A2(new_n224), .A3(new_n337), .ZN(new_n338));
  AOI21_X1  g152(.A(new_n224), .B1(new_n335), .B2(new_n337), .ZN(new_n339));
  NOR2_X1   g153(.A1(new_n338), .A2(new_n339), .ZN(new_n340));
  OAI211_X1 g154(.A(KEYINPUT17), .B(G131), .C1(new_n329), .C2(new_n330), .ZN(new_n341));
  NAND3_X1  g155(.A1(new_n334), .A2(new_n340), .A3(new_n341), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n327), .A2(new_n342), .ZN(new_n343));
  XNOR2_X1  g157(.A(G113), .B(G122), .ZN(new_n344));
  XNOR2_X1  g158(.A(new_n344), .B(new_n212), .ZN(new_n345));
  INV_X1    g159(.A(new_n345), .ZN(new_n346));
  NOR2_X1   g160(.A1(new_n343), .A2(new_n346), .ZN(new_n347));
  NAND3_X1  g161(.A1(new_n335), .A2(new_n224), .A3(new_n337), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n335), .A2(new_n337), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n349), .A2(G146), .ZN(new_n350));
  AND3_X1   g164(.A1(new_n341), .A2(new_n348), .A3(new_n350), .ZN(new_n351));
  AOI22_X1  g165(.A1(new_n351), .A2(new_n334), .B1(new_n313), .B2(new_n326), .ZN(new_n352));
  OAI21_X1  g166(.A(KEYINPUT88), .B1(new_n352), .B2(new_n345), .ZN(new_n353));
  INV_X1    g167(.A(KEYINPUT88), .ZN(new_n354));
  NAND3_X1  g168(.A1(new_n343), .A2(new_n354), .A3(new_n346), .ZN(new_n355));
  AOI21_X1  g169(.A(new_n347), .B1(new_n353), .B2(new_n355), .ZN(new_n356));
  OAI21_X1  g170(.A(new_n296), .B1(new_n356), .B2(G902), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n352), .A2(new_n345), .ZN(new_n358));
  AOI21_X1  g172(.A(new_n354), .B1(new_n343), .B2(new_n346), .ZN(new_n359));
  AOI211_X1 g173(.A(KEYINPUT88), .B(new_n345), .C1(new_n327), .C2(new_n342), .ZN(new_n360));
  OAI21_X1  g174(.A(new_n358), .B1(new_n359), .B2(new_n360), .ZN(new_n361));
  NAND3_X1  g175(.A1(new_n361), .A2(KEYINPUT89), .A3(new_n287), .ZN(new_n362));
  NAND3_X1  g176(.A1(new_n357), .A2(new_n362), .A3(G475), .ZN(new_n363));
  NOR2_X1   g177(.A1(G475), .A2(G902), .ZN(new_n364));
  NAND2_X1  g178(.A1(new_n331), .A2(new_n333), .ZN(new_n365));
  XOR2_X1   g179(.A(KEYINPUT86), .B(KEYINPUT19), .Z(new_n366));
  NAND3_X1  g180(.A1(new_n366), .A2(new_n317), .A3(new_n319), .ZN(new_n367));
  OR2_X1    g181(.A1(new_n367), .A2(KEYINPUT87), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n323), .A2(KEYINPUT19), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n367), .A2(KEYINPUT87), .ZN(new_n370));
  NAND3_X1  g184(.A1(new_n368), .A2(new_n369), .A3(new_n370), .ZN(new_n371));
  OAI211_X1 g185(.A(new_n365), .B(new_n350), .C1(new_n371), .C2(G146), .ZN(new_n372));
  AOI21_X1  g186(.A(new_n345), .B1(new_n372), .B2(new_n327), .ZN(new_n373));
  OAI21_X1  g187(.A(new_n364), .B1(new_n347), .B2(new_n373), .ZN(new_n374));
  XNOR2_X1  g188(.A(new_n374), .B(KEYINPUT20), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n363), .A2(new_n375), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n226), .A2(G128), .ZN(new_n377));
  INV_X1    g191(.A(G128), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n378), .A2(G143), .ZN(new_n379));
  NAND2_X1  g193(.A1(new_n377), .A2(new_n379), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n380), .A2(G134), .ZN(new_n381));
  NAND3_X1  g195(.A1(new_n377), .A2(new_n379), .A3(new_n189), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n381), .A2(new_n382), .ZN(new_n383));
  INV_X1    g197(.A(G122), .ZN(new_n384));
  OAI21_X1  g198(.A(KEYINPUT14), .B1(new_n384), .B2(G116), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n384), .A2(G116), .ZN(new_n386));
  NAND2_X1  g200(.A1(new_n385), .A2(new_n386), .ZN(new_n387));
  NOR3_X1   g201(.A1(new_n384), .A2(KEYINPUT14), .A3(G116), .ZN(new_n388));
  OAI21_X1  g202(.A(G107), .B1(new_n387), .B2(new_n388), .ZN(new_n389));
  NOR2_X1   g203(.A1(new_n384), .A2(G116), .ZN(new_n390));
  INV_X1    g204(.A(G116), .ZN(new_n391));
  NOR2_X1   g205(.A1(new_n391), .A2(G122), .ZN(new_n392));
  NOR2_X1   g206(.A1(new_n390), .A2(new_n392), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n393), .A2(new_n210), .ZN(new_n394));
  NAND3_X1  g208(.A1(new_n383), .A2(new_n389), .A3(new_n394), .ZN(new_n395));
  INV_X1    g209(.A(KEYINPUT90), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n395), .A2(new_n396), .ZN(new_n397));
  OAI21_X1  g211(.A(G107), .B1(new_n390), .B2(new_n392), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n394), .A2(new_n398), .ZN(new_n399));
  INV_X1    g213(.A(KEYINPUT13), .ZN(new_n400));
  OAI21_X1  g214(.A(new_n379), .B1(new_n377), .B2(new_n400), .ZN(new_n401));
  AOI21_X1  g215(.A(KEYINPUT13), .B1(new_n226), .B2(G128), .ZN(new_n402));
  OAI21_X1  g216(.A(G134), .B1(new_n401), .B2(new_n402), .ZN(new_n403));
  NAND3_X1  g217(.A1(new_n399), .A2(new_n382), .A3(new_n403), .ZN(new_n404));
  NAND4_X1  g218(.A1(new_n383), .A2(new_n389), .A3(KEYINPUT90), .A4(new_n394), .ZN(new_n405));
  NAND3_X1  g219(.A1(new_n397), .A2(new_n404), .A3(new_n405), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n297), .A2(G217), .ZN(new_n407));
  OAI21_X1  g221(.A(new_n406), .B1(new_n291), .B2(new_n407), .ZN(new_n408));
  NAND2_X1  g222(.A1(new_n408), .A2(KEYINPUT91), .ZN(new_n409));
  INV_X1    g223(.A(KEYINPUT91), .ZN(new_n410));
  OAI211_X1 g224(.A(new_n406), .B(new_n410), .C1(new_n291), .C2(new_n407), .ZN(new_n411));
  NOR2_X1   g225(.A1(new_n291), .A2(new_n407), .ZN(new_n412));
  NAND4_X1  g226(.A1(new_n397), .A2(new_n412), .A3(new_n405), .A4(new_n404), .ZN(new_n413));
  NAND3_X1  g227(.A1(new_n409), .A2(new_n411), .A3(new_n413), .ZN(new_n414));
  NAND3_X1  g228(.A1(new_n414), .A2(KEYINPUT92), .A3(new_n287), .ZN(new_n415));
  INV_X1    g229(.A(G478), .ZN(new_n416));
  NOR2_X1   g230(.A1(new_n416), .A2(KEYINPUT15), .ZN(new_n417));
  INV_X1    g231(.A(new_n417), .ZN(new_n418));
  XNOR2_X1  g232(.A(new_n415), .B(new_n418), .ZN(new_n419));
  INV_X1    g233(.A(new_n419), .ZN(new_n420));
  NOR2_X1   g234(.A1(new_n376), .A2(new_n420), .ZN(new_n421));
  AND2_X1   g235(.A1(new_n297), .A2(G952), .ZN(new_n422));
  NAND2_X1  g236(.A1(G234), .A2(G237), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n422), .A2(new_n423), .ZN(new_n424));
  XNOR2_X1  g238(.A(new_n424), .B(KEYINPUT93), .ZN(new_n425));
  XNOR2_X1  g239(.A(KEYINPUT21), .B(G898), .ZN(new_n426));
  INV_X1    g240(.A(new_n426), .ZN(new_n427));
  NAND3_X1  g241(.A1(new_n423), .A2(G902), .A3(G953), .ZN(new_n428));
  OAI21_X1  g242(.A(new_n425), .B1(new_n427), .B2(new_n428), .ZN(new_n429));
  OAI21_X1  g243(.A(G214), .B1(G237), .B2(G902), .ZN(new_n430));
  INV_X1    g244(.A(new_n430), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n240), .A2(G125), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n249), .A2(new_n318), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n432), .A2(new_n433), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n297), .A2(G224), .ZN(new_n435));
  XNOR2_X1  g249(.A(new_n435), .B(KEYINPUT84), .ZN(new_n436));
  NAND2_X1  g250(.A1(new_n436), .A2(KEYINPUT7), .ZN(new_n437));
  INV_X1    g251(.A(new_n437), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n434), .A2(new_n438), .ZN(new_n439));
  NAND3_X1  g253(.A1(new_n432), .A2(new_n433), .A3(new_n437), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n439), .A2(new_n440), .ZN(new_n441));
  INV_X1    g255(.A(G119), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n442), .A2(G116), .ZN(new_n443));
  OAI21_X1  g257(.A(G113), .B1(new_n443), .B2(KEYINPUT5), .ZN(new_n444));
  OAI21_X1  g258(.A(KEYINPUT65), .B1(new_n442), .B2(G116), .ZN(new_n445));
  INV_X1    g259(.A(KEYINPUT65), .ZN(new_n446));
  NAND3_X1  g260(.A1(new_n446), .A2(new_n391), .A3(G119), .ZN(new_n447));
  AOI22_X1  g261(.A1(new_n445), .A2(new_n447), .B1(G116), .B2(new_n442), .ZN(new_n448));
  AOI21_X1  g262(.A(new_n444), .B1(new_n448), .B2(KEYINPUT5), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n445), .A2(new_n447), .ZN(new_n450));
  INV_X1    g264(.A(G113), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n451), .A2(KEYINPUT2), .ZN(new_n452));
  INV_X1    g266(.A(KEYINPUT2), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n453), .A2(G113), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n452), .A2(new_n454), .ZN(new_n455));
  AND3_X1   g269(.A1(new_n450), .A2(new_n443), .A3(new_n455), .ZN(new_n456));
  NOR2_X1   g270(.A1(new_n449), .A2(new_n456), .ZN(new_n457));
  OAI21_X1  g271(.A(new_n457), .B1(new_n256), .B2(new_n257), .ZN(new_n458));
  OAI21_X1  g272(.A(new_n222), .B1(new_n449), .B2(new_n456), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  XNOR2_X1  g274(.A(G110), .B(G122), .ZN(new_n461));
  XNOR2_X1  g275(.A(new_n461), .B(KEYINPUT8), .ZN(new_n462));
  AOI21_X1  g276(.A(new_n441), .B1(new_n460), .B2(new_n462), .ZN(new_n463));
  AOI21_X1  g277(.A(new_n455), .B1(new_n450), .B2(new_n443), .ZN(new_n464));
  INV_X1    g278(.A(KEYINPUT66), .ZN(new_n465));
  NOR3_X1   g279(.A1(new_n456), .A2(new_n464), .A3(new_n465), .ZN(new_n466));
  AOI21_X1  g280(.A(new_n446), .B1(new_n391), .B2(G119), .ZN(new_n467));
  NOR3_X1   g281(.A1(new_n442), .A2(KEYINPUT65), .A3(G116), .ZN(new_n468));
  OAI21_X1  g282(.A(new_n443), .B1(new_n467), .B2(new_n468), .ZN(new_n469));
  INV_X1    g283(.A(new_n455), .ZN(new_n470));
  NAND2_X1  g284(.A1(new_n469), .A2(new_n470), .ZN(new_n471));
  NAND2_X1  g285(.A1(new_n448), .A2(new_n455), .ZN(new_n472));
  AOI21_X1  g286(.A(KEYINPUT66), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  NOR2_X1   g287(.A1(new_n466), .A2(new_n473), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n235), .A2(new_n242), .ZN(new_n475));
  OAI211_X1 g289(.A(new_n461), .B(new_n458), .C1(new_n474), .C2(new_n475), .ZN(new_n476));
  AOI21_X1  g290(.A(G902), .B1(new_n463), .B2(new_n476), .ZN(new_n477));
  INV_X1    g291(.A(new_n461), .ZN(new_n478));
  INV_X1    g292(.A(new_n458), .ZN(new_n479));
  OAI21_X1  g293(.A(new_n465), .B1(new_n456), .B2(new_n464), .ZN(new_n480));
  NAND3_X1  g294(.A1(new_n471), .A2(new_n472), .A3(KEYINPUT66), .ZN(new_n481));
  AOI21_X1  g295(.A(new_n475), .B1(new_n480), .B2(new_n481), .ZN(new_n482));
  OAI21_X1  g296(.A(new_n478), .B1(new_n479), .B2(new_n482), .ZN(new_n483));
  INV_X1    g297(.A(KEYINPUT82), .ZN(new_n484));
  INV_X1    g298(.A(KEYINPUT6), .ZN(new_n485));
  NOR2_X1   g299(.A1(new_n484), .A2(new_n485), .ZN(new_n486));
  NAND3_X1  g300(.A1(new_n483), .A2(new_n476), .A3(new_n486), .ZN(new_n487));
  XNOR2_X1  g301(.A(new_n436), .B(KEYINPUT83), .ZN(new_n488));
  XNOR2_X1  g302(.A(new_n434), .B(new_n488), .ZN(new_n489));
  OAI221_X1 g303(.A(new_n478), .B1(new_n484), .B2(new_n485), .C1(new_n479), .C2(new_n482), .ZN(new_n490));
  NAND3_X1  g304(.A1(new_n487), .A2(new_n489), .A3(new_n490), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n477), .A2(new_n491), .ZN(new_n492));
  OAI21_X1  g306(.A(G210), .B1(G237), .B2(G902), .ZN(new_n493));
  INV_X1    g307(.A(new_n493), .ZN(new_n494));
  NAND2_X1  g308(.A1(new_n492), .A2(new_n494), .ZN(new_n495));
  NAND3_X1  g309(.A1(new_n477), .A2(new_n491), .A3(new_n493), .ZN(new_n496));
  AOI21_X1  g310(.A(new_n431), .B1(new_n495), .B2(new_n496), .ZN(new_n497));
  AND4_X1   g311(.A1(new_n295), .A2(new_n421), .A3(new_n429), .A4(new_n497), .ZN(new_n498));
  NOR2_X1   g312(.A1(G472), .A2(G902), .ZN(new_n499));
  INV_X1    g313(.A(new_n474), .ZN(new_n500));
  OAI21_X1  g314(.A(new_n240), .B1(new_n198), .B2(new_n206), .ZN(new_n501));
  INV_X1    g315(.A(KEYINPUT30), .ZN(new_n502));
  NAND3_X1  g316(.A1(new_n201), .A2(new_n199), .A3(new_n205), .ZN(new_n503));
  OAI21_X1  g317(.A(G131), .B1(new_n190), .B2(new_n200), .ZN(new_n504));
  NAND3_X1  g318(.A1(new_n249), .A2(new_n503), .A3(new_n504), .ZN(new_n505));
  AND3_X1   g319(.A1(new_n501), .A2(new_n502), .A3(new_n505), .ZN(new_n506));
  AOI21_X1  g320(.A(new_n502), .B1(new_n501), .B2(new_n505), .ZN(new_n507));
  OAI21_X1  g321(.A(new_n500), .B1(new_n506), .B2(new_n507), .ZN(new_n508));
  AND2_X1   g322(.A1(new_n501), .A2(new_n505), .ZN(new_n509));
  AND3_X1   g323(.A1(new_n480), .A2(KEYINPUT67), .A3(new_n481), .ZN(new_n510));
  AOI21_X1  g324(.A(KEYINPUT67), .B1(new_n480), .B2(new_n481), .ZN(new_n511));
  OAI21_X1  g325(.A(new_n509), .B1(new_n510), .B2(new_n511), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n306), .A2(G210), .ZN(new_n513));
  XNOR2_X1  g327(.A(KEYINPUT69), .B(KEYINPUT27), .ZN(new_n514));
  XNOR2_X1  g328(.A(new_n513), .B(new_n514), .ZN(new_n515));
  XNOR2_X1  g329(.A(KEYINPUT26), .B(G101), .ZN(new_n516));
  XNOR2_X1  g330(.A(new_n515), .B(new_n516), .ZN(new_n517));
  NAND3_X1  g331(.A1(new_n508), .A2(new_n512), .A3(new_n517), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n518), .A2(KEYINPUT31), .ZN(new_n519));
  INV_X1    g333(.A(KEYINPUT31), .ZN(new_n520));
  NAND4_X1  g334(.A1(new_n508), .A2(new_n520), .A3(new_n512), .A4(new_n517), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n519), .A2(new_n521), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n501), .A2(new_n505), .ZN(new_n523));
  INV_X1    g337(.A(KEYINPUT67), .ZN(new_n524));
  OAI21_X1  g338(.A(new_n524), .B1(new_n466), .B2(new_n473), .ZN(new_n525));
  NAND3_X1  g339(.A1(new_n480), .A2(new_n481), .A3(KEYINPUT67), .ZN(new_n526));
  AOI21_X1  g340(.A(new_n523), .B1(new_n525), .B2(new_n526), .ZN(new_n527));
  NOR2_X1   g341(.A1(new_n509), .A2(new_n474), .ZN(new_n528));
  OAI21_X1  g342(.A(KEYINPUT28), .B1(new_n527), .B2(new_n528), .ZN(new_n529));
  INV_X1    g343(.A(KEYINPUT28), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n523), .A2(KEYINPUT70), .ZN(new_n531));
  INV_X1    g345(.A(KEYINPUT70), .ZN(new_n532));
  NAND3_X1  g346(.A1(new_n501), .A2(new_n532), .A3(new_n505), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n531), .A2(new_n533), .ZN(new_n534));
  NOR2_X1   g348(.A1(new_n510), .A2(new_n511), .ZN(new_n535));
  OAI21_X1  g349(.A(new_n530), .B1(new_n534), .B2(new_n535), .ZN(new_n536));
  AOI21_X1  g350(.A(new_n517), .B1(new_n529), .B2(new_n536), .ZN(new_n537));
  OAI21_X1  g351(.A(new_n499), .B1(new_n522), .B2(new_n537), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n538), .A2(KEYINPUT32), .ZN(new_n539));
  INV_X1    g353(.A(KEYINPUT32), .ZN(new_n540));
  OAI211_X1 g354(.A(new_n540), .B(new_n499), .C1(new_n522), .C2(new_n537), .ZN(new_n541));
  INV_X1    g355(.A(new_n533), .ZN(new_n542));
  AOI21_X1  g356(.A(new_n532), .B1(new_n501), .B2(new_n505), .ZN(new_n543));
  NOR2_X1   g357(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  NAND2_X1  g358(.A1(new_n525), .A2(new_n526), .ZN(new_n545));
  AOI21_X1  g359(.A(KEYINPUT28), .B1(new_n544), .B2(new_n545), .ZN(new_n546));
  NAND3_X1  g360(.A1(new_n525), .A2(new_n526), .A3(new_n523), .ZN(new_n547));
  AOI21_X1  g361(.A(new_n530), .B1(new_n512), .B2(new_n547), .ZN(new_n548));
  NOR2_X1   g362(.A1(new_n546), .A2(new_n548), .ZN(new_n549));
  AND2_X1   g363(.A1(new_n517), .A2(KEYINPUT29), .ZN(new_n550));
  AOI21_X1  g364(.A(G902), .B1(new_n549), .B2(new_n550), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n508), .A2(new_n512), .ZN(new_n552));
  NOR2_X1   g366(.A1(new_n552), .A2(new_n517), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n529), .A2(new_n536), .ZN(new_n554));
  AOI21_X1  g368(.A(new_n553), .B1(new_n554), .B2(new_n517), .ZN(new_n555));
  OAI21_X1  g369(.A(new_n551), .B1(new_n555), .B2(KEYINPUT29), .ZN(new_n556));
  AOI22_X1  g370(.A1(new_n539), .A2(new_n541), .B1(new_n556), .B2(G472), .ZN(new_n557));
  INV_X1    g371(.A(G217), .ZN(new_n558));
  AOI21_X1  g372(.A(new_n558), .B1(G234), .B2(new_n287), .ZN(new_n559));
  INV_X1    g373(.A(KEYINPUT25), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n560), .A2(KEYINPUT74), .ZN(new_n561));
  INV_X1    g375(.A(KEYINPUT72), .ZN(new_n562));
  INV_X1    g376(.A(KEYINPUT23), .ZN(new_n563));
  AND4_X1   g377(.A1(new_n562), .A2(new_n563), .A3(new_n378), .A4(G119), .ZN(new_n564));
  OAI21_X1  g378(.A(KEYINPUT23), .B1(new_n378), .B2(G119), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n565), .A2(new_n562), .ZN(new_n566));
  NOR2_X1   g380(.A1(new_n442), .A2(G128), .ZN(new_n567));
  INV_X1    g381(.A(new_n567), .ZN(new_n568));
  AOI21_X1  g382(.A(new_n564), .B1(new_n566), .B2(new_n568), .ZN(new_n569));
  INV_X1    g383(.A(KEYINPUT71), .ZN(new_n570));
  OAI21_X1  g384(.A(new_n570), .B1(new_n378), .B2(G119), .ZN(new_n571));
  NAND3_X1  g385(.A1(new_n442), .A2(KEYINPUT71), .A3(G128), .ZN(new_n572));
  AOI21_X1  g386(.A(new_n567), .B1(new_n571), .B2(new_n572), .ZN(new_n573));
  XNOR2_X1  g387(.A(KEYINPUT24), .B(G110), .ZN(new_n574));
  INV_X1    g388(.A(new_n574), .ZN(new_n575));
  AOI22_X1  g389(.A1(new_n569), .A2(G110), .B1(new_n573), .B2(new_n575), .ZN(new_n576));
  OAI21_X1  g390(.A(new_n576), .B1(new_n338), .B2(new_n339), .ZN(new_n577));
  INV_X1    g391(.A(G110), .ZN(new_n578));
  AOI21_X1  g392(.A(new_n567), .B1(new_n565), .B2(new_n562), .ZN(new_n579));
  OAI21_X1  g393(.A(new_n578), .B1(new_n579), .B2(new_n564), .ZN(new_n580));
  AND3_X1   g394(.A1(new_n442), .A2(KEYINPUT71), .A3(G128), .ZN(new_n581));
  AOI21_X1  g395(.A(KEYINPUT71), .B1(new_n442), .B2(G128), .ZN(new_n582));
  OAI21_X1  g396(.A(new_n568), .B1(new_n581), .B2(new_n582), .ZN(new_n583));
  NAND2_X1  g397(.A1(new_n583), .A2(new_n574), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n580), .A2(new_n584), .ZN(new_n585));
  NAND3_X1  g399(.A1(new_n350), .A2(new_n585), .A3(new_n325), .ZN(new_n586));
  XNOR2_X1  g400(.A(KEYINPUT22), .B(G137), .ZN(new_n587));
  NAND3_X1  g401(.A1(new_n297), .A2(G221), .A3(G234), .ZN(new_n588));
  XNOR2_X1  g402(.A(new_n587), .B(new_n588), .ZN(new_n589));
  AND3_X1   g403(.A1(new_n577), .A2(new_n586), .A3(new_n589), .ZN(new_n590));
  AOI21_X1  g404(.A(new_n589), .B1(new_n577), .B2(new_n586), .ZN(new_n591));
  NOR2_X1   g405(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  AOI21_X1  g406(.A(new_n561), .B1(new_n592), .B2(new_n287), .ZN(new_n593));
  INV_X1    g407(.A(new_n561), .ZN(new_n594));
  NOR4_X1   g408(.A1(new_n590), .A2(new_n591), .A3(G902), .A4(new_n594), .ZN(new_n595));
  OAI21_X1  g409(.A(new_n559), .B1(new_n593), .B2(new_n595), .ZN(new_n596));
  NAND2_X1  g410(.A1(new_n596), .A2(KEYINPUT75), .ZN(new_n597));
  INV_X1    g411(.A(KEYINPUT75), .ZN(new_n598));
  OAI211_X1 g412(.A(new_n598), .B(new_n559), .C1(new_n593), .C2(new_n595), .ZN(new_n599));
  AND2_X1   g413(.A1(new_n597), .A2(new_n599), .ZN(new_n600));
  NOR2_X1   g414(.A1(new_n559), .A2(G902), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n592), .A2(new_n601), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n600), .A2(new_n602), .ZN(new_n603));
  NOR2_X1   g417(.A1(new_n557), .A2(new_n603), .ZN(new_n604));
  NAND2_X1  g418(.A1(new_n498), .A2(new_n604), .ZN(new_n605));
  XNOR2_X1  g419(.A(new_n605), .B(G101), .ZN(G3));
  OAI21_X1  g420(.A(new_n287), .B1(new_n522), .B2(new_n537), .ZN(new_n607));
  AOI21_X1  g421(.A(KEYINPUT94), .B1(new_n607), .B2(G472), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n607), .A2(G472), .ZN(new_n609));
  NAND2_X1  g423(.A1(new_n609), .A2(new_n538), .ZN(new_n610));
  AOI21_X1  g424(.A(new_n608), .B1(new_n610), .B2(KEYINPUT94), .ZN(new_n611));
  INV_X1    g425(.A(new_n603), .ZN(new_n612));
  AND2_X1   g426(.A1(new_n611), .A2(new_n612), .ZN(new_n613));
  NAND2_X1  g427(.A1(new_n613), .A2(new_n295), .ZN(new_n614));
  INV_X1    g428(.A(new_n614), .ZN(new_n615));
  AND3_X1   g429(.A1(new_n408), .A2(KEYINPUT33), .A3(new_n413), .ZN(new_n616));
  INV_X1    g430(.A(KEYINPUT33), .ZN(new_n617));
  AOI21_X1  g431(.A(new_n616), .B1(new_n414), .B2(new_n617), .ZN(new_n618));
  NOR2_X1   g432(.A1(new_n416), .A2(G902), .ZN(new_n619));
  NAND2_X1  g433(.A1(new_n414), .A2(new_n287), .ZN(new_n620));
  AOI22_X1  g434(.A1(new_n618), .A2(new_n619), .B1(new_n620), .B2(new_n416), .ZN(new_n621));
  AOI21_X1  g435(.A(new_n621), .B1(new_n363), .B2(new_n375), .ZN(new_n622));
  INV_X1    g436(.A(new_n622), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n497), .A2(new_n429), .ZN(new_n624));
  NOR2_X1   g438(.A1(new_n623), .A2(new_n624), .ZN(new_n625));
  NAND2_X1  g439(.A1(new_n615), .A2(new_n625), .ZN(new_n626));
  XOR2_X1   g440(.A(KEYINPUT34), .B(G104), .Z(new_n627));
  XNOR2_X1  g441(.A(new_n626), .B(new_n627), .ZN(G6));
  AND2_X1   g442(.A1(new_n363), .A2(new_n375), .ZN(new_n629));
  NAND2_X1  g443(.A1(new_n629), .A2(new_n420), .ZN(new_n630));
  NOR2_X1   g444(.A1(new_n630), .A2(new_n624), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n615), .A2(new_n631), .ZN(new_n632));
  XOR2_X1   g446(.A(KEYINPUT35), .B(G107), .Z(new_n633));
  XNOR2_X1  g447(.A(new_n632), .B(new_n633), .ZN(G9));
  NAND2_X1  g448(.A1(new_n577), .A2(new_n586), .ZN(new_n635));
  INV_X1    g449(.A(new_n589), .ZN(new_n636));
  NOR2_X1   g450(.A1(new_n636), .A2(KEYINPUT36), .ZN(new_n637));
  XNOR2_X1  g451(.A(new_n635), .B(new_n637), .ZN(new_n638));
  NAND2_X1  g452(.A1(new_n638), .A2(new_n601), .ZN(new_n639));
  NAND3_X1  g453(.A1(new_n597), .A2(new_n599), .A3(new_n639), .ZN(new_n640));
  INV_X1    g454(.A(KEYINPUT95), .ZN(new_n641));
  NAND2_X1  g455(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  NAND4_X1  g456(.A1(new_n597), .A2(KEYINPUT95), .A3(new_n599), .A4(new_n639), .ZN(new_n643));
  NAND2_X1  g457(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  INV_X1    g458(.A(new_n644), .ZN(new_n645));
  NAND2_X1  g459(.A1(new_n645), .A2(new_n611), .ZN(new_n646));
  INV_X1    g460(.A(KEYINPUT96), .ZN(new_n647));
  NAND2_X1  g461(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  NAND3_X1  g462(.A1(new_n645), .A2(new_n611), .A3(KEYINPUT96), .ZN(new_n649));
  NAND3_X1  g463(.A1(new_n498), .A2(new_n648), .A3(new_n649), .ZN(new_n650));
  XOR2_X1   g464(.A(KEYINPUT37), .B(G110), .Z(new_n651));
  XNOR2_X1  g465(.A(new_n650), .B(new_n651), .ZN(G12));
  NAND2_X1  g466(.A1(new_n289), .A2(new_n294), .ZN(new_n653));
  NOR3_X1   g467(.A1(new_n653), .A2(new_n644), .A3(new_n557), .ZN(new_n654));
  NOR2_X1   g468(.A1(new_n428), .A2(G900), .ZN(new_n655));
  XOR2_X1   g469(.A(new_n655), .B(KEYINPUT97), .Z(new_n656));
  NAND2_X1  g470(.A1(new_n656), .A2(new_n425), .ZN(new_n657));
  NAND3_X1  g471(.A1(new_n629), .A2(new_n420), .A3(new_n657), .ZN(new_n658));
  AND3_X1   g472(.A1(new_n477), .A2(new_n491), .A3(new_n493), .ZN(new_n659));
  AOI21_X1  g473(.A(new_n493), .B1(new_n477), .B2(new_n491), .ZN(new_n660));
  OAI21_X1  g474(.A(new_n430), .B1(new_n659), .B2(new_n660), .ZN(new_n661));
  NOR2_X1   g475(.A1(new_n658), .A2(new_n661), .ZN(new_n662));
  NAND2_X1  g476(.A1(new_n654), .A2(new_n662), .ZN(new_n663));
  XNOR2_X1  g477(.A(new_n663), .B(G128), .ZN(G30));
  XNOR2_X1  g478(.A(KEYINPUT99), .B(KEYINPUT39), .ZN(new_n665));
  XNOR2_X1  g479(.A(new_n657), .B(new_n665), .ZN(new_n666));
  NOR2_X1   g480(.A1(new_n653), .A2(new_n666), .ZN(new_n667));
  INV_X1    g481(.A(new_n667), .ZN(new_n668));
  OR2_X1    g482(.A1(new_n668), .A2(KEYINPUT40), .ZN(new_n669));
  NAND2_X1  g483(.A1(new_n668), .A2(KEYINPUT40), .ZN(new_n670));
  AOI21_X1  g484(.A(new_n419), .B1(new_n363), .B2(new_n375), .ZN(new_n671));
  NAND2_X1  g485(.A1(new_n552), .A2(new_n517), .ZN(new_n672));
  INV_X1    g486(.A(new_n517), .ZN(new_n673));
  NAND3_X1  g487(.A1(new_n673), .A2(new_n512), .A3(new_n547), .ZN(new_n674));
  NAND3_X1  g488(.A1(new_n672), .A2(new_n287), .A3(new_n674), .ZN(new_n675));
  NAND2_X1  g489(.A1(new_n675), .A2(G472), .ZN(new_n676));
  AND2_X1   g490(.A1(new_n529), .A2(new_n536), .ZN(new_n677));
  OAI211_X1 g491(.A(new_n519), .B(new_n521), .C1(new_n677), .C2(new_n517), .ZN(new_n678));
  AOI21_X1  g492(.A(new_n540), .B1(new_n678), .B2(new_n499), .ZN(new_n679));
  INV_X1    g493(.A(new_n541), .ZN(new_n680));
  OAI21_X1  g494(.A(new_n676), .B1(new_n679), .B2(new_n680), .ZN(new_n681));
  INV_X1    g495(.A(new_n681), .ZN(new_n682));
  NAND2_X1  g496(.A1(new_n495), .A2(new_n496), .ZN(new_n683));
  XNOR2_X1  g497(.A(KEYINPUT98), .B(KEYINPUT38), .ZN(new_n684));
  XNOR2_X1  g498(.A(new_n683), .B(new_n684), .ZN(new_n685));
  NOR4_X1   g499(.A1(new_n682), .A2(new_n685), .A3(new_n431), .A4(new_n640), .ZN(new_n686));
  NAND4_X1  g500(.A1(new_n669), .A2(new_n670), .A3(new_n671), .A4(new_n686), .ZN(new_n687));
  XOR2_X1   g501(.A(new_n687), .B(KEYINPUT100), .Z(new_n688));
  XNOR2_X1  g502(.A(new_n688), .B(G143), .ZN(G45));
  INV_X1    g503(.A(new_n621), .ZN(new_n690));
  NAND4_X1  g504(.A1(new_n376), .A2(new_n497), .A3(new_n690), .A4(new_n657), .ZN(new_n691));
  NAND2_X1  g505(.A1(new_n691), .A2(KEYINPUT101), .ZN(new_n692));
  NOR2_X1   g506(.A1(new_n644), .A2(new_n557), .ZN(new_n693));
  INV_X1    g507(.A(KEYINPUT101), .ZN(new_n694));
  NAND4_X1  g508(.A1(new_n622), .A2(new_n694), .A3(new_n497), .A4(new_n657), .ZN(new_n695));
  NAND4_X1  g509(.A1(new_n692), .A2(new_n295), .A3(new_n693), .A4(new_n695), .ZN(new_n696));
  INV_X1    g510(.A(KEYINPUT102), .ZN(new_n697));
  NAND2_X1  g511(.A1(new_n696), .A2(new_n697), .ZN(new_n698));
  NAND4_X1  g512(.A1(new_n654), .A2(KEYINPUT102), .A3(new_n695), .A4(new_n692), .ZN(new_n699));
  NAND2_X1  g513(.A1(new_n698), .A2(new_n699), .ZN(new_n700));
  XNOR2_X1  g514(.A(KEYINPUT103), .B(G146), .ZN(new_n701));
  XNOR2_X1  g515(.A(new_n700), .B(new_n701), .ZN(G48));
  NAND2_X1  g516(.A1(new_n286), .A2(new_n287), .ZN(new_n703));
  NAND2_X1  g517(.A1(new_n703), .A2(G469), .ZN(new_n704));
  NAND3_X1  g518(.A1(new_n704), .A2(new_n294), .A3(new_n288), .ZN(new_n705));
  NOR3_X1   g519(.A1(new_n557), .A2(new_n603), .A3(new_n705), .ZN(new_n706));
  NAND2_X1  g520(.A1(new_n625), .A2(new_n706), .ZN(new_n707));
  XNOR2_X1  g521(.A(KEYINPUT41), .B(G113), .ZN(new_n708));
  XNOR2_X1  g522(.A(new_n707), .B(new_n708), .ZN(G15));
  NAND2_X1  g523(.A1(new_n631), .A2(new_n706), .ZN(new_n710));
  XNOR2_X1  g524(.A(new_n710), .B(G116), .ZN(G18));
  INV_X1    g525(.A(KEYINPUT104), .ZN(new_n712));
  OAI21_X1  g526(.A(new_n712), .B1(new_n705), .B2(new_n661), .ZN(new_n713));
  AOI21_X1  g527(.A(new_n282), .B1(new_n286), .B2(new_n287), .ZN(new_n714));
  AOI211_X1 g528(.A(G469), .B(G902), .C1(new_n284), .C2(new_n285), .ZN(new_n715));
  NOR3_X1   g529(.A1(new_n714), .A2(new_n715), .A3(new_n293), .ZN(new_n716));
  NAND3_X1  g530(.A1(new_n716), .A2(new_n497), .A3(KEYINPUT104), .ZN(new_n717));
  NAND2_X1  g531(.A1(new_n713), .A2(new_n717), .ZN(new_n718));
  NAND4_X1  g532(.A1(new_n693), .A2(new_n421), .A3(new_n718), .A4(new_n429), .ZN(new_n719));
  XNOR2_X1  g533(.A(new_n719), .B(G119), .ZN(G21));
  OAI21_X1  g534(.A(new_n673), .B1(new_n546), .B2(new_n548), .ZN(new_n721));
  NAND3_X1  g535(.A1(new_n721), .A2(new_n519), .A3(new_n521), .ZN(new_n722));
  AOI22_X1  g536(.A1(new_n607), .A2(G472), .B1(new_n722), .B2(new_n499), .ZN(new_n723));
  AND2_X1   g537(.A1(new_n612), .A2(new_n723), .ZN(new_n724));
  AND2_X1   g538(.A1(new_n671), .A2(new_n497), .ZN(new_n725));
  NAND4_X1  g539(.A1(new_n724), .A2(new_n429), .A3(new_n716), .A4(new_n725), .ZN(new_n726));
  XNOR2_X1  g540(.A(new_n726), .B(G122), .ZN(G24));
  INV_X1    g541(.A(KEYINPUT106), .ZN(new_n728));
  INV_X1    g542(.A(new_n657), .ZN(new_n729));
  AOI211_X1 g543(.A(new_n621), .B(new_n729), .C1(new_n363), .C2(new_n375), .ZN(new_n730));
  NAND2_X1  g544(.A1(new_n722), .A2(new_n499), .ZN(new_n731));
  AND4_X1   g545(.A1(KEYINPUT105), .A2(new_n640), .A3(new_n609), .A4(new_n731), .ZN(new_n732));
  AOI21_X1  g546(.A(KEYINPUT105), .B1(new_n723), .B2(new_n640), .ZN(new_n733));
  OAI21_X1  g547(.A(new_n730), .B1(new_n732), .B2(new_n733), .ZN(new_n734));
  AND2_X1   g548(.A1(new_n713), .A2(new_n717), .ZN(new_n735));
  OAI21_X1  g549(.A(new_n728), .B1(new_n734), .B2(new_n735), .ZN(new_n736));
  NAND2_X1  g550(.A1(new_n723), .A2(new_n640), .ZN(new_n737));
  INV_X1    g551(.A(KEYINPUT105), .ZN(new_n738));
  NAND2_X1  g552(.A1(new_n737), .A2(new_n738), .ZN(new_n739));
  NAND3_X1  g553(.A1(new_n723), .A2(KEYINPUT105), .A3(new_n640), .ZN(new_n740));
  NAND2_X1  g554(.A1(new_n739), .A2(new_n740), .ZN(new_n741));
  NAND4_X1  g555(.A1(new_n741), .A2(new_n718), .A3(KEYINPUT106), .A4(new_n730), .ZN(new_n742));
  NAND2_X1  g556(.A1(new_n736), .A2(new_n742), .ZN(new_n743));
  XNOR2_X1  g557(.A(new_n743), .B(G125), .ZN(G27));
  INV_X1    g558(.A(KEYINPUT108), .ZN(new_n745));
  XNOR2_X1  g559(.A(new_n269), .B(KEYINPUT107), .ZN(new_n746));
  NAND3_X1  g560(.A1(new_n746), .A2(G469), .A3(new_n277), .ZN(new_n747));
  NOR2_X1   g561(.A1(new_n282), .A2(new_n287), .ZN(new_n748));
  NOR2_X1   g562(.A1(new_n715), .A2(new_n748), .ZN(new_n749));
  AOI21_X1  g563(.A(new_n293), .B1(new_n747), .B2(new_n749), .ZN(new_n750));
  NOR2_X1   g564(.A1(new_n683), .A2(new_n431), .ZN(new_n751));
  NAND3_X1  g565(.A1(new_n604), .A2(new_n750), .A3(new_n751), .ZN(new_n752));
  INV_X1    g566(.A(new_n730), .ZN(new_n753));
  OAI21_X1  g567(.A(new_n745), .B1(new_n752), .B2(new_n753), .ZN(new_n754));
  INV_X1    g568(.A(KEYINPUT42), .ZN(new_n755));
  OR2_X1    g569(.A1(new_n754), .A2(new_n755), .ZN(new_n756));
  NAND2_X1  g570(.A1(new_n754), .A2(new_n755), .ZN(new_n757));
  NAND2_X1  g571(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  XNOR2_X1  g572(.A(new_n758), .B(new_n199), .ZN(G33));
  INV_X1    g573(.A(KEYINPUT109), .ZN(new_n760));
  AOI21_X1  g574(.A(new_n752), .B1(new_n760), .B2(new_n658), .ZN(new_n761));
  OAI21_X1  g575(.A(new_n761), .B1(new_n760), .B2(new_n658), .ZN(new_n762));
  XNOR2_X1  g576(.A(new_n762), .B(G134), .ZN(G36));
  AOI21_X1  g577(.A(KEYINPUT45), .B1(new_n269), .B2(new_n277), .ZN(new_n764));
  AND2_X1   g578(.A1(new_n746), .A2(new_n277), .ZN(new_n765));
  AOI211_X1 g579(.A(new_n282), .B(new_n764), .C1(new_n765), .C2(KEYINPUT45), .ZN(new_n766));
  NOR2_X1   g580(.A1(new_n766), .A2(new_n748), .ZN(new_n767));
  NOR2_X1   g581(.A1(new_n767), .A2(KEYINPUT46), .ZN(new_n768));
  OR2_X1    g582(.A1(new_n768), .A2(KEYINPUT110), .ZN(new_n769));
  NAND2_X1  g583(.A1(new_n768), .A2(KEYINPUT110), .ZN(new_n770));
  AOI21_X1  g584(.A(new_n715), .B1(new_n767), .B2(KEYINPUT46), .ZN(new_n771));
  NAND3_X1  g585(.A1(new_n769), .A2(new_n770), .A3(new_n771), .ZN(new_n772));
  NAND2_X1  g586(.A1(new_n772), .A2(new_n294), .ZN(new_n773));
  NOR2_X1   g587(.A1(new_n773), .A2(new_n666), .ZN(new_n774));
  NAND2_X1  g588(.A1(new_n629), .A2(new_n690), .ZN(new_n775));
  XNOR2_X1  g589(.A(new_n775), .B(KEYINPUT43), .ZN(new_n776));
  AOI211_X1 g590(.A(new_n611), .B(new_n776), .C1(new_n600), .C2(new_n639), .ZN(new_n777));
  OR2_X1    g591(.A1(new_n777), .A2(KEYINPUT44), .ZN(new_n778));
  INV_X1    g592(.A(new_n751), .ZN(new_n779));
  AOI21_X1  g593(.A(new_n779), .B1(new_n777), .B2(KEYINPUT44), .ZN(new_n780));
  AND3_X1   g594(.A1(new_n774), .A2(new_n778), .A3(new_n780), .ZN(new_n781));
  XNOR2_X1  g595(.A(new_n781), .B(new_n194), .ZN(G39));
  AND4_X1   g596(.A1(new_n557), .A2(new_n730), .A3(new_n603), .A4(new_n751), .ZN(new_n783));
  INV_X1    g597(.A(new_n783), .ZN(new_n784));
  INV_X1    g598(.A(KEYINPUT47), .ZN(new_n785));
  NAND2_X1  g599(.A1(new_n773), .A2(new_n785), .ZN(new_n786));
  NAND3_X1  g600(.A1(new_n772), .A2(KEYINPUT47), .A3(new_n294), .ZN(new_n787));
  AOI21_X1  g601(.A(new_n784), .B1(new_n786), .B2(new_n787), .ZN(new_n788));
  XNOR2_X1  g602(.A(new_n788), .B(new_n316), .ZN(G42));
  INV_X1    g603(.A(KEYINPUT51), .ZN(new_n790));
  NOR2_X1   g604(.A1(new_n779), .A2(new_n705), .ZN(new_n791));
  NOR2_X1   g605(.A1(new_n603), .A2(new_n425), .ZN(new_n792));
  NAND3_X1  g606(.A1(new_n791), .A2(new_n682), .A3(new_n792), .ZN(new_n793));
  NOR3_X1   g607(.A1(new_n793), .A2(new_n376), .A3(new_n690), .ZN(new_n794));
  NOR2_X1   g608(.A1(new_n776), .A2(new_n425), .ZN(new_n795));
  AND2_X1   g609(.A1(new_n795), .A2(new_n791), .ZN(new_n796));
  AOI21_X1  g610(.A(new_n794), .B1(new_n796), .B2(new_n741), .ZN(new_n797));
  NAND2_X1  g611(.A1(new_n795), .A2(new_n724), .ZN(new_n798));
  NAND3_X1  g612(.A1(new_n685), .A2(new_n431), .A3(new_n716), .ZN(new_n799));
  NOR2_X1   g613(.A1(new_n798), .A2(new_n799), .ZN(new_n800));
  AND2_X1   g614(.A1(new_n800), .A2(KEYINPUT50), .ZN(new_n801));
  NOR2_X1   g615(.A1(new_n800), .A2(KEYINPUT50), .ZN(new_n802));
  OAI21_X1  g616(.A(new_n797), .B1(new_n801), .B2(new_n802), .ZN(new_n803));
  XOR2_X1   g617(.A(new_n803), .B(KEYINPUT114), .Z(new_n804));
  INV_X1    g618(.A(new_n798), .ZN(new_n805));
  NAND2_X1  g619(.A1(new_n805), .A2(new_n751), .ZN(new_n806));
  AND2_X1   g620(.A1(new_n786), .A2(new_n787), .ZN(new_n807));
  NOR2_X1   g621(.A1(new_n714), .A2(new_n715), .ZN(new_n808));
  NAND2_X1  g622(.A1(new_n808), .A2(new_n293), .ZN(new_n809));
  AOI21_X1  g623(.A(new_n806), .B1(new_n807), .B2(new_n809), .ZN(new_n810));
  OAI21_X1  g624(.A(new_n790), .B1(new_n804), .B2(new_n810), .ZN(new_n811));
  OR3_X1    g625(.A1(new_n810), .A2(new_n790), .A3(new_n803), .ZN(new_n812));
  NAND2_X1  g626(.A1(new_n805), .A2(new_n718), .ZN(new_n813));
  XNOR2_X1  g627(.A(new_n813), .B(KEYINPUT115), .ZN(new_n814));
  NAND2_X1  g628(.A1(new_n796), .A2(new_n604), .ZN(new_n815));
  XNOR2_X1  g629(.A(new_n815), .B(KEYINPUT48), .ZN(new_n816));
  OR2_X1    g630(.A1(new_n793), .A2(new_n623), .ZN(new_n817));
  AND4_X1   g631(.A1(new_n422), .A2(new_n814), .A3(new_n816), .A4(new_n817), .ZN(new_n818));
  NAND3_X1  g632(.A1(new_n811), .A2(new_n812), .A3(new_n818), .ZN(new_n819));
  AND3_X1   g633(.A1(new_n756), .A2(new_n762), .A3(new_n757), .ZN(new_n820));
  OAI211_X1 g634(.A(new_n613), .B(new_n295), .C1(new_n631), .C2(new_n625), .ZN(new_n821));
  NAND3_X1  g635(.A1(new_n650), .A2(new_n719), .A3(new_n821), .ZN(new_n822));
  NAND4_X1  g636(.A1(new_n605), .A2(new_n707), .A3(new_n710), .A4(new_n726), .ZN(new_n823));
  NOR2_X1   g637(.A1(new_n822), .A2(new_n823), .ZN(new_n824));
  NAND2_X1  g638(.A1(new_n654), .A2(new_n421), .ZN(new_n825));
  NAND3_X1  g639(.A1(new_n741), .A2(new_n622), .A3(new_n750), .ZN(new_n826));
  NAND2_X1  g640(.A1(new_n825), .A2(new_n826), .ZN(new_n827));
  NAND3_X1  g641(.A1(new_n827), .A2(new_n657), .A3(new_n751), .ZN(new_n828));
  AND3_X1   g642(.A1(new_n820), .A2(new_n824), .A3(new_n828), .ZN(new_n829));
  INV_X1    g643(.A(KEYINPUT52), .ZN(new_n830));
  INV_X1    g644(.A(new_n700), .ZN(new_n831));
  NAND4_X1  g645(.A1(new_n597), .A2(new_n599), .A3(new_n639), .A4(new_n657), .ZN(new_n832));
  INV_X1    g646(.A(new_n832), .ZN(new_n833));
  NAND4_X1  g647(.A1(new_n681), .A2(new_n671), .A3(new_n497), .A4(new_n833), .ZN(new_n834));
  INV_X1    g648(.A(new_n750), .ZN(new_n835));
  OAI21_X1  g649(.A(KEYINPUT112), .B1(new_n834), .B2(new_n835), .ZN(new_n836));
  INV_X1    g650(.A(KEYINPUT112), .ZN(new_n837));
  NAND2_X1  g651(.A1(new_n539), .A2(new_n541), .ZN(new_n838));
  AOI21_X1  g652(.A(new_n832), .B1(new_n838), .B2(new_n676), .ZN(new_n839));
  NAND4_X1  g653(.A1(new_n725), .A2(new_n837), .A3(new_n750), .A4(new_n839), .ZN(new_n840));
  AOI22_X1  g654(.A1(new_n836), .A2(new_n840), .B1(new_n654), .B2(new_n662), .ZN(new_n841));
  NAND2_X1  g655(.A1(new_n841), .A2(new_n743), .ZN(new_n842));
  OAI21_X1  g656(.A(new_n830), .B1(new_n831), .B2(new_n842), .ZN(new_n843));
  AND2_X1   g657(.A1(new_n841), .A2(new_n743), .ZN(new_n844));
  NAND3_X1  g658(.A1(new_n844), .A2(KEYINPUT52), .A3(new_n700), .ZN(new_n845));
  NAND2_X1  g659(.A1(new_n843), .A2(new_n845), .ZN(new_n846));
  NAND2_X1  g660(.A1(new_n829), .A2(new_n846), .ZN(new_n847));
  NAND3_X1  g661(.A1(new_n820), .A2(new_n824), .A3(new_n828), .ZN(new_n848));
  AOI21_X1  g662(.A(KEYINPUT52), .B1(new_n844), .B2(new_n700), .ZN(new_n849));
  AND4_X1   g663(.A1(KEYINPUT52), .A2(new_n700), .A3(new_n743), .A4(new_n841), .ZN(new_n850));
  OAI21_X1  g664(.A(KEYINPUT113), .B1(new_n849), .B2(new_n850), .ZN(new_n851));
  INV_X1    g665(.A(KEYINPUT113), .ZN(new_n852));
  NAND3_X1  g666(.A1(new_n843), .A2(new_n845), .A3(new_n852), .ZN(new_n853));
  AOI21_X1  g667(.A(new_n848), .B1(new_n851), .B2(new_n853), .ZN(new_n854));
  MUX2_X1   g668(.A(new_n847), .B(new_n854), .S(KEYINPUT53), .Z(new_n855));
  NAND2_X1  g669(.A1(new_n855), .A2(KEYINPUT54), .ZN(new_n856));
  INV_X1    g670(.A(KEYINPUT54), .ZN(new_n857));
  NAND3_X1  g671(.A1(new_n829), .A2(KEYINPUT53), .A3(new_n846), .ZN(new_n858));
  OAI211_X1 g672(.A(new_n857), .B(new_n858), .C1(new_n854), .C2(KEYINPUT53), .ZN(new_n859));
  NAND2_X1  g673(.A1(new_n856), .A2(new_n859), .ZN(new_n860));
  OAI22_X1  g674(.A1(new_n819), .A2(new_n860), .B1(G952), .B2(G953), .ZN(new_n861));
  NOR4_X1   g675(.A1(new_n775), .A2(new_n603), .A3(new_n293), .A4(new_n431), .ZN(new_n862));
  NOR2_X1   g676(.A1(new_n862), .A2(KEYINPUT111), .ZN(new_n863));
  NAND2_X1  g677(.A1(new_n862), .A2(KEYINPUT111), .ZN(new_n864));
  XNOR2_X1  g678(.A(new_n808), .B(KEYINPUT49), .ZN(new_n865));
  NAND4_X1  g679(.A1(new_n864), .A2(new_n685), .A3(new_n682), .A4(new_n865), .ZN(new_n866));
  OAI21_X1  g680(.A(new_n861), .B1(new_n863), .B2(new_n866), .ZN(G75));
  OAI21_X1  g681(.A(new_n858), .B1(new_n854), .B2(KEYINPUT53), .ZN(new_n868));
  INV_X1    g682(.A(new_n868), .ZN(new_n869));
  NOR2_X1   g683(.A1(new_n869), .A2(new_n287), .ZN(new_n870));
  AOI21_X1  g684(.A(KEYINPUT56), .B1(new_n870), .B2(G210), .ZN(new_n871));
  NAND2_X1  g685(.A1(new_n487), .A2(new_n490), .ZN(new_n872));
  XNOR2_X1  g686(.A(new_n872), .B(new_n489), .ZN(new_n873));
  XOR2_X1   g687(.A(new_n873), .B(KEYINPUT55), .Z(new_n874));
  INV_X1    g688(.A(new_n874), .ZN(new_n875));
  NAND2_X1  g689(.A1(new_n871), .A2(new_n875), .ZN(new_n876));
  NOR2_X1   g690(.A1(new_n297), .A2(G952), .ZN(new_n877));
  INV_X1    g691(.A(new_n877), .ZN(new_n878));
  NAND2_X1  g692(.A1(new_n876), .A2(new_n878), .ZN(new_n879));
  INV_X1    g693(.A(KEYINPUT116), .ZN(new_n880));
  OAI21_X1  g694(.A(new_n880), .B1(new_n871), .B2(new_n875), .ZN(new_n881));
  INV_X1    g695(.A(new_n871), .ZN(new_n882));
  NAND3_X1  g696(.A1(new_n882), .A2(KEYINPUT116), .A3(new_n874), .ZN(new_n883));
  AOI21_X1  g697(.A(new_n879), .B1(new_n881), .B2(new_n883), .ZN(G51));
  NAND2_X1  g698(.A1(new_n868), .A2(KEYINPUT54), .ZN(new_n885));
  NAND3_X1  g699(.A1(new_n885), .A2(KEYINPUT117), .A3(new_n859), .ZN(new_n886));
  INV_X1    g700(.A(KEYINPUT117), .ZN(new_n887));
  NAND3_X1  g701(.A1(new_n868), .A2(new_n887), .A3(KEYINPUT54), .ZN(new_n888));
  XNOR2_X1  g702(.A(new_n748), .B(KEYINPUT57), .ZN(new_n889));
  NAND3_X1  g703(.A1(new_n886), .A2(new_n888), .A3(new_n889), .ZN(new_n890));
  INV_X1    g704(.A(KEYINPUT118), .ZN(new_n891));
  NAND2_X1  g705(.A1(new_n890), .A2(new_n891), .ZN(new_n892));
  NAND4_X1  g706(.A1(new_n886), .A2(KEYINPUT118), .A3(new_n888), .A4(new_n889), .ZN(new_n893));
  NAND3_X1  g707(.A1(new_n892), .A2(new_n286), .A3(new_n893), .ZN(new_n894));
  NAND2_X1  g708(.A1(new_n870), .A2(new_n766), .ZN(new_n895));
  AOI21_X1  g709(.A(new_n877), .B1(new_n894), .B2(new_n895), .ZN(G54));
  NAND3_X1  g710(.A1(new_n870), .A2(KEYINPUT58), .A3(G475), .ZN(new_n897));
  NOR2_X1   g711(.A1(new_n347), .A2(new_n373), .ZN(new_n898));
  AND2_X1   g712(.A1(new_n897), .A2(new_n898), .ZN(new_n899));
  NOR2_X1   g713(.A1(new_n897), .A2(new_n898), .ZN(new_n900));
  NOR3_X1   g714(.A1(new_n899), .A2(new_n900), .A3(new_n877), .ZN(G60));
  NAND2_X1  g715(.A1(G478), .A2(G902), .ZN(new_n902));
  XNOR2_X1  g716(.A(new_n902), .B(KEYINPUT59), .ZN(new_n903));
  AND4_X1   g717(.A1(new_n618), .A2(new_n886), .A3(new_n888), .A4(new_n903), .ZN(new_n904));
  AOI21_X1  g718(.A(new_n618), .B1(new_n860), .B2(new_n903), .ZN(new_n905));
  NOR3_X1   g719(.A1(new_n904), .A2(new_n905), .A3(new_n877), .ZN(G63));
  NAND2_X1  g720(.A1(G217), .A2(G902), .ZN(new_n907));
  XNOR2_X1  g721(.A(new_n907), .B(KEYINPUT60), .ZN(new_n908));
  NOR2_X1   g722(.A1(new_n869), .A2(new_n908), .ZN(new_n909));
  NAND2_X1  g723(.A1(new_n909), .A2(new_n638), .ZN(new_n910));
  XOR2_X1   g724(.A(new_n592), .B(KEYINPUT119), .Z(new_n911));
  INV_X1    g725(.A(new_n911), .ZN(new_n912));
  OAI211_X1 g726(.A(new_n910), .B(new_n878), .C1(new_n909), .C2(new_n912), .ZN(new_n913));
  INV_X1    g727(.A(KEYINPUT61), .ZN(new_n914));
  XNOR2_X1  g728(.A(new_n913), .B(new_n914), .ZN(G66));
  AND3_X1   g729(.A1(new_n427), .A2(G224), .A3(G953), .ZN(new_n916));
  AOI21_X1  g730(.A(new_n916), .B1(new_n824), .B2(new_n297), .ZN(new_n917));
  OAI21_X1  g731(.A(new_n872), .B1(G898), .B2(new_n297), .ZN(new_n918));
  XNOR2_X1  g732(.A(new_n917), .B(new_n918), .ZN(G69));
  INV_X1    g733(.A(G900), .ZN(new_n920));
  OAI21_X1  g734(.A(G953), .B1(new_n265), .B2(new_n920), .ZN(new_n921));
  NOR2_X1   g735(.A1(new_n921), .A2(KEYINPUT124), .ZN(new_n922));
  XNOR2_X1  g736(.A(new_n922), .B(KEYINPUT125), .ZN(new_n923));
  NAND3_X1  g737(.A1(new_n774), .A2(new_n604), .A3(new_n725), .ZN(new_n924));
  AND2_X1   g738(.A1(new_n743), .A2(new_n663), .ZN(new_n925));
  AND3_X1   g739(.A1(new_n924), .A2(new_n700), .A3(new_n925), .ZN(new_n926));
  INV_X1    g740(.A(new_n820), .ZN(new_n927));
  NOR2_X1   g741(.A1(new_n781), .A2(new_n927), .ZN(new_n928));
  OAI211_X1 g742(.A(new_n926), .B(new_n928), .C1(new_n807), .C2(new_n784), .ZN(new_n929));
  NAND2_X1  g743(.A1(new_n929), .A2(new_n297), .ZN(new_n930));
  XNOR2_X1  g744(.A(new_n371), .B(KEYINPUT122), .ZN(new_n931));
  NOR2_X1   g745(.A1(new_n506), .A2(new_n507), .ZN(new_n932));
  XNOR2_X1  g746(.A(new_n931), .B(new_n932), .ZN(new_n933));
  XOR2_X1   g747(.A(KEYINPUT120), .B(KEYINPUT121), .Z(new_n934));
  XNOR2_X1  g748(.A(new_n933), .B(new_n934), .ZN(new_n935));
  AOI21_X1  g749(.A(new_n935), .B1(new_n920), .B2(G953), .ZN(new_n936));
  AOI22_X1  g750(.A1(new_n930), .A2(new_n936), .B1(KEYINPUT124), .B2(new_n921), .ZN(new_n937));
  NAND2_X1  g751(.A1(new_n630), .A2(new_n623), .ZN(new_n938));
  NAND4_X1  g752(.A1(new_n667), .A2(new_n938), .A3(new_n604), .A4(new_n751), .ZN(new_n939));
  XNOR2_X1  g753(.A(new_n939), .B(KEYINPUT123), .ZN(new_n940));
  NOR3_X1   g754(.A1(new_n781), .A2(new_n788), .A3(new_n940), .ZN(new_n941));
  NAND3_X1  g755(.A1(new_n688), .A2(new_n700), .A3(new_n925), .ZN(new_n942));
  OR2_X1    g756(.A1(new_n942), .A2(KEYINPUT62), .ZN(new_n943));
  NAND2_X1  g757(.A1(new_n942), .A2(KEYINPUT62), .ZN(new_n944));
  NAND3_X1  g758(.A1(new_n941), .A2(new_n943), .A3(new_n944), .ZN(new_n945));
  NAND3_X1  g759(.A1(new_n945), .A2(new_n297), .A3(new_n935), .ZN(new_n946));
  AOI21_X1  g760(.A(new_n923), .B1(new_n937), .B2(new_n946), .ZN(new_n947));
  NAND3_X1  g761(.A1(new_n924), .A2(new_n700), .A3(new_n925), .ZN(new_n948));
  NOR4_X1   g762(.A1(new_n948), .A2(new_n781), .A3(new_n788), .A4(new_n927), .ZN(new_n949));
  OAI21_X1  g763(.A(new_n936), .B1(new_n949), .B2(G953), .ZN(new_n950));
  NAND2_X1  g764(.A1(new_n921), .A2(KEYINPUT124), .ZN(new_n951));
  AND4_X1   g765(.A1(new_n946), .A2(new_n950), .A3(new_n951), .A4(new_n923), .ZN(new_n952));
  NOR2_X1   g766(.A1(new_n947), .A2(new_n952), .ZN(G72));
  NAND2_X1  g767(.A1(G472), .A2(G902), .ZN(new_n954));
  XOR2_X1   g768(.A(new_n954), .B(KEYINPUT63), .Z(new_n955));
  INV_X1    g769(.A(new_n824), .ZN(new_n956));
  OAI21_X1  g770(.A(new_n955), .B1(new_n929), .B2(new_n956), .ZN(new_n957));
  XNOR2_X1  g771(.A(new_n553), .B(KEYINPUT126), .ZN(new_n958));
  AOI21_X1  g772(.A(new_n877), .B1(new_n957), .B2(new_n958), .ZN(new_n959));
  INV_X1    g773(.A(new_n553), .ZN(new_n960));
  NAND4_X1  g774(.A1(new_n855), .A2(new_n960), .A3(new_n672), .A4(new_n955), .ZN(new_n961));
  OAI21_X1  g775(.A(new_n955), .B1(new_n945), .B2(new_n956), .ZN(new_n962));
  NAND3_X1  g776(.A1(new_n962), .A2(new_n517), .A3(new_n552), .ZN(new_n963));
  AND3_X1   g777(.A1(new_n959), .A2(new_n961), .A3(new_n963), .ZN(G57));
endmodule


