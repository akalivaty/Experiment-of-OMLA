//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 1 0 1 1 0 0 0 0 1 0 1 0 0 1 1 1 1 1 0 0 1 1 1 0 1 1 0 1 0 0 1 1 1 0 1 1 0 1 0 1 1 1 0 1 1 1 0 0 0 1 0 1 1 1 1 1 1 0 0 0 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:36:15 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n241, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1237, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1246, new_n1247,
    new_n1248, new_n1249, new_n1250, new_n1251, new_n1252, new_n1253,
    new_n1254, new_n1255, new_n1257, new_n1258, new_n1259, new_n1260,
    new_n1261, new_n1262, new_n1263, new_n1264, new_n1265, new_n1266,
    new_n1267, new_n1268, new_n1269, new_n1271, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1316, new_n1317,
    new_n1318, new_n1319, new_n1320, new_n1321, new_n1322, new_n1323,
    new_n1324, new_n1325, new_n1326, new_n1327, new_n1328, new_n1329,
    new_n1330, new_n1331;
  INV_X1    g0000(.A(KEYINPUT64), .ZN(new_n201));
  INV_X1    g0001(.A(G58), .ZN(new_n202));
  INV_X1    g0002(.A(G68), .ZN(new_n203));
  NAND3_X1  g0003(.A1(new_n201), .A2(new_n202), .A3(new_n203), .ZN(new_n204));
  OAI21_X1  g0004(.A(KEYINPUT64), .B1(G58), .B2(G68), .ZN(new_n205));
  NAND2_X1  g0005(.A1(new_n204), .A2(new_n205), .ZN(new_n206));
  INV_X1    g0006(.A(new_n206), .ZN(new_n207));
  NOR3_X1   g0007(.A1(new_n207), .A2(G50), .A3(G77), .ZN(G353));
  OAI21_X1  g0008(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0009(.A1(new_n207), .A2(G50), .ZN(new_n210));
  NAND2_X1  g0010(.A1(G1), .A2(G13), .ZN(new_n211));
  INV_X1    g0011(.A(G20), .ZN(new_n212));
  NOR2_X1   g0012(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  INV_X1    g0013(.A(new_n213), .ZN(new_n214));
  INV_X1    g0014(.A(G1), .ZN(new_n215));
  NOR3_X1   g0015(.A1(new_n215), .A2(new_n212), .A3(G13), .ZN(new_n216));
  OAI211_X1 g0016(.A(new_n216), .B(G250), .C1(G257), .C2(G264), .ZN(new_n217));
  INV_X1    g0017(.A(KEYINPUT0), .ZN(new_n218));
  OAI22_X1  g0018(.A1(new_n210), .A2(new_n214), .B1(new_n217), .B2(new_n218), .ZN(new_n219));
  AOI22_X1  g0019(.A1(G87), .A2(G250), .B1(G107), .B2(G264), .ZN(new_n220));
  NAND2_X1  g0020(.A1(G97), .A2(G257), .ZN(new_n221));
  NAND2_X1  g0021(.A1(G68), .A2(G238), .ZN(new_n222));
  NAND3_X1  g0022(.A1(new_n220), .A2(new_n221), .A3(new_n222), .ZN(new_n223));
  AOI22_X1  g0023(.A1(G50), .A2(G226), .B1(G77), .B2(G244), .ZN(new_n224));
  INV_X1    g0024(.A(G116), .ZN(new_n225));
  INV_X1    g0025(.A(G270), .ZN(new_n226));
  OAI21_X1  g0026(.A(new_n224), .B1(new_n225), .B2(new_n226), .ZN(new_n227));
  AOI211_X1 g0027(.A(new_n223), .B(new_n227), .C1(G58), .C2(G232), .ZN(new_n228));
  AOI21_X1  g0028(.A(new_n228), .B1(G1), .B2(G20), .ZN(new_n229));
  XOR2_X1   g0029(.A(new_n229), .B(KEYINPUT1), .Z(new_n230));
  AOI211_X1 g0030(.A(new_n219), .B(new_n230), .C1(new_n218), .C2(new_n217), .ZN(G361));
  XNOR2_X1  g0031(.A(G238), .B(G244), .ZN(new_n232));
  INV_X1    g0032(.A(G232), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n232), .B(new_n233), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n234), .B(KEYINPUT2), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n235), .B(G226), .ZN(new_n236));
  XNOR2_X1  g0036(.A(G250), .B(G257), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n237), .B(G264), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n238), .B(new_n226), .ZN(new_n239));
  XOR2_X1   g0039(.A(new_n236), .B(new_n239), .Z(G358));
  XNOR2_X1  g0040(.A(G68), .B(G77), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n241), .B(KEYINPUT65), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n242), .B(G50), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n243), .B(new_n202), .ZN(new_n244));
  XNOR2_X1  g0044(.A(G87), .B(G97), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n245), .B(KEYINPUT66), .ZN(new_n246));
  INV_X1    g0046(.A(G107), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n246), .B(new_n247), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n248), .B(new_n225), .ZN(new_n249));
  XNOR2_X1  g0049(.A(new_n244), .B(new_n249), .ZN(G351));
  NAND3_X1  g0050(.A1(new_n215), .A2(G13), .A3(G20), .ZN(new_n251));
  NOR2_X1   g0051(.A1(new_n251), .A2(G77), .ZN(new_n252));
  XOR2_X1   g0052(.A(KEYINPUT15), .B(G87), .Z(new_n253));
  NAND3_X1  g0053(.A1(new_n253), .A2(new_n212), .A3(G33), .ZN(new_n254));
  INV_X1    g0054(.A(G77), .ZN(new_n255));
  OAI21_X1  g0055(.A(KEYINPUT69), .B1(new_n212), .B2(new_n255), .ZN(new_n256));
  OAI21_X1  g0056(.A(KEYINPUT67), .B1(G20), .B2(G33), .ZN(new_n257));
  INV_X1    g0057(.A(new_n257), .ZN(new_n258));
  NOR3_X1   g0058(.A1(KEYINPUT67), .A2(G20), .A3(G33), .ZN(new_n259));
  OR2_X1    g0059(.A1(new_n258), .A2(new_n259), .ZN(new_n260));
  XNOR2_X1  g0060(.A(KEYINPUT8), .B(G58), .ZN(new_n261));
  INV_X1    g0061(.A(new_n261), .ZN(new_n262));
  AOI22_X1  g0062(.A1(new_n254), .A2(new_n256), .B1(new_n260), .B2(new_n262), .ZN(new_n263));
  INV_X1    g0063(.A(KEYINPUT69), .ZN(new_n264));
  OAI21_X1  g0064(.A(new_n263), .B1(new_n264), .B2(new_n254), .ZN(new_n265));
  NAND3_X1  g0065(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n266));
  NAND2_X1  g0066(.A1(new_n266), .A2(new_n211), .ZN(new_n267));
  AOI21_X1  g0067(.A(new_n252), .B1(new_n265), .B2(new_n267), .ZN(new_n268));
  AOI21_X1  g0068(.A(new_n267), .B1(new_n215), .B2(G20), .ZN(new_n269));
  INV_X1    g0069(.A(new_n269), .ZN(new_n270));
  OAI21_X1  g0070(.A(new_n268), .B1(new_n255), .B2(new_n270), .ZN(new_n271));
  XNOR2_X1  g0071(.A(KEYINPUT3), .B(G33), .ZN(new_n272));
  NAND2_X1  g0072(.A1(G238), .A2(G1698), .ZN(new_n273));
  OAI21_X1  g0073(.A(new_n273), .B1(new_n233), .B2(G1698), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n272), .A2(new_n274), .ZN(new_n275));
  OAI21_X1  g0075(.A(new_n275), .B1(new_n247), .B2(new_n272), .ZN(new_n276));
  XNOR2_X1  g0076(.A(new_n276), .B(KEYINPUT68), .ZN(new_n277));
  NAND2_X1  g0077(.A1(G33), .A2(G41), .ZN(new_n278));
  NAND3_X1  g0078(.A1(new_n278), .A2(G1), .A3(G13), .ZN(new_n279));
  INV_X1    g0079(.A(new_n279), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n277), .A2(new_n280), .ZN(new_n281));
  OAI21_X1  g0081(.A(new_n215), .B1(G41), .B2(G45), .ZN(new_n282));
  INV_X1    g0082(.A(G274), .ZN(new_n283));
  NOR2_X1   g0083(.A1(new_n282), .A2(new_n283), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n279), .A2(new_n282), .ZN(new_n285));
  INV_X1    g0085(.A(new_n285), .ZN(new_n286));
  AOI21_X1  g0086(.A(new_n284), .B1(new_n286), .B2(G244), .ZN(new_n287));
  AND2_X1   g0087(.A1(new_n281), .A2(new_n287), .ZN(new_n288));
  OAI211_X1 g0088(.A(new_n271), .B(KEYINPUT70), .C1(new_n288), .C2(G169), .ZN(new_n289));
  INV_X1    g0089(.A(G179), .ZN(new_n290));
  NAND2_X1  g0090(.A1(new_n288), .A2(new_n290), .ZN(new_n291));
  INV_X1    g0091(.A(KEYINPUT70), .ZN(new_n292));
  AOI21_X1  g0092(.A(G169), .B1(new_n281), .B2(new_n287), .ZN(new_n293));
  NOR2_X1   g0093(.A1(new_n270), .A2(new_n255), .ZN(new_n294));
  AOI211_X1 g0094(.A(new_n252), .B(new_n294), .C1(new_n265), .C2(new_n267), .ZN(new_n295));
  OAI21_X1  g0095(.A(new_n292), .B1(new_n293), .B2(new_n295), .ZN(new_n296));
  NAND3_X1  g0096(.A1(new_n289), .A2(new_n291), .A3(new_n296), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n288), .A2(G190), .ZN(new_n298));
  INV_X1    g0098(.A(G200), .ZN(new_n299));
  OAI211_X1 g0099(.A(new_n298), .B(new_n295), .C1(new_n299), .C2(new_n288), .ZN(new_n300));
  AND2_X1   g0100(.A1(new_n297), .A2(new_n300), .ZN(new_n301));
  INV_X1    g0101(.A(new_n284), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n286), .A2(G226), .ZN(new_n303));
  INV_X1    g0103(.A(G33), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n304), .A2(KEYINPUT3), .ZN(new_n305));
  INV_X1    g0105(.A(KEYINPUT3), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n306), .A2(G33), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n305), .A2(new_n307), .ZN(new_n308));
  NOR2_X1   g0108(.A1(new_n308), .A2(G1698), .ZN(new_n309));
  AOI22_X1  g0109(.A1(new_n309), .A2(G222), .B1(G77), .B2(new_n308), .ZN(new_n310));
  NAND3_X1  g0110(.A1(new_n272), .A2(G223), .A3(G1698), .ZN(new_n311));
  AND2_X1   g0111(.A1(new_n310), .A2(new_n311), .ZN(new_n312));
  OAI211_X1 g0112(.A(new_n302), .B(new_n303), .C1(new_n312), .C2(new_n279), .ZN(new_n313));
  INV_X1    g0113(.A(G190), .ZN(new_n314));
  NOR2_X1   g0114(.A1(new_n313), .A2(new_n314), .ZN(new_n315));
  AOI21_X1  g0115(.A(new_n315), .B1(G200), .B2(new_n313), .ZN(new_n316));
  OAI21_X1  g0116(.A(G20), .B1(new_n207), .B2(G50), .ZN(new_n317));
  NAND3_X1  g0117(.A1(new_n262), .A2(new_n212), .A3(G33), .ZN(new_n318));
  INV_X1    g0118(.A(G150), .ZN(new_n319));
  NOR2_X1   g0119(.A1(new_n258), .A2(new_n259), .ZN(new_n320));
  OAI211_X1 g0120(.A(new_n317), .B(new_n318), .C1(new_n319), .C2(new_n320), .ZN(new_n321));
  INV_X1    g0121(.A(G50), .ZN(new_n322));
  INV_X1    g0122(.A(new_n251), .ZN(new_n323));
  AOI22_X1  g0123(.A1(new_n321), .A2(new_n267), .B1(new_n322), .B2(new_n323), .ZN(new_n324));
  OAI21_X1  g0124(.A(new_n324), .B1(new_n322), .B2(new_n270), .ZN(new_n325));
  INV_X1    g0125(.A(KEYINPUT9), .ZN(new_n326));
  OR2_X1    g0126(.A1(new_n325), .A2(new_n326), .ZN(new_n327));
  AND3_X1   g0127(.A1(new_n325), .A2(KEYINPUT71), .A3(new_n326), .ZN(new_n328));
  AOI21_X1  g0128(.A(KEYINPUT71), .B1(new_n325), .B2(new_n326), .ZN(new_n329));
  OAI211_X1 g0129(.A(new_n316), .B(new_n327), .C1(new_n328), .C2(new_n329), .ZN(new_n330));
  INV_X1    g0130(.A(KEYINPUT10), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n330), .A2(new_n331), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n325), .A2(new_n326), .ZN(new_n333));
  INV_X1    g0133(.A(KEYINPUT71), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n333), .A2(new_n334), .ZN(new_n335));
  NAND3_X1  g0135(.A1(new_n325), .A2(KEYINPUT71), .A3(new_n326), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n335), .A2(new_n336), .ZN(new_n337));
  NAND4_X1  g0137(.A1(new_n337), .A2(KEYINPUT10), .A3(new_n327), .A4(new_n316), .ZN(new_n338));
  INV_X1    g0138(.A(G169), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n313), .A2(new_n339), .ZN(new_n340));
  OAI211_X1 g0140(.A(new_n325), .B(new_n340), .C1(G179), .C2(new_n313), .ZN(new_n341));
  NAND4_X1  g0141(.A1(new_n301), .A2(new_n332), .A3(new_n338), .A4(new_n341), .ZN(new_n342));
  INV_X1    g0142(.A(KEYINPUT72), .ZN(new_n343));
  NAND2_X1  g0143(.A1(new_n342), .A2(new_n343), .ZN(new_n344));
  NOR2_X1   g0144(.A1(new_n320), .A2(new_n322), .ZN(new_n345));
  NAND3_X1  g0145(.A1(new_n212), .A2(G33), .A3(G77), .ZN(new_n346));
  OAI21_X1  g0146(.A(new_n346), .B1(new_n212), .B2(G68), .ZN(new_n347));
  OAI21_X1  g0147(.A(new_n267), .B1(new_n345), .B2(new_n347), .ZN(new_n348));
  INV_X1    g0148(.A(KEYINPUT11), .ZN(new_n349));
  XNOR2_X1  g0149(.A(new_n348), .B(new_n349), .ZN(new_n350));
  NAND4_X1  g0150(.A1(new_n215), .A2(new_n203), .A3(G13), .A4(G20), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n351), .A2(KEYINPUT74), .ZN(new_n352));
  XOR2_X1   g0152(.A(new_n352), .B(KEYINPUT12), .Z(new_n353));
  NAND2_X1  g0153(.A1(new_n269), .A2(G68), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n353), .A2(new_n354), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n355), .A2(KEYINPUT75), .ZN(new_n356));
  INV_X1    g0156(.A(KEYINPUT75), .ZN(new_n357));
  NAND3_X1  g0157(.A1(new_n353), .A2(new_n357), .A3(new_n354), .ZN(new_n358));
  AOI21_X1  g0158(.A(new_n350), .B1(new_n356), .B2(new_n358), .ZN(new_n359));
  NAND4_X1  g0159(.A1(new_n305), .A2(new_n307), .A3(G232), .A4(G1698), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n360), .A2(KEYINPUT73), .ZN(new_n361));
  INV_X1    g0161(.A(KEYINPUT73), .ZN(new_n362));
  NAND4_X1  g0162(.A1(new_n272), .A2(new_n362), .A3(G232), .A4(G1698), .ZN(new_n363));
  INV_X1    g0163(.A(G1698), .ZN(new_n364));
  NAND3_X1  g0164(.A1(new_n272), .A2(G226), .A3(new_n364), .ZN(new_n365));
  NAND2_X1  g0165(.A1(G33), .A2(G97), .ZN(new_n366));
  NAND4_X1  g0166(.A1(new_n361), .A2(new_n363), .A3(new_n365), .A4(new_n366), .ZN(new_n367));
  AOI21_X1  g0167(.A(new_n284), .B1(new_n367), .B2(new_n280), .ZN(new_n368));
  INV_X1    g0168(.A(KEYINPUT13), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n286), .A2(G238), .ZN(new_n370));
  AND3_X1   g0170(.A1(new_n368), .A2(new_n369), .A3(new_n370), .ZN(new_n371));
  AOI21_X1  g0171(.A(new_n369), .B1(new_n368), .B2(new_n370), .ZN(new_n372));
  OAI21_X1  g0172(.A(G200), .B1(new_n371), .B2(new_n372), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n368), .A2(new_n370), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n374), .A2(KEYINPUT13), .ZN(new_n375));
  NAND3_X1  g0175(.A1(new_n368), .A2(new_n369), .A3(new_n370), .ZN(new_n376));
  NAND3_X1  g0176(.A1(new_n375), .A2(G190), .A3(new_n376), .ZN(new_n377));
  AND3_X1   g0177(.A1(new_n359), .A2(new_n373), .A3(new_n377), .ZN(new_n378));
  OAI21_X1  g0178(.A(G169), .B1(new_n371), .B2(new_n372), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n379), .A2(KEYINPUT14), .ZN(new_n380));
  NAND3_X1  g0180(.A1(new_n375), .A2(G179), .A3(new_n376), .ZN(new_n381));
  INV_X1    g0181(.A(KEYINPUT14), .ZN(new_n382));
  OAI211_X1 g0182(.A(new_n382), .B(G169), .C1(new_n371), .C2(new_n372), .ZN(new_n383));
  NAND3_X1  g0183(.A1(new_n380), .A2(new_n381), .A3(new_n383), .ZN(new_n384));
  INV_X1    g0184(.A(new_n359), .ZN(new_n385));
  AOI21_X1  g0185(.A(new_n378), .B1(new_n384), .B2(new_n385), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n344), .A2(new_n386), .ZN(new_n387));
  NOR2_X1   g0187(.A1(new_n202), .A2(new_n203), .ZN(new_n388));
  OR2_X1    g0188(.A1(new_n206), .A2(new_n388), .ZN(new_n389));
  AOI22_X1  g0189(.A1(new_n389), .A2(G20), .B1(G159), .B2(new_n260), .ZN(new_n390));
  INV_X1    g0190(.A(KEYINPUT7), .ZN(new_n391));
  NOR3_X1   g0191(.A1(new_n272), .A2(new_n391), .A3(G20), .ZN(new_n392));
  INV_X1    g0192(.A(KEYINPUT76), .ZN(new_n393));
  AND3_X1   g0193(.A1(new_n305), .A2(new_n307), .A3(new_n393), .ZN(new_n394));
  AOI21_X1  g0194(.A(new_n393), .B1(new_n305), .B2(new_n307), .ZN(new_n395));
  OAI21_X1  g0195(.A(new_n212), .B1(new_n394), .B2(new_n395), .ZN(new_n396));
  AOI21_X1  g0196(.A(new_n392), .B1(new_n396), .B2(new_n391), .ZN(new_n397));
  OAI211_X1 g0197(.A(KEYINPUT16), .B(new_n390), .C1(new_n397), .C2(new_n203), .ZN(new_n398));
  INV_X1    g0198(.A(KEYINPUT16), .ZN(new_n399));
  OAI21_X1  g0199(.A(G20), .B1(new_n206), .B2(new_n388), .ZN(new_n400));
  INV_X1    g0200(.A(G159), .ZN(new_n401));
  OAI21_X1  g0201(.A(new_n400), .B1(new_n401), .B2(new_n320), .ZN(new_n402));
  OAI21_X1  g0202(.A(new_n391), .B1(new_n272), .B2(G20), .ZN(new_n403));
  NAND3_X1  g0203(.A1(new_n308), .A2(KEYINPUT7), .A3(new_n212), .ZN(new_n404));
  AOI21_X1  g0204(.A(new_n203), .B1(new_n403), .B2(new_n404), .ZN(new_n405));
  OAI21_X1  g0205(.A(new_n399), .B1(new_n402), .B2(new_n405), .ZN(new_n406));
  NAND3_X1  g0206(.A1(new_n398), .A2(new_n267), .A3(new_n406), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n261), .A2(new_n251), .ZN(new_n408));
  OAI21_X1  g0208(.A(new_n408), .B1(new_n269), .B2(new_n261), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n407), .A2(new_n409), .ZN(new_n410));
  OAI21_X1  g0210(.A(KEYINPUT78), .B1(new_n285), .B2(new_n233), .ZN(new_n411));
  INV_X1    g0211(.A(KEYINPUT78), .ZN(new_n412));
  NAND4_X1  g0212(.A1(new_n279), .A2(new_n282), .A3(new_n412), .A4(G232), .ZN(new_n413));
  NAND3_X1  g0213(.A1(new_n411), .A2(new_n302), .A3(new_n413), .ZN(new_n414));
  INV_X1    g0214(.A(KEYINPUT79), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n414), .A2(new_n415), .ZN(new_n416));
  NAND4_X1  g0216(.A1(new_n411), .A2(KEYINPUT79), .A3(new_n302), .A4(new_n413), .ZN(new_n417));
  NAND4_X1  g0217(.A1(new_n305), .A2(new_n307), .A3(G223), .A4(new_n364), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n418), .A2(KEYINPUT77), .ZN(new_n419));
  INV_X1    g0219(.A(KEYINPUT77), .ZN(new_n420));
  NAND4_X1  g0220(.A1(new_n272), .A2(new_n420), .A3(G223), .A4(new_n364), .ZN(new_n421));
  NAND3_X1  g0221(.A1(new_n272), .A2(G226), .A3(G1698), .ZN(new_n422));
  NAND2_X1  g0222(.A1(G33), .A2(G87), .ZN(new_n423));
  NAND4_X1  g0223(.A1(new_n419), .A2(new_n421), .A3(new_n422), .A4(new_n423), .ZN(new_n424));
  AOI22_X1  g0224(.A1(new_n416), .A2(new_n417), .B1(new_n280), .B2(new_n424), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n424), .A2(new_n280), .ZN(new_n426));
  AND2_X1   g0226(.A1(new_n411), .A2(new_n413), .ZN(new_n427));
  NAND3_X1  g0227(.A1(new_n426), .A2(new_n302), .A3(new_n427), .ZN(new_n428));
  AOI22_X1  g0228(.A1(new_n425), .A2(new_n314), .B1(new_n428), .B2(new_n299), .ZN(new_n429));
  OAI21_X1  g0229(.A(KEYINPUT17), .B1(new_n410), .B2(new_n429), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n428), .A2(new_n299), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n416), .A2(new_n417), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n432), .A2(new_n426), .ZN(new_n433));
  OAI21_X1  g0233(.A(new_n431), .B1(new_n433), .B2(G190), .ZN(new_n434));
  INV_X1    g0234(.A(KEYINPUT17), .ZN(new_n435));
  NAND4_X1  g0235(.A1(new_n434), .A2(new_n435), .A3(new_n407), .A4(new_n409), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n430), .A2(new_n436), .ZN(new_n437));
  INV_X1    g0237(.A(KEYINPUT80), .ZN(new_n438));
  INV_X1    g0238(.A(KEYINPUT18), .ZN(new_n439));
  AOI22_X1  g0239(.A1(new_n425), .A2(new_n290), .B1(new_n428), .B2(new_n339), .ZN(new_n440));
  AOI211_X1 g0240(.A(new_n438), .B(new_n439), .C1(new_n410), .C2(new_n440), .ZN(new_n441));
  NAND2_X1  g0241(.A1(new_n438), .A2(new_n439), .ZN(new_n442));
  NAND2_X1  g0242(.A1(KEYINPUT80), .A2(KEYINPUT18), .ZN(new_n443));
  NAND4_X1  g0243(.A1(new_n410), .A2(new_n440), .A3(new_n442), .A4(new_n443), .ZN(new_n444));
  INV_X1    g0244(.A(new_n444), .ZN(new_n445));
  NOR2_X1   g0245(.A1(new_n441), .A2(new_n445), .ZN(new_n446));
  OAI211_X1 g0246(.A(new_n437), .B(new_n446), .C1(new_n342), .C2(new_n343), .ZN(new_n447));
  NOR2_X1   g0247(.A1(new_n387), .A2(new_n447), .ZN(new_n448));
  NAND4_X1  g0248(.A1(new_n305), .A2(new_n307), .A3(G244), .A4(G1698), .ZN(new_n449));
  NAND4_X1  g0249(.A1(new_n305), .A2(new_n307), .A3(G238), .A4(new_n364), .ZN(new_n450));
  NOR2_X1   g0250(.A1(new_n304), .A2(new_n225), .ZN(new_n451));
  INV_X1    g0251(.A(new_n451), .ZN(new_n452));
  NAND3_X1  g0252(.A1(new_n449), .A2(new_n450), .A3(new_n452), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n453), .A2(KEYINPUT85), .ZN(new_n454));
  INV_X1    g0254(.A(KEYINPUT85), .ZN(new_n455));
  NAND4_X1  g0255(.A1(new_n449), .A2(new_n450), .A3(new_n455), .A4(new_n452), .ZN(new_n456));
  NAND3_X1  g0256(.A1(new_n454), .A2(new_n280), .A3(new_n456), .ZN(new_n457));
  INV_X1    g0257(.A(G45), .ZN(new_n458));
  NOR2_X1   g0258(.A1(new_n458), .A2(G1), .ZN(new_n459));
  NOR2_X1   g0259(.A1(new_n280), .A2(new_n459), .ZN(new_n460));
  AOI22_X1  g0260(.A1(new_n460), .A2(G250), .B1(G274), .B2(new_n459), .ZN(new_n461));
  AND3_X1   g0261(.A1(new_n457), .A2(KEYINPUT86), .A3(new_n461), .ZN(new_n462));
  AOI21_X1  g0262(.A(KEYINPUT86), .B1(new_n457), .B2(new_n461), .ZN(new_n463));
  OAI21_X1  g0263(.A(new_n290), .B1(new_n462), .B2(new_n463), .ZN(new_n464));
  NAND2_X1  g0264(.A1(new_n457), .A2(new_n461), .ZN(new_n465));
  INV_X1    g0265(.A(KEYINPUT86), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  NAND3_X1  g0267(.A1(new_n457), .A2(KEYINPUT86), .A3(new_n461), .ZN(new_n468));
  NAND3_X1  g0268(.A1(new_n467), .A2(new_n339), .A3(new_n468), .ZN(new_n469));
  NAND3_X1  g0269(.A1(new_n272), .A2(new_n212), .A3(G68), .ZN(new_n470));
  INV_X1    g0270(.A(KEYINPUT19), .ZN(new_n471));
  OAI21_X1  g0271(.A(new_n212), .B1(new_n366), .B2(new_n471), .ZN(new_n472));
  NOR2_X1   g0272(.A1(G97), .A2(G107), .ZN(new_n473));
  INV_X1    g0273(.A(G87), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n473), .A2(new_n474), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n472), .A2(new_n475), .ZN(new_n476));
  OAI21_X1  g0276(.A(new_n471), .B1(new_n366), .B2(G20), .ZN(new_n477));
  NAND3_X1  g0277(.A1(new_n470), .A2(new_n476), .A3(new_n477), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n478), .A2(new_n267), .ZN(new_n479));
  INV_X1    g0279(.A(new_n253), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n480), .A2(new_n323), .ZN(new_n481));
  INV_X1    g0281(.A(new_n267), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n215), .A2(G33), .ZN(new_n483));
  NAND3_X1  g0283(.A1(new_n482), .A2(new_n251), .A3(new_n483), .ZN(new_n484));
  OAI211_X1 g0284(.A(new_n479), .B(new_n481), .C1(new_n480), .C2(new_n484), .ZN(new_n485));
  NAND3_X1  g0285(.A1(new_n464), .A2(new_n469), .A3(new_n485), .ZN(new_n486));
  OAI21_X1  g0286(.A(G190), .B1(new_n462), .B2(new_n463), .ZN(new_n487));
  NAND3_X1  g0287(.A1(new_n467), .A2(G200), .A3(new_n468), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n479), .A2(new_n481), .ZN(new_n489));
  INV_X1    g0289(.A(new_n484), .ZN(new_n490));
  AOI21_X1  g0290(.A(new_n489), .B1(G87), .B2(new_n490), .ZN(new_n491));
  NAND3_X1  g0291(.A1(new_n487), .A2(new_n488), .A3(new_n491), .ZN(new_n492));
  INV_X1    g0292(.A(KEYINPUT87), .ZN(new_n493));
  AND3_X1   g0293(.A1(new_n486), .A2(new_n492), .A3(new_n493), .ZN(new_n494));
  AOI21_X1  g0294(.A(new_n493), .B1(new_n486), .B2(new_n492), .ZN(new_n495));
  NOR2_X1   g0295(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  INV_X1    g0296(.A(KEYINPUT24), .ZN(new_n497));
  NAND4_X1  g0297(.A1(new_n305), .A2(new_n307), .A3(new_n212), .A4(G87), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n498), .A2(KEYINPUT22), .ZN(new_n499));
  INV_X1    g0299(.A(KEYINPUT22), .ZN(new_n500));
  NAND4_X1  g0300(.A1(new_n272), .A2(new_n500), .A3(new_n212), .A4(G87), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n499), .A2(new_n501), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n451), .A2(new_n212), .ZN(new_n503));
  NOR2_X1   g0303(.A1(new_n212), .A2(G107), .ZN(new_n504));
  XNOR2_X1  g0304(.A(new_n504), .B(KEYINPUT23), .ZN(new_n505));
  AND4_X1   g0305(.A1(new_n497), .A2(new_n502), .A3(new_n503), .A4(new_n505), .ZN(new_n506));
  AOI22_X1  g0306(.A1(new_n499), .A2(new_n501), .B1(new_n212), .B2(new_n451), .ZN(new_n507));
  AOI21_X1  g0307(.A(new_n497), .B1(new_n507), .B2(new_n505), .ZN(new_n508));
  OAI21_X1  g0308(.A(new_n267), .B1(new_n506), .B2(new_n508), .ZN(new_n509));
  NOR2_X1   g0309(.A1(new_n484), .A2(new_n247), .ZN(new_n510));
  INV_X1    g0310(.A(new_n510), .ZN(new_n511));
  NOR2_X1   g0311(.A1(new_n251), .A2(G107), .ZN(new_n512));
  XNOR2_X1  g0312(.A(new_n512), .B(KEYINPUT25), .ZN(new_n513));
  NAND3_X1  g0313(.A1(new_n509), .A2(new_n511), .A3(new_n513), .ZN(new_n514));
  NAND4_X1  g0314(.A1(new_n305), .A2(new_n307), .A3(G257), .A4(G1698), .ZN(new_n515));
  NAND4_X1  g0315(.A1(new_n305), .A2(new_n307), .A3(G250), .A4(new_n364), .ZN(new_n516));
  NAND2_X1  g0316(.A1(G33), .A2(G294), .ZN(new_n517));
  NAND3_X1  g0317(.A1(new_n515), .A2(new_n516), .A3(new_n517), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n518), .A2(new_n280), .ZN(new_n519));
  INV_X1    g0319(.A(G41), .ZN(new_n520));
  OAI211_X1 g0320(.A(new_n215), .B(G45), .C1(new_n520), .C2(KEYINPUT5), .ZN(new_n521));
  INV_X1    g0321(.A(KEYINPUT5), .ZN(new_n522));
  NOR2_X1   g0322(.A1(new_n522), .A2(G41), .ZN(new_n523));
  OAI211_X1 g0323(.A(G264), .B(new_n279), .C1(new_n521), .C2(new_n523), .ZN(new_n524));
  INV_X1    g0324(.A(KEYINPUT84), .ZN(new_n525));
  OAI21_X1  g0325(.A(new_n525), .B1(new_n522), .B2(G41), .ZN(new_n526));
  NAND3_X1  g0326(.A1(new_n520), .A2(KEYINPUT84), .A3(KEYINPUT5), .ZN(new_n527));
  AOI21_X1  g0327(.A(new_n283), .B1(new_n526), .B2(new_n527), .ZN(new_n528));
  INV_X1    g0328(.A(KEYINPUT83), .ZN(new_n529));
  NOR2_X1   g0329(.A1(new_n521), .A2(new_n529), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n522), .A2(G41), .ZN(new_n531));
  AOI21_X1  g0331(.A(KEYINPUT83), .B1(new_n459), .B2(new_n531), .ZN(new_n532));
  OAI211_X1 g0332(.A(new_n279), .B(new_n528), .C1(new_n530), .C2(new_n532), .ZN(new_n533));
  NAND3_X1  g0333(.A1(new_n519), .A2(new_n524), .A3(new_n533), .ZN(new_n534));
  NAND2_X1  g0334(.A1(new_n534), .A2(new_n339), .ZN(new_n535));
  OR2_X1    g0335(.A1(new_n534), .A2(G179), .ZN(new_n536));
  NAND3_X1  g0336(.A1(new_n514), .A2(new_n535), .A3(new_n536), .ZN(new_n537));
  NAND3_X1  g0337(.A1(new_n502), .A2(new_n503), .A3(new_n505), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n538), .A2(KEYINPUT24), .ZN(new_n539));
  NAND3_X1  g0339(.A1(new_n507), .A2(new_n497), .A3(new_n505), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  AOI21_X1  g0341(.A(new_n510), .B1(new_n541), .B2(new_n267), .ZN(new_n542));
  NAND4_X1  g0342(.A1(new_n519), .A2(new_n314), .A3(new_n533), .A4(new_n524), .ZN(new_n543));
  NOR2_X1   g0343(.A1(new_n543), .A2(KEYINPUT90), .ZN(new_n544));
  INV_X1    g0344(.A(new_n544), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n534), .A2(new_n299), .ZN(new_n546));
  NAND3_X1  g0346(.A1(new_n546), .A2(KEYINPUT90), .A3(new_n543), .ZN(new_n547));
  NAND4_X1  g0347(.A1(new_n542), .A2(new_n545), .A3(new_n513), .A4(new_n547), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n537), .A2(new_n548), .ZN(new_n549));
  INV_X1    g0349(.A(KEYINPUT91), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  NAND3_X1  g0351(.A1(new_n537), .A2(new_n548), .A3(KEYINPUT91), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  NAND4_X1  g0353(.A1(new_n215), .A2(new_n225), .A3(G13), .A4(G20), .ZN(new_n554));
  XNOR2_X1  g0354(.A(new_n554), .B(KEYINPUT88), .ZN(new_n555));
  NAND4_X1  g0355(.A1(new_n482), .A2(G116), .A3(new_n251), .A4(new_n483), .ZN(new_n556));
  AOI22_X1  g0356(.A1(new_n266), .A2(new_n211), .B1(G20), .B2(new_n225), .ZN(new_n557));
  NAND2_X1  g0357(.A1(G33), .A2(G283), .ZN(new_n558));
  INV_X1    g0358(.A(G97), .ZN(new_n559));
  OAI211_X1 g0359(.A(new_n558), .B(new_n212), .C1(G33), .C2(new_n559), .ZN(new_n560));
  AND3_X1   g0360(.A1(new_n557), .A2(KEYINPUT20), .A3(new_n560), .ZN(new_n561));
  AOI21_X1  g0361(.A(KEYINPUT20), .B1(new_n557), .B2(new_n560), .ZN(new_n562));
  OAI211_X1 g0362(.A(new_n555), .B(new_n556), .C1(new_n561), .C2(new_n562), .ZN(new_n563));
  NAND4_X1  g0363(.A1(new_n305), .A2(new_n307), .A3(G257), .A4(new_n364), .ZN(new_n564));
  NAND4_X1  g0364(.A1(new_n305), .A2(new_n307), .A3(G264), .A4(G1698), .ZN(new_n565));
  INV_X1    g0365(.A(G303), .ZN(new_n566));
  OAI211_X1 g0366(.A(new_n564), .B(new_n565), .C1(new_n566), .C2(new_n272), .ZN(new_n567));
  AND2_X1   g0367(.A1(new_n567), .A2(new_n280), .ZN(new_n568));
  OAI211_X1 g0368(.A(G270), .B(new_n279), .C1(new_n521), .C2(new_n523), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n533), .A2(new_n569), .ZN(new_n570));
  OAI211_X1 g0370(.A(G169), .B(new_n563), .C1(new_n568), .C2(new_n570), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n571), .A2(KEYINPUT89), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n567), .A2(new_n280), .ZN(new_n573));
  NAND3_X1  g0373(.A1(new_n573), .A2(new_n533), .A3(new_n569), .ZN(new_n574));
  INV_X1    g0374(.A(KEYINPUT89), .ZN(new_n575));
  NAND4_X1  g0375(.A1(new_n574), .A2(new_n575), .A3(G169), .A4(new_n563), .ZN(new_n576));
  INV_X1    g0376(.A(KEYINPUT21), .ZN(new_n577));
  NAND3_X1  g0377(.A1(new_n572), .A2(new_n576), .A3(new_n577), .ZN(new_n578));
  OAI211_X1 g0378(.A(KEYINPUT21), .B(G169), .C1(new_n568), .C2(new_n570), .ZN(new_n579));
  NAND4_X1  g0379(.A1(new_n573), .A2(G179), .A3(new_n533), .A4(new_n569), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n581), .A2(new_n563), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n578), .A2(new_n582), .ZN(new_n583));
  INV_X1    g0383(.A(new_n583), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n574), .A2(G200), .ZN(new_n585));
  INV_X1    g0385(.A(new_n563), .ZN(new_n586));
  OAI211_X1 g0386(.A(new_n585), .B(new_n586), .C1(new_n314), .C2(new_n574), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n584), .A2(new_n587), .ZN(new_n588));
  AOI21_X1  g0388(.A(KEYINPUT7), .B1(new_n308), .B2(new_n212), .ZN(new_n589));
  OAI21_X1  g0389(.A(G107), .B1(new_n392), .B2(new_n589), .ZN(new_n590));
  NAND3_X1  g0390(.A1(new_n247), .A2(KEYINPUT6), .A3(G97), .ZN(new_n591));
  XOR2_X1   g0391(.A(G97), .B(G107), .Z(new_n592));
  OAI21_X1  g0392(.A(new_n591), .B1(new_n592), .B2(KEYINPUT6), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n593), .A2(G20), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n260), .A2(G77), .ZN(new_n595));
  NAND3_X1  g0395(.A1(new_n590), .A2(new_n594), .A3(new_n595), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n596), .A2(new_n267), .ZN(new_n597));
  NOR2_X1   g0397(.A1(new_n251), .A2(G97), .ZN(new_n598));
  NOR2_X1   g0398(.A1(new_n598), .A2(KEYINPUT81), .ZN(new_n599));
  INV_X1    g0399(.A(new_n599), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n598), .A2(KEYINPUT81), .ZN(new_n601));
  OAI21_X1  g0401(.A(new_n601), .B1(new_n484), .B2(new_n559), .ZN(new_n602));
  INV_X1    g0402(.A(new_n602), .ZN(new_n603));
  NAND3_X1  g0403(.A1(new_n597), .A2(new_n600), .A3(new_n603), .ZN(new_n604));
  NAND4_X1  g0404(.A1(new_n305), .A2(new_n307), .A3(G244), .A4(new_n364), .ZN(new_n605));
  NAND2_X1  g0405(.A1(KEYINPUT82), .A2(KEYINPUT4), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n605), .A2(new_n606), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n607), .A2(new_n558), .ZN(new_n608));
  NAND4_X1  g0408(.A1(new_n305), .A2(new_n307), .A3(G250), .A4(G1698), .ZN(new_n609));
  OR2_X1    g0409(.A1(KEYINPUT82), .A2(KEYINPUT4), .ZN(new_n610));
  OAI211_X1 g0410(.A(new_n609), .B(new_n610), .C1(new_n605), .C2(new_n606), .ZN(new_n611));
  OAI21_X1  g0411(.A(new_n280), .B1(new_n608), .B2(new_n611), .ZN(new_n612));
  OAI211_X1 g0412(.A(G257), .B(new_n279), .C1(new_n521), .C2(new_n523), .ZN(new_n613));
  NAND3_X1  g0413(.A1(new_n612), .A2(new_n533), .A3(new_n613), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n614), .A2(new_n339), .ZN(new_n615));
  NAND4_X1  g0415(.A1(new_n612), .A2(new_n290), .A3(new_n533), .A4(new_n613), .ZN(new_n616));
  NAND3_X1  g0416(.A1(new_n604), .A2(new_n615), .A3(new_n616), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n614), .A2(G200), .ZN(new_n618));
  AOI21_X1  g0418(.A(new_n602), .B1(new_n596), .B2(new_n267), .ZN(new_n619));
  NAND4_X1  g0419(.A1(new_n612), .A2(G190), .A3(new_n533), .A4(new_n613), .ZN(new_n620));
  NAND4_X1  g0420(.A1(new_n618), .A2(new_n600), .A3(new_n619), .A4(new_n620), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n617), .A2(new_n621), .ZN(new_n622));
  NOR2_X1   g0422(.A1(new_n588), .A2(new_n622), .ZN(new_n623));
  AND4_X1   g0423(.A1(new_n448), .A2(new_n496), .A3(new_n553), .A4(new_n623), .ZN(G372));
  OR2_X1    g0424(.A1(new_n297), .A2(new_n378), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n384), .A2(new_n385), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n627), .A2(new_n437), .ZN(new_n628));
  INV_X1    g0428(.A(KEYINPUT94), .ZN(new_n629));
  AND3_X1   g0429(.A1(new_n410), .A2(new_n629), .A3(new_n440), .ZN(new_n630));
  AOI21_X1  g0430(.A(new_n629), .B1(new_n410), .B2(new_n440), .ZN(new_n631));
  OAI21_X1  g0431(.A(new_n439), .B1(new_n630), .B2(new_n631), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n410), .A2(new_n440), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n633), .A2(KEYINPUT94), .ZN(new_n634));
  NAND3_X1  g0434(.A1(new_n410), .A2(new_n629), .A3(new_n440), .ZN(new_n635));
  NAND3_X1  g0435(.A1(new_n634), .A2(KEYINPUT18), .A3(new_n635), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n632), .A2(new_n636), .ZN(new_n637));
  INV_X1    g0437(.A(new_n637), .ZN(new_n638));
  INV_X1    g0438(.A(KEYINPUT95), .ZN(new_n639));
  NAND3_X1  g0439(.A1(new_n628), .A2(new_n638), .A3(new_n639), .ZN(new_n640));
  AOI22_X1  g0440(.A1(new_n625), .A2(new_n626), .B1(new_n430), .B2(new_n436), .ZN(new_n641));
  OAI21_X1  g0441(.A(KEYINPUT95), .B1(new_n641), .B2(new_n637), .ZN(new_n642));
  AND2_X1   g0442(.A1(new_n332), .A2(new_n338), .ZN(new_n643));
  NAND3_X1  g0443(.A1(new_n640), .A2(new_n642), .A3(new_n643), .ZN(new_n644));
  AND2_X1   g0444(.A1(new_n644), .A2(new_n341), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n465), .A2(new_n339), .ZN(new_n646));
  NAND3_X1  g0446(.A1(new_n464), .A2(new_n485), .A3(new_n646), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n465), .A2(G200), .ZN(new_n648));
  NAND3_X1  g0448(.A1(new_n487), .A2(new_n491), .A3(new_n648), .ZN(new_n649));
  INV_X1    g0449(.A(new_n617), .ZN(new_n650));
  INV_X1    g0450(.A(KEYINPUT26), .ZN(new_n651));
  NAND4_X1  g0451(.A1(new_n647), .A2(new_n649), .A3(new_n650), .A4(new_n651), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n652), .A2(new_n647), .ZN(new_n653));
  INV_X1    g0453(.A(new_n653), .ZN(new_n654));
  NOR3_X1   g0454(.A1(new_n494), .A2(new_n495), .A3(new_n617), .ZN(new_n655));
  OAI21_X1  g0455(.A(new_n654), .B1(new_n655), .B2(new_n651), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n647), .A2(new_n649), .ZN(new_n657));
  NAND4_X1  g0457(.A1(new_n547), .A2(new_n509), .A3(new_n511), .A4(new_n513), .ZN(new_n658));
  OAI211_X1 g0458(.A(new_n617), .B(new_n621), .C1(new_n658), .C2(new_n544), .ZN(new_n659));
  NOR2_X1   g0459(.A1(new_n657), .A2(new_n659), .ZN(new_n660));
  INV_X1    g0460(.A(KEYINPUT92), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n583), .A2(new_n661), .ZN(new_n662));
  NAND3_X1  g0462(.A1(new_n578), .A2(KEYINPUT92), .A3(new_n582), .ZN(new_n663));
  NAND3_X1  g0463(.A1(new_n662), .A2(new_n537), .A3(new_n663), .ZN(new_n664));
  INV_X1    g0464(.A(KEYINPUT93), .ZN(new_n665));
  AND3_X1   g0465(.A1(new_n660), .A2(new_n664), .A3(new_n665), .ZN(new_n666));
  AOI21_X1  g0466(.A(new_n665), .B1(new_n660), .B2(new_n664), .ZN(new_n667));
  NOR2_X1   g0467(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  OAI21_X1  g0468(.A(new_n448), .B1(new_n656), .B2(new_n668), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n645), .A2(new_n669), .ZN(G369));
  XOR2_X1   g0470(.A(KEYINPUT96), .B(KEYINPUT27), .Z(new_n671));
  INV_X1    g0471(.A(G13), .ZN(new_n672));
  NOR3_X1   g0472(.A1(new_n672), .A2(G1), .A3(G20), .ZN(new_n673));
  OR2_X1    g0473(.A1(new_n671), .A2(new_n673), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n671), .A2(new_n673), .ZN(new_n675));
  NAND3_X1  g0475(.A1(new_n674), .A2(G213), .A3(new_n675), .ZN(new_n676));
  INV_X1    g0476(.A(G343), .ZN(new_n677));
  NOR2_X1   g0477(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  NOR2_X1   g0478(.A1(new_n537), .A2(new_n678), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n514), .A2(new_n678), .ZN(new_n680));
  INV_X1    g0480(.A(new_n680), .ZN(new_n681));
  AOI21_X1  g0481(.A(new_n681), .B1(new_n551), .B2(new_n552), .ZN(new_n682));
  INV_X1    g0482(.A(new_n678), .ZN(new_n683));
  NOR2_X1   g0483(.A1(new_n537), .A2(new_n683), .ZN(new_n684));
  OAI21_X1  g0484(.A(KEYINPUT97), .B1(new_n682), .B2(new_n684), .ZN(new_n685));
  AND3_X1   g0485(.A1(new_n537), .A2(new_n548), .A3(KEYINPUT91), .ZN(new_n686));
  AOI21_X1  g0486(.A(KEYINPUT91), .B1(new_n537), .B2(new_n548), .ZN(new_n687));
  OAI21_X1  g0487(.A(new_n680), .B1(new_n686), .B2(new_n687), .ZN(new_n688));
  INV_X1    g0488(.A(KEYINPUT97), .ZN(new_n689));
  INV_X1    g0489(.A(new_n684), .ZN(new_n690));
  NAND3_X1  g0490(.A1(new_n688), .A2(new_n689), .A3(new_n690), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n685), .A2(new_n691), .ZN(new_n692));
  NOR2_X1   g0492(.A1(new_n584), .A2(new_n678), .ZN(new_n693));
  AOI21_X1  g0493(.A(new_n679), .B1(new_n692), .B2(new_n693), .ZN(new_n694));
  NOR2_X1   g0494(.A1(new_n683), .A2(new_n586), .ZN(new_n695));
  OR2_X1    g0495(.A1(new_n588), .A2(new_n695), .ZN(new_n696));
  NAND2_X1  g0496(.A1(new_n662), .A2(new_n663), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n697), .A2(new_n695), .ZN(new_n698));
  NAND2_X1  g0498(.A1(new_n696), .A2(new_n698), .ZN(new_n699));
  INV_X1    g0499(.A(new_n699), .ZN(new_n700));
  INV_X1    g0500(.A(G330), .ZN(new_n701));
  NOR2_X1   g0501(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  NAND2_X1  g0502(.A1(new_n702), .A2(new_n692), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n694), .A2(new_n703), .ZN(G399));
  INV_X1    g0504(.A(new_n216), .ZN(new_n705));
  NOR2_X1   g0505(.A1(new_n705), .A2(G41), .ZN(new_n706));
  INV_X1    g0506(.A(new_n706), .ZN(new_n707));
  NOR2_X1   g0507(.A1(new_n475), .A2(G116), .ZN(new_n708));
  NAND3_X1  g0508(.A1(new_n707), .A2(G1), .A3(new_n708), .ZN(new_n709));
  OAI21_X1  g0509(.A(new_n709), .B1(new_n210), .B2(new_n707), .ZN(new_n710));
  XNOR2_X1  g0510(.A(new_n710), .B(KEYINPUT28), .ZN(new_n711));
  OAI21_X1  g0511(.A(new_n683), .B1(new_n668), .B2(new_n656), .ZN(new_n712));
  INV_X1    g0512(.A(KEYINPUT29), .ZN(new_n713));
  NAND2_X1  g0513(.A1(new_n712), .A2(new_n713), .ZN(new_n714));
  INV_X1    g0514(.A(new_n647), .ZN(new_n715));
  NAND2_X1  g0515(.A1(new_n584), .A2(new_n537), .ZN(new_n716));
  AOI21_X1  g0516(.A(new_n715), .B1(new_n660), .B2(new_n716), .ZN(new_n717));
  OAI21_X1  g0517(.A(KEYINPUT26), .B1(new_n657), .B2(new_n617), .ZN(new_n718));
  NAND2_X1  g0518(.A1(new_n486), .A2(new_n492), .ZN(new_n719));
  NAND2_X1  g0519(.A1(new_n719), .A2(KEYINPUT87), .ZN(new_n720));
  NAND3_X1  g0520(.A1(new_n486), .A2(new_n492), .A3(new_n493), .ZN(new_n721));
  NAND4_X1  g0521(.A1(new_n720), .A2(new_n651), .A3(new_n721), .A4(new_n650), .ZN(new_n722));
  NAND3_X1  g0522(.A1(new_n717), .A2(new_n718), .A3(new_n722), .ZN(new_n723));
  NAND3_X1  g0523(.A1(new_n723), .A2(KEYINPUT29), .A3(new_n683), .ZN(new_n724));
  NAND2_X1  g0524(.A1(new_n724), .A2(KEYINPUT99), .ZN(new_n725));
  INV_X1    g0525(.A(KEYINPUT99), .ZN(new_n726));
  NAND4_X1  g0526(.A1(new_n723), .A2(new_n726), .A3(KEYINPUT29), .A4(new_n683), .ZN(new_n727));
  NAND3_X1  g0527(.A1(new_n714), .A2(new_n725), .A3(new_n727), .ZN(new_n728));
  NAND4_X1  g0528(.A1(new_n496), .A2(new_n553), .A3(new_n623), .A4(new_n683), .ZN(new_n729));
  AND2_X1   g0529(.A1(new_n612), .A2(new_n613), .ZN(new_n730));
  NOR2_X1   g0530(.A1(new_n580), .A2(new_n534), .ZN(new_n731));
  OAI211_X1 g0531(.A(new_n730), .B(new_n731), .C1(new_n462), .C2(new_n463), .ZN(new_n732));
  INV_X1    g0532(.A(KEYINPUT30), .ZN(new_n733));
  NAND2_X1  g0533(.A1(new_n732), .A2(new_n733), .ZN(new_n734));
  NAND2_X1  g0534(.A1(new_n467), .A2(new_n468), .ZN(new_n735));
  NAND4_X1  g0535(.A1(new_n735), .A2(KEYINPUT30), .A3(new_n730), .A4(new_n731), .ZN(new_n736));
  AND2_X1   g0536(.A1(new_n614), .A2(new_n290), .ZN(new_n737));
  NAND4_X1  g0537(.A1(new_n737), .A2(new_n465), .A3(new_n534), .A4(new_n574), .ZN(new_n738));
  NAND3_X1  g0538(.A1(new_n734), .A2(new_n736), .A3(new_n738), .ZN(new_n739));
  NAND2_X1  g0539(.A1(new_n739), .A2(new_n678), .ZN(new_n740));
  INV_X1    g0540(.A(KEYINPUT31), .ZN(new_n741));
  NAND3_X1  g0541(.A1(new_n740), .A2(KEYINPUT98), .A3(new_n741), .ZN(new_n742));
  NAND3_X1  g0542(.A1(new_n739), .A2(KEYINPUT31), .A3(new_n678), .ZN(new_n743));
  NAND2_X1  g0543(.A1(new_n740), .A2(new_n741), .ZN(new_n744));
  INV_X1    g0544(.A(KEYINPUT98), .ZN(new_n745));
  NAND2_X1  g0545(.A1(new_n744), .A2(new_n745), .ZN(new_n746));
  NAND4_X1  g0546(.A1(new_n729), .A2(new_n742), .A3(new_n743), .A4(new_n746), .ZN(new_n747));
  NAND2_X1  g0547(.A1(new_n747), .A2(G330), .ZN(new_n748));
  NAND2_X1  g0548(.A1(new_n728), .A2(new_n748), .ZN(new_n749));
  INV_X1    g0549(.A(new_n749), .ZN(new_n750));
  OAI21_X1  g0550(.A(new_n711), .B1(new_n750), .B2(G1), .ZN(G364));
  INV_X1    g0551(.A(new_n702), .ZN(new_n752));
  NOR2_X1   g0552(.A1(new_n672), .A2(G20), .ZN(new_n753));
  NAND2_X1  g0553(.A1(new_n753), .A2(G45), .ZN(new_n754));
  NAND3_X1  g0554(.A1(new_n707), .A2(G1), .A3(new_n754), .ZN(new_n755));
  NAND2_X1  g0555(.A1(new_n700), .A2(new_n701), .ZN(new_n756));
  NAND3_X1  g0556(.A1(new_n752), .A2(new_n755), .A3(new_n756), .ZN(new_n757));
  INV_X1    g0557(.A(new_n755), .ZN(new_n758));
  NAND2_X1  g0558(.A1(new_n244), .A2(G45), .ZN(new_n759));
  NOR2_X1   g0559(.A1(new_n394), .A2(new_n395), .ZN(new_n760));
  NOR2_X1   g0560(.A1(new_n760), .A2(new_n705), .ZN(new_n761));
  OAI211_X1 g0561(.A(new_n759), .B(new_n761), .C1(G45), .C2(new_n210), .ZN(new_n762));
  XNOR2_X1  g0562(.A(G355), .B(KEYINPUT100), .ZN(new_n763));
  NAND3_X1  g0563(.A1(new_n763), .A2(new_n216), .A3(new_n272), .ZN(new_n764));
  OAI211_X1 g0564(.A(new_n762), .B(new_n764), .C1(G116), .C2(new_n216), .ZN(new_n765));
  INV_X1    g0565(.A(KEYINPUT101), .ZN(new_n766));
  AND2_X1   g0566(.A1(new_n765), .A2(new_n766), .ZN(new_n767));
  NOR2_X1   g0567(.A1(G13), .A2(G33), .ZN(new_n768));
  INV_X1    g0568(.A(new_n768), .ZN(new_n769));
  NOR2_X1   g0569(.A1(new_n769), .A2(G20), .ZN(new_n770));
  AOI21_X1  g0570(.A(new_n211), .B1(G20), .B2(new_n339), .ZN(new_n771));
  NOR2_X1   g0571(.A1(new_n770), .A2(new_n771), .ZN(new_n772));
  OAI21_X1  g0572(.A(new_n772), .B1(new_n765), .B2(new_n766), .ZN(new_n773));
  OAI21_X1  g0573(.A(new_n758), .B1(new_n767), .B2(new_n773), .ZN(new_n774));
  XOR2_X1   g0574(.A(new_n774), .B(KEYINPUT102), .Z(new_n775));
  NOR2_X1   g0575(.A1(new_n212), .A2(G190), .ZN(new_n776));
  NOR2_X1   g0576(.A1(G179), .A2(G200), .ZN(new_n777));
  NAND2_X1  g0577(.A1(new_n776), .A2(new_n777), .ZN(new_n778));
  INV_X1    g0578(.A(new_n778), .ZN(new_n779));
  NAND2_X1  g0579(.A1(new_n779), .A2(G159), .ZN(new_n780));
  XNOR2_X1  g0580(.A(new_n780), .B(KEYINPUT32), .ZN(new_n781));
  NOR2_X1   g0581(.A1(new_n299), .A2(G179), .ZN(new_n782));
  NAND2_X1  g0582(.A1(new_n782), .A2(new_n776), .ZN(new_n783));
  NOR2_X1   g0583(.A1(new_n212), .A2(new_n314), .ZN(new_n784));
  NOR2_X1   g0584(.A1(new_n290), .A2(G200), .ZN(new_n785));
  NAND2_X1  g0585(.A1(new_n784), .A2(new_n785), .ZN(new_n786));
  OAI221_X1 g0586(.A(new_n272), .B1(new_n783), .B2(new_n247), .C1(new_n202), .C2(new_n786), .ZN(new_n787));
  NOR2_X1   g0587(.A1(new_n212), .A2(new_n290), .ZN(new_n788));
  NAND3_X1  g0588(.A1(new_n788), .A2(new_n314), .A3(G200), .ZN(new_n789));
  AOI21_X1  g0589(.A(new_n212), .B1(new_n777), .B2(G190), .ZN(new_n790));
  OAI22_X1  g0590(.A1(new_n789), .A2(new_n203), .B1(new_n790), .B2(new_n559), .ZN(new_n791));
  NOR2_X1   g0591(.A1(new_n787), .A2(new_n791), .ZN(new_n792));
  NAND2_X1  g0592(.A1(new_n776), .A2(new_n785), .ZN(new_n793));
  AND2_X1   g0593(.A1(new_n784), .A2(new_n782), .ZN(new_n794));
  OR2_X1    g0594(.A1(new_n794), .A2(KEYINPUT104), .ZN(new_n795));
  NAND2_X1  g0595(.A1(new_n794), .A2(KEYINPUT104), .ZN(new_n796));
  NAND2_X1  g0596(.A1(new_n795), .A2(new_n796), .ZN(new_n797));
  OAI221_X1 g0597(.A(new_n792), .B1(new_n255), .B2(new_n793), .C1(new_n474), .C2(new_n797), .ZN(new_n798));
  NAND3_X1  g0598(.A1(new_n788), .A2(G190), .A3(G200), .ZN(new_n799));
  INV_X1    g0599(.A(KEYINPUT103), .ZN(new_n800));
  NAND2_X1  g0600(.A1(new_n799), .A2(new_n800), .ZN(new_n801));
  INV_X1    g0601(.A(new_n801), .ZN(new_n802));
  NOR2_X1   g0602(.A1(new_n799), .A2(new_n800), .ZN(new_n803));
  NOR2_X1   g0603(.A1(new_n802), .A2(new_n803), .ZN(new_n804));
  INV_X1    g0604(.A(new_n804), .ZN(new_n805));
  AOI211_X1 g0605(.A(new_n781), .B(new_n798), .C1(G50), .C2(new_n805), .ZN(new_n806));
  AND2_X1   g0606(.A1(new_n805), .A2(G326), .ZN(new_n807));
  INV_X1    g0607(.A(new_n786), .ZN(new_n808));
  AOI22_X1  g0608(.A1(G322), .A2(new_n808), .B1(new_n779), .B2(G329), .ZN(new_n809));
  OAI21_X1  g0609(.A(new_n809), .B1(new_n797), .B2(new_n566), .ZN(new_n810));
  INV_X1    g0610(.A(G283), .ZN(new_n811));
  NOR2_X1   g0611(.A1(new_n783), .A2(new_n811), .ZN(new_n812));
  INV_X1    g0612(.A(new_n790), .ZN(new_n813));
  AOI21_X1  g0613(.A(new_n272), .B1(new_n813), .B2(G294), .ZN(new_n814));
  INV_X1    g0614(.A(G311), .ZN(new_n815));
  XOR2_X1   g0615(.A(KEYINPUT33), .B(G317), .Z(new_n816));
  OAI221_X1 g0616(.A(new_n814), .B1(new_n815), .B2(new_n793), .C1(new_n789), .C2(new_n816), .ZN(new_n817));
  NOR4_X1   g0617(.A1(new_n807), .A2(new_n810), .A3(new_n812), .A4(new_n817), .ZN(new_n818));
  OAI21_X1  g0618(.A(new_n771), .B1(new_n806), .B2(new_n818), .ZN(new_n819));
  INV_X1    g0619(.A(new_n770), .ZN(new_n820));
  OAI21_X1  g0620(.A(new_n819), .B1(new_n699), .B2(new_n820), .ZN(new_n821));
  OAI21_X1  g0621(.A(new_n757), .B1(new_n775), .B2(new_n821), .ZN(G396));
  NAND2_X1  g0622(.A1(new_n271), .A2(new_n678), .ZN(new_n823));
  NAND3_X1  g0623(.A1(new_n297), .A2(new_n300), .A3(new_n823), .ZN(new_n824));
  OAI21_X1  g0624(.A(new_n824), .B1(new_n297), .B2(new_n823), .ZN(new_n825));
  XNOR2_X1  g0625(.A(new_n712), .B(new_n825), .ZN(new_n826));
  INV_X1    g0626(.A(new_n748), .ZN(new_n827));
  AOI21_X1  g0627(.A(KEYINPUT105), .B1(new_n826), .B2(new_n827), .ZN(new_n828));
  NOR2_X1   g0628(.A1(new_n826), .A2(new_n827), .ZN(new_n829));
  NOR2_X1   g0629(.A1(new_n828), .A2(new_n829), .ZN(new_n830));
  NAND3_X1  g0630(.A1(new_n826), .A2(KEYINPUT105), .A3(new_n827), .ZN(new_n831));
  NAND3_X1  g0631(.A1(new_n830), .A2(new_n755), .A3(new_n831), .ZN(new_n832));
  INV_X1    g0632(.A(new_n783), .ZN(new_n833));
  NAND2_X1  g0633(.A1(new_n833), .A2(G87), .ZN(new_n834));
  OAI221_X1 g0634(.A(new_n834), .B1(new_n815), .B2(new_n778), .C1(new_n797), .C2(new_n247), .ZN(new_n835));
  OAI21_X1  g0635(.A(new_n308), .B1(new_n793), .B2(new_n225), .ZN(new_n836));
  OAI22_X1  g0636(.A1(new_n789), .A2(new_n811), .B1(new_n790), .B2(new_n559), .ZN(new_n837));
  NOR3_X1   g0637(.A1(new_n835), .A2(new_n836), .A3(new_n837), .ZN(new_n838));
  INV_X1    g0638(.A(G294), .ZN(new_n839));
  OAI221_X1 g0639(.A(new_n838), .B1(new_n839), .B2(new_n786), .C1(new_n566), .C2(new_n804), .ZN(new_n840));
  OAI22_X1  g0640(.A1(new_n789), .A2(new_n319), .B1(new_n793), .B2(new_n401), .ZN(new_n841));
  AOI21_X1  g0641(.A(new_n841), .B1(new_n805), .B2(G137), .ZN(new_n842));
  INV_X1    g0642(.A(G143), .ZN(new_n843));
  OAI21_X1  g0643(.A(new_n842), .B1(new_n843), .B2(new_n786), .ZN(new_n844));
  XNOR2_X1  g0644(.A(new_n844), .B(KEYINPUT34), .ZN(new_n845));
  INV_X1    g0645(.A(G132), .ZN(new_n846));
  OAI22_X1  g0646(.A1(new_n846), .A2(new_n778), .B1(new_n790), .B2(new_n202), .ZN(new_n847));
  INV_X1    g0647(.A(new_n797), .ZN(new_n848));
  AOI21_X1  g0648(.A(new_n847), .B1(new_n848), .B2(G50), .ZN(new_n849));
  OAI211_X1 g0649(.A(new_n845), .B(new_n849), .C1(new_n203), .C2(new_n783), .ZN(new_n850));
  INV_X1    g0650(.A(new_n760), .ZN(new_n851));
  OAI21_X1  g0651(.A(new_n840), .B1(new_n850), .B2(new_n851), .ZN(new_n852));
  NOR2_X1   g0652(.A1(new_n771), .A2(new_n768), .ZN(new_n853));
  AOI22_X1  g0653(.A1(new_n852), .A2(new_n771), .B1(new_n255), .B2(new_n853), .ZN(new_n854));
  OAI211_X1 g0654(.A(new_n854), .B(new_n758), .C1(new_n769), .C2(new_n825), .ZN(new_n855));
  NAND2_X1  g0655(.A1(new_n832), .A2(new_n855), .ZN(G384));
  NAND2_X1  g0656(.A1(new_n637), .A2(new_n676), .ZN(new_n857));
  OAI211_X1 g0657(.A(new_n683), .B(new_n825), .C1(new_n668), .C2(new_n656), .ZN(new_n858));
  NOR2_X1   g0658(.A1(new_n297), .A2(new_n678), .ZN(new_n859));
  INV_X1    g0659(.A(new_n859), .ZN(new_n860));
  NAND2_X1  g0660(.A1(new_n858), .A2(new_n860), .ZN(new_n861));
  NAND3_X1  g0661(.A1(new_n633), .A2(KEYINPUT80), .A3(KEYINPUT18), .ZN(new_n862));
  NAND3_X1  g0662(.A1(new_n437), .A2(new_n862), .A3(new_n444), .ZN(new_n863));
  OAI21_X1  g0663(.A(new_n390), .B1(new_n397), .B2(new_n203), .ZN(new_n864));
  NAND2_X1  g0664(.A1(new_n864), .A2(new_n399), .ZN(new_n865));
  NAND3_X1  g0665(.A1(new_n865), .A2(new_n267), .A3(new_n398), .ZN(new_n866));
  AOI21_X1  g0666(.A(new_n676), .B1(new_n866), .B2(new_n409), .ZN(new_n867));
  NAND3_X1  g0667(.A1(new_n432), .A2(new_n290), .A3(new_n426), .ZN(new_n868));
  NAND2_X1  g0668(.A1(new_n428), .A2(new_n339), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n868), .A2(new_n869), .ZN(new_n870));
  AOI22_X1  g0670(.A1(new_n866), .A2(new_n409), .B1(new_n870), .B2(new_n676), .ZN(new_n871));
  NOR2_X1   g0671(.A1(new_n410), .A2(new_n429), .ZN(new_n872));
  OAI21_X1  g0672(.A(KEYINPUT37), .B1(new_n871), .B2(new_n872), .ZN(new_n873));
  NAND3_X1  g0673(.A1(new_n434), .A2(new_n407), .A3(new_n409), .ZN(new_n874));
  INV_X1    g0674(.A(new_n676), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n410), .A2(new_n875), .ZN(new_n876));
  INV_X1    g0676(.A(KEYINPUT37), .ZN(new_n877));
  NAND4_X1  g0677(.A1(new_n874), .A2(new_n633), .A3(new_n876), .A4(new_n877), .ZN(new_n878));
  AOI22_X1  g0678(.A1(new_n863), .A2(new_n867), .B1(new_n873), .B2(new_n878), .ZN(new_n879));
  OAI21_X1  g0679(.A(KEYINPUT108), .B1(new_n879), .B2(KEYINPUT38), .ZN(new_n880));
  INV_X1    g0680(.A(KEYINPUT108), .ZN(new_n881));
  INV_X1    g0681(.A(KEYINPUT38), .ZN(new_n882));
  INV_X1    g0682(.A(new_n867), .ZN(new_n883));
  AOI21_X1  g0683(.A(new_n883), .B1(new_n446), .B2(new_n437), .ZN(new_n884));
  AND2_X1   g0684(.A1(new_n873), .A2(new_n878), .ZN(new_n885));
  OAI211_X1 g0685(.A(new_n881), .B(new_n882), .C1(new_n884), .C2(new_n885), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n879), .A2(KEYINPUT38), .ZN(new_n887));
  NAND3_X1  g0687(.A1(new_n880), .A2(new_n886), .A3(new_n887), .ZN(new_n888));
  NOR2_X1   g0688(.A1(new_n626), .A2(new_n683), .ZN(new_n889));
  INV_X1    g0689(.A(new_n889), .ZN(new_n890));
  INV_X1    g0690(.A(KEYINPUT107), .ZN(new_n891));
  INV_X1    g0691(.A(new_n378), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n385), .A2(new_n678), .ZN(new_n893));
  AND4_X1   g0693(.A1(new_n891), .A2(new_n626), .A3(new_n892), .A4(new_n893), .ZN(new_n894));
  AOI21_X1  g0694(.A(new_n891), .B1(new_n386), .B2(new_n893), .ZN(new_n895));
  OAI21_X1  g0695(.A(new_n890), .B1(new_n894), .B2(new_n895), .ZN(new_n896));
  NAND3_X1  g0696(.A1(new_n861), .A2(new_n888), .A3(new_n896), .ZN(new_n897));
  NAND3_X1  g0697(.A1(new_n632), .A2(new_n636), .A3(new_n437), .ZN(new_n898));
  INV_X1    g0698(.A(new_n876), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n898), .A2(new_n899), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n874), .A2(new_n876), .ZN(new_n901));
  NOR3_X1   g0701(.A1(new_n901), .A2(new_n630), .A3(new_n631), .ZN(new_n902));
  OAI21_X1  g0702(.A(new_n878), .B1(new_n902), .B2(new_n877), .ZN(new_n903));
  AOI21_X1  g0703(.A(KEYINPUT38), .B1(new_n900), .B2(new_n903), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n863), .A2(new_n867), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n873), .A2(new_n878), .ZN(new_n906));
  AND3_X1   g0706(.A1(new_n905), .A2(KEYINPUT38), .A3(new_n906), .ZN(new_n907));
  NOR3_X1   g0707(.A1(new_n904), .A2(KEYINPUT39), .A3(new_n907), .ZN(new_n908));
  AOI21_X1  g0708(.A(new_n908), .B1(KEYINPUT39), .B2(new_n888), .ZN(new_n909));
  NOR2_X1   g0709(.A1(new_n626), .A2(new_n678), .ZN(new_n910));
  INV_X1    g0710(.A(new_n910), .ZN(new_n911));
  OAI211_X1 g0711(.A(new_n857), .B(new_n897), .C1(new_n909), .C2(new_n911), .ZN(new_n912));
  NAND4_X1  g0712(.A1(new_n714), .A2(new_n448), .A3(new_n725), .A4(new_n727), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n913), .A2(new_n645), .ZN(new_n914));
  XOR2_X1   g0714(.A(new_n912), .B(new_n914), .Z(new_n915));
  INV_X1    g0715(.A(KEYINPUT40), .ZN(new_n916));
  AND3_X1   g0716(.A1(new_n880), .A2(new_n886), .A3(new_n887), .ZN(new_n917));
  NAND3_X1  g0717(.A1(new_n729), .A2(new_n744), .A3(new_n743), .ZN(new_n918));
  NAND3_X1  g0718(.A1(new_n918), .A2(new_n896), .A3(new_n825), .ZN(new_n919));
  OAI21_X1  g0719(.A(new_n916), .B1(new_n917), .B2(new_n919), .ZN(new_n920));
  AND3_X1   g0720(.A1(new_n918), .A2(new_n896), .A3(new_n825), .ZN(new_n921));
  AND2_X1   g0721(.A1(new_n900), .A2(new_n903), .ZN(new_n922));
  OAI21_X1  g0722(.A(new_n887), .B1(new_n922), .B2(KEYINPUT38), .ZN(new_n923));
  NAND3_X1  g0723(.A1(new_n921), .A2(KEYINPUT40), .A3(new_n923), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n920), .A2(new_n924), .ZN(new_n925));
  AND2_X1   g0725(.A1(new_n448), .A2(new_n918), .ZN(new_n926));
  XNOR2_X1  g0726(.A(new_n925), .B(new_n926), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n927), .A2(G330), .ZN(new_n928));
  XNOR2_X1  g0728(.A(new_n915), .B(new_n928), .ZN(new_n929));
  OAI21_X1  g0729(.A(new_n929), .B1(new_n215), .B2(new_n753), .ZN(new_n930));
  XNOR2_X1  g0730(.A(new_n593), .B(KEYINPUT106), .ZN(new_n931));
  AOI21_X1  g0731(.A(new_n225), .B1(new_n931), .B2(KEYINPUT35), .ZN(new_n932));
  OAI211_X1 g0732(.A(new_n932), .B(new_n213), .C1(KEYINPUT35), .C2(new_n931), .ZN(new_n933));
  XNOR2_X1  g0733(.A(new_n933), .B(KEYINPUT36), .ZN(new_n934));
  OAI21_X1  g0734(.A(G77), .B1(new_n202), .B2(new_n203), .ZN(new_n935));
  OAI22_X1  g0735(.A1(new_n210), .A2(new_n935), .B1(G50), .B2(new_n203), .ZN(new_n936));
  NAND3_X1  g0736(.A1(new_n936), .A2(G1), .A3(new_n672), .ZN(new_n937));
  NAND3_X1  g0737(.A1(new_n930), .A2(new_n934), .A3(new_n937), .ZN(G367));
  INV_X1    g0738(.A(new_n793), .ZN(new_n939));
  AOI22_X1  g0739(.A1(G50), .A2(new_n939), .B1(new_n779), .B2(G137), .ZN(new_n940));
  OAI21_X1  g0740(.A(new_n940), .B1(new_n797), .B2(new_n202), .ZN(new_n941));
  OAI21_X1  g0741(.A(new_n272), .B1(new_n786), .B2(new_n319), .ZN(new_n942));
  NOR2_X1   g0742(.A1(new_n790), .A2(new_n203), .ZN(new_n943));
  INV_X1    g0743(.A(new_n943), .ZN(new_n944));
  OAI21_X1  g0744(.A(new_n944), .B1(new_n401), .B2(new_n789), .ZN(new_n945));
  NOR3_X1   g0745(.A1(new_n941), .A2(new_n942), .A3(new_n945), .ZN(new_n946));
  OAI221_X1 g0746(.A(new_n946), .B1(new_n255), .B2(new_n783), .C1(new_n843), .C2(new_n804), .ZN(new_n947));
  XNOR2_X1  g0747(.A(new_n947), .B(KEYINPUT115), .ZN(new_n948));
  AOI21_X1  g0748(.A(KEYINPUT114), .B1(new_n848), .B2(G116), .ZN(new_n949));
  XNOR2_X1  g0749(.A(new_n949), .B(KEYINPUT46), .ZN(new_n950));
  OAI21_X1  g0750(.A(new_n851), .B1(new_n839), .B2(new_n789), .ZN(new_n951));
  AOI22_X1  g0751(.A1(G97), .A2(new_n833), .B1(new_n779), .B2(G317), .ZN(new_n952));
  OAI221_X1 g0752(.A(new_n952), .B1(new_n811), .B2(new_n793), .C1(new_n566), .C2(new_n786), .ZN(new_n953));
  AOI211_X1 g0753(.A(new_n951), .B(new_n953), .C1(G311), .C2(new_n805), .ZN(new_n954));
  OAI211_X1 g0754(.A(new_n950), .B(new_n954), .C1(new_n247), .C2(new_n790), .ZN(new_n955));
  NAND2_X1  g0755(.A1(new_n948), .A2(new_n955), .ZN(new_n956));
  XNOR2_X1  g0756(.A(new_n956), .B(KEYINPUT47), .ZN(new_n957));
  AOI21_X1  g0757(.A(new_n755), .B1(new_n957), .B2(new_n771), .ZN(new_n958));
  INV_X1    g0758(.A(new_n761), .ZN(new_n959));
  OAI221_X1 g0759(.A(new_n772), .B1(new_n216), .B2(new_n480), .C1(new_n239), .C2(new_n959), .ZN(new_n960));
  NOR2_X1   g0760(.A1(new_n491), .A2(new_n683), .ZN(new_n961));
  XNOR2_X1  g0761(.A(new_n961), .B(KEYINPUT109), .ZN(new_n962));
  OR2_X1    g0762(.A1(new_n962), .A2(new_n657), .ZN(new_n963));
  NAND2_X1  g0763(.A1(new_n962), .A2(new_n715), .ZN(new_n964));
  NAND2_X1  g0764(.A1(new_n963), .A2(new_n964), .ZN(new_n965));
  OAI211_X1 g0765(.A(new_n958), .B(new_n960), .C1(new_n820), .C2(new_n965), .ZN(new_n966));
  NAND2_X1  g0766(.A1(new_n754), .A2(G1), .ZN(new_n967));
  INV_X1    g0767(.A(KEYINPUT44), .ZN(new_n968));
  INV_X1    g0768(.A(new_n622), .ZN(new_n969));
  NAND2_X1  g0769(.A1(new_n604), .A2(new_n678), .ZN(new_n970));
  NAND2_X1  g0770(.A1(new_n969), .A2(new_n970), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n650), .A2(new_n678), .ZN(new_n972));
  NAND2_X1  g0772(.A1(new_n971), .A2(new_n972), .ZN(new_n973));
  OAI21_X1  g0773(.A(new_n968), .B1(new_n694), .B2(new_n973), .ZN(new_n974));
  NOR3_X1   g0774(.A1(new_n682), .A2(KEYINPUT97), .A3(new_n684), .ZN(new_n975));
  AOI21_X1  g0775(.A(new_n689), .B1(new_n688), .B2(new_n690), .ZN(new_n976));
  OAI21_X1  g0776(.A(new_n693), .B1(new_n975), .B2(new_n976), .ZN(new_n977));
  INV_X1    g0777(.A(new_n679), .ZN(new_n978));
  NAND2_X1  g0778(.A1(new_n977), .A2(new_n978), .ZN(new_n979));
  INV_X1    g0779(.A(new_n973), .ZN(new_n980));
  NAND3_X1  g0780(.A1(new_n979), .A2(KEYINPUT44), .A3(new_n980), .ZN(new_n981));
  NAND2_X1  g0781(.A1(new_n974), .A2(new_n981), .ZN(new_n982));
  NAND3_X1  g0782(.A1(new_n977), .A2(new_n978), .A3(new_n973), .ZN(new_n983));
  INV_X1    g0783(.A(KEYINPUT45), .ZN(new_n984));
  NAND2_X1  g0784(.A1(new_n983), .A2(new_n984), .ZN(new_n985));
  NAND3_X1  g0785(.A1(new_n694), .A2(KEYINPUT45), .A3(new_n973), .ZN(new_n986));
  NAND2_X1  g0786(.A1(new_n985), .A2(new_n986), .ZN(new_n987));
  AND3_X1   g0787(.A1(new_n982), .A2(new_n987), .A3(new_n703), .ZN(new_n988));
  AOI21_X1  g0788(.A(new_n703), .B1(new_n982), .B2(new_n987), .ZN(new_n989));
  NOR2_X1   g0789(.A1(new_n988), .A2(new_n989), .ZN(new_n990));
  NOR2_X1   g0790(.A1(new_n692), .A2(new_n693), .ZN(new_n991));
  INV_X1    g0791(.A(new_n693), .ZN(new_n992));
  AOI21_X1  g0792(.A(new_n992), .B1(new_n685), .B2(new_n691), .ZN(new_n993));
  NOR2_X1   g0793(.A1(new_n991), .A2(new_n993), .ZN(new_n994));
  NAND2_X1  g0794(.A1(new_n994), .A2(new_n702), .ZN(new_n995));
  OAI21_X1  g0795(.A(new_n752), .B1(new_n991), .B2(new_n993), .ZN(new_n996));
  NAND2_X1  g0796(.A1(new_n995), .A2(new_n996), .ZN(new_n997));
  NOR2_X1   g0797(.A1(new_n997), .A2(new_n749), .ZN(new_n998));
  AOI21_X1  g0798(.A(KEYINPUT113), .B1(new_n990), .B2(new_n998), .ZN(new_n999));
  AOI21_X1  g0799(.A(KEYINPUT44), .B1(new_n979), .B2(new_n980), .ZN(new_n1000));
  AOI211_X1 g0800(.A(new_n968), .B(new_n973), .C1(new_n977), .C2(new_n978), .ZN(new_n1001));
  AOI21_X1  g0801(.A(KEYINPUT45), .B1(new_n694), .B2(new_n973), .ZN(new_n1002));
  NOR4_X1   g0802(.A1(new_n993), .A2(new_n984), .A3(new_n679), .A4(new_n980), .ZN(new_n1003));
  OAI22_X1  g0803(.A1(new_n1000), .A2(new_n1001), .B1(new_n1002), .B2(new_n1003), .ZN(new_n1004));
  INV_X1    g0804(.A(new_n703), .ZN(new_n1005));
  NAND2_X1  g0805(.A1(new_n1004), .A2(new_n1005), .ZN(new_n1006));
  NAND3_X1  g0806(.A1(new_n982), .A2(new_n987), .A3(new_n703), .ZN(new_n1007));
  NAND4_X1  g0807(.A1(new_n1006), .A2(new_n998), .A3(KEYINPUT113), .A4(new_n1007), .ZN(new_n1008));
  INV_X1    g0808(.A(new_n1008), .ZN(new_n1009));
  OAI21_X1  g0809(.A(new_n750), .B1(new_n999), .B2(new_n1009), .ZN(new_n1010));
  XNOR2_X1  g0810(.A(new_n706), .B(KEYINPUT41), .ZN(new_n1011));
  AOI21_X1  g0811(.A(new_n967), .B1(new_n1010), .B2(new_n1011), .ZN(new_n1012));
  OAI21_X1  g0812(.A(KEYINPUT42), .B1(new_n977), .B2(new_n980), .ZN(new_n1013));
  INV_X1    g0813(.A(KEYINPUT42), .ZN(new_n1014));
  NAND3_X1  g0814(.A1(new_n993), .A2(new_n1014), .A3(new_n973), .ZN(new_n1015));
  OAI21_X1  g0815(.A(new_n617), .B1(new_n971), .B2(new_n537), .ZN(new_n1016));
  XOR2_X1   g0816(.A(new_n1016), .B(KEYINPUT110), .Z(new_n1017));
  OAI211_X1 g0817(.A(new_n1013), .B(new_n1015), .C1(new_n678), .C2(new_n1017), .ZN(new_n1018));
  INV_X1    g0818(.A(new_n965), .ZN(new_n1019));
  INV_X1    g0819(.A(KEYINPUT43), .ZN(new_n1020));
  NAND2_X1  g0820(.A1(new_n1019), .A2(new_n1020), .ZN(new_n1021));
  NAND2_X1  g0821(.A1(new_n1021), .A2(KEYINPUT111), .ZN(new_n1022));
  OAI21_X1  g0822(.A(new_n1022), .B1(new_n1020), .B2(new_n1019), .ZN(new_n1023));
  NAND3_X1  g0823(.A1(new_n965), .A2(KEYINPUT111), .A3(KEYINPUT43), .ZN(new_n1024));
  NAND3_X1  g0824(.A1(new_n1018), .A2(new_n1023), .A3(new_n1024), .ZN(new_n1025));
  AOI21_X1  g0825(.A(new_n1021), .B1(new_n1018), .B2(KEYINPUT111), .ZN(new_n1026));
  NOR2_X1   g0826(.A1(new_n1026), .A2(KEYINPUT112), .ZN(new_n1027));
  INV_X1    g0827(.A(KEYINPUT112), .ZN(new_n1028));
  AOI211_X1 g0828(.A(new_n1028), .B(new_n1021), .C1(new_n1018), .C2(KEYINPUT111), .ZN(new_n1029));
  OAI21_X1  g0829(.A(new_n1025), .B1(new_n1027), .B2(new_n1029), .ZN(new_n1030));
  NOR2_X1   g0830(.A1(new_n703), .A2(new_n980), .ZN(new_n1031));
  XOR2_X1   g0831(.A(new_n1030), .B(new_n1031), .Z(new_n1032));
  OAI21_X1  g0832(.A(new_n966), .B1(new_n1012), .B2(new_n1032), .ZN(G387));
  INV_X1    g0833(.A(new_n789), .ZN(new_n1034));
  AOI22_X1  g0834(.A1(new_n1034), .A2(G311), .B1(new_n939), .B2(G303), .ZN(new_n1035));
  INV_X1    g0835(.A(G317), .ZN(new_n1036));
  INV_X1    g0836(.A(G322), .ZN(new_n1037));
  OAI221_X1 g0837(.A(new_n1035), .B1(new_n1036), .B2(new_n786), .C1(new_n804), .C2(new_n1037), .ZN(new_n1038));
  XNOR2_X1  g0838(.A(new_n1038), .B(KEYINPUT48), .ZN(new_n1039));
  OAI221_X1 g0839(.A(new_n1039), .B1(new_n811), .B2(new_n790), .C1(new_n839), .C2(new_n797), .ZN(new_n1040));
  INV_X1    g0840(.A(KEYINPUT49), .ZN(new_n1041));
  OR2_X1    g0841(.A1(new_n1040), .A2(new_n1041), .ZN(new_n1042));
  NAND2_X1  g0842(.A1(new_n779), .A2(G326), .ZN(new_n1043));
  NAND2_X1  g0843(.A1(new_n1040), .A2(new_n1041), .ZN(new_n1044));
  AOI21_X1  g0844(.A(new_n760), .B1(G116), .B2(new_n833), .ZN(new_n1045));
  NAND4_X1  g0845(.A1(new_n1042), .A2(new_n1043), .A3(new_n1044), .A4(new_n1045), .ZN(new_n1046));
  AOI22_X1  g0846(.A1(G97), .A2(new_n833), .B1(new_n779), .B2(G150), .ZN(new_n1047));
  OAI221_X1 g0847(.A(new_n1047), .B1(new_n203), .B2(new_n793), .C1(new_n797), .C2(new_n255), .ZN(new_n1048));
  OAI221_X1 g0848(.A(new_n760), .B1(new_n261), .B2(new_n789), .C1(new_n480), .C2(new_n790), .ZN(new_n1049));
  NOR2_X1   g0849(.A1(new_n1048), .A2(new_n1049), .ZN(new_n1050));
  OAI221_X1 g0850(.A(new_n1050), .B1(new_n322), .B2(new_n786), .C1(new_n401), .C2(new_n804), .ZN(new_n1051));
  NAND2_X1  g0851(.A1(new_n1046), .A2(new_n1051), .ZN(new_n1052));
  NAND2_X1  g0852(.A1(new_n262), .A2(new_n322), .ZN(new_n1053));
  AOI211_X1 g0853(.A(G116), .B(new_n475), .C1(new_n1053), .C2(KEYINPUT50), .ZN(new_n1054));
  NAND2_X1  g0854(.A1(G68), .A2(G77), .ZN(new_n1055));
  OR2_X1    g0855(.A1(new_n1053), .A2(KEYINPUT50), .ZN(new_n1056));
  NAND4_X1  g0856(.A1(new_n1054), .A2(new_n458), .A3(new_n1055), .A4(new_n1056), .ZN(new_n1057));
  AOI21_X1  g0857(.A(new_n959), .B1(new_n236), .B2(G45), .ZN(new_n1058));
  NOR3_X1   g0858(.A1(new_n708), .A2(new_n705), .A3(new_n308), .ZN(new_n1059));
  OAI21_X1  g0859(.A(new_n1057), .B1(new_n1058), .B2(new_n1059), .ZN(new_n1060));
  OAI21_X1  g0860(.A(new_n1060), .B1(G107), .B2(new_n216), .ZN(new_n1061));
  AOI22_X1  g0861(.A1(new_n1052), .A2(new_n771), .B1(new_n772), .B2(new_n1061), .ZN(new_n1062));
  OAI211_X1 g0862(.A(new_n1062), .B(new_n758), .C1(new_n692), .C2(new_n820), .ZN(new_n1063));
  INV_X1    g0863(.A(new_n967), .ZN(new_n1064));
  INV_X1    g0864(.A(new_n997), .ZN(new_n1065));
  OAI21_X1  g0865(.A(new_n706), .B1(new_n1065), .B2(new_n750), .ZN(new_n1066));
  OAI221_X1 g0866(.A(new_n1063), .B1(new_n1064), .B2(new_n997), .C1(new_n1066), .C2(new_n998), .ZN(G393));
  NOR3_X1   g0867(.A1(new_n988), .A2(new_n989), .A3(new_n1064), .ZN(new_n1068));
  NAND2_X1  g0868(.A1(new_n249), .A2(new_n761), .ZN(new_n1069));
  OAI211_X1 g0869(.A(new_n1069), .B(new_n772), .C1(new_n559), .C2(new_n216), .ZN(new_n1070));
  XOR2_X1   g0870(.A(new_n1070), .B(KEYINPUT116), .Z(new_n1071));
  OAI221_X1 g0871(.A(new_n760), .B1(new_n322), .B2(new_n789), .C1(new_n255), .C2(new_n790), .ZN(new_n1072));
  OAI221_X1 g0872(.A(new_n834), .B1(new_n261), .B2(new_n793), .C1(new_n797), .C2(new_n203), .ZN(new_n1073));
  INV_X1    g0873(.A(KEYINPUT51), .ZN(new_n1074));
  OAI22_X1  g0874(.A1(new_n804), .A2(new_n319), .B1(new_n401), .B2(new_n786), .ZN(new_n1075));
  AOI211_X1 g0875(.A(new_n1072), .B(new_n1073), .C1(new_n1074), .C2(new_n1075), .ZN(new_n1076));
  OAI221_X1 g0876(.A(new_n1076), .B1(new_n1074), .B2(new_n1075), .C1(new_n843), .C2(new_n778), .ZN(new_n1077));
  OAI22_X1  g0877(.A1(new_n804), .A2(new_n1036), .B1(new_n815), .B2(new_n786), .ZN(new_n1078));
  XNOR2_X1  g0878(.A(new_n1078), .B(KEYINPUT52), .ZN(new_n1079));
  OAI22_X1  g0879(.A1(new_n789), .A2(new_n566), .B1(new_n790), .B2(new_n225), .ZN(new_n1080));
  OAI221_X1 g0880(.A(new_n308), .B1(new_n783), .B2(new_n247), .C1(new_n839), .C2(new_n793), .ZN(new_n1081));
  AOI211_X1 g0881(.A(new_n1080), .B(new_n1081), .C1(new_n848), .C2(G283), .ZN(new_n1082));
  OAI211_X1 g0882(.A(new_n1079), .B(new_n1082), .C1(new_n1037), .C2(new_n778), .ZN(new_n1083));
  NAND2_X1  g0883(.A1(new_n1077), .A2(new_n1083), .ZN(new_n1084));
  AOI21_X1  g0884(.A(new_n755), .B1(new_n1084), .B2(new_n771), .ZN(new_n1085));
  OAI211_X1 g0885(.A(new_n1071), .B(new_n1085), .C1(new_n820), .C2(new_n973), .ZN(new_n1086));
  INV_X1    g0886(.A(new_n1086), .ZN(new_n1087));
  NAND3_X1  g0887(.A1(new_n1006), .A2(new_n998), .A3(new_n1007), .ZN(new_n1088));
  INV_X1    g0888(.A(KEYINPUT113), .ZN(new_n1089));
  NAND2_X1  g0889(.A1(new_n1088), .A2(new_n1089), .ZN(new_n1090));
  AOI21_X1  g0890(.A(new_n707), .B1(new_n1090), .B2(new_n1008), .ZN(new_n1091));
  OR2_X1    g0891(.A1(new_n990), .A2(new_n998), .ZN(new_n1092));
  AOI211_X1 g0892(.A(new_n1068), .B(new_n1087), .C1(new_n1091), .C2(new_n1092), .ZN(new_n1093));
  INV_X1    g0893(.A(new_n1093), .ZN(G390));
  INV_X1    g0894(.A(KEYINPUT117), .ZN(new_n1095));
  NAND2_X1  g0895(.A1(new_n386), .A2(new_n893), .ZN(new_n1096));
  NAND2_X1  g0896(.A1(new_n1096), .A2(KEYINPUT107), .ZN(new_n1097));
  NAND3_X1  g0897(.A1(new_n386), .A2(new_n891), .A3(new_n893), .ZN(new_n1098));
  AOI21_X1  g0898(.A(new_n889), .B1(new_n1097), .B2(new_n1098), .ZN(new_n1099));
  NAND3_X1  g0899(.A1(new_n723), .A2(new_n683), .A3(new_n825), .ZN(new_n1100));
  AOI21_X1  g0900(.A(new_n1099), .B1(new_n1100), .B2(new_n860), .ZN(new_n1101));
  OAI21_X1  g0901(.A(new_n911), .B1(new_n904), .B2(new_n907), .ZN(new_n1102));
  OR2_X1    g0902(.A1(new_n1101), .A2(new_n1102), .ZN(new_n1103));
  AND2_X1   g0903(.A1(new_n825), .A2(G330), .ZN(new_n1104));
  NAND3_X1  g0904(.A1(new_n747), .A2(new_n896), .A3(new_n1104), .ZN(new_n1105));
  INV_X1    g0905(.A(new_n1105), .ZN(new_n1106));
  AOI21_X1  g0906(.A(new_n910), .B1(new_n861), .B2(new_n896), .ZN(new_n1107));
  NAND2_X1  g0907(.A1(new_n888), .A2(KEYINPUT39), .ZN(new_n1108));
  INV_X1    g0908(.A(KEYINPUT39), .ZN(new_n1109));
  OAI211_X1 g0909(.A(new_n1109), .B(new_n887), .C1(new_n922), .C2(KEYINPUT38), .ZN(new_n1110));
  NAND2_X1  g0910(.A1(new_n1108), .A2(new_n1110), .ZN(new_n1111));
  OAI211_X1 g0911(.A(new_n1103), .B(new_n1106), .C1(new_n1107), .C2(new_n1111), .ZN(new_n1112));
  NOR2_X1   g0912(.A1(new_n1101), .A2(new_n1102), .ZN(new_n1113));
  AND3_X1   g0913(.A1(new_n662), .A2(new_n537), .A3(new_n663), .ZN(new_n1114));
  NAND4_X1  g0914(.A1(new_n969), .A2(new_n548), .A3(new_n647), .A4(new_n649), .ZN(new_n1115));
  OAI21_X1  g0915(.A(KEYINPUT93), .B1(new_n1114), .B2(new_n1115), .ZN(new_n1116));
  NAND3_X1  g0916(.A1(new_n660), .A2(new_n664), .A3(new_n665), .ZN(new_n1117));
  NAND2_X1  g0917(.A1(new_n1116), .A2(new_n1117), .ZN(new_n1118));
  NAND3_X1  g0918(.A1(new_n720), .A2(new_n721), .A3(new_n650), .ZN(new_n1119));
  AOI21_X1  g0919(.A(new_n653), .B1(new_n1119), .B2(KEYINPUT26), .ZN(new_n1120));
  AOI21_X1  g0920(.A(new_n678), .B1(new_n1118), .B2(new_n1120), .ZN(new_n1121));
  AOI21_X1  g0921(.A(new_n859), .B1(new_n1121), .B2(new_n825), .ZN(new_n1122));
  OAI21_X1  g0922(.A(new_n911), .B1(new_n1122), .B2(new_n1099), .ZN(new_n1123));
  AOI21_X1  g0923(.A(new_n1113), .B1(new_n1123), .B2(new_n909), .ZN(new_n1124));
  AND3_X1   g0924(.A1(new_n918), .A2(new_n896), .A3(new_n1104), .ZN(new_n1125));
  OAI21_X1  g0925(.A(new_n1112), .B1(new_n1124), .B2(new_n1125), .ZN(new_n1126));
  AOI21_X1  g0926(.A(new_n896), .B1(new_n747), .B2(new_n1104), .ZN(new_n1127));
  OAI21_X1  g0927(.A(new_n861), .B1(new_n1125), .B2(new_n1127), .ZN(new_n1128));
  NAND2_X1  g0928(.A1(new_n918), .A2(new_n1104), .ZN(new_n1129));
  NAND2_X1  g0929(.A1(new_n1129), .A2(new_n1099), .ZN(new_n1130));
  AND2_X1   g0930(.A1(new_n1100), .A2(new_n860), .ZN(new_n1131));
  NAND3_X1  g0931(.A1(new_n1130), .A2(new_n1131), .A3(new_n1105), .ZN(new_n1132));
  AND2_X1   g0932(.A1(new_n1128), .A2(new_n1132), .ZN(new_n1133));
  NAND3_X1  g0933(.A1(new_n448), .A2(G330), .A3(new_n918), .ZN(new_n1134));
  NAND3_X1  g0934(.A1(new_n913), .A2(new_n645), .A3(new_n1134), .ZN(new_n1135));
  NOR2_X1   g0935(.A1(new_n1133), .A2(new_n1135), .ZN(new_n1136));
  OAI21_X1  g0936(.A(new_n1095), .B1(new_n1126), .B2(new_n1136), .ZN(new_n1137));
  AOI21_X1  g0937(.A(new_n707), .B1(new_n1126), .B2(new_n1136), .ZN(new_n1138));
  OAI21_X1  g0938(.A(new_n1103), .B1(new_n1107), .B2(new_n1111), .ZN(new_n1139));
  INV_X1    g0939(.A(new_n1125), .ZN(new_n1140));
  NAND2_X1  g0940(.A1(new_n1139), .A2(new_n1140), .ZN(new_n1141));
  NAND2_X1  g0941(.A1(new_n1128), .A2(new_n1132), .ZN(new_n1142));
  NAND4_X1  g0942(.A1(new_n1142), .A2(new_n645), .A3(new_n913), .A4(new_n1134), .ZN(new_n1143));
  NAND4_X1  g0943(.A1(new_n1141), .A2(new_n1143), .A3(KEYINPUT117), .A4(new_n1112), .ZN(new_n1144));
  NAND3_X1  g0944(.A1(new_n1137), .A2(new_n1138), .A3(new_n1144), .ZN(new_n1145));
  NOR2_X1   g0945(.A1(new_n797), .A2(new_n319), .ZN(new_n1146));
  XNOR2_X1  g0946(.A(KEYINPUT118), .B(KEYINPUT53), .ZN(new_n1147));
  XNOR2_X1  g0947(.A(new_n1146), .B(new_n1147), .ZN(new_n1148));
  NAND2_X1  g0948(.A1(new_n808), .A2(G132), .ZN(new_n1149));
  NAND2_X1  g0949(.A1(new_n805), .A2(G128), .ZN(new_n1150));
  INV_X1    g0950(.A(G125), .ZN(new_n1151));
  OAI22_X1  g0951(.A1(new_n783), .A2(new_n322), .B1(new_n778), .B2(new_n1151), .ZN(new_n1152));
  INV_X1    g0952(.A(G137), .ZN(new_n1153));
  OAI221_X1 g0953(.A(new_n272), .B1(new_n790), .B2(new_n401), .C1(new_n789), .C2(new_n1153), .ZN(new_n1154));
  XOR2_X1   g0954(.A(KEYINPUT54), .B(G143), .Z(new_n1155));
  AOI211_X1 g0955(.A(new_n1152), .B(new_n1154), .C1(new_n939), .C2(new_n1155), .ZN(new_n1156));
  NAND4_X1  g0956(.A1(new_n1148), .A2(new_n1149), .A3(new_n1150), .A4(new_n1156), .ZN(new_n1157));
  AOI22_X1  g0957(.A1(new_n805), .A2(G283), .B1(G107), .B2(new_n1034), .ZN(new_n1158));
  OAI21_X1  g0958(.A(new_n1158), .B1(new_n559), .B2(new_n793), .ZN(new_n1159));
  OR2_X1    g0959(.A1(new_n1159), .A2(KEYINPUT119), .ZN(new_n1160));
  NAND2_X1  g0960(.A1(new_n1159), .A2(KEYINPUT119), .ZN(new_n1161));
  OAI22_X1  g0961(.A1(new_n783), .A2(new_n203), .B1(new_n778), .B2(new_n839), .ZN(new_n1162));
  OAI21_X1  g0962(.A(new_n308), .B1(new_n1162), .B2(KEYINPUT120), .ZN(new_n1163));
  NOR2_X1   g0963(.A1(new_n797), .A2(new_n474), .ZN(new_n1164));
  AOI211_X1 g0964(.A(new_n1163), .B(new_n1164), .C1(KEYINPUT120), .C2(new_n1162), .ZN(new_n1165));
  NAND3_X1  g0965(.A1(new_n1160), .A2(new_n1161), .A3(new_n1165), .ZN(new_n1166));
  OAI22_X1  g0966(.A1(new_n786), .A2(new_n225), .B1(new_n790), .B2(new_n255), .ZN(new_n1167));
  XNOR2_X1  g0967(.A(new_n1167), .B(KEYINPUT121), .ZN(new_n1168));
  OAI21_X1  g0968(.A(new_n1157), .B1(new_n1166), .B2(new_n1168), .ZN(new_n1169));
  NAND2_X1  g0969(.A1(new_n1169), .A2(new_n771), .ZN(new_n1170));
  INV_X1    g0970(.A(new_n853), .ZN(new_n1171));
  OAI21_X1  g0971(.A(new_n1170), .B1(new_n262), .B2(new_n1171), .ZN(new_n1172));
  AOI211_X1 g0972(.A(new_n755), .B(new_n1172), .C1(new_n909), .C2(new_n768), .ZN(new_n1173));
  AOI21_X1  g0973(.A(new_n1173), .B1(new_n1126), .B2(new_n967), .ZN(new_n1174));
  NAND2_X1  g0974(.A1(new_n1145), .A2(new_n1174), .ZN(G378));
  NAND2_X1  g0975(.A1(new_n325), .A2(new_n875), .ZN(new_n1176));
  NAND3_X1  g0976(.A1(new_n643), .A2(new_n341), .A3(new_n1176), .ZN(new_n1177));
  INV_X1    g0977(.A(KEYINPUT55), .ZN(new_n1178));
  NAND3_X1  g0978(.A1(new_n332), .A2(new_n338), .A3(new_n341), .ZN(new_n1179));
  NAND3_X1  g0979(.A1(new_n1179), .A2(new_n325), .A3(new_n875), .ZN(new_n1180));
  AND3_X1   g0980(.A1(new_n1177), .A2(new_n1178), .A3(new_n1180), .ZN(new_n1181));
  AOI21_X1  g0981(.A(new_n1178), .B1(new_n1177), .B2(new_n1180), .ZN(new_n1182));
  INV_X1    g0982(.A(KEYINPUT56), .ZN(new_n1183));
  OR3_X1    g0983(.A1(new_n1181), .A2(new_n1182), .A3(new_n1183), .ZN(new_n1184));
  OAI21_X1  g0984(.A(new_n1183), .B1(new_n1181), .B2(new_n1182), .ZN(new_n1185));
  NAND2_X1  g0985(.A1(new_n1184), .A2(new_n1185), .ZN(new_n1186));
  INV_X1    g0986(.A(new_n1186), .ZN(new_n1187));
  NAND2_X1  g0987(.A1(new_n1187), .A2(new_n768), .ZN(new_n1188));
  NAND2_X1  g0988(.A1(new_n853), .A2(new_n322), .ZN(new_n1189));
  NAND2_X1  g0989(.A1(new_n833), .A2(G58), .ZN(new_n1190));
  OAI211_X1 g0990(.A(new_n1190), .B(new_n520), .C1(new_n811), .C2(new_n778), .ZN(new_n1191));
  AOI211_X1 g0991(.A(new_n760), .B(new_n1191), .C1(new_n848), .C2(G77), .ZN(new_n1192));
  XNOR2_X1  g0992(.A(new_n1192), .B(KEYINPUT122), .ZN(new_n1193));
  OAI221_X1 g0993(.A(new_n944), .B1(new_n559), .B2(new_n789), .C1(new_n480), .C2(new_n793), .ZN(new_n1194));
  AOI21_X1  g0994(.A(new_n1194), .B1(G116), .B2(new_n805), .ZN(new_n1195));
  OAI211_X1 g0995(.A(new_n1193), .B(new_n1195), .C1(new_n247), .C2(new_n786), .ZN(new_n1196));
  XNOR2_X1  g0996(.A(new_n1196), .B(KEYINPUT58), .ZN(new_n1197));
  AOI21_X1  g0997(.A(G41), .B1(new_n760), .B2(G33), .ZN(new_n1198));
  AOI22_X1  g0998(.A1(new_n808), .A2(G128), .B1(new_n813), .B2(G150), .ZN(new_n1199));
  OAI21_X1  g0999(.A(new_n1199), .B1(new_n846), .B2(new_n789), .ZN(new_n1200));
  AOI21_X1  g1000(.A(new_n1200), .B1(new_n848), .B2(new_n1155), .ZN(new_n1201));
  OAI221_X1 g1001(.A(new_n1201), .B1(new_n1151), .B2(new_n804), .C1(new_n1153), .C2(new_n793), .ZN(new_n1202));
  XNOR2_X1  g1002(.A(new_n1202), .B(KEYINPUT59), .ZN(new_n1203));
  AOI21_X1  g1003(.A(G41), .B1(new_n779), .B2(G124), .ZN(new_n1204));
  OAI211_X1 g1004(.A(new_n1204), .B(new_n304), .C1(new_n401), .C2(new_n783), .ZN(new_n1205));
  XOR2_X1   g1005(.A(new_n1205), .B(KEYINPUT123), .Z(new_n1206));
  OAI221_X1 g1006(.A(new_n1197), .B1(G50), .B2(new_n1198), .C1(new_n1203), .C2(new_n1206), .ZN(new_n1207));
  AOI21_X1  g1007(.A(new_n755), .B1(new_n1207), .B2(new_n771), .ZN(new_n1208));
  NAND3_X1  g1008(.A1(new_n1188), .A2(new_n1189), .A3(new_n1208), .ZN(new_n1209));
  INV_X1    g1009(.A(new_n1209), .ZN(new_n1210));
  AND3_X1   g1010(.A1(new_n920), .A2(new_n924), .A3(G330), .ZN(new_n1211));
  NOR2_X1   g1011(.A1(new_n912), .A2(new_n1211), .ZN(new_n1212));
  NAND3_X1  g1012(.A1(new_n920), .A2(new_n924), .A3(G330), .ZN(new_n1213));
  AOI21_X1  g1013(.A(new_n1099), .B1(new_n858), .B2(new_n860), .ZN(new_n1214));
  AOI22_X1  g1014(.A1(new_n1111), .A2(new_n910), .B1(new_n1214), .B2(new_n888), .ZN(new_n1215));
  AOI21_X1  g1015(.A(new_n1213), .B1(new_n1215), .B2(new_n857), .ZN(new_n1216));
  OAI21_X1  g1016(.A(new_n1186), .B1(new_n1212), .B2(new_n1216), .ZN(new_n1217));
  NAND2_X1  g1017(.A1(new_n912), .A2(new_n1211), .ZN(new_n1218));
  NAND3_X1  g1018(.A1(new_n1215), .A2(new_n1213), .A3(new_n857), .ZN(new_n1219));
  NAND3_X1  g1019(.A1(new_n1218), .A2(new_n1219), .A3(new_n1187), .ZN(new_n1220));
  NAND2_X1  g1020(.A1(new_n1217), .A2(new_n1220), .ZN(new_n1221));
  AOI21_X1  g1021(.A(new_n1210), .B1(new_n1221), .B2(new_n967), .ZN(new_n1222));
  INV_X1    g1022(.A(new_n1112), .ZN(new_n1223));
  OAI211_X1 g1023(.A(new_n1108), .B(new_n1110), .C1(new_n1214), .C2(new_n910), .ZN(new_n1224));
  AOI21_X1  g1024(.A(new_n1125), .B1(new_n1224), .B2(new_n1103), .ZN(new_n1225));
  OAI21_X1  g1025(.A(new_n1136), .B1(new_n1223), .B2(new_n1225), .ZN(new_n1226));
  INV_X1    g1026(.A(new_n1135), .ZN(new_n1227));
  AOI22_X1  g1027(.A1(new_n1217), .A2(new_n1220), .B1(new_n1226), .B2(new_n1227), .ZN(new_n1228));
  OAI21_X1  g1028(.A(new_n706), .B1(new_n1228), .B2(KEYINPUT57), .ZN(new_n1229));
  AND3_X1   g1029(.A1(new_n1218), .A2(new_n1219), .A3(new_n1187), .ZN(new_n1230));
  AOI21_X1  g1030(.A(new_n1187), .B1(new_n1218), .B2(new_n1219), .ZN(new_n1231));
  AOI21_X1  g1031(.A(new_n1143), .B1(new_n1141), .B2(new_n1112), .ZN(new_n1232));
  OAI22_X1  g1032(.A1(new_n1230), .A2(new_n1231), .B1(new_n1232), .B2(new_n1135), .ZN(new_n1233));
  INV_X1    g1033(.A(KEYINPUT57), .ZN(new_n1234));
  NOR2_X1   g1034(.A1(new_n1233), .A2(new_n1234), .ZN(new_n1235));
  OAI21_X1  g1035(.A(new_n1222), .B1(new_n1229), .B2(new_n1235), .ZN(G375));
  NAND2_X1  g1036(.A1(new_n779), .A2(G128), .ZN(new_n1237));
  OAI211_X1 g1037(.A(new_n1190), .B(new_n1237), .C1(new_n1153), .C2(new_n786), .ZN(new_n1238));
  AOI21_X1  g1038(.A(new_n851), .B1(new_n1034), .B2(new_n1155), .ZN(new_n1239));
  OAI21_X1  g1039(.A(new_n1239), .B1(new_n322), .B2(new_n790), .ZN(new_n1240));
  AOI211_X1 g1040(.A(new_n1238), .B(new_n1240), .C1(G159), .C2(new_n848), .ZN(new_n1241));
  OAI221_X1 g1041(.A(new_n1241), .B1(new_n846), .B2(new_n804), .C1(new_n319), .C2(new_n793), .ZN(new_n1242));
  NOR2_X1   g1042(.A1(new_n797), .A2(new_n559), .ZN(new_n1243));
  OAI21_X1  g1043(.A(new_n308), .B1(new_n789), .B2(new_n225), .ZN(new_n1244));
  OAI22_X1  g1044(.A1(new_n480), .A2(new_n790), .B1(new_n255), .B2(new_n783), .ZN(new_n1245));
  OAI22_X1  g1045(.A1(new_n793), .A2(new_n247), .B1(new_n778), .B2(new_n566), .ZN(new_n1246));
  NOR4_X1   g1046(.A1(new_n1243), .A2(new_n1244), .A3(new_n1245), .A4(new_n1246), .ZN(new_n1247));
  OAI221_X1 g1047(.A(new_n1247), .B1(new_n811), .B2(new_n786), .C1(new_n839), .C2(new_n804), .ZN(new_n1248));
  NAND2_X1  g1048(.A1(new_n1242), .A2(new_n1248), .ZN(new_n1249));
  NAND2_X1  g1049(.A1(new_n1249), .A2(new_n771), .ZN(new_n1250));
  OAI21_X1  g1050(.A(new_n1250), .B1(G68), .B2(new_n1171), .ZN(new_n1251));
  AOI211_X1 g1051(.A(new_n755), .B(new_n1251), .C1(new_n1099), .C2(new_n768), .ZN(new_n1252));
  AOI21_X1  g1052(.A(new_n1252), .B1(new_n1142), .B2(new_n967), .ZN(new_n1253));
  OAI21_X1  g1053(.A(new_n1011), .B1(new_n1227), .B2(new_n1142), .ZN(new_n1254));
  OAI21_X1  g1054(.A(new_n1253), .B1(new_n1254), .B2(new_n1136), .ZN(new_n1255));
  XOR2_X1   g1055(.A(new_n1255), .B(KEYINPUT124), .Z(G381));
  INV_X1    g1056(.A(KEYINPUT125), .ZN(new_n1257));
  NAND3_X1  g1057(.A1(new_n1145), .A2(new_n1257), .A3(new_n1174), .ZN(new_n1258));
  INV_X1    g1058(.A(new_n1258), .ZN(new_n1259));
  AOI21_X1  g1059(.A(new_n1257), .B1(new_n1145), .B2(new_n1174), .ZN(new_n1260));
  NOR2_X1   g1060(.A1(new_n1259), .A2(new_n1260), .ZN(new_n1261));
  NOR2_X1   g1061(.A1(new_n1261), .A2(G375), .ZN(new_n1262));
  XNOR2_X1  g1062(.A(new_n1030), .B(new_n1031), .ZN(new_n1263));
  INV_X1    g1063(.A(new_n1011), .ZN(new_n1264));
  NAND2_X1  g1064(.A1(new_n1090), .A2(new_n1008), .ZN(new_n1265));
  AOI21_X1  g1065(.A(new_n1264), .B1(new_n1265), .B2(new_n750), .ZN(new_n1266));
  OAI21_X1  g1066(.A(new_n1263), .B1(new_n1266), .B2(new_n967), .ZN(new_n1267));
  AND3_X1   g1067(.A1(new_n1267), .A2(new_n1093), .A3(new_n966), .ZN(new_n1268));
  NOR4_X1   g1068(.A1(G381), .A2(G396), .A3(G384), .A4(G393), .ZN(new_n1269));
  NAND3_X1  g1069(.A1(new_n1262), .A2(new_n1268), .A3(new_n1269), .ZN(G407));
  NAND2_X1  g1070(.A1(new_n1262), .A2(new_n677), .ZN(new_n1271));
  NAND3_X1  g1071(.A1(G407), .A2(G213), .A3(new_n1271), .ZN(G409));
  OAI21_X1  g1072(.A(new_n1222), .B1(new_n1264), .B2(new_n1233), .ZN(new_n1273));
  OAI21_X1  g1073(.A(new_n1273), .B1(new_n1259), .B2(new_n1260), .ZN(new_n1274));
  OAI211_X1 g1074(.A(G378), .B(new_n1222), .C1(new_n1229), .C2(new_n1235), .ZN(new_n1275));
  AOI22_X1  g1075(.A1(new_n1274), .A2(new_n1275), .B1(G213), .B2(new_n677), .ZN(new_n1276));
  NAND3_X1  g1076(.A1(new_n1133), .A2(KEYINPUT60), .A3(new_n1135), .ZN(new_n1277));
  INV_X1    g1077(.A(KEYINPUT126), .ZN(new_n1278));
  XNOR2_X1  g1078(.A(new_n1277), .B(new_n1278), .ZN(new_n1279));
  NOR2_X1   g1079(.A1(new_n1227), .A2(new_n1142), .ZN(new_n1280));
  OAI211_X1 g1080(.A(new_n706), .B(new_n1143), .C1(new_n1280), .C2(KEYINPUT60), .ZN(new_n1281));
  OAI21_X1  g1081(.A(new_n1253), .B1(new_n1279), .B2(new_n1281), .ZN(new_n1282));
  NAND3_X1  g1082(.A1(new_n1282), .A2(new_n855), .A3(new_n832), .ZN(new_n1283));
  OAI211_X1 g1083(.A(G384), .B(new_n1253), .C1(new_n1279), .C2(new_n1281), .ZN(new_n1284));
  NAND2_X1  g1084(.A1(new_n1283), .A2(new_n1284), .ZN(new_n1285));
  NAND2_X1  g1085(.A1(new_n677), .A2(G213), .ZN(new_n1286));
  INV_X1    g1086(.A(G2897), .ZN(new_n1287));
  NOR2_X1   g1087(.A1(new_n1286), .A2(new_n1287), .ZN(new_n1288));
  NAND2_X1  g1088(.A1(new_n1285), .A2(new_n1288), .ZN(new_n1289));
  OAI211_X1 g1089(.A(new_n1283), .B(new_n1284), .C1(new_n1287), .C2(new_n1286), .ZN(new_n1290));
  NAND2_X1  g1090(.A1(new_n1289), .A2(new_n1290), .ZN(new_n1291));
  OR2_X1    g1091(.A1(new_n1276), .A2(new_n1291), .ZN(new_n1292));
  NAND2_X1  g1092(.A1(new_n1274), .A2(new_n1275), .ZN(new_n1293));
  INV_X1    g1093(.A(new_n1285), .ZN(new_n1294));
  NAND3_X1  g1094(.A1(new_n1293), .A2(new_n1286), .A3(new_n1294), .ZN(new_n1295));
  NAND2_X1  g1095(.A1(new_n1295), .A2(KEYINPUT62), .ZN(new_n1296));
  INV_X1    g1096(.A(KEYINPUT61), .ZN(new_n1297));
  INV_X1    g1097(.A(KEYINPUT62), .ZN(new_n1298));
  NAND3_X1  g1098(.A1(new_n1276), .A2(new_n1298), .A3(new_n1294), .ZN(new_n1299));
  NAND4_X1  g1099(.A1(new_n1292), .A2(new_n1296), .A3(new_n1297), .A4(new_n1299), .ZN(new_n1300));
  XOR2_X1   g1100(.A(G393), .B(G396), .Z(new_n1301));
  AOI21_X1  g1101(.A(new_n1093), .B1(new_n1267), .B2(new_n966), .ZN(new_n1302));
  OAI21_X1  g1102(.A(new_n1301), .B1(new_n1268), .B2(new_n1302), .ZN(new_n1303));
  NAND2_X1  g1103(.A1(G387), .A2(G390), .ZN(new_n1304));
  NAND3_X1  g1104(.A1(new_n1267), .A2(new_n1093), .A3(new_n966), .ZN(new_n1305));
  INV_X1    g1105(.A(new_n1301), .ZN(new_n1306));
  NAND3_X1  g1106(.A1(new_n1304), .A2(new_n1305), .A3(new_n1306), .ZN(new_n1307));
  NAND2_X1  g1107(.A1(new_n1303), .A2(new_n1307), .ZN(new_n1308));
  NAND2_X1  g1108(.A1(new_n1300), .A2(new_n1308), .ZN(new_n1309));
  AND3_X1   g1109(.A1(new_n1276), .A2(KEYINPUT63), .A3(new_n1294), .ZN(new_n1310));
  NOR2_X1   g1110(.A1(new_n1310), .A2(new_n1308), .ZN(new_n1311));
  OAI21_X1  g1111(.A(KEYINPUT63), .B1(new_n1276), .B2(new_n1291), .ZN(new_n1312));
  AOI21_X1  g1112(.A(KEYINPUT61), .B1(new_n1312), .B2(new_n1295), .ZN(new_n1313));
  NAND2_X1  g1113(.A1(new_n1311), .A2(new_n1313), .ZN(new_n1314));
  NAND2_X1  g1114(.A1(new_n1309), .A2(new_n1314), .ZN(G405));
  OAI21_X1  g1115(.A(new_n967), .B1(new_n1230), .B2(new_n1231), .ZN(new_n1316));
  NAND2_X1  g1116(.A1(new_n1316), .A2(new_n1209), .ZN(new_n1317));
  AOI21_X1  g1117(.A(new_n707), .B1(new_n1233), .B2(new_n1234), .ZN(new_n1318));
  NAND2_X1  g1118(.A1(new_n1228), .A2(KEYINPUT57), .ZN(new_n1319));
  AOI21_X1  g1119(.A(new_n1317), .B1(new_n1318), .B2(new_n1319), .ZN(new_n1320));
  OAI211_X1 g1120(.A(new_n1275), .B(new_n1285), .C1(new_n1261), .C2(new_n1320), .ZN(new_n1321));
  INV_X1    g1121(.A(new_n1321), .ZN(new_n1322));
  NAND2_X1  g1122(.A1(G378), .A2(KEYINPUT125), .ZN(new_n1323));
  NAND2_X1  g1123(.A1(new_n1323), .A2(new_n1258), .ZN(new_n1324));
  NAND2_X1  g1124(.A1(G375), .A2(new_n1324), .ZN(new_n1325));
  AOI21_X1  g1125(.A(new_n1285), .B1(new_n1325), .B2(new_n1275), .ZN(new_n1326));
  NOR2_X1   g1126(.A1(new_n1322), .A2(new_n1326), .ZN(new_n1327));
  INV_X1    g1127(.A(KEYINPUT127), .ZN(new_n1328));
  AND3_X1   g1128(.A1(new_n1327), .A2(new_n1328), .A3(new_n1308), .ZN(new_n1329));
  AOI21_X1  g1129(.A(new_n1328), .B1(new_n1327), .B2(new_n1308), .ZN(new_n1330));
  NOR2_X1   g1130(.A1(new_n1327), .A2(new_n1308), .ZN(new_n1331));
  NOR3_X1   g1131(.A1(new_n1329), .A2(new_n1330), .A3(new_n1331), .ZN(G402));
endmodule


