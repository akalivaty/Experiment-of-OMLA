

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302,
         n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313,
         n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324,
         n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335,
         n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346,
         n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357,
         n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368,
         n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379,
         n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390,
         n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
         n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412,
         n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423,
         n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
         n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445,
         n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456,
         n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467,
         n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478,
         n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489,
         n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500,
         n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511,
         n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588,
         n589, n590, n591, n592, n593;

  XNOR2_X1 U324 ( .A(n399), .B(n398), .ZN(n400) );
  XNOR2_X1 U325 ( .A(n411), .B(n410), .ZN(n415) );
  INV_X1 U326 ( .A(KEYINPUT77), .ZN(n396) );
  XNOR2_X1 U327 ( .A(n397), .B(n396), .ZN(n398) );
  INV_X1 U328 ( .A(n432), .ZN(n408) );
  XNOR2_X1 U329 ( .A(n409), .B(n408), .ZN(n410) );
  XNOR2_X1 U330 ( .A(KEYINPUT64), .B(KEYINPUT48), .ZN(n426) );
  NOR2_X1 U331 ( .A1(n525), .A2(n445), .ZN(n579) );
  XNOR2_X1 U332 ( .A(n427), .B(n426), .ZN(n537) );
  XOR2_X1 U333 ( .A(n464), .B(n463), .Z(n539) );
  XNOR2_X1 U334 ( .A(n466), .B(G190GAT), .ZN(n467) );
  XNOR2_X1 U335 ( .A(n468), .B(n467), .ZN(G1351GAT) );
  XOR2_X1 U336 ( .A(KEYINPUT85), .B(KEYINPUT9), .Z(n293) );
  XNOR2_X1 U337 ( .A(G162GAT), .B(G106GAT), .ZN(n292) );
  XOR2_X1 U338 ( .A(n293), .B(n292), .Z(n316) );
  INV_X1 U339 ( .A(KEYINPUT65), .ZN(n294) );
  NAND2_X1 U340 ( .A1(KEYINPUT11), .A2(n294), .ZN(n297) );
  INV_X1 U341 ( .A(KEYINPUT11), .ZN(n295) );
  NAND2_X1 U342 ( .A1(n295), .A2(KEYINPUT65), .ZN(n296) );
  NAND2_X1 U343 ( .A1(n297), .A2(n296), .ZN(n299) );
  NAND2_X1 U344 ( .A1(G232GAT), .A2(G233GAT), .ZN(n298) );
  XNOR2_X1 U345 ( .A(n299), .B(n298), .ZN(n301) );
  INV_X1 U346 ( .A(KEYINPUT10), .ZN(n300) );
  XOR2_X1 U347 ( .A(n301), .B(n300), .Z(n305) );
  XNOR2_X1 U348 ( .A(G43GAT), .B(KEYINPUT7), .ZN(n302) );
  XNOR2_X1 U349 ( .A(n302), .B(KEYINPUT8), .ZN(n354) );
  XNOR2_X1 U350 ( .A(G36GAT), .B(G190GAT), .ZN(n303) );
  XNOR2_X1 U351 ( .A(n303), .B(G218GAT), .ZN(n438) );
  XNOR2_X1 U352 ( .A(n354), .B(n438), .ZN(n304) );
  XNOR2_X1 U353 ( .A(n305), .B(n304), .ZN(n312) );
  INV_X1 U354 ( .A(KEYINPUT78), .ZN(n306) );
  NAND2_X1 U355 ( .A1(n306), .A2(G92GAT), .ZN(n309) );
  INV_X1 U356 ( .A(G92GAT), .ZN(n307) );
  NAND2_X1 U357 ( .A1(n307), .A2(KEYINPUT78), .ZN(n308) );
  NAND2_X1 U358 ( .A1(n309), .A2(n308), .ZN(n311) );
  XNOR2_X1 U359 ( .A(G99GAT), .B(G85GAT), .ZN(n310) );
  XNOR2_X1 U360 ( .A(n311), .B(n310), .ZN(n399) );
  XNOR2_X1 U361 ( .A(n312), .B(n399), .ZN(n314) );
  XOR2_X1 U362 ( .A(G50GAT), .B(KEYINPUT84), .Z(n319) );
  XOR2_X1 U363 ( .A(G29GAT), .B(G134GAT), .Z(n343) );
  XNOR2_X1 U364 ( .A(n319), .B(n343), .ZN(n313) );
  XNOR2_X1 U365 ( .A(n314), .B(n313), .ZN(n315) );
  XNOR2_X1 U366 ( .A(n316), .B(n315), .ZN(n552) );
  INV_X1 U367 ( .A(n552), .ZN(n566) );
  XOR2_X1 U368 ( .A(G211GAT), .B(KEYINPUT94), .Z(n318) );
  XNOR2_X1 U369 ( .A(G22GAT), .B(KEYINPUT22), .ZN(n317) );
  XNOR2_X1 U370 ( .A(n318), .B(n317), .ZN(n323) );
  XOR2_X1 U371 ( .A(KEYINPUT24), .B(G218GAT), .Z(n321) );
  XOR2_X1 U372 ( .A(G197GAT), .B(KEYINPUT21), .Z(n433) );
  XNOR2_X1 U373 ( .A(n319), .B(n433), .ZN(n320) );
  XNOR2_X1 U374 ( .A(n321), .B(n320), .ZN(n322) );
  XOR2_X1 U375 ( .A(n323), .B(n322), .Z(n325) );
  NAND2_X1 U376 ( .A1(G228GAT), .A2(G233GAT), .ZN(n324) );
  XNOR2_X1 U377 ( .A(n325), .B(n324), .ZN(n329) );
  XOR2_X1 U378 ( .A(KEYINPUT23), .B(KEYINPUT93), .Z(n327) );
  XNOR2_X1 U379 ( .A(G148GAT), .B(G155GAT), .ZN(n326) );
  XNOR2_X1 U380 ( .A(n327), .B(n326), .ZN(n328) );
  XOR2_X1 U381 ( .A(n329), .B(n328), .Z(n334) );
  XOR2_X1 U382 ( .A(KEYINPUT2), .B(KEYINPUT3), .Z(n331) );
  XNOR2_X1 U383 ( .A(G141GAT), .B(G162GAT), .ZN(n330) );
  XNOR2_X1 U384 ( .A(n331), .B(n330), .ZN(n349) );
  XNOR2_X1 U385 ( .A(G106GAT), .B(G78GAT), .ZN(n332) );
  XNOR2_X1 U386 ( .A(n332), .B(G204GAT), .ZN(n413) );
  XNOR2_X1 U387 ( .A(n349), .B(n413), .ZN(n333) );
  XNOR2_X1 U388 ( .A(n334), .B(n333), .ZN(n475) );
  XOR2_X1 U389 ( .A(KEYINPUT95), .B(KEYINPUT98), .Z(n336) );
  XNOR2_X1 U390 ( .A(KEYINPUT96), .B(KEYINPUT4), .ZN(n335) );
  XNOR2_X1 U391 ( .A(n336), .B(n335), .ZN(n353) );
  XOR2_X1 U392 ( .A(KEYINPUT97), .B(KEYINPUT6), .Z(n338) );
  XNOR2_X1 U393 ( .A(KEYINPUT1), .B(KEYINPUT5), .ZN(n337) );
  XNOR2_X1 U394 ( .A(n338), .B(n337), .ZN(n339) );
  XOR2_X1 U395 ( .A(n339), .B(G57GAT), .Z(n341) );
  XOR2_X1 U396 ( .A(G120GAT), .B(G148GAT), .Z(n412) );
  XNOR2_X1 U397 ( .A(n412), .B(G85GAT), .ZN(n340) );
  XNOR2_X1 U398 ( .A(n341), .B(n340), .ZN(n347) );
  XNOR2_X1 U399 ( .A(G1GAT), .B(G127GAT), .ZN(n342) );
  XNOR2_X1 U400 ( .A(n342), .B(G155GAT), .ZN(n386) );
  XOR2_X1 U401 ( .A(n386), .B(n343), .Z(n345) );
  NAND2_X1 U402 ( .A1(G225GAT), .A2(G233GAT), .ZN(n344) );
  XNOR2_X1 U403 ( .A(n345), .B(n344), .ZN(n346) );
  XOR2_X1 U404 ( .A(n347), .B(n346), .Z(n351) );
  XNOR2_X1 U405 ( .A(G113GAT), .B(KEYINPUT0), .ZN(n348) );
  XNOR2_X1 U406 ( .A(n348), .B(KEYINPUT88), .ZN(n456) );
  XNOR2_X1 U407 ( .A(n456), .B(n349), .ZN(n350) );
  XNOR2_X1 U408 ( .A(n351), .B(n350), .ZN(n352) );
  XOR2_X1 U409 ( .A(n353), .B(n352), .Z(n481) );
  XNOR2_X1 U410 ( .A(KEYINPUT99), .B(n481), .ZN(n525) );
  XOR2_X1 U411 ( .A(n354), .B(G8GAT), .Z(n356) );
  NAND2_X1 U412 ( .A1(G229GAT), .A2(G233GAT), .ZN(n355) );
  XNOR2_X1 U413 ( .A(n356), .B(n355), .ZN(n360) );
  XOR2_X1 U414 ( .A(KEYINPUT29), .B(KEYINPUT67), .Z(n358) );
  XNOR2_X1 U415 ( .A(KEYINPUT71), .B(KEYINPUT73), .ZN(n357) );
  XNOR2_X1 U416 ( .A(n358), .B(n357), .ZN(n359) );
  XNOR2_X1 U417 ( .A(n360), .B(n359), .ZN(n364) );
  XOR2_X1 U418 ( .A(KEYINPUT69), .B(G113GAT), .Z(n362) );
  XNOR2_X1 U419 ( .A(G169GAT), .B(G141GAT), .ZN(n361) );
  XNOR2_X1 U420 ( .A(n362), .B(n361), .ZN(n363) );
  XNOR2_X1 U421 ( .A(n364), .B(n363), .ZN(n369) );
  XOR2_X1 U422 ( .A(G50GAT), .B(G36GAT), .Z(n367) );
  XNOR2_X1 U423 ( .A(G22GAT), .B(G15GAT), .ZN(n365) );
  XNOR2_X1 U424 ( .A(n365), .B(KEYINPUT72), .ZN(n388) );
  XNOR2_X1 U425 ( .A(G197GAT), .B(n388), .ZN(n366) );
  XNOR2_X1 U426 ( .A(n367), .B(n366), .ZN(n368) );
  XOR2_X1 U427 ( .A(n369), .B(n368), .Z(n374) );
  XOR2_X1 U428 ( .A(G1GAT), .B(KEYINPUT70), .Z(n371) );
  XNOR2_X1 U429 ( .A(KEYINPUT30), .B(KEYINPUT68), .ZN(n370) );
  XNOR2_X1 U430 ( .A(n371), .B(n370), .ZN(n372) );
  XNOR2_X1 U431 ( .A(n372), .B(G29GAT), .ZN(n373) );
  XNOR2_X1 U432 ( .A(n374), .B(n373), .ZN(n580) );
  XNOR2_X1 U433 ( .A(n552), .B(KEYINPUT105), .ZN(n375) );
  XNOR2_X1 U434 ( .A(n375), .B(KEYINPUT36), .ZN(n591) );
  XOR2_X1 U435 ( .A(KEYINPUT74), .B(KEYINPUT75), .Z(n377) );
  XNOR2_X1 U436 ( .A(G71GAT), .B(KEYINPUT13), .ZN(n376) );
  XNOR2_X1 U437 ( .A(n377), .B(n376), .ZN(n378) );
  XOR2_X1 U438 ( .A(G57GAT), .B(n378), .Z(n401) );
  XOR2_X1 U439 ( .A(KEYINPUT87), .B(KEYINPUT15), .Z(n380) );
  XNOR2_X1 U440 ( .A(KEYINPUT14), .B(KEYINPUT12), .ZN(n379) );
  XNOR2_X1 U441 ( .A(n380), .B(n379), .ZN(n381) );
  XNOR2_X1 U442 ( .A(n401), .B(n381), .ZN(n392) );
  XOR2_X1 U443 ( .A(KEYINPUT86), .B(G211GAT), .Z(n383) );
  XNOR2_X1 U444 ( .A(G8GAT), .B(G183GAT), .ZN(n382) );
  XNOR2_X1 U445 ( .A(n383), .B(n382), .ZN(n436) );
  XOR2_X1 U446 ( .A(n436), .B(G64GAT), .Z(n385) );
  NAND2_X1 U447 ( .A1(G231GAT), .A2(G233GAT), .ZN(n384) );
  XNOR2_X1 U448 ( .A(n385), .B(n384), .ZN(n387) );
  XOR2_X1 U449 ( .A(n387), .B(n386), .Z(n390) );
  XNOR2_X1 U450 ( .A(n388), .B(G78GAT), .ZN(n389) );
  XNOR2_X1 U451 ( .A(n390), .B(n389), .ZN(n391) );
  XNOR2_X1 U452 ( .A(n392), .B(n391), .ZN(n563) );
  NOR2_X1 U453 ( .A1(n591), .A2(n563), .ZN(n394) );
  XNOR2_X1 U454 ( .A(KEYINPUT66), .B(KEYINPUT45), .ZN(n393) );
  XNOR2_X1 U455 ( .A(n394), .B(n393), .ZN(n395) );
  NAND2_X1 U456 ( .A1(n580), .A2(n395), .ZN(n416) );
  NAND2_X1 U457 ( .A1(G230GAT), .A2(G233GAT), .ZN(n397) );
  XNOR2_X1 U458 ( .A(n401), .B(n400), .ZN(n411) );
  XOR2_X1 U459 ( .A(KEYINPUT81), .B(KEYINPUT79), .Z(n403) );
  XNOR2_X1 U460 ( .A(KEYINPUT31), .B(KEYINPUT82), .ZN(n402) );
  XNOR2_X1 U461 ( .A(n403), .B(n402), .ZN(n407) );
  XOR2_X1 U462 ( .A(KEYINPUT32), .B(KEYINPUT80), .Z(n405) );
  XNOR2_X1 U463 ( .A(KEYINPUT33), .B(KEYINPUT76), .ZN(n404) );
  XNOR2_X1 U464 ( .A(n405), .B(n404), .ZN(n406) );
  XOR2_X1 U465 ( .A(n407), .B(n406), .Z(n409) );
  XOR2_X1 U466 ( .A(G176GAT), .B(G64GAT), .Z(n432) );
  XNOR2_X1 U467 ( .A(n413), .B(n412), .ZN(n414) );
  XNOR2_X1 U468 ( .A(n415), .B(n414), .ZN(n418) );
  NOR2_X1 U469 ( .A1(n416), .A2(n418), .ZN(n417) );
  XNOR2_X1 U470 ( .A(n417), .B(KEYINPUT119), .ZN(n425) );
  XNOR2_X1 U471 ( .A(KEYINPUT41), .B(n418), .ZN(n559) );
  NOR2_X1 U472 ( .A1(n559), .A2(n580), .ZN(n420) );
  XOR2_X1 U473 ( .A(KEYINPUT118), .B(KEYINPUT46), .Z(n419) );
  XNOR2_X1 U474 ( .A(n420), .B(n419), .ZN(n422) );
  INV_X1 U475 ( .A(n563), .ZN(n588) );
  XNOR2_X1 U476 ( .A(KEYINPUT117), .B(n588), .ZN(n576) );
  AND2_X1 U477 ( .A1(n576), .A2(n566), .ZN(n421) );
  AND2_X1 U478 ( .A1(n422), .A2(n421), .ZN(n423) );
  XNOR2_X1 U479 ( .A(n423), .B(KEYINPUT47), .ZN(n424) );
  AND2_X1 U480 ( .A1(n425), .A2(n424), .ZN(n427) );
  XNOR2_X1 U481 ( .A(KEYINPUT91), .B(KEYINPUT17), .ZN(n428) );
  XNOR2_X1 U482 ( .A(n428), .B(KEYINPUT19), .ZN(n429) );
  XOR2_X1 U483 ( .A(n429), .B(KEYINPUT90), .Z(n431) );
  XNOR2_X1 U484 ( .A(G169GAT), .B(KEYINPUT18), .ZN(n430) );
  XNOR2_X1 U485 ( .A(n431), .B(n430), .ZN(n460) );
  XNOR2_X1 U486 ( .A(n433), .B(n432), .ZN(n442) );
  XOR2_X1 U487 ( .A(G92GAT), .B(KEYINPUT100), .Z(n435) );
  NAND2_X1 U488 ( .A1(G226GAT), .A2(G233GAT), .ZN(n434) );
  XNOR2_X1 U489 ( .A(n435), .B(n434), .ZN(n437) );
  XOR2_X1 U490 ( .A(n437), .B(n436), .Z(n440) );
  XNOR2_X1 U491 ( .A(G204GAT), .B(n438), .ZN(n439) );
  XNOR2_X1 U492 ( .A(n440), .B(n439), .ZN(n441) );
  XNOR2_X1 U493 ( .A(n442), .B(n441), .ZN(n443) );
  XNOR2_X1 U494 ( .A(n460), .B(n443), .ZN(n474) );
  NOR2_X1 U495 ( .A1(n537), .A2(n474), .ZN(n444) );
  XOR2_X1 U496 ( .A(KEYINPUT54), .B(n444), .Z(n445) );
  NAND2_X1 U497 ( .A1(n475), .A2(n579), .ZN(n446) );
  XNOR2_X1 U498 ( .A(n446), .B(KEYINPUT55), .ZN(n447) );
  XNOR2_X1 U499 ( .A(n447), .B(KEYINPUT124), .ZN(n465) );
  XOR2_X1 U500 ( .A(G176GAT), .B(G183GAT), .Z(n449) );
  XNOR2_X1 U501 ( .A(KEYINPUT92), .B(KEYINPUT89), .ZN(n448) );
  XNOR2_X1 U502 ( .A(n449), .B(n448), .ZN(n464) );
  XOR2_X1 U503 ( .A(G99GAT), .B(G134GAT), .Z(n451) );
  XNOR2_X1 U504 ( .A(G43GAT), .B(G190GAT), .ZN(n450) );
  XNOR2_X1 U505 ( .A(n451), .B(n450), .ZN(n455) );
  XOR2_X1 U506 ( .A(KEYINPUT20), .B(G127GAT), .Z(n453) );
  XNOR2_X1 U507 ( .A(G15GAT), .B(G120GAT), .ZN(n452) );
  XNOR2_X1 U508 ( .A(n453), .B(n452), .ZN(n454) );
  XOR2_X1 U509 ( .A(n455), .B(n454), .Z(n462) );
  XOR2_X1 U510 ( .A(n456), .B(G71GAT), .Z(n458) );
  NAND2_X1 U511 ( .A1(G227GAT), .A2(G233GAT), .ZN(n457) );
  XNOR2_X1 U512 ( .A(n458), .B(n457), .ZN(n459) );
  XNOR2_X1 U513 ( .A(n460), .B(n459), .ZN(n461) );
  XNOR2_X1 U514 ( .A(n462), .B(n461), .ZN(n463) );
  NAND2_X1 U515 ( .A1(n465), .A2(n539), .ZN(n575) );
  NOR2_X1 U516 ( .A1(n566), .A2(n575), .ZN(n468) );
  INV_X1 U517 ( .A(KEYINPUT58), .ZN(n466) );
  NOR2_X1 U518 ( .A1(n580), .A2(n418), .ZN(n469) );
  XOR2_X1 U519 ( .A(KEYINPUT83), .B(n469), .Z(n499) );
  INV_X1 U520 ( .A(n539), .ZN(n471) );
  XOR2_X1 U521 ( .A(n475), .B(KEYINPUT28), .Z(n532) );
  XOR2_X1 U522 ( .A(KEYINPUT27), .B(n474), .Z(n473) );
  NAND2_X1 U523 ( .A1(n525), .A2(n473), .ZN(n556) );
  NOR2_X1 U524 ( .A1(n532), .A2(n556), .ZN(n538) );
  XOR2_X1 U525 ( .A(n538), .B(KEYINPUT101), .Z(n470) );
  NAND2_X1 U526 ( .A1(n471), .A2(n470), .ZN(n484) );
  NOR2_X1 U527 ( .A1(n475), .A2(n539), .ZN(n472) );
  XNOR2_X1 U528 ( .A(n472), .B(KEYINPUT26), .ZN(n578) );
  NAND2_X1 U529 ( .A1(n473), .A2(n578), .ZN(n480) );
  INV_X1 U530 ( .A(n474), .ZN(n527) );
  NAND2_X1 U531 ( .A1(n527), .A2(n539), .ZN(n476) );
  NAND2_X1 U532 ( .A1(n476), .A2(n475), .ZN(n477) );
  XNOR2_X1 U533 ( .A(n477), .B(KEYINPUT25), .ZN(n478) );
  XOR2_X1 U534 ( .A(KEYINPUT102), .B(n478), .Z(n479) );
  NAND2_X1 U535 ( .A1(n480), .A2(n479), .ZN(n482) );
  NAND2_X1 U536 ( .A1(n482), .A2(n481), .ZN(n483) );
  NAND2_X1 U537 ( .A1(n484), .A2(n483), .ZN(n485) );
  XNOR2_X1 U538 ( .A(n485), .B(KEYINPUT103), .ZN(n496) );
  NOR2_X1 U539 ( .A1(n552), .A2(n563), .ZN(n486) );
  XOR2_X1 U540 ( .A(KEYINPUT16), .B(n486), .Z(n487) );
  NOR2_X1 U541 ( .A1(n496), .A2(n487), .ZN(n510) );
  AND2_X1 U542 ( .A1(n499), .A2(n510), .ZN(n494) );
  NAND2_X1 U543 ( .A1(n525), .A2(n494), .ZN(n488) );
  XNOR2_X1 U544 ( .A(n488), .B(KEYINPUT34), .ZN(n489) );
  XNOR2_X1 U545 ( .A(G1GAT), .B(n489), .ZN(G1324GAT) );
  NAND2_X1 U546 ( .A1(n494), .A2(n527), .ZN(n490) );
  XNOR2_X1 U547 ( .A(n490), .B(G8GAT), .ZN(G1325GAT) );
  XOR2_X1 U548 ( .A(KEYINPUT104), .B(KEYINPUT35), .Z(n492) );
  NAND2_X1 U549 ( .A1(n494), .A2(n539), .ZN(n491) );
  XNOR2_X1 U550 ( .A(n492), .B(n491), .ZN(n493) );
  XNOR2_X1 U551 ( .A(G15GAT), .B(n493), .ZN(G1326GAT) );
  NAND2_X1 U552 ( .A1(n494), .A2(n532), .ZN(n495) );
  XNOR2_X1 U553 ( .A(n495), .B(G22GAT), .ZN(G1327GAT) );
  XOR2_X1 U554 ( .A(G29GAT), .B(KEYINPUT39), .Z(n503) );
  XOR2_X1 U555 ( .A(KEYINPUT38), .B(KEYINPUT106), .Z(n501) );
  NOR2_X1 U556 ( .A1(n591), .A2(n496), .ZN(n497) );
  NAND2_X1 U557 ( .A1(n563), .A2(n497), .ZN(n498) );
  XNOR2_X1 U558 ( .A(KEYINPUT37), .B(n498), .ZN(n522) );
  NAND2_X1 U559 ( .A1(n499), .A2(n522), .ZN(n500) );
  XNOR2_X1 U560 ( .A(n501), .B(n500), .ZN(n508) );
  NAND2_X1 U561 ( .A1(n508), .A2(n525), .ZN(n502) );
  XNOR2_X1 U562 ( .A(n503), .B(n502), .ZN(G1328GAT) );
  NAND2_X1 U563 ( .A1(n508), .A2(n527), .ZN(n504) );
  XNOR2_X1 U564 ( .A(n504), .B(G36GAT), .ZN(G1329GAT) );
  XOR2_X1 U565 ( .A(KEYINPUT40), .B(KEYINPUT107), .Z(n506) );
  NAND2_X1 U566 ( .A1(n508), .A2(n539), .ZN(n505) );
  XNOR2_X1 U567 ( .A(n506), .B(n505), .ZN(n507) );
  XNOR2_X1 U568 ( .A(G43GAT), .B(n507), .ZN(G1330GAT) );
  NAND2_X1 U569 ( .A1(n508), .A2(n532), .ZN(n509) );
  XNOR2_X1 U570 ( .A(n509), .B(G50GAT), .ZN(G1331GAT) );
  XNOR2_X1 U571 ( .A(KEYINPUT108), .B(n559), .ZN(n569) );
  INV_X1 U572 ( .A(n580), .ZN(n541) );
  NOR2_X1 U573 ( .A1(n569), .A2(n541), .ZN(n523) );
  AND2_X1 U574 ( .A1(n523), .A2(n510), .ZN(n518) );
  NAND2_X1 U575 ( .A1(n518), .A2(n525), .ZN(n511) );
  XNOR2_X1 U576 ( .A(KEYINPUT42), .B(n511), .ZN(n512) );
  XNOR2_X1 U577 ( .A(G57GAT), .B(n512), .ZN(G1332GAT) );
  XOR2_X1 U578 ( .A(KEYINPUT109), .B(KEYINPUT110), .Z(n514) );
  NAND2_X1 U579 ( .A1(n518), .A2(n527), .ZN(n513) );
  XNOR2_X1 U580 ( .A(n514), .B(n513), .ZN(n515) );
  XNOR2_X1 U581 ( .A(G64GAT), .B(n515), .ZN(G1333GAT) );
  XOR2_X1 U582 ( .A(G71GAT), .B(KEYINPUT111), .Z(n517) );
  NAND2_X1 U583 ( .A1(n518), .A2(n539), .ZN(n516) );
  XNOR2_X1 U584 ( .A(n517), .B(n516), .ZN(G1334GAT) );
  XOR2_X1 U585 ( .A(KEYINPUT112), .B(KEYINPUT43), .Z(n520) );
  NAND2_X1 U586 ( .A1(n518), .A2(n532), .ZN(n519) );
  XNOR2_X1 U587 ( .A(n520), .B(n519), .ZN(n521) );
  XNOR2_X1 U588 ( .A(G78GAT), .B(n521), .ZN(G1335GAT) );
  NAND2_X1 U589 ( .A1(n523), .A2(n522), .ZN(n524) );
  XNOR2_X1 U590 ( .A(n524), .B(KEYINPUT113), .ZN(n533) );
  NAND2_X1 U591 ( .A1(n525), .A2(n533), .ZN(n526) );
  XNOR2_X1 U592 ( .A(n526), .B(G85GAT), .ZN(G1336GAT) );
  NAND2_X1 U593 ( .A1(n533), .A2(n527), .ZN(n528) );
  XNOR2_X1 U594 ( .A(n528), .B(G92GAT), .ZN(G1337GAT) );
  XOR2_X1 U595 ( .A(KEYINPUT114), .B(KEYINPUT115), .Z(n530) );
  NAND2_X1 U596 ( .A1(n533), .A2(n539), .ZN(n529) );
  XNOR2_X1 U597 ( .A(n530), .B(n529), .ZN(n531) );
  XNOR2_X1 U598 ( .A(G99GAT), .B(n531), .ZN(G1338GAT) );
  XOR2_X1 U599 ( .A(KEYINPUT116), .B(KEYINPUT44), .Z(n535) );
  NAND2_X1 U600 ( .A1(n533), .A2(n532), .ZN(n534) );
  XNOR2_X1 U601 ( .A(n535), .B(n534), .ZN(n536) );
  XOR2_X1 U602 ( .A(G106GAT), .B(n536), .Z(G1339GAT) );
  NAND2_X1 U603 ( .A1(n539), .A2(n538), .ZN(n540) );
  NOR2_X1 U604 ( .A1(n537), .A2(n540), .ZN(n553) );
  NAND2_X1 U605 ( .A1(n541), .A2(n553), .ZN(n542) );
  XNOR2_X1 U606 ( .A(n542), .B(KEYINPUT120), .ZN(n543) );
  XNOR2_X1 U607 ( .A(G113GAT), .B(n543), .ZN(G1340GAT) );
  INV_X1 U608 ( .A(n553), .ZN(n548) );
  NOR2_X1 U609 ( .A1(n548), .A2(n569), .ZN(n547) );
  XOR2_X1 U610 ( .A(KEYINPUT121), .B(KEYINPUT122), .Z(n545) );
  XNOR2_X1 U611 ( .A(G120GAT), .B(KEYINPUT49), .ZN(n544) );
  XNOR2_X1 U612 ( .A(n545), .B(n544), .ZN(n546) );
  XNOR2_X1 U613 ( .A(n547), .B(n546), .ZN(G1341GAT) );
  NOR2_X1 U614 ( .A1(n576), .A2(n548), .ZN(n550) );
  XNOR2_X1 U615 ( .A(KEYINPUT123), .B(KEYINPUT50), .ZN(n549) );
  XNOR2_X1 U616 ( .A(n550), .B(n549), .ZN(n551) );
  XNOR2_X1 U617 ( .A(G127GAT), .B(n551), .ZN(G1342GAT) );
  XOR2_X1 U618 ( .A(G134GAT), .B(KEYINPUT51), .Z(n555) );
  NAND2_X1 U619 ( .A1(n553), .A2(n552), .ZN(n554) );
  XNOR2_X1 U620 ( .A(n555), .B(n554), .ZN(G1343GAT) );
  NOR2_X1 U621 ( .A1(n537), .A2(n556), .ZN(n557) );
  NAND2_X1 U622 ( .A1(n557), .A2(n578), .ZN(n565) );
  NOR2_X1 U623 ( .A1(n580), .A2(n565), .ZN(n558) );
  XOR2_X1 U624 ( .A(G141GAT), .B(n558), .Z(G1344GAT) );
  NOR2_X1 U625 ( .A1(n559), .A2(n565), .ZN(n561) );
  XNOR2_X1 U626 ( .A(KEYINPUT53), .B(KEYINPUT52), .ZN(n560) );
  XNOR2_X1 U627 ( .A(n561), .B(n560), .ZN(n562) );
  XNOR2_X1 U628 ( .A(G148GAT), .B(n562), .ZN(G1345GAT) );
  NOR2_X1 U629 ( .A1(n563), .A2(n565), .ZN(n564) );
  XOR2_X1 U630 ( .A(G155GAT), .B(n564), .Z(G1346GAT) );
  NOR2_X1 U631 ( .A1(n566), .A2(n565), .ZN(n567) );
  XOR2_X1 U632 ( .A(G162GAT), .B(n567), .Z(G1347GAT) );
  NOR2_X1 U633 ( .A1(n580), .A2(n575), .ZN(n568) );
  XOR2_X1 U634 ( .A(G169GAT), .B(n568), .Z(G1348GAT) );
  NOR2_X1 U635 ( .A1(n569), .A2(n575), .ZN(n574) );
  XOR2_X1 U636 ( .A(KEYINPUT57), .B(KEYINPUT126), .Z(n571) );
  XNOR2_X1 U637 ( .A(G176GAT), .B(KEYINPUT125), .ZN(n570) );
  XNOR2_X1 U638 ( .A(n571), .B(n570), .ZN(n572) );
  XNOR2_X1 U639 ( .A(KEYINPUT56), .B(n572), .ZN(n573) );
  XNOR2_X1 U640 ( .A(n574), .B(n573), .ZN(G1349GAT) );
  NOR2_X1 U641 ( .A1(n576), .A2(n575), .ZN(n577) );
  XOR2_X1 U642 ( .A(G183GAT), .B(n577), .Z(G1350GAT) );
  NAND2_X1 U643 ( .A1(n579), .A2(n578), .ZN(n590) );
  NOR2_X1 U644 ( .A1(n580), .A2(n590), .ZN(n582) );
  XNOR2_X1 U645 ( .A(KEYINPUT60), .B(KEYINPUT59), .ZN(n581) );
  XNOR2_X1 U646 ( .A(n582), .B(n581), .ZN(n583) );
  XNOR2_X1 U647 ( .A(G197GAT), .B(n583), .ZN(G1352GAT) );
  XOR2_X1 U648 ( .A(KEYINPUT127), .B(KEYINPUT61), .Z(n585) );
  INV_X1 U649 ( .A(n590), .ZN(n587) );
  NAND2_X1 U650 ( .A1(n587), .A2(n418), .ZN(n584) );
  XNOR2_X1 U651 ( .A(n585), .B(n584), .ZN(n586) );
  XOR2_X1 U652 ( .A(G204GAT), .B(n586), .Z(G1353GAT) );
  NAND2_X1 U653 ( .A1(n588), .A2(n587), .ZN(n589) );
  XNOR2_X1 U654 ( .A(n589), .B(G211GAT), .ZN(G1354GAT) );
  NOR2_X1 U655 ( .A1(n591), .A2(n590), .ZN(n592) );
  XOR2_X1 U656 ( .A(KEYINPUT62), .B(n592), .Z(n593) );
  XNOR2_X1 U657 ( .A(G218GAT), .B(n593), .ZN(G1355GAT) );
endmodule

