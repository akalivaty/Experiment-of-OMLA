//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 1 1 1 1 1 1 1 0 0 0 0 0 0 0 1 1 1 0 1 0 0 0 1 1 0 1 1 0 1 0 1 1 1 1 0 0 0 0 0 0 1 0 0 0 0 0 0 0 1 0 0 1 0 0 1 0 1 1 0 0 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:30:37 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n448, new_n449, new_n452, new_n453, new_n454, new_n455,
    new_n458, new_n459, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n498, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n516, new_n517, new_n518, new_n519,
    new_n520, new_n521, new_n522, new_n523, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n531, new_n532, new_n533, new_n534, new_n535,
    new_n536, new_n537, new_n538, new_n539, new_n540, new_n541, new_n542,
    new_n545, new_n546, new_n548, new_n549, new_n550, new_n551, new_n552,
    new_n553, new_n554, new_n555, new_n556, new_n557, new_n558, new_n559,
    new_n560, new_n561, new_n562, new_n566, new_n567, new_n568, new_n569,
    new_n571, new_n572, new_n573, new_n574, new_n575, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n601, new_n604,
    new_n606, new_n607, new_n608, new_n609, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1190,
    new_n1191, new_n1192;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  XOR2_X1   g002(.A(KEYINPUT64), .B(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  XOR2_X1   g011(.A(KEYINPUT65), .B(G96), .Z(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  INV_X1    g022(.A(G567), .ZN(new_n448));
  NOR2_X1   g023(.A1(new_n446), .A2(new_n448), .ZN(new_n449));
  XOR2_X1   g024(.A(new_n449), .B(KEYINPUT66), .Z(G234));
  NAND3_X1  g025(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g026(.A1(G221), .A2(G220), .A3(G218), .A4(G219), .ZN(new_n452));
  XNOR2_X1  g027(.A(new_n452), .B(KEYINPUT2), .ZN(new_n453));
  NOR4_X1   g028(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n454));
  NAND2_X1  g029(.A1(new_n453), .A2(new_n454), .ZN(new_n455));
  XNOR2_X1  g030(.A(new_n455), .B(KEYINPUT67), .ZN(G261));
  INV_X1    g031(.A(G261), .ZN(G325));
  INV_X1    g032(.A(G2106), .ZN(new_n458));
  OAI22_X1  g033(.A1(new_n453), .A2(new_n458), .B1(new_n448), .B2(new_n454), .ZN(new_n459));
  INV_X1    g034(.A(new_n459), .ZN(G319));
  INV_X1    g035(.A(KEYINPUT68), .ZN(new_n461));
  INV_X1    g036(.A(KEYINPUT3), .ZN(new_n462));
  OAI21_X1  g037(.A(new_n461), .B1(new_n462), .B2(G2104), .ZN(new_n463));
  INV_X1    g038(.A(G2104), .ZN(new_n464));
  NAND3_X1  g039(.A1(new_n464), .A2(KEYINPUT68), .A3(KEYINPUT3), .ZN(new_n465));
  INV_X1    g040(.A(G2105), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n462), .A2(G2104), .ZN(new_n467));
  NAND4_X1  g042(.A1(new_n463), .A2(new_n465), .A3(new_n466), .A4(new_n467), .ZN(new_n468));
  INV_X1    g043(.A(G137), .ZN(new_n469));
  NOR2_X1   g044(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n464), .A2(KEYINPUT3), .ZN(new_n471));
  NAND3_X1  g046(.A1(new_n471), .A2(new_n467), .A3(G125), .ZN(new_n472));
  NAND2_X1  g047(.A1(G113), .A2(G2104), .ZN(new_n473));
  AOI21_X1  g048(.A(new_n466), .B1(new_n472), .B2(new_n473), .ZN(new_n474));
  NOR2_X1   g049(.A1(new_n464), .A2(G2105), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n475), .A2(G101), .ZN(new_n476));
  INV_X1    g051(.A(new_n476), .ZN(new_n477));
  NOR3_X1   g052(.A1(new_n470), .A2(new_n474), .A3(new_n477), .ZN(G160));
  NAND4_X1  g053(.A1(new_n463), .A2(new_n465), .A3(G2105), .A4(new_n467), .ZN(new_n479));
  INV_X1    g054(.A(G124), .ZN(new_n480));
  NOR2_X1   g055(.A1(new_n466), .A2(G112), .ZN(new_n481));
  OAI21_X1  g056(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n482));
  OAI22_X1  g057(.A1(new_n479), .A2(new_n480), .B1(new_n481), .B2(new_n482), .ZN(new_n483));
  INV_X1    g058(.A(new_n468), .ZN(new_n484));
  AOI21_X1  g059(.A(new_n483), .B1(new_n484), .B2(G136), .ZN(G162));
  INV_X1    g060(.A(G138), .ZN(new_n486));
  NOR2_X1   g061(.A1(new_n486), .A2(G2105), .ZN(new_n487));
  NAND4_X1  g062(.A1(new_n463), .A2(new_n465), .A3(new_n487), .A4(new_n467), .ZN(new_n488));
  AND2_X1   g063(.A1(new_n471), .A2(new_n467), .ZN(new_n489));
  NOR3_X1   g064(.A1(new_n486), .A2(KEYINPUT4), .A3(G2105), .ZN(new_n490));
  AOI22_X1  g065(.A1(new_n488), .A2(KEYINPUT4), .B1(new_n489), .B2(new_n490), .ZN(new_n491));
  OR2_X1    g066(.A1(G102), .A2(G2105), .ZN(new_n492));
  OAI211_X1 g067(.A(new_n492), .B(G2104), .C1(G114), .C2(new_n466), .ZN(new_n493));
  INV_X1    g068(.A(G126), .ZN(new_n494));
  OAI21_X1  g069(.A(new_n493), .B1(new_n479), .B2(new_n494), .ZN(new_n495));
  OR2_X1    g070(.A1(new_n491), .A2(new_n495), .ZN(new_n496));
  INV_X1    g071(.A(new_n496), .ZN(G164));
  XNOR2_X1  g072(.A(KEYINPUT5), .B(G543), .ZN(new_n498));
  AOI22_X1  g073(.A1(new_n498), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n499));
  INV_X1    g074(.A(G651), .ZN(new_n500));
  NOR2_X1   g075(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  OR2_X1    g076(.A1(KEYINPUT6), .A2(G651), .ZN(new_n502));
  NAND2_X1  g077(.A1(KEYINPUT6), .A2(G651), .ZN(new_n503));
  NAND2_X1  g078(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  NAND2_X1  g079(.A1(new_n504), .A2(G543), .ZN(new_n505));
  INV_X1    g080(.A(G50), .ZN(new_n506));
  NOR2_X1   g081(.A1(KEYINPUT5), .A2(G543), .ZN(new_n507));
  AND2_X1   g082(.A1(KEYINPUT5), .A2(G543), .ZN(new_n508));
  AND2_X1   g083(.A1(KEYINPUT6), .A2(G651), .ZN(new_n509));
  NOR2_X1   g084(.A1(KEYINPUT6), .A2(G651), .ZN(new_n510));
  OAI22_X1  g085(.A1(new_n507), .A2(new_n508), .B1(new_n509), .B2(new_n510), .ZN(new_n511));
  XOR2_X1   g086(.A(KEYINPUT69), .B(G88), .Z(new_n512));
  OAI22_X1  g087(.A1(new_n505), .A2(new_n506), .B1(new_n511), .B2(new_n512), .ZN(new_n513));
  OR2_X1    g088(.A1(new_n501), .A2(new_n513), .ZN(G303));
  INV_X1    g089(.A(G303), .ZN(G166));
  NAND3_X1  g090(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n516));
  XNOR2_X1  g091(.A(new_n516), .B(KEYINPUT7), .ZN(new_n517));
  XOR2_X1   g092(.A(KEYINPUT70), .B(G51), .Z(new_n518));
  OAI21_X1  g093(.A(new_n517), .B1(new_n505), .B2(new_n518), .ZN(new_n519));
  NOR2_X1   g094(.A1(new_n508), .A2(new_n507), .ZN(new_n520));
  NAND2_X1  g095(.A1(new_n504), .A2(G89), .ZN(new_n521));
  NAND2_X1  g096(.A1(G63), .A2(G651), .ZN(new_n522));
  AOI21_X1  g097(.A(new_n520), .B1(new_n521), .B2(new_n522), .ZN(new_n523));
  NOR2_X1   g098(.A1(new_n519), .A2(new_n523), .ZN(G168));
  AOI22_X1  g099(.A1(new_n498), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n525));
  NOR2_X1   g100(.A1(new_n525), .A2(new_n500), .ZN(new_n526));
  INV_X1    g101(.A(G52), .ZN(new_n527));
  INV_X1    g102(.A(G90), .ZN(new_n528));
  OAI22_X1  g103(.A1(new_n505), .A2(new_n527), .B1(new_n511), .B2(new_n528), .ZN(new_n529));
  NOR2_X1   g104(.A1(new_n526), .A2(new_n529), .ZN(G171));
  NAND2_X1  g105(.A1(G68), .A2(G543), .ZN(new_n531));
  INV_X1    g106(.A(G56), .ZN(new_n532));
  OAI21_X1  g107(.A(new_n531), .B1(new_n520), .B2(new_n532), .ZN(new_n533));
  AOI21_X1  g108(.A(KEYINPUT71), .B1(new_n533), .B2(G651), .ZN(new_n534));
  INV_X1    g109(.A(G43), .ZN(new_n535));
  INV_X1    g110(.A(G81), .ZN(new_n536));
  OAI22_X1  g111(.A1(new_n505), .A2(new_n535), .B1(new_n511), .B2(new_n536), .ZN(new_n537));
  NOR2_X1   g112(.A1(new_n534), .A2(new_n537), .ZN(new_n538));
  NAND3_X1  g113(.A1(new_n533), .A2(KEYINPUT71), .A3(G651), .ZN(new_n539));
  NAND2_X1  g114(.A1(new_n538), .A2(new_n539), .ZN(new_n540));
  INV_X1    g115(.A(new_n540), .ZN(new_n541));
  NAND2_X1  g116(.A1(new_n541), .A2(G860), .ZN(new_n542));
  XNOR2_X1  g117(.A(new_n542), .B(KEYINPUT72), .ZN(G153));
  NAND4_X1  g118(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g119(.A1(G1), .A2(G3), .ZN(new_n545));
  XNOR2_X1  g120(.A(new_n545), .B(KEYINPUT8), .ZN(new_n546));
  NAND4_X1  g121(.A1(G319), .A2(G483), .A3(G661), .A4(new_n546), .ZN(G188));
  INV_X1    g122(.A(KEYINPUT73), .ZN(new_n548));
  NAND2_X1  g123(.A1(new_n511), .A2(new_n548), .ZN(new_n549));
  NAND3_X1  g124(.A1(new_n504), .A2(new_n498), .A3(KEYINPUT73), .ZN(new_n550));
  NAND3_X1  g125(.A1(new_n549), .A2(G91), .A3(new_n550), .ZN(new_n551));
  INV_X1    g126(.A(G543), .ZN(new_n552));
  AOI21_X1  g127(.A(new_n552), .B1(new_n502), .B2(new_n503), .ZN(new_n553));
  INV_X1    g128(.A(KEYINPUT9), .ZN(new_n554));
  NAND3_X1  g129(.A1(new_n553), .A2(new_n554), .A3(G53), .ZN(new_n555));
  OAI211_X1 g130(.A(G53), .B(G543), .C1(new_n509), .C2(new_n510), .ZN(new_n556));
  NAND2_X1  g131(.A1(new_n556), .A2(KEYINPUT9), .ZN(new_n557));
  NAND2_X1  g132(.A1(new_n555), .A2(new_n557), .ZN(new_n558));
  NAND2_X1  g133(.A1(G78), .A2(G543), .ZN(new_n559));
  XNOR2_X1  g134(.A(KEYINPUT74), .B(G65), .ZN(new_n560));
  OAI21_X1  g135(.A(new_n559), .B1(new_n520), .B2(new_n560), .ZN(new_n561));
  NAND2_X1  g136(.A1(new_n561), .A2(G651), .ZN(new_n562));
  NAND3_X1  g137(.A1(new_n551), .A2(new_n558), .A3(new_n562), .ZN(G299));
  INV_X1    g138(.A(G171), .ZN(G301));
  INV_X1    g139(.A(G168), .ZN(G286));
  NAND3_X1  g140(.A1(new_n549), .A2(G87), .A3(new_n550), .ZN(new_n566));
  INV_X1    g141(.A(G74), .ZN(new_n567));
  NAND2_X1  g142(.A1(new_n520), .A2(new_n567), .ZN(new_n568));
  AOI22_X1  g143(.A1(new_n568), .A2(G651), .B1(new_n553), .B2(G49), .ZN(new_n569));
  NAND2_X1  g144(.A1(new_n566), .A2(new_n569), .ZN(G288));
  NAND3_X1  g145(.A1(new_n549), .A2(G86), .A3(new_n550), .ZN(new_n571));
  OAI21_X1  g146(.A(G61), .B1(new_n508), .B2(new_n507), .ZN(new_n572));
  NAND2_X1  g147(.A1(G73), .A2(G543), .ZN(new_n573));
  NAND2_X1  g148(.A1(new_n572), .A2(new_n573), .ZN(new_n574));
  AOI22_X1  g149(.A1(new_n574), .A2(G651), .B1(G48), .B2(new_n553), .ZN(new_n575));
  NAND2_X1  g150(.A1(new_n571), .A2(new_n575), .ZN(G305));
  AOI22_X1  g151(.A1(new_n498), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n577));
  NOR2_X1   g152(.A1(new_n577), .A2(new_n500), .ZN(new_n578));
  INV_X1    g153(.A(G47), .ZN(new_n579));
  INV_X1    g154(.A(G85), .ZN(new_n580));
  OAI22_X1  g155(.A1(new_n505), .A2(new_n579), .B1(new_n511), .B2(new_n580), .ZN(new_n581));
  INV_X1    g156(.A(KEYINPUT75), .ZN(new_n582));
  OR3_X1    g157(.A1(new_n578), .A2(new_n581), .A3(new_n582), .ZN(new_n583));
  OAI21_X1  g158(.A(new_n582), .B1(new_n578), .B2(new_n581), .ZN(new_n584));
  NAND2_X1  g159(.A1(new_n583), .A2(new_n584), .ZN(G290));
  INV_X1    g160(.A(G868), .ZN(new_n586));
  NOR2_X1   g161(.A1(G171), .A2(new_n586), .ZN(new_n587));
  XNOR2_X1  g162(.A(new_n587), .B(KEYINPUT76), .ZN(new_n588));
  NAND2_X1  g163(.A1(G79), .A2(G543), .ZN(new_n589));
  INV_X1    g164(.A(G66), .ZN(new_n590));
  OAI21_X1  g165(.A(new_n589), .B1(new_n520), .B2(new_n590), .ZN(new_n591));
  AOI22_X1  g166(.A1(new_n591), .A2(G651), .B1(G54), .B2(new_n553), .ZN(new_n592));
  INV_X1    g167(.A(new_n592), .ZN(new_n593));
  NAND3_X1  g168(.A1(new_n549), .A2(G92), .A3(new_n550), .ZN(new_n594));
  INV_X1    g169(.A(KEYINPUT10), .ZN(new_n595));
  OR2_X1    g170(.A1(new_n594), .A2(new_n595), .ZN(new_n596));
  NAND2_X1  g171(.A1(new_n594), .A2(new_n595), .ZN(new_n597));
  AOI21_X1  g172(.A(new_n593), .B1(new_n596), .B2(new_n597), .ZN(new_n598));
  OAI21_X1  g173(.A(new_n588), .B1(G868), .B2(new_n598), .ZN(G284));
  OAI21_X1  g174(.A(new_n588), .B1(G868), .B2(new_n598), .ZN(G321));
  NAND2_X1  g175(.A1(G299), .A2(new_n586), .ZN(new_n601));
  OAI21_X1  g176(.A(new_n601), .B1(new_n586), .B2(G168), .ZN(G297));
  OAI21_X1  g177(.A(new_n601), .B1(new_n586), .B2(G168), .ZN(G280));
  INV_X1    g178(.A(G559), .ZN(new_n604));
  OAI21_X1  g179(.A(new_n598), .B1(new_n604), .B2(G860), .ZN(G148));
  NAND2_X1  g180(.A1(new_n540), .A2(new_n586), .ZN(new_n606));
  NAND2_X1  g181(.A1(new_n596), .A2(new_n597), .ZN(new_n607));
  NAND2_X1  g182(.A1(new_n607), .A2(new_n592), .ZN(new_n608));
  NOR2_X1   g183(.A1(new_n608), .A2(G559), .ZN(new_n609));
  OAI21_X1  g184(.A(new_n606), .B1(new_n609), .B2(new_n586), .ZN(G323));
  XNOR2_X1  g185(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g186(.A1(new_n489), .A2(new_n475), .ZN(new_n612));
  XNOR2_X1  g187(.A(new_n612), .B(KEYINPUT12), .ZN(new_n613));
  XNOR2_X1  g188(.A(new_n613), .B(KEYINPUT13), .ZN(new_n614));
  XNOR2_X1  g189(.A(new_n614), .B(G2100), .ZN(new_n615));
  AND2_X1   g190(.A1(new_n484), .A2(G135), .ZN(new_n616));
  INV_X1    g191(.A(G123), .ZN(new_n617));
  NOR2_X1   g192(.A1(new_n466), .A2(G111), .ZN(new_n618));
  OAI21_X1  g193(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n619));
  OAI22_X1  g194(.A1(new_n479), .A2(new_n617), .B1(new_n618), .B2(new_n619), .ZN(new_n620));
  NOR2_X1   g195(.A1(new_n616), .A2(new_n620), .ZN(new_n621));
  INV_X1    g196(.A(new_n621), .ZN(new_n622));
  OR2_X1    g197(.A1(new_n622), .A2(G2096), .ZN(new_n623));
  NAND2_X1  g198(.A1(new_n622), .A2(G2096), .ZN(new_n624));
  NAND3_X1  g199(.A1(new_n615), .A2(new_n623), .A3(new_n624), .ZN(G156));
  XNOR2_X1  g200(.A(KEYINPUT15), .B(G2435), .ZN(new_n626));
  XNOR2_X1  g201(.A(new_n626), .B(G2438), .ZN(new_n627));
  XNOR2_X1  g202(.A(G2427), .B(G2430), .ZN(new_n628));
  NAND2_X1  g203(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  NAND2_X1  g204(.A1(new_n629), .A2(KEYINPUT14), .ZN(new_n630));
  AND2_X1   g205(.A1(new_n630), .A2(KEYINPUT77), .ZN(new_n631));
  NOR2_X1   g206(.A1(new_n630), .A2(KEYINPUT77), .ZN(new_n632));
  OAI22_X1  g207(.A1(new_n631), .A2(new_n632), .B1(new_n627), .B2(new_n628), .ZN(new_n633));
  XOR2_X1   g208(.A(G2443), .B(G2446), .Z(new_n634));
  XNOR2_X1  g209(.A(new_n633), .B(new_n634), .ZN(new_n635));
  XNOR2_X1  g210(.A(G2451), .B(G2454), .ZN(new_n636));
  XNOR2_X1  g211(.A(new_n636), .B(KEYINPUT16), .ZN(new_n637));
  XNOR2_X1  g212(.A(new_n635), .B(new_n637), .ZN(new_n638));
  XOR2_X1   g213(.A(G1341), .B(G1348), .Z(new_n639));
  OAI21_X1  g214(.A(G14), .B1(new_n638), .B2(new_n639), .ZN(new_n640));
  NAND2_X1  g215(.A1(new_n638), .A2(new_n639), .ZN(new_n641));
  INV_X1    g216(.A(KEYINPUT78), .ZN(new_n642));
  NAND2_X1  g217(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  NAND3_X1  g218(.A1(new_n638), .A2(KEYINPUT78), .A3(new_n639), .ZN(new_n644));
  AOI21_X1  g219(.A(new_n640), .B1(new_n643), .B2(new_n644), .ZN(G401));
  XOR2_X1   g220(.A(G2072), .B(G2078), .Z(new_n646));
  INV_X1    g221(.A(new_n646), .ZN(new_n647));
  XNOR2_X1  g222(.A(G2067), .B(G2678), .ZN(new_n648));
  XOR2_X1   g223(.A(G2084), .B(G2090), .Z(new_n649));
  NAND3_X1  g224(.A1(new_n647), .A2(new_n648), .A3(new_n649), .ZN(new_n650));
  XNOR2_X1  g225(.A(new_n650), .B(KEYINPUT18), .ZN(new_n651));
  XNOR2_X1  g226(.A(KEYINPUT79), .B(KEYINPUT17), .ZN(new_n652));
  XNOR2_X1  g227(.A(new_n646), .B(new_n652), .ZN(new_n653));
  INV_X1    g228(.A(new_n649), .ZN(new_n654));
  NOR3_X1   g229(.A1(new_n653), .A2(new_n648), .A3(new_n654), .ZN(new_n655));
  OAI21_X1  g230(.A(new_n654), .B1(new_n647), .B2(new_n648), .ZN(new_n656));
  AOI21_X1  g231(.A(new_n656), .B1(new_n653), .B2(new_n648), .ZN(new_n657));
  NOR3_X1   g232(.A1(new_n651), .A2(new_n655), .A3(new_n657), .ZN(new_n658));
  XNOR2_X1  g233(.A(G2096), .B(G2100), .ZN(new_n659));
  XNOR2_X1  g234(.A(new_n658), .B(new_n659), .ZN(G227));
  XOR2_X1   g235(.A(G1971), .B(G1976), .Z(new_n661));
  XNOR2_X1  g236(.A(new_n661), .B(KEYINPUT19), .ZN(new_n662));
  XOR2_X1   g237(.A(G1956), .B(G2474), .Z(new_n663));
  XOR2_X1   g238(.A(G1961), .B(G1966), .Z(new_n664));
  AND2_X1   g239(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  NAND2_X1  g240(.A1(new_n662), .A2(new_n665), .ZN(new_n666));
  INV_X1    g241(.A(KEYINPUT20), .ZN(new_n667));
  XNOR2_X1  g242(.A(new_n666), .B(new_n667), .ZN(new_n668));
  NOR2_X1   g243(.A1(new_n663), .A2(new_n664), .ZN(new_n669));
  NOR2_X1   g244(.A1(new_n665), .A2(new_n669), .ZN(new_n670));
  MUX2_X1   g245(.A(new_n670), .B(new_n669), .S(new_n662), .Z(new_n671));
  NOR2_X1   g246(.A1(new_n668), .A2(new_n671), .ZN(new_n672));
  XNOR2_X1  g247(.A(new_n672), .B(G1981), .ZN(new_n673));
  XNOR2_X1  g248(.A(new_n673), .B(G1986), .ZN(new_n674));
  XNOR2_X1  g249(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n675));
  XNOR2_X1  g250(.A(new_n675), .B(KEYINPUT80), .ZN(new_n676));
  NAND2_X1  g251(.A1(new_n674), .A2(new_n676), .ZN(new_n677));
  INV_X1    g252(.A(G1986), .ZN(new_n678));
  XNOR2_X1  g253(.A(new_n673), .B(new_n678), .ZN(new_n679));
  INV_X1    g254(.A(new_n676), .ZN(new_n680));
  NAND2_X1  g255(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  NAND2_X1  g256(.A1(new_n677), .A2(new_n681), .ZN(new_n682));
  XNOR2_X1  g257(.A(G1991), .B(G1996), .ZN(new_n683));
  INV_X1    g258(.A(new_n683), .ZN(new_n684));
  NAND2_X1  g259(.A1(new_n682), .A2(new_n684), .ZN(new_n685));
  NAND3_X1  g260(.A1(new_n677), .A2(new_n681), .A3(new_n683), .ZN(new_n686));
  NAND2_X1  g261(.A1(new_n685), .A2(new_n686), .ZN(G229));
  INV_X1    g262(.A(G16), .ZN(new_n688));
  NOR2_X1   g263(.A1(G171), .A2(new_n688), .ZN(new_n689));
  AOI21_X1  g264(.A(new_n689), .B1(G5), .B2(new_n688), .ZN(new_n690));
  INV_X1    g265(.A(G1961), .ZN(new_n691));
  INV_X1    g266(.A(G2084), .ZN(new_n692));
  INV_X1    g267(.A(G29), .ZN(new_n693));
  INV_X1    g268(.A(KEYINPUT24), .ZN(new_n694));
  OAI21_X1  g269(.A(new_n693), .B1(new_n694), .B2(G34), .ZN(new_n695));
  OR2_X1    g270(.A1(new_n695), .A2(KEYINPUT89), .ZN(new_n696));
  NAND2_X1  g271(.A1(new_n695), .A2(KEYINPUT89), .ZN(new_n697));
  NAND2_X1  g272(.A1(new_n694), .A2(G34), .ZN(new_n698));
  NAND3_X1  g273(.A1(new_n696), .A2(new_n697), .A3(new_n698), .ZN(new_n699));
  INV_X1    g274(.A(G160), .ZN(new_n700));
  OAI21_X1  g275(.A(new_n699), .B1(new_n700), .B2(new_n693), .ZN(new_n701));
  OAI22_X1  g276(.A1(new_n690), .A2(new_n691), .B1(new_n692), .B2(new_n701), .ZN(new_n702));
  OAI21_X1  g277(.A(KEYINPUT91), .B1(G16), .B2(G21), .ZN(new_n703));
  NAND2_X1  g278(.A1(G168), .A2(G16), .ZN(new_n704));
  MUX2_X1   g279(.A(KEYINPUT91), .B(new_n703), .S(new_n704), .Z(new_n705));
  XOR2_X1   g280(.A(KEYINPUT92), .B(G1966), .Z(new_n706));
  XNOR2_X1  g281(.A(new_n705), .B(new_n706), .ZN(new_n707));
  NOR2_X1   g282(.A1(G4), .A2(G16), .ZN(new_n708));
  AOI21_X1  g283(.A(new_n708), .B1(new_n598), .B2(G16), .ZN(new_n709));
  AOI211_X1 g284(.A(new_n702), .B(new_n707), .C1(G1348), .C2(new_n709), .ZN(new_n710));
  NAND2_X1  g285(.A1(new_n693), .A2(G27), .ZN(new_n711));
  XNOR2_X1  g286(.A(new_n711), .B(KEYINPUT96), .ZN(new_n712));
  OAI21_X1  g287(.A(new_n712), .B1(G164), .B2(new_n693), .ZN(new_n713));
  XOR2_X1   g288(.A(KEYINPUT97), .B(G2078), .Z(new_n714));
  XNOR2_X1  g289(.A(new_n713), .B(new_n714), .ZN(new_n715));
  NAND2_X1  g290(.A1(new_n688), .A2(G19), .ZN(new_n716));
  OAI21_X1  g291(.A(new_n716), .B1(new_n541), .B2(new_n688), .ZN(new_n717));
  XOR2_X1   g292(.A(new_n717), .B(G1341), .Z(new_n718));
  NAND3_X1  g293(.A1(new_n710), .A2(new_n715), .A3(new_n718), .ZN(new_n719));
  AOI22_X1  g294(.A1(new_n690), .A2(new_n691), .B1(new_n692), .B2(new_n701), .ZN(new_n720));
  INV_X1    g295(.A(KEYINPUT90), .ZN(new_n721));
  OAI21_X1  g296(.A(new_n721), .B1(G29), .B2(G32), .ZN(new_n722));
  NAND3_X1  g297(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n723));
  INV_X1    g298(.A(KEYINPUT26), .ZN(new_n724));
  OR2_X1    g299(.A1(new_n723), .A2(new_n724), .ZN(new_n725));
  NAND2_X1  g300(.A1(new_n723), .A2(new_n724), .ZN(new_n726));
  AOI22_X1  g301(.A1(new_n725), .A2(new_n726), .B1(G105), .B2(new_n475), .ZN(new_n727));
  INV_X1    g302(.A(G129), .ZN(new_n728));
  OAI21_X1  g303(.A(new_n727), .B1(new_n479), .B2(new_n728), .ZN(new_n729));
  AND2_X1   g304(.A1(new_n484), .A2(G141), .ZN(new_n730));
  NOR2_X1   g305(.A1(new_n729), .A2(new_n730), .ZN(new_n731));
  NAND2_X1  g306(.A1(new_n731), .A2(G29), .ZN(new_n732));
  MUX2_X1   g307(.A(new_n721), .B(new_n722), .S(new_n732), .Z(new_n733));
  XNOR2_X1  g308(.A(KEYINPUT27), .B(G1996), .ZN(new_n734));
  OAI21_X1  g309(.A(new_n720), .B1(new_n733), .B2(new_n734), .ZN(new_n735));
  INV_X1    g310(.A(KEYINPUT95), .ZN(new_n736));
  OR2_X1    g311(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  NAND2_X1  g312(.A1(new_n735), .A2(new_n736), .ZN(new_n738));
  NAND2_X1  g313(.A1(new_n693), .A2(G35), .ZN(new_n739));
  OAI21_X1  g314(.A(new_n739), .B1(G162), .B2(new_n693), .ZN(new_n740));
  XNOR2_X1  g315(.A(new_n740), .B(KEYINPUT29), .ZN(new_n741));
  NOR2_X1   g316(.A1(new_n741), .A2(G2090), .ZN(new_n742));
  OAI211_X1 g317(.A(new_n737), .B(new_n738), .C1(KEYINPUT98), .C2(new_n742), .ZN(new_n743));
  NAND2_X1  g318(.A1(new_n733), .A2(new_n734), .ZN(new_n744));
  XOR2_X1   g319(.A(KEYINPUT31), .B(G11), .Z(new_n745));
  INV_X1    g320(.A(KEYINPUT30), .ZN(new_n746));
  OAI21_X1  g321(.A(new_n693), .B1(new_n746), .B2(G28), .ZN(new_n747));
  INV_X1    g322(.A(new_n747), .ZN(new_n748));
  OR2_X1    g323(.A1(new_n748), .A2(KEYINPUT93), .ZN(new_n749));
  AOI22_X1  g324(.A1(new_n748), .A2(KEYINPUT93), .B1(new_n746), .B2(G28), .ZN(new_n750));
  AOI21_X1  g325(.A(new_n745), .B1(new_n749), .B2(new_n750), .ZN(new_n751));
  OAI21_X1  g326(.A(new_n751), .B1(new_n622), .B2(new_n693), .ZN(new_n752));
  XOR2_X1   g327(.A(new_n752), .B(KEYINPUT94), .Z(new_n753));
  OAI211_X1 g328(.A(new_n744), .B(new_n753), .C1(G1348), .C2(new_n709), .ZN(new_n754));
  NAND2_X1  g329(.A1(new_n693), .A2(G26), .ZN(new_n755));
  XOR2_X1   g330(.A(new_n755), .B(KEYINPUT28), .Z(new_n756));
  OR2_X1    g331(.A1(G104), .A2(G2105), .ZN(new_n757));
  OAI211_X1 g332(.A(new_n757), .B(G2104), .C1(G116), .C2(new_n466), .ZN(new_n758));
  INV_X1    g333(.A(G128), .ZN(new_n759));
  OAI21_X1  g334(.A(new_n758), .B1(new_n479), .B2(new_n759), .ZN(new_n760));
  AOI21_X1  g335(.A(new_n760), .B1(new_n484), .B2(G140), .ZN(new_n761));
  XOR2_X1   g336(.A(new_n761), .B(KEYINPUT84), .Z(new_n762));
  AOI21_X1  g337(.A(new_n756), .B1(new_n762), .B2(G29), .ZN(new_n763));
  XNOR2_X1  g338(.A(new_n763), .B(G2067), .ZN(new_n764));
  NAND2_X1  g339(.A1(new_n742), .A2(KEYINPUT98), .ZN(new_n765));
  NAND2_X1  g340(.A1(new_n764), .A2(new_n765), .ZN(new_n766));
  NOR4_X1   g341(.A1(new_n719), .A2(new_n743), .A3(new_n754), .A4(new_n766), .ZN(new_n767));
  NAND2_X1  g342(.A1(G299), .A2(G16), .ZN(new_n768));
  NAND2_X1  g343(.A1(new_n688), .A2(G20), .ZN(new_n769));
  XNOR2_X1  g344(.A(new_n769), .B(KEYINPUT99), .ZN(new_n770));
  XNOR2_X1  g345(.A(new_n770), .B(KEYINPUT23), .ZN(new_n771));
  NAND2_X1  g346(.A1(new_n768), .A2(new_n771), .ZN(new_n772));
  XNOR2_X1  g347(.A(new_n772), .B(KEYINPUT100), .ZN(new_n773));
  INV_X1    g348(.A(G1956), .ZN(new_n774));
  XNOR2_X1  g349(.A(new_n773), .B(new_n774), .ZN(new_n775));
  NAND2_X1  g350(.A1(new_n693), .A2(G33), .ZN(new_n776));
  NAND3_X1  g351(.A1(new_n466), .A2(G103), .A3(G2104), .ZN(new_n777));
  INV_X1    g352(.A(KEYINPUT86), .ZN(new_n778));
  XNOR2_X1  g353(.A(new_n777), .B(new_n778), .ZN(new_n779));
  OR2_X1    g354(.A1(new_n779), .A2(KEYINPUT85), .ZN(new_n780));
  NAND2_X1  g355(.A1(new_n779), .A2(KEYINPUT85), .ZN(new_n781));
  NAND2_X1  g356(.A1(new_n780), .A2(new_n781), .ZN(new_n782));
  INV_X1    g357(.A(KEYINPUT25), .ZN(new_n783));
  NAND2_X1  g358(.A1(new_n782), .A2(new_n783), .ZN(new_n784));
  INV_X1    g359(.A(G139), .ZN(new_n785));
  NOR2_X1   g360(.A1(new_n468), .A2(new_n785), .ZN(new_n786));
  XNOR2_X1  g361(.A(new_n786), .B(KEYINPUT87), .ZN(new_n787));
  NAND3_X1  g362(.A1(new_n780), .A2(KEYINPUT25), .A3(new_n781), .ZN(new_n788));
  NAND3_X1  g363(.A1(new_n784), .A2(new_n787), .A3(new_n788), .ZN(new_n789));
  INV_X1    g364(.A(KEYINPUT88), .ZN(new_n790));
  XNOR2_X1  g365(.A(new_n789), .B(new_n790), .ZN(new_n791));
  AOI22_X1  g366(.A1(new_n489), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n792));
  OR2_X1    g367(.A1(new_n792), .A2(new_n466), .ZN(new_n793));
  NAND2_X1  g368(.A1(new_n791), .A2(new_n793), .ZN(new_n794));
  INV_X1    g369(.A(new_n794), .ZN(new_n795));
  OAI21_X1  g370(.A(new_n776), .B1(new_n795), .B2(new_n693), .ZN(new_n796));
  AND2_X1   g371(.A1(new_n796), .A2(G2072), .ZN(new_n797));
  AOI211_X1 g372(.A(new_n775), .B(new_n797), .C1(G2090), .C2(new_n741), .ZN(new_n798));
  OAI211_X1 g373(.A(new_n767), .B(new_n798), .C1(G2072), .C2(new_n796), .ZN(new_n799));
  NAND2_X1  g374(.A1(new_n688), .A2(G22), .ZN(new_n800));
  OAI21_X1  g375(.A(new_n800), .B1(G166), .B2(new_n688), .ZN(new_n801));
  INV_X1    g376(.A(G1971), .ZN(new_n802));
  XNOR2_X1  g377(.A(new_n801), .B(new_n802), .ZN(new_n803));
  AND2_X1   g378(.A1(new_n688), .A2(G6), .ZN(new_n804));
  AOI21_X1  g379(.A(new_n804), .B1(G305), .B2(G16), .ZN(new_n805));
  XOR2_X1   g380(.A(KEYINPUT32), .B(G1981), .Z(new_n806));
  OR2_X1    g381(.A1(new_n805), .A2(new_n806), .ZN(new_n807));
  NOR2_X1   g382(.A1(G16), .A2(G23), .ZN(new_n808));
  XNOR2_X1  g383(.A(new_n808), .B(KEYINPUT83), .ZN(new_n809));
  OAI21_X1  g384(.A(new_n809), .B1(G288), .B2(new_n688), .ZN(new_n810));
  XNOR2_X1  g385(.A(KEYINPUT33), .B(G1976), .ZN(new_n811));
  OR2_X1    g386(.A1(new_n810), .A2(new_n811), .ZN(new_n812));
  AOI22_X1  g387(.A1(new_n806), .A2(new_n805), .B1(new_n810), .B2(new_n811), .ZN(new_n813));
  NAND4_X1  g388(.A1(new_n803), .A2(new_n807), .A3(new_n812), .A4(new_n813), .ZN(new_n814));
  OR2_X1    g389(.A1(new_n814), .A2(KEYINPUT34), .ZN(new_n815));
  NAND2_X1  g390(.A1(new_n814), .A2(KEYINPUT34), .ZN(new_n816));
  NAND2_X1  g391(.A1(new_n688), .A2(G24), .ZN(new_n817));
  INV_X1    g392(.A(G290), .ZN(new_n818));
  OAI21_X1  g393(.A(new_n817), .B1(new_n818), .B2(new_n688), .ZN(new_n819));
  XOR2_X1   g394(.A(KEYINPUT82), .B(G1986), .Z(new_n820));
  XNOR2_X1  g395(.A(new_n819), .B(new_n820), .ZN(new_n821));
  NAND2_X1  g396(.A1(new_n693), .A2(G25), .ZN(new_n822));
  INV_X1    g397(.A(G119), .ZN(new_n823));
  NOR2_X1   g398(.A1(new_n479), .A2(new_n823), .ZN(new_n824));
  INV_X1    g399(.A(KEYINPUT81), .ZN(new_n825));
  XNOR2_X1  g400(.A(new_n824), .B(new_n825), .ZN(new_n826));
  OAI21_X1  g401(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n827));
  INV_X1    g402(.A(G107), .ZN(new_n828));
  AOI21_X1  g403(.A(new_n827), .B1(new_n828), .B2(G2105), .ZN(new_n829));
  AOI21_X1  g404(.A(new_n829), .B1(new_n484), .B2(G131), .ZN(new_n830));
  NAND2_X1  g405(.A1(new_n826), .A2(new_n830), .ZN(new_n831));
  INV_X1    g406(.A(new_n831), .ZN(new_n832));
  OAI21_X1  g407(.A(new_n822), .B1(new_n832), .B2(new_n693), .ZN(new_n833));
  XOR2_X1   g408(.A(KEYINPUT35), .B(G1991), .Z(new_n834));
  XNOR2_X1  g409(.A(new_n833), .B(new_n834), .ZN(new_n835));
  NAND4_X1  g410(.A1(new_n815), .A2(new_n816), .A3(new_n821), .A4(new_n835), .ZN(new_n836));
  XOR2_X1   g411(.A(new_n836), .B(KEYINPUT36), .Z(new_n837));
  NOR2_X1   g412(.A1(new_n799), .A2(new_n837), .ZN(G311));
  INV_X1    g413(.A(G311), .ZN(G150));
  NAND2_X1  g414(.A1(new_n598), .A2(G559), .ZN(new_n840));
  XOR2_X1   g415(.A(new_n840), .B(KEYINPUT38), .Z(new_n841));
  NAND2_X1  g416(.A1(G80), .A2(G543), .ZN(new_n842));
  INV_X1    g417(.A(G67), .ZN(new_n843));
  OAI21_X1  g418(.A(new_n842), .B1(new_n520), .B2(new_n843), .ZN(new_n844));
  AOI21_X1  g419(.A(new_n500), .B1(new_n844), .B2(KEYINPUT101), .ZN(new_n845));
  OAI21_X1  g420(.A(new_n845), .B1(KEYINPUT101), .B2(new_n844), .ZN(new_n846));
  INV_X1    g421(.A(new_n511), .ZN(new_n847));
  AOI22_X1  g422(.A1(new_n847), .A2(G93), .B1(G55), .B2(new_n553), .ZN(new_n848));
  NAND2_X1  g423(.A1(new_n846), .A2(new_n848), .ZN(new_n849));
  OR2_X1    g424(.A1(new_n849), .A2(new_n540), .ZN(new_n850));
  NAND2_X1  g425(.A1(new_n849), .A2(new_n540), .ZN(new_n851));
  NAND2_X1  g426(.A1(new_n850), .A2(new_n851), .ZN(new_n852));
  XNOR2_X1  g427(.A(new_n841), .B(new_n852), .ZN(new_n853));
  AND2_X1   g428(.A1(new_n853), .A2(KEYINPUT39), .ZN(new_n854));
  NOR2_X1   g429(.A1(new_n853), .A2(KEYINPUT39), .ZN(new_n855));
  NOR3_X1   g430(.A1(new_n854), .A2(new_n855), .A3(G860), .ZN(new_n856));
  NAND2_X1  g431(.A1(new_n849), .A2(G860), .ZN(new_n857));
  XNOR2_X1  g432(.A(new_n857), .B(KEYINPUT37), .ZN(new_n858));
  OR2_X1    g433(.A1(new_n856), .A2(new_n858), .ZN(G145));
  XNOR2_X1  g434(.A(new_n831), .B(KEYINPUT102), .ZN(new_n860));
  XNOR2_X1  g435(.A(new_n860), .B(new_n613), .ZN(new_n861));
  INV_X1    g436(.A(G130), .ZN(new_n862));
  NOR2_X1   g437(.A1(new_n466), .A2(G118), .ZN(new_n863));
  OAI21_X1  g438(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n864));
  OAI22_X1  g439(.A1(new_n479), .A2(new_n862), .B1(new_n863), .B2(new_n864), .ZN(new_n865));
  AOI21_X1  g440(.A(new_n865), .B1(new_n484), .B2(G142), .ZN(new_n866));
  XNOR2_X1  g441(.A(new_n861), .B(new_n866), .ZN(new_n867));
  INV_X1    g442(.A(new_n867), .ZN(new_n868));
  XNOR2_X1  g443(.A(new_n762), .B(G164), .ZN(new_n869));
  NOR2_X1   g444(.A1(new_n794), .A2(new_n869), .ZN(new_n870));
  INV_X1    g445(.A(new_n870), .ZN(new_n871));
  NAND2_X1  g446(.A1(new_n794), .A2(new_n869), .ZN(new_n872));
  AOI21_X1  g447(.A(new_n731), .B1(new_n871), .B2(new_n872), .ZN(new_n873));
  INV_X1    g448(.A(new_n872), .ZN(new_n874));
  INV_X1    g449(.A(new_n731), .ZN(new_n875));
  NOR3_X1   g450(.A1(new_n874), .A2(new_n875), .A3(new_n870), .ZN(new_n876));
  OAI22_X1  g451(.A1(new_n868), .A2(KEYINPUT103), .B1(new_n873), .B2(new_n876), .ZN(new_n877));
  XNOR2_X1  g452(.A(new_n700), .B(new_n621), .ZN(new_n878));
  XNOR2_X1  g453(.A(new_n878), .B(G162), .ZN(new_n879));
  INV_X1    g454(.A(new_n879), .ZN(new_n880));
  OAI21_X1  g455(.A(new_n875), .B1(new_n874), .B2(new_n870), .ZN(new_n881));
  NAND3_X1  g456(.A1(new_n871), .A2(new_n731), .A3(new_n872), .ZN(new_n882));
  INV_X1    g457(.A(KEYINPUT103), .ZN(new_n883));
  NAND4_X1  g458(.A1(new_n881), .A2(new_n882), .A3(new_n867), .A4(new_n883), .ZN(new_n884));
  NAND3_X1  g459(.A1(new_n877), .A2(new_n880), .A3(new_n884), .ZN(new_n885));
  INV_X1    g460(.A(G37), .ZN(new_n886));
  OAI21_X1  g461(.A(new_n867), .B1(new_n873), .B2(new_n876), .ZN(new_n887));
  NAND3_X1  g462(.A1(new_n868), .A2(new_n882), .A3(new_n881), .ZN(new_n888));
  NAND3_X1  g463(.A1(new_n887), .A2(new_n888), .A3(new_n879), .ZN(new_n889));
  NAND3_X1  g464(.A1(new_n885), .A2(new_n886), .A3(new_n889), .ZN(new_n890));
  XNOR2_X1  g465(.A(new_n890), .B(KEYINPUT40), .ZN(G395));
  XNOR2_X1  g466(.A(new_n852), .B(new_n609), .ZN(new_n892));
  AND2_X1   g467(.A1(new_n608), .A2(G299), .ZN(new_n893));
  NOR2_X1   g468(.A1(new_n608), .A2(G299), .ZN(new_n894));
  NOR2_X1   g469(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  NOR2_X1   g470(.A1(new_n892), .A2(new_n895), .ZN(new_n896));
  NAND2_X1  g471(.A1(new_n895), .A2(KEYINPUT41), .ZN(new_n897));
  INV_X1    g472(.A(KEYINPUT41), .ZN(new_n898));
  OAI21_X1  g473(.A(new_n898), .B1(new_n893), .B2(new_n894), .ZN(new_n899));
  NAND2_X1  g474(.A1(new_n897), .A2(new_n899), .ZN(new_n900));
  AOI21_X1  g475(.A(new_n896), .B1(new_n892), .B2(new_n900), .ZN(new_n901));
  INV_X1    g476(.A(KEYINPUT42), .ZN(new_n902));
  OR2_X1    g477(.A1(new_n901), .A2(new_n902), .ZN(new_n903));
  XNOR2_X1  g478(.A(G290), .B(G305), .ZN(new_n904));
  XOR2_X1   g479(.A(G303), .B(G288), .Z(new_n905));
  XNOR2_X1  g480(.A(new_n904), .B(new_n905), .ZN(new_n906));
  INV_X1    g481(.A(new_n906), .ZN(new_n907));
  NOR2_X1   g482(.A1(new_n907), .A2(KEYINPUT104), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n901), .A2(new_n902), .ZN(new_n909));
  AND3_X1   g484(.A1(new_n903), .A2(new_n908), .A3(new_n909), .ZN(new_n910));
  AOI21_X1  g485(.A(new_n908), .B1(new_n903), .B2(new_n909), .ZN(new_n911));
  OAI21_X1  g486(.A(G868), .B1(new_n910), .B2(new_n911), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n849), .A2(new_n586), .ZN(new_n913));
  NAND2_X1  g488(.A1(new_n912), .A2(new_n913), .ZN(G295));
  NAND2_X1  g489(.A1(new_n912), .A2(new_n913), .ZN(G331));
  INV_X1    g490(.A(KEYINPUT44), .ZN(new_n916));
  XNOR2_X1  g491(.A(KEYINPUT105), .B(KEYINPUT43), .ZN(new_n917));
  XNOR2_X1  g492(.A(G171), .B(KEYINPUT106), .ZN(new_n918));
  NAND3_X1  g493(.A1(new_n850), .A2(new_n851), .A3(new_n918), .ZN(new_n919));
  INV_X1    g494(.A(new_n919), .ZN(new_n920));
  AOI21_X1  g495(.A(new_n918), .B1(new_n850), .B2(new_n851), .ZN(new_n921));
  OAI21_X1  g496(.A(G286), .B1(new_n920), .B2(new_n921), .ZN(new_n922));
  INV_X1    g497(.A(new_n918), .ZN(new_n923));
  NAND2_X1  g498(.A1(new_n852), .A2(new_n923), .ZN(new_n924));
  NAND3_X1  g499(.A1(new_n924), .A2(G168), .A3(new_n919), .ZN(new_n925));
  NAND3_X1  g500(.A1(new_n922), .A2(new_n895), .A3(new_n925), .ZN(new_n926));
  AND2_X1   g501(.A1(new_n922), .A2(new_n925), .ZN(new_n927));
  OAI21_X1  g502(.A(new_n926), .B1(new_n927), .B2(new_n900), .ZN(new_n928));
  NAND2_X1  g503(.A1(new_n928), .A2(KEYINPUT107), .ZN(new_n929));
  INV_X1    g504(.A(KEYINPUT107), .ZN(new_n930));
  OAI211_X1 g505(.A(new_n930), .B(new_n926), .C1(new_n927), .C2(new_n900), .ZN(new_n931));
  NAND3_X1  g506(.A1(new_n929), .A2(new_n906), .A3(new_n931), .ZN(new_n932));
  OAI211_X1 g507(.A(new_n907), .B(new_n926), .C1(new_n927), .C2(new_n900), .ZN(new_n933));
  NAND2_X1  g508(.A1(new_n933), .A2(new_n886), .ZN(new_n934));
  INV_X1    g509(.A(new_n934), .ZN(new_n935));
  AOI21_X1  g510(.A(new_n917), .B1(new_n932), .B2(new_n935), .ZN(new_n936));
  INV_X1    g511(.A(KEYINPUT108), .ZN(new_n937));
  OAI211_X1 g512(.A(new_n937), .B(new_n926), .C1(new_n927), .C2(new_n900), .ZN(new_n938));
  NAND4_X1  g513(.A1(new_n922), .A2(new_n925), .A3(KEYINPUT108), .A4(new_n895), .ZN(new_n939));
  AND2_X1   g514(.A1(new_n939), .A2(new_n906), .ZN(new_n940));
  NAND2_X1  g515(.A1(new_n938), .A2(new_n940), .ZN(new_n941));
  NAND3_X1  g516(.A1(new_n941), .A2(new_n886), .A3(new_n933), .ZN(new_n942));
  INV_X1    g517(.A(new_n917), .ZN(new_n943));
  NOR2_X1   g518(.A1(new_n942), .A2(new_n943), .ZN(new_n944));
  OAI21_X1  g519(.A(new_n916), .B1(new_n936), .B2(new_n944), .ZN(new_n945));
  AOI21_X1  g520(.A(new_n916), .B1(new_n942), .B2(KEYINPUT43), .ZN(new_n946));
  NAND3_X1  g521(.A1(new_n932), .A2(new_n935), .A3(new_n917), .ZN(new_n947));
  AND3_X1   g522(.A1(new_n946), .A2(KEYINPUT109), .A3(new_n947), .ZN(new_n948));
  AOI21_X1  g523(.A(KEYINPUT109), .B1(new_n946), .B2(new_n947), .ZN(new_n949));
  OAI21_X1  g524(.A(new_n945), .B1(new_n948), .B2(new_n949), .ZN(G397));
  INV_X1    g525(.A(G1384), .ZN(new_n951));
  OAI21_X1  g526(.A(new_n951), .B1(new_n491), .B2(new_n495), .ZN(new_n952));
  INV_X1    g527(.A(KEYINPUT45), .ZN(new_n953));
  NAND2_X1  g528(.A1(new_n952), .A2(new_n953), .ZN(new_n954));
  NAND2_X1  g529(.A1(new_n472), .A2(new_n473), .ZN(new_n955));
  NAND2_X1  g530(.A1(new_n955), .A2(G2105), .ZN(new_n956));
  AND2_X1   g531(.A1(new_n465), .A2(new_n467), .ZN(new_n957));
  NAND4_X1  g532(.A1(new_n957), .A2(G137), .A3(new_n466), .A4(new_n463), .ZN(new_n958));
  NAND4_X1  g533(.A1(new_n956), .A2(new_n958), .A3(G40), .A4(new_n476), .ZN(new_n959));
  NOR2_X1   g534(.A1(new_n954), .A2(new_n959), .ZN(new_n960));
  INV_X1    g535(.A(G1996), .ZN(new_n961));
  NAND2_X1  g536(.A1(new_n960), .A2(new_n961), .ZN(new_n962));
  XOR2_X1   g537(.A(new_n962), .B(KEYINPUT110), .Z(new_n963));
  NOR2_X1   g538(.A1(new_n963), .A2(new_n875), .ZN(new_n964));
  INV_X1    g539(.A(new_n960), .ZN(new_n965));
  INV_X1    g540(.A(G2067), .ZN(new_n966));
  XNOR2_X1  g541(.A(new_n762), .B(new_n966), .ZN(new_n967));
  NAND2_X1  g542(.A1(new_n875), .A2(G1996), .ZN(new_n968));
  AOI21_X1  g543(.A(new_n965), .B1(new_n967), .B2(new_n968), .ZN(new_n969));
  NOR2_X1   g544(.A1(new_n964), .A2(new_n969), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n832), .A2(new_n834), .ZN(new_n971));
  INV_X1    g546(.A(new_n971), .ZN(new_n972));
  NOR2_X1   g547(.A1(new_n832), .A2(new_n834), .ZN(new_n973));
  OAI21_X1  g548(.A(new_n960), .B1(new_n972), .B2(new_n973), .ZN(new_n974));
  NAND2_X1  g549(.A1(new_n970), .A2(new_n974), .ZN(new_n975));
  INV_X1    g550(.A(KEYINPUT126), .ZN(new_n976));
  NAND2_X1  g551(.A1(new_n975), .A2(new_n976), .ZN(new_n977));
  NAND2_X1  g552(.A1(new_n818), .A2(new_n678), .ZN(new_n978));
  NOR2_X1   g553(.A1(new_n978), .A2(new_n965), .ZN(new_n979));
  XNOR2_X1  g554(.A(new_n979), .B(KEYINPUT127), .ZN(new_n980));
  XOR2_X1   g555(.A(new_n980), .B(KEYINPUT48), .Z(new_n981));
  NAND3_X1  g556(.A1(new_n970), .A2(KEYINPUT126), .A3(new_n974), .ZN(new_n982));
  NAND3_X1  g557(.A1(new_n977), .A2(new_n981), .A3(new_n982), .ZN(new_n983));
  INV_X1    g558(.A(new_n967), .ZN(new_n984));
  OAI21_X1  g559(.A(new_n960), .B1(new_n984), .B2(new_n875), .ZN(new_n985));
  AND2_X1   g560(.A1(new_n963), .A2(KEYINPUT46), .ZN(new_n986));
  NOR2_X1   g561(.A1(new_n963), .A2(KEYINPUT46), .ZN(new_n987));
  OAI21_X1  g562(.A(new_n985), .B1(new_n986), .B2(new_n987), .ZN(new_n988));
  XNOR2_X1  g563(.A(new_n988), .B(KEYINPUT47), .ZN(new_n989));
  NOR3_X1   g564(.A1(new_n964), .A2(new_n969), .A3(new_n971), .ZN(new_n990));
  NOR2_X1   g565(.A1(new_n762), .A2(G2067), .ZN(new_n991));
  OAI21_X1  g566(.A(new_n960), .B1(new_n990), .B2(new_n991), .ZN(new_n992));
  AND3_X1   g567(.A1(new_n983), .A2(new_n989), .A3(new_n992), .ZN(new_n993));
  NAND2_X1  g568(.A1(G290), .A2(G1986), .ZN(new_n994));
  AOI21_X1  g569(.A(new_n965), .B1(new_n978), .B2(new_n994), .ZN(new_n995));
  NOR2_X1   g570(.A1(new_n975), .A2(new_n995), .ZN(new_n996));
  INV_X1    g571(.A(G8), .ZN(new_n997));
  NOR2_X1   g572(.A1(G168), .A2(new_n997), .ZN(new_n998));
  INV_X1    g573(.A(new_n998), .ZN(new_n999));
  NAND2_X1  g574(.A1(new_n952), .A2(KEYINPUT50), .ZN(new_n1000));
  INV_X1    g575(.A(G40), .ZN(new_n1001));
  NOR4_X1   g576(.A1(new_n470), .A2(new_n474), .A3(new_n1001), .A4(new_n477), .ZN(new_n1002));
  NOR2_X1   g577(.A1(KEYINPUT50), .A2(G1384), .ZN(new_n1003));
  OAI21_X1  g578(.A(new_n1003), .B1(new_n491), .B2(new_n495), .ZN(new_n1004));
  NAND4_X1  g579(.A1(new_n1000), .A2(new_n692), .A3(new_n1002), .A4(new_n1004), .ZN(new_n1005));
  NAND2_X1  g580(.A1(new_n1005), .A2(KEYINPUT118), .ZN(new_n1006));
  AND2_X1   g581(.A1(new_n952), .A2(new_n953), .ZN(new_n1007));
  OAI211_X1 g582(.A(KEYINPUT45), .B(new_n951), .C1(new_n491), .C2(new_n495), .ZN(new_n1008));
  NAND2_X1  g583(.A1(new_n1002), .A2(new_n1008), .ZN(new_n1009));
  OAI21_X1  g584(.A(new_n706), .B1(new_n1007), .B2(new_n1009), .ZN(new_n1010));
  AOI21_X1  g585(.A(new_n959), .B1(new_n496), .B2(new_n1003), .ZN(new_n1011));
  INV_X1    g586(.A(KEYINPUT118), .ZN(new_n1012));
  NAND4_X1  g587(.A1(new_n1011), .A2(new_n1012), .A3(new_n692), .A4(new_n1000), .ZN(new_n1013));
  NAND3_X1  g588(.A1(new_n1006), .A2(new_n1010), .A3(new_n1013), .ZN(new_n1014));
  NAND2_X1  g589(.A1(new_n1014), .A2(KEYINPUT122), .ZN(new_n1015));
  INV_X1    g590(.A(KEYINPUT122), .ZN(new_n1016));
  NAND4_X1  g591(.A1(new_n1006), .A2(new_n1010), .A3(new_n1013), .A4(new_n1016), .ZN(new_n1017));
  AOI21_X1  g592(.A(new_n999), .B1(new_n1015), .B2(new_n1017), .ZN(new_n1018));
  NAND3_X1  g593(.A1(new_n1015), .A2(G168), .A3(new_n1017), .ZN(new_n1019));
  AND2_X1   g594(.A1(KEYINPUT51), .A2(G8), .ZN(new_n1020));
  NAND2_X1  g595(.A1(new_n1019), .A2(new_n1020), .ZN(new_n1021));
  NAND2_X1  g596(.A1(new_n1014), .A2(G8), .ZN(new_n1022));
  NOR2_X1   g597(.A1(new_n998), .A2(KEYINPUT51), .ZN(new_n1023));
  NAND2_X1  g598(.A1(new_n1022), .A2(new_n1023), .ZN(new_n1024));
  AOI21_X1  g599(.A(new_n1018), .B1(new_n1021), .B2(new_n1024), .ZN(new_n1025));
  INV_X1    g600(.A(KEYINPUT62), .ZN(new_n1026));
  OAI21_X1  g601(.A(KEYINPUT124), .B1(new_n1025), .B2(new_n1026), .ZN(new_n1027));
  INV_X1    g602(.A(KEYINPUT117), .ZN(new_n1028));
  AND2_X1   g603(.A1(new_n1002), .A2(new_n1008), .ZN(new_n1029));
  AOI21_X1  g604(.A(G1971), .B1(new_n1029), .B2(new_n954), .ZN(new_n1030));
  INV_X1    g605(.A(G2090), .ZN(new_n1031));
  AND4_X1   g606(.A1(new_n1031), .A2(new_n1000), .A3(new_n1002), .A4(new_n1004), .ZN(new_n1032));
  OAI21_X1  g607(.A(new_n1028), .B1(new_n1030), .B2(new_n1032), .ZN(new_n1033));
  OAI21_X1  g608(.A(new_n802), .B1(new_n1007), .B2(new_n1009), .ZN(new_n1034));
  NAND3_X1  g609(.A1(new_n1011), .A2(new_n1031), .A3(new_n1000), .ZN(new_n1035));
  NAND3_X1  g610(.A1(new_n1034), .A2(new_n1035), .A3(KEYINPUT117), .ZN(new_n1036));
  NAND3_X1  g611(.A1(new_n1033), .A2(G8), .A3(new_n1036), .ZN(new_n1037));
  NAND2_X1  g612(.A1(G303), .A2(G8), .ZN(new_n1038));
  XNOR2_X1  g613(.A(new_n1038), .B(KEYINPUT55), .ZN(new_n1039));
  NAND2_X1  g614(.A1(new_n1037), .A2(new_n1039), .ZN(new_n1040));
  AND2_X1   g615(.A1(new_n952), .A2(KEYINPUT50), .ZN(new_n1041));
  NAND2_X1  g616(.A1(new_n1002), .A2(new_n1004), .ZN(new_n1042));
  NOR2_X1   g617(.A1(new_n1041), .A2(new_n1042), .ZN(new_n1043));
  AOI22_X1  g618(.A1(new_n1034), .A2(KEYINPUT111), .B1(new_n1043), .B2(new_n1031), .ZN(new_n1044));
  INV_X1    g619(.A(KEYINPUT111), .ZN(new_n1045));
  NAND2_X1  g620(.A1(new_n1030), .A2(new_n1045), .ZN(new_n1046));
  NAND2_X1  g621(.A1(new_n1044), .A2(new_n1046), .ZN(new_n1047));
  INV_X1    g622(.A(new_n1039), .ZN(new_n1048));
  NAND3_X1  g623(.A1(new_n1047), .A2(G8), .A3(new_n1048), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n553), .A2(G48), .ZN(new_n1050));
  NAND3_X1  g625(.A1(new_n504), .A2(new_n498), .A3(G86), .ZN(new_n1051));
  INV_X1    g626(.A(new_n573), .ZN(new_n1052));
  AOI21_X1  g627(.A(new_n1052), .B1(new_n498), .B2(G61), .ZN(new_n1053));
  OAI211_X1 g628(.A(new_n1050), .B(new_n1051), .C1(new_n1053), .C2(new_n500), .ZN(new_n1054));
  NAND2_X1  g629(.A1(new_n1054), .A2(G1981), .ZN(new_n1055));
  NAND2_X1  g630(.A1(new_n1055), .A2(KEYINPUT113), .ZN(new_n1056));
  INV_X1    g631(.A(G1981), .ZN(new_n1057));
  NAND3_X1  g632(.A1(new_n571), .A2(new_n575), .A3(new_n1057), .ZN(new_n1058));
  INV_X1    g633(.A(KEYINPUT113), .ZN(new_n1059));
  NAND3_X1  g634(.A1(new_n1054), .A2(new_n1059), .A3(G1981), .ZN(new_n1060));
  NAND4_X1  g635(.A1(new_n1056), .A2(KEYINPUT49), .A3(new_n1058), .A4(new_n1060), .ZN(new_n1061));
  NOR2_X1   g636(.A1(new_n952), .A2(new_n959), .ZN(new_n1062));
  NOR2_X1   g637(.A1(new_n1062), .A2(new_n997), .ZN(new_n1063));
  NAND2_X1  g638(.A1(new_n1061), .A2(new_n1063), .ZN(new_n1064));
  XOR2_X1   g639(.A(KEYINPUT114), .B(KEYINPUT49), .Z(new_n1065));
  NAND2_X1  g640(.A1(new_n1060), .A2(new_n1058), .ZN(new_n1066));
  AOI21_X1  g641(.A(new_n1059), .B1(new_n1054), .B2(G1981), .ZN(new_n1067));
  OAI21_X1  g642(.A(new_n1065), .B1(new_n1066), .B2(new_n1067), .ZN(new_n1068));
  INV_X1    g643(.A(KEYINPUT115), .ZN(new_n1069));
  NAND2_X1  g644(.A1(new_n1068), .A2(new_n1069), .ZN(new_n1070));
  OAI211_X1 g645(.A(KEYINPUT115), .B(new_n1065), .C1(new_n1066), .C2(new_n1067), .ZN(new_n1071));
  AOI21_X1  g646(.A(new_n1064), .B1(new_n1070), .B2(new_n1071), .ZN(new_n1072));
  INV_X1    g647(.A(KEYINPUT112), .ZN(new_n1073));
  NAND3_X1  g648(.A1(new_n566), .A2(G1976), .A3(new_n569), .ZN(new_n1074));
  OAI211_X1 g649(.A(new_n1074), .B(G8), .C1(new_n952), .C2(new_n959), .ZN(new_n1075));
  NAND2_X1  g650(.A1(new_n1075), .A2(KEYINPUT52), .ZN(new_n1076));
  INV_X1    g651(.A(new_n1075), .ZN(new_n1077));
  INV_X1    g652(.A(G1976), .ZN(new_n1078));
  AOI21_X1  g653(.A(KEYINPUT52), .B1(G288), .B2(new_n1078), .ZN(new_n1079));
  AND4_X1   g654(.A1(new_n1073), .A2(new_n1076), .A3(new_n1077), .A4(new_n1079), .ZN(new_n1080));
  AOI22_X1  g655(.A1(new_n1073), .A2(new_n1076), .B1(new_n1077), .B2(new_n1079), .ZN(new_n1081));
  NOR3_X1   g656(.A1(new_n1072), .A2(new_n1080), .A3(new_n1081), .ZN(new_n1082));
  INV_X1    g657(.A(G2078), .ZN(new_n1083));
  NAND4_X1  g658(.A1(new_n954), .A2(new_n1083), .A3(new_n1002), .A4(new_n1008), .ZN(new_n1084));
  INV_X1    g659(.A(KEYINPUT53), .ZN(new_n1085));
  NAND2_X1  g660(.A1(new_n1084), .A2(new_n1085), .ZN(new_n1086));
  NAND4_X1  g661(.A1(new_n1029), .A2(KEYINPUT53), .A3(new_n1083), .A4(new_n954), .ZN(new_n1087));
  OAI21_X1  g662(.A(new_n691), .B1(new_n1041), .B2(new_n1042), .ZN(new_n1088));
  NAND3_X1  g663(.A1(new_n1086), .A2(new_n1087), .A3(new_n1088), .ZN(new_n1089));
  AND2_X1   g664(.A1(new_n1089), .A2(G171), .ZN(new_n1090));
  NAND4_X1  g665(.A1(new_n1040), .A2(new_n1049), .A3(new_n1082), .A4(new_n1090), .ZN(new_n1091));
  AOI21_X1  g666(.A(new_n1091), .B1(new_n1025), .B2(new_n1026), .ZN(new_n1092));
  INV_X1    g667(.A(KEYINPUT124), .ZN(new_n1093));
  AOI22_X1  g668(.A1(new_n1019), .A2(new_n1020), .B1(new_n1022), .B2(new_n1023), .ZN(new_n1094));
  OAI211_X1 g669(.A(new_n1093), .B(KEYINPUT62), .C1(new_n1094), .C2(new_n1018), .ZN(new_n1095));
  AND3_X1   g670(.A1(new_n1027), .A2(new_n1092), .A3(new_n1095), .ZN(new_n1096));
  NOR2_X1   g671(.A1(new_n1022), .A2(G286), .ZN(new_n1097));
  NAND4_X1  g672(.A1(new_n1040), .A2(new_n1049), .A3(new_n1082), .A4(new_n1097), .ZN(new_n1098));
  INV_X1    g673(.A(KEYINPUT63), .ZN(new_n1099));
  NAND2_X1  g674(.A1(new_n1098), .A2(new_n1099), .ZN(new_n1100));
  NAND2_X1  g675(.A1(new_n1047), .A2(G8), .ZN(new_n1101));
  NAND2_X1  g676(.A1(new_n1101), .A2(new_n1039), .ZN(new_n1102));
  NOR3_X1   g677(.A1(new_n1022), .A2(new_n1099), .A3(G286), .ZN(new_n1103));
  NAND4_X1  g678(.A1(new_n1102), .A2(new_n1049), .A3(new_n1082), .A4(new_n1103), .ZN(new_n1104));
  NAND2_X1  g679(.A1(new_n1100), .A2(new_n1104), .ZN(new_n1105));
  NOR2_X1   g680(.A1(G288), .A2(G1976), .ZN(new_n1106));
  INV_X1    g681(.A(new_n1106), .ZN(new_n1107));
  OAI21_X1  g682(.A(new_n1058), .B1(new_n1072), .B2(new_n1107), .ZN(new_n1108));
  AOI211_X1 g683(.A(new_n997), .B(new_n1062), .C1(new_n1108), .C2(KEYINPUT116), .ZN(new_n1109));
  INV_X1    g684(.A(KEYINPUT116), .ZN(new_n1110));
  OAI211_X1 g685(.A(new_n1110), .B(new_n1058), .C1(new_n1072), .C2(new_n1107), .ZN(new_n1111));
  INV_X1    g686(.A(new_n1049), .ZN(new_n1112));
  AOI22_X1  g687(.A1(new_n1109), .A2(new_n1111), .B1(new_n1112), .B2(new_n1082), .ZN(new_n1113));
  OAI21_X1  g688(.A(new_n774), .B1(new_n1041), .B2(new_n1042), .ZN(new_n1114));
  INV_X1    g689(.A(KEYINPUT57), .ZN(new_n1115));
  XNOR2_X1  g690(.A(G299), .B(new_n1115), .ZN(new_n1116));
  XNOR2_X1  g691(.A(KEYINPUT56), .B(G2072), .ZN(new_n1117));
  NAND4_X1  g692(.A1(new_n954), .A2(new_n1002), .A3(new_n1008), .A4(new_n1117), .ZN(new_n1118));
  AND3_X1   g693(.A1(new_n1114), .A2(new_n1116), .A3(new_n1118), .ZN(new_n1119));
  INV_X1    g694(.A(G1348), .ZN(new_n1120));
  OAI21_X1  g695(.A(new_n1120), .B1(new_n1041), .B2(new_n1042), .ZN(new_n1121));
  NOR3_X1   g696(.A1(new_n952), .A2(new_n959), .A3(G2067), .ZN(new_n1122));
  INV_X1    g697(.A(new_n1122), .ZN(new_n1123));
  AOI21_X1  g698(.A(new_n608), .B1(new_n1121), .B2(new_n1123), .ZN(new_n1124));
  INV_X1    g699(.A(new_n1124), .ZN(new_n1125));
  OR2_X1    g700(.A1(new_n1125), .A2(KEYINPUT119), .ZN(new_n1126));
  AOI21_X1  g701(.A(new_n1116), .B1(new_n1114), .B2(new_n1118), .ZN(new_n1127));
  AOI21_X1  g702(.A(new_n1127), .B1(new_n1125), .B2(KEYINPUT119), .ZN(new_n1128));
  AOI21_X1  g703(.A(new_n1119), .B1(new_n1126), .B2(new_n1128), .ZN(new_n1129));
  AND3_X1   g704(.A1(new_n1121), .A2(new_n608), .A3(new_n1123), .ZN(new_n1130));
  OAI21_X1  g705(.A(KEYINPUT60), .B1(new_n1130), .B2(new_n1124), .ZN(new_n1131));
  INV_X1    g706(.A(new_n1116), .ZN(new_n1132));
  INV_X1    g707(.A(new_n1118), .ZN(new_n1133));
  AOI21_X1  g708(.A(G1956), .B1(new_n1011), .B2(new_n1000), .ZN(new_n1134));
  OAI21_X1  g709(.A(new_n1132), .B1(new_n1133), .B2(new_n1134), .ZN(new_n1135));
  NAND3_X1  g710(.A1(new_n1114), .A2(new_n1116), .A3(new_n1118), .ZN(new_n1136));
  NAND3_X1  g711(.A1(new_n1135), .A2(KEYINPUT61), .A3(new_n1136), .ZN(new_n1137));
  INV_X1    g712(.A(KEYINPUT60), .ZN(new_n1138));
  NAND4_X1  g713(.A1(new_n1121), .A2(new_n1138), .A3(new_n598), .A4(new_n1123), .ZN(new_n1139));
  NAND3_X1  g714(.A1(new_n1131), .A2(new_n1137), .A3(new_n1139), .ZN(new_n1140));
  INV_X1    g715(.A(KEYINPUT61), .ZN(new_n1141));
  OAI21_X1  g716(.A(new_n1141), .B1(new_n1119), .B2(new_n1127), .ZN(new_n1142));
  INV_X1    g717(.A(KEYINPUT121), .ZN(new_n1143));
  NAND2_X1  g718(.A1(new_n1142), .A2(new_n1143), .ZN(new_n1144));
  OAI211_X1 g719(.A(KEYINPUT121), .B(new_n1141), .C1(new_n1119), .C2(new_n1127), .ZN(new_n1145));
  AOI21_X1  g720(.A(new_n1140), .B1(new_n1144), .B2(new_n1145), .ZN(new_n1146));
  NAND4_X1  g721(.A1(new_n954), .A2(new_n961), .A3(new_n1002), .A4(new_n1008), .ZN(new_n1147));
  INV_X1    g722(.A(KEYINPUT120), .ZN(new_n1148));
  XOR2_X1   g723(.A(KEYINPUT58), .B(G1341), .Z(new_n1149));
  OAI21_X1  g724(.A(new_n1149), .B1(new_n952), .B2(new_n959), .ZN(new_n1150));
  AND3_X1   g725(.A1(new_n1147), .A2(new_n1148), .A3(new_n1150), .ZN(new_n1151));
  AOI21_X1  g726(.A(new_n1148), .B1(new_n1147), .B2(new_n1150), .ZN(new_n1152));
  OAI21_X1  g727(.A(new_n541), .B1(new_n1151), .B2(new_n1152), .ZN(new_n1153));
  NAND2_X1  g728(.A1(new_n1153), .A2(KEYINPUT59), .ZN(new_n1154));
  INV_X1    g729(.A(KEYINPUT59), .ZN(new_n1155));
  OAI211_X1 g730(.A(new_n1155), .B(new_n541), .C1(new_n1151), .C2(new_n1152), .ZN(new_n1156));
  NAND2_X1  g731(.A1(new_n1154), .A2(new_n1156), .ZN(new_n1157));
  AOI21_X1  g732(.A(new_n1129), .B1(new_n1146), .B2(new_n1157), .ZN(new_n1158));
  AND3_X1   g733(.A1(new_n1040), .A2(new_n1049), .A3(new_n1082), .ZN(new_n1159));
  AND2_X1   g734(.A1(new_n1086), .A2(new_n1087), .ZN(new_n1160));
  INV_X1    g735(.A(KEYINPUT123), .ZN(new_n1161));
  XOR2_X1   g736(.A(G171), .B(KEYINPUT54), .Z(new_n1162));
  OAI211_X1 g737(.A(new_n1160), .B(new_n1088), .C1(new_n1161), .C2(new_n1162), .ZN(new_n1163));
  NAND3_X1  g738(.A1(new_n1086), .A2(new_n1087), .A3(new_n1161), .ZN(new_n1164));
  INV_X1    g739(.A(new_n1162), .ZN(new_n1165));
  NAND3_X1  g740(.A1(new_n1089), .A2(new_n1164), .A3(new_n1165), .ZN(new_n1166));
  NAND2_X1  g741(.A1(new_n1163), .A2(new_n1166), .ZN(new_n1167));
  OAI211_X1 g742(.A(new_n1159), .B(new_n1167), .C1(new_n1018), .C2(new_n1094), .ZN(new_n1168));
  OAI211_X1 g743(.A(new_n1105), .B(new_n1113), .C1(new_n1158), .C2(new_n1168), .ZN(new_n1169));
  OAI211_X1 g744(.A(KEYINPUT125), .B(new_n996), .C1(new_n1096), .C2(new_n1169), .ZN(new_n1170));
  INV_X1    g745(.A(new_n1170), .ZN(new_n1171));
  NAND3_X1  g746(.A1(new_n1027), .A2(new_n1092), .A3(new_n1095), .ZN(new_n1172));
  NAND2_X1  g747(.A1(new_n1112), .A2(new_n1082), .ZN(new_n1173));
  NAND2_X1  g748(.A1(new_n1108), .A2(KEYINPUT116), .ZN(new_n1174));
  NAND2_X1  g749(.A1(new_n1174), .A2(new_n1063), .ZN(new_n1175));
  INV_X1    g750(.A(new_n1111), .ZN(new_n1176));
  OAI21_X1  g751(.A(new_n1173), .B1(new_n1175), .B2(new_n1176), .ZN(new_n1177));
  NAND4_X1  g752(.A1(new_n1167), .A2(new_n1049), .A3(new_n1082), .A4(new_n1040), .ZN(new_n1178));
  NOR2_X1   g753(.A1(new_n1025), .A2(new_n1178), .ZN(new_n1179));
  NAND2_X1  g754(.A1(new_n1144), .A2(new_n1145), .ZN(new_n1180));
  AND3_X1   g755(.A1(new_n1131), .A2(new_n1137), .A3(new_n1139), .ZN(new_n1181));
  NAND3_X1  g756(.A1(new_n1180), .A2(new_n1181), .A3(new_n1157), .ZN(new_n1182));
  INV_X1    g757(.A(new_n1129), .ZN(new_n1183));
  NAND2_X1  g758(.A1(new_n1182), .A2(new_n1183), .ZN(new_n1184));
  AOI21_X1  g759(.A(new_n1177), .B1(new_n1179), .B2(new_n1184), .ZN(new_n1185));
  NAND3_X1  g760(.A1(new_n1172), .A2(new_n1185), .A3(new_n1105), .ZN(new_n1186));
  AOI21_X1  g761(.A(KEYINPUT125), .B1(new_n1186), .B2(new_n996), .ZN(new_n1187));
  OAI21_X1  g762(.A(new_n993), .B1(new_n1171), .B2(new_n1187), .ZN(G329));
  assign    G231 = 1'b0;
  NOR2_X1   g763(.A1(G227), .A2(new_n459), .ZN(new_n1190));
  NAND3_X1  g764(.A1(new_n685), .A2(new_n686), .A3(new_n1190), .ZN(new_n1191));
  NOR2_X1   g765(.A1(new_n1191), .A2(G401), .ZN(new_n1192));
  OAI211_X1 g766(.A(new_n1192), .B(new_n890), .C1(new_n936), .C2(new_n944), .ZN(G225));
  INV_X1    g767(.A(G225), .ZN(G308));
endmodule


