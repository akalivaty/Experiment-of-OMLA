//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 0 0 1 0 0 0 1 0 1 1 1 1 0 0 1 1 1 0 1 0 1 1 0 0 0 0 1 0 0 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 0 0 1 1 0 1 0 0 1 0 1 1 1 1 0 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:21:17 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n663, new_n664, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n695, new_n696,
    new_n697, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n726, new_n727, new_n728,
    new_n729, new_n731, new_n732, new_n733, new_n734, new_n736, new_n738,
    new_n739, new_n740, new_n741, new_n742, new_n743, new_n744, new_n745,
    new_n746, new_n747, new_n748, new_n749, new_n750, new_n751, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n761,
    new_n762, new_n763, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n819, new_n820,
    new_n822, new_n823, new_n825, new_n826, new_n827, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n913, new_n914, new_n915, new_n916,
    new_n918, new_n919, new_n920, new_n921, new_n922, new_n923, new_n924,
    new_n925, new_n926, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n939, new_n940,
    new_n942, new_n943, new_n944, new_n945, new_n946, new_n948, new_n949,
    new_n950, new_n951, new_n953, new_n954, new_n955, new_n956, new_n957,
    new_n958, new_n959, new_n960, new_n961, new_n962, new_n963, new_n964,
    new_n965, new_n967, new_n968, new_n969, new_n970, new_n971, new_n973,
    new_n974, new_n975, new_n976, new_n977, new_n978, new_n980, new_n981,
    new_n982, new_n983, new_n984;
  XNOR2_X1  g000(.A(G15gat), .B(G22gat), .ZN(new_n202));
  INV_X1    g001(.A(KEYINPUT16), .ZN(new_n203));
  AOI21_X1  g002(.A(G1gat), .B1(new_n202), .B2(new_n203), .ZN(new_n204));
  INV_X1    g003(.A(G8gat), .ZN(new_n205));
  NAND2_X1  g004(.A1(new_n204), .A2(new_n205), .ZN(new_n206));
  INV_X1    g005(.A(new_n206), .ZN(new_n207));
  NOR2_X1   g006(.A1(new_n204), .A2(new_n205), .ZN(new_n208));
  XOR2_X1   g007(.A(G15gat), .B(G22gat), .Z(new_n209));
  OAI22_X1  g008(.A1(new_n207), .A2(new_n208), .B1(KEYINPUT89), .B2(new_n209), .ZN(new_n210));
  INV_X1    g009(.A(KEYINPUT14), .ZN(new_n211));
  INV_X1    g010(.A(G29gat), .ZN(new_n212));
  INV_X1    g011(.A(G36gat), .ZN(new_n213));
  NAND3_X1  g012(.A1(new_n211), .A2(new_n212), .A3(new_n213), .ZN(new_n214));
  OAI21_X1  g013(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n215));
  AOI22_X1  g014(.A1(new_n214), .A2(new_n215), .B1(G29gat), .B2(G36gat), .ZN(new_n216));
  INV_X1    g015(.A(KEYINPUT15), .ZN(new_n217));
  XOR2_X1   g016(.A(G43gat), .B(G50gat), .Z(new_n218));
  OR3_X1    g017(.A1(new_n216), .A2(new_n217), .A3(new_n218), .ZN(new_n219));
  NAND2_X1  g018(.A1(new_n218), .A2(new_n217), .ZN(new_n220));
  XNOR2_X1  g019(.A(G43gat), .B(G50gat), .ZN(new_n221));
  NAND2_X1  g020(.A1(new_n221), .A2(KEYINPUT15), .ZN(new_n222));
  NAND3_X1  g021(.A1(new_n220), .A2(new_n222), .A3(new_n216), .ZN(new_n223));
  NAND2_X1  g022(.A1(new_n219), .A2(new_n223), .ZN(new_n224));
  INV_X1    g023(.A(G1gat), .ZN(new_n225));
  OAI21_X1  g024(.A(new_n225), .B1(new_n209), .B2(KEYINPUT16), .ZN(new_n226));
  NAND2_X1  g025(.A1(new_n226), .A2(G8gat), .ZN(new_n227));
  NOR2_X1   g026(.A1(new_n209), .A2(KEYINPUT89), .ZN(new_n228));
  NAND3_X1  g027(.A1(new_n227), .A2(new_n228), .A3(new_n206), .ZN(new_n229));
  NAND3_X1  g028(.A1(new_n210), .A2(new_n224), .A3(new_n229), .ZN(new_n230));
  INV_X1    g029(.A(KEYINPUT90), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n230), .A2(new_n231), .ZN(new_n232));
  NAND4_X1  g031(.A1(new_n210), .A2(KEYINPUT90), .A3(new_n224), .A4(new_n229), .ZN(new_n233));
  NAND2_X1  g032(.A1(new_n232), .A2(new_n233), .ZN(new_n234));
  NAND2_X1  g033(.A1(new_n210), .A2(new_n229), .ZN(new_n235));
  INV_X1    g034(.A(new_n235), .ZN(new_n236));
  OAI21_X1  g035(.A(new_n234), .B1(new_n224), .B2(new_n236), .ZN(new_n237));
  NAND2_X1  g036(.A1(G229gat), .A2(G233gat), .ZN(new_n238));
  XOR2_X1   g037(.A(new_n238), .B(KEYINPUT13), .Z(new_n239));
  NAND2_X1  g038(.A1(new_n237), .A2(new_n239), .ZN(new_n240));
  INV_X1    g039(.A(KEYINPUT91), .ZN(new_n241));
  NAND3_X1  g040(.A1(new_n219), .A2(KEYINPUT17), .A3(new_n223), .ZN(new_n242));
  INV_X1    g041(.A(KEYINPUT17), .ZN(new_n243));
  NAND2_X1  g042(.A1(new_n224), .A2(new_n243), .ZN(new_n244));
  NAND3_X1  g043(.A1(new_n235), .A2(new_n242), .A3(new_n244), .ZN(new_n245));
  NAND4_X1  g044(.A1(new_n234), .A2(new_n241), .A3(new_n238), .A4(new_n245), .ZN(new_n246));
  AOI21_X1  g045(.A(KEYINPUT18), .B1(new_n246), .B2(KEYINPUT92), .ZN(new_n247));
  AOI21_X1  g046(.A(KEYINPUT91), .B1(KEYINPUT92), .B2(KEYINPUT18), .ZN(new_n248));
  AND2_X1   g047(.A1(new_n244), .A2(new_n242), .ZN(new_n249));
  AOI22_X1  g048(.A1(new_n232), .A2(new_n233), .B1(new_n249), .B2(new_n235), .ZN(new_n250));
  AOI21_X1  g049(.A(new_n248), .B1(new_n250), .B2(new_n238), .ZN(new_n251));
  OAI21_X1  g050(.A(new_n240), .B1(new_n247), .B2(new_n251), .ZN(new_n252));
  XNOR2_X1  g051(.A(G113gat), .B(G141gat), .ZN(new_n253));
  INV_X1    g052(.A(G197gat), .ZN(new_n254));
  XNOR2_X1  g053(.A(new_n253), .B(new_n254), .ZN(new_n255));
  XNOR2_X1  g054(.A(KEYINPUT11), .B(G169gat), .ZN(new_n256));
  XNOR2_X1  g055(.A(new_n255), .B(new_n256), .ZN(new_n257));
  XOR2_X1   g056(.A(new_n257), .B(KEYINPUT12), .Z(new_n258));
  NAND2_X1  g057(.A1(new_n252), .A2(new_n258), .ZN(new_n259));
  INV_X1    g058(.A(new_n258), .ZN(new_n260));
  OAI211_X1 g059(.A(new_n240), .B(new_n260), .C1(new_n247), .C2(new_n251), .ZN(new_n261));
  NAND2_X1  g060(.A1(new_n259), .A2(new_n261), .ZN(new_n262));
  INV_X1    g061(.A(new_n262), .ZN(new_n263));
  INV_X1    g062(.A(KEYINPUT7), .ZN(new_n264));
  NOR2_X1   g063(.A1(new_n264), .A2(KEYINPUT96), .ZN(new_n265));
  INV_X1    g064(.A(new_n265), .ZN(new_n266));
  NAND2_X1  g065(.A1(G85gat), .A2(G92gat), .ZN(new_n267));
  INV_X1    g066(.A(KEYINPUT97), .ZN(new_n268));
  INV_X1    g067(.A(KEYINPUT96), .ZN(new_n269));
  OAI211_X1 g068(.A(new_n267), .B(new_n268), .C1(new_n269), .C2(KEYINPUT7), .ZN(new_n270));
  INV_X1    g069(.A(new_n270), .ZN(new_n271));
  NAND2_X1  g070(.A1(new_n264), .A2(KEYINPUT96), .ZN(new_n272));
  AOI21_X1  g071(.A(new_n268), .B1(new_n272), .B2(new_n267), .ZN(new_n273));
  OAI21_X1  g072(.A(new_n266), .B1(new_n271), .B2(new_n273), .ZN(new_n274));
  NAND2_X1  g073(.A1(G99gat), .A2(G106gat), .ZN(new_n275));
  INV_X1    g074(.A(G85gat), .ZN(new_n276));
  INV_X1    g075(.A(G92gat), .ZN(new_n277));
  AOI22_X1  g076(.A1(KEYINPUT8), .A2(new_n275), .B1(new_n276), .B2(new_n277), .ZN(new_n278));
  OAI21_X1  g077(.A(new_n267), .B1(new_n269), .B2(KEYINPUT7), .ZN(new_n279));
  NAND2_X1  g078(.A1(new_n279), .A2(KEYINPUT97), .ZN(new_n280));
  NAND3_X1  g079(.A1(new_n280), .A2(new_n265), .A3(new_n270), .ZN(new_n281));
  NAND3_X1  g080(.A1(new_n274), .A2(new_n278), .A3(new_n281), .ZN(new_n282));
  XNOR2_X1  g081(.A(G99gat), .B(G106gat), .ZN(new_n283));
  INV_X1    g082(.A(new_n283), .ZN(new_n284));
  NAND2_X1  g083(.A1(new_n282), .A2(new_n284), .ZN(new_n285));
  NAND4_X1  g084(.A1(new_n274), .A2(new_n283), .A3(new_n281), .A4(new_n278), .ZN(new_n286));
  NAND2_X1  g085(.A1(G71gat), .A2(G78gat), .ZN(new_n287));
  INV_X1    g086(.A(G71gat), .ZN(new_n288));
  INV_X1    g087(.A(G78gat), .ZN(new_n289));
  NAND2_X1  g088(.A1(new_n288), .A2(new_n289), .ZN(new_n290));
  XNOR2_X1  g089(.A(G57gat), .B(G64gat), .ZN(new_n291));
  INV_X1    g090(.A(KEYINPUT9), .ZN(new_n292));
  OAI211_X1 g091(.A(new_n287), .B(new_n290), .C1(new_n291), .C2(new_n292), .ZN(new_n293));
  AND2_X1   g092(.A1(G71gat), .A2(G78gat), .ZN(new_n294));
  NOR2_X1   g093(.A1(G71gat), .A2(G78gat), .ZN(new_n295));
  OAI21_X1  g094(.A(KEYINPUT93), .B1(new_n294), .B2(new_n295), .ZN(new_n296));
  INV_X1    g095(.A(KEYINPUT93), .ZN(new_n297));
  NAND3_X1  g096(.A1(new_n290), .A2(new_n297), .A3(new_n287), .ZN(new_n298));
  NAND2_X1  g097(.A1(new_n296), .A2(new_n298), .ZN(new_n299));
  NAND2_X1  g098(.A1(new_n287), .A2(new_n292), .ZN(new_n300));
  INV_X1    g099(.A(G64gat), .ZN(new_n301));
  AND2_X1   g100(.A1(new_n301), .A2(G57gat), .ZN(new_n302));
  NOR2_X1   g101(.A1(new_n301), .A2(G57gat), .ZN(new_n303));
  OAI21_X1  g102(.A(new_n300), .B1(new_n302), .B2(new_n303), .ZN(new_n304));
  OAI21_X1  g103(.A(new_n293), .B1(new_n299), .B2(new_n304), .ZN(new_n305));
  AND3_X1   g104(.A1(new_n285), .A2(new_n286), .A3(new_n305), .ZN(new_n306));
  NAND2_X1  g105(.A1(new_n305), .A2(KEYINPUT94), .ZN(new_n307));
  XOR2_X1   g106(.A(G57gat), .B(G64gat), .Z(new_n308));
  NAND4_X1  g107(.A1(new_n308), .A2(new_n296), .A3(new_n298), .A4(new_n300), .ZN(new_n309));
  INV_X1    g108(.A(KEYINPUT94), .ZN(new_n310));
  NAND3_X1  g109(.A1(new_n309), .A2(new_n310), .A3(new_n293), .ZN(new_n311));
  AOI22_X1  g110(.A1(new_n285), .A2(new_n286), .B1(new_n307), .B2(new_n311), .ZN(new_n312));
  NAND2_X1  g111(.A1(G230gat), .A2(G233gat), .ZN(new_n313));
  NOR3_X1   g112(.A1(new_n306), .A2(new_n312), .A3(new_n313), .ZN(new_n314));
  AND2_X1   g113(.A1(new_n314), .A2(KEYINPUT99), .ZN(new_n315));
  XNOR2_X1  g114(.A(G120gat), .B(G148gat), .ZN(new_n316));
  XNOR2_X1  g115(.A(G176gat), .B(G204gat), .ZN(new_n317));
  XNOR2_X1  g116(.A(new_n316), .B(new_n317), .ZN(new_n318));
  INV_X1    g117(.A(new_n318), .ZN(new_n319));
  OAI21_X1  g118(.A(new_n319), .B1(new_n314), .B2(KEYINPUT99), .ZN(new_n320));
  INV_X1    g119(.A(new_n313), .ZN(new_n321));
  INV_X1    g120(.A(KEYINPUT10), .ZN(new_n322));
  OAI21_X1  g121(.A(new_n322), .B1(new_n306), .B2(new_n312), .ZN(new_n323));
  AND2_X1   g122(.A1(new_n285), .A2(new_n286), .ZN(new_n324));
  NAND3_X1  g123(.A1(new_n307), .A2(KEYINPUT95), .A3(new_n311), .ZN(new_n325));
  INV_X1    g124(.A(KEYINPUT95), .ZN(new_n326));
  AND3_X1   g125(.A1(new_n309), .A2(new_n310), .A3(new_n293), .ZN(new_n327));
  AOI21_X1  g126(.A(new_n310), .B1(new_n309), .B2(new_n293), .ZN(new_n328));
  OAI21_X1  g127(.A(new_n326), .B1(new_n327), .B2(new_n328), .ZN(new_n329));
  NAND4_X1  g128(.A1(new_n324), .A2(KEYINPUT10), .A3(new_n325), .A4(new_n329), .ZN(new_n330));
  AOI21_X1  g129(.A(new_n321), .B1(new_n323), .B2(new_n330), .ZN(new_n331));
  NOR3_X1   g130(.A1(new_n315), .A2(new_n320), .A3(new_n331), .ZN(new_n332));
  INV_X1    g131(.A(new_n332), .ZN(new_n333));
  OAI21_X1  g132(.A(new_n318), .B1(new_n331), .B2(new_n314), .ZN(new_n334));
  NAND2_X1  g133(.A1(new_n333), .A2(new_n334), .ZN(new_n335));
  NOR2_X1   g134(.A1(new_n263), .A2(new_n335), .ZN(new_n336));
  INV_X1    g135(.A(new_n336), .ZN(new_n337));
  NAND2_X1  g136(.A1(new_n307), .A2(new_n311), .ZN(new_n338));
  OR2_X1    g137(.A1(new_n338), .A2(KEYINPUT21), .ZN(new_n339));
  XNOR2_X1  g138(.A(new_n339), .B(G211gat), .ZN(new_n340));
  INV_X1    g139(.A(new_n340), .ZN(new_n341));
  AND2_X1   g140(.A1(new_n329), .A2(new_n325), .ZN(new_n342));
  AOI21_X1  g141(.A(new_n236), .B1(new_n342), .B2(KEYINPUT21), .ZN(new_n343));
  INV_X1    g142(.A(G183gat), .ZN(new_n344));
  NAND2_X1  g143(.A1(new_n343), .A2(new_n344), .ZN(new_n345));
  INV_X1    g144(.A(new_n345), .ZN(new_n346));
  NOR2_X1   g145(.A1(new_n343), .A2(new_n344), .ZN(new_n347));
  XNOR2_X1  g146(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n348));
  INV_X1    g147(.A(new_n348), .ZN(new_n349));
  NOR3_X1   g148(.A1(new_n346), .A2(new_n347), .A3(new_n349), .ZN(new_n350));
  NAND2_X1  g149(.A1(new_n342), .A2(KEYINPUT21), .ZN(new_n351));
  NAND2_X1  g150(.A1(new_n351), .A2(new_n235), .ZN(new_n352));
  NAND2_X1  g151(.A1(new_n352), .A2(G183gat), .ZN(new_n353));
  AOI21_X1  g152(.A(new_n348), .B1(new_n353), .B2(new_n345), .ZN(new_n354));
  OAI21_X1  g153(.A(new_n341), .B1(new_n350), .B2(new_n354), .ZN(new_n355));
  OAI21_X1  g154(.A(new_n349), .B1(new_n346), .B2(new_n347), .ZN(new_n356));
  NAND3_X1  g155(.A1(new_n353), .A2(new_n345), .A3(new_n348), .ZN(new_n357));
  NAND3_X1  g156(.A1(new_n356), .A2(new_n357), .A3(new_n340), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n355), .A2(new_n358), .ZN(new_n359));
  XNOR2_X1  g158(.A(G127gat), .B(G155gat), .ZN(new_n360));
  NAND2_X1  g159(.A1(G231gat), .A2(G233gat), .ZN(new_n361));
  XNOR2_X1  g160(.A(new_n360), .B(new_n361), .ZN(new_n362));
  INV_X1    g161(.A(new_n362), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n359), .A2(new_n363), .ZN(new_n364));
  NAND3_X1  g163(.A1(new_n355), .A2(new_n362), .A3(new_n358), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n364), .A2(new_n365), .ZN(new_n366));
  NAND2_X1  g165(.A1(new_n285), .A2(new_n286), .ZN(new_n367));
  NAND2_X1  g166(.A1(new_n249), .A2(new_n367), .ZN(new_n368));
  NAND3_X1  g167(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n369));
  NAND2_X1  g168(.A1(new_n324), .A2(new_n224), .ZN(new_n370));
  NAND3_X1  g169(.A1(new_n368), .A2(new_n369), .A3(new_n370), .ZN(new_n371));
  XNOR2_X1  g170(.A(G190gat), .B(G218gat), .ZN(new_n372));
  INV_X1    g171(.A(new_n372), .ZN(new_n373));
  NAND2_X1  g172(.A1(new_n371), .A2(new_n373), .ZN(new_n374));
  INV_X1    g173(.A(KEYINPUT98), .ZN(new_n375));
  NAND4_X1  g174(.A1(new_n368), .A2(new_n369), .A3(new_n370), .A4(new_n372), .ZN(new_n376));
  NAND3_X1  g175(.A1(new_n374), .A2(new_n375), .A3(new_n376), .ZN(new_n377));
  INV_X1    g176(.A(new_n377), .ZN(new_n378));
  AOI21_X1  g177(.A(new_n375), .B1(new_n374), .B2(new_n376), .ZN(new_n379));
  XNOR2_X1  g178(.A(G134gat), .B(G162gat), .ZN(new_n380));
  AOI21_X1  g179(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n381));
  XOR2_X1   g180(.A(new_n380), .B(new_n381), .Z(new_n382));
  NOR3_X1   g181(.A1(new_n378), .A2(new_n379), .A3(new_n382), .ZN(new_n383));
  NAND2_X1  g182(.A1(new_n379), .A2(new_n382), .ZN(new_n384));
  INV_X1    g183(.A(new_n384), .ZN(new_n385));
  NOR2_X1   g184(.A1(new_n383), .A2(new_n385), .ZN(new_n386));
  INV_X1    g185(.A(new_n386), .ZN(new_n387));
  NAND2_X1  g186(.A1(new_n366), .A2(new_n387), .ZN(new_n388));
  INV_X1    g187(.A(KEYINPUT82), .ZN(new_n389));
  INV_X1    g188(.A(G148gat), .ZN(new_n390));
  NOR2_X1   g189(.A1(KEYINPUT79), .A2(G141gat), .ZN(new_n391));
  INV_X1    g190(.A(new_n391), .ZN(new_n392));
  NAND2_X1  g191(.A1(KEYINPUT79), .A2(G141gat), .ZN(new_n393));
  AOI21_X1  g192(.A(new_n390), .B1(new_n392), .B2(new_n393), .ZN(new_n394));
  INV_X1    g193(.A(G141gat), .ZN(new_n395));
  NAND2_X1  g194(.A1(new_n390), .A2(KEYINPUT80), .ZN(new_n396));
  INV_X1    g195(.A(KEYINPUT80), .ZN(new_n397));
  NAND2_X1  g196(.A1(new_n397), .A2(G148gat), .ZN(new_n398));
  AOI21_X1  g197(.A(new_n395), .B1(new_n396), .B2(new_n398), .ZN(new_n399));
  OAI21_X1  g198(.A(KEYINPUT81), .B1(new_n394), .B2(new_n399), .ZN(new_n400));
  AND2_X1   g199(.A1(KEYINPUT79), .A2(G141gat), .ZN(new_n401));
  OAI21_X1  g200(.A(G148gat), .B1(new_n401), .B2(new_n391), .ZN(new_n402));
  INV_X1    g201(.A(KEYINPUT81), .ZN(new_n403));
  XNOR2_X1  g202(.A(KEYINPUT80), .B(G148gat), .ZN(new_n404));
  OAI211_X1 g203(.A(new_n402), .B(new_n403), .C1(new_n395), .C2(new_n404), .ZN(new_n405));
  NAND2_X1  g204(.A1(new_n400), .A2(new_n405), .ZN(new_n406));
  NOR2_X1   g205(.A1(G155gat), .A2(G162gat), .ZN(new_n407));
  INV_X1    g206(.A(KEYINPUT2), .ZN(new_n408));
  NAND2_X1  g207(.A1(new_n407), .A2(new_n408), .ZN(new_n409));
  NAND2_X1  g208(.A1(G155gat), .A2(G162gat), .ZN(new_n410));
  NAND2_X1  g209(.A1(new_n409), .A2(new_n410), .ZN(new_n411));
  NAND2_X1  g210(.A1(new_n406), .A2(new_n411), .ZN(new_n412));
  XOR2_X1   g211(.A(new_n407), .B(KEYINPUT78), .Z(new_n413));
  INV_X1    g212(.A(new_n410), .ZN(new_n414));
  NAND2_X1  g213(.A1(new_n390), .A2(G141gat), .ZN(new_n415));
  NAND2_X1  g214(.A1(new_n395), .A2(G148gat), .ZN(new_n416));
  AOI21_X1  g215(.A(KEYINPUT2), .B1(new_n415), .B2(new_n416), .ZN(new_n417));
  NOR3_X1   g216(.A1(new_n413), .A2(new_n414), .A3(new_n417), .ZN(new_n418));
  INV_X1    g217(.A(new_n418), .ZN(new_n419));
  AOI21_X1  g218(.A(new_n389), .B1(new_n412), .B2(new_n419), .ZN(new_n420));
  AOI22_X1  g219(.A1(new_n400), .A2(new_n405), .B1(new_n410), .B2(new_n409), .ZN(new_n421));
  NOR3_X1   g220(.A1(new_n421), .A2(KEYINPUT82), .A3(new_n418), .ZN(new_n422));
  OAI21_X1  g221(.A(KEYINPUT3), .B1(new_n420), .B2(new_n422), .ZN(new_n423));
  INV_X1    g222(.A(KEYINPUT1), .ZN(new_n424));
  XNOR2_X1  g223(.A(G127gat), .B(G134gat), .ZN(new_n425));
  XNOR2_X1  g224(.A(KEYINPUT68), .B(G120gat), .ZN(new_n426));
  INV_X1    g225(.A(G113gat), .ZN(new_n427));
  NOR2_X1   g226(.A1(new_n426), .A2(new_n427), .ZN(new_n428));
  AND2_X1   g227(.A1(new_n427), .A2(G120gat), .ZN(new_n429));
  OAI211_X1 g228(.A(new_n424), .B(new_n425), .C1(new_n428), .C2(new_n429), .ZN(new_n430));
  XNOR2_X1  g229(.A(G113gat), .B(G120gat), .ZN(new_n431));
  NOR2_X1   g230(.A1(new_n431), .A2(KEYINPUT1), .ZN(new_n432));
  OR2_X1    g231(.A1(new_n432), .A2(new_n425), .ZN(new_n433));
  NAND2_X1  g232(.A1(new_n430), .A2(new_n433), .ZN(new_n434));
  NOR3_X1   g233(.A1(new_n421), .A2(KEYINPUT3), .A3(new_n418), .ZN(new_n435));
  INV_X1    g234(.A(new_n435), .ZN(new_n436));
  NAND3_X1  g235(.A1(new_n423), .A2(new_n434), .A3(new_n436), .ZN(new_n437));
  AND2_X1   g236(.A1(new_n430), .A2(new_n433), .ZN(new_n438));
  NAND3_X1  g237(.A1(new_n438), .A2(new_n412), .A3(new_n419), .ZN(new_n439));
  XNOR2_X1  g238(.A(new_n439), .B(KEYINPUT4), .ZN(new_n440));
  INV_X1    g239(.A(KEYINPUT5), .ZN(new_n441));
  NAND2_X1  g240(.A1(G225gat), .A2(G233gat), .ZN(new_n442));
  NAND4_X1  g241(.A1(new_n437), .A2(new_n440), .A3(new_n441), .A4(new_n442), .ZN(new_n443));
  INV_X1    g242(.A(KEYINPUT3), .ZN(new_n444));
  NAND3_X1  g243(.A1(new_n412), .A2(new_n419), .A3(new_n389), .ZN(new_n445));
  OAI21_X1  g244(.A(KEYINPUT82), .B1(new_n421), .B2(new_n418), .ZN(new_n446));
  AOI21_X1  g245(.A(new_n444), .B1(new_n445), .B2(new_n446), .ZN(new_n447));
  NOR3_X1   g246(.A1(new_n447), .A2(new_n438), .A3(new_n435), .ZN(new_n448));
  INV_X1    g247(.A(KEYINPUT4), .ZN(new_n449));
  XNOR2_X1  g248(.A(new_n439), .B(new_n449), .ZN(new_n450));
  INV_X1    g249(.A(new_n442), .ZN(new_n451));
  NOR3_X1   g250(.A1(new_n448), .A2(new_n450), .A3(new_n451), .ZN(new_n452));
  OAI211_X1 g251(.A(KEYINPUT83), .B(new_n434), .C1(new_n420), .C2(new_n422), .ZN(new_n453));
  AOI21_X1  g252(.A(new_n438), .B1(new_n445), .B2(new_n446), .ZN(new_n454));
  INV_X1    g253(.A(KEYINPUT83), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n439), .A2(new_n455), .ZN(new_n456));
  OAI211_X1 g255(.A(new_n453), .B(new_n451), .C1(new_n454), .C2(new_n456), .ZN(new_n457));
  NAND2_X1  g256(.A1(new_n457), .A2(KEYINPUT5), .ZN(new_n458));
  OAI21_X1  g257(.A(new_n443), .B1(new_n452), .B2(new_n458), .ZN(new_n459));
  XNOR2_X1  g258(.A(G1gat), .B(G29gat), .ZN(new_n460));
  XNOR2_X1  g259(.A(new_n460), .B(new_n276), .ZN(new_n461));
  XNOR2_X1  g260(.A(KEYINPUT0), .B(G57gat), .ZN(new_n462));
  XOR2_X1   g261(.A(new_n461), .B(new_n462), .Z(new_n463));
  NAND2_X1  g262(.A1(new_n459), .A2(new_n463), .ZN(new_n464));
  INV_X1    g263(.A(KEYINPUT6), .ZN(new_n465));
  INV_X1    g264(.A(new_n463), .ZN(new_n466));
  OAI211_X1 g265(.A(new_n443), .B(new_n466), .C1(new_n452), .C2(new_n458), .ZN(new_n467));
  NAND3_X1  g266(.A1(new_n464), .A2(new_n465), .A3(new_n467), .ZN(new_n468));
  NAND3_X1  g267(.A1(new_n459), .A2(KEYINPUT6), .A3(new_n463), .ZN(new_n469));
  NAND2_X1  g268(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  NAND2_X1  g269(.A1(G226gat), .A2(G233gat), .ZN(new_n471));
  XOR2_X1   g270(.A(new_n471), .B(KEYINPUT73), .Z(new_n472));
  XNOR2_X1  g271(.A(KEYINPUT27), .B(G183gat), .ZN(new_n473));
  INV_X1    g272(.A(new_n473), .ZN(new_n474));
  OAI21_X1  g273(.A(KEYINPUT28), .B1(new_n474), .B2(G190gat), .ZN(new_n475));
  NOR3_X1   g274(.A1(KEYINPUT67), .A2(G169gat), .A3(G176gat), .ZN(new_n476));
  AND2_X1   g275(.A1(G169gat), .A2(G176gat), .ZN(new_n477));
  OR3_X1    g276(.A1(new_n476), .A2(KEYINPUT26), .A3(new_n477), .ZN(new_n478));
  AOI22_X1  g277(.A1(new_n476), .A2(KEYINPUT26), .B1(G183gat), .B2(G190gat), .ZN(new_n479));
  INV_X1    g278(.A(KEYINPUT28), .ZN(new_n480));
  INV_X1    g279(.A(G190gat), .ZN(new_n481));
  NAND3_X1  g280(.A1(new_n473), .A2(new_n480), .A3(new_n481), .ZN(new_n482));
  NAND4_X1  g281(.A1(new_n475), .A2(new_n478), .A3(new_n479), .A4(new_n482), .ZN(new_n483));
  INV_X1    g282(.A(new_n483), .ZN(new_n484));
  NOR2_X1   g283(.A1(G169gat), .A2(G176gat), .ZN(new_n485));
  AOI21_X1  g284(.A(new_n477), .B1(KEYINPUT23), .B2(new_n485), .ZN(new_n486));
  NAND2_X1  g285(.A1(G183gat), .A2(G190gat), .ZN(new_n487));
  INV_X1    g286(.A(KEYINPUT24), .ZN(new_n488));
  NAND2_X1  g287(.A1(new_n487), .A2(new_n488), .ZN(new_n489));
  NAND2_X1  g288(.A1(new_n344), .A2(new_n481), .ZN(new_n490));
  NAND3_X1  g289(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n491));
  NAND3_X1  g290(.A1(new_n489), .A2(new_n490), .A3(new_n491), .ZN(new_n492));
  OAI21_X1  g291(.A(KEYINPUT66), .B1(new_n485), .B2(KEYINPUT23), .ZN(new_n493));
  INV_X1    g292(.A(KEYINPUT66), .ZN(new_n494));
  INV_X1    g293(.A(KEYINPUT23), .ZN(new_n495));
  OAI211_X1 g294(.A(new_n494), .B(new_n495), .C1(G169gat), .C2(G176gat), .ZN(new_n496));
  NAND4_X1  g295(.A1(new_n486), .A2(new_n492), .A3(new_n493), .A4(new_n496), .ZN(new_n497));
  INV_X1    g296(.A(KEYINPUT25), .ZN(new_n498));
  INV_X1    g297(.A(KEYINPUT65), .ZN(new_n499));
  NAND4_X1  g298(.A1(new_n486), .A2(new_n499), .A3(new_n493), .A4(new_n496), .ZN(new_n500));
  AOI21_X1  g299(.A(new_n497), .B1(new_n498), .B2(new_n500), .ZN(new_n501));
  INV_X1    g300(.A(new_n501), .ZN(new_n502));
  NAND3_X1  g301(.A1(new_n497), .A2(new_n500), .A3(new_n498), .ZN(new_n503));
  AOI21_X1  g302(.A(new_n484), .B1(new_n502), .B2(new_n503), .ZN(new_n504));
  OAI21_X1  g303(.A(new_n472), .B1(new_n504), .B2(KEYINPUT29), .ZN(new_n505));
  XNOR2_X1  g304(.A(G197gat), .B(G204gat), .ZN(new_n506));
  XNOR2_X1  g305(.A(KEYINPUT72), .B(G218gat), .ZN(new_n507));
  OAI21_X1  g306(.A(new_n506), .B1(new_n507), .B2(KEYINPUT22), .ZN(new_n508));
  NAND2_X1  g307(.A1(new_n508), .A2(G211gat), .ZN(new_n509));
  INV_X1    g308(.A(G211gat), .ZN(new_n510));
  NAND3_X1  g309(.A1(new_n506), .A2(KEYINPUT22), .A3(new_n510), .ZN(new_n511));
  NAND2_X1  g310(.A1(new_n509), .A2(new_n511), .ZN(new_n512));
  NAND2_X1  g311(.A1(new_n512), .A2(G218gat), .ZN(new_n513));
  INV_X1    g312(.A(G218gat), .ZN(new_n514));
  NAND3_X1  g313(.A1(new_n509), .A2(new_n514), .A3(new_n511), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n513), .A2(new_n515), .ZN(new_n516));
  INV_X1    g315(.A(new_n516), .ZN(new_n517));
  INV_X1    g316(.A(new_n503), .ZN(new_n518));
  OAI21_X1  g317(.A(new_n483), .B1(new_n518), .B2(new_n501), .ZN(new_n519));
  INV_X1    g318(.A(KEYINPUT76), .ZN(new_n520));
  XOR2_X1   g319(.A(new_n472), .B(KEYINPUT74), .Z(new_n521));
  AND3_X1   g320(.A1(new_n519), .A2(new_n520), .A3(new_n521), .ZN(new_n522));
  AOI21_X1  g321(.A(new_n520), .B1(new_n519), .B2(new_n521), .ZN(new_n523));
  OAI211_X1 g322(.A(new_n505), .B(new_n517), .C1(new_n522), .C2(new_n523), .ZN(new_n524));
  NOR2_X1   g323(.A1(new_n504), .A2(new_n472), .ZN(new_n525));
  XNOR2_X1  g324(.A(KEYINPUT75), .B(KEYINPUT29), .ZN(new_n526));
  INV_X1    g325(.A(new_n526), .ZN(new_n527));
  AOI21_X1  g326(.A(new_n521), .B1(new_n519), .B2(new_n527), .ZN(new_n528));
  OAI21_X1  g327(.A(new_n516), .B1(new_n525), .B2(new_n528), .ZN(new_n529));
  XNOR2_X1  g328(.A(G8gat), .B(G36gat), .ZN(new_n530));
  XNOR2_X1  g329(.A(new_n530), .B(KEYINPUT77), .ZN(new_n531));
  XNOR2_X1  g330(.A(G64gat), .B(G92gat), .ZN(new_n532));
  XOR2_X1   g331(.A(new_n531), .B(new_n532), .Z(new_n533));
  NAND3_X1  g332(.A1(new_n524), .A2(new_n529), .A3(new_n533), .ZN(new_n534));
  INV_X1    g333(.A(KEYINPUT30), .ZN(new_n535));
  NAND2_X1  g334(.A1(new_n534), .A2(new_n535), .ZN(new_n536));
  NAND2_X1  g335(.A1(new_n524), .A2(new_n529), .ZN(new_n537));
  INV_X1    g336(.A(new_n533), .ZN(new_n538));
  NAND2_X1  g337(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  NAND4_X1  g338(.A1(new_n524), .A2(KEYINPUT30), .A3(new_n529), .A4(new_n533), .ZN(new_n540));
  NAND3_X1  g339(.A1(new_n536), .A2(new_n539), .A3(new_n540), .ZN(new_n541));
  INV_X1    g340(.A(new_n541), .ZN(new_n542));
  NAND2_X1  g341(.A1(new_n470), .A2(new_n542), .ZN(new_n543));
  NAND2_X1  g342(.A1(new_n517), .A2(new_n527), .ZN(new_n544));
  AOI22_X1  g343(.A1(new_n544), .A2(new_n444), .B1(new_n412), .B2(new_n419), .ZN(new_n545));
  AOI21_X1  g344(.A(new_n517), .B1(new_n436), .B2(new_n527), .ZN(new_n546));
  INV_X1    g345(.A(G228gat), .ZN(new_n547));
  INV_X1    g346(.A(G233gat), .ZN(new_n548));
  OAI22_X1  g347(.A1(new_n545), .A2(new_n546), .B1(new_n547), .B2(new_n548), .ZN(new_n549));
  INV_X1    g348(.A(KEYINPUT29), .ZN(new_n550));
  NAND3_X1  g349(.A1(new_n513), .A2(new_n550), .A3(new_n515), .ZN(new_n551));
  AOI22_X1  g350(.A1(new_n444), .A2(new_n551), .B1(new_n445), .B2(new_n446), .ZN(new_n552));
  NAND2_X1  g351(.A1(G228gat), .A2(G233gat), .ZN(new_n553));
  OR3_X1    g352(.A1(new_n546), .A2(new_n552), .A3(new_n553), .ZN(new_n554));
  NAND2_X1  g353(.A1(new_n549), .A2(new_n554), .ZN(new_n555));
  XNOR2_X1  g354(.A(G78gat), .B(G106gat), .ZN(new_n556));
  XNOR2_X1  g355(.A(KEYINPUT31), .B(G50gat), .ZN(new_n557));
  XNOR2_X1  g356(.A(new_n556), .B(new_n557), .ZN(new_n558));
  NOR2_X1   g357(.A1(new_n558), .A2(G22gat), .ZN(new_n559));
  NAND2_X1  g358(.A1(KEYINPUT84), .A2(G22gat), .ZN(new_n560));
  INV_X1    g359(.A(new_n560), .ZN(new_n561));
  AOI21_X1  g360(.A(new_n559), .B1(new_n558), .B2(new_n561), .ZN(new_n562));
  NAND2_X1  g361(.A1(new_n555), .A2(new_n562), .ZN(new_n563));
  INV_X1    g362(.A(new_n562), .ZN(new_n564));
  NAND3_X1  g363(.A1(new_n549), .A2(new_n554), .A3(new_n564), .ZN(new_n565));
  NAND2_X1  g364(.A1(new_n563), .A2(new_n565), .ZN(new_n566));
  NAND2_X1  g365(.A1(new_n519), .A2(new_n438), .ZN(new_n567));
  NAND2_X1  g366(.A1(G227gat), .A2(G233gat), .ZN(new_n568));
  XOR2_X1   g367(.A(new_n568), .B(KEYINPUT64), .Z(new_n569));
  OAI211_X1 g368(.A(new_n434), .B(new_n483), .C1(new_n518), .C2(new_n501), .ZN(new_n570));
  NAND3_X1  g369(.A1(new_n567), .A2(new_n569), .A3(new_n570), .ZN(new_n571));
  INV_X1    g370(.A(KEYINPUT33), .ZN(new_n572));
  XNOR2_X1  g371(.A(G15gat), .B(G43gat), .ZN(new_n573));
  XNOR2_X1  g372(.A(G71gat), .B(G99gat), .ZN(new_n574));
  XOR2_X1   g373(.A(new_n573), .B(new_n574), .Z(new_n575));
  INV_X1    g374(.A(new_n575), .ZN(new_n576));
  OAI211_X1 g375(.A(new_n571), .B(KEYINPUT32), .C1(new_n572), .C2(new_n576), .ZN(new_n577));
  NOR2_X1   g376(.A1(new_n572), .A2(KEYINPUT32), .ZN(new_n578));
  INV_X1    g377(.A(new_n578), .ZN(new_n579));
  NAND2_X1  g378(.A1(new_n571), .A2(new_n579), .ZN(new_n580));
  AOI21_X1  g379(.A(KEYINPUT69), .B1(new_n580), .B2(new_n575), .ZN(new_n581));
  INV_X1    g380(.A(KEYINPUT69), .ZN(new_n582));
  AOI211_X1 g381(.A(new_n582), .B(new_n576), .C1(new_n571), .C2(new_n579), .ZN(new_n583));
  OAI21_X1  g382(.A(new_n577), .B1(new_n581), .B2(new_n583), .ZN(new_n584));
  NAND2_X1  g383(.A1(new_n567), .A2(new_n570), .ZN(new_n585));
  INV_X1    g384(.A(new_n569), .ZN(new_n586));
  NAND2_X1  g385(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  INV_X1    g386(.A(KEYINPUT34), .ZN(new_n588));
  NAND2_X1  g387(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  NAND3_X1  g388(.A1(new_n585), .A2(KEYINPUT34), .A3(new_n586), .ZN(new_n590));
  NAND2_X1  g389(.A1(new_n589), .A2(new_n590), .ZN(new_n591));
  INV_X1    g390(.A(new_n591), .ZN(new_n592));
  NAND2_X1  g391(.A1(new_n584), .A2(new_n592), .ZN(new_n593));
  OAI211_X1 g392(.A(new_n591), .B(new_n577), .C1(new_n581), .C2(new_n583), .ZN(new_n594));
  AND3_X1   g393(.A1(new_n566), .A2(new_n593), .A3(new_n594), .ZN(new_n595));
  INV_X1    g394(.A(new_n595), .ZN(new_n596));
  OAI21_X1  g395(.A(KEYINPUT35), .B1(new_n543), .B2(new_n596), .ZN(new_n597));
  INV_X1    g396(.A(KEYINPUT71), .ZN(new_n598));
  NAND3_X1  g397(.A1(new_n593), .A2(new_n598), .A3(new_n594), .ZN(new_n599));
  OR2_X1    g398(.A1(new_n594), .A2(new_n598), .ZN(new_n600));
  NAND2_X1  g399(.A1(new_n599), .A2(new_n600), .ZN(new_n601));
  NAND2_X1  g400(.A1(new_n601), .A2(KEYINPUT88), .ZN(new_n602));
  INV_X1    g401(.A(new_n566), .ZN(new_n603));
  NOR2_X1   g402(.A1(new_n603), .A2(new_n541), .ZN(new_n604));
  INV_X1    g403(.A(KEYINPUT88), .ZN(new_n605));
  NAND3_X1  g404(.A1(new_n599), .A2(new_n600), .A3(new_n605), .ZN(new_n606));
  NAND3_X1  g405(.A1(new_n602), .A2(new_n604), .A3(new_n606), .ZN(new_n607));
  INV_X1    g406(.A(KEYINPUT87), .ZN(new_n608));
  NAND2_X1  g407(.A1(new_n469), .A2(new_n608), .ZN(new_n609));
  NAND4_X1  g408(.A1(new_n459), .A2(KEYINPUT87), .A3(KEYINPUT6), .A4(new_n463), .ZN(new_n610));
  NAND3_X1  g409(.A1(new_n468), .A2(new_n609), .A3(new_n610), .ZN(new_n611));
  INV_X1    g410(.A(KEYINPUT35), .ZN(new_n612));
  NAND2_X1  g411(.A1(new_n611), .A2(new_n612), .ZN(new_n613));
  OAI21_X1  g412(.A(new_n597), .B1(new_n607), .B2(new_n613), .ZN(new_n614));
  NAND2_X1  g413(.A1(new_n543), .A2(new_n603), .ZN(new_n615));
  NAND3_X1  g414(.A1(new_n593), .A2(KEYINPUT36), .A3(new_n594), .ZN(new_n616));
  XOR2_X1   g415(.A(KEYINPUT70), .B(KEYINPUT36), .Z(new_n617));
  OAI21_X1  g416(.A(new_n616), .B1(new_n601), .B2(new_n617), .ZN(new_n618));
  OAI21_X1  g417(.A(new_n451), .B1(new_n448), .B2(new_n450), .ZN(new_n619));
  OAI21_X1  g418(.A(new_n453), .B1(new_n454), .B2(new_n456), .ZN(new_n620));
  NAND2_X1  g419(.A1(new_n620), .A2(new_n442), .ZN(new_n621));
  NAND3_X1  g420(.A1(new_n619), .A2(KEYINPUT39), .A3(new_n621), .ZN(new_n622));
  INV_X1    g421(.A(KEYINPUT39), .ZN(new_n623));
  OAI211_X1 g422(.A(new_n623), .B(new_n451), .C1(new_n448), .C2(new_n450), .ZN(new_n624));
  INV_X1    g423(.A(KEYINPUT85), .ZN(new_n625));
  AND3_X1   g424(.A1(new_n624), .A2(new_n625), .A3(new_n466), .ZN(new_n626));
  AOI21_X1  g425(.A(new_n625), .B1(new_n624), .B2(new_n466), .ZN(new_n627));
  OAI21_X1  g426(.A(new_n622), .B1(new_n626), .B2(new_n627), .ZN(new_n628));
  INV_X1    g427(.A(KEYINPUT40), .ZN(new_n629));
  NAND2_X1  g428(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  AND2_X1   g429(.A1(new_n464), .A2(new_n541), .ZN(new_n631));
  OAI211_X1 g430(.A(new_n622), .B(KEYINPUT40), .C1(new_n626), .C2(new_n627), .ZN(new_n632));
  NAND3_X1  g431(.A1(new_n630), .A2(new_n631), .A3(new_n632), .ZN(new_n633));
  NAND2_X1  g432(.A1(new_n633), .A2(new_n566), .ZN(new_n634));
  NAND2_X1  g433(.A1(new_n538), .A2(KEYINPUT37), .ZN(new_n635));
  NAND2_X1  g434(.A1(new_n539), .A2(new_n635), .ZN(new_n636));
  XOR2_X1   g435(.A(KEYINPUT86), .B(KEYINPUT38), .Z(new_n637));
  OAI21_X1  g436(.A(new_n517), .B1(new_n525), .B2(new_n528), .ZN(new_n638));
  OAI21_X1  g437(.A(new_n505), .B1(new_n522), .B2(new_n523), .ZN(new_n639));
  OAI211_X1 g438(.A(KEYINPUT37), .B(new_n638), .C1(new_n639), .C2(new_n517), .ZN(new_n640));
  NAND3_X1  g439(.A1(new_n636), .A2(new_n637), .A3(new_n640), .ZN(new_n641));
  AOI22_X1  g440(.A1(new_n539), .A2(new_n635), .B1(KEYINPUT37), .B2(new_n537), .ZN(new_n642));
  OAI211_X1 g441(.A(new_n641), .B(new_n534), .C1(new_n637), .C2(new_n642), .ZN(new_n643));
  NOR2_X1   g442(.A1(new_n611), .A2(new_n643), .ZN(new_n644));
  OAI211_X1 g443(.A(new_n615), .B(new_n618), .C1(new_n634), .C2(new_n644), .ZN(new_n645));
  AOI211_X1 g444(.A(new_n337), .B(new_n388), .C1(new_n614), .C2(new_n645), .ZN(new_n646));
  INV_X1    g445(.A(new_n470), .ZN(new_n647));
  NAND2_X1  g446(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  XNOR2_X1  g447(.A(new_n648), .B(G1gat), .ZN(G1324gat));
  AOI21_X1  g448(.A(new_n205), .B1(new_n646), .B2(new_n541), .ZN(new_n650));
  XNOR2_X1  g449(.A(new_n650), .B(KEYINPUT100), .ZN(new_n651));
  XOR2_X1   g450(.A(KEYINPUT16), .B(G8gat), .Z(new_n652));
  NAND3_X1  g451(.A1(new_n646), .A2(new_n541), .A3(new_n652), .ZN(new_n653));
  AND2_X1   g452(.A1(new_n653), .A2(KEYINPUT42), .ZN(new_n654));
  NOR2_X1   g453(.A1(new_n653), .A2(KEYINPUT42), .ZN(new_n655));
  OAI21_X1  g454(.A(new_n651), .B1(new_n654), .B2(new_n655), .ZN(G1325gat));
  AND2_X1   g455(.A1(new_n602), .A2(new_n606), .ZN(new_n657));
  AOI21_X1  g456(.A(G15gat), .B1(new_n646), .B2(new_n657), .ZN(new_n658));
  INV_X1    g457(.A(G15gat), .ZN(new_n659));
  NOR2_X1   g458(.A1(new_n618), .A2(new_n659), .ZN(new_n660));
  XNOR2_X1  g459(.A(new_n660), .B(KEYINPUT101), .ZN(new_n661));
  AOI21_X1  g460(.A(new_n658), .B1(new_n646), .B2(new_n661), .ZN(G1326gat));
  NAND2_X1  g461(.A1(new_n646), .A2(new_n603), .ZN(new_n663));
  XNOR2_X1  g462(.A(KEYINPUT43), .B(G22gat), .ZN(new_n664));
  XNOR2_X1  g463(.A(new_n663), .B(new_n664), .ZN(G1327gat));
  NAND2_X1  g464(.A1(new_n614), .A2(new_n645), .ZN(new_n666));
  NAND2_X1  g465(.A1(new_n666), .A2(new_n386), .ZN(new_n667));
  NOR3_X1   g466(.A1(new_n667), .A2(new_n337), .A3(new_n366), .ZN(new_n668));
  NAND3_X1  g467(.A1(new_n668), .A2(new_n212), .A3(new_n647), .ZN(new_n669));
  XNOR2_X1  g468(.A(new_n669), .B(KEYINPUT45), .ZN(new_n670));
  INV_X1    g469(.A(KEYINPUT104), .ZN(new_n671));
  NAND3_X1  g470(.A1(new_n614), .A2(new_n645), .A3(new_n671), .ZN(new_n672));
  INV_X1    g471(.A(new_n672), .ZN(new_n673));
  AOI21_X1  g472(.A(new_n671), .B1(new_n614), .B2(new_n645), .ZN(new_n674));
  NOR2_X1   g473(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  OAI21_X1  g474(.A(KEYINPUT105), .B1(new_n383), .B2(new_n385), .ZN(new_n676));
  INV_X1    g475(.A(new_n379), .ZN(new_n677));
  INV_X1    g476(.A(new_n382), .ZN(new_n678));
  NAND3_X1  g477(.A1(new_n677), .A2(new_n678), .A3(new_n377), .ZN(new_n679));
  INV_X1    g478(.A(KEYINPUT105), .ZN(new_n680));
  NAND3_X1  g479(.A1(new_n679), .A2(new_n680), .A3(new_n384), .ZN(new_n681));
  NAND2_X1  g480(.A1(new_n676), .A2(new_n681), .ZN(new_n682));
  INV_X1    g481(.A(KEYINPUT44), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  AOI21_X1  g483(.A(new_n387), .B1(new_n614), .B2(new_n645), .ZN(new_n685));
  OAI22_X1  g484(.A1(new_n675), .A2(new_n684), .B1(new_n683), .B2(new_n685), .ZN(new_n686));
  AND3_X1   g485(.A1(new_n364), .A2(KEYINPUT102), .A3(new_n365), .ZN(new_n687));
  AOI21_X1  g486(.A(KEYINPUT102), .B1(new_n364), .B2(new_n365), .ZN(new_n688));
  NOR2_X1   g487(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  NAND2_X1  g488(.A1(new_n689), .A2(new_n336), .ZN(new_n690));
  XOR2_X1   g489(.A(new_n690), .B(KEYINPUT103), .Z(new_n691));
  NAND2_X1  g490(.A1(new_n686), .A2(new_n691), .ZN(new_n692));
  OAI21_X1  g491(.A(G29gat), .B1(new_n692), .B2(new_n470), .ZN(new_n693));
  NAND2_X1  g492(.A1(new_n670), .A2(new_n693), .ZN(G1328gat));
  NAND3_X1  g493(.A1(new_n668), .A2(new_n213), .A3(new_n541), .ZN(new_n695));
  XOR2_X1   g494(.A(new_n695), .B(KEYINPUT46), .Z(new_n696));
  OAI21_X1  g495(.A(G36gat), .B1(new_n692), .B2(new_n542), .ZN(new_n697));
  NAND2_X1  g496(.A1(new_n696), .A2(new_n697), .ZN(G1329gat));
  INV_X1    g497(.A(G43gat), .ZN(new_n699));
  INV_X1    g498(.A(new_n668), .ZN(new_n700));
  INV_X1    g499(.A(new_n657), .ZN(new_n701));
  OAI21_X1  g500(.A(new_n699), .B1(new_n700), .B2(new_n701), .ZN(new_n702));
  NAND3_X1  g501(.A1(new_n686), .A2(G43gat), .A3(new_n691), .ZN(new_n703));
  OAI21_X1  g502(.A(new_n702), .B1(new_n703), .B2(new_n618), .ZN(new_n704));
  XNOR2_X1  g503(.A(new_n704), .B(KEYINPUT47), .ZN(G1330gat));
  INV_X1    g504(.A(KEYINPUT106), .ZN(new_n706));
  NAND4_X1  g505(.A1(new_n686), .A2(new_n706), .A3(new_n603), .A4(new_n691), .ZN(new_n707));
  NAND2_X1  g506(.A1(new_n666), .A2(KEYINPUT104), .ZN(new_n708));
  AOI21_X1  g507(.A(new_n684), .B1(new_n708), .B2(new_n672), .ZN(new_n709));
  NOR2_X1   g508(.A1(new_n685), .A2(new_n683), .ZN(new_n710));
  OAI211_X1 g509(.A(new_n603), .B(new_n691), .C1(new_n709), .C2(new_n710), .ZN(new_n711));
  NAND2_X1  g510(.A1(new_n711), .A2(KEYINPUT106), .ZN(new_n712));
  NAND3_X1  g511(.A1(new_n707), .A2(new_n712), .A3(G50gat), .ZN(new_n713));
  NOR3_X1   g512(.A1(new_n700), .A2(G50gat), .A3(new_n566), .ZN(new_n714));
  INV_X1    g513(.A(new_n714), .ZN(new_n715));
  NAND3_X1  g514(.A1(new_n713), .A2(KEYINPUT48), .A3(new_n715), .ZN(new_n716));
  AOI21_X1  g515(.A(new_n714), .B1(new_n711), .B2(G50gat), .ZN(new_n717));
  OAI21_X1  g516(.A(new_n716), .B1(KEYINPUT48), .B2(new_n717), .ZN(G1331gat));
  NAND2_X1  g517(.A1(new_n708), .A2(new_n672), .ZN(new_n719));
  INV_X1    g518(.A(new_n388), .ZN(new_n720));
  INV_X1    g519(.A(new_n335), .ZN(new_n721));
  NOR2_X1   g520(.A1(new_n262), .A2(new_n721), .ZN(new_n722));
  NAND3_X1  g521(.A1(new_n719), .A2(new_n720), .A3(new_n722), .ZN(new_n723));
  NOR2_X1   g522(.A1(new_n723), .A2(new_n470), .ZN(new_n724));
  XOR2_X1   g523(.A(new_n724), .B(G57gat), .Z(G1332gat));
  NOR2_X1   g524(.A1(new_n723), .A2(new_n542), .ZN(new_n726));
  NOR2_X1   g525(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n727));
  AND2_X1   g526(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n728));
  OAI21_X1  g527(.A(new_n726), .B1(new_n727), .B2(new_n728), .ZN(new_n729));
  OAI21_X1  g528(.A(new_n729), .B1(new_n726), .B2(new_n727), .ZN(G1333gat));
  XNOR2_X1  g529(.A(new_n657), .B(KEYINPUT107), .ZN(new_n731));
  OAI21_X1  g530(.A(new_n288), .B1(new_n723), .B2(new_n731), .ZN(new_n732));
  OR2_X1    g531(.A1(new_n618), .A2(new_n288), .ZN(new_n733));
  OAI21_X1  g532(.A(new_n732), .B1(new_n723), .B2(new_n733), .ZN(new_n734));
  XNOR2_X1  g533(.A(new_n734), .B(KEYINPUT50), .ZN(G1334gat));
  NOR2_X1   g534(.A1(new_n723), .A2(new_n566), .ZN(new_n736));
  XNOR2_X1  g535(.A(new_n736), .B(new_n289), .ZN(G1335gat));
  NOR3_X1   g536(.A1(new_n366), .A2(new_n262), .A3(new_n721), .ZN(new_n738));
  NAND2_X1  g537(.A1(new_n686), .A2(new_n738), .ZN(new_n739));
  NOR3_X1   g538(.A1(new_n739), .A2(new_n276), .A3(new_n470), .ZN(new_n740));
  NAND3_X1  g539(.A1(new_n666), .A2(KEYINPUT108), .A3(new_n386), .ZN(new_n741));
  NAND2_X1  g540(.A1(new_n741), .A2(new_n263), .ZN(new_n742));
  AND2_X1   g541(.A1(new_n364), .A2(new_n365), .ZN(new_n743));
  OAI21_X1  g542(.A(new_n743), .B1(new_n685), .B2(KEYINPUT108), .ZN(new_n744));
  OAI21_X1  g543(.A(KEYINPUT51), .B1(new_n742), .B2(new_n744), .ZN(new_n745));
  INV_X1    g544(.A(KEYINPUT108), .ZN(new_n746));
  NAND2_X1  g545(.A1(new_n667), .A2(new_n746), .ZN(new_n747));
  AOI21_X1  g546(.A(new_n262), .B1(new_n685), .B2(KEYINPUT108), .ZN(new_n748));
  INV_X1    g547(.A(KEYINPUT51), .ZN(new_n749));
  NAND4_X1  g548(.A1(new_n747), .A2(new_n748), .A3(new_n749), .A4(new_n743), .ZN(new_n750));
  NAND4_X1  g549(.A1(new_n745), .A2(new_n750), .A3(new_n647), .A4(new_n335), .ZN(new_n751));
  AOI21_X1  g550(.A(new_n740), .B1(new_n276), .B2(new_n751), .ZN(G1336gat));
  OAI211_X1 g551(.A(new_n541), .B(new_n738), .C1(new_n709), .C2(new_n710), .ZN(new_n753));
  NAND2_X1  g552(.A1(new_n753), .A2(G92gat), .ZN(new_n754));
  NAND4_X1  g553(.A1(new_n745), .A2(new_n750), .A3(new_n335), .A4(new_n541), .ZN(new_n755));
  OAI21_X1  g554(.A(new_n754), .B1(new_n755), .B2(G92gat), .ZN(new_n756));
  NAND2_X1  g555(.A1(new_n756), .A2(KEYINPUT52), .ZN(new_n757));
  INV_X1    g556(.A(KEYINPUT52), .ZN(new_n758));
  OAI211_X1 g557(.A(new_n754), .B(new_n758), .C1(new_n755), .C2(G92gat), .ZN(new_n759));
  NAND2_X1  g558(.A1(new_n757), .A2(new_n759), .ZN(G1337gat));
  OAI21_X1  g559(.A(G99gat), .B1(new_n739), .B2(new_n618), .ZN(new_n761));
  INV_X1    g560(.A(G99gat), .ZN(new_n762));
  NAND4_X1  g561(.A1(new_n745), .A2(new_n750), .A3(new_n762), .A4(new_n335), .ZN(new_n763));
  OAI21_X1  g562(.A(new_n761), .B1(new_n701), .B2(new_n763), .ZN(G1338gat));
  NAND4_X1  g563(.A1(new_n745), .A2(new_n750), .A3(new_n335), .A4(new_n603), .ZN(new_n765));
  INV_X1    g564(.A(G106gat), .ZN(new_n766));
  NAND2_X1  g565(.A1(new_n765), .A2(new_n766), .ZN(new_n767));
  NAND4_X1  g566(.A1(new_n686), .A2(G106gat), .A3(new_n603), .A4(new_n738), .ZN(new_n768));
  NAND2_X1  g567(.A1(new_n767), .A2(new_n768), .ZN(new_n769));
  XNOR2_X1  g568(.A(KEYINPUT109), .B(KEYINPUT53), .ZN(new_n770));
  INV_X1    g569(.A(new_n770), .ZN(new_n771));
  NAND2_X1  g570(.A1(new_n769), .A2(new_n771), .ZN(new_n772));
  NAND3_X1  g571(.A1(new_n767), .A2(new_n768), .A3(new_n770), .ZN(new_n773));
  NAND2_X1  g572(.A1(new_n772), .A2(new_n773), .ZN(G1339gat));
  INV_X1    g573(.A(new_n331), .ZN(new_n775));
  NAND3_X1  g574(.A1(new_n323), .A2(new_n321), .A3(new_n330), .ZN(new_n776));
  NAND3_X1  g575(.A1(new_n775), .A2(KEYINPUT54), .A3(new_n776), .ZN(new_n777));
  INV_X1    g576(.A(KEYINPUT54), .ZN(new_n778));
  AOI211_X1 g577(.A(KEYINPUT110), .B(new_n319), .C1(new_n331), .C2(new_n778), .ZN(new_n779));
  INV_X1    g578(.A(KEYINPUT110), .ZN(new_n780));
  NAND2_X1  g579(.A1(new_n367), .A2(new_n338), .ZN(new_n781));
  NAND3_X1  g580(.A1(new_n285), .A2(new_n286), .A3(new_n305), .ZN(new_n782));
  AOI21_X1  g581(.A(KEYINPUT10), .B1(new_n781), .B2(new_n782), .ZN(new_n783));
  NAND3_X1  g582(.A1(new_n329), .A2(new_n325), .A3(KEYINPUT10), .ZN(new_n784));
  NOR2_X1   g583(.A1(new_n784), .A2(new_n367), .ZN(new_n785));
  OAI211_X1 g584(.A(new_n778), .B(new_n313), .C1(new_n783), .C2(new_n785), .ZN(new_n786));
  AOI21_X1  g585(.A(new_n780), .B1(new_n786), .B2(new_n318), .ZN(new_n787));
  OAI211_X1 g586(.A(KEYINPUT55), .B(new_n777), .C1(new_n779), .C2(new_n787), .ZN(new_n788));
  NAND2_X1  g587(.A1(new_n788), .A2(new_n333), .ZN(new_n789));
  INV_X1    g588(.A(KEYINPUT111), .ZN(new_n790));
  NAND2_X1  g589(.A1(new_n789), .A2(new_n790), .ZN(new_n791));
  OAI21_X1  g590(.A(new_n777), .B1(new_n779), .B2(new_n787), .ZN(new_n792));
  INV_X1    g591(.A(KEYINPUT55), .ZN(new_n793));
  NAND2_X1  g592(.A1(new_n792), .A2(new_n793), .ZN(new_n794));
  NAND3_X1  g593(.A1(new_n788), .A2(KEYINPUT111), .A3(new_n333), .ZN(new_n795));
  NAND4_X1  g594(.A1(new_n791), .A2(new_n262), .A3(new_n794), .A4(new_n795), .ZN(new_n796));
  NOR2_X1   g595(.A1(new_n237), .A2(new_n239), .ZN(new_n797));
  NOR2_X1   g596(.A1(new_n250), .A2(new_n238), .ZN(new_n798));
  OAI21_X1  g597(.A(new_n257), .B1(new_n797), .B2(new_n798), .ZN(new_n799));
  AND2_X1   g598(.A1(new_n261), .A2(new_n799), .ZN(new_n800));
  NAND2_X1  g599(.A1(new_n800), .A2(new_n335), .ZN(new_n801));
  AOI21_X1  g600(.A(new_n682), .B1(new_n796), .B2(new_n801), .ZN(new_n802));
  NAND4_X1  g601(.A1(new_n791), .A2(new_n794), .A3(new_n795), .A4(new_n800), .ZN(new_n803));
  NOR3_X1   g602(.A1(new_n383), .A2(new_n385), .A3(KEYINPUT105), .ZN(new_n804));
  AOI21_X1  g603(.A(new_n680), .B1(new_n679), .B2(new_n384), .ZN(new_n805));
  NOR2_X1   g604(.A1(new_n804), .A2(new_n805), .ZN(new_n806));
  NOR2_X1   g605(.A1(new_n803), .A2(new_n806), .ZN(new_n807));
  OAI21_X1  g606(.A(new_n689), .B1(new_n802), .B2(new_n807), .ZN(new_n808));
  NAND3_X1  g607(.A1(new_n720), .A2(new_n263), .A3(new_n721), .ZN(new_n809));
  AOI21_X1  g608(.A(new_n470), .B1(new_n808), .B2(new_n809), .ZN(new_n810));
  INV_X1    g609(.A(new_n810), .ZN(new_n811));
  NOR2_X1   g610(.A1(new_n811), .A2(new_n607), .ZN(new_n812));
  INV_X1    g611(.A(new_n812), .ZN(new_n813));
  OAI21_X1  g612(.A(G113gat), .B1(new_n813), .B2(new_n263), .ZN(new_n814));
  NAND3_X1  g613(.A1(new_n810), .A2(new_n542), .A3(new_n595), .ZN(new_n815));
  INV_X1    g614(.A(new_n815), .ZN(new_n816));
  NAND3_X1  g615(.A1(new_n816), .A2(new_n427), .A3(new_n262), .ZN(new_n817));
  NAND2_X1  g616(.A1(new_n814), .A2(new_n817), .ZN(G1340gat));
  OAI21_X1  g617(.A(G120gat), .B1(new_n813), .B2(new_n721), .ZN(new_n819));
  OR2_X1    g618(.A1(new_n721), .A2(new_n426), .ZN(new_n820));
  OAI21_X1  g619(.A(new_n819), .B1(new_n815), .B2(new_n820), .ZN(G1341gat));
  AOI21_X1  g620(.A(G127gat), .B1(new_n816), .B2(new_n366), .ZN(new_n822));
  NOR2_X1   g621(.A1(new_n813), .A2(new_n689), .ZN(new_n823));
  AOI21_X1  g622(.A(new_n822), .B1(new_n823), .B2(G127gat), .ZN(G1342gat));
  NOR3_X1   g623(.A1(new_n815), .A2(G134gat), .A3(new_n387), .ZN(new_n825));
  XNOR2_X1  g624(.A(new_n825), .B(KEYINPUT56), .ZN(new_n826));
  OAI21_X1  g625(.A(G134gat), .B1(new_n813), .B2(new_n387), .ZN(new_n827));
  NAND2_X1  g626(.A1(new_n826), .A2(new_n827), .ZN(G1343gat));
  NOR2_X1   g627(.A1(new_n401), .A2(new_n391), .ZN(new_n829));
  INV_X1    g628(.A(new_n829), .ZN(new_n830));
  NAND3_X1  g629(.A1(new_n618), .A2(new_n647), .A3(new_n542), .ZN(new_n831));
  INV_X1    g630(.A(KEYINPUT112), .ZN(new_n832));
  NAND2_X1  g631(.A1(new_n776), .A2(KEYINPUT54), .ZN(new_n833));
  NOR2_X1   g632(.A1(new_n833), .A2(new_n331), .ZN(new_n834));
  AOI211_X1 g633(.A(KEYINPUT54), .B(new_n321), .C1(new_n323), .C2(new_n330), .ZN(new_n835));
  OAI21_X1  g634(.A(KEYINPUT110), .B1(new_n835), .B2(new_n319), .ZN(new_n836));
  NAND3_X1  g635(.A1(new_n786), .A2(new_n780), .A3(new_n318), .ZN(new_n837));
  AOI21_X1  g636(.A(new_n834), .B1(new_n836), .B2(new_n837), .ZN(new_n838));
  OAI21_X1  g637(.A(new_n832), .B1(new_n838), .B2(KEYINPUT55), .ZN(new_n839));
  AOI21_X1  g638(.A(new_n332), .B1(new_n838), .B2(KEYINPUT55), .ZN(new_n840));
  NAND3_X1  g639(.A1(new_n792), .A2(KEYINPUT112), .A3(new_n793), .ZN(new_n841));
  NAND4_X1  g640(.A1(new_n839), .A2(new_n840), .A3(new_n262), .A4(new_n841), .ZN(new_n842));
  AOI21_X1  g641(.A(new_n386), .B1(new_n842), .B2(new_n801), .ZN(new_n843));
  OAI21_X1  g642(.A(new_n743), .B1(new_n807), .B2(new_n843), .ZN(new_n844));
  NAND2_X1  g643(.A1(new_n844), .A2(new_n809), .ZN(new_n845));
  INV_X1    g644(.A(KEYINPUT57), .ZN(new_n846));
  NOR2_X1   g645(.A1(new_n566), .A2(new_n846), .ZN(new_n847));
  AOI21_X1  g646(.A(KEYINPUT113), .B1(new_n845), .B2(new_n847), .ZN(new_n848));
  INV_X1    g647(.A(KEYINPUT113), .ZN(new_n849));
  INV_X1    g648(.A(new_n847), .ZN(new_n850));
  AOI211_X1 g649(.A(new_n849), .B(new_n850), .C1(new_n844), .C2(new_n809), .ZN(new_n851));
  NOR2_X1   g650(.A1(new_n848), .A2(new_n851), .ZN(new_n852));
  NAND2_X1  g651(.A1(new_n808), .A2(new_n809), .ZN(new_n853));
  NAND2_X1  g652(.A1(new_n853), .A2(new_n603), .ZN(new_n854));
  NAND2_X1  g653(.A1(new_n854), .A2(new_n846), .ZN(new_n855));
  AOI21_X1  g654(.A(new_n831), .B1(new_n852), .B2(new_n855), .ZN(new_n856));
  AOI21_X1  g655(.A(new_n830), .B1(new_n856), .B2(new_n262), .ZN(new_n857));
  AND2_X1   g656(.A1(new_n618), .A2(new_n603), .ZN(new_n858));
  NAND2_X1  g657(.A1(new_n858), .A2(KEYINPUT114), .ZN(new_n859));
  OR2_X1    g658(.A1(new_n858), .A2(KEYINPUT114), .ZN(new_n860));
  NAND4_X1  g659(.A1(new_n853), .A2(new_n647), .A3(new_n859), .A4(new_n860), .ZN(new_n861));
  NOR4_X1   g660(.A1(new_n861), .A2(G141gat), .A3(new_n263), .A4(new_n541), .ZN(new_n862));
  OAI211_X1 g661(.A(KEYINPUT115), .B(KEYINPUT58), .C1(new_n857), .C2(new_n862), .ZN(new_n863));
  INV_X1    g662(.A(KEYINPUT115), .ZN(new_n864));
  INV_X1    g663(.A(new_n831), .ZN(new_n865));
  NAND2_X1  g664(.A1(new_n842), .A2(new_n801), .ZN(new_n866));
  NAND2_X1  g665(.A1(new_n866), .A2(new_n387), .ZN(new_n867));
  AND3_X1   g666(.A1(new_n788), .A2(KEYINPUT111), .A3(new_n333), .ZN(new_n868));
  AOI21_X1  g667(.A(KEYINPUT111), .B1(new_n788), .B2(new_n333), .ZN(new_n869));
  NOR2_X1   g668(.A1(new_n868), .A2(new_n869), .ZN(new_n870));
  NAND4_X1  g669(.A1(new_n870), .A2(new_n682), .A3(new_n794), .A4(new_n800), .ZN(new_n871));
  AOI21_X1  g670(.A(new_n366), .B1(new_n867), .B2(new_n871), .ZN(new_n872));
  NOR3_X1   g671(.A1(new_n388), .A2(new_n262), .A3(new_n335), .ZN(new_n873));
  OAI21_X1  g672(.A(new_n847), .B1(new_n872), .B2(new_n873), .ZN(new_n874));
  NAND2_X1  g673(.A1(new_n874), .A2(new_n849), .ZN(new_n875));
  NAND3_X1  g674(.A1(new_n845), .A2(KEYINPUT113), .A3(new_n847), .ZN(new_n876));
  NAND2_X1  g675(.A1(new_n875), .A2(new_n876), .ZN(new_n877));
  AOI21_X1  g676(.A(new_n566), .B1(new_n808), .B2(new_n809), .ZN(new_n878));
  NOR2_X1   g677(.A1(new_n878), .A2(KEYINPUT57), .ZN(new_n879));
  OAI211_X1 g678(.A(new_n262), .B(new_n865), .C1(new_n877), .C2(new_n879), .ZN(new_n880));
  AOI21_X1  g679(.A(new_n862), .B1(new_n880), .B2(new_n829), .ZN(new_n881));
  INV_X1    g680(.A(KEYINPUT58), .ZN(new_n882));
  OAI21_X1  g681(.A(new_n864), .B1(new_n881), .B2(new_n882), .ZN(new_n883));
  INV_X1    g682(.A(KEYINPUT116), .ZN(new_n884));
  NAND2_X1  g683(.A1(new_n861), .A2(new_n884), .ZN(new_n885));
  NOR2_X1   g684(.A1(new_n263), .A2(G141gat), .ZN(new_n886));
  NAND4_X1  g685(.A1(new_n810), .A2(KEYINPUT116), .A3(new_n859), .A4(new_n860), .ZN(new_n887));
  NAND4_X1  g686(.A1(new_n885), .A2(new_n542), .A3(new_n886), .A4(new_n887), .ZN(new_n888));
  OR2_X1    g687(.A1(new_n888), .A2(KEYINPUT117), .ZN(new_n889));
  AOI21_X1  g688(.A(KEYINPUT58), .B1(new_n880), .B2(new_n829), .ZN(new_n890));
  NAND2_X1  g689(.A1(new_n888), .A2(KEYINPUT117), .ZN(new_n891));
  NAND3_X1  g690(.A1(new_n889), .A2(new_n890), .A3(new_n891), .ZN(new_n892));
  NAND3_X1  g691(.A1(new_n863), .A2(new_n883), .A3(new_n892), .ZN(G1344gat));
  AND3_X1   g692(.A1(new_n885), .A2(new_n542), .A3(new_n887), .ZN(new_n894));
  INV_X1    g693(.A(new_n404), .ZN(new_n895));
  NAND3_X1  g694(.A1(new_n894), .A2(new_n895), .A3(new_n335), .ZN(new_n896));
  NOR2_X1   g695(.A1(new_n803), .A2(new_n387), .ZN(new_n897));
  OAI21_X1  g696(.A(new_n743), .B1(new_n897), .B2(new_n843), .ZN(new_n898));
  AOI21_X1  g697(.A(KEYINPUT57), .B1(new_n898), .B2(new_n809), .ZN(new_n899));
  AOI22_X1  g698(.A1(new_n854), .A2(KEYINPUT57), .B1(new_n603), .B2(new_n899), .ZN(new_n900));
  INV_X1    g699(.A(KEYINPUT119), .ZN(new_n901));
  NAND4_X1  g700(.A1(new_n900), .A2(new_n901), .A3(new_n335), .A4(new_n865), .ZN(new_n902));
  NAND4_X1  g701(.A1(new_n870), .A2(new_n386), .A3(new_n794), .A4(new_n800), .ZN(new_n903));
  AOI21_X1  g702(.A(new_n366), .B1(new_n867), .B2(new_n903), .ZN(new_n904));
  OAI211_X1 g703(.A(new_n846), .B(new_n603), .C1(new_n904), .C2(new_n873), .ZN(new_n905));
  OAI211_X1 g704(.A(new_n905), .B(new_n865), .C1(new_n878), .C2(new_n846), .ZN(new_n906));
  OAI21_X1  g705(.A(KEYINPUT119), .B1(new_n906), .B2(new_n721), .ZN(new_n907));
  NAND3_X1  g706(.A1(new_n902), .A2(G148gat), .A3(new_n907), .ZN(new_n908));
  XNOR2_X1  g707(.A(KEYINPUT118), .B(KEYINPUT59), .ZN(new_n909));
  AND2_X1   g708(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  AOI211_X1 g709(.A(KEYINPUT59), .B(new_n895), .C1(new_n856), .C2(new_n335), .ZN(new_n911));
  OAI21_X1  g710(.A(new_n896), .B1(new_n910), .B2(new_n911), .ZN(G1345gat));
  AOI21_X1  g711(.A(G155gat), .B1(new_n894), .B2(new_n366), .ZN(new_n913));
  INV_X1    g712(.A(G155gat), .ZN(new_n914));
  NOR2_X1   g713(.A1(new_n689), .A2(new_n914), .ZN(new_n915));
  XNOR2_X1  g714(.A(new_n915), .B(KEYINPUT120), .ZN(new_n916));
  AOI21_X1  g715(.A(new_n913), .B1(new_n856), .B2(new_n916), .ZN(G1346gat));
  OAI21_X1  g716(.A(new_n865), .B1(new_n877), .B2(new_n879), .ZN(new_n918));
  OAI21_X1  g717(.A(G162gat), .B1(new_n918), .B2(new_n806), .ZN(new_n919));
  INV_X1    g718(.A(KEYINPUT121), .ZN(new_n920));
  NAND4_X1  g719(.A1(new_n885), .A2(new_n542), .A3(new_n386), .A4(new_n887), .ZN(new_n921));
  OAI211_X1 g720(.A(new_n919), .B(new_n920), .C1(G162gat), .C2(new_n921), .ZN(new_n922));
  INV_X1    g721(.A(G162gat), .ZN(new_n923));
  AOI21_X1  g722(.A(new_n923), .B1(new_n856), .B2(new_n682), .ZN(new_n924));
  NOR2_X1   g723(.A1(new_n921), .A2(G162gat), .ZN(new_n925));
  OAI21_X1  g724(.A(KEYINPUT121), .B1(new_n924), .B2(new_n925), .ZN(new_n926));
  NAND2_X1  g725(.A1(new_n922), .A2(new_n926), .ZN(G1347gat));
  NOR2_X1   g726(.A1(new_n647), .A2(new_n542), .ZN(new_n928));
  NAND2_X1  g727(.A1(new_n853), .A2(new_n928), .ZN(new_n929));
  NOR3_X1   g728(.A1(new_n929), .A2(new_n603), .A3(new_n731), .ZN(new_n930));
  INV_X1    g729(.A(new_n930), .ZN(new_n931));
  OAI21_X1  g730(.A(G169gat), .B1(new_n931), .B2(new_n263), .ZN(new_n932));
  AND2_X1   g731(.A1(new_n853), .A2(new_n928), .ZN(new_n933));
  NAND2_X1  g732(.A1(new_n933), .A2(new_n595), .ZN(new_n934));
  INV_X1    g733(.A(new_n934), .ZN(new_n935));
  INV_X1    g734(.A(G169gat), .ZN(new_n936));
  NAND3_X1  g735(.A1(new_n935), .A2(new_n936), .A3(new_n262), .ZN(new_n937));
  NAND2_X1  g736(.A1(new_n932), .A2(new_n937), .ZN(G1348gat));
  AOI21_X1  g737(.A(G176gat), .B1(new_n935), .B2(new_n335), .ZN(new_n939));
  NOR2_X1   g738(.A1(new_n931), .A2(new_n721), .ZN(new_n940));
  AOI21_X1  g739(.A(new_n939), .B1(G176gat), .B2(new_n940), .ZN(G1349gat));
  NOR3_X1   g740(.A1(new_n934), .A2(new_n474), .A3(new_n743), .ZN(new_n942));
  INV_X1    g741(.A(new_n689), .ZN(new_n943));
  AOI21_X1  g742(.A(new_n344), .B1(new_n930), .B2(new_n943), .ZN(new_n944));
  NOR2_X1   g743(.A1(new_n942), .A2(new_n944), .ZN(new_n945));
  INV_X1    g744(.A(KEYINPUT60), .ZN(new_n946));
  XNOR2_X1  g745(.A(new_n945), .B(new_n946), .ZN(G1350gat));
  NAND3_X1  g746(.A1(new_n935), .A2(new_n481), .A3(new_n682), .ZN(new_n948));
  OAI21_X1  g747(.A(G190gat), .B1(new_n931), .B2(new_n387), .ZN(new_n949));
  AND2_X1   g748(.A1(new_n949), .A2(KEYINPUT61), .ZN(new_n950));
  NOR2_X1   g749(.A1(new_n949), .A2(KEYINPUT61), .ZN(new_n951));
  OAI21_X1  g750(.A(new_n948), .B1(new_n950), .B2(new_n951), .ZN(G1351gat));
  NAND2_X1  g751(.A1(new_n928), .A2(new_n618), .ZN(new_n953));
  XNOR2_X1  g752(.A(new_n953), .B(KEYINPUT124), .ZN(new_n954));
  OR2_X1    g753(.A1(new_n954), .A2(KEYINPUT125), .ZN(new_n955));
  NAND2_X1  g754(.A1(new_n954), .A2(KEYINPUT125), .ZN(new_n956));
  NAND3_X1  g755(.A1(new_n900), .A2(new_n955), .A3(new_n956), .ZN(new_n957));
  OAI21_X1  g756(.A(G197gat), .B1(new_n957), .B2(new_n263), .ZN(new_n958));
  NAND2_X1  g757(.A1(new_n933), .A2(new_n858), .ZN(new_n959));
  NAND2_X1  g758(.A1(new_n959), .A2(KEYINPUT122), .ZN(new_n960));
  INV_X1    g759(.A(KEYINPUT122), .ZN(new_n961));
  NAND3_X1  g760(.A1(new_n933), .A2(new_n961), .A3(new_n858), .ZN(new_n962));
  NAND4_X1  g761(.A1(new_n960), .A2(new_n254), .A3(new_n262), .A4(new_n962), .ZN(new_n963));
  AND2_X1   g762(.A1(new_n963), .A2(KEYINPUT123), .ZN(new_n964));
  NOR2_X1   g763(.A1(new_n963), .A2(KEYINPUT123), .ZN(new_n965));
  OAI21_X1  g764(.A(new_n958), .B1(new_n964), .B2(new_n965), .ZN(G1352gat));
  OR3_X1    g765(.A1(new_n957), .A2(KEYINPUT126), .A3(new_n721), .ZN(new_n967));
  OAI21_X1  g766(.A(KEYINPUT126), .B1(new_n957), .B2(new_n721), .ZN(new_n968));
  NAND3_X1  g767(.A1(new_n967), .A2(G204gat), .A3(new_n968), .ZN(new_n969));
  NOR3_X1   g768(.A1(new_n959), .A2(G204gat), .A3(new_n721), .ZN(new_n970));
  XNOR2_X1  g769(.A(new_n970), .B(KEYINPUT62), .ZN(new_n971));
  NAND2_X1  g770(.A1(new_n969), .A2(new_n971), .ZN(G1353gat));
  AND2_X1   g771(.A1(new_n960), .A2(new_n962), .ZN(new_n973));
  NAND3_X1  g772(.A1(new_n973), .A2(new_n510), .A3(new_n366), .ZN(new_n974));
  NAND3_X1  g773(.A1(new_n900), .A2(new_n366), .A3(new_n954), .ZN(new_n975));
  AOI21_X1  g774(.A(KEYINPUT63), .B1(new_n975), .B2(G211gat), .ZN(new_n976));
  NAND3_X1  g775(.A1(new_n975), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n977));
  INV_X1    g776(.A(new_n977), .ZN(new_n978));
  OAI21_X1  g777(.A(new_n974), .B1(new_n976), .B2(new_n978), .ZN(G1354gat));
  AOI21_X1  g778(.A(G218gat), .B1(new_n973), .B2(new_n682), .ZN(new_n980));
  INV_X1    g779(.A(KEYINPUT127), .ZN(new_n981));
  NAND2_X1  g780(.A1(new_n957), .A2(new_n981), .ZN(new_n982));
  OAI211_X1 g781(.A(new_n507), .B(new_n386), .C1(new_n957), .C2(new_n981), .ZN(new_n983));
  INV_X1    g782(.A(new_n983), .ZN(new_n984));
  AOI21_X1  g783(.A(new_n980), .B1(new_n982), .B2(new_n984), .ZN(G1355gat));
endmodule


