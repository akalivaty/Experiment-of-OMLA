//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 1 1 0 0 0 1 0 1 0 0 1 0 1 0 0 0 0 1 1 1 1 1 0 0 1 0 0 0 0 1 0 0 0 0 1 1 0 1 0 1 0 1 0 0 1 1 1 0 1 0 1 0 1 1 0 1 1 0 1 0 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:30:58 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n457, new_n458,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n483, new_n484, new_n485, new_n486,
    new_n487, new_n488, new_n489, new_n490, new_n491, new_n492, new_n493,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n532, new_n533, new_n534, new_n535, new_n536, new_n537, new_n538,
    new_n539, new_n540, new_n541, new_n542, new_n543, new_n544, new_n546,
    new_n547, new_n548, new_n549, new_n550, new_n551, new_n552, new_n553,
    new_n554, new_n555, new_n556, new_n557, new_n559, new_n560, new_n561,
    new_n562, new_n563, new_n566, new_n567, new_n568, new_n569, new_n570,
    new_n571, new_n572, new_n573, new_n574, new_n576, new_n578, new_n579,
    new_n581, new_n582, new_n583, new_n584, new_n585, new_n586, new_n587,
    new_n590, new_n591, new_n592, new_n594, new_n595, new_n596, new_n598,
    new_n599, new_n600, new_n601, new_n602, new_n603, new_n604, new_n606,
    new_n607, new_n608, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n629, new_n630,
    new_n633, new_n634, new_n636, new_n637, new_n638, new_n640, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1180, new_n1181, new_n1182;
  XOR2_X1   g000(.A(KEYINPUT64), .B(G452), .Z(G350));
  XNOR2_X1  g001(.A(KEYINPUT65), .B(G452), .ZN(G335));
  XNOR2_X1  g002(.A(KEYINPUT66), .B(G452), .ZN(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  XOR2_X1   g008(.A(KEYINPUT67), .B(G44), .Z(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G218), .A2(G220), .A3(G221), .A4(G219), .ZN(new_n450));
  XOR2_X1   g025(.A(new_n450), .B(KEYINPUT2), .Z(new_n451));
  NOR4_X1   g026(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n452));
  INV_X1    g027(.A(new_n452), .ZN(new_n453));
  NOR2_X1   g028(.A1(new_n451), .A2(new_n453), .ZN(G325));
  INV_X1    g029(.A(G325), .ZN(G261));
  AOI22_X1  g030(.A1(new_n451), .A2(G2106), .B1(G567), .B2(new_n453), .ZN(G319));
  INV_X1    g031(.A(G2104), .ZN(new_n457));
  AND3_X1   g032(.A1(new_n457), .A2(KEYINPUT70), .A3(KEYINPUT3), .ZN(new_n458));
  XNOR2_X1  g033(.A(KEYINPUT3), .B(G2104), .ZN(new_n459));
  INV_X1    g034(.A(KEYINPUT70), .ZN(new_n460));
  AOI21_X1  g035(.A(new_n458), .B1(new_n459), .B2(new_n460), .ZN(new_n461));
  INV_X1    g036(.A(G2105), .ZN(new_n462));
  NAND2_X1  g037(.A1(new_n462), .A2(G137), .ZN(new_n463));
  OAI21_X1  g038(.A(KEYINPUT71), .B1(new_n461), .B2(new_n463), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n457), .A2(KEYINPUT3), .ZN(new_n465));
  INV_X1    g040(.A(KEYINPUT3), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n466), .A2(G2104), .ZN(new_n467));
  NAND3_X1  g042(.A1(new_n465), .A2(new_n467), .A3(new_n460), .ZN(new_n468));
  NAND3_X1  g043(.A1(new_n457), .A2(KEYINPUT70), .A3(KEYINPUT3), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  INV_X1    g045(.A(KEYINPUT71), .ZN(new_n471));
  INV_X1    g046(.A(new_n463), .ZN(new_n472));
  NAND3_X1  g047(.A1(new_n470), .A2(new_n471), .A3(new_n472), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n464), .A2(new_n473), .ZN(new_n474));
  NOR2_X1   g049(.A1(new_n457), .A2(G2105), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n475), .A2(G101), .ZN(new_n476));
  AOI21_X1  g051(.A(KEYINPUT72), .B1(new_n474), .B2(new_n476), .ZN(new_n477));
  INV_X1    g052(.A(KEYINPUT72), .ZN(new_n478));
  INV_X1    g053(.A(new_n476), .ZN(new_n479));
  AOI211_X1 g054(.A(new_n478), .B(new_n479), .C1(new_n464), .C2(new_n473), .ZN(new_n480));
  NOR2_X1   g055(.A1(new_n477), .A2(new_n480), .ZN(new_n481));
  INV_X1    g056(.A(G113), .ZN(new_n482));
  OAI21_X1  g057(.A(KEYINPUT68), .B1(new_n482), .B2(new_n457), .ZN(new_n483));
  INV_X1    g058(.A(KEYINPUT68), .ZN(new_n484));
  NAND3_X1  g059(.A1(new_n484), .A2(G113), .A3(G2104), .ZN(new_n485));
  NAND2_X1  g060(.A1(new_n465), .A2(new_n467), .ZN(new_n486));
  INV_X1    g061(.A(G125), .ZN(new_n487));
  OAI211_X1 g062(.A(new_n483), .B(new_n485), .C1(new_n486), .C2(new_n487), .ZN(new_n488));
  INV_X1    g063(.A(KEYINPUT69), .ZN(new_n489));
  AND3_X1   g064(.A1(new_n488), .A2(new_n489), .A3(G2105), .ZN(new_n490));
  AOI21_X1  g065(.A(new_n489), .B1(new_n488), .B2(G2105), .ZN(new_n491));
  NOR2_X1   g066(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  NAND2_X1  g067(.A1(new_n481), .A2(new_n492), .ZN(new_n493));
  INV_X1    g068(.A(new_n493), .ZN(G160));
  OAI21_X1  g069(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n495));
  INV_X1    g070(.A(G112), .ZN(new_n496));
  AOI21_X1  g071(.A(new_n495), .B1(new_n496), .B2(G2105), .ZN(new_n497));
  NAND2_X1  g072(.A1(new_n470), .A2(G2105), .ZN(new_n498));
  INV_X1    g073(.A(new_n498), .ZN(new_n499));
  AOI21_X1  g074(.A(new_n497), .B1(new_n499), .B2(G124), .ZN(new_n500));
  NAND2_X1  g075(.A1(new_n470), .A2(new_n462), .ZN(new_n501));
  INV_X1    g076(.A(new_n501), .ZN(new_n502));
  NAND2_X1  g077(.A1(new_n502), .A2(G136), .ZN(new_n503));
  NAND2_X1  g078(.A1(new_n500), .A2(new_n503), .ZN(new_n504));
  INV_X1    g079(.A(new_n504), .ZN(G162));
  AND2_X1   g080(.A1(KEYINPUT4), .A2(G138), .ZN(new_n506));
  NAND3_X1  g081(.A1(new_n470), .A2(new_n462), .A3(new_n506), .ZN(new_n507));
  NAND3_X1  g082(.A1(new_n470), .A2(G126), .A3(G2105), .ZN(new_n508));
  OAI21_X1  g083(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n509));
  INV_X1    g084(.A(G114), .ZN(new_n510));
  AOI21_X1  g085(.A(new_n509), .B1(new_n510), .B2(G2105), .ZN(new_n511));
  INV_X1    g086(.A(KEYINPUT4), .ZN(new_n512));
  NAND4_X1  g087(.A1(new_n465), .A2(new_n467), .A3(G138), .A4(new_n462), .ZN(new_n513));
  AOI21_X1  g088(.A(new_n511), .B1(new_n512), .B2(new_n513), .ZN(new_n514));
  NAND3_X1  g089(.A1(new_n507), .A2(new_n508), .A3(new_n514), .ZN(new_n515));
  NAND2_X1  g090(.A1(new_n515), .A2(KEYINPUT73), .ZN(new_n516));
  INV_X1    g091(.A(KEYINPUT73), .ZN(new_n517));
  NAND4_X1  g092(.A1(new_n507), .A2(new_n508), .A3(new_n514), .A4(new_n517), .ZN(new_n518));
  NAND2_X1  g093(.A1(new_n516), .A2(new_n518), .ZN(new_n519));
  INV_X1    g094(.A(new_n519), .ZN(G164));
  AND2_X1   g095(.A1(KEYINPUT6), .A2(G651), .ZN(new_n521));
  NOR2_X1   g096(.A1(KEYINPUT6), .A2(G651), .ZN(new_n522));
  OR2_X1    g097(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  NAND2_X1  g098(.A1(new_n523), .A2(G543), .ZN(new_n524));
  INV_X1    g099(.A(G50), .ZN(new_n525));
  INV_X1    g100(.A(G88), .ZN(new_n526));
  NAND2_X1  g101(.A1(KEYINPUT5), .A2(G543), .ZN(new_n527));
  INV_X1    g102(.A(new_n527), .ZN(new_n528));
  NOR2_X1   g103(.A1(KEYINPUT5), .A2(G543), .ZN(new_n529));
  OAI22_X1  g104(.A1(new_n528), .A2(new_n529), .B1(new_n521), .B2(new_n522), .ZN(new_n530));
  OAI22_X1  g105(.A1(new_n524), .A2(new_n525), .B1(new_n526), .B2(new_n530), .ZN(new_n531));
  OR2_X1    g106(.A1(KEYINPUT5), .A2(G543), .ZN(new_n532));
  NAND2_X1  g107(.A1(new_n532), .A2(new_n527), .ZN(new_n533));
  NAND2_X1  g108(.A1(new_n533), .A2(G62), .ZN(new_n534));
  AOI22_X1  g109(.A1(new_n534), .A2(KEYINPUT74), .B1(G75), .B2(G543), .ZN(new_n535));
  INV_X1    g110(.A(KEYINPUT74), .ZN(new_n536));
  NAND3_X1  g111(.A1(new_n533), .A2(new_n536), .A3(G62), .ZN(new_n537));
  NAND2_X1  g112(.A1(new_n535), .A2(new_n537), .ZN(new_n538));
  NAND2_X1  g113(.A1(new_n538), .A2(G651), .ZN(new_n539));
  INV_X1    g114(.A(KEYINPUT75), .ZN(new_n540));
  NAND2_X1  g115(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  INV_X1    g116(.A(G651), .ZN(new_n542));
  AOI21_X1  g117(.A(new_n542), .B1(new_n535), .B2(new_n537), .ZN(new_n543));
  NAND2_X1  g118(.A1(new_n543), .A2(KEYINPUT75), .ZN(new_n544));
  AOI21_X1  g119(.A(new_n531), .B1(new_n541), .B2(new_n544), .ZN(G166));
  XOR2_X1   g120(.A(KEYINPUT77), .B(KEYINPUT7), .Z(new_n546));
  NAND3_X1  g121(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n547));
  XNOR2_X1  g122(.A(new_n546), .B(new_n547), .ZN(new_n548));
  INV_X1    g123(.A(KEYINPUT76), .ZN(new_n549));
  INV_X1    g124(.A(new_n533), .ZN(new_n550));
  NAND2_X1  g125(.A1(G63), .A2(G651), .ZN(new_n551));
  OAI21_X1  g126(.A(new_n549), .B1(new_n550), .B2(new_n551), .ZN(new_n552));
  NAND4_X1  g127(.A1(new_n533), .A2(KEYINPUT76), .A3(G63), .A4(G651), .ZN(new_n553));
  NAND3_X1  g128(.A1(new_n548), .A2(new_n552), .A3(new_n553), .ZN(new_n554));
  INV_X1    g129(.A(G51), .ZN(new_n555));
  INV_X1    g130(.A(G89), .ZN(new_n556));
  OAI22_X1  g131(.A1(new_n524), .A2(new_n555), .B1(new_n556), .B2(new_n530), .ZN(new_n557));
  NOR2_X1   g132(.A1(new_n554), .A2(new_n557), .ZN(G168));
  INV_X1    g133(.A(G52), .ZN(new_n559));
  INV_X1    g134(.A(G90), .ZN(new_n560));
  OAI22_X1  g135(.A1(new_n524), .A2(new_n559), .B1(new_n560), .B2(new_n530), .ZN(new_n561));
  AOI22_X1  g136(.A1(new_n533), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n562));
  NOR2_X1   g137(.A1(new_n562), .A2(new_n542), .ZN(new_n563));
  OR2_X1    g138(.A1(new_n561), .A2(new_n563), .ZN(G301));
  INV_X1    g139(.A(G301), .ZN(G171));
  AOI22_X1  g140(.A1(new_n533), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n566));
  NOR2_X1   g141(.A1(new_n566), .A2(new_n542), .ZN(new_n567));
  INV_X1    g142(.A(KEYINPUT78), .ZN(new_n568));
  XNOR2_X1  g143(.A(new_n567), .B(new_n568), .ZN(new_n569));
  AND2_X1   g144(.A1(new_n523), .A2(G543), .ZN(new_n570));
  INV_X1    g145(.A(new_n530), .ZN(new_n571));
  AOI22_X1  g146(.A1(new_n570), .A2(G43), .B1(G81), .B2(new_n571), .ZN(new_n572));
  NAND2_X1  g147(.A1(new_n569), .A2(new_n572), .ZN(new_n573));
  INV_X1    g148(.A(new_n573), .ZN(new_n574));
  NAND2_X1  g149(.A1(new_n574), .A2(G860), .ZN(G153));
  AND3_X1   g150(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n576));
  NAND2_X1  g151(.A1(new_n576), .A2(G36), .ZN(G176));
  NAND2_X1  g152(.A1(G1), .A2(G3), .ZN(new_n578));
  XNOR2_X1  g153(.A(new_n578), .B(KEYINPUT8), .ZN(new_n579));
  NAND2_X1  g154(.A1(new_n576), .A2(new_n579), .ZN(G188));
  INV_X1    g155(.A(KEYINPUT79), .ZN(new_n581));
  NAND3_X1  g156(.A1(new_n570), .A2(new_n581), .A3(G53), .ZN(new_n582));
  XNOR2_X1  g157(.A(new_n582), .B(KEYINPUT9), .ZN(new_n583));
  NAND2_X1  g158(.A1(G78), .A2(G543), .ZN(new_n584));
  INV_X1    g159(.A(G65), .ZN(new_n585));
  OAI21_X1  g160(.A(new_n584), .B1(new_n550), .B2(new_n585), .ZN(new_n586));
  AOI22_X1  g161(.A1(new_n586), .A2(G651), .B1(G91), .B2(new_n571), .ZN(new_n587));
  NAND2_X1  g162(.A1(new_n583), .A2(new_n587), .ZN(G299));
  INV_X1    g163(.A(G168), .ZN(G286));
  INV_X1    g164(.A(new_n531), .ZN(new_n590));
  INV_X1    g165(.A(new_n544), .ZN(new_n591));
  NOR2_X1   g166(.A1(new_n543), .A2(KEYINPUT75), .ZN(new_n592));
  OAI21_X1  g167(.A(new_n590), .B1(new_n591), .B2(new_n592), .ZN(G303));
  NAND2_X1  g168(.A1(new_n570), .A2(G49), .ZN(new_n594));
  NAND2_X1  g169(.A1(new_n571), .A2(G87), .ZN(new_n595));
  OAI21_X1  g170(.A(G651), .B1(new_n533), .B2(G74), .ZN(new_n596));
  NAND3_X1  g171(.A1(new_n594), .A2(new_n595), .A3(new_n596), .ZN(G288));
  INV_X1    g172(.A(G61), .ZN(new_n598));
  AOI21_X1  g173(.A(new_n598), .B1(new_n532), .B2(new_n527), .ZN(new_n599));
  NAND2_X1  g174(.A1(G73), .A2(G543), .ZN(new_n600));
  INV_X1    g175(.A(new_n600), .ZN(new_n601));
  OAI21_X1  g176(.A(G651), .B1(new_n599), .B2(new_n601), .ZN(new_n602));
  NAND3_X1  g177(.A1(new_n523), .A2(G86), .A3(new_n533), .ZN(new_n603));
  OAI211_X1 g178(.A(G48), .B(G543), .C1(new_n521), .C2(new_n522), .ZN(new_n604));
  NAND3_X1  g179(.A1(new_n602), .A2(new_n603), .A3(new_n604), .ZN(G305));
  XOR2_X1   g180(.A(KEYINPUT80), .B(G47), .Z(new_n606));
  AOI22_X1  g181(.A1(new_n570), .A2(new_n606), .B1(G85), .B2(new_n571), .ZN(new_n607));
  AOI22_X1  g182(.A1(new_n533), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n608));
  OAI21_X1  g183(.A(new_n607), .B1(new_n542), .B2(new_n608), .ZN(G290));
  NAND2_X1  g184(.A1(new_n571), .A2(G92), .ZN(new_n610));
  XOR2_X1   g185(.A(new_n610), .B(KEYINPUT10), .Z(new_n611));
  NAND2_X1  g186(.A1(new_n570), .A2(KEYINPUT81), .ZN(new_n612));
  INV_X1    g187(.A(G54), .ZN(new_n613));
  INV_X1    g188(.A(KEYINPUT81), .ZN(new_n614));
  AOI21_X1  g189(.A(new_n613), .B1(new_n524), .B2(new_n614), .ZN(new_n615));
  NAND2_X1  g190(.A1(G79), .A2(G543), .ZN(new_n616));
  INV_X1    g191(.A(G66), .ZN(new_n617));
  OAI21_X1  g192(.A(new_n616), .B1(new_n550), .B2(new_n617), .ZN(new_n618));
  AOI22_X1  g193(.A1(new_n612), .A2(new_n615), .B1(G651), .B2(new_n618), .ZN(new_n619));
  NAND2_X1  g194(.A1(new_n611), .A2(new_n619), .ZN(new_n620));
  INV_X1    g195(.A(new_n620), .ZN(new_n621));
  INV_X1    g196(.A(KEYINPUT82), .ZN(new_n622));
  NAND2_X1  g197(.A1(new_n621), .A2(new_n622), .ZN(new_n623));
  AOI21_X1  g198(.A(new_n622), .B1(new_n611), .B2(new_n619), .ZN(new_n624));
  INV_X1    g199(.A(new_n624), .ZN(new_n625));
  AOI21_X1  g200(.A(G868), .B1(new_n623), .B2(new_n625), .ZN(new_n626));
  AOI21_X1  g201(.A(new_n626), .B1(G868), .B2(G171), .ZN(G321));
  XNOR2_X1  g202(.A(G321), .B(KEYINPUT83), .ZN(G284));
  NAND2_X1  g203(.A1(G286), .A2(G868), .ZN(new_n629));
  INV_X1    g204(.A(G299), .ZN(new_n630));
  OAI21_X1  g205(.A(new_n629), .B1(new_n630), .B2(G868), .ZN(G297));
  OAI21_X1  g206(.A(new_n629), .B1(new_n630), .B2(G868), .ZN(G280));
  NAND2_X1  g207(.A1(new_n623), .A2(new_n625), .ZN(new_n633));
  INV_X1    g208(.A(G559), .ZN(new_n634));
  OAI21_X1  g209(.A(new_n633), .B1(new_n634), .B2(G860), .ZN(G148));
  NOR2_X1   g210(.A1(new_n574), .A2(G868), .ZN(new_n636));
  NAND2_X1  g211(.A1(new_n633), .A2(new_n634), .ZN(new_n637));
  AOI21_X1  g212(.A(new_n636), .B1(new_n637), .B2(G868), .ZN(new_n638));
  XOR2_X1   g213(.A(new_n638), .B(KEYINPUT84), .Z(G323));
  XNOR2_X1  g214(.A(KEYINPUT85), .B(KEYINPUT11), .ZN(new_n640));
  XNOR2_X1  g215(.A(G323), .B(new_n640), .ZN(G282));
  OAI21_X1  g216(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n642));
  INV_X1    g217(.A(G111), .ZN(new_n643));
  AOI22_X1  g218(.A1(new_n642), .A2(KEYINPUT86), .B1(new_n643), .B2(G2105), .ZN(new_n644));
  OAI21_X1  g219(.A(new_n644), .B1(KEYINPUT86), .B2(new_n642), .ZN(new_n645));
  INV_X1    g220(.A(G135), .ZN(new_n646));
  INV_X1    g221(.A(G123), .ZN(new_n647));
  OAI221_X1 g222(.A(new_n645), .B1(new_n501), .B2(new_n646), .C1(new_n647), .C2(new_n498), .ZN(new_n648));
  OR2_X1    g223(.A1(new_n648), .A2(G2096), .ZN(new_n649));
  NAND3_X1  g224(.A1(new_n462), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n650));
  XNOR2_X1  g225(.A(new_n650), .B(KEYINPUT12), .ZN(new_n651));
  XNOR2_X1  g226(.A(new_n651), .B(KEYINPUT13), .ZN(new_n652));
  XNOR2_X1  g227(.A(new_n652), .B(G2100), .ZN(new_n653));
  NAND2_X1  g228(.A1(new_n648), .A2(G2096), .ZN(new_n654));
  NAND3_X1  g229(.A1(new_n649), .A2(new_n653), .A3(new_n654), .ZN(new_n655));
  XNOR2_X1  g230(.A(new_n655), .B(KEYINPUT87), .ZN(G156));
  INV_X1    g231(.A(KEYINPUT14), .ZN(new_n657));
  XNOR2_X1  g232(.A(G2427), .B(G2438), .ZN(new_n658));
  XNOR2_X1  g233(.A(new_n658), .B(G2430), .ZN(new_n659));
  XNOR2_X1  g234(.A(KEYINPUT15), .B(G2435), .ZN(new_n660));
  AOI21_X1  g235(.A(new_n657), .B1(new_n659), .B2(new_n660), .ZN(new_n661));
  OAI21_X1  g236(.A(new_n661), .B1(new_n660), .B2(new_n659), .ZN(new_n662));
  XNOR2_X1  g237(.A(G2451), .B(G2454), .ZN(new_n663));
  XNOR2_X1  g238(.A(new_n663), .B(KEYINPUT16), .ZN(new_n664));
  XNOR2_X1  g239(.A(G1341), .B(G1348), .ZN(new_n665));
  XNOR2_X1  g240(.A(new_n664), .B(new_n665), .ZN(new_n666));
  XNOR2_X1  g241(.A(new_n662), .B(new_n666), .ZN(new_n667));
  XNOR2_X1  g242(.A(G2443), .B(G2446), .ZN(new_n668));
  OR2_X1    g243(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  NAND2_X1  g244(.A1(new_n667), .A2(new_n668), .ZN(new_n670));
  AND3_X1   g245(.A1(new_n669), .A2(G14), .A3(new_n670), .ZN(G401));
  XOR2_X1   g246(.A(G2084), .B(G2090), .Z(new_n672));
  XNOR2_X1  g247(.A(G2067), .B(G2678), .ZN(new_n673));
  NAND2_X1  g248(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  AND2_X1   g249(.A1(new_n674), .A2(KEYINPUT17), .ZN(new_n675));
  OR2_X1    g250(.A1(new_n672), .A2(new_n673), .ZN(new_n676));
  AOI21_X1  g251(.A(KEYINPUT18), .B1(new_n675), .B2(new_n676), .ZN(new_n677));
  XOR2_X1   g252(.A(G2072), .B(G2078), .Z(new_n678));
  AOI21_X1  g253(.A(new_n678), .B1(new_n674), .B2(KEYINPUT18), .ZN(new_n679));
  XNOR2_X1  g254(.A(new_n677), .B(new_n679), .ZN(new_n680));
  XNOR2_X1  g255(.A(G2096), .B(G2100), .ZN(new_n681));
  XNOR2_X1  g256(.A(new_n681), .B(KEYINPUT88), .ZN(new_n682));
  XNOR2_X1  g257(.A(new_n680), .B(new_n682), .ZN(G227));
  XOR2_X1   g258(.A(G1971), .B(G1976), .Z(new_n684));
  XNOR2_X1  g259(.A(new_n684), .B(KEYINPUT19), .ZN(new_n685));
  XOR2_X1   g260(.A(G1956), .B(G2474), .Z(new_n686));
  XOR2_X1   g261(.A(G1961), .B(G1966), .Z(new_n687));
  AND2_X1   g262(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  NAND2_X1  g263(.A1(new_n685), .A2(new_n688), .ZN(new_n689));
  XNOR2_X1  g264(.A(new_n689), .B(KEYINPUT20), .ZN(new_n690));
  NOR2_X1   g265(.A1(new_n686), .A2(new_n687), .ZN(new_n691));
  NOR3_X1   g266(.A1(new_n685), .A2(new_n688), .A3(new_n691), .ZN(new_n692));
  AOI21_X1  g267(.A(new_n692), .B1(new_n685), .B2(new_n691), .ZN(new_n693));
  NAND2_X1  g268(.A1(new_n690), .A2(new_n693), .ZN(new_n694));
  XNOR2_X1  g269(.A(G1981), .B(G1986), .ZN(new_n695));
  XNOR2_X1  g270(.A(new_n694), .B(new_n695), .ZN(new_n696));
  XOR2_X1   g271(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n697));
  XNOR2_X1  g272(.A(new_n697), .B(KEYINPUT89), .ZN(new_n698));
  XNOR2_X1  g273(.A(new_n696), .B(new_n698), .ZN(new_n699));
  XNOR2_X1  g274(.A(G1991), .B(G1996), .ZN(new_n700));
  XNOR2_X1  g275(.A(new_n699), .B(new_n700), .ZN(G229));
  NOR2_X1   g276(.A1(G4), .A2(G16), .ZN(new_n702));
  AOI21_X1  g277(.A(new_n702), .B1(new_n633), .B2(G16), .ZN(new_n703));
  INV_X1    g278(.A(G1348), .ZN(new_n704));
  XNOR2_X1  g279(.A(new_n703), .B(new_n704), .ZN(new_n705));
  INV_X1    g280(.A(G2084), .ZN(new_n706));
  INV_X1    g281(.A(G29), .ZN(new_n707));
  OAI21_X1  g282(.A(new_n707), .B1(KEYINPUT24), .B2(G34), .ZN(new_n708));
  AOI21_X1  g283(.A(new_n708), .B1(KEYINPUT24), .B2(G34), .ZN(new_n709));
  AOI21_X1  g284(.A(new_n709), .B1(new_n493), .B2(G29), .ZN(new_n710));
  OAI21_X1  g285(.A(new_n705), .B1(new_n706), .B2(new_n710), .ZN(new_n711));
  AOI21_X1  g286(.A(new_n711), .B1(new_n706), .B2(new_n710), .ZN(new_n712));
  XNOR2_X1  g287(.A(KEYINPUT96), .B(KEYINPUT28), .ZN(new_n713));
  NAND2_X1  g288(.A1(new_n707), .A2(G26), .ZN(new_n714));
  XNOR2_X1  g289(.A(new_n713), .B(new_n714), .ZN(new_n715));
  OR2_X1    g290(.A1(G104), .A2(G2105), .ZN(new_n716));
  OAI211_X1 g291(.A(new_n716), .B(G2104), .C1(G116), .C2(new_n462), .ZN(new_n717));
  INV_X1    g292(.A(G140), .ZN(new_n718));
  INV_X1    g293(.A(G128), .ZN(new_n719));
  OAI221_X1 g294(.A(new_n717), .B1(new_n501), .B2(new_n718), .C1(new_n719), .C2(new_n498), .ZN(new_n720));
  XNOR2_X1  g295(.A(new_n720), .B(KEYINPUT95), .ZN(new_n721));
  AOI21_X1  g296(.A(new_n715), .B1(new_n721), .B2(G29), .ZN(new_n722));
  XNOR2_X1  g297(.A(new_n722), .B(G2067), .ZN(new_n723));
  NOR2_X1   g298(.A1(G5), .A2(G16), .ZN(new_n724));
  XNOR2_X1  g299(.A(new_n724), .B(KEYINPUT99), .ZN(new_n725));
  INV_X1    g300(.A(G16), .ZN(new_n726));
  OAI21_X1  g301(.A(new_n725), .B1(G301), .B2(new_n726), .ZN(new_n727));
  INV_X1    g302(.A(G1961), .ZN(new_n728));
  NOR2_X1   g303(.A1(new_n727), .A2(new_n728), .ZN(new_n729));
  XOR2_X1   g304(.A(new_n729), .B(KEYINPUT100), .Z(new_n730));
  AOI22_X1  g305(.A1(new_n726), .A2(G21), .B1(KEYINPUT98), .B2(G1966), .ZN(new_n731));
  OAI21_X1  g306(.A(new_n731), .B1(G168), .B2(new_n726), .ZN(new_n732));
  NOR2_X1   g307(.A1(KEYINPUT98), .A2(G1966), .ZN(new_n733));
  XNOR2_X1  g308(.A(new_n732), .B(new_n733), .ZN(new_n734));
  NOR2_X1   g309(.A1(G162), .A2(new_n707), .ZN(new_n735));
  AOI21_X1  g310(.A(new_n735), .B1(new_n707), .B2(G35), .ZN(new_n736));
  XOR2_X1   g311(.A(KEYINPUT29), .B(G2090), .Z(new_n737));
  OAI211_X1 g312(.A(new_n730), .B(new_n734), .C1(new_n736), .C2(new_n737), .ZN(new_n738));
  NAND2_X1  g313(.A1(new_n726), .A2(G20), .ZN(new_n739));
  XOR2_X1   g314(.A(new_n739), .B(KEYINPUT23), .Z(new_n740));
  AOI21_X1  g315(.A(new_n740), .B1(G299), .B2(G16), .ZN(new_n741));
  XNOR2_X1  g316(.A(new_n741), .B(G1956), .ZN(new_n742));
  NAND2_X1  g317(.A1(new_n736), .A2(new_n737), .ZN(new_n743));
  NAND2_X1  g318(.A1(new_n742), .A2(new_n743), .ZN(new_n744));
  NAND2_X1  g319(.A1(new_n707), .A2(G33), .ZN(new_n745));
  NAND3_X1  g320(.A1(new_n462), .A2(G103), .A3(G2104), .ZN(new_n746));
  XOR2_X1   g321(.A(new_n746), .B(KEYINPUT25), .Z(new_n747));
  AOI22_X1  g322(.A1(new_n459), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n748));
  OAI21_X1  g323(.A(new_n747), .B1(new_n748), .B2(new_n462), .ZN(new_n749));
  AOI21_X1  g324(.A(new_n749), .B1(G139), .B2(new_n502), .ZN(new_n750));
  OAI21_X1  g325(.A(new_n745), .B1(new_n750), .B2(new_n707), .ZN(new_n751));
  XOR2_X1   g326(.A(new_n751), .B(G2072), .Z(new_n752));
  NAND2_X1  g327(.A1(new_n727), .A2(new_n728), .ZN(new_n753));
  XOR2_X1   g328(.A(KEYINPUT31), .B(G11), .Z(new_n754));
  NOR2_X1   g329(.A1(new_n648), .A2(new_n707), .ZN(new_n755));
  INV_X1    g330(.A(G28), .ZN(new_n756));
  OR2_X1    g331(.A1(new_n756), .A2(KEYINPUT30), .ZN(new_n757));
  AOI21_X1  g332(.A(G29), .B1(new_n756), .B2(KEYINPUT30), .ZN(new_n758));
  AOI211_X1 g333(.A(new_n754), .B(new_n755), .C1(new_n757), .C2(new_n758), .ZN(new_n759));
  NAND3_X1  g334(.A1(new_n752), .A2(new_n753), .A3(new_n759), .ZN(new_n760));
  NOR3_X1   g335(.A1(new_n738), .A2(new_n744), .A3(new_n760), .ZN(new_n761));
  NAND2_X1  g336(.A1(new_n726), .A2(G19), .ZN(new_n762));
  XOR2_X1   g337(.A(new_n762), .B(KEYINPUT93), .Z(new_n763));
  OAI21_X1  g338(.A(new_n763), .B1(new_n574), .B2(new_n726), .ZN(new_n764));
  XNOR2_X1  g339(.A(new_n764), .B(KEYINPUT94), .ZN(new_n765));
  XNOR2_X1  g340(.A(new_n765), .B(G1341), .ZN(new_n766));
  NAND2_X1  g341(.A1(new_n707), .A2(G27), .ZN(new_n767));
  OAI21_X1  g342(.A(new_n767), .B1(G164), .B2(new_n707), .ZN(new_n768));
  XOR2_X1   g343(.A(KEYINPUT101), .B(G2078), .Z(new_n769));
  XNOR2_X1  g344(.A(new_n768), .B(new_n769), .ZN(new_n770));
  AND4_X1   g345(.A1(new_n723), .A2(new_n761), .A3(new_n766), .A4(new_n770), .ZN(new_n771));
  NAND2_X1  g346(.A1(new_n707), .A2(G32), .ZN(new_n772));
  NAND3_X1  g347(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n773));
  INV_X1    g348(.A(KEYINPUT26), .ZN(new_n774));
  OR2_X1    g349(.A1(new_n773), .A2(new_n774), .ZN(new_n775));
  NAND2_X1  g350(.A1(new_n773), .A2(new_n774), .ZN(new_n776));
  AOI22_X1  g351(.A1(new_n775), .A2(new_n776), .B1(G105), .B2(new_n475), .ZN(new_n777));
  INV_X1    g352(.A(G141), .ZN(new_n778));
  INV_X1    g353(.A(G129), .ZN(new_n779));
  OAI221_X1 g354(.A(new_n777), .B1(new_n501), .B2(new_n778), .C1(new_n779), .C2(new_n498), .ZN(new_n780));
  INV_X1    g355(.A(KEYINPUT97), .ZN(new_n781));
  OR2_X1    g356(.A1(new_n780), .A2(new_n781), .ZN(new_n782));
  NAND2_X1  g357(.A1(new_n780), .A2(new_n781), .ZN(new_n783));
  NAND2_X1  g358(.A1(new_n782), .A2(new_n783), .ZN(new_n784));
  INV_X1    g359(.A(new_n784), .ZN(new_n785));
  OAI21_X1  g360(.A(new_n772), .B1(new_n785), .B2(new_n707), .ZN(new_n786));
  XNOR2_X1  g361(.A(new_n786), .B(KEYINPUT27), .ZN(new_n787));
  XNOR2_X1  g362(.A(new_n787), .B(G1996), .ZN(new_n788));
  NAND3_X1  g363(.A1(new_n712), .A2(new_n771), .A3(new_n788), .ZN(new_n789));
  XNOR2_X1  g364(.A(new_n789), .B(KEYINPUT102), .ZN(new_n790));
  NAND2_X1  g365(.A1(new_n726), .A2(G23), .ZN(new_n791));
  INV_X1    g366(.A(G288), .ZN(new_n792));
  OAI21_X1  g367(.A(new_n791), .B1(new_n792), .B2(new_n726), .ZN(new_n793));
  XNOR2_X1  g368(.A(new_n793), .B(KEYINPUT33), .ZN(new_n794));
  XNOR2_X1  g369(.A(new_n794), .B(G1976), .ZN(new_n795));
  NAND2_X1  g370(.A1(G166), .A2(G16), .ZN(new_n796));
  OAI21_X1  g371(.A(new_n796), .B1(G16), .B2(G22), .ZN(new_n797));
  INV_X1    g372(.A(G1971), .ZN(new_n798));
  OR2_X1    g373(.A1(new_n797), .A2(new_n798), .ZN(new_n799));
  NAND2_X1  g374(.A1(new_n797), .A2(new_n798), .ZN(new_n800));
  MUX2_X1   g375(.A(G6), .B(G305), .S(G16), .Z(new_n801));
  XNOR2_X1  g376(.A(KEYINPUT32), .B(G1981), .ZN(new_n802));
  XNOR2_X1  g377(.A(new_n802), .B(KEYINPUT92), .ZN(new_n803));
  XNOR2_X1  g378(.A(new_n801), .B(new_n803), .ZN(new_n804));
  NAND4_X1  g379(.A1(new_n795), .A2(new_n799), .A3(new_n800), .A4(new_n804), .ZN(new_n805));
  OR2_X1    g380(.A1(new_n805), .A2(KEYINPUT34), .ZN(new_n806));
  NAND2_X1  g381(.A1(new_n805), .A2(KEYINPUT34), .ZN(new_n807));
  NAND2_X1  g382(.A1(new_n707), .A2(G25), .ZN(new_n808));
  NAND2_X1  g383(.A1(new_n502), .A2(G131), .ZN(new_n809));
  NAND2_X1  g384(.A1(new_n499), .A2(G119), .ZN(new_n810));
  OR2_X1    g385(.A1(G95), .A2(G2105), .ZN(new_n811));
  OAI211_X1 g386(.A(new_n811), .B(G2104), .C1(G107), .C2(new_n462), .ZN(new_n812));
  NAND3_X1  g387(.A1(new_n809), .A2(new_n810), .A3(new_n812), .ZN(new_n813));
  INV_X1    g388(.A(new_n813), .ZN(new_n814));
  OAI21_X1  g389(.A(new_n808), .B1(new_n814), .B2(new_n707), .ZN(new_n815));
  XNOR2_X1  g390(.A(new_n815), .B(KEYINPUT90), .ZN(new_n816));
  XOR2_X1   g391(.A(KEYINPUT35), .B(G1991), .Z(new_n817));
  XNOR2_X1  g392(.A(new_n816), .B(new_n817), .ZN(new_n818));
  NOR2_X1   g393(.A1(G16), .A2(G24), .ZN(new_n819));
  XNOR2_X1  g394(.A(G290), .B(KEYINPUT91), .ZN(new_n820));
  AOI21_X1  g395(.A(new_n819), .B1(new_n820), .B2(G16), .ZN(new_n821));
  XOR2_X1   g396(.A(new_n821), .B(G1986), .Z(new_n822));
  NAND4_X1  g397(.A1(new_n806), .A2(new_n807), .A3(new_n818), .A4(new_n822), .ZN(new_n823));
  XNOR2_X1  g398(.A(new_n823), .B(KEYINPUT36), .ZN(new_n824));
  NAND2_X1  g399(.A1(new_n790), .A2(new_n824), .ZN(G150));
  INV_X1    g400(.A(G150), .ZN(G311));
  INV_X1    g401(.A(G55), .ZN(new_n827));
  INV_X1    g402(.A(G93), .ZN(new_n828));
  OAI22_X1  g403(.A1(new_n524), .A2(new_n827), .B1(new_n828), .B2(new_n530), .ZN(new_n829));
  AOI22_X1  g404(.A1(new_n533), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n830));
  NOR2_X1   g405(.A1(new_n830), .A2(new_n542), .ZN(new_n831));
  NOR2_X1   g406(.A1(new_n829), .A2(new_n831), .ZN(new_n832));
  OAI21_X1  g407(.A(new_n573), .B1(KEYINPUT103), .B2(new_n832), .ZN(new_n833));
  NAND2_X1  g408(.A1(new_n832), .A2(KEYINPUT103), .ZN(new_n834));
  XOR2_X1   g409(.A(new_n833), .B(new_n834), .Z(new_n835));
  XNOR2_X1  g410(.A(new_n835), .B(KEYINPUT38), .ZN(new_n836));
  NAND2_X1  g411(.A1(new_n633), .A2(G559), .ZN(new_n837));
  XNOR2_X1  g412(.A(new_n836), .B(new_n837), .ZN(new_n838));
  INV_X1    g413(.A(KEYINPUT39), .ZN(new_n839));
  AOI21_X1  g414(.A(G860), .B1(new_n838), .B2(new_n839), .ZN(new_n840));
  OAI21_X1  g415(.A(new_n840), .B1(new_n839), .B2(new_n838), .ZN(new_n841));
  INV_X1    g416(.A(KEYINPUT104), .ZN(new_n842));
  XNOR2_X1  g417(.A(new_n841), .B(new_n842), .ZN(new_n843));
  OAI21_X1  g418(.A(G860), .B1(new_n829), .B2(new_n831), .ZN(new_n844));
  XOR2_X1   g419(.A(new_n844), .B(KEYINPUT37), .Z(new_n845));
  NAND2_X1  g420(.A1(new_n843), .A2(new_n845), .ZN(G145));
  XNOR2_X1  g421(.A(new_n721), .B(new_n750), .ZN(new_n847));
  NAND2_X1  g422(.A1(new_n499), .A2(G130), .ZN(new_n848));
  NOR2_X1   g423(.A1(new_n462), .A2(G118), .ZN(new_n849));
  OAI21_X1  g424(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n850));
  OAI21_X1  g425(.A(new_n848), .B1(new_n849), .B2(new_n850), .ZN(new_n851));
  AOI21_X1  g426(.A(new_n851), .B1(G142), .B2(new_n502), .ZN(new_n852));
  XNOR2_X1  g427(.A(new_n852), .B(new_n651), .ZN(new_n853));
  XOR2_X1   g428(.A(new_n847), .B(new_n853), .Z(new_n854));
  XNOR2_X1  g429(.A(new_n784), .B(new_n515), .ZN(new_n855));
  XNOR2_X1  g430(.A(new_n855), .B(new_n813), .ZN(new_n856));
  NAND2_X1  g431(.A1(new_n854), .A2(new_n856), .ZN(new_n857));
  XNOR2_X1  g432(.A(new_n855), .B(new_n814), .ZN(new_n858));
  XNOR2_X1  g433(.A(new_n847), .B(new_n853), .ZN(new_n859));
  NAND2_X1  g434(.A1(new_n858), .A2(new_n859), .ZN(new_n860));
  NAND2_X1  g435(.A1(new_n857), .A2(new_n860), .ZN(new_n861));
  XNOR2_X1  g436(.A(new_n504), .B(new_n648), .ZN(new_n862));
  XNOR2_X1  g437(.A(new_n862), .B(new_n493), .ZN(new_n863));
  INV_X1    g438(.A(new_n863), .ZN(new_n864));
  OAI21_X1  g439(.A(KEYINPUT105), .B1(new_n861), .B2(new_n864), .ZN(new_n865));
  INV_X1    g440(.A(KEYINPUT105), .ZN(new_n866));
  NAND4_X1  g441(.A1(new_n857), .A2(new_n860), .A3(new_n866), .A4(new_n863), .ZN(new_n867));
  NAND2_X1  g442(.A1(new_n865), .A2(new_n867), .ZN(new_n868));
  AOI21_X1  g443(.A(G37), .B1(new_n861), .B2(new_n864), .ZN(new_n869));
  AND3_X1   g444(.A1(new_n868), .A2(KEYINPUT106), .A3(new_n869), .ZN(new_n870));
  AOI21_X1  g445(.A(KEYINPUT106), .B1(new_n868), .B2(new_n869), .ZN(new_n871));
  XNOR2_X1  g446(.A(KEYINPUT107), .B(KEYINPUT40), .ZN(new_n872));
  INV_X1    g447(.A(new_n872), .ZN(new_n873));
  NOR3_X1   g448(.A1(new_n870), .A2(new_n871), .A3(new_n873), .ZN(new_n874));
  NAND2_X1  g449(.A1(new_n868), .A2(new_n869), .ZN(new_n875));
  INV_X1    g450(.A(KEYINPUT106), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n875), .A2(new_n876), .ZN(new_n877));
  NAND3_X1  g452(.A1(new_n868), .A2(KEYINPUT106), .A3(new_n869), .ZN(new_n878));
  AOI21_X1  g453(.A(new_n872), .B1(new_n877), .B2(new_n878), .ZN(new_n879));
  NOR2_X1   g454(.A1(new_n874), .A2(new_n879), .ZN(G395));
  XNOR2_X1  g455(.A(new_n835), .B(new_n637), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n630), .A2(new_n620), .ZN(new_n882));
  INV_X1    g457(.A(KEYINPUT108), .ZN(new_n883));
  NAND2_X1  g458(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  NAND2_X1  g459(.A1(new_n621), .A2(G299), .ZN(new_n885));
  XNOR2_X1  g460(.A(new_n884), .B(new_n885), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n881), .A2(new_n886), .ZN(new_n887));
  AOI21_X1  g462(.A(KEYINPUT109), .B1(new_n621), .B2(G299), .ZN(new_n888));
  XOR2_X1   g463(.A(new_n888), .B(new_n882), .Z(new_n889));
  INV_X1    g464(.A(KEYINPUT41), .ZN(new_n890));
  AND2_X1   g465(.A1(new_n889), .A2(new_n890), .ZN(new_n891));
  NOR2_X1   g466(.A1(new_n886), .A2(new_n890), .ZN(new_n892));
  NOR2_X1   g467(.A1(new_n891), .A2(new_n892), .ZN(new_n893));
  OAI21_X1  g468(.A(new_n887), .B1(new_n893), .B2(new_n881), .ZN(new_n894));
  XNOR2_X1  g469(.A(G288), .B(KEYINPUT110), .ZN(new_n895));
  XNOR2_X1  g470(.A(G303), .B(new_n895), .ZN(new_n896));
  XNOR2_X1  g471(.A(G290), .B(G305), .ZN(new_n897));
  XNOR2_X1  g472(.A(new_n896), .B(new_n897), .ZN(new_n898));
  XOR2_X1   g473(.A(new_n898), .B(KEYINPUT42), .Z(new_n899));
  XNOR2_X1  g474(.A(new_n894), .B(new_n899), .ZN(new_n900));
  NAND2_X1  g475(.A1(new_n900), .A2(G868), .ZN(new_n901));
  OAI21_X1  g476(.A(new_n901), .B1(G868), .B2(new_n832), .ZN(G295));
  OAI21_X1  g477(.A(new_n901), .B1(G868), .B2(new_n832), .ZN(G331));
  XNOR2_X1  g478(.A(G171), .B(G168), .ZN(new_n904));
  OR2_X1    g479(.A1(new_n835), .A2(new_n904), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n835), .A2(new_n904), .ZN(new_n906));
  NAND3_X1  g481(.A1(new_n905), .A2(new_n886), .A3(new_n906), .ZN(new_n907));
  OR2_X1    g482(.A1(new_n907), .A2(KEYINPUT111), .ZN(new_n908));
  INV_X1    g483(.A(new_n898), .ZN(new_n909));
  OR2_X1    g484(.A1(new_n886), .A2(KEYINPUT41), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n905), .A2(new_n906), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n889), .A2(KEYINPUT41), .ZN(new_n912));
  AND3_X1   g487(.A1(new_n910), .A2(new_n911), .A3(new_n912), .ZN(new_n913));
  NAND2_X1  g488(.A1(new_n907), .A2(KEYINPUT111), .ZN(new_n914));
  OAI211_X1 g489(.A(new_n908), .B(new_n909), .C1(new_n913), .C2(new_n914), .ZN(new_n915));
  INV_X1    g490(.A(KEYINPUT43), .ZN(new_n916));
  INV_X1    g491(.A(G37), .ZN(new_n917));
  OAI21_X1  g492(.A(new_n911), .B1(new_n891), .B2(new_n892), .ZN(new_n918));
  NAND3_X1  g493(.A1(new_n918), .A2(new_n898), .A3(new_n907), .ZN(new_n919));
  NAND4_X1  g494(.A1(new_n915), .A2(new_n916), .A3(new_n917), .A4(new_n919), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n919), .A2(new_n917), .ZN(new_n921));
  AOI21_X1  g496(.A(new_n898), .B1(new_n918), .B2(new_n907), .ZN(new_n922));
  OAI21_X1  g497(.A(KEYINPUT43), .B1(new_n921), .B2(new_n922), .ZN(new_n923));
  NAND2_X1  g498(.A1(new_n920), .A2(new_n923), .ZN(new_n924));
  OAI21_X1  g499(.A(new_n916), .B1(new_n921), .B2(new_n922), .ZN(new_n925));
  NAND3_X1  g500(.A1(new_n915), .A2(new_n917), .A3(new_n919), .ZN(new_n926));
  OAI21_X1  g501(.A(new_n925), .B1(new_n926), .B2(new_n916), .ZN(new_n927));
  MUX2_X1   g502(.A(new_n924), .B(new_n927), .S(KEYINPUT44), .Z(G397));
  INV_X1    g503(.A(G1996), .ZN(new_n929));
  XNOR2_X1  g504(.A(new_n784), .B(new_n929), .ZN(new_n930));
  INV_X1    g505(.A(G2067), .ZN(new_n931));
  XNOR2_X1  g506(.A(new_n721), .B(new_n931), .ZN(new_n932));
  NAND2_X1  g507(.A1(new_n930), .A2(new_n932), .ZN(new_n933));
  XOR2_X1   g508(.A(new_n813), .B(new_n817), .Z(new_n934));
  NOR2_X1   g509(.A1(new_n933), .A2(new_n934), .ZN(new_n935));
  INV_X1    g510(.A(new_n935), .ZN(new_n936));
  NOR2_X1   g511(.A1(G290), .A2(G1986), .ZN(new_n937));
  AND2_X1   g512(.A1(G290), .A2(G1986), .ZN(new_n938));
  OR3_X1    g513(.A1(new_n936), .A2(new_n937), .A3(new_n938), .ZN(new_n939));
  AOI21_X1  g514(.A(new_n471), .B1(new_n470), .B2(new_n472), .ZN(new_n940));
  AOI211_X1 g515(.A(KEYINPUT71), .B(new_n463), .C1(new_n468), .C2(new_n469), .ZN(new_n941));
  OAI21_X1  g516(.A(new_n476), .B1(new_n940), .B2(new_n941), .ZN(new_n942));
  NAND2_X1  g517(.A1(new_n942), .A2(new_n478), .ZN(new_n943));
  OAI211_X1 g518(.A(KEYINPUT72), .B(new_n476), .C1(new_n940), .C2(new_n941), .ZN(new_n944));
  NAND4_X1  g519(.A1(new_n943), .A2(G40), .A3(new_n944), .A4(new_n492), .ZN(new_n945));
  INV_X1    g520(.A(G1384), .ZN(new_n946));
  NAND2_X1  g521(.A1(new_n515), .A2(new_n946), .ZN(new_n947));
  INV_X1    g522(.A(KEYINPUT45), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n947), .A2(new_n948), .ZN(new_n949));
  NOR2_X1   g524(.A1(new_n945), .A2(new_n949), .ZN(new_n950));
  NAND2_X1  g525(.A1(new_n939), .A2(new_n950), .ZN(new_n951));
  INV_X1    g526(.A(new_n951), .ZN(new_n952));
  AND2_X1   g527(.A1(new_n515), .A2(new_n946), .ZN(new_n953));
  NAND4_X1  g528(.A1(new_n481), .A2(G40), .A3(new_n492), .A4(new_n953), .ZN(new_n954));
  INV_X1    g529(.A(G86), .ZN(new_n955));
  OAI21_X1  g530(.A(new_n604), .B1(new_n530), .B2(new_n955), .ZN(new_n956));
  OAI21_X1  g531(.A(G61), .B1(new_n528), .B2(new_n529), .ZN(new_n957));
  AOI21_X1  g532(.A(new_n542), .B1(new_n957), .B2(new_n600), .ZN(new_n958));
  OAI21_X1  g533(.A(G1981), .B1(new_n956), .B2(new_n958), .ZN(new_n959));
  INV_X1    g534(.A(G1981), .ZN(new_n960));
  NAND4_X1  g535(.A1(new_n602), .A2(new_n603), .A3(new_n960), .A4(new_n604), .ZN(new_n961));
  AND3_X1   g536(.A1(new_n959), .A2(KEYINPUT49), .A3(new_n961), .ZN(new_n962));
  AOI21_X1  g537(.A(KEYINPUT49), .B1(new_n959), .B2(new_n961), .ZN(new_n963));
  NOR2_X1   g538(.A1(new_n962), .A2(new_n963), .ZN(new_n964));
  OAI211_X1 g539(.A(G8), .B(new_n964), .C1(new_n945), .C2(new_n947), .ZN(new_n965));
  INV_X1    g540(.A(KEYINPUT115), .ZN(new_n966));
  XNOR2_X1  g541(.A(new_n965), .B(new_n966), .ZN(new_n967));
  INV_X1    g542(.A(G1976), .ZN(new_n968));
  AND3_X1   g543(.A1(new_n967), .A2(new_n968), .A3(new_n792), .ZN(new_n969));
  XOR2_X1   g544(.A(new_n961), .B(KEYINPUT116), .Z(new_n970));
  OAI211_X1 g545(.A(G8), .B(new_n954), .C1(new_n969), .C2(new_n970), .ZN(new_n971));
  INV_X1    g546(.A(G8), .ZN(new_n972));
  AND4_X1   g547(.A1(G40), .A2(new_n943), .A3(new_n944), .A4(new_n492), .ZN(new_n973));
  NAND3_X1  g548(.A1(new_n519), .A2(KEYINPUT45), .A3(new_n946), .ZN(new_n974));
  NAND3_X1  g549(.A1(new_n973), .A2(new_n949), .A3(new_n974), .ZN(new_n975));
  INV_X1    g550(.A(G1966), .ZN(new_n976));
  NAND2_X1  g551(.A1(new_n975), .A2(new_n976), .ZN(new_n977));
  NOR2_X1   g552(.A1(new_n947), .A2(KEYINPUT50), .ZN(new_n978));
  NOR2_X1   g553(.A1(new_n945), .A2(new_n978), .ZN(new_n979));
  NAND2_X1  g554(.A1(new_n519), .A2(new_n946), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n980), .A2(KEYINPUT50), .ZN(new_n981));
  NAND3_X1  g556(.A1(new_n979), .A2(new_n981), .A3(new_n706), .ZN(new_n982));
  AOI21_X1  g557(.A(new_n972), .B1(new_n977), .B2(new_n982), .ZN(new_n983));
  NAND2_X1  g558(.A1(new_n792), .A2(G1976), .ZN(new_n984));
  AOI21_X1  g559(.A(KEYINPUT52), .B1(G288), .B2(new_n968), .ZN(new_n985));
  NAND4_X1  g560(.A1(new_n954), .A2(G8), .A3(new_n984), .A4(new_n985), .ZN(new_n986));
  OAI211_X1 g561(.A(G8), .B(new_n984), .C1(new_n945), .C2(new_n947), .ZN(new_n987));
  NAND2_X1  g562(.A1(new_n987), .A2(KEYINPUT52), .ZN(new_n988));
  AND2_X1   g563(.A1(new_n986), .A2(new_n988), .ZN(new_n989));
  NAND4_X1  g564(.A1(new_n983), .A2(new_n989), .A3(new_n967), .A4(G168), .ZN(new_n990));
  NAND3_X1  g565(.A1(G303), .A2(KEYINPUT55), .A3(G8), .ZN(new_n991));
  INV_X1    g566(.A(KEYINPUT55), .ZN(new_n992));
  OAI21_X1  g567(.A(new_n992), .B1(G166), .B2(new_n972), .ZN(new_n993));
  NAND2_X1  g568(.A1(new_n991), .A2(new_n993), .ZN(new_n994));
  XNOR2_X1  g569(.A(KEYINPUT112), .B(G1971), .ZN(new_n995));
  INV_X1    g570(.A(new_n995), .ZN(new_n996));
  NAND3_X1  g571(.A1(new_n515), .A2(KEYINPUT45), .A3(new_n946), .ZN(new_n997));
  NAND4_X1  g572(.A1(new_n481), .A2(G40), .A3(new_n492), .A4(new_n997), .ZN(new_n998));
  AOI21_X1  g573(.A(KEYINPUT45), .B1(new_n519), .B2(new_n946), .ZN(new_n999));
  OAI21_X1  g574(.A(new_n996), .B1(new_n998), .B2(new_n999), .ZN(new_n1000));
  XNOR2_X1  g575(.A(KEYINPUT113), .B(G2090), .ZN(new_n1001));
  NAND3_X1  g576(.A1(new_n979), .A2(new_n981), .A3(new_n1001), .ZN(new_n1002));
  NAND2_X1  g577(.A1(new_n1000), .A2(new_n1002), .ZN(new_n1003));
  AOI21_X1  g578(.A(new_n994), .B1(new_n1003), .B2(G8), .ZN(new_n1004));
  OAI21_X1  g579(.A(KEYINPUT63), .B1(new_n990), .B2(new_n1004), .ZN(new_n1005));
  NAND2_X1  g580(.A1(new_n947), .A2(KEYINPUT50), .ZN(new_n1006));
  INV_X1    g581(.A(new_n1006), .ZN(new_n1007));
  NOR2_X1   g582(.A1(new_n945), .A2(new_n1007), .ZN(new_n1008));
  INV_X1    g583(.A(KEYINPUT50), .ZN(new_n1009));
  NAND3_X1  g584(.A1(new_n519), .A2(new_n1009), .A3(new_n946), .ZN(new_n1010));
  NAND3_X1  g585(.A1(new_n1008), .A2(new_n1001), .A3(new_n1010), .ZN(new_n1011));
  NAND2_X1  g586(.A1(new_n1000), .A2(new_n1011), .ZN(new_n1012));
  AOI21_X1  g587(.A(new_n994), .B1(new_n1012), .B2(G8), .ZN(new_n1013));
  NOR2_X1   g588(.A1(new_n1013), .A2(KEYINPUT63), .ZN(new_n1014));
  AND2_X1   g589(.A1(new_n983), .A2(G168), .ZN(new_n1015));
  INV_X1    g590(.A(new_n997), .ZN(new_n1016));
  NOR2_X1   g591(.A1(new_n945), .A2(new_n1016), .ZN(new_n1017));
  NAND2_X1  g592(.A1(new_n980), .A2(new_n948), .ZN(new_n1018));
  AOI21_X1  g593(.A(new_n995), .B1(new_n1017), .B2(new_n1018), .ZN(new_n1019));
  AOI21_X1  g594(.A(new_n1009), .B1(new_n519), .B2(new_n946), .ZN(new_n1020));
  INV_X1    g595(.A(new_n1001), .ZN(new_n1021));
  NOR4_X1   g596(.A1(new_n1020), .A2(new_n945), .A3(new_n978), .A4(new_n1021), .ZN(new_n1022));
  OAI211_X1 g597(.A(G8), .B(new_n994), .C1(new_n1019), .C2(new_n1022), .ZN(new_n1023));
  NAND2_X1  g598(.A1(new_n1023), .A2(KEYINPUT114), .ZN(new_n1024));
  INV_X1    g599(.A(KEYINPUT114), .ZN(new_n1025));
  NAND4_X1  g600(.A1(new_n1003), .A2(new_n1025), .A3(G8), .A4(new_n994), .ZN(new_n1026));
  AOI22_X1  g601(.A1(new_n1014), .A2(new_n1015), .B1(new_n1024), .B2(new_n1026), .ZN(new_n1027));
  AND2_X1   g602(.A1(new_n965), .A2(new_n966), .ZN(new_n1028));
  NOR2_X1   g603(.A1(new_n965), .A2(new_n966), .ZN(new_n1029));
  OAI211_X1 g604(.A(new_n988), .B(new_n986), .C1(new_n1028), .C2(new_n1029), .ZN(new_n1030));
  OAI211_X1 g605(.A(new_n971), .B(new_n1005), .C1(new_n1027), .C2(new_n1030), .ZN(new_n1031));
  INV_X1    g606(.A(KEYINPUT120), .ZN(new_n1032));
  NAND2_X1  g607(.A1(new_n1032), .A2(KEYINPUT51), .ZN(new_n1033));
  AOI211_X1 g608(.A(new_n948), .B(G1384), .C1(new_n516), .C2(new_n518), .ZN(new_n1034));
  AOI21_X1  g609(.A(KEYINPUT45), .B1(new_n515), .B2(new_n946), .ZN(new_n1035));
  NOR3_X1   g610(.A1(new_n1034), .A2(new_n945), .A3(new_n1035), .ZN(new_n1036));
  OAI211_X1 g611(.A(new_n982), .B(G168), .C1(G1966), .C2(new_n1036), .ZN(new_n1037));
  INV_X1    g612(.A(KEYINPUT51), .ZN(new_n1038));
  AOI21_X1  g613(.A(new_n972), .B1(KEYINPUT120), .B2(new_n1038), .ZN(new_n1039));
  AOI21_X1  g614(.A(new_n1033), .B1(new_n1037), .B2(new_n1039), .ZN(new_n1040));
  INV_X1    g615(.A(new_n1040), .ZN(new_n1041));
  NAND3_X1  g616(.A1(new_n1037), .A2(new_n1039), .A3(new_n1033), .ZN(new_n1042));
  AOI211_X1 g617(.A(new_n972), .B(G168), .C1(new_n977), .C2(new_n982), .ZN(new_n1043));
  INV_X1    g618(.A(new_n1043), .ZN(new_n1044));
  NAND3_X1  g619(.A1(new_n1041), .A2(new_n1042), .A3(new_n1044), .ZN(new_n1045));
  INV_X1    g620(.A(KEYINPUT54), .ZN(new_n1046));
  INV_X1    g621(.A(KEYINPUT121), .ZN(new_n1047));
  AOI21_X1  g622(.A(G1961), .B1(new_n979), .B2(new_n981), .ZN(new_n1048));
  INV_X1    g623(.A(KEYINPUT53), .ZN(new_n1049));
  NOR3_X1   g624(.A1(new_n1035), .A2(new_n1049), .A3(G2078), .ZN(new_n1050));
  AND3_X1   g625(.A1(new_n973), .A2(new_n974), .A3(new_n1050), .ZN(new_n1051));
  OAI21_X1  g626(.A(new_n1047), .B1(new_n1048), .B2(new_n1051), .ZN(new_n1052));
  NAND3_X1  g627(.A1(new_n973), .A2(new_n974), .A3(new_n1050), .ZN(new_n1053));
  NOR3_X1   g628(.A1(new_n1020), .A2(new_n945), .A3(new_n978), .ZN(new_n1054));
  OAI211_X1 g629(.A(new_n1053), .B(KEYINPUT121), .C1(new_n1054), .C2(G1961), .ZN(new_n1055));
  NAND2_X1  g630(.A1(new_n1052), .A2(new_n1055), .ZN(new_n1056));
  XOR2_X1   g631(.A(KEYINPUT122), .B(KEYINPUT53), .Z(new_n1057));
  NAND2_X1  g632(.A1(new_n1017), .A2(new_n1018), .ZN(new_n1058));
  OAI21_X1  g633(.A(new_n1057), .B1(new_n1058), .B2(G2078), .ZN(new_n1059));
  AOI21_X1  g634(.A(G301), .B1(new_n1056), .B2(new_n1059), .ZN(new_n1060));
  NAND2_X1  g635(.A1(new_n488), .A2(G2105), .ZN(new_n1061));
  INV_X1    g636(.A(G2078), .ZN(new_n1062));
  NAND3_X1  g637(.A1(new_n1061), .A2(G40), .A3(new_n1062), .ZN(new_n1063));
  NOR4_X1   g638(.A1(new_n1016), .A2(new_n1035), .A3(new_n1049), .A4(new_n1063), .ZN(new_n1064));
  INV_X1    g639(.A(KEYINPUT123), .ZN(new_n1065));
  OAI21_X1  g640(.A(new_n1065), .B1(new_n477), .B2(new_n480), .ZN(new_n1066));
  NAND2_X1  g641(.A1(new_n481), .A2(KEYINPUT123), .ZN(new_n1067));
  NAND3_X1  g642(.A1(new_n1064), .A2(new_n1066), .A3(new_n1067), .ZN(new_n1068));
  OAI21_X1  g643(.A(new_n1068), .B1(new_n1054), .B2(G1961), .ZN(new_n1069));
  INV_X1    g644(.A(new_n1057), .ZN(new_n1070));
  NOR3_X1   g645(.A1(new_n999), .A2(new_n945), .A3(new_n1016), .ZN(new_n1071));
  AOI21_X1  g646(.A(new_n1070), .B1(new_n1071), .B2(new_n1062), .ZN(new_n1072));
  NOR3_X1   g647(.A1(new_n1069), .A2(new_n1072), .A3(G171), .ZN(new_n1073));
  OAI21_X1  g648(.A(new_n1046), .B1(new_n1060), .B2(new_n1073), .ZN(new_n1074));
  AOI21_X1  g649(.A(new_n972), .B1(new_n1000), .B2(new_n1011), .ZN(new_n1075));
  OAI211_X1 g650(.A(new_n989), .B(new_n967), .C1(new_n1075), .C2(new_n994), .ZN(new_n1076));
  AOI21_X1  g651(.A(new_n1076), .B1(new_n1024), .B2(new_n1026), .ZN(new_n1077));
  INV_X1    g652(.A(KEYINPUT124), .ZN(new_n1078));
  OAI21_X1  g653(.A(new_n1078), .B1(new_n1069), .B2(new_n1072), .ZN(new_n1079));
  INV_X1    g654(.A(new_n1048), .ZN(new_n1080));
  NAND4_X1  g655(.A1(new_n1059), .A2(new_n1080), .A3(KEYINPUT124), .A4(new_n1068), .ZN(new_n1081));
  NAND3_X1  g656(.A1(new_n1079), .A2(G171), .A3(new_n1081), .ZN(new_n1082));
  NAND3_X1  g657(.A1(new_n1056), .A2(G301), .A3(new_n1059), .ZN(new_n1083));
  NAND3_X1  g658(.A1(new_n1082), .A2(new_n1083), .A3(KEYINPUT54), .ZN(new_n1084));
  AND4_X1   g659(.A1(new_n1045), .A2(new_n1074), .A3(new_n1077), .A4(new_n1084), .ZN(new_n1085));
  INV_X1    g660(.A(G1956), .ZN(new_n1086));
  NAND4_X1  g661(.A1(new_n481), .A2(G40), .A3(new_n492), .A4(new_n1006), .ZN(new_n1087));
  INV_X1    g662(.A(new_n1010), .ZN(new_n1088));
  OAI21_X1  g663(.A(new_n1086), .B1(new_n1087), .B2(new_n1088), .ZN(new_n1089));
  NOR2_X1   g664(.A1(G299), .A2(KEYINPUT57), .ZN(new_n1090));
  INV_X1    g665(.A(KEYINPUT57), .ZN(new_n1091));
  AOI21_X1  g666(.A(new_n1091), .B1(new_n583), .B2(new_n587), .ZN(new_n1092));
  NOR2_X1   g667(.A1(new_n1090), .A2(new_n1092), .ZN(new_n1093));
  XNOR2_X1  g668(.A(KEYINPUT56), .B(G2072), .ZN(new_n1094));
  NAND3_X1  g669(.A1(new_n1017), .A2(new_n1018), .A3(new_n1094), .ZN(new_n1095));
  NAND3_X1  g670(.A1(new_n1089), .A2(new_n1093), .A3(new_n1095), .ZN(new_n1096));
  AOI21_X1  g671(.A(new_n1093), .B1(new_n1089), .B2(new_n1095), .ZN(new_n1097));
  INV_X1    g672(.A(KEYINPUT118), .ZN(new_n1098));
  OAI21_X1  g673(.A(new_n1096), .B1(new_n1097), .B2(new_n1098), .ZN(new_n1099));
  NAND4_X1  g674(.A1(new_n1089), .A2(new_n1093), .A3(new_n1095), .A4(KEYINPUT118), .ZN(new_n1100));
  NAND3_X1  g675(.A1(new_n1099), .A2(KEYINPUT61), .A3(new_n1100), .ZN(new_n1101));
  INV_X1    g676(.A(KEYINPUT119), .ZN(new_n1102));
  NAND2_X1  g677(.A1(new_n1101), .A2(new_n1102), .ZN(new_n1103));
  INV_X1    g678(.A(KEYINPUT59), .ZN(new_n1104));
  NAND3_X1  g679(.A1(new_n1017), .A2(new_n1018), .A3(new_n929), .ZN(new_n1105));
  XOR2_X1   g680(.A(KEYINPUT58), .B(G1341), .Z(new_n1106));
  OAI21_X1  g681(.A(new_n1106), .B1(new_n945), .B2(new_n947), .ZN(new_n1107));
  NAND2_X1  g682(.A1(new_n1105), .A2(new_n1107), .ZN(new_n1108));
  NOR2_X1   g683(.A1(new_n573), .A2(KEYINPUT117), .ZN(new_n1109));
  AOI21_X1  g684(.A(new_n1104), .B1(new_n1108), .B2(new_n1109), .ZN(new_n1110));
  INV_X1    g685(.A(new_n1109), .ZN(new_n1111));
  AOI211_X1 g686(.A(KEYINPUT59), .B(new_n1111), .C1(new_n1105), .C2(new_n1107), .ZN(new_n1112));
  NOR2_X1   g687(.A1(new_n1110), .A2(new_n1112), .ZN(new_n1113));
  OR2_X1    g688(.A1(new_n1090), .A2(new_n1092), .ZN(new_n1114));
  AOI21_X1  g689(.A(G1956), .B1(new_n1008), .B2(new_n1010), .ZN(new_n1115));
  INV_X1    g690(.A(new_n1094), .ZN(new_n1116));
  NOR4_X1   g691(.A1(new_n999), .A2(new_n945), .A3(new_n1016), .A4(new_n1116), .ZN(new_n1117));
  OAI21_X1  g692(.A(new_n1114), .B1(new_n1115), .B2(new_n1117), .ZN(new_n1118));
  AOI21_X1  g693(.A(KEYINPUT61), .B1(new_n1118), .B2(new_n1096), .ZN(new_n1119));
  NAND3_X1  g694(.A1(new_n973), .A2(new_n931), .A3(new_n953), .ZN(new_n1120));
  INV_X1    g695(.A(new_n1120), .ZN(new_n1121));
  AOI21_X1  g696(.A(G1348), .B1(new_n979), .B2(new_n981), .ZN(new_n1122));
  OAI211_X1 g697(.A(KEYINPUT60), .B(new_n633), .C1(new_n1121), .C2(new_n1122), .ZN(new_n1123));
  NAND2_X1  g698(.A1(new_n953), .A2(new_n1009), .ZN(new_n1124));
  NAND4_X1  g699(.A1(new_n481), .A2(new_n1124), .A3(G40), .A4(new_n492), .ZN(new_n1125));
  OAI21_X1  g700(.A(new_n704), .B1(new_n1125), .B2(new_n1020), .ZN(new_n1126));
  INV_X1    g701(.A(KEYINPUT60), .ZN(new_n1127));
  NAND3_X1  g702(.A1(new_n623), .A2(new_n1127), .A3(new_n625), .ZN(new_n1128));
  NOR2_X1   g703(.A1(new_n620), .A2(KEYINPUT82), .ZN(new_n1129));
  OAI21_X1  g704(.A(KEYINPUT60), .B1(new_n1129), .B2(new_n624), .ZN(new_n1130));
  NAND4_X1  g705(.A1(new_n1126), .A2(new_n1128), .A3(new_n1130), .A4(new_n1120), .ZN(new_n1131));
  NAND2_X1  g706(.A1(new_n1123), .A2(new_n1131), .ZN(new_n1132));
  NOR3_X1   g707(.A1(new_n1113), .A2(new_n1119), .A3(new_n1132), .ZN(new_n1133));
  NAND4_X1  g708(.A1(new_n1099), .A2(new_n1100), .A3(KEYINPUT119), .A4(KEYINPUT61), .ZN(new_n1134));
  NAND3_X1  g709(.A1(new_n1103), .A2(new_n1133), .A3(new_n1134), .ZN(new_n1135));
  AOI22_X1  g710(.A1(new_n1126), .A2(new_n1120), .B1(new_n625), .B2(new_n623), .ZN(new_n1136));
  AOI21_X1  g711(.A(new_n1097), .B1(new_n1136), .B2(new_n1096), .ZN(new_n1137));
  NAND2_X1  g712(.A1(new_n1135), .A2(new_n1137), .ZN(new_n1138));
  AOI21_X1  g713(.A(new_n1031), .B1(new_n1085), .B2(new_n1138), .ZN(new_n1139));
  INV_X1    g714(.A(KEYINPUT125), .ZN(new_n1140));
  INV_X1    g715(.A(new_n1042), .ZN(new_n1141));
  NOR4_X1   g716(.A1(new_n1141), .A2(new_n1040), .A3(new_n1043), .A4(KEYINPUT62), .ZN(new_n1142));
  NAND2_X1  g717(.A1(new_n1024), .A2(new_n1026), .ZN(new_n1143));
  NOR2_X1   g718(.A1(new_n1013), .A2(new_n1030), .ZN(new_n1144));
  NAND3_X1  g719(.A1(new_n1060), .A2(new_n1143), .A3(new_n1144), .ZN(new_n1145));
  OAI21_X1  g720(.A(new_n1140), .B1(new_n1142), .B2(new_n1145), .ZN(new_n1146));
  INV_X1    g721(.A(KEYINPUT62), .ZN(new_n1147));
  NAND4_X1  g722(.A1(new_n1041), .A2(new_n1147), .A3(new_n1044), .A4(new_n1042), .ZN(new_n1148));
  NAND4_X1  g723(.A1(new_n1148), .A2(new_n1077), .A3(KEYINPUT125), .A4(new_n1060), .ZN(new_n1149));
  INV_X1    g724(.A(KEYINPUT126), .ZN(new_n1150));
  NOR3_X1   g725(.A1(new_n1141), .A2(new_n1040), .A3(new_n1043), .ZN(new_n1151));
  OAI21_X1  g726(.A(new_n1150), .B1(new_n1151), .B2(new_n1147), .ZN(new_n1152));
  NAND3_X1  g727(.A1(new_n1045), .A2(KEYINPUT126), .A3(KEYINPUT62), .ZN(new_n1153));
  NAND4_X1  g728(.A1(new_n1146), .A2(new_n1149), .A3(new_n1152), .A4(new_n1153), .ZN(new_n1154));
  AOI21_X1  g729(.A(new_n952), .B1(new_n1139), .B2(new_n1154), .ZN(new_n1155));
  NAND2_X1  g730(.A1(new_n932), .A2(new_n785), .ZN(new_n1156));
  NAND2_X1  g731(.A1(new_n1156), .A2(new_n950), .ZN(new_n1157));
  NOR3_X1   g732(.A1(new_n945), .A2(G1996), .A3(new_n949), .ZN(new_n1158));
  NAND2_X1  g733(.A1(new_n1158), .A2(KEYINPUT46), .ZN(new_n1159));
  OR2_X1    g734(.A1(new_n1158), .A2(KEYINPUT46), .ZN(new_n1160));
  NAND3_X1  g735(.A1(new_n1157), .A2(new_n1159), .A3(new_n1160), .ZN(new_n1161));
  XNOR2_X1  g736(.A(new_n1161), .B(KEYINPUT47), .ZN(new_n1162));
  NAND2_X1  g737(.A1(new_n936), .A2(new_n950), .ZN(new_n1163));
  NAND2_X1  g738(.A1(new_n950), .A2(new_n937), .ZN(new_n1164));
  XNOR2_X1  g739(.A(new_n1164), .B(KEYINPUT48), .ZN(new_n1165));
  NAND2_X1  g740(.A1(new_n814), .A2(new_n817), .ZN(new_n1166));
  OAI22_X1  g741(.A1(new_n933), .A2(new_n1166), .B1(G2067), .B2(new_n721), .ZN(new_n1167));
  AOI22_X1  g742(.A1(new_n1163), .A2(new_n1165), .B1(new_n950), .B2(new_n1167), .ZN(new_n1168));
  NAND2_X1  g743(.A1(new_n1162), .A2(new_n1168), .ZN(new_n1169));
  OAI21_X1  g744(.A(KEYINPUT127), .B1(new_n1155), .B2(new_n1169), .ZN(new_n1170));
  NAND2_X1  g745(.A1(new_n1085), .A2(new_n1138), .ZN(new_n1171));
  INV_X1    g746(.A(new_n1031), .ZN(new_n1172));
  NAND3_X1  g747(.A1(new_n1171), .A2(new_n1154), .A3(new_n1172), .ZN(new_n1173));
  NAND2_X1  g748(.A1(new_n1173), .A2(new_n951), .ZN(new_n1174));
  INV_X1    g749(.A(KEYINPUT127), .ZN(new_n1175));
  INV_X1    g750(.A(new_n1169), .ZN(new_n1176));
  NAND3_X1  g751(.A1(new_n1174), .A2(new_n1175), .A3(new_n1176), .ZN(new_n1177));
  NAND2_X1  g752(.A1(new_n1170), .A2(new_n1177), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g753(.A(G319), .ZN(new_n1180));
  OR4_X1    g754(.A1(new_n1180), .A2(G229), .A3(G401), .A4(G227), .ZN(new_n1181));
  AOI21_X1  g755(.A(new_n1181), .B1(new_n920), .B2(new_n923), .ZN(new_n1182));
  OAI21_X1  g756(.A(new_n1182), .B1(new_n871), .B2(new_n870), .ZN(G225));
  INV_X1    g757(.A(G225), .ZN(G308));
endmodule


