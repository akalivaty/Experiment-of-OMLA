//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 0 1 0 0 0 0 0 1 1 1 0 0 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 1 1 0 0 1 0 1 1 1 1 1 1 0 1 0 0 0 1 1 1 1 1 1 0 1 1 0 1 1 0 1 1 0 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:22:13 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n707, new_n708, new_n709, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n720, new_n721, new_n722, new_n724, new_n725, new_n726, new_n728,
    new_n729, new_n730, new_n731, new_n732, new_n733, new_n734, new_n735,
    new_n737, new_n738, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n753, new_n754, new_n755, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n783, new_n784, new_n785, new_n786, new_n787, new_n788, new_n789,
    new_n790, new_n791, new_n792, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n903, new_n904, new_n905,
    new_n906, new_n908, new_n909, new_n910, new_n911, new_n912, new_n913,
    new_n914, new_n915, new_n916, new_n917, new_n918, new_n919, new_n920,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n976, new_n977, new_n978, new_n979, new_n980,
    new_n981, new_n982, new_n983, new_n984, new_n985;
  XOR2_X1   g000(.A(KEYINPUT22), .B(G137), .Z(new_n187));
  INV_X1    g001(.A(G953), .ZN(new_n188));
  AND3_X1   g002(.A1(new_n188), .A2(G221), .A3(G234), .ZN(new_n189));
  XNOR2_X1  g003(.A(new_n187), .B(new_n189), .ZN(new_n190));
  INV_X1    g004(.A(new_n190), .ZN(new_n191));
  INV_X1    g005(.A(G128), .ZN(new_n192));
  OAI211_X1 g006(.A(KEYINPUT74), .B(KEYINPUT23), .C1(new_n192), .C2(G119), .ZN(new_n193));
  OAI21_X1  g007(.A(new_n193), .B1(KEYINPUT74), .B2(KEYINPUT23), .ZN(new_n194));
  INV_X1    g008(.A(G119), .ZN(new_n195));
  NOR2_X1   g009(.A1(new_n195), .A2(G128), .ZN(new_n196));
  MUX2_X1   g010(.A(new_n193), .B(new_n194), .S(new_n196), .Z(new_n197));
  NAND2_X1  g011(.A1(new_n197), .A2(G110), .ZN(new_n198));
  INV_X1    g012(.A(KEYINPUT73), .ZN(new_n199));
  AOI21_X1  g013(.A(new_n199), .B1(new_n195), .B2(G128), .ZN(new_n200));
  MUX2_X1   g014(.A(new_n200), .B(new_n199), .S(new_n196), .Z(new_n201));
  XOR2_X1   g015(.A(KEYINPUT24), .B(G110), .Z(new_n202));
  NAND2_X1  g016(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  INV_X1    g017(.A(G140), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n204), .A2(G125), .ZN(new_n205));
  NOR2_X1   g019(.A1(new_n205), .A2(KEYINPUT16), .ZN(new_n206));
  XNOR2_X1  g020(.A(G125), .B(G140), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n207), .A2(KEYINPUT75), .ZN(new_n208));
  OR2_X1    g022(.A1(new_n205), .A2(KEYINPUT75), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  AOI21_X1  g024(.A(new_n206), .B1(new_n210), .B2(KEYINPUT16), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n211), .A2(G146), .ZN(new_n212));
  INV_X1    g026(.A(new_n212), .ZN(new_n213));
  NOR2_X1   g027(.A1(new_n211), .A2(G146), .ZN(new_n214));
  OAI211_X1 g028(.A(new_n198), .B(new_n203), .C1(new_n213), .C2(new_n214), .ZN(new_n215));
  INV_X1    g029(.A(G146), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n207), .A2(new_n216), .ZN(new_n217));
  NOR2_X1   g031(.A1(new_n197), .A2(G110), .ZN(new_n218));
  NOR2_X1   g032(.A1(new_n201), .A2(new_n202), .ZN(new_n219));
  OAI211_X1 g033(.A(new_n212), .B(new_n217), .C1(new_n218), .C2(new_n219), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n215), .A2(new_n220), .ZN(new_n221));
  AOI21_X1  g035(.A(new_n191), .B1(new_n221), .B2(KEYINPUT76), .ZN(new_n222));
  OAI21_X1  g036(.A(new_n222), .B1(KEYINPUT76), .B2(new_n221), .ZN(new_n223));
  INV_X1    g037(.A(KEYINPUT76), .ZN(new_n224));
  NAND4_X1  g038(.A1(new_n215), .A2(new_n224), .A3(new_n220), .A4(new_n191), .ZN(new_n225));
  AND2_X1   g039(.A1(new_n223), .A2(new_n225), .ZN(new_n226));
  OAI21_X1  g040(.A(KEYINPUT25), .B1(new_n226), .B2(G902), .ZN(new_n227));
  INV_X1    g041(.A(G217), .ZN(new_n228));
  INV_X1    g042(.A(G902), .ZN(new_n229));
  AOI21_X1  g043(.A(new_n228), .B1(G234), .B2(new_n229), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n223), .A2(new_n225), .ZN(new_n231));
  INV_X1    g045(.A(KEYINPUT25), .ZN(new_n232));
  NAND3_X1  g046(.A1(new_n231), .A2(new_n232), .A3(new_n229), .ZN(new_n233));
  NAND3_X1  g047(.A1(new_n227), .A2(new_n230), .A3(new_n233), .ZN(new_n234));
  NOR2_X1   g048(.A1(new_n230), .A2(G902), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n231), .A2(new_n235), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n234), .A2(new_n236), .ZN(new_n237));
  AND2_X1   g051(.A1(KEYINPUT64), .A2(G143), .ZN(new_n238));
  NOR2_X1   g052(.A1(KEYINPUT64), .A2(G143), .ZN(new_n239));
  OAI21_X1  g053(.A(G146), .B1(new_n238), .B2(new_n239), .ZN(new_n240));
  INV_X1    g054(.A(G143), .ZN(new_n241));
  NOR2_X1   g055(.A1(new_n241), .A2(G146), .ZN(new_n242));
  INV_X1    g056(.A(new_n242), .ZN(new_n243));
  AND4_X1   g057(.A1(KEYINPUT0), .A2(new_n240), .A3(G128), .A4(new_n243), .ZN(new_n244));
  XNOR2_X1  g058(.A(KEYINPUT0), .B(G128), .ZN(new_n245));
  OR2_X1    g059(.A1(KEYINPUT64), .A2(G143), .ZN(new_n246));
  NAND2_X1  g060(.A1(KEYINPUT64), .A2(G143), .ZN(new_n247));
  NAND3_X1  g061(.A1(new_n246), .A2(new_n216), .A3(new_n247), .ZN(new_n248));
  NOR2_X1   g062(.A1(new_n216), .A2(G143), .ZN(new_n249));
  INV_X1    g063(.A(new_n249), .ZN(new_n250));
  AOI21_X1  g064(.A(new_n245), .B1(new_n248), .B2(new_n250), .ZN(new_n251));
  NOR2_X1   g065(.A1(new_n244), .A2(new_n251), .ZN(new_n252));
  INV_X1    g066(.A(KEYINPUT11), .ZN(new_n253));
  AND2_X1   g067(.A1(KEYINPUT65), .A2(G134), .ZN(new_n254));
  NOR2_X1   g068(.A1(KEYINPUT65), .A2(G134), .ZN(new_n255));
  OAI21_X1  g069(.A(G137), .B1(new_n254), .B2(new_n255), .ZN(new_n256));
  INV_X1    g070(.A(G134), .ZN(new_n257));
  NOR2_X1   g071(.A1(new_n257), .A2(G137), .ZN(new_n258));
  INV_X1    g072(.A(new_n258), .ZN(new_n259));
  AOI21_X1  g073(.A(new_n253), .B1(new_n256), .B2(new_n259), .ZN(new_n260));
  NOR2_X1   g074(.A1(new_n254), .A2(new_n255), .ZN(new_n261));
  INV_X1    g075(.A(G137), .ZN(new_n262));
  AOI21_X1  g076(.A(KEYINPUT11), .B1(new_n261), .B2(new_n262), .ZN(new_n263));
  OAI21_X1  g077(.A(G131), .B1(new_n260), .B2(new_n263), .ZN(new_n264));
  INV_X1    g078(.A(G131), .ZN(new_n265));
  XNOR2_X1  g079(.A(KEYINPUT65), .B(G134), .ZN(new_n266));
  OAI21_X1  g080(.A(new_n253), .B1(new_n266), .B2(G137), .ZN(new_n267));
  AOI21_X1  g081(.A(new_n258), .B1(new_n266), .B2(G137), .ZN(new_n268));
  OAI211_X1 g082(.A(new_n265), .B(new_n267), .C1(new_n268), .C2(new_n253), .ZN(new_n269));
  AND3_X1   g083(.A1(new_n264), .A2(new_n269), .A3(KEYINPUT68), .ZN(new_n270));
  AOI21_X1  g084(.A(KEYINPUT68), .B1(new_n264), .B2(new_n269), .ZN(new_n271));
  OAI21_X1  g085(.A(new_n252), .B1(new_n270), .B2(new_n271), .ZN(new_n272));
  INV_X1    g086(.A(G116), .ZN(new_n273));
  OAI21_X1  g087(.A(KEYINPUT66), .B1(new_n273), .B2(G119), .ZN(new_n274));
  INV_X1    g088(.A(KEYINPUT66), .ZN(new_n275));
  NAND3_X1  g089(.A1(new_n275), .A2(new_n195), .A3(G116), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n273), .A2(G119), .ZN(new_n277));
  NAND3_X1  g091(.A1(new_n274), .A2(new_n276), .A3(new_n277), .ZN(new_n278));
  XNOR2_X1  g092(.A(KEYINPUT2), .B(G113), .ZN(new_n279));
  OR2_X1    g093(.A1(new_n278), .A2(new_n279), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n278), .A2(new_n279), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n280), .A2(new_n281), .ZN(new_n282));
  INV_X1    g096(.A(KEYINPUT67), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n282), .A2(new_n283), .ZN(new_n284));
  NAND3_X1  g098(.A1(new_n280), .A2(new_n281), .A3(KEYINPUT67), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n284), .A2(new_n285), .ZN(new_n286));
  INV_X1    g100(.A(KEYINPUT1), .ZN(new_n287));
  OAI21_X1  g101(.A(G128), .B1(new_n242), .B2(new_n287), .ZN(new_n288));
  NOR3_X1   g102(.A1(new_n238), .A2(new_n239), .A3(G146), .ZN(new_n289));
  OAI21_X1  g103(.A(new_n288), .B1(new_n289), .B2(new_n249), .ZN(new_n290));
  NAND4_X1  g104(.A1(new_n240), .A2(new_n287), .A3(G128), .A4(new_n243), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n290), .A2(new_n291), .ZN(new_n292));
  NOR2_X1   g106(.A1(new_n266), .A2(G137), .ZN(new_n293));
  NOR2_X1   g107(.A1(new_n262), .A2(G134), .ZN(new_n294));
  OAI21_X1  g108(.A(G131), .B1(new_n293), .B2(new_n294), .ZN(new_n295));
  NAND3_X1  g109(.A1(new_n269), .A2(new_n292), .A3(new_n295), .ZN(new_n296));
  NAND2_X1  g110(.A1(new_n296), .A2(KEYINPUT69), .ZN(new_n297));
  INV_X1    g111(.A(KEYINPUT69), .ZN(new_n298));
  NAND4_X1  g112(.A1(new_n269), .A2(new_n292), .A3(new_n298), .A4(new_n295), .ZN(new_n299));
  NAND4_X1  g113(.A1(new_n272), .A2(new_n286), .A3(new_n297), .A4(new_n299), .ZN(new_n300));
  INV_X1    g114(.A(new_n300), .ZN(new_n301));
  INV_X1    g115(.A(new_n252), .ZN(new_n302));
  INV_X1    g116(.A(KEYINPUT68), .ZN(new_n303));
  NOR3_X1   g117(.A1(new_n260), .A2(new_n263), .A3(G131), .ZN(new_n304));
  INV_X1    g118(.A(KEYINPUT65), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n305), .A2(new_n257), .ZN(new_n306));
  NAND2_X1  g120(.A1(KEYINPUT65), .A2(G134), .ZN(new_n307));
  AOI21_X1  g121(.A(new_n262), .B1(new_n306), .B2(new_n307), .ZN(new_n308));
  OAI21_X1  g122(.A(KEYINPUT11), .B1(new_n308), .B2(new_n258), .ZN(new_n309));
  AOI21_X1  g123(.A(new_n265), .B1(new_n309), .B2(new_n267), .ZN(new_n310));
  OAI21_X1  g124(.A(new_n303), .B1(new_n304), .B2(new_n310), .ZN(new_n311));
  NAND3_X1  g125(.A1(new_n264), .A2(new_n269), .A3(KEYINPUT68), .ZN(new_n312));
  AOI21_X1  g126(.A(new_n302), .B1(new_n311), .B2(new_n312), .ZN(new_n313));
  NAND2_X1  g127(.A1(new_n297), .A2(new_n299), .ZN(new_n314));
  OAI21_X1  g128(.A(KEYINPUT30), .B1(new_n313), .B2(new_n314), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n264), .A2(new_n269), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n316), .A2(new_n252), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n317), .A2(new_n296), .ZN(new_n318));
  OR2_X1    g132(.A1(new_n318), .A2(KEYINPUT30), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n315), .A2(new_n319), .ZN(new_n320));
  INV_X1    g134(.A(new_n286), .ZN(new_n321));
  AOI21_X1  g135(.A(new_n301), .B1(new_n320), .B2(new_n321), .ZN(new_n322));
  INV_X1    g136(.A(G237), .ZN(new_n323));
  NAND3_X1  g137(.A1(new_n323), .A2(new_n188), .A3(G210), .ZN(new_n324));
  INV_X1    g138(.A(G101), .ZN(new_n325));
  XNOR2_X1  g139(.A(new_n324), .B(new_n325), .ZN(new_n326));
  XNOR2_X1  g140(.A(KEYINPUT26), .B(KEYINPUT27), .ZN(new_n327));
  XOR2_X1   g141(.A(new_n326), .B(new_n327), .Z(new_n328));
  OAI21_X1  g142(.A(KEYINPUT70), .B1(new_n322), .B2(new_n328), .ZN(new_n329));
  AND2_X1   g143(.A1(new_n286), .A2(new_n296), .ZN(new_n330));
  AOI21_X1  g144(.A(KEYINPUT28), .B1(new_n330), .B2(new_n272), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n318), .A2(new_n321), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n300), .A2(new_n332), .ZN(new_n333));
  AOI21_X1  g147(.A(new_n331), .B1(new_n333), .B2(KEYINPUT28), .ZN(new_n334));
  AOI21_X1  g148(.A(KEYINPUT29), .B1(new_n334), .B2(new_n328), .ZN(new_n335));
  INV_X1    g149(.A(KEYINPUT70), .ZN(new_n336));
  INV_X1    g150(.A(new_n328), .ZN(new_n337));
  AOI21_X1  g151(.A(new_n286), .B1(new_n315), .B2(new_n319), .ZN(new_n338));
  OAI211_X1 g152(.A(new_n336), .B(new_n337), .C1(new_n338), .C2(new_n301), .ZN(new_n339));
  NAND3_X1  g153(.A1(new_n329), .A2(new_n335), .A3(new_n339), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n340), .A2(KEYINPUT71), .ZN(new_n341));
  INV_X1    g155(.A(KEYINPUT72), .ZN(new_n342));
  OAI21_X1  g156(.A(new_n321), .B1(new_n313), .B2(new_n314), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n343), .A2(new_n300), .ZN(new_n344));
  AOI21_X1  g158(.A(new_n331), .B1(new_n344), .B2(KEYINPUT28), .ZN(new_n345));
  AND2_X1   g159(.A1(new_n328), .A2(KEYINPUT29), .ZN(new_n346));
  AOI211_X1 g160(.A(new_n342), .B(G902), .C1(new_n345), .C2(new_n346), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n344), .A2(KEYINPUT28), .ZN(new_n348));
  INV_X1    g162(.A(new_n331), .ZN(new_n349));
  NAND3_X1  g163(.A1(new_n348), .A2(new_n349), .A3(new_n346), .ZN(new_n350));
  AOI21_X1  g164(.A(KEYINPUT72), .B1(new_n350), .B2(new_n229), .ZN(new_n351));
  NOR2_X1   g165(.A1(new_n347), .A2(new_n351), .ZN(new_n352));
  INV_X1    g166(.A(KEYINPUT71), .ZN(new_n353));
  NAND4_X1  g167(.A1(new_n329), .A2(new_n335), .A3(new_n353), .A4(new_n339), .ZN(new_n354));
  NAND3_X1  g168(.A1(new_n341), .A2(new_n352), .A3(new_n354), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n355), .A2(G472), .ZN(new_n356));
  NOR2_X1   g170(.A1(G472), .A2(G902), .ZN(new_n357));
  INV_X1    g171(.A(KEYINPUT31), .ZN(new_n358));
  NAND3_X1  g172(.A1(new_n322), .A2(new_n358), .A3(new_n328), .ZN(new_n359));
  INV_X1    g173(.A(KEYINPUT28), .ZN(new_n360));
  AOI21_X1  g174(.A(new_n360), .B1(new_n300), .B2(new_n332), .ZN(new_n361));
  OAI21_X1  g175(.A(new_n337), .B1(new_n361), .B2(new_n331), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n359), .A2(new_n362), .ZN(new_n363));
  AOI21_X1  g177(.A(new_n358), .B1(new_n322), .B2(new_n328), .ZN(new_n364));
  OAI21_X1  g178(.A(new_n357), .B1(new_n363), .B2(new_n364), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n365), .A2(KEYINPUT32), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n322), .A2(new_n328), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n367), .A2(KEYINPUT31), .ZN(new_n368));
  NAND3_X1  g182(.A1(new_n368), .A2(new_n359), .A3(new_n362), .ZN(new_n369));
  INV_X1    g183(.A(KEYINPUT32), .ZN(new_n370));
  NAND3_X1  g184(.A1(new_n369), .A2(new_n370), .A3(new_n357), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n366), .A2(new_n371), .ZN(new_n372));
  AOI21_X1  g186(.A(new_n237), .B1(new_n356), .B2(new_n372), .ZN(new_n373));
  INV_X1    g187(.A(new_n373), .ZN(new_n374));
  XNOR2_X1  g188(.A(G110), .B(G140), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n188), .A2(G227), .ZN(new_n376));
  XNOR2_X1  g190(.A(new_n375), .B(new_n376), .ZN(new_n377));
  AND2_X1   g191(.A1(KEYINPUT77), .A2(G107), .ZN(new_n378));
  NOR2_X1   g192(.A1(KEYINPUT77), .A2(G107), .ZN(new_n379));
  NOR3_X1   g193(.A1(new_n378), .A2(new_n379), .A3(G104), .ZN(new_n380));
  INV_X1    g194(.A(G104), .ZN(new_n381));
  NOR2_X1   g195(.A1(new_n381), .A2(G107), .ZN(new_n382));
  OAI21_X1  g196(.A(G101), .B1(new_n380), .B2(new_n382), .ZN(new_n383));
  INV_X1    g197(.A(KEYINPUT3), .ZN(new_n384));
  OAI211_X1 g198(.A(new_n384), .B(G104), .C1(new_n378), .C2(new_n379), .ZN(new_n385));
  OAI21_X1  g199(.A(KEYINPUT3), .B1(new_n381), .B2(G107), .ZN(new_n386));
  NAND2_X1  g200(.A1(new_n381), .A2(G107), .ZN(new_n387));
  NAND4_X1  g201(.A1(new_n385), .A2(new_n325), .A3(new_n386), .A4(new_n387), .ZN(new_n388));
  INV_X1    g202(.A(KEYINPUT78), .ZN(new_n389));
  AND3_X1   g203(.A1(new_n383), .A2(new_n388), .A3(new_n389), .ZN(new_n390));
  AOI21_X1  g204(.A(new_n389), .B1(new_n383), .B2(new_n388), .ZN(new_n391));
  OAI211_X1 g205(.A(KEYINPUT10), .B(new_n292), .C1(new_n390), .C2(new_n391), .ZN(new_n392));
  INV_X1    g206(.A(KEYINPUT10), .ZN(new_n393));
  AOI21_X1  g207(.A(new_n192), .B1(new_n248), .B2(KEYINPUT1), .ZN(new_n394));
  XNOR2_X1  g208(.A(KEYINPUT64), .B(G143), .ZN(new_n395));
  AOI21_X1  g209(.A(new_n242), .B1(new_n395), .B2(G146), .ZN(new_n396));
  OAI21_X1  g210(.A(new_n291), .B1(new_n394), .B2(new_n396), .ZN(new_n397));
  INV_X1    g211(.A(new_n397), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n383), .A2(new_n388), .ZN(new_n399));
  OAI21_X1  g213(.A(new_n393), .B1(new_n398), .B2(new_n399), .ZN(new_n400));
  NAND3_X1  g214(.A1(new_n385), .A2(new_n386), .A3(new_n387), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n401), .A2(G101), .ZN(new_n402));
  NAND3_X1  g216(.A1(new_n402), .A2(KEYINPUT4), .A3(new_n388), .ZN(new_n403));
  INV_X1    g217(.A(KEYINPUT4), .ZN(new_n404));
  NAND3_X1  g218(.A1(new_n401), .A2(new_n404), .A3(G101), .ZN(new_n405));
  NAND3_X1  g219(.A1(new_n403), .A2(new_n252), .A3(new_n405), .ZN(new_n406));
  NAND3_X1  g220(.A1(new_n392), .A2(new_n400), .A3(new_n406), .ZN(new_n407));
  NAND2_X1  g221(.A1(new_n311), .A2(new_n312), .ZN(new_n408));
  OAI21_X1  g222(.A(new_n377), .B1(new_n407), .B2(new_n408), .ZN(new_n409));
  INV_X1    g223(.A(KEYINPUT79), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n409), .A2(new_n410), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n407), .A2(new_n408), .ZN(new_n412));
  NOR2_X1   g226(.A1(new_n270), .A2(new_n271), .ZN(new_n413));
  NAND4_X1  g227(.A1(new_n413), .A2(new_n400), .A3(new_n406), .A4(new_n392), .ZN(new_n414));
  NAND3_X1  g228(.A1(new_n414), .A2(KEYINPUT79), .A3(new_n377), .ZN(new_n415));
  NAND3_X1  g229(.A1(new_n411), .A2(new_n412), .A3(new_n415), .ZN(new_n416));
  INV_X1    g230(.A(KEYINPUT80), .ZN(new_n417));
  INV_X1    g231(.A(new_n377), .ZN(new_n418));
  NAND3_X1  g232(.A1(new_n399), .A2(new_n290), .A3(new_n291), .ZN(new_n419));
  OAI21_X1  g233(.A(new_n419), .B1(new_n398), .B2(new_n399), .ZN(new_n420));
  AOI21_X1  g234(.A(KEYINPUT12), .B1(new_n408), .B2(new_n420), .ZN(new_n421));
  AND3_X1   g235(.A1(new_n420), .A2(KEYINPUT12), .A3(new_n316), .ZN(new_n422));
  NOR2_X1   g236(.A1(new_n421), .A2(new_n422), .ZN(new_n423));
  INV_X1    g237(.A(new_n414), .ZN(new_n424));
  OAI21_X1  g238(.A(new_n418), .B1(new_n423), .B2(new_n424), .ZN(new_n425));
  AND3_X1   g239(.A1(new_n416), .A2(new_n417), .A3(new_n425), .ZN(new_n426));
  AOI21_X1  g240(.A(new_n417), .B1(new_n416), .B2(new_n425), .ZN(new_n427));
  NOR2_X1   g241(.A1(new_n426), .A2(new_n427), .ZN(new_n428));
  OAI211_X1 g242(.A(KEYINPUT81), .B(G469), .C1(new_n428), .C2(G902), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n416), .A2(new_n425), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n430), .A2(KEYINPUT80), .ZN(new_n431));
  NAND3_X1  g245(.A1(new_n416), .A2(new_n417), .A3(new_n425), .ZN(new_n432));
  NAND3_X1  g246(.A1(new_n431), .A2(G469), .A3(new_n432), .ZN(new_n433));
  INV_X1    g247(.A(KEYINPUT81), .ZN(new_n434));
  INV_X1    g248(.A(G469), .ZN(new_n435));
  NOR2_X1   g249(.A1(new_n435), .A2(new_n229), .ZN(new_n436));
  INV_X1    g250(.A(new_n436), .ZN(new_n437));
  NAND3_X1  g251(.A1(new_n433), .A2(new_n434), .A3(new_n437), .ZN(new_n438));
  AND2_X1   g252(.A1(new_n412), .A2(new_n414), .ZN(new_n439));
  OAI22_X1  g253(.A1(new_n439), .A2(new_n377), .B1(new_n423), .B2(new_n409), .ZN(new_n440));
  NAND3_X1  g254(.A1(new_n440), .A2(new_n435), .A3(new_n229), .ZN(new_n441));
  NAND3_X1  g255(.A1(new_n429), .A2(new_n438), .A3(new_n441), .ZN(new_n442));
  INV_X1    g256(.A(KEYINPUT5), .ZN(new_n443));
  NAND3_X1  g257(.A1(new_n443), .A2(new_n195), .A3(G116), .ZN(new_n444));
  OAI211_X1 g258(.A(G113), .B(new_n444), .C1(new_n278), .C2(new_n443), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n445), .A2(new_n280), .ZN(new_n446));
  INV_X1    g260(.A(KEYINPUT84), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n446), .A2(new_n447), .ZN(new_n448));
  INV_X1    g262(.A(new_n399), .ZN(new_n449));
  NAND3_X1  g263(.A1(new_n445), .A2(new_n280), .A3(KEYINPUT84), .ZN(new_n450));
  NAND3_X1  g264(.A1(new_n448), .A2(new_n449), .A3(new_n450), .ZN(new_n451));
  INV_X1    g265(.A(KEYINPUT85), .ZN(new_n452));
  INV_X1    g266(.A(new_n446), .ZN(new_n453));
  OAI211_X1 g267(.A(new_n451), .B(new_n452), .C1(new_n449), .C2(new_n453), .ZN(new_n454));
  XOR2_X1   g268(.A(G110), .B(G122), .Z(new_n455));
  NAND2_X1  g269(.A1(new_n455), .A2(KEYINPUT8), .ZN(new_n456));
  NAND4_X1  g270(.A1(new_n448), .A2(KEYINPUT85), .A3(new_n449), .A4(new_n450), .ZN(new_n457));
  OR2_X1    g271(.A1(new_n455), .A2(KEYINPUT8), .ZN(new_n458));
  NAND4_X1  g272(.A1(new_n454), .A2(new_n456), .A3(new_n457), .A4(new_n458), .ZN(new_n459));
  INV_X1    g273(.A(KEYINPUT87), .ZN(new_n460));
  OAI21_X1  g274(.A(G125), .B1(new_n244), .B2(new_n251), .ZN(new_n461));
  INV_X1    g275(.A(G125), .ZN(new_n462));
  NAND3_X1  g276(.A1(new_n290), .A2(new_n462), .A3(new_n291), .ZN(new_n463));
  AND3_X1   g277(.A1(new_n461), .A2(KEYINPUT86), .A3(new_n463), .ZN(new_n464));
  XNOR2_X1  g278(.A(KEYINPUT83), .B(G224), .ZN(new_n465));
  NAND2_X1  g279(.A1(new_n465), .A2(new_n188), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n466), .A2(KEYINPUT7), .ZN(new_n467));
  OAI21_X1  g281(.A(new_n467), .B1(new_n463), .B2(KEYINPUT86), .ZN(new_n468));
  OAI21_X1  g282(.A(new_n460), .B1(new_n464), .B2(new_n468), .ZN(new_n469));
  NAND4_X1  g283(.A1(new_n284), .A2(new_n403), .A3(new_n285), .A4(new_n405), .ZN(new_n470));
  OAI21_X1  g284(.A(new_n453), .B1(new_n390), .B2(new_n391), .ZN(new_n471));
  INV_X1    g285(.A(new_n455), .ZN(new_n472));
  NAND3_X1  g286(.A1(new_n470), .A2(new_n471), .A3(new_n472), .ZN(new_n473));
  AND2_X1   g287(.A1(new_n469), .A2(new_n473), .ZN(new_n474));
  OR3_X1    g288(.A1(new_n464), .A2(new_n460), .A3(new_n468), .ZN(new_n475));
  AND2_X1   g289(.A1(new_n461), .A2(new_n463), .ZN(new_n476));
  NAND3_X1  g290(.A1(new_n476), .A2(KEYINPUT7), .A3(new_n466), .ZN(new_n477));
  NAND4_X1  g291(.A1(new_n459), .A2(new_n474), .A3(new_n475), .A4(new_n477), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n470), .A2(new_n471), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n479), .A2(new_n455), .ZN(new_n480));
  NAND3_X1  g294(.A1(new_n480), .A2(KEYINPUT6), .A3(new_n473), .ZN(new_n481));
  INV_X1    g295(.A(KEYINPUT6), .ZN(new_n482));
  NAND3_X1  g296(.A1(new_n479), .A2(new_n482), .A3(new_n455), .ZN(new_n483));
  XNOR2_X1  g297(.A(new_n466), .B(KEYINPUT82), .ZN(new_n484));
  XNOR2_X1  g298(.A(new_n476), .B(new_n484), .ZN(new_n485));
  NAND3_X1  g299(.A1(new_n481), .A2(new_n483), .A3(new_n485), .ZN(new_n486));
  NAND3_X1  g300(.A1(new_n478), .A2(new_n486), .A3(new_n229), .ZN(new_n487));
  OAI21_X1  g301(.A(G210), .B1(G237), .B2(G902), .ZN(new_n488));
  INV_X1    g302(.A(new_n488), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n487), .A2(new_n489), .ZN(new_n490));
  INV_X1    g304(.A(KEYINPUT88), .ZN(new_n491));
  NAND4_X1  g305(.A1(new_n478), .A2(new_n486), .A3(new_n229), .A4(new_n488), .ZN(new_n492));
  NAND3_X1  g306(.A1(new_n490), .A2(new_n491), .A3(new_n492), .ZN(new_n493));
  NAND3_X1  g307(.A1(new_n487), .A2(KEYINPUT88), .A3(new_n489), .ZN(new_n494));
  NAND2_X1  g308(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  NAND2_X1  g309(.A1(G234), .A2(G237), .ZN(new_n496));
  NAND3_X1  g310(.A1(new_n496), .A2(G952), .A3(new_n188), .ZN(new_n497));
  INV_X1    g311(.A(new_n497), .ZN(new_n498));
  XOR2_X1   g312(.A(KEYINPUT21), .B(G898), .Z(new_n499));
  INV_X1    g313(.A(new_n499), .ZN(new_n500));
  NAND3_X1  g314(.A1(new_n496), .A2(G902), .A3(G953), .ZN(new_n501));
  INV_X1    g315(.A(new_n501), .ZN(new_n502));
  AOI21_X1  g316(.A(new_n498), .B1(new_n500), .B2(new_n502), .ZN(new_n503));
  OAI21_X1  g317(.A(G214), .B1(G237), .B2(G902), .ZN(new_n504));
  INV_X1    g318(.A(new_n504), .ZN(new_n505));
  NOR3_X1   g319(.A1(new_n495), .A2(new_n503), .A3(new_n505), .ZN(new_n506));
  NOR2_X1   g320(.A1(new_n241), .A2(G128), .ZN(new_n507));
  AOI21_X1  g321(.A(new_n507), .B1(new_n395), .B2(G128), .ZN(new_n508));
  XNOR2_X1  g322(.A(new_n508), .B(new_n266), .ZN(new_n509));
  OR2_X1    g323(.A1(new_n378), .A2(new_n379), .ZN(new_n510));
  XNOR2_X1  g324(.A(G116), .B(G122), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  INV_X1    g326(.A(KEYINPUT96), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  NAND3_X1  g328(.A1(new_n510), .A2(new_n511), .A3(KEYINPUT96), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  INV_X1    g330(.A(KEYINPUT14), .ZN(new_n517));
  NAND2_X1  g331(.A1(new_n511), .A2(new_n517), .ZN(new_n518));
  NAND3_X1  g332(.A1(new_n273), .A2(KEYINPUT14), .A3(G122), .ZN(new_n519));
  NAND3_X1  g333(.A1(new_n518), .A2(G107), .A3(new_n519), .ZN(new_n520));
  NAND3_X1  g334(.A1(new_n509), .A2(new_n516), .A3(new_n520), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n521), .A2(KEYINPUT97), .ZN(new_n522));
  INV_X1    g336(.A(KEYINPUT97), .ZN(new_n523));
  NAND4_X1  g337(.A1(new_n509), .A2(new_n516), .A3(new_n523), .A4(new_n520), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n522), .A2(new_n524), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n508), .A2(new_n266), .ZN(new_n526));
  INV_X1    g340(.A(new_n526), .ZN(new_n527));
  OAI21_X1  g341(.A(G128), .B1(new_n238), .B2(new_n239), .ZN(new_n528));
  XNOR2_X1  g342(.A(KEYINPUT93), .B(KEYINPUT13), .ZN(new_n529));
  INV_X1    g343(.A(new_n507), .ZN(new_n530));
  NAND3_X1  g344(.A1(new_n528), .A2(new_n529), .A3(new_n530), .ZN(new_n531));
  INV_X1    g345(.A(KEYINPUT13), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n532), .A2(KEYINPUT93), .ZN(new_n533));
  INV_X1    g347(.A(KEYINPUT93), .ZN(new_n534));
  NAND2_X1  g348(.A1(new_n534), .A2(KEYINPUT13), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n533), .A2(new_n535), .ZN(new_n536));
  NAND3_X1  g350(.A1(new_n536), .A2(new_n395), .A3(G128), .ZN(new_n537));
  NAND3_X1  g351(.A1(new_n531), .A2(G134), .A3(new_n537), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n538), .A2(KEYINPUT94), .ZN(new_n539));
  INV_X1    g353(.A(KEYINPUT94), .ZN(new_n540));
  NAND4_X1  g354(.A1(new_n531), .A2(new_n537), .A3(new_n540), .A4(G134), .ZN(new_n541));
  AOI21_X1  g355(.A(new_n527), .B1(new_n539), .B2(new_n541), .ZN(new_n542));
  INV_X1    g356(.A(new_n512), .ZN(new_n543));
  NOR2_X1   g357(.A1(new_n510), .A2(new_n511), .ZN(new_n544));
  OAI21_X1  g358(.A(KEYINPUT92), .B1(new_n543), .B2(new_n544), .ZN(new_n545));
  OR2_X1    g359(.A1(new_n510), .A2(new_n511), .ZN(new_n546));
  INV_X1    g360(.A(KEYINPUT92), .ZN(new_n547));
  NAND3_X1  g361(.A1(new_n546), .A2(new_n547), .A3(new_n512), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n545), .A2(new_n548), .ZN(new_n549));
  AND3_X1   g363(.A1(new_n542), .A2(KEYINPUT95), .A3(new_n549), .ZN(new_n550));
  AOI21_X1  g364(.A(KEYINPUT95), .B1(new_n542), .B2(new_n549), .ZN(new_n551));
  OAI21_X1  g365(.A(new_n525), .B1(new_n550), .B2(new_n551), .ZN(new_n552));
  XOR2_X1   g366(.A(KEYINPUT9), .B(G234), .Z(new_n553));
  INV_X1    g367(.A(new_n553), .ZN(new_n554));
  NOR3_X1   g368(.A1(new_n554), .A2(new_n228), .A3(G953), .ZN(new_n555));
  INV_X1    g369(.A(new_n555), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n552), .A2(new_n556), .ZN(new_n557));
  OAI211_X1 g371(.A(new_n525), .B(new_n555), .C1(new_n550), .C2(new_n551), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n557), .A2(new_n558), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n559), .A2(new_n229), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n560), .A2(KEYINPUT98), .ZN(new_n561));
  INV_X1    g375(.A(G478), .ZN(new_n562));
  INV_X1    g376(.A(KEYINPUT99), .ZN(new_n563));
  NOR2_X1   g377(.A1(new_n563), .A2(KEYINPUT15), .ZN(new_n564));
  INV_X1    g378(.A(new_n564), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n563), .A2(KEYINPUT15), .ZN(new_n566));
  AOI21_X1  g380(.A(new_n562), .B1(new_n565), .B2(new_n566), .ZN(new_n567));
  INV_X1    g381(.A(KEYINPUT98), .ZN(new_n568));
  NAND3_X1  g382(.A1(new_n559), .A2(new_n568), .A3(new_n229), .ZN(new_n569));
  NAND3_X1  g383(.A1(new_n561), .A2(new_n567), .A3(new_n569), .ZN(new_n570));
  NOR2_X1   g384(.A1(new_n560), .A2(new_n567), .ZN(new_n571));
  INV_X1    g385(.A(new_n571), .ZN(new_n572));
  NAND2_X1  g386(.A1(new_n570), .A2(new_n572), .ZN(new_n573));
  XNOR2_X1  g387(.A(G113), .B(G122), .ZN(new_n574));
  XNOR2_X1  g388(.A(new_n574), .B(new_n381), .ZN(new_n575));
  INV_X1    g389(.A(new_n575), .ZN(new_n576));
  INV_X1    g390(.A(KEYINPUT19), .ZN(new_n577));
  NAND2_X1  g391(.A1(new_n207), .A2(new_n577), .ZN(new_n578));
  OAI21_X1  g392(.A(new_n578), .B1(new_n210), .B2(new_n577), .ZN(new_n579));
  OAI21_X1  g393(.A(new_n212), .B1(G146), .B2(new_n579), .ZN(new_n580));
  INV_X1    g394(.A(KEYINPUT89), .ZN(new_n581));
  NAND3_X1  g395(.A1(new_n323), .A2(new_n188), .A3(G214), .ZN(new_n582));
  INV_X1    g396(.A(new_n582), .ZN(new_n583));
  NOR2_X1   g397(.A1(new_n238), .A2(new_n239), .ZN(new_n584));
  OAI21_X1  g398(.A(new_n581), .B1(new_n583), .B2(new_n584), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n583), .A2(G143), .ZN(new_n586));
  NAND3_X1  g400(.A1(new_n395), .A2(KEYINPUT89), .A3(new_n582), .ZN(new_n587));
  NAND3_X1  g401(.A1(new_n585), .A2(new_n586), .A3(new_n587), .ZN(new_n588));
  NAND2_X1  g402(.A1(new_n588), .A2(G131), .ZN(new_n589));
  OR2_X1    g403(.A1(new_n588), .A2(G131), .ZN(new_n590));
  AOI21_X1  g404(.A(new_n580), .B1(new_n589), .B2(new_n590), .ZN(new_n591));
  INV_X1    g405(.A(KEYINPUT18), .ZN(new_n592));
  NOR3_X1   g406(.A1(new_n592), .A2(new_n265), .A3(KEYINPUT90), .ZN(new_n593));
  OR2_X1    g407(.A1(new_n588), .A2(new_n593), .ZN(new_n594));
  OAI21_X1  g408(.A(new_n217), .B1(new_n210), .B2(new_n216), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n588), .A2(new_n593), .ZN(new_n596));
  NAND3_X1  g410(.A1(new_n594), .A2(new_n595), .A3(new_n596), .ZN(new_n597));
  INV_X1    g411(.A(new_n597), .ZN(new_n598));
  OAI21_X1  g412(.A(new_n576), .B1(new_n591), .B2(new_n598), .ZN(new_n599));
  NOR2_X1   g413(.A1(new_n213), .A2(new_n214), .ZN(new_n600));
  INV_X1    g414(.A(KEYINPUT17), .ZN(new_n601));
  NAND3_X1  g415(.A1(new_n590), .A2(new_n601), .A3(new_n589), .ZN(new_n602));
  NAND3_X1  g416(.A1(new_n588), .A2(KEYINPUT17), .A3(G131), .ZN(new_n603));
  NAND3_X1  g417(.A1(new_n600), .A2(new_n602), .A3(new_n603), .ZN(new_n604));
  XNOR2_X1  g418(.A(new_n575), .B(KEYINPUT91), .ZN(new_n605));
  NAND3_X1  g419(.A1(new_n604), .A2(new_n597), .A3(new_n605), .ZN(new_n606));
  NAND2_X1  g420(.A1(new_n599), .A2(new_n606), .ZN(new_n607));
  INV_X1    g421(.A(G475), .ZN(new_n608));
  NAND3_X1  g422(.A1(new_n607), .A2(new_n608), .A3(new_n229), .ZN(new_n609));
  INV_X1    g423(.A(KEYINPUT20), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n609), .A2(new_n610), .ZN(new_n611));
  INV_X1    g425(.A(new_n606), .ZN(new_n612));
  AOI21_X1  g426(.A(new_n575), .B1(new_n604), .B2(new_n597), .ZN(new_n613));
  OAI21_X1  g427(.A(new_n229), .B1(new_n612), .B2(new_n613), .ZN(new_n614));
  NAND2_X1  g428(.A1(new_n614), .A2(G475), .ZN(new_n615));
  NAND4_X1  g429(.A1(new_n607), .A2(KEYINPUT20), .A3(new_n608), .A4(new_n229), .ZN(new_n616));
  NAND3_X1  g430(.A1(new_n611), .A2(new_n615), .A3(new_n616), .ZN(new_n617));
  NOR2_X1   g431(.A1(new_n573), .A2(new_n617), .ZN(new_n618));
  INV_X1    g432(.A(G221), .ZN(new_n619));
  AOI21_X1  g433(.A(new_n619), .B1(new_n553), .B2(new_n229), .ZN(new_n620));
  INV_X1    g434(.A(new_n620), .ZN(new_n621));
  NAND4_X1  g435(.A1(new_n442), .A2(new_n506), .A3(new_n618), .A4(new_n621), .ZN(new_n622));
  NOR2_X1   g436(.A1(new_n374), .A2(new_n622), .ZN(new_n623));
  XNOR2_X1  g437(.A(new_n623), .B(new_n325), .ZN(G3));
  INV_X1    g438(.A(new_n237), .ZN(new_n625));
  OAI21_X1  g439(.A(new_n229), .B1(new_n363), .B2(new_n364), .ZN(new_n626));
  AOI22_X1  g440(.A1(new_n626), .A2(G472), .B1(new_n369), .B2(new_n357), .ZN(new_n627));
  NAND4_X1  g441(.A1(new_n625), .A2(new_n442), .A3(new_n621), .A4(new_n627), .ZN(new_n628));
  XNOR2_X1  g442(.A(new_n628), .B(KEYINPUT100), .ZN(new_n629));
  OAI21_X1  g443(.A(KEYINPUT33), .B1(new_n555), .B2(KEYINPUT101), .ZN(new_n630));
  INV_X1    g444(.A(new_n630), .ZN(new_n631));
  AND3_X1   g445(.A1(new_n557), .A2(new_n558), .A3(new_n631), .ZN(new_n632));
  AOI21_X1  g446(.A(new_n631), .B1(new_n557), .B2(new_n558), .ZN(new_n633));
  NOR2_X1   g447(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  NAND4_X1  g448(.A1(new_n634), .A2(KEYINPUT102), .A3(G478), .A4(new_n229), .ZN(new_n635));
  NAND2_X1  g449(.A1(new_n559), .A2(new_n630), .ZN(new_n636));
  NAND3_X1  g450(.A1(new_n557), .A2(new_n558), .A3(new_n631), .ZN(new_n637));
  NAND4_X1  g451(.A1(new_n636), .A2(G478), .A3(new_n229), .A4(new_n637), .ZN(new_n638));
  INV_X1    g452(.A(KEYINPUT102), .ZN(new_n639));
  NAND2_X1  g453(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  NAND3_X1  g454(.A1(new_n561), .A2(new_n562), .A3(new_n569), .ZN(new_n641));
  NAND3_X1  g455(.A1(new_n635), .A2(new_n640), .A3(new_n641), .ZN(new_n642));
  NAND2_X1  g456(.A1(new_n642), .A2(new_n617), .ZN(new_n643));
  NAND2_X1  g457(.A1(new_n490), .A2(new_n492), .ZN(new_n644));
  INV_X1    g458(.A(new_n503), .ZN(new_n645));
  NAND3_X1  g459(.A1(new_n644), .A2(new_n645), .A3(new_n504), .ZN(new_n646));
  NOR3_X1   g460(.A1(new_n629), .A2(new_n643), .A3(new_n646), .ZN(new_n647));
  XNOR2_X1  g461(.A(KEYINPUT34), .B(G104), .ZN(new_n648));
  XNOR2_X1  g462(.A(new_n647), .B(new_n648), .ZN(G6));
  INV_X1    g463(.A(KEYINPUT103), .ZN(new_n650));
  AND3_X1   g464(.A1(new_n611), .A2(new_n615), .A3(new_n616), .ZN(new_n651));
  AOI21_X1  g465(.A(new_n568), .B1(new_n559), .B2(new_n229), .ZN(new_n652));
  AOI211_X1 g466(.A(KEYINPUT98), .B(G902), .C1(new_n557), .C2(new_n558), .ZN(new_n653));
  INV_X1    g467(.A(new_n567), .ZN(new_n654));
  NOR3_X1   g468(.A1(new_n652), .A2(new_n653), .A3(new_n654), .ZN(new_n655));
  OAI21_X1  g469(.A(new_n651), .B1(new_n655), .B2(new_n571), .ZN(new_n656));
  OAI21_X1  g470(.A(new_n650), .B1(new_n656), .B2(new_n646), .ZN(new_n657));
  AOI21_X1  g471(.A(new_n617), .B1(new_n570), .B2(new_n572), .ZN(new_n658));
  AOI211_X1 g472(.A(new_n503), .B(new_n505), .C1(new_n490), .C2(new_n492), .ZN(new_n659));
  NAND3_X1  g473(.A1(new_n658), .A2(new_n659), .A3(KEYINPUT103), .ZN(new_n660));
  AOI21_X1  g474(.A(new_n629), .B1(new_n657), .B2(new_n660), .ZN(new_n661));
  XNOR2_X1  g475(.A(KEYINPUT35), .B(G107), .ZN(new_n662));
  XNOR2_X1  g476(.A(new_n661), .B(new_n662), .ZN(G9));
  INV_X1    g477(.A(new_n627), .ZN(new_n664));
  NOR2_X1   g478(.A1(new_n191), .A2(KEYINPUT36), .ZN(new_n665));
  XNOR2_X1  g479(.A(new_n221), .B(new_n665), .ZN(new_n666));
  NAND2_X1  g480(.A1(new_n666), .A2(new_n235), .ZN(new_n667));
  AND2_X1   g481(.A1(new_n234), .A2(new_n667), .ZN(new_n668));
  OAI21_X1  g482(.A(KEYINPUT104), .B1(new_n664), .B2(new_n668), .ZN(new_n669));
  NAND2_X1  g483(.A1(new_n234), .A2(new_n667), .ZN(new_n670));
  INV_X1    g484(.A(KEYINPUT104), .ZN(new_n671));
  NAND3_X1  g485(.A1(new_n627), .A2(new_n670), .A3(new_n671), .ZN(new_n672));
  NAND2_X1  g486(.A1(new_n669), .A2(new_n672), .ZN(new_n673));
  NOR2_X1   g487(.A1(new_n673), .A2(new_n622), .ZN(new_n674));
  XNOR2_X1  g488(.A(KEYINPUT37), .B(G110), .ZN(new_n675));
  XNOR2_X1  g489(.A(new_n674), .B(new_n675), .ZN(G12));
  AOI21_X1  g490(.A(new_n668), .B1(new_n356), .B2(new_n372), .ZN(new_n677));
  INV_X1    g491(.A(new_n441), .ZN(new_n678));
  AOI21_X1  g492(.A(new_n436), .B1(new_n428), .B2(G469), .ZN(new_n679));
  AOI21_X1  g493(.A(new_n678), .B1(new_n679), .B2(new_n434), .ZN(new_n680));
  AOI21_X1  g494(.A(new_n620), .B1(new_n680), .B2(new_n429), .ZN(new_n681));
  NAND2_X1  g495(.A1(new_n644), .A2(new_n504), .ZN(new_n682));
  INV_X1    g496(.A(new_n682), .ZN(new_n683));
  OR3_X1    g497(.A1(new_n501), .A2(KEYINPUT105), .A3(G900), .ZN(new_n684));
  OAI21_X1  g498(.A(KEYINPUT105), .B1(new_n501), .B2(G900), .ZN(new_n685));
  NAND3_X1  g499(.A1(new_n684), .A2(new_n497), .A3(new_n685), .ZN(new_n686));
  INV_X1    g500(.A(new_n686), .ZN(new_n687));
  NOR2_X1   g501(.A1(new_n656), .A2(new_n687), .ZN(new_n688));
  NAND4_X1  g502(.A1(new_n677), .A2(new_n681), .A3(new_n683), .A4(new_n688), .ZN(new_n689));
  XNOR2_X1  g503(.A(new_n689), .B(G128), .ZN(G30));
  XOR2_X1   g504(.A(new_n686), .B(KEYINPUT39), .Z(new_n691));
  INV_X1    g505(.A(new_n691), .ZN(new_n692));
  NAND2_X1  g506(.A1(new_n681), .A2(new_n692), .ZN(new_n693));
  NAND2_X1  g507(.A1(new_n693), .A2(KEYINPUT40), .ZN(new_n694));
  NAND2_X1  g508(.A1(new_n442), .A2(new_n621), .ZN(new_n695));
  OR3_X1    g509(.A1(new_n695), .A2(KEYINPUT40), .A3(new_n691), .ZN(new_n696));
  XOR2_X1   g510(.A(KEYINPUT106), .B(KEYINPUT38), .Z(new_n697));
  XNOR2_X1  g511(.A(new_n495), .B(new_n697), .ZN(new_n698));
  NOR2_X1   g512(.A1(new_n322), .A2(new_n337), .ZN(new_n699));
  OAI21_X1  g513(.A(new_n229), .B1(new_n344), .B2(new_n328), .ZN(new_n700));
  OAI21_X1  g514(.A(G472), .B1(new_n699), .B2(new_n700), .ZN(new_n701));
  NAND2_X1  g515(.A1(new_n372), .A2(new_n701), .ZN(new_n702));
  AND4_X1   g516(.A1(new_n573), .A2(new_n698), .A3(new_n617), .A4(new_n702), .ZN(new_n703));
  NOR2_X1   g517(.A1(new_n670), .A2(new_n505), .ZN(new_n704));
  NAND4_X1  g518(.A1(new_n694), .A2(new_n696), .A3(new_n703), .A4(new_n704), .ZN(new_n705));
  XNOR2_X1  g519(.A(new_n705), .B(new_n584), .ZN(G45));
  NOR2_X1   g520(.A1(new_n643), .A2(new_n687), .ZN(new_n707));
  NAND4_X1  g521(.A1(new_n677), .A2(new_n681), .A3(new_n683), .A4(new_n707), .ZN(new_n708));
  XOR2_X1   g522(.A(KEYINPUT107), .B(G146), .Z(new_n709));
  XNOR2_X1  g523(.A(new_n708), .B(new_n709), .ZN(G48));
  NOR2_X1   g524(.A1(new_n643), .A2(new_n646), .ZN(new_n711));
  NAND2_X1  g525(.A1(new_n440), .A2(new_n229), .ZN(new_n712));
  NAND2_X1  g526(.A1(new_n712), .A2(G469), .ZN(new_n713));
  AND2_X1   g527(.A1(new_n713), .A2(new_n441), .ZN(new_n714));
  NAND2_X1  g528(.A1(new_n714), .A2(new_n621), .ZN(new_n715));
  INV_X1    g529(.A(new_n715), .ZN(new_n716));
  NAND3_X1  g530(.A1(new_n373), .A2(new_n711), .A3(new_n716), .ZN(new_n717));
  XNOR2_X1  g531(.A(KEYINPUT41), .B(G113), .ZN(new_n718));
  XNOR2_X1  g532(.A(new_n717), .B(new_n718), .ZN(G15));
  NAND2_X1  g533(.A1(new_n657), .A2(new_n660), .ZN(new_n720));
  NAND2_X1  g534(.A1(new_n356), .A2(new_n372), .ZN(new_n721));
  NAND4_X1  g535(.A1(new_n720), .A2(new_n721), .A3(new_n625), .A4(new_n716), .ZN(new_n722));
  XNOR2_X1  g536(.A(new_n722), .B(G116), .ZN(G18));
  NOR3_X1   g537(.A1(new_n715), .A2(new_n573), .A3(new_n617), .ZN(new_n724));
  NAND4_X1  g538(.A1(new_n721), .A2(new_n659), .A3(new_n670), .A4(new_n724), .ZN(new_n725));
  XOR2_X1   g539(.A(KEYINPUT108), .B(G119), .Z(new_n726));
  XNOR2_X1  g540(.A(new_n725), .B(new_n726), .ZN(G21));
  NAND2_X1  g541(.A1(new_n626), .A2(G472), .ZN(new_n728));
  OAI21_X1  g542(.A(new_n359), .B1(new_n328), .B2(new_n345), .ZN(new_n729));
  OAI21_X1  g543(.A(new_n357), .B1(new_n729), .B2(new_n364), .ZN(new_n730));
  NAND2_X1  g544(.A1(new_n728), .A2(new_n730), .ZN(new_n731));
  NOR2_X1   g545(.A1(new_n731), .A2(new_n237), .ZN(new_n732));
  NAND2_X1  g546(.A1(new_n573), .A2(new_n617), .ZN(new_n733));
  NOR2_X1   g547(.A1(new_n733), .A2(new_n715), .ZN(new_n734));
  NAND3_X1  g548(.A1(new_n732), .A2(new_n659), .A3(new_n734), .ZN(new_n735));
  XNOR2_X1  g549(.A(new_n735), .B(G122), .ZN(G24));
  NOR2_X1   g550(.A1(new_n668), .A2(new_n731), .ZN(new_n737));
  NAND4_X1  g551(.A1(new_n737), .A2(new_n707), .A3(new_n683), .A4(new_n716), .ZN(new_n738));
  XNOR2_X1  g552(.A(new_n738), .B(G125), .ZN(G27));
  OAI211_X1 g553(.A(new_n441), .B(new_n437), .C1(new_n435), .C2(new_n430), .ZN(new_n740));
  AND2_X1   g554(.A1(new_n740), .A2(new_n621), .ZN(new_n741));
  AOI21_X1  g555(.A(new_n505), .B1(new_n493), .B2(new_n494), .ZN(new_n742));
  NAND2_X1  g556(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  INV_X1    g557(.A(new_n743), .ZN(new_n744));
  NAND3_X1  g558(.A1(new_n373), .A2(new_n707), .A3(new_n744), .ZN(new_n745));
  INV_X1    g559(.A(KEYINPUT42), .ZN(new_n746));
  NAND2_X1  g560(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  AOI22_X1  g561(.A1(new_n355), .A2(G472), .B1(new_n366), .B2(new_n371), .ZN(new_n748));
  NOR3_X1   g562(.A1(new_n748), .A2(new_n743), .A3(new_n237), .ZN(new_n749));
  NAND3_X1  g563(.A1(new_n749), .A2(KEYINPUT42), .A3(new_n707), .ZN(new_n750));
  NAND2_X1  g564(.A1(new_n747), .A2(new_n750), .ZN(new_n751));
  XNOR2_X1  g565(.A(new_n751), .B(G131), .ZN(G33));
  NAND2_X1  g566(.A1(new_n688), .A2(KEYINPUT109), .ZN(new_n753));
  OR2_X1    g567(.A1(new_n688), .A2(KEYINPUT109), .ZN(new_n754));
  NAND3_X1  g568(.A1(new_n749), .A2(new_n753), .A3(new_n754), .ZN(new_n755));
  XNOR2_X1  g569(.A(new_n755), .B(G134), .ZN(G36));
  OAI21_X1  g570(.A(G469), .B1(new_n428), .B2(KEYINPUT45), .ZN(new_n757));
  NAND2_X1  g571(.A1(new_n757), .A2(KEYINPUT110), .ZN(new_n758));
  NAND3_X1  g572(.A1(new_n416), .A2(KEYINPUT45), .A3(new_n425), .ZN(new_n759));
  INV_X1    g573(.A(KEYINPUT110), .ZN(new_n760));
  OAI211_X1 g574(.A(new_n760), .B(G469), .C1(new_n428), .C2(KEYINPUT45), .ZN(new_n761));
  NAND3_X1  g575(.A1(new_n758), .A2(new_n759), .A3(new_n761), .ZN(new_n762));
  NAND2_X1  g576(.A1(new_n762), .A2(new_n437), .ZN(new_n763));
  INV_X1    g577(.A(KEYINPUT46), .ZN(new_n764));
  NAND2_X1  g578(.A1(new_n763), .A2(new_n764), .ZN(new_n765));
  NAND3_X1  g579(.A1(new_n762), .A2(KEYINPUT46), .A3(new_n437), .ZN(new_n766));
  NAND3_X1  g580(.A1(new_n765), .A2(new_n441), .A3(new_n766), .ZN(new_n767));
  NAND2_X1  g581(.A1(new_n767), .A2(new_n621), .ZN(new_n768));
  NAND2_X1  g582(.A1(new_n642), .A2(new_n651), .ZN(new_n769));
  NAND2_X1  g583(.A1(new_n769), .A2(KEYINPUT43), .ZN(new_n770));
  INV_X1    g584(.A(KEYINPUT43), .ZN(new_n771));
  NAND3_X1  g585(.A1(new_n642), .A2(new_n771), .A3(new_n651), .ZN(new_n772));
  NAND4_X1  g586(.A1(new_n770), .A2(new_n664), .A3(new_n670), .A4(new_n772), .ZN(new_n773));
  INV_X1    g587(.A(KEYINPUT44), .ZN(new_n774));
  AND2_X1   g588(.A1(new_n773), .A2(new_n774), .ZN(new_n775));
  NOR3_X1   g589(.A1(new_n768), .A2(new_n691), .A3(new_n775), .ZN(new_n776));
  OAI21_X1  g590(.A(new_n742), .B1(new_n773), .B2(new_n774), .ZN(new_n777));
  INV_X1    g591(.A(KEYINPUT111), .ZN(new_n778));
  XNOR2_X1  g592(.A(new_n777), .B(new_n778), .ZN(new_n779));
  NAND2_X1  g593(.A1(new_n776), .A2(new_n779), .ZN(new_n780));
  XNOR2_X1  g594(.A(KEYINPUT112), .B(G137), .ZN(new_n781));
  XNOR2_X1  g595(.A(new_n780), .B(new_n781), .ZN(G39));
  INV_X1    g596(.A(KEYINPUT47), .ZN(new_n783));
  NAND2_X1  g597(.A1(new_n783), .A2(KEYINPUT113), .ZN(new_n784));
  NAND2_X1  g598(.A1(new_n768), .A2(new_n784), .ZN(new_n785));
  INV_X1    g599(.A(new_n784), .ZN(new_n786));
  NOR2_X1   g600(.A1(new_n783), .A2(KEYINPUT113), .ZN(new_n787));
  OAI211_X1 g601(.A(new_n767), .B(new_n621), .C1(new_n786), .C2(new_n787), .ZN(new_n788));
  NOR2_X1   g602(.A1(new_n721), .A2(new_n625), .ZN(new_n789));
  INV_X1    g603(.A(new_n742), .ZN(new_n790));
  NOR3_X1   g604(.A1(new_n643), .A2(new_n790), .A3(new_n687), .ZN(new_n791));
  NAND4_X1  g605(.A1(new_n785), .A2(new_n788), .A3(new_n789), .A4(new_n791), .ZN(new_n792));
  XNOR2_X1  g606(.A(new_n792), .B(G140), .ZN(G42));
  XOR2_X1   g607(.A(new_n714), .B(KEYINPUT49), .Z(new_n794));
  NOR3_X1   g608(.A1(new_n794), .A2(new_n698), .A3(new_n237), .ZN(new_n795));
  INV_X1    g609(.A(new_n702), .ZN(new_n796));
  NOR3_X1   g610(.A1(new_n769), .A2(new_n620), .A3(new_n505), .ZN(new_n797));
  NAND3_X1  g611(.A1(new_n795), .A2(new_n796), .A3(new_n797), .ZN(new_n798));
  XNOR2_X1  g612(.A(new_n769), .B(new_n771), .ZN(new_n799));
  AND3_X1   g613(.A1(new_n799), .A2(new_n498), .A3(new_n732), .ZN(new_n800));
  INV_X1    g614(.A(new_n800), .ZN(new_n801));
  NAND2_X1  g615(.A1(new_n785), .A2(new_n788), .ZN(new_n802));
  NAND2_X1  g616(.A1(new_n714), .A2(new_n620), .ZN(new_n803));
  AOI211_X1 g617(.A(new_n790), .B(new_n801), .C1(new_n802), .C2(new_n803), .ZN(new_n804));
  NOR2_X1   g618(.A1(new_n698), .A2(new_n504), .ZN(new_n805));
  NAND3_X1  g619(.A1(new_n800), .A2(new_n716), .A3(new_n805), .ZN(new_n806));
  INV_X1    g620(.A(KEYINPUT50), .ZN(new_n807));
  NAND2_X1  g621(.A1(new_n806), .A2(new_n807), .ZN(new_n808));
  NAND4_X1  g622(.A1(new_n800), .A2(KEYINPUT50), .A3(new_n716), .A4(new_n805), .ZN(new_n809));
  NAND2_X1  g623(.A1(new_n808), .A2(new_n809), .ZN(new_n810));
  AND2_X1   g624(.A1(new_n799), .A2(new_n498), .ZN(new_n811));
  INV_X1    g625(.A(KEYINPUT116), .ZN(new_n812));
  NOR2_X1   g626(.A1(new_n790), .A2(new_n715), .ZN(new_n813));
  AND3_X1   g627(.A1(new_n811), .A2(new_n812), .A3(new_n813), .ZN(new_n814));
  AOI21_X1  g628(.A(new_n812), .B1(new_n811), .B2(new_n813), .ZN(new_n815));
  OAI21_X1  g629(.A(new_n737), .B1(new_n814), .B2(new_n815), .ZN(new_n816));
  NAND4_X1  g630(.A1(new_n796), .A2(new_n813), .A3(new_n625), .A4(new_n498), .ZN(new_n817));
  OR2_X1    g631(.A1(new_n817), .A2(KEYINPUT117), .ZN(new_n818));
  INV_X1    g632(.A(new_n642), .ZN(new_n819));
  NAND2_X1  g633(.A1(new_n817), .A2(KEYINPUT117), .ZN(new_n820));
  NAND4_X1  g634(.A1(new_n818), .A2(new_n651), .A3(new_n819), .A4(new_n820), .ZN(new_n821));
  NAND3_X1  g635(.A1(new_n810), .A2(new_n816), .A3(new_n821), .ZN(new_n822));
  INV_X1    g636(.A(KEYINPUT118), .ZN(new_n823));
  INV_X1    g637(.A(KEYINPUT51), .ZN(new_n824));
  OAI22_X1  g638(.A1(new_n804), .A2(new_n822), .B1(new_n823), .B2(new_n824), .ZN(new_n825));
  NAND2_X1  g639(.A1(new_n802), .A2(new_n803), .ZN(new_n826));
  NAND3_X1  g640(.A1(new_n826), .A2(new_n742), .A3(new_n800), .ZN(new_n827));
  AND3_X1   g641(.A1(new_n810), .A2(new_n821), .A3(new_n816), .ZN(new_n828));
  NOR2_X1   g642(.A1(new_n823), .A2(new_n824), .ZN(new_n829));
  NAND3_X1  g643(.A1(new_n827), .A2(new_n828), .A3(new_n829), .ZN(new_n830));
  NAND2_X1  g644(.A1(new_n823), .A2(new_n824), .ZN(new_n831));
  NAND2_X1  g645(.A1(new_n818), .A2(new_n820), .ZN(new_n832));
  OAI211_X1 g646(.A(G952), .B(new_n188), .C1(new_n832), .C2(new_n643), .ZN(new_n833));
  NOR2_X1   g647(.A1(new_n814), .A2(new_n815), .ZN(new_n834));
  OR3_X1    g648(.A1(new_n834), .A2(KEYINPUT48), .A3(new_n374), .ZN(new_n835));
  OAI21_X1  g649(.A(KEYINPUT48), .B1(new_n834), .B2(new_n374), .ZN(new_n836));
  AOI21_X1  g650(.A(new_n833), .B1(new_n835), .B2(new_n836), .ZN(new_n837));
  NAND4_X1  g651(.A1(new_n825), .A2(new_n830), .A3(new_n831), .A4(new_n837), .ZN(new_n838));
  INV_X1    g652(.A(KEYINPUT53), .ZN(new_n839));
  NAND4_X1  g653(.A1(new_n717), .A2(new_n722), .A3(new_n725), .A4(new_n735), .ZN(new_n840));
  AOI21_X1  g654(.A(new_n622), .B1(new_n673), .B2(new_n374), .ZN(new_n841));
  AND3_X1   g655(.A1(new_n642), .A2(KEYINPUT114), .A3(new_n617), .ZN(new_n842));
  AOI21_X1  g656(.A(KEYINPUT114), .B1(new_n642), .B2(new_n617), .ZN(new_n843));
  NOR3_X1   g657(.A1(new_n842), .A2(new_n843), .A3(new_n658), .ZN(new_n844));
  INV_X1    g658(.A(new_n506), .ZN(new_n845));
  NOR3_X1   g659(.A1(new_n844), .A2(new_n845), .A3(new_n628), .ZN(new_n846));
  NOR3_X1   g660(.A1(new_n840), .A2(new_n841), .A3(new_n846), .ZN(new_n847));
  NOR3_X1   g661(.A1(new_n695), .A2(new_n748), .A3(new_n668), .ZN(new_n848));
  NAND3_X1  g662(.A1(new_n618), .A2(new_n686), .A3(new_n742), .ZN(new_n849));
  OR2_X1    g663(.A1(new_n849), .A2(KEYINPUT115), .ZN(new_n850));
  NAND2_X1  g664(.A1(new_n849), .A2(KEYINPUT115), .ZN(new_n851));
  NAND3_X1  g665(.A1(new_n848), .A2(new_n850), .A3(new_n851), .ZN(new_n852));
  NAND3_X1  g666(.A1(new_n737), .A2(new_n707), .A3(new_n744), .ZN(new_n853));
  AND3_X1   g667(.A1(new_n754), .A2(new_n373), .A3(new_n744), .ZN(new_n854));
  AOI22_X1  g668(.A1(new_n747), .A2(new_n750), .B1(new_n854), .B2(new_n753), .ZN(new_n855));
  NAND4_X1  g669(.A1(new_n847), .A2(new_n852), .A3(new_n853), .A4(new_n855), .ZN(new_n856));
  OAI211_X1 g670(.A(new_n848), .B(new_n683), .C1(new_n688), .C2(new_n707), .ZN(new_n857));
  INV_X1    g671(.A(KEYINPUT52), .ZN(new_n858));
  NOR2_X1   g672(.A1(new_n670), .A2(new_n687), .ZN(new_n859));
  NOR2_X1   g673(.A1(new_n733), .A2(new_n682), .ZN(new_n860));
  NAND4_X1  g674(.A1(new_n702), .A2(new_n859), .A3(new_n741), .A4(new_n860), .ZN(new_n861));
  NAND4_X1  g675(.A1(new_n857), .A2(new_n858), .A3(new_n738), .A4(new_n861), .ZN(new_n862));
  NAND4_X1  g676(.A1(new_n689), .A2(new_n708), .A3(new_n738), .A4(new_n861), .ZN(new_n863));
  NAND2_X1  g677(.A1(new_n863), .A2(KEYINPUT52), .ZN(new_n864));
  NAND2_X1  g678(.A1(new_n862), .A2(new_n864), .ZN(new_n865));
  OAI21_X1  g679(.A(new_n839), .B1(new_n856), .B2(new_n865), .ZN(new_n866));
  AND4_X1   g680(.A1(new_n717), .A2(new_n722), .A3(new_n725), .A4(new_n735), .ZN(new_n867));
  INV_X1    g681(.A(new_n622), .ZN(new_n868));
  AND2_X1   g682(.A1(new_n669), .A2(new_n672), .ZN(new_n869));
  OAI21_X1  g683(.A(new_n868), .B1(new_n869), .B2(new_n373), .ZN(new_n870));
  OR3_X1    g684(.A1(new_n844), .A2(new_n845), .A3(new_n628), .ZN(new_n871));
  NAND4_X1  g685(.A1(new_n867), .A2(new_n870), .A3(new_n871), .A4(new_n852), .ZN(new_n872));
  AOI21_X1  g686(.A(KEYINPUT42), .B1(new_n749), .B2(new_n707), .ZN(new_n873));
  AND4_X1   g687(.A1(KEYINPUT42), .A2(new_n373), .A3(new_n707), .A4(new_n744), .ZN(new_n874));
  OAI211_X1 g688(.A(new_n755), .B(new_n853), .C1(new_n873), .C2(new_n874), .ZN(new_n875));
  NOR2_X1   g689(.A1(new_n872), .A2(new_n875), .ZN(new_n876));
  AND2_X1   g690(.A1(new_n862), .A2(new_n864), .ZN(new_n877));
  NAND3_X1  g691(.A1(new_n876), .A2(new_n877), .A3(KEYINPUT53), .ZN(new_n878));
  AND3_X1   g692(.A1(new_n866), .A2(new_n878), .A3(KEYINPUT54), .ZN(new_n879));
  AOI21_X1  g693(.A(KEYINPUT54), .B1(new_n866), .B2(new_n878), .ZN(new_n880));
  NOR2_X1   g694(.A1(new_n879), .A2(new_n880), .ZN(new_n881));
  NOR3_X1   g695(.A1(new_n801), .A2(new_n682), .A3(new_n715), .ZN(new_n882));
  NOR3_X1   g696(.A1(new_n838), .A2(new_n881), .A3(new_n882), .ZN(new_n883));
  NOR2_X1   g697(.A1(G952), .A2(G953), .ZN(new_n884));
  XOR2_X1   g698(.A(new_n884), .B(KEYINPUT119), .Z(new_n885));
  OAI21_X1  g699(.A(new_n798), .B1(new_n883), .B2(new_n885), .ZN(G75));
  AOI21_X1  g700(.A(new_n229), .B1(new_n866), .B2(new_n878), .ZN(new_n887));
  AOI21_X1  g701(.A(KEYINPUT56), .B1(new_n887), .B2(G210), .ZN(new_n888));
  NAND2_X1  g702(.A1(new_n481), .A2(new_n483), .ZN(new_n889));
  XNOR2_X1  g703(.A(new_n889), .B(new_n485), .ZN(new_n890));
  XOR2_X1   g704(.A(new_n890), .B(KEYINPUT55), .Z(new_n891));
  INV_X1    g705(.A(new_n891), .ZN(new_n892));
  AND2_X1   g706(.A1(new_n888), .A2(new_n892), .ZN(new_n893));
  NOR2_X1   g707(.A1(new_n888), .A2(new_n892), .ZN(new_n894));
  NOR2_X1   g708(.A1(new_n188), .A2(G952), .ZN(new_n895));
  NOR3_X1   g709(.A1(new_n893), .A2(new_n894), .A3(new_n895), .ZN(G51));
  XNOR2_X1  g710(.A(new_n436), .B(KEYINPUT57), .ZN(new_n897));
  NAND2_X1  g711(.A1(new_n881), .A2(new_n897), .ZN(new_n898));
  NAND2_X1  g712(.A1(new_n898), .A2(new_n440), .ZN(new_n899));
  XOR2_X1   g713(.A(new_n762), .B(KEYINPUT120), .Z(new_n900));
  NAND2_X1  g714(.A1(new_n887), .A2(new_n900), .ZN(new_n901));
  AOI21_X1  g715(.A(new_n895), .B1(new_n899), .B2(new_n901), .ZN(G54));
  NAND3_X1  g716(.A1(new_n887), .A2(KEYINPUT58), .A3(G475), .ZN(new_n903));
  INV_X1    g717(.A(new_n607), .ZN(new_n904));
  AND2_X1   g718(.A1(new_n903), .A2(new_n904), .ZN(new_n905));
  NOR2_X1   g719(.A1(new_n903), .A2(new_n904), .ZN(new_n906));
  NOR3_X1   g720(.A1(new_n905), .A2(new_n906), .A3(new_n895), .ZN(G60));
  NAND2_X1  g721(.A1(new_n866), .A2(new_n878), .ZN(new_n908));
  INV_X1    g722(.A(KEYINPUT54), .ZN(new_n909));
  NAND2_X1  g723(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  NAND3_X1  g724(.A1(new_n866), .A2(new_n878), .A3(KEYINPUT54), .ZN(new_n911));
  NAND2_X1  g725(.A1(G478), .A2(G902), .ZN(new_n912));
  XNOR2_X1  g726(.A(new_n912), .B(KEYINPUT59), .ZN(new_n913));
  NAND3_X1  g727(.A1(new_n910), .A2(new_n911), .A3(new_n913), .ZN(new_n914));
  INV_X1    g728(.A(new_n634), .ZN(new_n915));
  AOI21_X1  g729(.A(new_n895), .B1(new_n914), .B2(new_n915), .ZN(new_n916));
  NAND4_X1  g730(.A1(new_n910), .A2(new_n634), .A3(new_n911), .A4(new_n913), .ZN(new_n917));
  INV_X1    g731(.A(KEYINPUT121), .ZN(new_n918));
  NAND2_X1  g732(.A1(new_n917), .A2(new_n918), .ZN(new_n919));
  NAND4_X1  g733(.A1(new_n881), .A2(KEYINPUT121), .A3(new_n634), .A4(new_n913), .ZN(new_n920));
  AND3_X1   g734(.A1(new_n916), .A2(new_n919), .A3(new_n920), .ZN(G63));
  INV_X1    g735(.A(KEYINPUT61), .ZN(new_n922));
  NAND2_X1  g736(.A1(G217), .A2(G902), .ZN(new_n923));
  XNOR2_X1  g737(.A(new_n923), .B(KEYINPUT60), .ZN(new_n924));
  AOI21_X1  g738(.A(new_n924), .B1(new_n866), .B2(new_n878), .ZN(new_n925));
  AOI21_X1  g739(.A(new_n895), .B1(new_n925), .B2(new_n666), .ZN(new_n926));
  INV_X1    g740(.A(new_n924), .ZN(new_n927));
  AOI21_X1  g741(.A(KEYINPUT53), .B1(new_n876), .B2(new_n877), .ZN(new_n928));
  NOR4_X1   g742(.A1(new_n865), .A2(new_n872), .A3(new_n839), .A4(new_n875), .ZN(new_n929));
  OAI21_X1  g743(.A(new_n927), .B1(new_n928), .B2(new_n929), .ZN(new_n930));
  NAND2_X1  g744(.A1(new_n930), .A2(new_n226), .ZN(new_n931));
  AOI211_X1 g745(.A(KEYINPUT122), .B(new_n922), .C1(new_n926), .C2(new_n931), .ZN(new_n932));
  OAI211_X1 g746(.A(new_n666), .B(new_n927), .C1(new_n928), .C2(new_n929), .ZN(new_n933));
  INV_X1    g747(.A(new_n895), .ZN(new_n934));
  OAI211_X1 g748(.A(new_n933), .B(new_n934), .C1(new_n231), .C2(new_n925), .ZN(new_n935));
  INV_X1    g749(.A(KEYINPUT122), .ZN(new_n936));
  AOI21_X1  g750(.A(KEYINPUT61), .B1(new_n935), .B2(new_n936), .ZN(new_n937));
  NOR2_X1   g751(.A1(new_n932), .A2(new_n937), .ZN(G66));
  AOI21_X1  g752(.A(new_n188), .B1(new_n499), .B2(new_n465), .ZN(new_n939));
  INV_X1    g753(.A(new_n847), .ZN(new_n940));
  AOI21_X1  g754(.A(new_n939), .B1(new_n940), .B2(new_n188), .ZN(new_n941));
  MUX2_X1   g755(.A(new_n939), .B(new_n941), .S(KEYINPUT123), .Z(new_n942));
  OAI21_X1  g756(.A(new_n889), .B1(G898), .B2(new_n188), .ZN(new_n943));
  XOR2_X1   g757(.A(new_n942), .B(new_n943), .Z(G69));
  NOR4_X1   g758(.A1(new_n693), .A2(new_n844), .A3(new_n374), .A4(new_n790), .ZN(new_n945));
  AOI22_X1  g759(.A1(new_n776), .A2(new_n779), .B1(KEYINPUT124), .B2(new_n945), .ZN(new_n946));
  INV_X1    g760(.A(KEYINPUT62), .ZN(new_n947));
  INV_X1    g761(.A(new_n705), .ZN(new_n948));
  NAND2_X1  g762(.A1(new_n857), .A2(new_n738), .ZN(new_n949));
  OAI21_X1  g763(.A(new_n947), .B1(new_n948), .B2(new_n949), .ZN(new_n950));
  NAND4_X1  g764(.A1(new_n705), .A2(KEYINPUT62), .A3(new_n738), .A4(new_n857), .ZN(new_n951));
  NAND2_X1  g765(.A1(new_n950), .A2(new_n951), .ZN(new_n952));
  OR2_X1    g766(.A1(new_n945), .A2(KEYINPUT124), .ZN(new_n953));
  NAND4_X1  g767(.A1(new_n946), .A2(new_n952), .A3(new_n792), .A4(new_n953), .ZN(new_n954));
  NAND2_X1  g768(.A1(new_n954), .A2(new_n188), .ZN(new_n955));
  XNOR2_X1  g769(.A(new_n320), .B(new_n579), .ZN(new_n956));
  NAND2_X1  g770(.A1(new_n955), .A2(new_n956), .ZN(new_n957));
  INV_X1    g771(.A(new_n956), .ZN(new_n958));
  NAND2_X1  g772(.A1(G900), .A2(G953), .ZN(new_n959));
  INV_X1    g773(.A(new_n855), .ZN(new_n960));
  AOI21_X1  g774(.A(new_n960), .B1(new_n776), .B2(new_n779), .ZN(new_n961));
  INV_X1    g775(.A(new_n949), .ZN(new_n962));
  NOR2_X1   g776(.A1(new_n768), .A2(new_n691), .ZN(new_n963));
  NAND3_X1  g777(.A1(new_n963), .A2(new_n373), .A3(new_n860), .ZN(new_n964));
  NAND4_X1  g778(.A1(new_n961), .A2(new_n792), .A3(new_n962), .A4(new_n964), .ZN(new_n965));
  OAI211_X1 g779(.A(new_n958), .B(new_n959), .C1(new_n965), .C2(G953), .ZN(new_n966));
  NAND2_X1  g780(.A1(new_n957), .A2(new_n966), .ZN(new_n967));
  AOI21_X1  g781(.A(new_n188), .B1(G227), .B2(G900), .ZN(new_n968));
  NAND2_X1  g782(.A1(new_n967), .A2(new_n968), .ZN(new_n969));
  NAND2_X1  g783(.A1(new_n957), .A2(KEYINPUT125), .ZN(new_n970));
  INV_X1    g784(.A(KEYINPUT125), .ZN(new_n971));
  NAND3_X1  g785(.A1(new_n955), .A2(new_n971), .A3(new_n956), .ZN(new_n972));
  NAND3_X1  g786(.A1(new_n970), .A2(new_n966), .A3(new_n972), .ZN(new_n973));
  XNOR2_X1  g787(.A(new_n968), .B(KEYINPUT126), .ZN(new_n974));
  OAI21_X1  g788(.A(new_n969), .B1(new_n973), .B2(new_n974), .ZN(G72));
  NAND2_X1  g789(.A1(G472), .A2(G902), .ZN(new_n976));
  XOR2_X1   g790(.A(new_n976), .B(KEYINPUT63), .Z(new_n977));
  OAI21_X1  g791(.A(new_n977), .B1(new_n965), .B2(new_n940), .ZN(new_n978));
  NAND3_X1  g792(.A1(new_n978), .A2(new_n322), .A3(new_n337), .ZN(new_n979));
  OAI21_X1  g793(.A(new_n977), .B1(new_n954), .B2(new_n940), .ZN(new_n980));
  NAND2_X1  g794(.A1(new_n980), .A2(new_n699), .ZN(new_n981));
  NAND3_X1  g795(.A1(new_n979), .A2(new_n981), .A3(new_n934), .ZN(new_n982));
  NAND3_X1  g796(.A1(new_n329), .A2(new_n367), .A3(new_n339), .ZN(new_n983));
  NAND2_X1  g797(.A1(new_n983), .A2(new_n977), .ZN(new_n984));
  XOR2_X1   g798(.A(new_n984), .B(KEYINPUT127), .Z(new_n985));
  AOI21_X1  g799(.A(new_n982), .B1(new_n908), .B2(new_n985), .ZN(G57));
endmodule


