

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n523, n524, n525, n526,
         n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537,
         n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548,
         n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559,
         n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570,
         n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581,
         n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592,
         n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603,
         n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614,
         n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625,
         n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636,
         n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647,
         n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658,
         n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669,
         n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680,
         n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691,
         n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702,
         n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713,
         n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724,
         n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735,
         n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746,
         n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757,
         n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768,
         n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, n779,
         n780, n781, n782, n783, n784, n785, n786, n787, n788, n789, n790,
         n791, n792, n793, n794, n795, n796, n797, n798, n799, n800, n801,
         n802, n803, n804, n805, n806, n807, n808, n809, n810, n811, n812,
         n813, n814, n815, n816, n817, n818, n819, n820, n821, n822, n823,
         n824, n825, n826, n827, n828, n829, n830, n831, n832, n833, n834,
         n835, n836, n837, n838, n839, n840, n841, n842, n843, n844, n845,
         n846, n847, n848, n849, n850, n851, n852, n853, n854, n855, n856,
         n857, n858, n859, n860, n861, n862, n863, n864, n865, n866, n867,
         n868, n869, n870, n871, n872, n873, n874, n875, n876, n877, n878,
         n879, n880, n881, n882, n883, n884, n885, n886, n887, n888, n889,
         n890, n891, n892, n893, n894, n895, n896, n897, n898, n899, n900,
         n901, n902, n903, n904, n905, n906, n907, n908, n909, n910, n911,
         n912, n913, n914, n915, n916, n917, n918, n919, n920, n921, n922,
         n923, n924, n925, n926, n927, n928, n929, n930, n931, n932, n933,
         n934, n935, n936, n937, n938, n939, n940, n941, n942, n943, n944,
         n945, n946, n947, n948, n949, n950, n951, n952, n953, n954, n955,
         n956, n957, n958, n959, n960, n961, n962, n963, n964, n965, n966,
         n967, n968, n969, n970, n971, n972, n973, n974, n975, n976, n977,
         n978, n979, n980, n981, n982, n983, n984, n985, n986, n987, n988,
         n989, n990, n991, n992, n993, n994, n995, n996, n997, n998, n999,
         n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009,
         n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019,
         n1020, n1021;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NOR2_X1 U555 ( .A1(G2104), .A2(n530), .ZN(n886) );
  NAND2_X1 U556 ( .A1(n719), .A2(n718), .ZN(n758) );
  BUF_X1 U557 ( .A(n886), .Z(n523) );
  NOR2_X1 U558 ( .A1(n964), .A2(n724), .ZN(n731) );
  INV_X1 U559 ( .A(n758), .ZN(n725) );
  NOR2_X1 U560 ( .A1(n749), .A2(n748), .ZN(n750) );
  NAND2_X1 U561 ( .A1(n886), .A2(G126), .ZN(n524) );
  NOR2_X1 U562 ( .A1(G651), .A2(n637), .ZN(n657) );
  INV_X1 U563 ( .A(G2105), .ZN(n530) );
  XOR2_X1 U564 ( .A(n524), .B(KEYINPUT87), .Z(n526) );
  AND2_X1 U565 ( .A1(G2105), .A2(G2104), .ZN(n885) );
  NAND2_X1 U566 ( .A1(n885), .A2(G114), .ZN(n525) );
  NAND2_X1 U567 ( .A1(n526), .A2(n525), .ZN(n527) );
  XNOR2_X1 U568 ( .A(n527), .B(KEYINPUT88), .ZN(n534) );
  XNOR2_X1 U569 ( .A(KEYINPUT65), .B(KEYINPUT17), .ZN(n529) );
  NOR2_X1 U570 ( .A1(G2105), .A2(G2104), .ZN(n528) );
  XNOR2_X2 U571 ( .A(n529), .B(n528), .ZN(n891) );
  NAND2_X1 U572 ( .A1(G138), .A2(n891), .ZN(n532) );
  AND2_X1 U573 ( .A1(n530), .A2(G2104), .ZN(n889) );
  NAND2_X1 U574 ( .A1(G102), .A2(n889), .ZN(n531) );
  NAND2_X1 U575 ( .A1(n532), .A2(n531), .ZN(n533) );
  NOR2_X1 U576 ( .A1(n534), .A2(n533), .ZN(n535) );
  XOR2_X1 U577 ( .A(KEYINPUT89), .B(n535), .Z(G164) );
  NOR2_X1 U578 ( .A1(G651), .A2(G543), .ZN(n653) );
  NAND2_X1 U579 ( .A1(G91), .A2(n653), .ZN(n537) );
  XOR2_X1 U580 ( .A(KEYINPUT0), .B(G543), .Z(n637) );
  INV_X1 U581 ( .A(G651), .ZN(n538) );
  NOR2_X1 U582 ( .A1(n637), .A2(n538), .ZN(n649) );
  NAND2_X1 U583 ( .A1(G78), .A2(n649), .ZN(n536) );
  NAND2_X1 U584 ( .A1(n537), .A2(n536), .ZN(n542) );
  NOR2_X1 U585 ( .A1(G543), .A2(n538), .ZN(n539) );
  XOR2_X1 U586 ( .A(KEYINPUT1), .B(n539), .Z(n650) );
  NAND2_X1 U587 ( .A1(G65), .A2(n650), .ZN(n540) );
  XNOR2_X1 U588 ( .A(KEYINPUT69), .B(n540), .ZN(n541) );
  NOR2_X1 U589 ( .A1(n542), .A2(n541), .ZN(n544) );
  NAND2_X1 U590 ( .A1(n657), .A2(G53), .ZN(n543) );
  NAND2_X1 U591 ( .A1(n544), .A2(n543), .ZN(G299) );
  XNOR2_X1 U592 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  XOR2_X1 U593 ( .A(G2427), .B(G2435), .Z(n546) );
  XNOR2_X1 U594 ( .A(G2454), .B(G2443), .ZN(n545) );
  XNOR2_X1 U595 ( .A(n546), .B(n545), .ZN(n553) );
  XOR2_X1 U596 ( .A(G2451), .B(KEYINPUT105), .Z(n548) );
  XNOR2_X1 U597 ( .A(G2430), .B(G2438), .ZN(n547) );
  XNOR2_X1 U598 ( .A(n548), .B(n547), .ZN(n549) );
  XOR2_X1 U599 ( .A(n549), .B(G2446), .Z(n551) );
  XNOR2_X1 U600 ( .A(G1341), .B(G1348), .ZN(n550) );
  XNOR2_X1 U601 ( .A(n551), .B(n550), .ZN(n552) );
  XNOR2_X1 U602 ( .A(n553), .B(n552), .ZN(n554) );
  AND2_X1 U603 ( .A1(n554), .A2(G14), .ZN(G401) );
  AND2_X1 U604 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U605 ( .A(G57), .ZN(G237) );
  NAND2_X1 U606 ( .A1(n653), .A2(G89), .ZN(n555) );
  XNOR2_X1 U607 ( .A(n555), .B(KEYINPUT4), .ZN(n557) );
  NAND2_X1 U608 ( .A1(G76), .A2(n649), .ZN(n556) );
  NAND2_X1 U609 ( .A1(n557), .A2(n556), .ZN(n558) );
  XNOR2_X1 U610 ( .A(n558), .B(KEYINPUT5), .ZN(n563) );
  NAND2_X1 U611 ( .A1(G63), .A2(n650), .ZN(n560) );
  NAND2_X1 U612 ( .A1(G51), .A2(n657), .ZN(n559) );
  NAND2_X1 U613 ( .A1(n560), .A2(n559), .ZN(n561) );
  XOR2_X1 U614 ( .A(KEYINPUT6), .B(n561), .Z(n562) );
  NAND2_X1 U615 ( .A1(n563), .A2(n562), .ZN(n564) );
  XNOR2_X1 U616 ( .A(n564), .B(KEYINPUT7), .ZN(G168) );
  XNOR2_X1 U617 ( .A(G168), .B(KEYINPUT8), .ZN(n565) );
  XNOR2_X1 U618 ( .A(n565), .B(KEYINPUT75), .ZN(G286) );
  NAND2_X1 U619 ( .A1(G7), .A2(G661), .ZN(n566) );
  XNOR2_X1 U620 ( .A(n566), .B(KEYINPUT10), .ZN(n567) );
  XNOR2_X1 U621 ( .A(KEYINPUT70), .B(n567), .ZN(G223) );
  XOR2_X1 U622 ( .A(KEYINPUT11), .B(KEYINPUT72), .Z(n569) );
  XNOR2_X1 U623 ( .A(KEYINPUT71), .B(G223), .ZN(n833) );
  NAND2_X1 U624 ( .A1(n833), .A2(G567), .ZN(n568) );
  XNOR2_X1 U625 ( .A(n569), .B(n568), .ZN(G234) );
  NAND2_X1 U626 ( .A1(n650), .A2(G56), .ZN(n570) );
  XOR2_X1 U627 ( .A(KEYINPUT14), .B(n570), .Z(n577) );
  NAND2_X1 U628 ( .A1(n653), .A2(G81), .ZN(n571) );
  XNOR2_X1 U629 ( .A(n571), .B(KEYINPUT12), .ZN(n573) );
  NAND2_X1 U630 ( .A1(G68), .A2(n649), .ZN(n572) );
  NAND2_X1 U631 ( .A1(n573), .A2(n572), .ZN(n574) );
  XNOR2_X1 U632 ( .A(KEYINPUT13), .B(n574), .ZN(n575) );
  XNOR2_X1 U633 ( .A(KEYINPUT73), .B(n575), .ZN(n576) );
  NOR2_X1 U634 ( .A1(n577), .A2(n576), .ZN(n578) );
  XNOR2_X1 U635 ( .A(n578), .B(KEYINPUT74), .ZN(n580) );
  NAND2_X1 U636 ( .A1(G43), .A2(n657), .ZN(n579) );
  NAND2_X1 U637 ( .A1(n580), .A2(n579), .ZN(n964) );
  INV_X1 U638 ( .A(G860), .ZN(n619) );
  OR2_X1 U639 ( .A1(n964), .A2(n619), .ZN(G153) );
  NAND2_X1 U640 ( .A1(n653), .A2(G90), .ZN(n581) );
  XNOR2_X1 U641 ( .A(n581), .B(KEYINPUT68), .ZN(n583) );
  NAND2_X1 U642 ( .A1(G77), .A2(n649), .ZN(n582) );
  NAND2_X1 U643 ( .A1(n583), .A2(n582), .ZN(n584) );
  XNOR2_X1 U644 ( .A(n584), .B(KEYINPUT9), .ZN(n586) );
  NAND2_X1 U645 ( .A1(G64), .A2(n650), .ZN(n585) );
  NAND2_X1 U646 ( .A1(n586), .A2(n585), .ZN(n589) );
  NAND2_X1 U647 ( .A1(G52), .A2(n657), .ZN(n587) );
  XNOR2_X1 U648 ( .A(KEYINPUT67), .B(n587), .ZN(n588) );
  NOR2_X1 U649 ( .A1(n589), .A2(n588), .ZN(G171) );
  INV_X1 U650 ( .A(G171), .ZN(G301) );
  NAND2_X1 U651 ( .A1(G868), .A2(G301), .ZN(n598) );
  NAND2_X1 U652 ( .A1(G92), .A2(n653), .ZN(n591) );
  NAND2_X1 U653 ( .A1(G79), .A2(n649), .ZN(n590) );
  NAND2_X1 U654 ( .A1(n591), .A2(n590), .ZN(n595) );
  NAND2_X1 U655 ( .A1(G66), .A2(n650), .ZN(n593) );
  NAND2_X1 U656 ( .A1(G54), .A2(n657), .ZN(n592) );
  NAND2_X1 U657 ( .A1(n593), .A2(n592), .ZN(n594) );
  NOR2_X1 U658 ( .A1(n595), .A2(n594), .ZN(n596) );
  XOR2_X1 U659 ( .A(KEYINPUT15), .B(n596), .Z(n953) );
  OR2_X1 U660 ( .A1(n953), .A2(G868), .ZN(n597) );
  NAND2_X1 U661 ( .A1(n598), .A2(n597), .ZN(G284) );
  INV_X1 U662 ( .A(G868), .ZN(n668) );
  NOR2_X1 U663 ( .A1(G286), .A2(n668), .ZN(n600) );
  NOR2_X1 U664 ( .A1(G868), .A2(G299), .ZN(n599) );
  NOR2_X1 U665 ( .A1(n600), .A2(n599), .ZN(G297) );
  NAND2_X1 U666 ( .A1(n619), .A2(G559), .ZN(n601) );
  NAND2_X1 U667 ( .A1(n601), .A2(n953), .ZN(n602) );
  XNOR2_X1 U668 ( .A(n602), .B(KEYINPUT76), .ZN(n603) );
  XNOR2_X1 U669 ( .A(KEYINPUT16), .B(n603), .ZN(G148) );
  NOR2_X1 U670 ( .A1(G868), .A2(n964), .ZN(n606) );
  NAND2_X1 U671 ( .A1(G868), .A2(n953), .ZN(n604) );
  NOR2_X1 U672 ( .A1(G559), .A2(n604), .ZN(n605) );
  NOR2_X1 U673 ( .A1(n606), .A2(n605), .ZN(G282) );
  NAND2_X1 U674 ( .A1(G99), .A2(n889), .ZN(n608) );
  NAND2_X1 U675 ( .A1(G111), .A2(n885), .ZN(n607) );
  NAND2_X1 U676 ( .A1(n608), .A2(n607), .ZN(n609) );
  XNOR2_X1 U677 ( .A(KEYINPUT78), .B(n609), .ZN(n615) );
  NAND2_X1 U678 ( .A1(n523), .A2(G123), .ZN(n610) );
  XNOR2_X1 U679 ( .A(n610), .B(KEYINPUT18), .ZN(n612) );
  NAND2_X1 U680 ( .A1(G135), .A2(n891), .ZN(n611) );
  NAND2_X1 U681 ( .A1(n612), .A2(n611), .ZN(n613) );
  XOR2_X1 U682 ( .A(KEYINPUT77), .B(n613), .Z(n614) );
  NOR2_X1 U683 ( .A1(n615), .A2(n614), .ZN(n922) );
  XNOR2_X1 U684 ( .A(n922), .B(G2096), .ZN(n617) );
  INV_X1 U685 ( .A(G2100), .ZN(n616) );
  NAND2_X1 U686 ( .A1(n617), .A2(n616), .ZN(G156) );
  NAND2_X1 U687 ( .A1(G559), .A2(n953), .ZN(n618) );
  XOR2_X1 U688 ( .A(n964), .B(n618), .Z(n666) );
  NAND2_X1 U689 ( .A1(n619), .A2(n666), .ZN(n627) );
  NAND2_X1 U690 ( .A1(G93), .A2(n653), .ZN(n621) );
  NAND2_X1 U691 ( .A1(G67), .A2(n650), .ZN(n620) );
  NAND2_X1 U692 ( .A1(n621), .A2(n620), .ZN(n624) );
  NAND2_X1 U693 ( .A1(G80), .A2(n649), .ZN(n622) );
  XNOR2_X1 U694 ( .A(KEYINPUT79), .B(n622), .ZN(n623) );
  NOR2_X1 U695 ( .A1(n624), .A2(n623), .ZN(n626) );
  NAND2_X1 U696 ( .A1(n657), .A2(G55), .ZN(n625) );
  NAND2_X1 U697 ( .A1(n626), .A2(n625), .ZN(n669) );
  XNOR2_X1 U698 ( .A(n627), .B(n669), .ZN(G145) );
  NAND2_X1 U699 ( .A1(G73), .A2(n649), .ZN(n628) );
  XNOR2_X1 U700 ( .A(n628), .B(KEYINPUT2), .ZN(n635) );
  NAND2_X1 U701 ( .A1(G61), .A2(n650), .ZN(n630) );
  NAND2_X1 U702 ( .A1(G48), .A2(n657), .ZN(n629) );
  NAND2_X1 U703 ( .A1(n630), .A2(n629), .ZN(n633) );
  NAND2_X1 U704 ( .A1(n653), .A2(G86), .ZN(n631) );
  XOR2_X1 U705 ( .A(KEYINPUT80), .B(n631), .Z(n632) );
  NOR2_X1 U706 ( .A1(n633), .A2(n632), .ZN(n634) );
  NAND2_X1 U707 ( .A1(n635), .A2(n634), .ZN(n636) );
  XOR2_X1 U708 ( .A(KEYINPUT81), .B(n636), .Z(G305) );
  NAND2_X1 U709 ( .A1(G49), .A2(n657), .ZN(n639) );
  NAND2_X1 U710 ( .A1(G87), .A2(n637), .ZN(n638) );
  NAND2_X1 U711 ( .A1(n639), .A2(n638), .ZN(n640) );
  NOR2_X1 U712 ( .A1(n650), .A2(n640), .ZN(n642) );
  NAND2_X1 U713 ( .A1(G651), .A2(G74), .ZN(n641) );
  NAND2_X1 U714 ( .A1(n642), .A2(n641), .ZN(G288) );
  NAND2_X1 U715 ( .A1(G88), .A2(n653), .ZN(n644) );
  NAND2_X1 U716 ( .A1(G75), .A2(n649), .ZN(n643) );
  NAND2_X1 U717 ( .A1(n644), .A2(n643), .ZN(n648) );
  NAND2_X1 U718 ( .A1(G62), .A2(n650), .ZN(n646) );
  NAND2_X1 U719 ( .A1(G50), .A2(n657), .ZN(n645) );
  NAND2_X1 U720 ( .A1(n646), .A2(n645), .ZN(n647) );
  NOR2_X1 U721 ( .A1(n648), .A2(n647), .ZN(G166) );
  INV_X1 U722 ( .A(G166), .ZN(G303) );
  NAND2_X1 U723 ( .A1(G72), .A2(n649), .ZN(n652) );
  NAND2_X1 U724 ( .A1(G60), .A2(n650), .ZN(n651) );
  NAND2_X1 U725 ( .A1(n652), .A2(n651), .ZN(n656) );
  NAND2_X1 U726 ( .A1(n653), .A2(G85), .ZN(n654) );
  XOR2_X1 U727 ( .A(KEYINPUT66), .B(n654), .Z(n655) );
  NOR2_X1 U728 ( .A1(n656), .A2(n655), .ZN(n659) );
  NAND2_X1 U729 ( .A1(n657), .A2(G47), .ZN(n658) );
  NAND2_X1 U730 ( .A1(n659), .A2(n658), .ZN(G290) );
  INV_X1 U731 ( .A(G299), .ZN(n945) );
  XNOR2_X1 U732 ( .A(n945), .B(G305), .ZN(n660) );
  XNOR2_X1 U733 ( .A(n660), .B(n669), .ZN(n661) );
  XNOR2_X1 U734 ( .A(KEYINPUT19), .B(n661), .ZN(n663) );
  XNOR2_X1 U735 ( .A(G288), .B(KEYINPUT82), .ZN(n662) );
  XNOR2_X1 U736 ( .A(n663), .B(n662), .ZN(n664) );
  XNOR2_X1 U737 ( .A(n664), .B(G303), .ZN(n665) );
  XNOR2_X1 U738 ( .A(n665), .B(G290), .ZN(n903) );
  XOR2_X1 U739 ( .A(n903), .B(n666), .Z(n667) );
  NOR2_X1 U740 ( .A1(n668), .A2(n667), .ZN(n671) );
  NOR2_X1 U741 ( .A1(G868), .A2(n669), .ZN(n670) );
  NOR2_X1 U742 ( .A1(n671), .A2(n670), .ZN(G295) );
  NAND2_X1 U743 ( .A1(G2084), .A2(G2078), .ZN(n672) );
  XNOR2_X1 U744 ( .A(n672), .B(KEYINPUT20), .ZN(n673) );
  XNOR2_X1 U745 ( .A(KEYINPUT83), .B(n673), .ZN(n674) );
  NAND2_X1 U746 ( .A1(n674), .A2(G2090), .ZN(n675) );
  XNOR2_X1 U747 ( .A(KEYINPUT21), .B(n675), .ZN(n676) );
  NAND2_X1 U748 ( .A1(n676), .A2(G2072), .ZN(G158) );
  NAND2_X1 U749 ( .A1(G120), .A2(G69), .ZN(n677) );
  NOR2_X1 U750 ( .A1(G237), .A2(n677), .ZN(n678) );
  NAND2_X1 U751 ( .A1(G108), .A2(n678), .ZN(n838) );
  NAND2_X1 U752 ( .A1(G567), .A2(n838), .ZN(n679) );
  XNOR2_X1 U753 ( .A(n679), .B(KEYINPUT85), .ZN(n685) );
  XOR2_X1 U754 ( .A(KEYINPUT22), .B(KEYINPUT84), .Z(n681) );
  NAND2_X1 U755 ( .A1(G132), .A2(G82), .ZN(n680) );
  XNOR2_X1 U756 ( .A(n681), .B(n680), .ZN(n682) );
  NAND2_X1 U757 ( .A1(n682), .A2(G96), .ZN(n683) );
  OR2_X1 U758 ( .A1(G218), .A2(n683), .ZN(n839) );
  AND2_X1 U759 ( .A1(G2106), .A2(n839), .ZN(n684) );
  NOR2_X1 U760 ( .A1(n685), .A2(n684), .ZN(G319) );
  INV_X1 U761 ( .A(G319), .ZN(n687) );
  NAND2_X1 U762 ( .A1(G483), .A2(G661), .ZN(n686) );
  NOR2_X1 U763 ( .A1(n687), .A2(n686), .ZN(n837) );
  NAND2_X1 U764 ( .A1(n837), .A2(G36), .ZN(n688) );
  XNOR2_X1 U765 ( .A(KEYINPUT86), .B(n688), .ZN(G176) );
  XOR2_X1 U766 ( .A(KEYINPUT64), .B(KEYINPUT23), .Z(n690) );
  NAND2_X1 U767 ( .A1(G101), .A2(n889), .ZN(n689) );
  XNOR2_X1 U768 ( .A(n690), .B(n689), .ZN(n692) );
  NAND2_X1 U769 ( .A1(n891), .A2(G137), .ZN(n691) );
  NAND2_X1 U770 ( .A1(n692), .A2(n691), .ZN(n696) );
  NAND2_X1 U771 ( .A1(G113), .A2(n885), .ZN(n694) );
  NAND2_X1 U772 ( .A1(G125), .A2(n523), .ZN(n693) );
  NAND2_X1 U773 ( .A1(n694), .A2(n693), .ZN(n695) );
  NOR2_X1 U774 ( .A1(n696), .A2(n695), .ZN(G160) );
  NOR2_X1 U775 ( .A1(G164), .A2(G1384), .ZN(n718) );
  NAND2_X1 U776 ( .A1(G160), .A2(G40), .ZN(n717) );
  NOR2_X1 U777 ( .A1(n718), .A2(n717), .ZN(n828) );
  INV_X1 U778 ( .A(n828), .ZN(n716) );
  NAND2_X1 U779 ( .A1(G117), .A2(n885), .ZN(n698) );
  NAND2_X1 U780 ( .A1(G129), .A2(n523), .ZN(n697) );
  NAND2_X1 U781 ( .A1(n698), .A2(n697), .ZN(n701) );
  NAND2_X1 U782 ( .A1(n889), .A2(G105), .ZN(n699) );
  XOR2_X1 U783 ( .A(KEYINPUT38), .B(n699), .Z(n700) );
  NOR2_X1 U784 ( .A1(n701), .A2(n700), .ZN(n702) );
  XNOR2_X1 U785 ( .A(n702), .B(KEYINPUT94), .ZN(n704) );
  NAND2_X1 U786 ( .A1(G141), .A2(n891), .ZN(n703) );
  NAND2_X1 U787 ( .A1(n704), .A2(n703), .ZN(n881) );
  NAND2_X1 U788 ( .A1(G1996), .A2(n881), .ZN(n714) );
  NAND2_X1 U789 ( .A1(G107), .A2(n885), .ZN(n706) );
  NAND2_X1 U790 ( .A1(G119), .A2(n523), .ZN(n705) );
  NAND2_X1 U791 ( .A1(n706), .A2(n705), .ZN(n707) );
  XNOR2_X1 U792 ( .A(KEYINPUT92), .B(n707), .ZN(n710) );
  NAND2_X1 U793 ( .A1(G95), .A2(n889), .ZN(n708) );
  XNOR2_X1 U794 ( .A(KEYINPUT93), .B(n708), .ZN(n709) );
  NOR2_X1 U795 ( .A1(n710), .A2(n709), .ZN(n712) );
  NAND2_X1 U796 ( .A1(n891), .A2(G131), .ZN(n711) );
  NAND2_X1 U797 ( .A1(n712), .A2(n711), .ZN(n880) );
  NAND2_X1 U798 ( .A1(G1991), .A2(n880), .ZN(n713) );
  NAND2_X1 U799 ( .A1(n714), .A2(n713), .ZN(n921) );
  XNOR2_X1 U800 ( .A(G1986), .B(G290), .ZN(n948) );
  NOR2_X1 U801 ( .A1(n921), .A2(n948), .ZN(n715) );
  NOR2_X1 U802 ( .A1(n716), .A2(n715), .ZN(n805) );
  INV_X1 U803 ( .A(n717), .ZN(n719) );
  NAND2_X1 U804 ( .A1(n725), .A2(G1996), .ZN(n720) );
  XNOR2_X1 U805 ( .A(n720), .B(KEYINPUT26), .ZN(n723) );
  AND2_X1 U806 ( .A1(n758), .A2(G1341), .ZN(n721) );
  XNOR2_X1 U807 ( .A(KEYINPUT97), .B(n721), .ZN(n722) );
  NAND2_X1 U808 ( .A1(n723), .A2(n722), .ZN(n724) );
  NAND2_X1 U809 ( .A1(n731), .A2(n953), .ZN(n729) );
  NOR2_X1 U810 ( .A1(G2067), .A2(n758), .ZN(n727) );
  NOR2_X1 U811 ( .A1(n725), .A2(G1348), .ZN(n726) );
  NOR2_X1 U812 ( .A1(n727), .A2(n726), .ZN(n728) );
  NAND2_X1 U813 ( .A1(n729), .A2(n728), .ZN(n730) );
  XNOR2_X1 U814 ( .A(n730), .B(KEYINPUT98), .ZN(n733) );
  OR2_X1 U815 ( .A1(n731), .A2(n953), .ZN(n732) );
  NAND2_X1 U816 ( .A1(n733), .A2(n732), .ZN(n738) );
  NAND2_X1 U817 ( .A1(n725), .A2(G2072), .ZN(n734) );
  XNOR2_X1 U818 ( .A(n734), .B(KEYINPUT27), .ZN(n736) );
  AND2_X1 U819 ( .A1(G1956), .A2(n758), .ZN(n735) );
  NOR2_X1 U820 ( .A1(n736), .A2(n735), .ZN(n739) );
  NAND2_X1 U821 ( .A1(n945), .A2(n739), .ZN(n737) );
  NAND2_X1 U822 ( .A1(n738), .A2(n737), .ZN(n742) );
  NOR2_X1 U823 ( .A1(n945), .A2(n739), .ZN(n740) );
  XOR2_X1 U824 ( .A(n740), .B(KEYINPUT28), .Z(n741) );
  NAND2_X1 U825 ( .A1(n742), .A2(n741), .ZN(n743) );
  XNOR2_X1 U826 ( .A(KEYINPUT29), .B(n743), .ZN(n749) );
  XOR2_X1 U827 ( .A(G2078), .B(KEYINPUT25), .Z(n998) );
  NOR2_X1 U828 ( .A1(n998), .A2(n758), .ZN(n745) );
  NOR2_X1 U829 ( .A1(n725), .A2(G1961), .ZN(n744) );
  NOR2_X1 U830 ( .A1(n745), .A2(n744), .ZN(n746) );
  XOR2_X1 U831 ( .A(KEYINPUT95), .B(n746), .Z(n754) );
  NOR2_X1 U832 ( .A1(n754), .A2(G301), .ZN(n747) );
  XNOR2_X1 U833 ( .A(n747), .B(KEYINPUT96), .ZN(n748) );
  XNOR2_X1 U834 ( .A(KEYINPUT99), .B(n750), .ZN(n771) );
  NAND2_X1 U835 ( .A1(G8), .A2(n758), .ZN(n792) );
  NOR2_X1 U836 ( .A1(G1966), .A2(n792), .ZN(n774) );
  NOR2_X1 U837 ( .A1(G2084), .A2(n758), .ZN(n770) );
  NOR2_X1 U838 ( .A1(n774), .A2(n770), .ZN(n751) );
  NAND2_X1 U839 ( .A1(G8), .A2(n751), .ZN(n752) );
  XNOR2_X1 U840 ( .A(KEYINPUT30), .B(n752), .ZN(n753) );
  NOR2_X1 U841 ( .A1(G168), .A2(n753), .ZN(n756) );
  AND2_X1 U842 ( .A1(G301), .A2(n754), .ZN(n755) );
  NOR2_X1 U843 ( .A1(n756), .A2(n755), .ZN(n757) );
  XOR2_X1 U844 ( .A(KEYINPUT31), .B(n757), .Z(n772) );
  NOR2_X1 U845 ( .A1(G2090), .A2(n758), .ZN(n759) );
  XNOR2_X1 U846 ( .A(n759), .B(KEYINPUT100), .ZN(n761) );
  NOR2_X1 U847 ( .A1(n792), .A2(G1971), .ZN(n760) );
  NOR2_X1 U848 ( .A1(n761), .A2(n760), .ZN(n762) );
  NAND2_X1 U849 ( .A1(n762), .A2(G303), .ZN(n764) );
  AND2_X1 U850 ( .A1(n772), .A2(n764), .ZN(n763) );
  NAND2_X1 U851 ( .A1(n771), .A2(n763), .ZN(n768) );
  INV_X1 U852 ( .A(n764), .ZN(n765) );
  OR2_X1 U853 ( .A1(n765), .A2(G286), .ZN(n766) );
  AND2_X1 U854 ( .A1(G8), .A2(n766), .ZN(n767) );
  NAND2_X1 U855 ( .A1(n768), .A2(n767), .ZN(n769) );
  XNOR2_X1 U856 ( .A(n769), .B(KEYINPUT32), .ZN(n778) );
  NAND2_X1 U857 ( .A1(G8), .A2(n770), .ZN(n776) );
  AND2_X1 U858 ( .A1(n772), .A2(n771), .ZN(n773) );
  NOR2_X1 U859 ( .A1(n774), .A2(n773), .ZN(n775) );
  NAND2_X1 U860 ( .A1(n776), .A2(n775), .ZN(n777) );
  NAND2_X1 U861 ( .A1(n778), .A2(n777), .ZN(n788) );
  NOR2_X1 U862 ( .A1(G2090), .A2(G303), .ZN(n779) );
  NAND2_X1 U863 ( .A1(G8), .A2(n779), .ZN(n780) );
  NAND2_X1 U864 ( .A1(n788), .A2(n780), .ZN(n781) );
  AND2_X1 U865 ( .A1(n781), .A2(n792), .ZN(n785) );
  NOR2_X1 U866 ( .A1(G1981), .A2(G305), .ZN(n782) );
  XOR2_X1 U867 ( .A(n782), .B(KEYINPUT24), .Z(n783) );
  NOR2_X1 U868 ( .A1(n792), .A2(n783), .ZN(n784) );
  NOR2_X1 U869 ( .A1(n785), .A2(n784), .ZN(n803) );
  NOR2_X1 U870 ( .A1(G1976), .A2(G288), .ZN(n786) );
  XOR2_X1 U871 ( .A(KEYINPUT101), .B(n786), .Z(n790) );
  NOR2_X1 U872 ( .A1(G1971), .A2(G303), .ZN(n787) );
  NOR2_X1 U873 ( .A1(n790), .A2(n787), .ZN(n954) );
  NAND2_X1 U874 ( .A1(n788), .A2(n954), .ZN(n798) );
  INV_X1 U875 ( .A(n792), .ZN(n789) );
  NAND2_X1 U876 ( .A1(G1976), .A2(G288), .ZN(n944) );
  AND2_X1 U877 ( .A1(n789), .A2(n944), .ZN(n796) );
  NAND2_X1 U878 ( .A1(KEYINPUT33), .A2(n790), .ZN(n791) );
  NOR2_X1 U879 ( .A1(n792), .A2(n791), .ZN(n793) );
  XNOR2_X1 U880 ( .A(n793), .B(KEYINPUT102), .ZN(n795) );
  XOR2_X1 U881 ( .A(G1981), .B(G305), .Z(n957) );
  INV_X1 U882 ( .A(n957), .ZN(n794) );
  NOR2_X1 U883 ( .A1(n795), .A2(n794), .ZN(n799) );
  AND2_X1 U884 ( .A1(n796), .A2(n799), .ZN(n797) );
  AND2_X1 U885 ( .A1(n798), .A2(n797), .ZN(n801) );
  AND2_X1 U886 ( .A1(n799), .A2(KEYINPUT33), .ZN(n800) );
  NOR2_X1 U887 ( .A1(n801), .A2(n800), .ZN(n802) );
  AND2_X1 U888 ( .A1(n803), .A2(n802), .ZN(n804) );
  NOR2_X1 U889 ( .A1(n805), .A2(n804), .ZN(n817) );
  XNOR2_X1 U890 ( .A(G2067), .B(KEYINPUT37), .ZN(n824) );
  NAND2_X1 U891 ( .A1(n891), .A2(G140), .ZN(n806) );
  XNOR2_X1 U892 ( .A(n806), .B(KEYINPUT90), .ZN(n808) );
  NAND2_X1 U893 ( .A1(G104), .A2(n889), .ZN(n807) );
  NAND2_X1 U894 ( .A1(n808), .A2(n807), .ZN(n809) );
  XNOR2_X1 U895 ( .A(KEYINPUT34), .B(n809), .ZN(n815) );
  NAND2_X1 U896 ( .A1(n885), .A2(G116), .ZN(n810) );
  XOR2_X1 U897 ( .A(KEYINPUT91), .B(n810), .Z(n812) );
  NAND2_X1 U898 ( .A1(n523), .A2(G128), .ZN(n811) );
  NAND2_X1 U899 ( .A1(n812), .A2(n811), .ZN(n813) );
  XOR2_X1 U900 ( .A(KEYINPUT35), .B(n813), .Z(n814) );
  NOR2_X1 U901 ( .A1(n815), .A2(n814), .ZN(n816) );
  XNOR2_X1 U902 ( .A(KEYINPUT36), .B(n816), .ZN(n900) );
  NOR2_X1 U903 ( .A1(n824), .A2(n900), .ZN(n926) );
  NAND2_X1 U904 ( .A1(n926), .A2(n828), .ZN(n822) );
  NAND2_X1 U905 ( .A1(n817), .A2(n822), .ZN(n831) );
  NOR2_X1 U906 ( .A1(G1996), .A2(n881), .ZN(n931) );
  NOR2_X1 U907 ( .A1(G1986), .A2(G290), .ZN(n818) );
  NOR2_X1 U908 ( .A1(G1991), .A2(n880), .ZN(n920) );
  NOR2_X1 U909 ( .A1(n818), .A2(n920), .ZN(n819) );
  NOR2_X1 U910 ( .A1(n921), .A2(n819), .ZN(n820) );
  NOR2_X1 U911 ( .A1(n931), .A2(n820), .ZN(n821) );
  XNOR2_X1 U912 ( .A(n821), .B(KEYINPUT39), .ZN(n823) );
  NAND2_X1 U913 ( .A1(n823), .A2(n822), .ZN(n825) );
  NAND2_X1 U914 ( .A1(n824), .A2(n900), .ZN(n927) );
  NAND2_X1 U915 ( .A1(n825), .A2(n927), .ZN(n826) );
  XOR2_X1 U916 ( .A(KEYINPUT103), .B(n826), .Z(n827) );
  NAND2_X1 U917 ( .A1(n828), .A2(n827), .ZN(n829) );
  XNOR2_X1 U918 ( .A(n829), .B(KEYINPUT104), .ZN(n830) );
  NAND2_X1 U919 ( .A1(n831), .A2(n830), .ZN(n832) );
  XNOR2_X1 U920 ( .A(KEYINPUT40), .B(n832), .ZN(G329) );
  NAND2_X1 U921 ( .A1(G2106), .A2(n833), .ZN(G217) );
  NAND2_X1 U922 ( .A1(G15), .A2(G2), .ZN(n834) );
  XOR2_X1 U923 ( .A(KEYINPUT106), .B(n834), .Z(n835) );
  NAND2_X1 U924 ( .A1(G661), .A2(n835), .ZN(G259) );
  NAND2_X1 U925 ( .A1(G3), .A2(G1), .ZN(n836) );
  NAND2_X1 U926 ( .A1(n837), .A2(n836), .ZN(G188) );
  XNOR2_X1 U927 ( .A(G69), .B(KEYINPUT107), .ZN(G235) );
  INV_X1 U929 ( .A(G132), .ZN(G219) );
  INV_X1 U930 ( .A(G120), .ZN(G236) );
  INV_X1 U931 ( .A(G96), .ZN(G221) );
  INV_X1 U932 ( .A(G82), .ZN(G220) );
  NOR2_X1 U933 ( .A1(n839), .A2(n838), .ZN(n840) );
  XNOR2_X1 U934 ( .A(KEYINPUT108), .B(n840), .ZN(G325) );
  INV_X1 U935 ( .A(G325), .ZN(G261) );
  XOR2_X1 U936 ( .A(G1976), .B(G1981), .Z(n842) );
  XNOR2_X1 U937 ( .A(G1966), .B(G1971), .ZN(n841) );
  XNOR2_X1 U938 ( .A(n842), .B(n841), .ZN(n843) );
  XOR2_X1 U939 ( .A(n843), .B(G2474), .Z(n845) );
  XNOR2_X1 U940 ( .A(G1996), .B(G1991), .ZN(n844) );
  XNOR2_X1 U941 ( .A(n845), .B(n844), .ZN(n849) );
  XOR2_X1 U942 ( .A(KEYINPUT41), .B(G1986), .Z(n847) );
  XNOR2_X1 U943 ( .A(G1956), .B(G1961), .ZN(n846) );
  XNOR2_X1 U944 ( .A(n847), .B(n846), .ZN(n848) );
  XNOR2_X1 U945 ( .A(n849), .B(n848), .ZN(G229) );
  XOR2_X1 U946 ( .A(KEYINPUT42), .B(G2090), .Z(n851) );
  XNOR2_X1 U947 ( .A(G2072), .B(G2078), .ZN(n850) );
  XNOR2_X1 U948 ( .A(n851), .B(n850), .ZN(n852) );
  XOR2_X1 U949 ( .A(n852), .B(G2100), .Z(n854) );
  XNOR2_X1 U950 ( .A(G2067), .B(G2084), .ZN(n853) );
  XNOR2_X1 U951 ( .A(n854), .B(n853), .ZN(n858) );
  XOR2_X1 U952 ( .A(G2096), .B(KEYINPUT43), .Z(n856) );
  XNOR2_X1 U953 ( .A(KEYINPUT109), .B(G2678), .ZN(n855) );
  XNOR2_X1 U954 ( .A(n856), .B(n855), .ZN(n857) );
  XOR2_X1 U955 ( .A(n858), .B(n857), .Z(G227) );
  NAND2_X1 U956 ( .A1(G124), .A2(n523), .ZN(n859) );
  XNOR2_X1 U957 ( .A(n859), .B(KEYINPUT44), .ZN(n862) );
  NAND2_X1 U958 ( .A1(G112), .A2(n885), .ZN(n860) );
  XNOR2_X1 U959 ( .A(n860), .B(KEYINPUT110), .ZN(n861) );
  NAND2_X1 U960 ( .A1(n862), .A2(n861), .ZN(n866) );
  NAND2_X1 U961 ( .A1(G100), .A2(n889), .ZN(n864) );
  NAND2_X1 U962 ( .A1(G136), .A2(n891), .ZN(n863) );
  NAND2_X1 U963 ( .A1(n864), .A2(n863), .ZN(n865) );
  NOR2_X1 U964 ( .A1(n866), .A2(n865), .ZN(G162) );
  XOR2_X1 U965 ( .A(KEYINPUT46), .B(KEYINPUT113), .Z(n868) );
  XNOR2_X1 U966 ( .A(KEYINPUT114), .B(KEYINPUT48), .ZN(n867) );
  XNOR2_X1 U967 ( .A(n868), .B(n867), .ZN(n877) );
  NAND2_X1 U968 ( .A1(G103), .A2(n889), .ZN(n870) );
  NAND2_X1 U969 ( .A1(G139), .A2(n891), .ZN(n869) );
  NAND2_X1 U970 ( .A1(n870), .A2(n869), .ZN(n876) );
  NAND2_X1 U971 ( .A1(G115), .A2(n885), .ZN(n872) );
  NAND2_X1 U972 ( .A1(G127), .A2(n523), .ZN(n871) );
  NAND2_X1 U973 ( .A1(n872), .A2(n871), .ZN(n873) );
  XOR2_X1 U974 ( .A(KEYINPUT47), .B(n873), .Z(n874) );
  XNOR2_X1 U975 ( .A(KEYINPUT112), .B(n874), .ZN(n875) );
  NOR2_X1 U976 ( .A1(n876), .A2(n875), .ZN(n914) );
  XOR2_X1 U977 ( .A(n877), .B(n914), .Z(n879) );
  XNOR2_X1 U978 ( .A(G160), .B(G164), .ZN(n878) );
  XNOR2_X1 U979 ( .A(n879), .B(n878), .ZN(n884) );
  XNOR2_X1 U980 ( .A(G162), .B(n880), .ZN(n882) );
  XNOR2_X1 U981 ( .A(n882), .B(n881), .ZN(n883) );
  XOR2_X1 U982 ( .A(n884), .B(n883), .Z(n899) );
  NAND2_X1 U983 ( .A1(G118), .A2(n885), .ZN(n888) );
  NAND2_X1 U984 ( .A1(G130), .A2(n523), .ZN(n887) );
  NAND2_X1 U985 ( .A1(n888), .A2(n887), .ZN(n896) );
  NAND2_X1 U986 ( .A1(n889), .A2(G106), .ZN(n890) );
  XOR2_X1 U987 ( .A(KEYINPUT111), .B(n890), .Z(n893) );
  NAND2_X1 U988 ( .A1(n891), .A2(G142), .ZN(n892) );
  NAND2_X1 U989 ( .A1(n893), .A2(n892), .ZN(n894) );
  XOR2_X1 U990 ( .A(KEYINPUT45), .B(n894), .Z(n895) );
  NOR2_X1 U991 ( .A1(n896), .A2(n895), .ZN(n897) );
  XNOR2_X1 U992 ( .A(n922), .B(n897), .ZN(n898) );
  XNOR2_X1 U993 ( .A(n899), .B(n898), .ZN(n901) );
  XNOR2_X1 U994 ( .A(n901), .B(n900), .ZN(n902) );
  NOR2_X1 U995 ( .A1(G37), .A2(n902), .ZN(G395) );
  XOR2_X1 U996 ( .A(n903), .B(G286), .Z(n905) );
  XNOR2_X1 U997 ( .A(n953), .B(G171), .ZN(n904) );
  XNOR2_X1 U998 ( .A(n905), .B(n904), .ZN(n906) );
  XNOR2_X1 U999 ( .A(n906), .B(n964), .ZN(n907) );
  NOR2_X1 U1000 ( .A1(G37), .A2(n907), .ZN(G397) );
  NOR2_X1 U1001 ( .A1(G229), .A2(G227), .ZN(n908) );
  XOR2_X1 U1002 ( .A(KEYINPUT49), .B(n908), .Z(n909) );
  NAND2_X1 U1003 ( .A1(G319), .A2(n909), .ZN(n910) );
  NOR2_X1 U1004 ( .A1(G401), .A2(n910), .ZN(n913) );
  NOR2_X1 U1005 ( .A1(G395), .A2(G397), .ZN(n911) );
  XOR2_X1 U1006 ( .A(KEYINPUT115), .B(n911), .Z(n912) );
  NAND2_X1 U1007 ( .A1(n913), .A2(n912), .ZN(G225) );
  INV_X1 U1008 ( .A(G225), .ZN(G308) );
  INV_X1 U1009 ( .A(G108), .ZN(G238) );
  XNOR2_X1 U1010 ( .A(KEYINPUT118), .B(KEYINPUT50), .ZN(n918) );
  XNOR2_X1 U1011 ( .A(G2072), .B(n914), .ZN(n916) );
  XNOR2_X1 U1012 ( .A(G164), .B(G2078), .ZN(n915) );
  NAND2_X1 U1013 ( .A1(n916), .A2(n915), .ZN(n917) );
  XNOR2_X1 U1014 ( .A(n918), .B(n917), .ZN(n937) );
  XOR2_X1 U1015 ( .A(G2084), .B(G160), .Z(n919) );
  NOR2_X1 U1016 ( .A1(n920), .A2(n919), .ZN(n924) );
  NOR2_X1 U1017 ( .A1(n922), .A2(n921), .ZN(n923) );
  NAND2_X1 U1018 ( .A1(n924), .A2(n923), .ZN(n925) );
  NOR2_X1 U1019 ( .A1(n926), .A2(n925), .ZN(n928) );
  NAND2_X1 U1020 ( .A1(n928), .A2(n927), .ZN(n934) );
  XOR2_X1 U1021 ( .A(G2090), .B(G162), .Z(n929) );
  XNOR2_X1 U1022 ( .A(KEYINPUT116), .B(n929), .ZN(n930) );
  NOR2_X1 U1023 ( .A1(n931), .A2(n930), .ZN(n932) );
  XNOR2_X1 U1024 ( .A(KEYINPUT51), .B(n932), .ZN(n933) );
  NOR2_X1 U1025 ( .A1(n934), .A2(n933), .ZN(n935) );
  XNOR2_X1 U1026 ( .A(n935), .B(KEYINPUT117), .ZN(n936) );
  NOR2_X1 U1027 ( .A1(n937), .A2(n936), .ZN(n938) );
  XNOR2_X1 U1028 ( .A(KEYINPUT52), .B(n938), .ZN(n940) );
  INV_X1 U1029 ( .A(KEYINPUT55), .ZN(n939) );
  NAND2_X1 U1030 ( .A1(n940), .A2(n939), .ZN(n941) );
  NAND2_X1 U1031 ( .A1(n941), .A2(G29), .ZN(n942) );
  XNOR2_X1 U1032 ( .A(KEYINPUT119), .B(n942), .ZN(n1020) );
  NAND2_X1 U1033 ( .A1(G1971), .A2(G303), .ZN(n943) );
  NAND2_X1 U1034 ( .A1(n944), .A2(n943), .ZN(n952) );
  XNOR2_X1 U1035 ( .A(G1956), .B(n945), .ZN(n946) );
  XNOR2_X1 U1036 ( .A(n946), .B(KEYINPUT122), .ZN(n950) );
  XNOR2_X1 U1037 ( .A(G1961), .B(G301), .ZN(n947) );
  NOR2_X1 U1038 ( .A1(n948), .A2(n947), .ZN(n949) );
  NAND2_X1 U1039 ( .A1(n950), .A2(n949), .ZN(n951) );
  NOR2_X1 U1040 ( .A1(n952), .A2(n951), .ZN(n963) );
  XNOR2_X1 U1041 ( .A(n953), .B(G1348), .ZN(n955) );
  NAND2_X1 U1042 ( .A1(n955), .A2(n954), .ZN(n961) );
  XOR2_X1 U1043 ( .A(G1966), .B(G168), .Z(n956) );
  XNOR2_X1 U1044 ( .A(KEYINPUT121), .B(n956), .ZN(n958) );
  NAND2_X1 U1045 ( .A1(n958), .A2(n957), .ZN(n959) );
  XOR2_X1 U1046 ( .A(KEYINPUT57), .B(n959), .Z(n960) );
  NOR2_X1 U1047 ( .A1(n961), .A2(n960), .ZN(n962) );
  NAND2_X1 U1048 ( .A1(n963), .A2(n962), .ZN(n966) );
  XNOR2_X1 U1049 ( .A(G1341), .B(n964), .ZN(n965) );
  NOR2_X1 U1050 ( .A1(n966), .A2(n965), .ZN(n968) );
  XOR2_X1 U1051 ( .A(KEYINPUT56), .B(G16), .Z(n967) );
  NOR2_X1 U1052 ( .A1(n968), .A2(n967), .ZN(n1017) );
  XNOR2_X1 U1053 ( .A(G1348), .B(KEYINPUT59), .ZN(n969) );
  XNOR2_X1 U1054 ( .A(n969), .B(G4), .ZN(n973) );
  XNOR2_X1 U1055 ( .A(G1341), .B(G19), .ZN(n971) );
  XNOR2_X1 U1056 ( .A(G6), .B(G1981), .ZN(n970) );
  NOR2_X1 U1057 ( .A1(n971), .A2(n970), .ZN(n972) );
  NAND2_X1 U1058 ( .A1(n973), .A2(n972), .ZN(n976) );
  XOR2_X1 U1059 ( .A(KEYINPUT123), .B(G1956), .Z(n974) );
  XNOR2_X1 U1060 ( .A(G20), .B(n974), .ZN(n975) );
  NOR2_X1 U1061 ( .A1(n976), .A2(n975), .ZN(n977) );
  XNOR2_X1 U1062 ( .A(KEYINPUT60), .B(n977), .ZN(n978) );
  XNOR2_X1 U1063 ( .A(n978), .B(KEYINPUT124), .ZN(n982) );
  XNOR2_X1 U1064 ( .A(G1966), .B(G21), .ZN(n980) );
  XNOR2_X1 U1065 ( .A(G5), .B(G1961), .ZN(n979) );
  NOR2_X1 U1066 ( .A1(n980), .A2(n979), .ZN(n981) );
  NAND2_X1 U1067 ( .A1(n982), .A2(n981), .ZN(n991) );
  XNOR2_X1 U1068 ( .A(G1971), .B(G22), .ZN(n984) );
  XNOR2_X1 U1069 ( .A(G24), .B(G1986), .ZN(n983) );
  NOR2_X1 U1070 ( .A1(n984), .A2(n983), .ZN(n987) );
  XNOR2_X1 U1071 ( .A(G1976), .B(KEYINPUT125), .ZN(n985) );
  XNOR2_X1 U1072 ( .A(n985), .B(G23), .ZN(n986) );
  NAND2_X1 U1073 ( .A1(n987), .A2(n986), .ZN(n988) );
  XOR2_X1 U1074 ( .A(KEYINPUT58), .B(n988), .Z(n989) );
  XOR2_X1 U1075 ( .A(KEYINPUT126), .B(n989), .Z(n990) );
  NOR2_X1 U1076 ( .A1(n991), .A2(n990), .ZN(n992) );
  XOR2_X1 U1077 ( .A(KEYINPUT61), .B(n992), .Z(n993) );
  NOR2_X1 U1078 ( .A1(G16), .A2(n993), .ZN(n1014) );
  XNOR2_X1 U1079 ( .A(G2084), .B(G34), .ZN(n994) );
  XNOR2_X1 U1080 ( .A(n994), .B(KEYINPUT54), .ZN(n1010) );
  XNOR2_X1 U1081 ( .A(G2090), .B(G35), .ZN(n1007) );
  XOR2_X1 U1082 ( .A(G1991), .B(G25), .Z(n995) );
  NAND2_X1 U1083 ( .A1(n995), .A2(G28), .ZN(n1004) );
  XNOR2_X1 U1084 ( .A(G1996), .B(G32), .ZN(n997) );
  XNOR2_X1 U1085 ( .A(G33), .B(G2072), .ZN(n996) );
  NOR2_X1 U1086 ( .A1(n997), .A2(n996), .ZN(n1002) );
  XNOR2_X1 U1087 ( .A(G2067), .B(G26), .ZN(n1000) );
  XNOR2_X1 U1088 ( .A(G27), .B(n998), .ZN(n999) );
  NOR2_X1 U1089 ( .A1(n1000), .A2(n999), .ZN(n1001) );
  NAND2_X1 U1090 ( .A1(n1002), .A2(n1001), .ZN(n1003) );
  NOR2_X1 U1091 ( .A1(n1004), .A2(n1003), .ZN(n1005) );
  XNOR2_X1 U1092 ( .A(KEYINPUT53), .B(n1005), .ZN(n1006) );
  NOR2_X1 U1093 ( .A1(n1007), .A2(n1006), .ZN(n1008) );
  XOR2_X1 U1094 ( .A(KEYINPUT120), .B(n1008), .Z(n1009) );
  NOR2_X1 U1095 ( .A1(n1010), .A2(n1009), .ZN(n1011) );
  XOR2_X1 U1096 ( .A(KEYINPUT55), .B(n1011), .Z(n1012) );
  NOR2_X1 U1097 ( .A1(G29), .A2(n1012), .ZN(n1013) );
  NOR2_X1 U1098 ( .A1(n1014), .A2(n1013), .ZN(n1015) );
  NAND2_X1 U1099 ( .A1(G11), .A2(n1015), .ZN(n1016) );
  NOR2_X1 U1100 ( .A1(n1017), .A2(n1016), .ZN(n1018) );
  XNOR2_X1 U1101 ( .A(n1018), .B(KEYINPUT127), .ZN(n1019) );
  NOR2_X1 U1102 ( .A1(n1020), .A2(n1019), .ZN(n1021) );
  XNOR2_X1 U1103 ( .A(KEYINPUT62), .B(n1021), .ZN(G311) );
  INV_X1 U1104 ( .A(G311), .ZN(G150) );
endmodule

