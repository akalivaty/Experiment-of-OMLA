

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303,
         n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314,
         n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325,
         n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336,
         n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347,
         n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358,
         n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369,
         n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380,
         n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391,
         n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402,
         n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413,
         n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424,
         n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435,
         n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446,
         n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457,
         n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468,
         n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479,
         n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490,
         n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501,
         n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512,
         n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589,
         n590, n591;

  XNOR2_X1 U325 ( .A(n370), .B(n369), .ZN(n517) );
  XOR2_X1 U326 ( .A(G92GAT), .B(n425), .Z(n293) );
  INV_X1 U327 ( .A(KEYINPUT25), .ZN(n408) );
  XNOR2_X1 U328 ( .A(n409), .B(n408), .ZN(n410) );
  XNOR2_X1 U329 ( .A(KEYINPUT69), .B(KEYINPUT8), .ZN(n300) );
  XNOR2_X1 U330 ( .A(n308), .B(n307), .ZN(n309) );
  XNOR2_X1 U331 ( .A(n310), .B(n309), .ZN(n311) );
  NOR2_X1 U332 ( .A1(n414), .A2(n413), .ZN(n415) );
  NOR2_X1 U333 ( .A1(n589), .A2(n416), .ZN(n418) );
  XOR2_X1 U334 ( .A(KEYINPUT36), .B(n557), .Z(n589) );
  NOR2_X1 U335 ( .A1(n570), .A2(n569), .ZN(n572) );
  XNOR2_X1 U336 ( .A(n455), .B(KEYINPUT38), .ZN(n499) );
  XNOR2_X1 U337 ( .A(G43GAT), .B(KEYINPUT40), .ZN(n456) );
  XNOR2_X1 U338 ( .A(n457), .B(n456), .ZN(G1330GAT) );
  XOR2_X1 U339 ( .A(KEYINPUT79), .B(KEYINPUT10), .Z(n295) );
  XNOR2_X1 U340 ( .A(G99GAT), .B(KEYINPUT77), .ZN(n294) );
  XNOR2_X1 U341 ( .A(n295), .B(n294), .ZN(n316) );
  INV_X1 U342 ( .A(KEYINPUT7), .ZN(n296) );
  NAND2_X1 U343 ( .A1(G29GAT), .A2(n296), .ZN(n299) );
  INV_X1 U344 ( .A(G29GAT), .ZN(n297) );
  NAND2_X1 U345 ( .A1(n297), .A2(KEYINPUT7), .ZN(n298) );
  NAND2_X1 U346 ( .A1(n299), .A2(n298), .ZN(n301) );
  XNOR2_X1 U347 ( .A(n301), .B(n300), .ZN(n425) );
  NAND2_X1 U348 ( .A1(G232GAT), .A2(G233GAT), .ZN(n302) );
  XNOR2_X1 U349 ( .A(n293), .B(n302), .ZN(n310) );
  XOR2_X1 U350 ( .A(KEYINPUT66), .B(G85GAT), .Z(n304) );
  XNOR2_X1 U351 ( .A(G218GAT), .B(G106GAT), .ZN(n303) );
  XNOR2_X1 U352 ( .A(n304), .B(n303), .ZN(n308) );
  XOR2_X1 U353 ( .A(KEYINPUT78), .B(KEYINPUT65), .Z(n306) );
  XNOR2_X1 U354 ( .A(KEYINPUT11), .B(KEYINPUT9), .ZN(n305) );
  XNOR2_X1 U355 ( .A(n306), .B(n305), .ZN(n307) );
  XOR2_X1 U356 ( .A(G36GAT), .B(G190GAT), .Z(n357) );
  XOR2_X1 U357 ( .A(n311), .B(n357), .Z(n314) );
  XOR2_X1 U358 ( .A(G43GAT), .B(G134GAT), .Z(n390) );
  XNOR2_X1 U359 ( .A(G50GAT), .B(KEYINPUT76), .ZN(n312) );
  XNOR2_X1 U360 ( .A(n312), .B(G162GAT), .ZN(n376) );
  XNOR2_X1 U361 ( .A(n390), .B(n376), .ZN(n313) );
  XNOR2_X1 U362 ( .A(n314), .B(n313), .ZN(n315) );
  XNOR2_X1 U363 ( .A(n316), .B(n315), .ZN(n557) );
  XOR2_X1 U364 ( .A(G8GAT), .B(G211GAT), .Z(n354) );
  XOR2_X1 U365 ( .A(G57GAT), .B(KEYINPUT13), .Z(n445) );
  XOR2_X1 U366 ( .A(n354), .B(n445), .Z(n318) );
  XOR2_X1 U367 ( .A(G1GAT), .B(KEYINPUT70), .Z(n422) );
  XOR2_X1 U368 ( .A(G15GAT), .B(G127GAT), .Z(n389) );
  XNOR2_X1 U369 ( .A(n422), .B(n389), .ZN(n317) );
  XNOR2_X1 U370 ( .A(n318), .B(n317), .ZN(n323) );
  XNOR2_X1 U371 ( .A(G22GAT), .B(G155GAT), .ZN(n319) );
  XNOR2_X1 U372 ( .A(n319), .B(G78GAT), .ZN(n381) );
  XOR2_X1 U373 ( .A(n381), .B(KEYINPUT82), .Z(n321) );
  NAND2_X1 U374 ( .A1(G231GAT), .A2(G233GAT), .ZN(n320) );
  XNOR2_X1 U375 ( .A(n321), .B(n320), .ZN(n322) );
  XOR2_X1 U376 ( .A(n323), .B(n322), .Z(n331) );
  XOR2_X1 U377 ( .A(KEYINPUT12), .B(G64GAT), .Z(n325) );
  XNOR2_X1 U378 ( .A(G183GAT), .B(G71GAT), .ZN(n324) );
  XNOR2_X1 U379 ( .A(n325), .B(n324), .ZN(n329) );
  XOR2_X1 U380 ( .A(KEYINPUT15), .B(KEYINPUT14), .Z(n327) );
  XNOR2_X1 U381 ( .A(KEYINPUT81), .B(KEYINPUT80), .ZN(n326) );
  XNOR2_X1 U382 ( .A(n327), .B(n326), .ZN(n328) );
  XNOR2_X1 U383 ( .A(n329), .B(n328), .ZN(n330) );
  XOR2_X1 U384 ( .A(n331), .B(n330), .Z(n553) );
  INV_X1 U385 ( .A(n553), .ZN(n586) );
  XOR2_X1 U386 ( .A(KEYINPUT93), .B(KEYINPUT5), .Z(n333) );
  XNOR2_X1 U387 ( .A(G1GAT), .B(KEYINPUT91), .ZN(n332) );
  XNOR2_X1 U388 ( .A(n333), .B(n332), .ZN(n338) );
  XNOR2_X1 U389 ( .A(G141GAT), .B(KEYINPUT3), .ZN(n334) );
  XNOR2_X1 U390 ( .A(n334), .B(KEYINPUT2), .ZN(n373) );
  XOR2_X1 U391 ( .A(n373), .B(KEYINPUT4), .Z(n336) );
  NAND2_X1 U392 ( .A1(G225GAT), .A2(G233GAT), .ZN(n335) );
  XNOR2_X1 U393 ( .A(n336), .B(n335), .ZN(n337) );
  XNOR2_X1 U394 ( .A(n338), .B(n337), .ZN(n353) );
  XOR2_X1 U395 ( .A(G148GAT), .B(G155GAT), .Z(n340) );
  XNOR2_X1 U396 ( .A(G127GAT), .B(G120GAT), .ZN(n339) );
  XNOR2_X1 U397 ( .A(n340), .B(n339), .ZN(n344) );
  XOR2_X1 U398 ( .A(KEYINPUT92), .B(G57GAT), .Z(n342) );
  XNOR2_X1 U399 ( .A(KEYINPUT6), .B(KEYINPUT1), .ZN(n341) );
  XNOR2_X1 U400 ( .A(n342), .B(n341), .ZN(n343) );
  XOR2_X1 U401 ( .A(n344), .B(n343), .Z(n351) );
  XOR2_X1 U402 ( .A(G85GAT), .B(G162GAT), .Z(n348) );
  XOR2_X1 U403 ( .A(KEYINPUT84), .B(KEYINPUT0), .Z(n346) );
  XNOR2_X1 U404 ( .A(G113GAT), .B(KEYINPUT83), .ZN(n345) );
  XNOR2_X1 U405 ( .A(n346), .B(n345), .ZN(n395) );
  XNOR2_X1 U406 ( .A(G29GAT), .B(n395), .ZN(n347) );
  XNOR2_X1 U407 ( .A(n348), .B(n347), .ZN(n349) );
  XNOR2_X1 U408 ( .A(G134GAT), .B(n349), .ZN(n350) );
  XNOR2_X1 U409 ( .A(n351), .B(n350), .ZN(n352) );
  XNOR2_X1 U410 ( .A(n353), .B(n352), .ZN(n544) );
  XNOR2_X1 U411 ( .A(n354), .B(KEYINPUT94), .ZN(n355) );
  XNOR2_X1 U412 ( .A(n355), .B(KEYINPUT95), .ZN(n356) );
  XOR2_X1 U413 ( .A(n357), .B(n356), .Z(n359) );
  NAND2_X1 U414 ( .A1(G226GAT), .A2(G233GAT), .ZN(n358) );
  XNOR2_X1 U415 ( .A(n359), .B(n358), .ZN(n361) );
  XNOR2_X1 U416 ( .A(G204GAT), .B(G92GAT), .ZN(n360) );
  XNOR2_X1 U417 ( .A(n360), .B(G64GAT), .ZN(n444) );
  XOR2_X1 U418 ( .A(n361), .B(n444), .Z(n370) );
  XOR2_X1 U419 ( .A(KEYINPUT85), .B(KEYINPUT17), .Z(n363) );
  XNOR2_X1 U420 ( .A(KEYINPUT18), .B(KEYINPUT19), .ZN(n362) );
  XNOR2_X1 U421 ( .A(n363), .B(n362), .ZN(n364) );
  XOR2_X1 U422 ( .A(n364), .B(G183GAT), .Z(n366) );
  XNOR2_X1 U423 ( .A(G169GAT), .B(G176GAT), .ZN(n365) );
  XNOR2_X1 U424 ( .A(n366), .B(n365), .ZN(n401) );
  XOR2_X1 U425 ( .A(KEYINPUT89), .B(KEYINPUT21), .Z(n368) );
  XNOR2_X1 U426 ( .A(G197GAT), .B(G218GAT), .ZN(n367) );
  XNOR2_X1 U427 ( .A(n368), .B(n367), .ZN(n382) );
  XNOR2_X1 U428 ( .A(n401), .B(n382), .ZN(n369) );
  XOR2_X1 U429 ( .A(n517), .B(KEYINPUT27), .Z(n404) );
  XNOR2_X1 U430 ( .A(KEYINPUT28), .B(KEYINPUT67), .ZN(n387) );
  XOR2_X1 U431 ( .A(KEYINPUT88), .B(KEYINPUT24), .Z(n372) );
  XNOR2_X1 U432 ( .A(KEYINPUT23), .B(KEYINPUT22), .ZN(n371) );
  XNOR2_X1 U433 ( .A(n372), .B(n371), .ZN(n386) );
  XOR2_X1 U434 ( .A(G106GAT), .B(G148GAT), .Z(n450) );
  XOR2_X1 U435 ( .A(n450), .B(n373), .Z(n375) );
  XNOR2_X1 U436 ( .A(KEYINPUT90), .B(G204GAT), .ZN(n374) );
  XNOR2_X1 U437 ( .A(n375), .B(n374), .ZN(n380) );
  XOR2_X1 U438 ( .A(G211GAT), .B(n376), .Z(n378) );
  NAND2_X1 U439 ( .A1(G228GAT), .A2(G233GAT), .ZN(n377) );
  XNOR2_X1 U440 ( .A(n378), .B(n377), .ZN(n379) );
  XOR2_X1 U441 ( .A(n380), .B(n379), .Z(n384) );
  XNOR2_X1 U442 ( .A(n382), .B(n381), .ZN(n383) );
  XNOR2_X1 U443 ( .A(n384), .B(n383), .ZN(n385) );
  XNOR2_X1 U444 ( .A(n386), .B(n385), .ZN(n473) );
  XNOR2_X1 U445 ( .A(n387), .B(n473), .ZN(n522) );
  NOR2_X1 U446 ( .A1(n404), .A2(n522), .ZN(n388) );
  NAND2_X1 U447 ( .A1(n544), .A2(n388), .ZN(n528) );
  XNOR2_X1 U448 ( .A(n390), .B(n389), .ZN(n399) );
  XOR2_X1 U449 ( .A(KEYINPUT86), .B(KEYINPUT20), .Z(n392) );
  NAND2_X1 U450 ( .A1(G227GAT), .A2(G233GAT), .ZN(n391) );
  XNOR2_X1 U451 ( .A(n392), .B(n391), .ZN(n393) );
  XOR2_X1 U452 ( .A(n393), .B(G190GAT), .Z(n397) );
  XNOR2_X1 U453 ( .A(G99GAT), .B(G71GAT), .ZN(n394) );
  XNOR2_X1 U454 ( .A(n394), .B(G120GAT), .ZN(n446) );
  XNOR2_X1 U455 ( .A(n395), .B(n446), .ZN(n396) );
  XNOR2_X1 U456 ( .A(n397), .B(n396), .ZN(n398) );
  XNOR2_X1 U457 ( .A(n399), .B(n398), .ZN(n400) );
  XNOR2_X1 U458 ( .A(n401), .B(n400), .ZN(n530) );
  XOR2_X1 U459 ( .A(KEYINPUT87), .B(n530), .Z(n402) );
  NOR2_X1 U460 ( .A1(n528), .A2(n402), .ZN(n414) );
  NOR2_X1 U461 ( .A1(n530), .A2(n473), .ZN(n403) );
  XNOR2_X1 U462 ( .A(KEYINPUT26), .B(n403), .ZN(n576) );
  INV_X1 U463 ( .A(n576), .ZN(n405) );
  NOR2_X1 U464 ( .A1(n405), .A2(n404), .ZN(n543) );
  NAND2_X1 U465 ( .A1(n517), .A2(n530), .ZN(n406) );
  XNOR2_X1 U466 ( .A(n406), .B(KEYINPUT96), .ZN(n407) );
  NAND2_X1 U467 ( .A1(n407), .A2(n473), .ZN(n409) );
  XNOR2_X1 U468 ( .A(KEYINPUT97), .B(n410), .ZN(n411) );
  NOR2_X1 U469 ( .A1(n543), .A2(n411), .ZN(n412) );
  NOR2_X1 U470 ( .A1(n544), .A2(n412), .ZN(n413) );
  XOR2_X1 U471 ( .A(KEYINPUT98), .B(n415), .Z(n482) );
  NAND2_X1 U472 ( .A1(n586), .A2(n482), .ZN(n416) );
  XNOR2_X1 U473 ( .A(KEYINPUT102), .B(KEYINPUT37), .ZN(n417) );
  XNOR2_X1 U474 ( .A(n418), .B(n417), .ZN(n513) );
  XOR2_X1 U475 ( .A(G141GAT), .B(G22GAT), .Z(n420) );
  XNOR2_X1 U476 ( .A(G36GAT), .B(G197GAT), .ZN(n419) );
  XNOR2_X1 U477 ( .A(n420), .B(n419), .ZN(n421) );
  XOR2_X1 U478 ( .A(n421), .B(G43GAT), .Z(n424) );
  XNOR2_X1 U479 ( .A(n422), .B(G50GAT), .ZN(n423) );
  XNOR2_X1 U480 ( .A(n424), .B(n423), .ZN(n429) );
  XOR2_X1 U481 ( .A(n425), .B(KEYINPUT29), .Z(n427) );
  NAND2_X1 U482 ( .A1(G229GAT), .A2(G233GAT), .ZN(n426) );
  XNOR2_X1 U483 ( .A(n427), .B(n426), .ZN(n428) );
  XOR2_X1 U484 ( .A(n429), .B(n428), .Z(n437) );
  XOR2_X1 U485 ( .A(G8GAT), .B(G15GAT), .Z(n431) );
  XNOR2_X1 U486 ( .A(G169GAT), .B(G113GAT), .ZN(n430) );
  XNOR2_X1 U487 ( .A(n431), .B(n430), .ZN(n435) );
  XOR2_X1 U488 ( .A(KEYINPUT72), .B(KEYINPUT71), .Z(n433) );
  XNOR2_X1 U489 ( .A(KEYINPUT68), .B(KEYINPUT30), .ZN(n432) );
  XNOR2_X1 U490 ( .A(n433), .B(n432), .ZN(n434) );
  XNOR2_X1 U491 ( .A(n435), .B(n434), .ZN(n436) );
  XOR2_X1 U492 ( .A(n437), .B(n436), .Z(n546) );
  XOR2_X1 U493 ( .A(KEYINPUT73), .B(G85GAT), .Z(n439) );
  XNOR2_X1 U494 ( .A(G176GAT), .B(G78GAT), .ZN(n438) );
  XNOR2_X1 U495 ( .A(n439), .B(n438), .ZN(n443) );
  XOR2_X1 U496 ( .A(KEYINPUT74), .B(KEYINPUT33), .Z(n441) );
  XNOR2_X1 U497 ( .A(KEYINPUT75), .B(KEYINPUT32), .ZN(n440) );
  XNOR2_X1 U498 ( .A(n441), .B(n440), .ZN(n442) );
  XNOR2_X1 U499 ( .A(n443), .B(n442), .ZN(n454) );
  XOR2_X1 U500 ( .A(n445), .B(n444), .Z(n452) );
  XOR2_X1 U501 ( .A(n446), .B(KEYINPUT31), .Z(n448) );
  NAND2_X1 U502 ( .A1(G230GAT), .A2(G233GAT), .ZN(n447) );
  XNOR2_X1 U503 ( .A(n448), .B(n447), .ZN(n449) );
  XNOR2_X1 U504 ( .A(n450), .B(n449), .ZN(n451) );
  XNOR2_X1 U505 ( .A(n452), .B(n451), .ZN(n453) );
  XOR2_X1 U506 ( .A(n454), .B(n453), .Z(n583) );
  NAND2_X1 U507 ( .A1(n546), .A2(n583), .ZN(n484) );
  NOR2_X1 U508 ( .A1(n513), .A2(n484), .ZN(n455) );
  NAND2_X1 U509 ( .A1(n499), .A2(n530), .ZN(n457) );
  INV_X1 U510 ( .A(n546), .ZN(n578) );
  XOR2_X1 U511 ( .A(KEYINPUT121), .B(KEYINPUT55), .Z(n476) );
  INV_X1 U512 ( .A(n557), .ZN(n570) );
  XNOR2_X1 U513 ( .A(n553), .B(KEYINPUT112), .ZN(n565) );
  XNOR2_X1 U514 ( .A(n583), .B(KEYINPUT64), .ZN(n459) );
  INV_X1 U515 ( .A(KEYINPUT41), .ZN(n458) );
  XNOR2_X1 U516 ( .A(n459), .B(n458), .ZN(n559) );
  NOR2_X1 U517 ( .A1(n578), .A2(n559), .ZN(n460) );
  XNOR2_X1 U518 ( .A(n460), .B(KEYINPUT46), .ZN(n461) );
  NOR2_X1 U519 ( .A1(n565), .A2(n461), .ZN(n462) );
  NAND2_X1 U520 ( .A1(n570), .A2(n462), .ZN(n463) );
  XNOR2_X1 U521 ( .A(n463), .B(KEYINPUT47), .ZN(n469) );
  NOR2_X1 U522 ( .A1(n586), .A2(n589), .ZN(n465) );
  XOR2_X1 U523 ( .A(KEYINPUT45), .B(KEYINPUT113), .Z(n464) );
  XNOR2_X1 U524 ( .A(n465), .B(n464), .ZN(n466) );
  NAND2_X1 U525 ( .A1(n466), .A2(n583), .ZN(n467) );
  NOR2_X1 U526 ( .A1(n546), .A2(n467), .ZN(n468) );
  NOR2_X1 U527 ( .A1(n469), .A2(n468), .ZN(n470) );
  XNOR2_X1 U528 ( .A(n470), .B(KEYINPUT48), .ZN(n527) );
  XOR2_X1 U529 ( .A(KEYINPUT120), .B(n517), .Z(n471) );
  NOR2_X1 U530 ( .A1(n527), .A2(n471), .ZN(n472) );
  XNOR2_X1 U531 ( .A(n472), .B(KEYINPUT54), .ZN(n574) );
  INV_X1 U532 ( .A(n544), .ZN(n575) );
  AND2_X1 U533 ( .A1(n575), .A2(n473), .ZN(n474) );
  NAND2_X1 U534 ( .A1(n574), .A2(n474), .ZN(n475) );
  XNOR2_X1 U535 ( .A(n476), .B(n475), .ZN(n477) );
  NAND2_X1 U536 ( .A1(n477), .A2(n530), .ZN(n569) );
  NOR2_X1 U537 ( .A1(n578), .A2(n569), .ZN(n478) );
  XNOR2_X1 U538 ( .A(G169GAT), .B(n478), .ZN(n480) );
  INV_X1 U539 ( .A(KEYINPUT122), .ZN(n479) );
  XNOR2_X1 U540 ( .A(n480), .B(n479), .ZN(G1348GAT) );
  NOR2_X1 U541 ( .A1(n586), .A2(n557), .ZN(n481) );
  XNOR2_X1 U542 ( .A(KEYINPUT16), .B(n481), .ZN(n483) );
  NAND2_X1 U543 ( .A1(n483), .A2(n482), .ZN(n501) );
  NOR2_X1 U544 ( .A1(n484), .A2(n501), .ZN(n492) );
  NAND2_X1 U545 ( .A1(n492), .A2(n544), .ZN(n485) );
  XNOR2_X1 U546 ( .A(n485), .B(KEYINPUT34), .ZN(n486) );
  XNOR2_X1 U547 ( .A(G1GAT), .B(n486), .ZN(G1324GAT) );
  XOR2_X1 U548 ( .A(G8GAT), .B(KEYINPUT99), .Z(n488) );
  NAND2_X1 U549 ( .A1(n492), .A2(n517), .ZN(n487) );
  XNOR2_X1 U550 ( .A(n488), .B(n487), .ZN(G1325GAT) );
  XOR2_X1 U551 ( .A(KEYINPUT100), .B(KEYINPUT35), .Z(n490) );
  NAND2_X1 U552 ( .A1(n492), .A2(n530), .ZN(n489) );
  XNOR2_X1 U553 ( .A(n490), .B(n489), .ZN(n491) );
  XNOR2_X1 U554 ( .A(G15GAT), .B(n491), .ZN(G1326GAT) );
  XOR2_X1 U555 ( .A(G22GAT), .B(KEYINPUT101), .Z(n494) );
  NAND2_X1 U556 ( .A1(n492), .A2(n522), .ZN(n493) );
  XNOR2_X1 U557 ( .A(n494), .B(n493), .ZN(G1327GAT) );
  XOR2_X1 U558 ( .A(G29GAT), .B(KEYINPUT39), .Z(n496) );
  NAND2_X1 U559 ( .A1(n544), .A2(n499), .ZN(n495) );
  XNOR2_X1 U560 ( .A(n496), .B(n495), .ZN(G1328GAT) );
  XOR2_X1 U561 ( .A(G36GAT), .B(KEYINPUT103), .Z(n498) );
  NAND2_X1 U562 ( .A1(n517), .A2(n499), .ZN(n497) );
  XNOR2_X1 U563 ( .A(n498), .B(n497), .ZN(G1329GAT) );
  NAND2_X1 U564 ( .A1(n499), .A2(n522), .ZN(n500) );
  XNOR2_X1 U565 ( .A(n500), .B(G50GAT), .ZN(G1331GAT) );
  XNOR2_X1 U566 ( .A(G57GAT), .B(KEYINPUT42), .ZN(n503) );
  INV_X1 U567 ( .A(n559), .ZN(n549) );
  NAND2_X1 U568 ( .A1(n578), .A2(n549), .ZN(n512) );
  NOR2_X1 U569 ( .A1(n512), .A2(n501), .ZN(n508) );
  NAND2_X1 U570 ( .A1(n544), .A2(n508), .ZN(n502) );
  XNOR2_X1 U571 ( .A(n503), .B(n502), .ZN(G1332GAT) );
  XOR2_X1 U572 ( .A(KEYINPUT104), .B(KEYINPUT105), .Z(n505) );
  NAND2_X1 U573 ( .A1(n508), .A2(n517), .ZN(n504) );
  XNOR2_X1 U574 ( .A(n505), .B(n504), .ZN(n506) );
  XNOR2_X1 U575 ( .A(G64GAT), .B(n506), .ZN(G1333GAT) );
  NAND2_X1 U576 ( .A1(n530), .A2(n508), .ZN(n507) );
  XNOR2_X1 U577 ( .A(n507), .B(G71GAT), .ZN(G1334GAT) );
  XOR2_X1 U578 ( .A(KEYINPUT43), .B(KEYINPUT106), .Z(n510) );
  NAND2_X1 U579 ( .A1(n508), .A2(n522), .ZN(n509) );
  XNOR2_X1 U580 ( .A(n510), .B(n509), .ZN(n511) );
  XNOR2_X1 U581 ( .A(G78GAT), .B(n511), .ZN(G1335GAT) );
  XOR2_X1 U582 ( .A(KEYINPUT107), .B(KEYINPUT108), .Z(n515) );
  NOR2_X1 U583 ( .A1(n513), .A2(n512), .ZN(n523) );
  NAND2_X1 U584 ( .A1(n523), .A2(n544), .ZN(n514) );
  XNOR2_X1 U585 ( .A(n515), .B(n514), .ZN(n516) );
  XNOR2_X1 U586 ( .A(G85GAT), .B(n516), .ZN(G1336GAT) );
  XOR2_X1 U587 ( .A(G92GAT), .B(KEYINPUT109), .Z(n519) );
  NAND2_X1 U588 ( .A1(n523), .A2(n517), .ZN(n518) );
  XNOR2_X1 U589 ( .A(n519), .B(n518), .ZN(G1337GAT) );
  NAND2_X1 U590 ( .A1(n530), .A2(n523), .ZN(n520) );
  XNOR2_X1 U591 ( .A(n520), .B(KEYINPUT110), .ZN(n521) );
  XNOR2_X1 U592 ( .A(G99GAT), .B(n521), .ZN(G1338GAT) );
  XOR2_X1 U593 ( .A(KEYINPUT44), .B(KEYINPUT111), .Z(n525) );
  NAND2_X1 U594 ( .A1(n523), .A2(n522), .ZN(n524) );
  XNOR2_X1 U595 ( .A(n525), .B(n524), .ZN(n526) );
  XNOR2_X1 U596 ( .A(G106GAT), .B(n526), .ZN(G1339GAT) );
  XOR2_X1 U597 ( .A(G113GAT), .B(KEYINPUT115), .Z(n533) );
  NOR2_X1 U598 ( .A1(n527), .A2(n528), .ZN(n529) );
  NAND2_X1 U599 ( .A1(n530), .A2(n529), .ZN(n531) );
  XOR2_X1 U600 ( .A(KEYINPUT114), .B(n531), .Z(n539) );
  NAND2_X1 U601 ( .A1(n539), .A2(n546), .ZN(n532) );
  XNOR2_X1 U602 ( .A(n533), .B(n532), .ZN(G1340GAT) );
  XOR2_X1 U603 ( .A(KEYINPUT49), .B(KEYINPUT116), .Z(n535) );
  NAND2_X1 U604 ( .A1(n539), .A2(n549), .ZN(n534) );
  XNOR2_X1 U605 ( .A(n535), .B(n534), .ZN(n536) );
  XNOR2_X1 U606 ( .A(G120GAT), .B(n536), .ZN(G1341GAT) );
  NAND2_X1 U607 ( .A1(n539), .A2(n565), .ZN(n537) );
  XNOR2_X1 U608 ( .A(n537), .B(KEYINPUT50), .ZN(n538) );
  XNOR2_X1 U609 ( .A(G127GAT), .B(n538), .ZN(G1342GAT) );
  XOR2_X1 U610 ( .A(KEYINPUT117), .B(KEYINPUT51), .Z(n541) );
  NAND2_X1 U611 ( .A1(n539), .A2(n557), .ZN(n540) );
  XNOR2_X1 U612 ( .A(n541), .B(n540), .ZN(n542) );
  XOR2_X1 U613 ( .A(G134GAT), .B(n542), .Z(G1343GAT) );
  NAND2_X1 U614 ( .A1(n544), .A2(n543), .ZN(n545) );
  NOR2_X1 U615 ( .A1(n527), .A2(n545), .ZN(n556) );
  NAND2_X1 U616 ( .A1(n546), .A2(n556), .ZN(n547) );
  XNOR2_X1 U617 ( .A(n547), .B(KEYINPUT118), .ZN(n548) );
  XNOR2_X1 U618 ( .A(G141GAT), .B(n548), .ZN(G1344GAT) );
  XOR2_X1 U619 ( .A(KEYINPUT53), .B(KEYINPUT52), .Z(n551) );
  NAND2_X1 U620 ( .A1(n556), .A2(n549), .ZN(n550) );
  XNOR2_X1 U621 ( .A(n551), .B(n550), .ZN(n552) );
  XNOR2_X1 U622 ( .A(G148GAT), .B(n552), .ZN(G1345GAT) );
  XOR2_X1 U623 ( .A(G155GAT), .B(KEYINPUT119), .Z(n555) );
  NAND2_X1 U624 ( .A1(n556), .A2(n553), .ZN(n554) );
  XNOR2_X1 U625 ( .A(n555), .B(n554), .ZN(G1346GAT) );
  NAND2_X1 U626 ( .A1(n557), .A2(n556), .ZN(n558) );
  XNOR2_X1 U627 ( .A(n558), .B(G162GAT), .ZN(G1347GAT) );
  NOR2_X1 U628 ( .A1(n559), .A2(n569), .ZN(n564) );
  XOR2_X1 U629 ( .A(KEYINPUT57), .B(KEYINPUT124), .Z(n561) );
  XNOR2_X1 U630 ( .A(G176GAT), .B(KEYINPUT56), .ZN(n560) );
  XNOR2_X1 U631 ( .A(n561), .B(n560), .ZN(n562) );
  XNOR2_X1 U632 ( .A(KEYINPUT123), .B(n562), .ZN(n563) );
  XNOR2_X1 U633 ( .A(n564), .B(n563), .ZN(G1349GAT) );
  XOR2_X1 U634 ( .A(G183GAT), .B(KEYINPUT125), .Z(n568) );
  INV_X1 U635 ( .A(n569), .ZN(n566) );
  NAND2_X1 U636 ( .A1(n566), .A2(n565), .ZN(n567) );
  XNOR2_X1 U637 ( .A(n568), .B(n567), .ZN(G1350GAT) );
  XNOR2_X1 U638 ( .A(KEYINPUT126), .B(KEYINPUT58), .ZN(n571) );
  XNOR2_X1 U639 ( .A(n572), .B(n571), .ZN(n573) );
  XOR2_X1 U640 ( .A(G190GAT), .B(n573), .Z(G1351GAT) );
  AND2_X1 U641 ( .A1(n575), .A2(n574), .ZN(n577) );
  NAND2_X1 U642 ( .A1(n577), .A2(n576), .ZN(n588) );
  NOR2_X1 U643 ( .A1(n588), .A2(n578), .ZN(n582) );
  XOR2_X1 U644 ( .A(KEYINPUT59), .B(KEYINPUT127), .Z(n580) );
  XNOR2_X1 U645 ( .A(G197GAT), .B(KEYINPUT60), .ZN(n579) );
  XNOR2_X1 U646 ( .A(n580), .B(n579), .ZN(n581) );
  XNOR2_X1 U647 ( .A(n582), .B(n581), .ZN(G1352GAT) );
  NOR2_X1 U648 ( .A1(n583), .A2(n588), .ZN(n585) );
  XNOR2_X1 U649 ( .A(G204GAT), .B(KEYINPUT61), .ZN(n584) );
  XNOR2_X1 U650 ( .A(n585), .B(n584), .ZN(G1353GAT) );
  NOR2_X1 U651 ( .A1(n586), .A2(n588), .ZN(n587) );
  XOR2_X1 U652 ( .A(G211GAT), .B(n587), .Z(G1354GAT) );
  NOR2_X1 U653 ( .A1(n589), .A2(n588), .ZN(n590) );
  XOR2_X1 U654 ( .A(KEYINPUT62), .B(n590), .Z(n591) );
  XNOR2_X1 U655 ( .A(G218GAT), .B(n591), .ZN(G1355GAT) );
endmodule

