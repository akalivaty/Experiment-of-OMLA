//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 0 0 1 1 1 0 1 1 0 0 1 0 1 0 0 0 0 0 1 0 1 0 0 0 1 1 0 1 1 0 0 0 0 1 1 1 0 1 1 1 0 1 1 0 1 1 0 0 0 1 0 0 1 1 1 1 0 0 0 1 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:28:23 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n442, new_n443, new_n444, new_n446, new_n450, new_n452, new_n455,
    new_n456, new_n457, new_n460, new_n461, new_n462, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n528, new_n529, new_n530, new_n531, new_n532, new_n533,
    new_n534, new_n535, new_n536, new_n537, new_n538, new_n539, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n561, new_n563, new_n564, new_n566, new_n567,
    new_n568, new_n569, new_n570, new_n571, new_n572, new_n573, new_n574,
    new_n575, new_n578, new_n579, new_n580, new_n581, new_n582, new_n584,
    new_n585, new_n586, new_n587, new_n588, new_n589, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n616,
    new_n619, new_n620, new_n622, new_n623, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n824, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1183, new_n1184,
    new_n1185;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  XNOR2_X1  g013(.A(KEYINPUT64), .B(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  XOR2_X1   g015(.A(KEYINPUT65), .B(G108), .Z(G238));
  INV_X1    g016(.A(G2072), .ZN(new_n442));
  INV_X1    g017(.A(G2078), .ZN(new_n443));
  NOR2_X1   g018(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  NAND3_X1  g019(.A1(new_n444), .A2(G2084), .A3(G2090), .ZN(G158));
  NAND3_X1  g020(.A1(G2), .A2(G15), .A3(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT66), .Z(G259));
  BUF_X1    g022(.A(G452), .Z(G391));
  AND2_X1   g023(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g024(.A1(G7), .A2(G661), .ZN(new_n450));
  XOR2_X1   g025(.A(new_n450), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g026(.A1(G7), .A2(G567), .A3(G661), .ZN(new_n452));
  XOR2_X1   g027(.A(new_n452), .B(KEYINPUT67), .Z(G234));
  NAND3_X1  g028(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g029(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n455));
  XOR2_X1   g030(.A(new_n455), .B(KEYINPUT2), .Z(new_n456));
  OR4_X1    g031(.A1(G237), .A2(G238), .A3(G235), .A4(G236), .ZN(new_n457));
  NOR2_X1   g032(.A1(new_n456), .A2(new_n457), .ZN(G325));
  INV_X1    g033(.A(G325), .ZN(G261));
  NAND2_X1  g034(.A1(new_n456), .A2(G2106), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n457), .A2(G567), .ZN(new_n461));
  NAND2_X1  g036(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  INV_X1    g037(.A(new_n462), .ZN(G319));
  INV_X1    g038(.A(G2105), .ZN(new_n464));
  AND2_X1   g039(.A1(new_n464), .A2(G2104), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n465), .A2(G101), .ZN(new_n466));
  XNOR2_X1  g041(.A(KEYINPUT3), .B(G2104), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n467), .A2(new_n464), .ZN(new_n468));
  INV_X1    g043(.A(G137), .ZN(new_n469));
  OAI21_X1  g044(.A(new_n466), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  AND2_X1   g045(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n471));
  NOR2_X1   g046(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n472));
  OAI21_X1  g047(.A(G125), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  INV_X1    g048(.A(KEYINPUT68), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n473), .A2(new_n474), .ZN(new_n475));
  OAI211_X1 g050(.A(KEYINPUT68), .B(G125), .C1(new_n471), .C2(new_n472), .ZN(new_n476));
  NAND2_X1  g051(.A1(G113), .A2(G2104), .ZN(new_n477));
  NAND3_X1  g052(.A1(new_n475), .A2(new_n476), .A3(new_n477), .ZN(new_n478));
  AOI21_X1  g053(.A(new_n470), .B1(new_n478), .B2(G2105), .ZN(G160));
  OR2_X1    g054(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n480));
  NAND2_X1  g055(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n481));
  AOI21_X1  g056(.A(G2105), .B1(new_n480), .B2(new_n481), .ZN(new_n482));
  NAND2_X1  g057(.A1(new_n482), .A2(G136), .ZN(new_n483));
  AOI21_X1  g058(.A(new_n464), .B1(new_n480), .B2(new_n481), .ZN(new_n484));
  NAND2_X1  g059(.A1(new_n484), .A2(G124), .ZN(new_n485));
  OR2_X1    g060(.A1(G100), .A2(G2105), .ZN(new_n486));
  OAI211_X1 g061(.A(new_n486), .B(G2104), .C1(G112), .C2(new_n464), .ZN(new_n487));
  NAND3_X1  g062(.A1(new_n483), .A2(new_n485), .A3(new_n487), .ZN(new_n488));
  INV_X1    g063(.A(new_n488), .ZN(G162));
  INV_X1    g064(.A(G138), .ZN(new_n490));
  NOR2_X1   g065(.A1(new_n490), .A2(G2105), .ZN(new_n491));
  INV_X1    g066(.A(KEYINPUT4), .ZN(new_n492));
  OAI211_X1 g067(.A(new_n491), .B(new_n492), .C1(new_n472), .C2(new_n471), .ZN(new_n493));
  INV_X1    g068(.A(new_n493), .ZN(new_n494));
  AOI21_X1  g069(.A(new_n492), .B1(new_n467), .B2(new_n491), .ZN(new_n495));
  NOR2_X1   g070(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  OR2_X1    g071(.A1(new_n464), .A2(G114), .ZN(new_n497));
  OAI21_X1  g072(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n498));
  INV_X1    g073(.A(new_n498), .ZN(new_n499));
  NAND2_X1  g074(.A1(new_n497), .A2(new_n499), .ZN(new_n500));
  NAND2_X1  g075(.A1(new_n467), .A2(G2105), .ZN(new_n501));
  INV_X1    g076(.A(G126), .ZN(new_n502));
  OAI21_X1  g077(.A(new_n500), .B1(new_n501), .B2(new_n502), .ZN(new_n503));
  OAI21_X1  g078(.A(KEYINPUT69), .B1(new_n496), .B2(new_n503), .ZN(new_n504));
  OAI21_X1  g079(.A(new_n491), .B1(new_n471), .B2(new_n472), .ZN(new_n505));
  NAND2_X1  g080(.A1(new_n505), .A2(KEYINPUT4), .ZN(new_n506));
  NAND2_X1  g081(.A1(new_n506), .A2(new_n493), .ZN(new_n507));
  INV_X1    g082(.A(KEYINPUT69), .ZN(new_n508));
  AOI22_X1  g083(.A1(new_n484), .A2(G126), .B1(new_n497), .B2(new_n499), .ZN(new_n509));
  NAND3_X1  g084(.A1(new_n507), .A2(new_n508), .A3(new_n509), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n504), .A2(new_n510), .ZN(new_n511));
  INV_X1    g086(.A(new_n511), .ZN(G164));
  XNOR2_X1  g087(.A(KEYINPUT5), .B(G543), .ZN(new_n513));
  AOI22_X1  g088(.A1(new_n513), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n514));
  INV_X1    g089(.A(G651), .ZN(new_n515));
  OR2_X1    g090(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  INV_X1    g091(.A(G50), .ZN(new_n517));
  XNOR2_X1  g092(.A(KEYINPUT6), .B(G651), .ZN(new_n518));
  NAND2_X1  g093(.A1(new_n518), .A2(G543), .ZN(new_n519));
  NAND2_X1  g094(.A1(new_n518), .A2(new_n513), .ZN(new_n520));
  NAND2_X1  g095(.A1(new_n520), .A2(KEYINPUT70), .ZN(new_n521));
  INV_X1    g096(.A(KEYINPUT70), .ZN(new_n522));
  NAND3_X1  g097(.A1(new_n518), .A2(new_n513), .A3(new_n522), .ZN(new_n523));
  NAND2_X1  g098(.A1(new_n521), .A2(new_n523), .ZN(new_n524));
  INV_X1    g099(.A(G88), .ZN(new_n525));
  OAI221_X1 g100(.A(new_n516), .B1(new_n517), .B2(new_n519), .C1(new_n524), .C2(new_n525), .ZN(G303));
  INV_X1    g101(.A(G303), .ZN(G166));
  AND2_X1   g102(.A1(new_n518), .A2(G543), .ZN(new_n528));
  XOR2_X1   g103(.A(KEYINPUT71), .B(KEYINPUT7), .Z(new_n529));
  NAND3_X1  g104(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n530));
  NAND2_X1  g105(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  XNOR2_X1  g106(.A(KEYINPUT71), .B(KEYINPUT7), .ZN(new_n532));
  INV_X1    g107(.A(new_n530), .ZN(new_n533));
  NAND2_X1  g108(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  AOI22_X1  g109(.A1(G51), .A2(new_n528), .B1(new_n531), .B2(new_n534), .ZN(new_n535));
  NAND3_X1  g110(.A1(new_n513), .A2(G63), .A3(G651), .ZN(new_n536));
  NAND2_X1  g111(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  NAND3_X1  g112(.A1(new_n521), .A2(G89), .A3(new_n523), .ZN(new_n538));
  INV_X1    g113(.A(new_n538), .ZN(new_n539));
  NOR2_X1   g114(.A1(new_n537), .A2(new_n539), .ZN(G168));
  NAND3_X1  g115(.A1(new_n521), .A2(G90), .A3(new_n523), .ZN(new_n541));
  NAND2_X1  g116(.A1(new_n528), .A2(G52), .ZN(new_n542));
  NAND2_X1  g117(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  INV_X1    g118(.A(KEYINPUT72), .ZN(new_n544));
  NAND2_X1  g119(.A1(new_n543), .A2(new_n544), .ZN(new_n545));
  NAND3_X1  g120(.A1(new_n541), .A2(KEYINPUT72), .A3(new_n542), .ZN(new_n546));
  NAND2_X1  g121(.A1(new_n545), .A2(new_n546), .ZN(new_n547));
  AOI22_X1  g122(.A1(new_n513), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n548));
  OR2_X1    g123(.A1(new_n548), .A2(new_n515), .ZN(new_n549));
  NAND2_X1  g124(.A1(new_n547), .A2(new_n549), .ZN(G301));
  INV_X1    g125(.A(G301), .ZN(G171));
  NAND2_X1  g126(.A1(G68), .A2(G543), .ZN(new_n552));
  XOR2_X1   g127(.A(KEYINPUT5), .B(G543), .Z(new_n553));
  INV_X1    g128(.A(G56), .ZN(new_n554));
  OAI21_X1  g129(.A(new_n552), .B1(new_n553), .B2(new_n554), .ZN(new_n555));
  AOI22_X1  g130(.A1(new_n555), .A2(G651), .B1(new_n528), .B2(G43), .ZN(new_n556));
  INV_X1    g131(.A(G81), .ZN(new_n557));
  OAI21_X1  g132(.A(new_n556), .B1(new_n557), .B2(new_n524), .ZN(new_n558));
  INV_X1    g133(.A(new_n558), .ZN(new_n559));
  NAND2_X1  g134(.A1(new_n559), .A2(G860), .ZN(G153));
  NAND4_X1  g135(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(new_n561));
  XNOR2_X1  g136(.A(new_n561), .B(KEYINPUT73), .ZN(G176));
  NAND2_X1  g137(.A1(G1), .A2(G3), .ZN(new_n563));
  XNOR2_X1  g138(.A(new_n563), .B(KEYINPUT8), .ZN(new_n564));
  NAND4_X1  g139(.A1(G319), .A2(G483), .A3(G661), .A4(new_n564), .ZN(G188));
  INV_X1    g140(.A(G53), .ZN(new_n566));
  OAI21_X1  g141(.A(KEYINPUT9), .B1(new_n519), .B2(new_n566), .ZN(new_n567));
  INV_X1    g142(.A(KEYINPUT9), .ZN(new_n568));
  NAND4_X1  g143(.A1(new_n518), .A2(new_n568), .A3(G53), .A4(G543), .ZN(new_n569));
  NAND2_X1  g144(.A1(new_n567), .A2(new_n569), .ZN(new_n570));
  NAND3_X1  g145(.A1(new_n521), .A2(G91), .A3(new_n523), .ZN(new_n571));
  NAND2_X1  g146(.A1(G78), .A2(G543), .ZN(new_n572));
  XNOR2_X1  g147(.A(KEYINPUT74), .B(G65), .ZN(new_n573));
  OAI21_X1  g148(.A(new_n572), .B1(new_n553), .B2(new_n573), .ZN(new_n574));
  NAND2_X1  g149(.A1(new_n574), .A2(G651), .ZN(new_n575));
  NAND3_X1  g150(.A1(new_n570), .A2(new_n571), .A3(new_n575), .ZN(G299));
  INV_X1    g151(.A(G168), .ZN(G286));
  INV_X1    g152(.A(new_n524), .ZN(new_n578));
  NAND2_X1  g153(.A1(new_n578), .A2(G87), .ZN(new_n579));
  OAI21_X1  g154(.A(G651), .B1(new_n513), .B2(G74), .ZN(new_n580));
  XOR2_X1   g155(.A(new_n580), .B(KEYINPUT75), .Z(new_n581));
  NAND2_X1  g156(.A1(new_n528), .A2(G49), .ZN(new_n582));
  NAND3_X1  g157(.A1(new_n579), .A2(new_n581), .A3(new_n582), .ZN(G288));
  NAND2_X1  g158(.A1(new_n578), .A2(G86), .ZN(new_n584));
  NAND2_X1  g159(.A1(G73), .A2(G543), .ZN(new_n585));
  XNOR2_X1  g160(.A(new_n585), .B(KEYINPUT76), .ZN(new_n586));
  INV_X1    g161(.A(G61), .ZN(new_n587));
  OAI21_X1  g162(.A(new_n586), .B1(new_n553), .B2(new_n587), .ZN(new_n588));
  AOI22_X1  g163(.A1(new_n588), .A2(G651), .B1(G48), .B2(new_n528), .ZN(new_n589));
  NAND2_X1  g164(.A1(new_n584), .A2(new_n589), .ZN(G305));
  XOR2_X1   g165(.A(KEYINPUT77), .B(G85), .Z(new_n591));
  NAND2_X1  g166(.A1(new_n578), .A2(new_n591), .ZN(new_n592));
  NAND2_X1  g167(.A1(G72), .A2(G543), .ZN(new_n593));
  INV_X1    g168(.A(G60), .ZN(new_n594));
  OAI21_X1  g169(.A(new_n593), .B1(new_n553), .B2(new_n594), .ZN(new_n595));
  AOI22_X1  g170(.A1(new_n595), .A2(G651), .B1(new_n528), .B2(G47), .ZN(new_n596));
  NAND2_X1  g171(.A1(new_n592), .A2(new_n596), .ZN(new_n597));
  NAND2_X1  g172(.A1(new_n597), .A2(KEYINPUT78), .ZN(new_n598));
  INV_X1    g173(.A(KEYINPUT78), .ZN(new_n599));
  NAND3_X1  g174(.A1(new_n592), .A2(new_n599), .A3(new_n596), .ZN(new_n600));
  NAND2_X1  g175(.A1(new_n598), .A2(new_n600), .ZN(G290));
  INV_X1    g176(.A(KEYINPUT10), .ZN(new_n602));
  INV_X1    g177(.A(G92), .ZN(new_n603));
  OAI21_X1  g178(.A(new_n602), .B1(new_n524), .B2(new_n603), .ZN(new_n604));
  NAND4_X1  g179(.A1(new_n521), .A2(KEYINPUT10), .A3(G92), .A4(new_n523), .ZN(new_n605));
  NAND2_X1  g180(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  NAND2_X1  g181(.A1(G79), .A2(G543), .ZN(new_n607));
  XNOR2_X1  g182(.A(KEYINPUT79), .B(G66), .ZN(new_n608));
  OAI21_X1  g183(.A(new_n607), .B1(new_n553), .B2(new_n608), .ZN(new_n609));
  AOI22_X1  g184(.A1(new_n609), .A2(G651), .B1(new_n528), .B2(G54), .ZN(new_n610));
  NAND2_X1  g185(.A1(new_n606), .A2(new_n610), .ZN(new_n611));
  INV_X1    g186(.A(G868), .ZN(new_n612));
  NAND2_X1  g187(.A1(new_n611), .A2(new_n612), .ZN(new_n613));
  OAI21_X1  g188(.A(new_n613), .B1(G171), .B2(new_n612), .ZN(G321));
  XOR2_X1   g189(.A(G321), .B(KEYINPUT80), .Z(G284));
  NAND2_X1  g190(.A1(G299), .A2(new_n612), .ZN(new_n616));
  OAI21_X1  g191(.A(new_n616), .B1(G168), .B2(new_n612), .ZN(G297));
  OAI21_X1  g192(.A(new_n616), .B1(G168), .B2(new_n612), .ZN(G280));
  INV_X1    g193(.A(new_n611), .ZN(new_n619));
  XNOR2_X1  g194(.A(KEYINPUT81), .B(G559), .ZN(new_n620));
  OAI21_X1  g195(.A(new_n619), .B1(G860), .B2(new_n620), .ZN(G148));
  NAND2_X1  g196(.A1(new_n558), .A2(new_n612), .ZN(new_n622));
  AND2_X1   g197(.A1(new_n619), .A2(new_n620), .ZN(new_n623));
  OAI21_X1  g198(.A(new_n622), .B1(new_n623), .B2(new_n612), .ZN(G323));
  XNOR2_X1  g199(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g200(.A1(new_n467), .A2(new_n465), .ZN(new_n626));
  XOR2_X1   g201(.A(KEYINPUT82), .B(KEYINPUT12), .Z(new_n627));
  XNOR2_X1  g202(.A(new_n626), .B(new_n627), .ZN(new_n628));
  XNOR2_X1  g203(.A(new_n628), .B(KEYINPUT13), .ZN(new_n629));
  INV_X1    g204(.A(G2100), .ZN(new_n630));
  OR2_X1    g205(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  NAND2_X1  g206(.A1(new_n629), .A2(new_n630), .ZN(new_n632));
  AOI22_X1  g207(.A1(G123), .A2(new_n484), .B1(new_n482), .B2(G135), .ZN(new_n633));
  OAI21_X1  g208(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n634));
  INV_X1    g209(.A(KEYINPUT83), .ZN(new_n635));
  INV_X1    g210(.A(G111), .ZN(new_n636));
  AOI22_X1  g211(.A1(new_n634), .A2(new_n635), .B1(new_n636), .B2(G2105), .ZN(new_n637));
  OAI21_X1  g212(.A(new_n637), .B1(new_n635), .B2(new_n634), .ZN(new_n638));
  NAND2_X1  g213(.A1(new_n633), .A2(new_n638), .ZN(new_n639));
  XOR2_X1   g214(.A(new_n639), .B(G2096), .Z(new_n640));
  NAND3_X1  g215(.A1(new_n631), .A2(new_n632), .A3(new_n640), .ZN(G156));
  XOR2_X1   g216(.A(KEYINPUT15), .B(G2435), .Z(new_n642));
  XNOR2_X1  g217(.A(new_n642), .B(G2438), .ZN(new_n643));
  XOR2_X1   g218(.A(G2427), .B(G2430), .Z(new_n644));
  OR2_X1    g219(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  XOR2_X1   g220(.A(KEYINPUT85), .B(KEYINPUT14), .Z(new_n646));
  NAND2_X1  g221(.A1(new_n643), .A2(new_n644), .ZN(new_n647));
  NAND3_X1  g222(.A1(new_n645), .A2(new_n646), .A3(new_n647), .ZN(new_n648));
  XOR2_X1   g223(.A(G1341), .B(G1348), .Z(new_n649));
  XNOR2_X1  g224(.A(KEYINPUT84), .B(KEYINPUT16), .ZN(new_n650));
  XNOR2_X1  g225(.A(new_n649), .B(new_n650), .ZN(new_n651));
  XNOR2_X1  g226(.A(new_n648), .B(new_n651), .ZN(new_n652));
  INV_X1    g227(.A(new_n652), .ZN(new_n653));
  XOR2_X1   g228(.A(G2443), .B(G2446), .Z(new_n654));
  XNOR2_X1  g229(.A(G2451), .B(G2454), .ZN(new_n655));
  XNOR2_X1  g230(.A(new_n654), .B(new_n655), .ZN(new_n656));
  INV_X1    g231(.A(new_n656), .ZN(new_n657));
  OAI21_X1  g232(.A(G14), .B1(new_n653), .B2(new_n657), .ZN(new_n658));
  AOI21_X1  g233(.A(new_n658), .B1(new_n657), .B2(new_n653), .ZN(G401));
  XOR2_X1   g234(.A(G2084), .B(G2090), .Z(new_n660));
  INV_X1    g235(.A(new_n660), .ZN(new_n661));
  XNOR2_X1  g236(.A(G2072), .B(G2078), .ZN(new_n662));
  XNOR2_X1  g237(.A(G2067), .B(G2678), .ZN(new_n663));
  OAI21_X1  g238(.A(new_n661), .B1(new_n662), .B2(new_n663), .ZN(new_n664));
  INV_X1    g239(.A(new_n664), .ZN(new_n665));
  INV_X1    g240(.A(KEYINPUT86), .ZN(new_n666));
  XNOR2_X1  g241(.A(new_n662), .B(KEYINPUT17), .ZN(new_n667));
  AOI22_X1  g242(.A1(new_n665), .A2(new_n666), .B1(new_n663), .B2(new_n667), .ZN(new_n668));
  OAI21_X1  g243(.A(new_n668), .B1(new_n666), .B2(new_n665), .ZN(new_n669));
  XOR2_X1   g244(.A(new_n669), .B(KEYINPUT87), .Z(new_n670));
  NOR3_X1   g245(.A1(new_n667), .A2(new_n663), .A3(new_n661), .ZN(new_n671));
  XNOR2_X1  g246(.A(new_n671), .B(KEYINPUT88), .ZN(new_n672));
  NAND3_X1  g247(.A1(new_n660), .A2(new_n663), .A3(new_n662), .ZN(new_n673));
  XOR2_X1   g248(.A(new_n673), .B(KEYINPUT18), .Z(new_n674));
  NAND3_X1  g249(.A1(new_n670), .A2(new_n672), .A3(new_n674), .ZN(new_n675));
  XOR2_X1   g250(.A(G2096), .B(G2100), .Z(new_n676));
  XNOR2_X1  g251(.A(new_n675), .B(new_n676), .ZN(G227));
  XOR2_X1   g252(.A(G1961), .B(G1966), .Z(new_n678));
  XNOR2_X1  g253(.A(new_n678), .B(KEYINPUT90), .ZN(new_n679));
  XNOR2_X1  g254(.A(G1956), .B(G2474), .ZN(new_n680));
  XNOR2_X1  g255(.A(new_n680), .B(KEYINPUT89), .ZN(new_n681));
  NAND2_X1  g256(.A1(new_n679), .A2(new_n681), .ZN(new_n682));
  XNOR2_X1  g257(.A(G1971), .B(G1976), .ZN(new_n683));
  XNOR2_X1  g258(.A(new_n683), .B(KEYINPUT19), .ZN(new_n684));
  NOR2_X1   g259(.A1(new_n682), .A2(new_n684), .ZN(new_n685));
  XOR2_X1   g260(.A(new_n685), .B(KEYINPUT20), .Z(new_n686));
  OR2_X1    g261(.A1(new_n679), .A2(new_n681), .ZN(new_n687));
  NAND3_X1  g262(.A1(new_n687), .A2(new_n684), .A3(new_n682), .ZN(new_n688));
  OAI211_X1 g263(.A(new_n686), .B(new_n688), .C1(new_n684), .C2(new_n687), .ZN(new_n689));
  XOR2_X1   g264(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n690));
  XNOR2_X1  g265(.A(new_n690), .B(KEYINPUT91), .ZN(new_n691));
  XNOR2_X1  g266(.A(new_n689), .B(new_n691), .ZN(new_n692));
  XNOR2_X1  g267(.A(G1981), .B(G1986), .ZN(new_n693));
  XNOR2_X1  g268(.A(new_n693), .B(KEYINPUT92), .ZN(new_n694));
  XNOR2_X1  g269(.A(new_n692), .B(new_n694), .ZN(new_n695));
  XNOR2_X1  g270(.A(G1991), .B(G1996), .ZN(new_n696));
  XNOR2_X1  g271(.A(new_n695), .B(new_n696), .ZN(G229));
  NAND2_X1  g272(.A1(new_n482), .A2(G139), .ZN(new_n698));
  XOR2_X1   g273(.A(new_n698), .B(KEYINPUT96), .Z(new_n699));
  NAND3_X1  g274(.A1(new_n464), .A2(G103), .A3(G2104), .ZN(new_n700));
  XOR2_X1   g275(.A(new_n700), .B(KEYINPUT25), .Z(new_n701));
  AOI22_X1  g276(.A1(new_n467), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n702));
  OAI211_X1 g277(.A(new_n699), .B(new_n701), .C1(new_n464), .C2(new_n702), .ZN(new_n703));
  MUX2_X1   g278(.A(G33), .B(new_n703), .S(G29), .Z(new_n704));
  XNOR2_X1  g279(.A(new_n704), .B(new_n442), .ZN(new_n705));
  NAND3_X1  g280(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n706));
  XOR2_X1   g281(.A(new_n706), .B(KEYINPUT26), .Z(new_n707));
  INV_X1    g282(.A(G129), .ZN(new_n708));
  OAI21_X1  g283(.A(new_n707), .B1(new_n501), .B2(new_n708), .ZN(new_n709));
  AOI22_X1  g284(.A1(new_n482), .A2(G141), .B1(G105), .B2(new_n465), .ZN(new_n710));
  INV_X1    g285(.A(new_n710), .ZN(new_n711));
  NOR2_X1   g286(.A1(new_n709), .A2(new_n711), .ZN(new_n712));
  INV_X1    g287(.A(G29), .ZN(new_n713));
  NOR2_X1   g288(.A1(new_n712), .A2(new_n713), .ZN(new_n714));
  AOI21_X1  g289(.A(new_n714), .B1(new_n713), .B2(G32), .ZN(new_n715));
  XOR2_X1   g290(.A(KEYINPUT27), .B(G1996), .Z(new_n716));
  XNOR2_X1  g291(.A(new_n716), .B(KEYINPUT97), .ZN(new_n717));
  INV_X1    g292(.A(KEYINPUT24), .ZN(new_n718));
  OAI21_X1  g293(.A(new_n713), .B1(new_n718), .B2(G34), .ZN(new_n719));
  AOI21_X1  g294(.A(new_n719), .B1(new_n718), .B2(G34), .ZN(new_n720));
  AOI21_X1  g295(.A(new_n720), .B1(G160), .B2(G29), .ZN(new_n721));
  AOI22_X1  g296(.A1(new_n715), .A2(new_n717), .B1(G2084), .B2(new_n721), .ZN(new_n722));
  NAND2_X1  g297(.A1(new_n705), .A2(new_n722), .ZN(new_n723));
  XOR2_X1   g298(.A(new_n723), .B(KEYINPUT98), .Z(new_n724));
  NOR2_X1   g299(.A1(G5), .A2(G16), .ZN(new_n725));
  XOR2_X1   g300(.A(new_n725), .B(KEYINPUT101), .Z(new_n726));
  INV_X1    g301(.A(G16), .ZN(new_n727));
  OAI21_X1  g302(.A(new_n726), .B1(G301), .B2(new_n727), .ZN(new_n728));
  XNOR2_X1  g303(.A(new_n728), .B(G1961), .ZN(new_n729));
  NAND2_X1  g304(.A1(new_n713), .A2(G27), .ZN(new_n730));
  OAI21_X1  g305(.A(new_n730), .B1(G164), .B2(new_n713), .ZN(new_n731));
  XOR2_X1   g306(.A(new_n731), .B(KEYINPUT102), .Z(new_n732));
  OAI21_X1  g307(.A(new_n729), .B1(new_n732), .B2(G2078), .ZN(new_n733));
  NOR2_X1   g308(.A1(G16), .A2(G19), .ZN(new_n734));
  AOI21_X1  g309(.A(new_n734), .B1(new_n559), .B2(G16), .ZN(new_n735));
  XOR2_X1   g310(.A(new_n735), .B(G1341), .Z(new_n736));
  INV_X1    g311(.A(new_n736), .ZN(new_n737));
  NOR2_X1   g312(.A1(new_n721), .A2(G2084), .ZN(new_n738));
  NAND2_X1  g313(.A1(new_n713), .A2(G35), .ZN(new_n739));
  OAI21_X1  g314(.A(new_n739), .B1(G162), .B2(new_n713), .ZN(new_n740));
  XNOR2_X1  g315(.A(KEYINPUT29), .B(G2090), .ZN(new_n741));
  XNOR2_X1  g316(.A(new_n740), .B(new_n741), .ZN(new_n742));
  XNOR2_X1  g317(.A(KEYINPUT31), .B(G11), .ZN(new_n743));
  XOR2_X1   g318(.A(KEYINPUT99), .B(G28), .Z(new_n744));
  AOI21_X1  g319(.A(G29), .B1(new_n744), .B2(KEYINPUT30), .ZN(new_n745));
  INV_X1    g320(.A(new_n745), .ZN(new_n746));
  OAI22_X1  g321(.A1(new_n746), .A2(KEYINPUT100), .B1(KEYINPUT30), .B2(new_n744), .ZN(new_n747));
  AND2_X1   g322(.A1(new_n746), .A2(KEYINPUT100), .ZN(new_n748));
  OAI221_X1 g323(.A(new_n743), .B1(new_n713), .B2(new_n639), .C1(new_n747), .C2(new_n748), .ZN(new_n749));
  INV_X1    g324(.A(new_n749), .ZN(new_n750));
  OAI21_X1  g325(.A(new_n750), .B1(new_n715), .B2(new_n717), .ZN(new_n751));
  NOR4_X1   g326(.A1(new_n737), .A2(new_n738), .A3(new_n742), .A4(new_n751), .ZN(new_n752));
  NAND2_X1  g327(.A1(new_n727), .A2(G21), .ZN(new_n753));
  OAI21_X1  g328(.A(new_n753), .B1(G168), .B2(new_n727), .ZN(new_n754));
  XNOR2_X1  g329(.A(new_n754), .B(G1966), .ZN(new_n755));
  NAND2_X1  g330(.A1(new_n727), .A2(G20), .ZN(new_n756));
  XOR2_X1   g331(.A(new_n756), .B(KEYINPUT23), .Z(new_n757));
  AOI21_X1  g332(.A(new_n757), .B1(G299), .B2(G16), .ZN(new_n758));
  INV_X1    g333(.A(G1956), .ZN(new_n759));
  XNOR2_X1  g334(.A(new_n758), .B(new_n759), .ZN(new_n760));
  NAND2_X1  g335(.A1(new_n713), .A2(G26), .ZN(new_n761));
  XNOR2_X1  g336(.A(new_n761), .B(KEYINPUT28), .ZN(new_n762));
  NAND2_X1  g337(.A1(new_n482), .A2(G140), .ZN(new_n763));
  NAND2_X1  g338(.A1(new_n484), .A2(G128), .ZN(new_n764));
  OR2_X1    g339(.A1(G104), .A2(G2105), .ZN(new_n765));
  OAI211_X1 g340(.A(new_n765), .B(G2104), .C1(G116), .C2(new_n464), .ZN(new_n766));
  NAND3_X1  g341(.A1(new_n763), .A2(new_n764), .A3(new_n766), .ZN(new_n767));
  INV_X1    g342(.A(new_n767), .ZN(new_n768));
  OAI21_X1  g343(.A(new_n762), .B1(new_n768), .B2(new_n713), .ZN(new_n769));
  XNOR2_X1  g344(.A(new_n769), .B(G2067), .ZN(new_n770));
  NOR3_X1   g345(.A1(new_n755), .A2(new_n760), .A3(new_n770), .ZN(new_n771));
  NOR2_X1   g346(.A1(G4), .A2(G16), .ZN(new_n772));
  AOI21_X1  g347(.A(new_n772), .B1(new_n619), .B2(G16), .ZN(new_n773));
  INV_X1    g348(.A(G1348), .ZN(new_n774));
  XNOR2_X1  g349(.A(new_n773), .B(new_n774), .ZN(new_n775));
  NAND2_X1  g350(.A1(new_n732), .A2(G2078), .ZN(new_n776));
  NAND4_X1  g351(.A1(new_n752), .A2(new_n771), .A3(new_n775), .A4(new_n776), .ZN(new_n777));
  NOR3_X1   g352(.A1(new_n724), .A2(new_n733), .A3(new_n777), .ZN(new_n778));
  INV_X1    g353(.A(new_n778), .ZN(new_n779));
  INV_X1    g354(.A(KEYINPUT36), .ZN(new_n780));
  NAND2_X1  g355(.A1(new_n727), .A2(G23), .ZN(new_n781));
  INV_X1    g356(.A(G288), .ZN(new_n782));
  OAI21_X1  g357(.A(new_n781), .B1(new_n782), .B2(new_n727), .ZN(new_n783));
  XNOR2_X1  g358(.A(KEYINPUT33), .B(G1976), .ZN(new_n784));
  XNOR2_X1  g359(.A(new_n783), .B(new_n784), .ZN(new_n785));
  INV_X1    g360(.A(KEYINPUT94), .ZN(new_n786));
  OR2_X1    g361(.A1(new_n785), .A2(new_n786), .ZN(new_n787));
  NAND2_X1  g362(.A1(new_n785), .A2(new_n786), .ZN(new_n788));
  NOR2_X1   g363(.A1(G6), .A2(G16), .ZN(new_n789));
  INV_X1    g364(.A(G305), .ZN(new_n790));
  AOI21_X1  g365(.A(new_n789), .B1(new_n790), .B2(G16), .ZN(new_n791));
  XOR2_X1   g366(.A(KEYINPUT32), .B(G1981), .Z(new_n792));
  XNOR2_X1  g367(.A(new_n791), .B(new_n792), .ZN(new_n793));
  NAND2_X1  g368(.A1(new_n727), .A2(G22), .ZN(new_n794));
  OAI21_X1  g369(.A(new_n794), .B1(G166), .B2(new_n727), .ZN(new_n795));
  INV_X1    g370(.A(G1971), .ZN(new_n796));
  XNOR2_X1  g371(.A(new_n795), .B(new_n796), .ZN(new_n797));
  AND2_X1   g372(.A1(new_n793), .A2(new_n797), .ZN(new_n798));
  NAND3_X1  g373(.A1(new_n787), .A2(new_n788), .A3(new_n798), .ZN(new_n799));
  NAND2_X1  g374(.A1(new_n799), .A2(KEYINPUT34), .ZN(new_n800));
  INV_X1    g375(.A(KEYINPUT95), .ZN(new_n801));
  NAND2_X1  g376(.A1(new_n800), .A2(new_n801), .ZN(new_n802));
  NAND3_X1  g377(.A1(new_n799), .A2(KEYINPUT95), .A3(KEYINPUT34), .ZN(new_n803));
  NAND2_X1  g378(.A1(new_n802), .A2(new_n803), .ZN(new_n804));
  NOR2_X1   g379(.A1(new_n799), .A2(KEYINPUT34), .ZN(new_n805));
  MUX2_X1   g380(.A(G24), .B(G290), .S(G16), .Z(new_n806));
  NOR2_X1   g381(.A1(new_n806), .A2(G1986), .ZN(new_n807));
  AND2_X1   g382(.A1(new_n806), .A2(G1986), .ZN(new_n808));
  NAND2_X1  g383(.A1(new_n482), .A2(G131), .ZN(new_n809));
  NAND2_X1  g384(.A1(new_n484), .A2(G119), .ZN(new_n810));
  NOR2_X1   g385(.A1(new_n464), .A2(G107), .ZN(new_n811));
  OAI21_X1  g386(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n812));
  OAI211_X1 g387(.A(new_n809), .B(new_n810), .C1(new_n811), .C2(new_n812), .ZN(new_n813));
  MUX2_X1   g388(.A(G25), .B(new_n813), .S(G29), .Z(new_n814));
  XNOR2_X1  g389(.A(KEYINPUT35), .B(G1991), .ZN(new_n815));
  XNOR2_X1  g390(.A(new_n815), .B(KEYINPUT93), .ZN(new_n816));
  XNOR2_X1  g391(.A(new_n814), .B(new_n816), .ZN(new_n817));
  OR2_X1    g392(.A1(new_n808), .A2(new_n817), .ZN(new_n818));
  NOR3_X1   g393(.A1(new_n805), .A2(new_n807), .A3(new_n818), .ZN(new_n819));
  AOI21_X1  g394(.A(new_n780), .B1(new_n804), .B2(new_n819), .ZN(new_n820));
  INV_X1    g395(.A(new_n820), .ZN(new_n821));
  NAND3_X1  g396(.A1(new_n804), .A2(new_n819), .A3(new_n780), .ZN(new_n822));
  AOI21_X1  g397(.A(new_n779), .B1(new_n821), .B2(new_n822), .ZN(G311));
  INV_X1    g398(.A(new_n822), .ZN(new_n824));
  OAI21_X1  g399(.A(new_n778), .B1(new_n824), .B2(new_n820), .ZN(G150));
  NAND2_X1  g400(.A1(G80), .A2(G543), .ZN(new_n826));
  INV_X1    g401(.A(G67), .ZN(new_n827));
  OAI21_X1  g402(.A(new_n826), .B1(new_n553), .B2(new_n827), .ZN(new_n828));
  AOI22_X1  g403(.A1(new_n828), .A2(G651), .B1(new_n528), .B2(G55), .ZN(new_n829));
  INV_X1    g404(.A(KEYINPUT103), .ZN(new_n830));
  NAND3_X1  g405(.A1(new_n521), .A2(G93), .A3(new_n523), .ZN(new_n831));
  AND3_X1   g406(.A1(new_n829), .A2(new_n830), .A3(new_n831), .ZN(new_n832));
  AOI21_X1  g407(.A(new_n830), .B1(new_n829), .B2(new_n831), .ZN(new_n833));
  NOR3_X1   g408(.A1(new_n832), .A2(new_n833), .A3(new_n558), .ZN(new_n834));
  NAND2_X1  g409(.A1(new_n829), .A2(new_n831), .ZN(new_n835));
  AND3_X1   g410(.A1(new_n558), .A2(new_n835), .A3(KEYINPUT103), .ZN(new_n836));
  NOR2_X1   g411(.A1(new_n834), .A2(new_n836), .ZN(new_n837));
  XNOR2_X1  g412(.A(new_n837), .B(KEYINPUT38), .ZN(new_n838));
  NAND2_X1  g413(.A1(new_n619), .A2(G559), .ZN(new_n839));
  XNOR2_X1  g414(.A(new_n838), .B(new_n839), .ZN(new_n840));
  AND2_X1   g415(.A1(new_n840), .A2(KEYINPUT39), .ZN(new_n841));
  NOR2_X1   g416(.A1(new_n840), .A2(KEYINPUT39), .ZN(new_n842));
  NOR3_X1   g417(.A1(new_n841), .A2(new_n842), .A3(G860), .ZN(new_n843));
  NAND2_X1  g418(.A1(new_n835), .A2(G860), .ZN(new_n844));
  XNOR2_X1  g419(.A(new_n844), .B(KEYINPUT37), .ZN(new_n845));
  OR2_X1    g420(.A1(new_n843), .A2(new_n845), .ZN(G145));
  NAND2_X1  g421(.A1(new_n507), .A2(new_n509), .ZN(new_n847));
  XNOR2_X1  g422(.A(new_n847), .B(new_n767), .ZN(new_n848));
  XNOR2_X1  g423(.A(new_n703), .B(new_n848), .ZN(new_n849));
  XNOR2_X1  g424(.A(new_n849), .B(new_n712), .ZN(new_n850));
  XNOR2_X1  g425(.A(new_n628), .B(new_n813), .ZN(new_n851));
  NAND2_X1  g426(.A1(new_n482), .A2(G142), .ZN(new_n852));
  NAND2_X1  g427(.A1(new_n484), .A2(G130), .ZN(new_n853));
  OR2_X1    g428(.A1(G106), .A2(G2105), .ZN(new_n854));
  OAI211_X1 g429(.A(new_n854), .B(G2104), .C1(G118), .C2(new_n464), .ZN(new_n855));
  NAND3_X1  g430(.A1(new_n852), .A2(new_n853), .A3(new_n855), .ZN(new_n856));
  XNOR2_X1  g431(.A(new_n851), .B(new_n856), .ZN(new_n857));
  NAND2_X1  g432(.A1(new_n857), .A2(KEYINPUT104), .ZN(new_n858));
  OR2_X1    g433(.A1(new_n850), .A2(new_n858), .ZN(new_n859));
  NAND2_X1  g434(.A1(new_n850), .A2(new_n858), .ZN(new_n860));
  XNOR2_X1  g435(.A(G160), .B(new_n488), .ZN(new_n861));
  XNOR2_X1  g436(.A(new_n861), .B(new_n639), .ZN(new_n862));
  NAND3_X1  g437(.A1(new_n859), .A2(new_n860), .A3(new_n862), .ZN(new_n863));
  AOI21_X1  g438(.A(new_n862), .B1(new_n850), .B2(new_n857), .ZN(new_n864));
  OAI21_X1  g439(.A(new_n864), .B1(new_n850), .B2(new_n857), .ZN(new_n865));
  INV_X1    g440(.A(G37), .ZN(new_n866));
  NAND3_X1  g441(.A1(new_n863), .A2(new_n865), .A3(new_n866), .ZN(new_n867));
  XNOR2_X1  g442(.A(new_n867), .B(KEYINPUT40), .ZN(G395));
  NAND2_X1  g443(.A1(new_n835), .A2(new_n612), .ZN(new_n869));
  AOI21_X1  g444(.A(G303), .B1(new_n598), .B2(new_n600), .ZN(new_n870));
  INV_X1    g445(.A(new_n870), .ZN(new_n871));
  NAND3_X1  g446(.A1(new_n598), .A2(G303), .A3(new_n600), .ZN(new_n872));
  NAND2_X1  g447(.A1(new_n790), .A2(G288), .ZN(new_n873));
  NAND2_X1  g448(.A1(new_n782), .A2(G305), .ZN(new_n874));
  NAND4_X1  g449(.A1(new_n871), .A2(new_n872), .A3(new_n873), .A4(new_n874), .ZN(new_n875));
  NAND2_X1  g450(.A1(new_n874), .A2(new_n873), .ZN(new_n876));
  INV_X1    g451(.A(new_n872), .ZN(new_n877));
  OAI21_X1  g452(.A(new_n876), .B1(new_n877), .B2(new_n870), .ZN(new_n878));
  NAND2_X1  g453(.A1(new_n875), .A2(new_n878), .ZN(new_n879));
  INV_X1    g454(.A(KEYINPUT105), .ZN(new_n880));
  OR2_X1    g455(.A1(new_n880), .A2(KEYINPUT42), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n880), .A2(KEYINPUT42), .ZN(new_n882));
  AOI21_X1  g457(.A(new_n879), .B1(new_n881), .B2(new_n882), .ZN(new_n883));
  INV_X1    g458(.A(KEYINPUT106), .ZN(new_n884));
  AOI22_X1  g459(.A1(new_n883), .A2(new_n884), .B1(KEYINPUT42), .B2(new_n879), .ZN(new_n885));
  OAI21_X1  g460(.A(new_n885), .B1(new_n884), .B2(new_n883), .ZN(new_n886));
  OR2_X1    g461(.A1(new_n834), .A2(new_n836), .ZN(new_n887));
  XNOR2_X1  g462(.A(new_n623), .B(new_n887), .ZN(new_n888));
  INV_X1    g463(.A(G299), .ZN(new_n889));
  AND3_X1   g464(.A1(new_n606), .A2(new_n889), .A3(new_n610), .ZN(new_n890));
  AOI21_X1  g465(.A(new_n889), .B1(new_n606), .B2(new_n610), .ZN(new_n891));
  NOR2_X1   g466(.A1(new_n890), .A2(new_n891), .ZN(new_n892));
  NOR2_X1   g467(.A1(new_n888), .A2(new_n892), .ZN(new_n893));
  INV_X1    g468(.A(KEYINPUT41), .ZN(new_n894));
  OAI21_X1  g469(.A(new_n894), .B1(new_n890), .B2(new_n891), .ZN(new_n895));
  NAND2_X1  g470(.A1(new_n611), .A2(G299), .ZN(new_n896));
  NAND3_X1  g471(.A1(new_n606), .A2(new_n889), .A3(new_n610), .ZN(new_n897));
  NAND3_X1  g472(.A1(new_n896), .A2(KEYINPUT41), .A3(new_n897), .ZN(new_n898));
  NAND2_X1  g473(.A1(new_n895), .A2(new_n898), .ZN(new_n899));
  AOI21_X1  g474(.A(new_n893), .B1(new_n888), .B2(new_n899), .ZN(new_n900));
  XNOR2_X1  g475(.A(new_n886), .B(new_n900), .ZN(new_n901));
  OAI21_X1  g476(.A(new_n869), .B1(new_n901), .B2(new_n612), .ZN(G295));
  OAI21_X1  g477(.A(new_n869), .B1(new_n901), .B2(new_n612), .ZN(G331));
  INV_X1    g478(.A(KEYINPUT107), .ZN(new_n904));
  NAND4_X1  g479(.A1(new_n535), .A2(new_n538), .A3(new_n904), .A4(new_n536), .ZN(new_n905));
  AND3_X1   g480(.A1(new_n541), .A2(KEYINPUT72), .A3(new_n542), .ZN(new_n906));
  AOI21_X1  g481(.A(KEYINPUT72), .B1(new_n541), .B2(new_n542), .ZN(new_n907));
  OAI211_X1 g482(.A(new_n549), .B(new_n905), .C1(new_n906), .C2(new_n907), .ZN(new_n908));
  OAI21_X1  g483(.A(KEYINPUT107), .B1(new_n537), .B2(new_n539), .ZN(new_n909));
  INV_X1    g484(.A(new_n909), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n908), .A2(new_n910), .ZN(new_n911));
  NAND4_X1  g486(.A1(new_n547), .A2(new_n909), .A3(new_n549), .A4(new_n905), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n911), .A2(new_n912), .ZN(new_n913));
  NAND2_X1  g488(.A1(new_n913), .A2(new_n887), .ZN(new_n914));
  NAND3_X1  g489(.A1(new_n837), .A2(new_n911), .A3(new_n912), .ZN(new_n915));
  NAND2_X1  g490(.A1(new_n914), .A2(new_n915), .ZN(new_n916));
  INV_X1    g491(.A(new_n899), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n916), .A2(new_n917), .ZN(new_n918));
  NAND3_X1  g493(.A1(new_n914), .A2(new_n892), .A3(new_n915), .ZN(new_n919));
  AOI21_X1  g494(.A(new_n879), .B1(new_n918), .B2(new_n919), .ZN(new_n920));
  OAI21_X1  g495(.A(KEYINPUT108), .B1(new_n920), .B2(G37), .ZN(new_n921));
  AND2_X1   g496(.A1(new_n875), .A2(new_n878), .ZN(new_n922));
  AND3_X1   g497(.A1(new_n914), .A2(new_n892), .A3(new_n915), .ZN(new_n923));
  AOI21_X1  g498(.A(new_n899), .B1(new_n914), .B2(new_n915), .ZN(new_n924));
  OAI21_X1  g499(.A(new_n922), .B1(new_n923), .B2(new_n924), .ZN(new_n925));
  INV_X1    g500(.A(KEYINPUT108), .ZN(new_n926));
  NAND3_X1  g501(.A1(new_n925), .A2(new_n926), .A3(new_n866), .ZN(new_n927));
  NAND3_X1  g502(.A1(new_n918), .A2(new_n879), .A3(new_n919), .ZN(new_n928));
  NAND3_X1  g503(.A1(new_n921), .A2(new_n927), .A3(new_n928), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n929), .A2(KEYINPUT43), .ZN(new_n930));
  AOI21_X1  g505(.A(new_n923), .B1(new_n918), .B2(KEYINPUT109), .ZN(new_n931));
  INV_X1    g506(.A(KEYINPUT109), .ZN(new_n932));
  NAND2_X1  g507(.A1(new_n924), .A2(new_n932), .ZN(new_n933));
  AOI21_X1  g508(.A(new_n879), .B1(new_n931), .B2(new_n933), .ZN(new_n934));
  INV_X1    g509(.A(new_n934), .ZN(new_n935));
  INV_X1    g510(.A(KEYINPUT43), .ZN(new_n936));
  NAND2_X1  g511(.A1(new_n928), .A2(new_n866), .ZN(new_n937));
  INV_X1    g512(.A(new_n937), .ZN(new_n938));
  NAND3_X1  g513(.A1(new_n935), .A2(new_n936), .A3(new_n938), .ZN(new_n939));
  INV_X1    g514(.A(KEYINPUT44), .ZN(new_n940));
  AND3_X1   g515(.A1(new_n930), .A2(new_n939), .A3(new_n940), .ZN(new_n941));
  OAI21_X1  g516(.A(KEYINPUT43), .B1(new_n934), .B2(new_n937), .ZN(new_n942));
  INV_X1    g517(.A(KEYINPUT110), .ZN(new_n943));
  NAND2_X1  g518(.A1(new_n942), .A2(new_n943), .ZN(new_n944));
  OAI211_X1 g519(.A(KEYINPUT110), .B(KEYINPUT43), .C1(new_n934), .C2(new_n937), .ZN(new_n945));
  OAI211_X1 g520(.A(new_n944), .B(new_n945), .C1(KEYINPUT43), .C2(new_n929), .ZN(new_n946));
  AOI21_X1  g521(.A(new_n941), .B1(new_n946), .B2(KEYINPUT44), .ZN(G397));
  NAND2_X1  g522(.A1(G303), .A2(G8), .ZN(new_n948));
  XNOR2_X1  g523(.A(new_n948), .B(KEYINPUT55), .ZN(new_n949));
  AOI21_X1  g524(.A(G1384), .B1(new_n504), .B2(new_n510), .ZN(new_n950));
  OAI21_X1  g525(.A(KEYINPUT113), .B1(new_n950), .B2(KEYINPUT45), .ZN(new_n951));
  INV_X1    g526(.A(G1384), .ZN(new_n952));
  AND3_X1   g527(.A1(new_n507), .A2(new_n508), .A3(new_n509), .ZN(new_n953));
  AOI21_X1  g528(.A(new_n508), .B1(new_n507), .B2(new_n509), .ZN(new_n954));
  OAI21_X1  g529(.A(new_n952), .B1(new_n953), .B2(new_n954), .ZN(new_n955));
  INV_X1    g530(.A(KEYINPUT113), .ZN(new_n956));
  INV_X1    g531(.A(KEYINPUT45), .ZN(new_n957));
  NAND3_X1  g532(.A1(new_n955), .A2(new_n956), .A3(new_n957), .ZN(new_n958));
  NAND2_X1  g533(.A1(new_n478), .A2(G2105), .ZN(new_n959));
  INV_X1    g534(.A(new_n470), .ZN(new_n960));
  NAND3_X1  g535(.A1(new_n959), .A2(G40), .A3(new_n960), .ZN(new_n961));
  AOI21_X1  g536(.A(G1384), .B1(new_n507), .B2(new_n509), .ZN(new_n962));
  AOI21_X1  g537(.A(new_n961), .B1(KEYINPUT45), .B2(new_n962), .ZN(new_n963));
  NAND3_X1  g538(.A1(new_n951), .A2(new_n958), .A3(new_n963), .ZN(new_n964));
  AND2_X1   g539(.A1(new_n964), .A2(new_n796), .ZN(new_n965));
  NAND2_X1  g540(.A1(new_n847), .A2(new_n952), .ZN(new_n966));
  AOI21_X1  g541(.A(new_n961), .B1(KEYINPUT50), .B2(new_n966), .ZN(new_n967));
  INV_X1    g542(.A(KEYINPUT121), .ZN(new_n968));
  INV_X1    g543(.A(KEYINPUT50), .ZN(new_n969));
  AOI21_X1  g544(.A(new_n968), .B1(new_n950), .B2(new_n969), .ZN(new_n970));
  OAI211_X1 g545(.A(new_n969), .B(new_n952), .C1(new_n953), .C2(new_n954), .ZN(new_n971));
  NOR2_X1   g546(.A1(new_n971), .A2(KEYINPUT121), .ZN(new_n972));
  OAI21_X1  g547(.A(new_n967), .B1(new_n970), .B2(new_n972), .ZN(new_n973));
  INV_X1    g548(.A(KEYINPUT122), .ZN(new_n974));
  AOI21_X1  g549(.A(G2090), .B1(new_n973), .B2(new_n974), .ZN(new_n975));
  INV_X1    g550(.A(new_n961), .ZN(new_n976));
  OAI21_X1  g551(.A(new_n976), .B1(new_n969), .B2(new_n962), .ZN(new_n977));
  NAND2_X1  g552(.A1(new_n971), .A2(KEYINPUT121), .ZN(new_n978));
  NAND4_X1  g553(.A1(new_n511), .A2(new_n968), .A3(new_n969), .A4(new_n952), .ZN(new_n979));
  AOI21_X1  g554(.A(new_n977), .B1(new_n978), .B2(new_n979), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n980), .A2(KEYINPUT122), .ZN(new_n981));
  AOI21_X1  g556(.A(new_n965), .B1(new_n975), .B2(new_n981), .ZN(new_n982));
  XOR2_X1   g557(.A(KEYINPUT115), .B(G8), .Z(new_n983));
  OAI21_X1  g558(.A(new_n949), .B1(new_n982), .B2(new_n983), .ZN(new_n984));
  INV_X1    g559(.A(new_n949), .ZN(new_n985));
  OAI211_X1 g560(.A(KEYINPUT50), .B(new_n952), .C1(new_n953), .C2(new_n954), .ZN(new_n986));
  NAND2_X1  g561(.A1(new_n966), .A2(new_n969), .ZN(new_n987));
  NAND2_X1  g562(.A1(new_n986), .A2(new_n987), .ZN(new_n988));
  NAND2_X1  g563(.A1(new_n988), .A2(new_n976), .ZN(new_n989));
  OR2_X1    g564(.A1(new_n989), .A2(G2090), .ZN(new_n990));
  INV_X1    g565(.A(KEYINPUT114), .ZN(new_n991));
  OAI21_X1  g566(.A(new_n990), .B1(new_n965), .B2(new_n991), .ZN(new_n992));
  AND3_X1   g567(.A1(new_n964), .A2(new_n991), .A3(new_n796), .ZN(new_n993));
  OAI211_X1 g568(.A(G8), .B(new_n985), .C1(new_n992), .C2(new_n993), .ZN(new_n994));
  INV_X1    g569(.A(KEYINPUT49), .ZN(new_n995));
  INV_X1    g570(.A(G1981), .ZN(new_n996));
  NOR2_X1   g571(.A1(new_n790), .A2(new_n996), .ZN(new_n997));
  NAND2_X1  g572(.A1(new_n996), .A2(KEYINPUT118), .ZN(new_n998));
  OR2_X1    g573(.A1(new_n996), .A2(KEYINPUT118), .ZN(new_n999));
  AOI21_X1  g574(.A(G305), .B1(new_n998), .B2(new_n999), .ZN(new_n1000));
  OAI21_X1  g575(.A(new_n995), .B1(new_n997), .B2(new_n1000), .ZN(new_n1001));
  NAND2_X1  g576(.A1(new_n999), .A2(new_n998), .ZN(new_n1002));
  NAND2_X1  g577(.A1(new_n790), .A2(new_n1002), .ZN(new_n1003));
  OAI211_X1 g578(.A(new_n1003), .B(KEYINPUT49), .C1(new_n996), .C2(new_n790), .ZN(new_n1004));
  NAND2_X1  g579(.A1(new_n976), .A2(new_n962), .ZN(new_n1005));
  INV_X1    g580(.A(new_n983), .ZN(new_n1006));
  NAND2_X1  g581(.A1(new_n1005), .A2(new_n1006), .ZN(new_n1007));
  NOR2_X1   g582(.A1(new_n1007), .A2(KEYINPUT116), .ZN(new_n1008));
  INV_X1    g583(.A(KEYINPUT116), .ZN(new_n1009));
  AOI21_X1  g584(.A(new_n1009), .B1(new_n1005), .B2(new_n1006), .ZN(new_n1010));
  OAI211_X1 g585(.A(new_n1001), .B(new_n1004), .C1(new_n1008), .C2(new_n1010), .ZN(new_n1011));
  NAND4_X1  g586(.A1(new_n579), .A2(new_n581), .A3(G1976), .A4(new_n582), .ZN(new_n1012));
  INV_X1    g587(.A(KEYINPUT117), .ZN(new_n1013));
  XNOR2_X1  g588(.A(new_n1012), .B(new_n1013), .ZN(new_n1014));
  INV_X1    g589(.A(G1976), .ZN(new_n1015));
  AOI21_X1  g590(.A(KEYINPUT52), .B1(G288), .B2(new_n1015), .ZN(new_n1016));
  OAI211_X1 g591(.A(new_n1014), .B(new_n1016), .C1(new_n1008), .C2(new_n1010), .ZN(new_n1017));
  NAND2_X1  g592(.A1(new_n1011), .A2(new_n1017), .ZN(new_n1018));
  INV_X1    g593(.A(KEYINPUT52), .ZN(new_n1019));
  XNOR2_X1  g594(.A(new_n1007), .B(KEYINPUT116), .ZN(new_n1020));
  AOI21_X1  g595(.A(new_n1019), .B1(new_n1020), .B2(new_n1014), .ZN(new_n1021));
  NOR2_X1   g596(.A1(new_n1018), .A2(new_n1021), .ZN(new_n1022));
  AOI21_X1  g597(.A(KEYINPUT45), .B1(new_n847), .B2(new_n952), .ZN(new_n1023));
  NOR2_X1   g598(.A1(new_n1023), .A2(new_n961), .ZN(new_n1024));
  OAI211_X1 g599(.A(KEYINPUT45), .B(new_n952), .C1(new_n953), .C2(new_n954), .ZN(new_n1025));
  AOI21_X1  g600(.A(G1966), .B1(new_n1024), .B2(new_n1025), .ZN(new_n1026));
  INV_X1    g601(.A(G2084), .ZN(new_n1027));
  NAND3_X1  g602(.A1(G160), .A2(G40), .A3(new_n1027), .ZN(new_n1028));
  AOI21_X1  g603(.A(new_n1028), .B1(new_n986), .B2(new_n987), .ZN(new_n1029));
  OAI21_X1  g604(.A(new_n1006), .B1(new_n1026), .B2(new_n1029), .ZN(new_n1030));
  INV_X1    g605(.A(new_n1030), .ZN(new_n1031));
  NAND2_X1  g606(.A1(new_n1031), .A2(G168), .ZN(new_n1032));
  INV_X1    g607(.A(new_n1032), .ZN(new_n1033));
  NAND4_X1  g608(.A1(new_n984), .A2(new_n994), .A3(new_n1022), .A4(new_n1033), .ZN(new_n1034));
  INV_X1    g609(.A(KEYINPUT63), .ZN(new_n1035));
  NAND2_X1  g610(.A1(new_n1034), .A2(new_n1035), .ZN(new_n1036));
  INV_X1    g611(.A(KEYINPUT119), .ZN(new_n1037));
  OAI21_X1  g612(.A(new_n1037), .B1(new_n1018), .B2(new_n1021), .ZN(new_n1038));
  OAI21_X1  g613(.A(new_n1014), .B1(new_n1008), .B2(new_n1010), .ZN(new_n1039));
  NAND2_X1  g614(.A1(new_n1039), .A2(KEYINPUT52), .ZN(new_n1040));
  NAND4_X1  g615(.A1(new_n1040), .A2(KEYINPUT119), .A3(new_n1011), .A4(new_n1017), .ZN(new_n1041));
  NAND2_X1  g616(.A1(new_n1038), .A2(new_n1041), .ZN(new_n1042));
  OAI21_X1  g617(.A(G8), .B1(new_n992), .B2(new_n993), .ZN(new_n1043));
  NAND2_X1  g618(.A1(new_n1043), .A2(new_n949), .ZN(new_n1044));
  NOR2_X1   g619(.A1(new_n1032), .A2(new_n1035), .ZN(new_n1045));
  NAND4_X1  g620(.A1(new_n1042), .A2(new_n1044), .A3(new_n994), .A4(new_n1045), .ZN(new_n1046));
  NAND2_X1  g621(.A1(new_n1036), .A2(new_n1046), .ZN(new_n1047));
  AOI21_X1  g622(.A(new_n994), .B1(new_n1038), .B2(new_n1041), .ZN(new_n1048));
  AND2_X1   g623(.A1(new_n1001), .A2(new_n1004), .ZN(new_n1049));
  NOR2_X1   g624(.A1(G288), .A2(G1976), .ZN(new_n1050));
  XOR2_X1   g625(.A(new_n1050), .B(KEYINPUT120), .Z(new_n1051));
  OAI21_X1  g626(.A(new_n1003), .B1(new_n1049), .B2(new_n1051), .ZN(new_n1052));
  AOI21_X1  g627(.A(new_n1048), .B1(new_n1020), .B2(new_n1052), .ZN(new_n1053));
  XNOR2_X1  g628(.A(KEYINPUT56), .B(G2072), .ZN(new_n1054));
  NAND4_X1  g629(.A1(new_n951), .A2(new_n958), .A3(new_n963), .A4(new_n1054), .ZN(new_n1055));
  XOR2_X1   g630(.A(G299), .B(KEYINPUT57), .Z(new_n1056));
  OAI211_X1 g631(.A(new_n1055), .B(new_n1056), .C1(new_n980), .C2(G1956), .ZN(new_n1057));
  NAND2_X1  g632(.A1(new_n973), .A2(new_n759), .ZN(new_n1058));
  AOI21_X1  g633(.A(new_n1056), .B1(new_n1058), .B2(new_n1055), .ZN(new_n1059));
  INV_X1    g634(.A(G2067), .ZN(new_n1060));
  NOR2_X1   g635(.A1(new_n961), .A2(new_n966), .ZN(new_n1061));
  AOI22_X1  g636(.A1(new_n989), .A2(new_n774), .B1(new_n1060), .B2(new_n1061), .ZN(new_n1062));
  NOR2_X1   g637(.A1(new_n1062), .A2(new_n611), .ZN(new_n1063));
  OAI21_X1  g638(.A(new_n1057), .B1(new_n1059), .B2(new_n1063), .ZN(new_n1064));
  INV_X1    g639(.A(KEYINPUT61), .ZN(new_n1065));
  INV_X1    g640(.A(new_n1057), .ZN(new_n1066));
  OAI21_X1  g641(.A(new_n1065), .B1(new_n1059), .B2(new_n1066), .ZN(new_n1067));
  OAI21_X1  g642(.A(new_n1055), .B1(new_n980), .B2(G1956), .ZN(new_n1068));
  INV_X1    g643(.A(new_n1056), .ZN(new_n1069));
  NAND2_X1  g644(.A1(new_n1068), .A2(new_n1069), .ZN(new_n1070));
  NAND3_X1  g645(.A1(new_n1070), .A2(KEYINPUT61), .A3(new_n1057), .ZN(new_n1071));
  NAND2_X1  g646(.A1(new_n1067), .A2(new_n1071), .ZN(new_n1072));
  NAND2_X1  g647(.A1(new_n1061), .A2(new_n1060), .ZN(new_n1073));
  AOI21_X1  g648(.A(new_n961), .B1(new_n986), .B2(new_n987), .ZN(new_n1074));
  OAI211_X1 g649(.A(KEYINPUT60), .B(new_n1073), .C1(new_n1074), .C2(G1348), .ZN(new_n1075));
  XNOR2_X1  g650(.A(new_n1075), .B(new_n611), .ZN(new_n1076));
  NOR2_X1   g651(.A1(new_n1062), .A2(KEYINPUT60), .ZN(new_n1077));
  INV_X1    g652(.A(KEYINPUT59), .ZN(new_n1078));
  INV_X1    g653(.A(G1996), .ZN(new_n1079));
  NAND4_X1  g654(.A1(new_n951), .A2(new_n1079), .A3(new_n958), .A4(new_n963), .ZN(new_n1080));
  XOR2_X1   g655(.A(KEYINPUT58), .B(G1341), .Z(new_n1081));
  NAND2_X1  g656(.A1(new_n1005), .A2(new_n1081), .ZN(new_n1082));
  NAND2_X1  g657(.A1(new_n1080), .A2(new_n1082), .ZN(new_n1083));
  AOI21_X1  g658(.A(new_n1078), .B1(new_n1083), .B2(new_n559), .ZN(new_n1084));
  AOI211_X1 g659(.A(KEYINPUT59), .B(new_n558), .C1(new_n1080), .C2(new_n1082), .ZN(new_n1085));
  OAI22_X1  g660(.A1(new_n1076), .A2(new_n1077), .B1(new_n1084), .B2(new_n1085), .ZN(new_n1086));
  OAI21_X1  g661(.A(new_n1064), .B1(new_n1072), .B2(new_n1086), .ZN(new_n1087));
  NAND2_X1  g662(.A1(new_n1030), .A2(KEYINPUT123), .ZN(new_n1088));
  INV_X1    g663(.A(KEYINPUT123), .ZN(new_n1089));
  OAI211_X1 g664(.A(new_n1089), .B(new_n1006), .C1(new_n1026), .C2(new_n1029), .ZN(new_n1090));
  NOR2_X1   g665(.A1(G168), .A2(new_n983), .ZN(new_n1091));
  NOR2_X1   g666(.A1(new_n1091), .A2(KEYINPUT51), .ZN(new_n1092));
  NAND3_X1  g667(.A1(new_n1088), .A2(new_n1090), .A3(new_n1092), .ZN(new_n1093));
  INV_X1    g668(.A(G8), .ZN(new_n1094));
  NAND2_X1  g669(.A1(new_n1024), .A2(new_n1025), .ZN(new_n1095));
  INV_X1    g670(.A(G1966), .ZN(new_n1096));
  NAND2_X1  g671(.A1(new_n1095), .A2(new_n1096), .ZN(new_n1097));
  INV_X1    g672(.A(new_n1028), .ZN(new_n1098));
  NAND2_X1  g673(.A1(new_n988), .A2(new_n1098), .ZN(new_n1099));
  AOI21_X1  g674(.A(new_n1094), .B1(new_n1097), .B2(new_n1099), .ZN(new_n1100));
  OAI21_X1  g675(.A(KEYINPUT51), .B1(new_n1100), .B2(new_n1091), .ZN(new_n1101));
  NAND2_X1  g676(.A1(new_n1093), .A2(new_n1101), .ZN(new_n1102));
  OAI21_X1  g677(.A(new_n1091), .B1(new_n1026), .B2(new_n1029), .ZN(new_n1103));
  NAND2_X1  g678(.A1(new_n1102), .A2(new_n1103), .ZN(new_n1104));
  XNOR2_X1  g679(.A(KEYINPUT124), .B(G1961), .ZN(new_n1105));
  INV_X1    g680(.A(new_n1095), .ZN(new_n1106));
  INV_X1    g681(.A(KEYINPUT53), .ZN(new_n1107));
  NOR2_X1   g682(.A1(new_n1107), .A2(G2078), .ZN(new_n1108));
  AOI22_X1  g683(.A1(new_n989), .A2(new_n1105), .B1(new_n1106), .B2(new_n1108), .ZN(new_n1109));
  NAND4_X1  g684(.A1(new_n951), .A2(new_n443), .A3(new_n958), .A4(new_n963), .ZN(new_n1110));
  NAND2_X1  g685(.A1(new_n1110), .A2(new_n1107), .ZN(new_n1111));
  NAND3_X1  g686(.A1(new_n1109), .A2(new_n1111), .A3(G301), .ZN(new_n1112));
  INV_X1    g687(.A(new_n1108), .ZN(new_n1113));
  INV_X1    g688(.A(KEYINPUT111), .ZN(new_n1114));
  AOI21_X1  g689(.A(KEYINPUT45), .B1(new_n966), .B2(new_n1114), .ZN(new_n1115));
  NAND2_X1  g690(.A1(new_n962), .A2(KEYINPUT111), .ZN(new_n1116));
  AOI21_X1  g691(.A(new_n1113), .B1(new_n1115), .B2(new_n1116), .ZN(new_n1117));
  AOI22_X1  g692(.A1(new_n989), .A2(new_n1105), .B1(new_n963), .B2(new_n1117), .ZN(new_n1118));
  AND2_X1   g693(.A1(new_n1111), .A2(new_n1118), .ZN(new_n1119));
  OAI211_X1 g694(.A(KEYINPUT54), .B(new_n1112), .C1(new_n1119), .C2(G301), .ZN(new_n1120));
  INV_X1    g695(.A(KEYINPUT54), .ZN(new_n1121));
  AND3_X1   g696(.A1(new_n1111), .A2(G301), .A3(new_n1118), .ZN(new_n1122));
  AOI21_X1  g697(.A(G301), .B1(new_n1109), .B2(new_n1111), .ZN(new_n1123));
  OAI21_X1  g698(.A(new_n1121), .B1(new_n1122), .B2(new_n1123), .ZN(new_n1124));
  AND3_X1   g699(.A1(new_n1104), .A2(new_n1120), .A3(new_n1124), .ZN(new_n1125));
  NAND2_X1  g700(.A1(new_n1104), .A2(KEYINPUT62), .ZN(new_n1126));
  INV_X1    g701(.A(new_n1123), .ZN(new_n1127));
  INV_X1    g702(.A(new_n1103), .ZN(new_n1128));
  AOI21_X1  g703(.A(new_n1128), .B1(new_n1093), .B2(new_n1101), .ZN(new_n1129));
  INV_X1    g704(.A(KEYINPUT62), .ZN(new_n1130));
  AOI21_X1  g705(.A(new_n1127), .B1(new_n1129), .B2(new_n1130), .ZN(new_n1131));
  AOI22_X1  g706(.A1(new_n1087), .A2(new_n1125), .B1(new_n1126), .B2(new_n1131), .ZN(new_n1132));
  NAND3_X1  g707(.A1(new_n984), .A2(new_n994), .A3(new_n1022), .ZN(new_n1133));
  OAI211_X1 g708(.A(new_n1047), .B(new_n1053), .C1(new_n1132), .C2(new_n1133), .ZN(new_n1134));
  AND2_X1   g709(.A1(new_n1115), .A2(new_n1116), .ZN(new_n1135));
  NAND2_X1  g710(.A1(new_n1135), .A2(new_n976), .ZN(new_n1136));
  XNOR2_X1  g711(.A(new_n767), .B(G2067), .ZN(new_n1137));
  AOI21_X1  g712(.A(new_n1137), .B1(new_n1079), .B2(new_n712), .ZN(new_n1138));
  NOR2_X1   g713(.A1(new_n1136), .A2(new_n1138), .ZN(new_n1139));
  INV_X1    g714(.A(KEYINPUT112), .ZN(new_n1140));
  INV_X1    g715(.A(new_n712), .ZN(new_n1141));
  NAND2_X1  g716(.A1(new_n1141), .A2(G1996), .ZN(new_n1142));
  OR3_X1    g717(.A1(new_n1136), .A2(new_n1140), .A3(new_n1142), .ZN(new_n1143));
  OAI21_X1  g718(.A(new_n1140), .B1(new_n1136), .B2(new_n1142), .ZN(new_n1144));
  AOI21_X1  g719(.A(new_n1139), .B1(new_n1143), .B2(new_n1144), .ZN(new_n1145));
  INV_X1    g720(.A(new_n1136), .ZN(new_n1146));
  NOR2_X1   g721(.A1(new_n813), .A2(new_n816), .ZN(new_n1147));
  AND2_X1   g722(.A1(new_n813), .A2(new_n816), .ZN(new_n1148));
  OAI21_X1  g723(.A(new_n1146), .B1(new_n1147), .B2(new_n1148), .ZN(new_n1149));
  AND2_X1   g724(.A1(new_n1145), .A2(new_n1149), .ZN(new_n1150));
  INV_X1    g725(.A(new_n1150), .ZN(new_n1151));
  XNOR2_X1  g726(.A(G290), .B(G1986), .ZN(new_n1152));
  AOI21_X1  g727(.A(new_n1151), .B1(new_n1146), .B2(new_n1152), .ZN(new_n1153));
  NAND2_X1  g728(.A1(new_n1134), .A2(new_n1153), .ZN(new_n1154));
  NAND2_X1  g729(.A1(new_n1145), .A2(new_n1147), .ZN(new_n1155));
  OAI21_X1  g730(.A(new_n1155), .B1(G2067), .B2(new_n767), .ZN(new_n1156));
  NAND2_X1  g731(.A1(new_n1156), .A2(new_n1146), .ZN(new_n1157));
  NOR3_X1   g732(.A1(new_n1136), .A2(G1986), .A3(G290), .ZN(new_n1158));
  XNOR2_X1  g733(.A(KEYINPUT126), .B(KEYINPUT48), .ZN(new_n1159));
  XNOR2_X1  g734(.A(new_n1158), .B(new_n1159), .ZN(new_n1160));
  NAND2_X1  g735(.A1(new_n1150), .A2(new_n1160), .ZN(new_n1161));
  AND2_X1   g736(.A1(new_n1157), .A2(new_n1161), .ZN(new_n1162));
  INV_X1    g737(.A(KEYINPUT127), .ZN(new_n1163));
  INV_X1    g738(.A(KEYINPUT125), .ZN(new_n1164));
  NOR2_X1   g739(.A1(new_n1136), .A2(G1996), .ZN(new_n1165));
  INV_X1    g740(.A(KEYINPUT46), .ZN(new_n1166));
  XNOR2_X1  g741(.A(new_n1165), .B(new_n1166), .ZN(new_n1167));
  OAI21_X1  g742(.A(new_n1146), .B1(new_n1141), .B2(new_n1137), .ZN(new_n1168));
  AOI21_X1  g743(.A(new_n1164), .B1(new_n1167), .B2(new_n1168), .ZN(new_n1169));
  INV_X1    g744(.A(new_n1169), .ZN(new_n1170));
  NAND3_X1  g745(.A1(new_n1167), .A2(new_n1164), .A3(new_n1168), .ZN(new_n1171));
  NAND3_X1  g746(.A1(new_n1170), .A2(KEYINPUT47), .A3(new_n1171), .ZN(new_n1172));
  INV_X1    g747(.A(KEYINPUT47), .ZN(new_n1173));
  INV_X1    g748(.A(new_n1171), .ZN(new_n1174));
  OAI21_X1  g749(.A(new_n1173), .B1(new_n1174), .B2(new_n1169), .ZN(new_n1175));
  NAND4_X1  g750(.A1(new_n1162), .A2(new_n1163), .A3(new_n1172), .A4(new_n1175), .ZN(new_n1176));
  NAND2_X1  g751(.A1(new_n1175), .A2(new_n1172), .ZN(new_n1177));
  NAND2_X1  g752(.A1(new_n1157), .A2(new_n1161), .ZN(new_n1178));
  OAI21_X1  g753(.A(KEYINPUT127), .B1(new_n1177), .B2(new_n1178), .ZN(new_n1179));
  NAND2_X1  g754(.A1(new_n1176), .A2(new_n1179), .ZN(new_n1180));
  NAND2_X1  g755(.A1(new_n1154), .A2(new_n1180), .ZN(G329));
  assign    G231 = 1'b0;
  OR3_X1    g756(.A1(G227), .A2(new_n462), .A3(G401), .ZN(new_n1183));
  NOR2_X1   g757(.A1(G229), .A2(new_n1183), .ZN(new_n1184));
  NAND2_X1  g758(.A1(new_n930), .A2(new_n939), .ZN(new_n1185));
  AND3_X1   g759(.A1(new_n1184), .A2(new_n867), .A3(new_n1185), .ZN(G308));
  NAND3_X1  g760(.A1(new_n1184), .A2(new_n867), .A3(new_n1185), .ZN(G225));
endmodule


