//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 1 0 1 1 1 0 0 0 0 0 0 1 0 0 1 1 1 1 1 1 1 1 0 0 0 1 1 1 1 0 0 0 0 1 1 0 0 0 0 1 1 0 0 1 1 1 1 1 0 1 1 0 1 0 1 1 1 0 0 1 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:42:07 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n241, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1087,
    new_n1088, new_n1089, new_n1090, new_n1091, new_n1092, new_n1093,
    new_n1094, new_n1095, new_n1096, new_n1097, new_n1098, new_n1099,
    new_n1100, new_n1101, new_n1102, new_n1103, new_n1104, new_n1105,
    new_n1107, new_n1108, new_n1109, new_n1110, new_n1111, new_n1112,
    new_n1113, new_n1114, new_n1115, new_n1116, new_n1117, new_n1118,
    new_n1119, new_n1120, new_n1121, new_n1122, new_n1123, new_n1124,
    new_n1125, new_n1126, new_n1127, new_n1128, new_n1129, new_n1130,
    new_n1131, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1186, new_n1187, new_n1188, new_n1189, new_n1190, new_n1191,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1249, new_n1250, new_n1251, new_n1252, new_n1253,
    new_n1254, new_n1255, new_n1256, new_n1257, new_n1258, new_n1259,
    new_n1260, new_n1261, new_n1262, new_n1263, new_n1264, new_n1265,
    new_n1266, new_n1268, new_n1269, new_n1270, new_n1271, new_n1272,
    new_n1273, new_n1274, new_n1275, new_n1276, new_n1277, new_n1278,
    new_n1279, new_n1280, new_n1281, new_n1283, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1342, new_n1343, new_n1344, new_n1345, new_n1346, new_n1347;
  NOR3_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G77), .ZN(new_n202));
  AND2_X1   g0002(.A1(new_n201), .A2(new_n202), .ZN(G353));
  OAI21_X1  g0003(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0004(.A(G1), .ZN(new_n205));
  INV_X1    g0005(.A(G20), .ZN(new_n206));
  NOR2_X1   g0006(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  XOR2_X1   g0007(.A(new_n207), .B(KEYINPUT64), .Z(new_n208));
  NOR2_X1   g0008(.A1(new_n208), .A2(G13), .ZN(new_n209));
  OAI211_X1 g0009(.A(new_n209), .B(G250), .C1(G257), .C2(G264), .ZN(new_n210));
  INV_X1    g0010(.A(KEYINPUT0), .ZN(new_n211));
  NAND2_X1  g0011(.A1(G1), .A2(G13), .ZN(new_n212));
  NOR2_X1   g0012(.A1(new_n212), .A2(new_n206), .ZN(new_n213));
  OAI21_X1  g0013(.A(G50), .B1(G58), .B2(G68), .ZN(new_n214));
  XOR2_X1   g0014(.A(new_n214), .B(KEYINPUT65), .Z(new_n215));
  AOI22_X1  g0015(.A1(new_n210), .A2(new_n211), .B1(new_n213), .B2(new_n215), .ZN(new_n216));
  OAI21_X1  g0016(.A(new_n216), .B1(new_n211), .B2(new_n210), .ZN(new_n217));
  AOI22_X1  g0017(.A1(G87), .A2(G250), .B1(G107), .B2(G264), .ZN(new_n218));
  INV_X1    g0018(.A(G58), .ZN(new_n219));
  INV_X1    g0019(.A(G232), .ZN(new_n220));
  INV_X1    g0020(.A(G97), .ZN(new_n221));
  INV_X1    g0021(.A(G257), .ZN(new_n222));
  OAI221_X1 g0022(.A(new_n218), .B1(new_n219), .B2(new_n220), .C1(new_n221), .C2(new_n222), .ZN(new_n223));
  NAND2_X1  g0023(.A1(new_n223), .A2(KEYINPUT66), .ZN(new_n224));
  AOI22_X1  g0024(.A1(G50), .A2(G226), .B1(G77), .B2(G244), .ZN(new_n225));
  AOI22_X1  g0025(.A1(G68), .A2(G238), .B1(G116), .B2(G270), .ZN(new_n226));
  NAND3_X1  g0026(.A1(new_n224), .A2(new_n225), .A3(new_n226), .ZN(new_n227));
  NOR2_X1   g0027(.A1(new_n223), .A2(KEYINPUT66), .ZN(new_n228));
  OAI21_X1  g0028(.A(new_n208), .B1(new_n227), .B2(new_n228), .ZN(new_n229));
  AND2_X1   g0029(.A1(new_n229), .A2(KEYINPUT1), .ZN(new_n230));
  NOR2_X1   g0030(.A1(new_n229), .A2(KEYINPUT1), .ZN(new_n231));
  NOR3_X1   g0031(.A1(new_n217), .A2(new_n230), .A3(new_n231), .ZN(G361));
  XNOR2_X1  g0032(.A(G238), .B(G244), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n233), .B(KEYINPUT2), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n234), .B(G226), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n235), .B(new_n220), .ZN(new_n236));
  XNOR2_X1  g0036(.A(G250), .B(G257), .ZN(new_n237));
  XNOR2_X1  g0037(.A(G264), .B(G270), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n236), .B(new_n239), .ZN(G358));
  XOR2_X1   g0040(.A(G68), .B(G77), .Z(new_n241));
  XNOR2_X1  g0041(.A(G50), .B(G58), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XOR2_X1   g0043(.A(G87), .B(G97), .Z(new_n244));
  XNOR2_X1  g0044(.A(G107), .B(G116), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n244), .B(new_n245), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n243), .B(new_n246), .ZN(G351));
  OR2_X1    g0047(.A1(KEYINPUT3), .A2(G33), .ZN(new_n248));
  NAND2_X1  g0048(.A1(KEYINPUT3), .A2(G33), .ZN(new_n249));
  NAND2_X1  g0049(.A1(new_n248), .A2(new_n249), .ZN(new_n250));
  AND2_X1   g0050(.A1(KEYINPUT68), .A2(G1698), .ZN(new_n251));
  NOR2_X1   g0051(.A1(KEYINPUT68), .A2(G1698), .ZN(new_n252));
  NOR2_X1   g0052(.A1(new_n251), .A2(new_n252), .ZN(new_n253));
  NAND3_X1  g0053(.A1(new_n250), .A2(new_n253), .A3(G222), .ZN(new_n254));
  INV_X1    g0054(.A(G223), .ZN(new_n255));
  NAND2_X1  g0055(.A1(new_n250), .A2(G1698), .ZN(new_n256));
  OAI221_X1 g0056(.A(new_n254), .B1(new_n202), .B2(new_n250), .C1(new_n255), .C2(new_n256), .ZN(new_n257));
  AOI21_X1  g0057(.A(new_n212), .B1(G33), .B2(G41), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n257), .A2(new_n258), .ZN(new_n259));
  OAI21_X1  g0059(.A(new_n205), .B1(G41), .B2(G45), .ZN(new_n260));
  INV_X1    g0060(.A(G274), .ZN(new_n261));
  NOR2_X1   g0061(.A1(new_n260), .A2(new_n261), .ZN(new_n262));
  INV_X1    g0062(.A(KEYINPUT67), .ZN(new_n263));
  OR2_X1    g0063(.A1(new_n260), .A2(new_n263), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n260), .A2(new_n263), .ZN(new_n265));
  AOI21_X1  g0065(.A(new_n258), .B1(new_n264), .B2(new_n265), .ZN(new_n266));
  AOI21_X1  g0066(.A(new_n262), .B1(new_n266), .B2(G226), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n259), .A2(new_n267), .ZN(new_n268));
  INV_X1    g0068(.A(new_n268), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n269), .A2(G190), .ZN(new_n270));
  INV_X1    g0070(.A(G150), .ZN(new_n271));
  NOR2_X1   g0071(.A1(G20), .A2(G33), .ZN(new_n272));
  INV_X1    g0072(.A(new_n272), .ZN(new_n273));
  OAI22_X1  g0073(.A1(new_n271), .A2(new_n273), .B1(new_n201), .B2(new_n206), .ZN(new_n274));
  XNOR2_X1  g0074(.A(KEYINPUT8), .B(G58), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n206), .A2(G33), .ZN(new_n276));
  NOR2_X1   g0076(.A1(new_n275), .A2(new_n276), .ZN(new_n277));
  OR2_X1    g0077(.A1(new_n274), .A2(new_n277), .ZN(new_n278));
  NAND3_X1  g0078(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n279));
  NAND2_X1  g0079(.A1(new_n279), .A2(new_n212), .ZN(new_n280));
  INV_X1    g0080(.A(KEYINPUT69), .ZN(new_n281));
  NAND2_X1  g0081(.A1(new_n280), .A2(new_n281), .ZN(new_n282));
  NAND3_X1  g0082(.A1(new_n279), .A2(KEYINPUT69), .A3(new_n212), .ZN(new_n283));
  AND2_X1   g0083(.A1(new_n282), .A2(new_n283), .ZN(new_n284));
  INV_X1    g0084(.A(G50), .ZN(new_n285));
  INV_X1    g0085(.A(G13), .ZN(new_n286));
  NOR2_X1   g0086(.A1(new_n286), .A2(G1), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n287), .A2(G20), .ZN(new_n288));
  INV_X1    g0088(.A(new_n288), .ZN(new_n289));
  AOI22_X1  g0089(.A1(new_n278), .A2(new_n284), .B1(new_n285), .B2(new_n289), .ZN(new_n290));
  NOR2_X1   g0090(.A1(new_n284), .A2(new_n289), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n205), .A2(G20), .ZN(new_n292));
  NAND3_X1  g0092(.A1(new_n291), .A2(G50), .A3(new_n292), .ZN(new_n293));
  NAND2_X1  g0093(.A1(new_n290), .A2(new_n293), .ZN(new_n294));
  INV_X1    g0094(.A(KEYINPUT9), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n294), .A2(new_n295), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n268), .A2(G200), .ZN(new_n297));
  NAND3_X1  g0097(.A1(new_n290), .A2(new_n293), .A3(KEYINPUT9), .ZN(new_n298));
  NAND4_X1  g0098(.A1(new_n270), .A2(new_n296), .A3(new_n297), .A4(new_n298), .ZN(new_n299));
  INV_X1    g0099(.A(KEYINPUT10), .ZN(new_n300));
  XNOR2_X1  g0100(.A(new_n299), .B(new_n300), .ZN(new_n301));
  INV_X1    g0101(.A(new_n294), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n269), .A2(G179), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n268), .A2(G169), .ZN(new_n304));
  AOI21_X1  g0104(.A(new_n302), .B1(new_n303), .B2(new_n304), .ZN(new_n305));
  NOR2_X1   g0105(.A1(new_n301), .A2(new_n305), .ZN(new_n306));
  OR3_X1    g0106(.A1(new_n273), .A2(KEYINPUT76), .A3(new_n285), .ZN(new_n307));
  INV_X1    g0107(.A(G68), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n308), .A2(G20), .ZN(new_n309));
  OAI21_X1  g0109(.A(KEYINPUT76), .B1(new_n273), .B2(new_n285), .ZN(new_n310));
  NAND3_X1  g0110(.A1(new_n206), .A2(G33), .A3(G77), .ZN(new_n311));
  NAND4_X1  g0111(.A1(new_n307), .A2(new_n309), .A3(new_n310), .A4(new_n311), .ZN(new_n312));
  AOI21_X1  g0112(.A(KEYINPUT11), .B1(new_n312), .B2(new_n284), .ZN(new_n313));
  NAND3_X1  g0113(.A1(new_n287), .A2(G20), .A3(new_n308), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n314), .A2(KEYINPUT12), .ZN(new_n315));
  OR2_X1    g0115(.A1(new_n314), .A2(KEYINPUT12), .ZN(new_n316));
  AOI21_X1  g0116(.A(new_n313), .B1(new_n315), .B2(new_n316), .ZN(new_n317));
  NAND3_X1  g0117(.A1(new_n312), .A2(KEYINPUT11), .A3(new_n284), .ZN(new_n318));
  NAND3_X1  g0118(.A1(new_n291), .A2(G68), .A3(new_n292), .ZN(new_n319));
  NAND3_X1  g0119(.A1(new_n317), .A2(new_n318), .A3(new_n319), .ZN(new_n320));
  NAND3_X1  g0120(.A1(new_n250), .A2(new_n253), .A3(G226), .ZN(new_n321));
  NAND2_X1  g0121(.A1(G33), .A2(G97), .ZN(new_n322));
  OAI211_X1 g0122(.A(new_n321), .B(new_n322), .C1(new_n220), .C2(new_n256), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n323), .A2(new_n258), .ZN(new_n324));
  AOI21_X1  g0124(.A(new_n262), .B1(new_n266), .B2(G238), .ZN(new_n325));
  XNOR2_X1  g0125(.A(KEYINPUT73), .B(KEYINPUT13), .ZN(new_n326));
  AND3_X1   g0126(.A1(new_n324), .A2(new_n325), .A3(new_n326), .ZN(new_n327));
  AOI21_X1  g0127(.A(new_n326), .B1(new_n324), .B2(new_n325), .ZN(new_n328));
  OAI21_X1  g0128(.A(G169), .B1(new_n327), .B2(new_n328), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n329), .A2(KEYINPUT14), .ZN(new_n330));
  INV_X1    g0130(.A(KEYINPUT14), .ZN(new_n331));
  OAI211_X1 g0131(.A(new_n331), .B(G169), .C1(new_n327), .C2(new_n328), .ZN(new_n332));
  INV_X1    g0132(.A(KEYINPUT13), .ZN(new_n333));
  AOI21_X1  g0133(.A(new_n333), .B1(new_n324), .B2(new_n325), .ZN(new_n334));
  INV_X1    g0134(.A(new_n334), .ZN(new_n335));
  NAND3_X1  g0135(.A1(new_n324), .A2(new_n325), .A3(new_n326), .ZN(new_n336));
  NAND3_X1  g0136(.A1(new_n335), .A2(G179), .A3(new_n336), .ZN(new_n337));
  NAND3_X1  g0137(.A1(new_n330), .A2(new_n332), .A3(new_n337), .ZN(new_n338));
  INV_X1    g0138(.A(KEYINPUT75), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n336), .A2(G190), .ZN(new_n340));
  OAI21_X1  g0140(.A(new_n339), .B1(new_n340), .B2(new_n334), .ZN(new_n341));
  NAND4_X1  g0141(.A1(new_n335), .A2(KEYINPUT75), .A3(G190), .A4(new_n336), .ZN(new_n342));
  AOI21_X1  g0142(.A(new_n320), .B1(new_n341), .B2(new_n342), .ZN(new_n343));
  OAI21_X1  g0143(.A(G200), .B1(new_n327), .B2(new_n328), .ZN(new_n344));
  INV_X1    g0144(.A(KEYINPUT74), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n344), .A2(new_n345), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n324), .A2(new_n325), .ZN(new_n347));
  INV_X1    g0147(.A(new_n326), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n347), .A2(new_n348), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n349), .A2(new_n336), .ZN(new_n350));
  NAND3_X1  g0150(.A1(new_n350), .A2(KEYINPUT74), .A3(G200), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n346), .A2(new_n351), .ZN(new_n352));
  AOI22_X1  g0152(.A1(new_n320), .A2(new_n338), .B1(new_n343), .B2(new_n352), .ZN(new_n353));
  NOR2_X1   g0153(.A1(new_n275), .A2(new_n273), .ZN(new_n354));
  XNOR2_X1  g0154(.A(KEYINPUT15), .B(G87), .ZN(new_n355));
  OAI22_X1  g0155(.A1(new_n355), .A2(new_n276), .B1(new_n206), .B2(new_n202), .ZN(new_n356));
  OAI21_X1  g0156(.A(new_n284), .B1(new_n354), .B2(new_n356), .ZN(new_n357));
  INV_X1    g0157(.A(KEYINPUT72), .ZN(new_n358));
  XNOR2_X1  g0158(.A(new_n357), .B(new_n358), .ZN(new_n359));
  AOI21_X1  g0159(.A(new_n202), .B1(new_n205), .B2(G20), .ZN(new_n360));
  AOI22_X1  g0160(.A1(new_n291), .A2(new_n360), .B1(new_n202), .B2(new_n289), .ZN(new_n361));
  AND2_X1   g0161(.A1(new_n359), .A2(new_n361), .ZN(new_n362));
  INV_X1    g0162(.A(new_n362), .ZN(new_n363));
  AND2_X1   g0163(.A1(KEYINPUT3), .A2(G33), .ZN(new_n364));
  NOR2_X1   g0164(.A1(KEYINPUT3), .A2(G33), .ZN(new_n365));
  OAI211_X1 g0165(.A(G238), .B(G1698), .C1(new_n364), .C2(new_n365), .ZN(new_n366));
  NAND3_X1  g0166(.A1(new_n248), .A2(G107), .A3(new_n249), .ZN(new_n367));
  OR2_X1    g0167(.A1(KEYINPUT68), .A2(G1698), .ZN(new_n368));
  NAND2_X1  g0168(.A1(KEYINPUT68), .A2(G1698), .ZN(new_n369));
  OAI211_X1 g0169(.A(new_n368), .B(new_n369), .C1(new_n364), .C2(new_n365), .ZN(new_n370));
  OAI211_X1 g0170(.A(new_n366), .B(new_n367), .C1(new_n370), .C2(new_n220), .ZN(new_n371));
  INV_X1    g0171(.A(KEYINPUT70), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n371), .A2(new_n372), .ZN(new_n373));
  NAND3_X1  g0173(.A1(new_n250), .A2(new_n253), .A3(G232), .ZN(new_n374));
  NAND4_X1  g0174(.A1(new_n374), .A2(KEYINPUT70), .A3(new_n366), .A4(new_n367), .ZN(new_n375));
  NAND3_X1  g0175(.A1(new_n373), .A2(new_n258), .A3(new_n375), .ZN(new_n376));
  INV_X1    g0176(.A(KEYINPUT71), .ZN(new_n377));
  AOI21_X1  g0177(.A(new_n262), .B1(new_n266), .B2(G244), .ZN(new_n378));
  AND3_X1   g0178(.A1(new_n376), .A2(new_n377), .A3(new_n378), .ZN(new_n379));
  AOI21_X1  g0179(.A(new_n377), .B1(new_n376), .B2(new_n378), .ZN(new_n380));
  INV_X1    g0180(.A(G169), .ZN(new_n381));
  NOR3_X1   g0181(.A1(new_n379), .A2(new_n380), .A3(new_n381), .ZN(new_n382));
  INV_X1    g0182(.A(G179), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n376), .A2(new_n378), .ZN(new_n384));
  NAND2_X1  g0184(.A1(new_n384), .A2(KEYINPUT71), .ZN(new_n385));
  NAND3_X1  g0185(.A1(new_n376), .A2(new_n377), .A3(new_n378), .ZN(new_n386));
  AOI21_X1  g0186(.A(new_n383), .B1(new_n385), .B2(new_n386), .ZN(new_n387));
  OAI21_X1  g0187(.A(new_n363), .B1(new_n382), .B2(new_n387), .ZN(new_n388));
  INV_X1    g0188(.A(G190), .ZN(new_n389));
  OAI21_X1  g0189(.A(new_n389), .B1(new_n379), .B2(new_n380), .ZN(new_n390));
  INV_X1    g0190(.A(G200), .ZN(new_n391));
  NAND3_X1  g0191(.A1(new_n385), .A2(new_n391), .A3(new_n386), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n390), .A2(new_n392), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n393), .A2(new_n362), .ZN(new_n394));
  NAND4_X1  g0194(.A1(new_n306), .A2(new_n353), .A3(new_n388), .A4(new_n394), .ZN(new_n395));
  AOI21_X1  g0195(.A(new_n275), .B1(new_n205), .B2(G20), .ZN(new_n396));
  AOI22_X1  g0196(.A1(new_n291), .A2(new_n396), .B1(new_n289), .B2(new_n275), .ZN(new_n397));
  INV_X1    g0197(.A(new_n397), .ZN(new_n398));
  INV_X1    g0198(.A(KEYINPUT78), .ZN(new_n399));
  NOR2_X1   g0199(.A1(new_n364), .A2(new_n365), .ZN(new_n400));
  AOI21_X1  g0200(.A(KEYINPUT7), .B1(new_n400), .B2(new_n206), .ZN(new_n401));
  INV_X1    g0201(.A(KEYINPUT7), .ZN(new_n402));
  NOR4_X1   g0202(.A1(new_n364), .A2(new_n365), .A3(new_n402), .A4(G20), .ZN(new_n403));
  OAI211_X1 g0203(.A(KEYINPUT77), .B(G68), .C1(new_n401), .C2(new_n403), .ZN(new_n404));
  NOR2_X1   g0204(.A1(new_n219), .A2(new_n308), .ZN(new_n405));
  NOR2_X1   g0205(.A1(G58), .A2(G68), .ZN(new_n406));
  OAI21_X1  g0206(.A(G20), .B1(new_n405), .B2(new_n406), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n272), .A2(G159), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n407), .A2(new_n408), .ZN(new_n409));
  INV_X1    g0209(.A(new_n409), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n404), .A2(new_n410), .ZN(new_n411));
  NAND3_X1  g0211(.A1(new_n248), .A2(new_n206), .A3(new_n249), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n412), .A2(new_n402), .ZN(new_n413));
  NAND3_X1  g0213(.A1(new_n400), .A2(KEYINPUT7), .A3(new_n206), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n413), .A2(new_n414), .ZN(new_n415));
  AOI21_X1  g0215(.A(KEYINPUT77), .B1(new_n415), .B2(G68), .ZN(new_n416));
  INV_X1    g0216(.A(KEYINPUT16), .ZN(new_n417));
  NOR3_X1   g0217(.A1(new_n411), .A2(new_n416), .A3(new_n417), .ZN(new_n418));
  AOI21_X1  g0218(.A(new_n308), .B1(new_n413), .B2(new_n414), .ZN(new_n419));
  OAI21_X1  g0219(.A(new_n417), .B1(new_n419), .B2(new_n409), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n420), .A2(new_n284), .ZN(new_n421));
  OAI21_X1  g0221(.A(new_n399), .B1(new_n418), .B2(new_n421), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n282), .A2(new_n283), .ZN(new_n423));
  OAI21_X1  g0223(.A(G68), .B1(new_n401), .B2(new_n403), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n424), .A2(new_n410), .ZN(new_n425));
  AOI21_X1  g0225(.A(new_n423), .B1(new_n425), .B2(new_n417), .ZN(new_n426));
  INV_X1    g0226(.A(KEYINPUT77), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n424), .A2(new_n427), .ZN(new_n428));
  NAND4_X1  g0228(.A1(new_n428), .A2(KEYINPUT16), .A3(new_n404), .A4(new_n410), .ZN(new_n429));
  NAND3_X1  g0229(.A1(new_n426), .A2(new_n429), .A3(KEYINPUT78), .ZN(new_n430));
  AOI21_X1  g0230(.A(new_n398), .B1(new_n422), .B2(new_n430), .ZN(new_n431));
  NAND3_X1  g0231(.A1(new_n250), .A2(G226), .A3(G1698), .ZN(new_n432));
  INV_X1    g0232(.A(G33), .ZN(new_n433));
  INV_X1    g0233(.A(G87), .ZN(new_n434));
  OAI221_X1 g0234(.A(new_n432), .B1(new_n433), .B2(new_n434), .C1(new_n255), .C2(new_n370), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n435), .A2(new_n258), .ZN(new_n436));
  AOI21_X1  g0236(.A(new_n262), .B1(new_n266), .B2(G232), .ZN(new_n437));
  AND3_X1   g0237(.A1(new_n436), .A2(new_n383), .A3(new_n437), .ZN(new_n438));
  AOI21_X1  g0238(.A(G169), .B1(new_n436), .B2(new_n437), .ZN(new_n439));
  NOR2_X1   g0239(.A1(new_n438), .A2(new_n439), .ZN(new_n440));
  INV_X1    g0240(.A(new_n440), .ZN(new_n441));
  OAI21_X1  g0241(.A(KEYINPUT18), .B1(new_n431), .B2(new_n441), .ZN(new_n442));
  AND3_X1   g0242(.A1(new_n426), .A2(new_n429), .A3(KEYINPUT78), .ZN(new_n443));
  AOI21_X1  g0243(.A(KEYINPUT78), .B1(new_n426), .B2(new_n429), .ZN(new_n444));
  OAI21_X1  g0244(.A(new_n397), .B1(new_n443), .B2(new_n444), .ZN(new_n445));
  INV_X1    g0245(.A(KEYINPUT18), .ZN(new_n446));
  NAND3_X1  g0246(.A1(new_n445), .A2(new_n440), .A3(new_n446), .ZN(new_n447));
  NAND2_X1  g0247(.A1(new_n436), .A2(new_n437), .ZN(new_n448));
  NAND2_X1  g0248(.A1(new_n448), .A2(new_n391), .ZN(new_n449));
  NAND3_X1  g0249(.A1(new_n436), .A2(new_n389), .A3(new_n437), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n449), .A2(new_n450), .ZN(new_n451));
  OAI211_X1 g0251(.A(new_n451), .B(new_n397), .C1(new_n443), .C2(new_n444), .ZN(new_n452));
  INV_X1    g0252(.A(KEYINPUT17), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n452), .A2(new_n453), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n422), .A2(new_n430), .ZN(new_n455));
  NAND4_X1  g0255(.A1(new_n455), .A2(KEYINPUT17), .A3(new_n397), .A4(new_n451), .ZN(new_n456));
  NAND4_X1  g0256(.A1(new_n442), .A2(new_n447), .A3(new_n454), .A4(new_n456), .ZN(new_n457));
  NOR2_X1   g0257(.A1(new_n395), .A2(new_n457), .ZN(new_n458));
  INV_X1    g0258(.A(KEYINPUT21), .ZN(new_n459));
  NAND2_X1  g0259(.A1(G33), .A2(G283), .ZN(new_n460));
  OAI21_X1  g0260(.A(new_n460), .B1(new_n221), .B2(G33), .ZN(new_n461));
  AND2_X1   g0261(.A1(new_n461), .A2(new_n206), .ZN(new_n462));
  INV_X1    g0262(.A(G116), .ZN(new_n463));
  NOR2_X1   g0263(.A1(new_n206), .A2(new_n463), .ZN(new_n464));
  OAI211_X1 g0264(.A(KEYINPUT20), .B(new_n280), .C1(new_n462), .C2(new_n464), .ZN(new_n465));
  INV_X1    g0265(.A(KEYINPUT20), .ZN(new_n466));
  AOI21_X1  g0266(.A(new_n464), .B1(new_n461), .B2(new_n206), .ZN(new_n467));
  INV_X1    g0267(.A(new_n280), .ZN(new_n468));
  OAI21_X1  g0268(.A(new_n466), .B1(new_n467), .B2(new_n468), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n465), .A2(new_n469), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n205), .A2(G33), .ZN(new_n471));
  NAND4_X1  g0271(.A1(new_n423), .A2(G116), .A3(new_n288), .A4(new_n471), .ZN(new_n472));
  NAND2_X1  g0272(.A1(new_n289), .A2(new_n463), .ZN(new_n473));
  AND3_X1   g0273(.A1(new_n470), .A2(new_n472), .A3(new_n473), .ZN(new_n474));
  INV_X1    g0274(.A(new_n258), .ZN(new_n475));
  INV_X1    g0275(.A(KEYINPUT5), .ZN(new_n476));
  INV_X1    g0276(.A(KEYINPUT81), .ZN(new_n477));
  OAI21_X1  g0277(.A(new_n476), .B1(new_n477), .B2(G41), .ZN(new_n478));
  INV_X1    g0278(.A(G41), .ZN(new_n479));
  NAND3_X1  g0279(.A1(new_n479), .A2(KEYINPUT81), .A3(KEYINPUT5), .ZN(new_n480));
  INV_X1    g0280(.A(G45), .ZN(new_n481));
  NOR2_X1   g0281(.A1(new_n481), .A2(G1), .ZN(new_n482));
  NAND3_X1  g0282(.A1(new_n478), .A2(new_n480), .A3(new_n482), .ZN(new_n483));
  NAND3_X1  g0283(.A1(new_n475), .A2(new_n483), .A3(G270), .ZN(new_n484));
  NAND4_X1  g0284(.A1(new_n478), .A2(new_n480), .A3(new_n482), .A4(G274), .ZN(new_n485));
  AND2_X1   g0285(.A1(new_n484), .A2(new_n485), .ZN(new_n486));
  OAI211_X1 g0286(.A(G264), .B(G1698), .C1(new_n364), .C2(new_n365), .ZN(new_n487));
  NAND3_X1  g0287(.A1(new_n248), .A2(G303), .A3(new_n249), .ZN(new_n488));
  OAI211_X1 g0288(.A(new_n487), .B(new_n488), .C1(new_n370), .C2(new_n222), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n489), .A2(new_n258), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n486), .A2(new_n490), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n491), .A2(G169), .ZN(new_n492));
  OAI21_X1  g0292(.A(new_n459), .B1(new_n474), .B2(new_n492), .ZN(new_n493));
  NOR2_X1   g0293(.A1(new_n491), .A2(G190), .ZN(new_n494));
  AOI21_X1  g0294(.A(G200), .B1(new_n486), .B2(new_n490), .ZN(new_n495));
  OAI21_X1  g0295(.A(new_n474), .B1(new_n494), .B2(new_n495), .ZN(new_n496));
  AOI21_X1  g0296(.A(new_n381), .B1(new_n486), .B2(new_n490), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n484), .A2(new_n485), .ZN(new_n498));
  AOI21_X1  g0298(.A(new_n498), .B1(new_n258), .B2(new_n489), .ZN(new_n499));
  AOI22_X1  g0299(.A1(new_n497), .A2(KEYINPUT21), .B1(new_n499), .B2(G179), .ZN(new_n500));
  OAI211_X1 g0300(.A(new_n493), .B(new_n496), .C1(new_n474), .C2(new_n500), .ZN(new_n501));
  INV_X1    g0301(.A(KEYINPUT85), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  NAND3_X1  g0303(.A1(new_n486), .A2(new_n490), .A3(G179), .ZN(new_n504));
  OAI21_X1  g0304(.A(new_n504), .B1(new_n492), .B2(new_n459), .ZN(new_n505));
  INV_X1    g0305(.A(new_n474), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  NAND4_X1  g0307(.A1(new_n507), .A2(KEYINPUT85), .A3(new_n496), .A4(new_n493), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n503), .A2(new_n508), .ZN(new_n509));
  INV_X1    g0309(.A(new_n355), .ZN(new_n510));
  NOR2_X1   g0310(.A1(new_n510), .A2(new_n288), .ZN(new_n511));
  NAND3_X1  g0311(.A1(new_n423), .A2(new_n288), .A3(new_n471), .ZN(new_n512));
  NOR2_X1   g0312(.A1(new_n512), .A2(new_n434), .ZN(new_n513));
  OAI211_X1 g0313(.A(new_n206), .B(G68), .C1(new_n364), .C2(new_n365), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n514), .A2(KEYINPUT83), .ZN(new_n515));
  INV_X1    g0315(.A(KEYINPUT83), .ZN(new_n516));
  NAND4_X1  g0316(.A1(new_n250), .A2(new_n516), .A3(new_n206), .A4(G68), .ZN(new_n517));
  NOR3_X1   g0317(.A1(G87), .A2(G97), .A3(G107), .ZN(new_n518));
  AOI21_X1  g0318(.A(G20), .B1(G33), .B2(G97), .ZN(new_n519));
  OAI21_X1  g0319(.A(KEYINPUT19), .B1(new_n518), .B2(new_n519), .ZN(new_n520));
  OR3_X1    g0320(.A1(new_n322), .A2(KEYINPUT19), .A3(G20), .ZN(new_n521));
  AOI22_X1  g0321(.A1(new_n515), .A2(new_n517), .B1(new_n520), .B2(new_n521), .ZN(new_n522));
  AOI21_X1  g0322(.A(new_n423), .B1(new_n522), .B2(KEYINPUT84), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n520), .A2(new_n521), .ZN(new_n524));
  AOI21_X1  g0324(.A(G20), .B1(new_n248), .B2(new_n249), .ZN(new_n525));
  AOI21_X1  g0325(.A(new_n516), .B1(new_n525), .B2(G68), .ZN(new_n526));
  NOR2_X1   g0326(.A1(new_n514), .A2(KEYINPUT83), .ZN(new_n527));
  OAI21_X1  g0327(.A(new_n524), .B1(new_n526), .B2(new_n527), .ZN(new_n528));
  INV_X1    g0328(.A(KEYINPUT84), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  AOI211_X1 g0330(.A(new_n511), .B(new_n513), .C1(new_n523), .C2(new_n530), .ZN(new_n531));
  OAI21_X1  g0331(.A(G250), .B1(new_n481), .B2(G1), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n482), .A2(G274), .ZN(new_n533));
  AOI21_X1  g0333(.A(new_n258), .B1(new_n532), .B2(new_n533), .ZN(new_n534));
  OAI211_X1 g0334(.A(G244), .B(G1698), .C1(new_n364), .C2(new_n365), .ZN(new_n535));
  NAND2_X1  g0335(.A1(G33), .A2(G116), .ZN(new_n536));
  INV_X1    g0336(.A(G238), .ZN(new_n537));
  OAI211_X1 g0337(.A(new_n535), .B(new_n536), .C1(new_n370), .C2(new_n537), .ZN(new_n538));
  AOI21_X1  g0338(.A(new_n534), .B1(new_n538), .B2(new_n258), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n539), .A2(new_n389), .ZN(new_n540));
  OAI21_X1  g0340(.A(new_n540), .B1(G200), .B2(new_n539), .ZN(new_n541));
  INV_X1    g0341(.A(new_n511), .ZN(new_n542));
  INV_X1    g0342(.A(new_n512), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n543), .A2(new_n510), .ZN(new_n544));
  OAI211_X1 g0344(.A(KEYINPUT84), .B(new_n524), .C1(new_n526), .C2(new_n527), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n545), .A2(new_n284), .ZN(new_n546));
  NOR2_X1   g0346(.A1(new_n522), .A2(KEYINPUT84), .ZN(new_n547));
  OAI211_X1 g0347(.A(new_n542), .B(new_n544), .C1(new_n546), .C2(new_n547), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n539), .A2(G179), .ZN(new_n549));
  OAI21_X1  g0349(.A(new_n549), .B1(new_n381), .B2(new_n539), .ZN(new_n550));
  AOI22_X1  g0350(.A1(new_n531), .A2(new_n541), .B1(new_n548), .B2(new_n550), .ZN(new_n551));
  INV_X1    g0351(.A(KEYINPUT82), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n272), .A2(G77), .ZN(new_n553));
  XNOR2_X1  g0353(.A(new_n553), .B(KEYINPUT79), .ZN(new_n554));
  AOI21_X1  g0354(.A(new_n554), .B1(new_n415), .B2(G107), .ZN(new_n555));
  INV_X1    g0355(.A(KEYINPUT6), .ZN(new_n556));
  INV_X1    g0356(.A(G107), .ZN(new_n557));
  NOR2_X1   g0357(.A1(new_n221), .A2(new_n557), .ZN(new_n558));
  NOR2_X1   g0358(.A1(G97), .A2(G107), .ZN(new_n559));
  OAI21_X1  g0359(.A(new_n556), .B1(new_n558), .B2(new_n559), .ZN(new_n560));
  NAND2_X1  g0360(.A1(KEYINPUT6), .A2(G97), .ZN(new_n561));
  OAI21_X1  g0361(.A(KEYINPUT80), .B1(new_n561), .B2(G107), .ZN(new_n562));
  INV_X1    g0362(.A(KEYINPUT80), .ZN(new_n563));
  NAND4_X1  g0363(.A1(new_n563), .A2(new_n557), .A3(KEYINPUT6), .A4(G97), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n562), .A2(new_n564), .ZN(new_n565));
  AOI21_X1  g0365(.A(new_n206), .B1(new_n560), .B2(new_n565), .ZN(new_n566));
  INV_X1    g0366(.A(new_n566), .ZN(new_n567));
  AOI21_X1  g0367(.A(new_n423), .B1(new_n555), .B2(new_n567), .ZN(new_n568));
  NOR2_X1   g0368(.A1(new_n288), .A2(G97), .ZN(new_n569));
  INV_X1    g0369(.A(new_n569), .ZN(new_n570));
  OAI21_X1  g0370(.A(new_n570), .B1(new_n512), .B2(new_n221), .ZN(new_n571));
  OAI21_X1  g0371(.A(new_n552), .B1(new_n568), .B2(new_n571), .ZN(new_n572));
  INV_X1    g0372(.A(new_n571), .ZN(new_n573));
  AOI21_X1  g0373(.A(new_n557), .B1(new_n413), .B2(new_n414), .ZN(new_n574));
  NOR3_X1   g0374(.A1(new_n574), .A2(new_n566), .A3(new_n554), .ZN(new_n575));
  OAI211_X1 g0375(.A(new_n573), .B(KEYINPUT82), .C1(new_n423), .C2(new_n575), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n475), .A2(new_n483), .ZN(new_n577));
  OAI21_X1  g0377(.A(new_n485), .B1(new_n577), .B2(new_n222), .ZN(new_n578));
  NAND3_X1  g0378(.A1(new_n250), .A2(new_n253), .A3(G244), .ZN(new_n579));
  INV_X1    g0379(.A(KEYINPUT4), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  NAND4_X1  g0381(.A1(new_n250), .A2(new_n253), .A3(KEYINPUT4), .A4(G244), .ZN(new_n582));
  OAI211_X1 g0382(.A(G250), .B(G1698), .C1(new_n364), .C2(new_n365), .ZN(new_n583));
  AND2_X1   g0383(.A1(new_n583), .A2(new_n460), .ZN(new_n584));
  NAND3_X1  g0384(.A1(new_n581), .A2(new_n582), .A3(new_n584), .ZN(new_n585));
  AOI21_X1  g0385(.A(new_n578), .B1(new_n585), .B2(new_n258), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n586), .A2(new_n383), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n583), .A2(new_n460), .ZN(new_n588));
  AOI21_X1  g0388(.A(new_n588), .B1(new_n580), .B2(new_n579), .ZN(new_n589));
  AOI21_X1  g0389(.A(new_n475), .B1(new_n589), .B2(new_n582), .ZN(new_n590));
  OAI21_X1  g0390(.A(new_n381), .B1(new_n590), .B2(new_n578), .ZN(new_n591));
  NAND4_X1  g0391(.A1(new_n572), .A2(new_n576), .A3(new_n587), .A4(new_n591), .ZN(new_n592));
  NOR2_X1   g0392(.A1(new_n568), .A2(new_n571), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n585), .A2(new_n258), .ZN(new_n594));
  INV_X1    g0394(.A(new_n578), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n594), .A2(new_n595), .ZN(new_n596));
  NOR2_X1   g0396(.A1(new_n596), .A2(G190), .ZN(new_n597));
  NOR2_X1   g0397(.A1(new_n586), .A2(G200), .ZN(new_n598));
  OAI21_X1  g0398(.A(new_n593), .B1(new_n597), .B2(new_n598), .ZN(new_n599));
  AND3_X1   g0399(.A1(new_n551), .A2(new_n592), .A3(new_n599), .ZN(new_n600));
  NOR2_X1   g0400(.A1(new_n512), .A2(new_n557), .ZN(new_n601));
  NAND3_X1  g0401(.A1(new_n287), .A2(G20), .A3(new_n557), .ZN(new_n602));
  XNOR2_X1  g0402(.A(new_n602), .B(KEYINPUT25), .ZN(new_n603));
  NOR2_X1   g0403(.A1(new_n601), .A2(new_n603), .ZN(new_n604));
  INV_X1    g0404(.A(KEYINPUT23), .ZN(new_n605));
  OAI21_X1  g0405(.A(new_n605), .B1(new_n206), .B2(G107), .ZN(new_n606));
  NAND3_X1  g0406(.A1(new_n557), .A2(KEYINPUT23), .A3(G20), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  NAND3_X1  g0408(.A1(new_n206), .A2(G33), .A3(G116), .ZN(new_n609));
  AND2_X1   g0409(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  INV_X1    g0410(.A(KEYINPUT22), .ZN(new_n611));
  AOI21_X1  g0411(.A(new_n611), .B1(new_n525), .B2(G87), .ZN(new_n612));
  OAI211_X1 g0412(.A(new_n206), .B(G87), .C1(new_n364), .C2(new_n365), .ZN(new_n613));
  NOR2_X1   g0413(.A1(new_n613), .A2(KEYINPUT22), .ZN(new_n614));
  OAI211_X1 g0414(.A(KEYINPUT24), .B(new_n610), .C1(new_n612), .C2(new_n614), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n615), .A2(new_n284), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n608), .A2(new_n609), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n613), .A2(KEYINPUT22), .ZN(new_n618));
  NAND4_X1  g0418(.A1(new_n250), .A2(new_n611), .A3(new_n206), .A4(G87), .ZN(new_n619));
  AOI21_X1  g0419(.A(new_n617), .B1(new_n618), .B2(new_n619), .ZN(new_n620));
  NOR2_X1   g0420(.A1(new_n620), .A2(KEYINPUT24), .ZN(new_n621));
  NOR3_X1   g0421(.A1(new_n616), .A2(new_n621), .A3(KEYINPUT86), .ZN(new_n622));
  INV_X1    g0422(.A(KEYINPUT86), .ZN(new_n623));
  AOI21_X1  g0423(.A(new_n423), .B1(new_n620), .B2(KEYINPUT24), .ZN(new_n624));
  OAI21_X1  g0424(.A(new_n610), .B1(new_n612), .B2(new_n614), .ZN(new_n625));
  INV_X1    g0425(.A(KEYINPUT24), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  AOI21_X1  g0427(.A(new_n623), .B1(new_n624), .B2(new_n627), .ZN(new_n628));
  OAI21_X1  g0428(.A(new_n604), .B1(new_n622), .B2(new_n628), .ZN(new_n629));
  OAI211_X1 g0429(.A(G257), .B(G1698), .C1(new_n364), .C2(new_n365), .ZN(new_n630));
  INV_X1    g0430(.A(KEYINPUT87), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n630), .A2(new_n631), .ZN(new_n632));
  NAND4_X1  g0432(.A1(new_n250), .A2(KEYINPUT87), .A3(G257), .A4(G1698), .ZN(new_n633));
  NAND3_X1  g0433(.A1(new_n250), .A2(new_n253), .A3(G250), .ZN(new_n634));
  NAND2_X1  g0434(.A1(G33), .A2(G294), .ZN(new_n635));
  NAND4_X1  g0435(.A1(new_n632), .A2(new_n633), .A3(new_n634), .A4(new_n635), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n636), .A2(new_n258), .ZN(new_n637));
  AND3_X1   g0437(.A1(new_n475), .A2(new_n483), .A3(G264), .ZN(new_n638));
  INV_X1    g0438(.A(new_n638), .ZN(new_n639));
  NAND3_X1  g0439(.A1(new_n637), .A2(new_n485), .A3(new_n639), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n640), .A2(G169), .ZN(new_n641));
  OAI21_X1  g0441(.A(new_n641), .B1(new_n383), .B2(new_n640), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n629), .A2(new_n642), .ZN(new_n643));
  OAI21_X1  g0443(.A(KEYINPUT86), .B1(new_n616), .B2(new_n621), .ZN(new_n644));
  NAND3_X1  g0444(.A1(new_n624), .A2(new_n627), .A3(new_n623), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  NAND4_X1  g0446(.A1(new_n637), .A2(new_n389), .A3(new_n485), .A4(new_n639), .ZN(new_n647));
  INV_X1    g0447(.A(new_n485), .ZN(new_n648));
  AOI211_X1 g0448(.A(new_n648), .B(new_n638), .C1(new_n636), .C2(new_n258), .ZN(new_n649));
  OAI21_X1  g0449(.A(new_n647), .B1(new_n649), .B2(G200), .ZN(new_n650));
  NAND3_X1  g0450(.A1(new_n646), .A2(new_n604), .A3(new_n650), .ZN(new_n651));
  AND2_X1   g0451(.A1(new_n643), .A2(new_n651), .ZN(new_n652));
  AND4_X1   g0452(.A1(new_n458), .A2(new_n509), .A3(new_n600), .A4(new_n652), .ZN(G372));
  NAND4_X1  g0453(.A1(new_n551), .A2(new_n651), .A3(new_n592), .A4(new_n599), .ZN(new_n654));
  INV_X1    g0454(.A(KEYINPUT88), .ZN(new_n655));
  INV_X1    g0455(.A(new_n604), .ZN(new_n656));
  AOI21_X1  g0456(.A(new_n656), .B1(new_n644), .B2(new_n645), .ZN(new_n657));
  AOI21_X1  g0457(.A(new_n638), .B1(new_n636), .B2(new_n258), .ZN(new_n658));
  AND3_X1   g0458(.A1(new_n658), .A2(G179), .A3(new_n485), .ZN(new_n659));
  AOI21_X1  g0459(.A(new_n381), .B1(new_n658), .B2(new_n485), .ZN(new_n660));
  NOR2_X1   g0460(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  OAI21_X1  g0461(.A(new_n655), .B1(new_n657), .B2(new_n661), .ZN(new_n662));
  NAND3_X1  g0462(.A1(new_n629), .A2(new_n642), .A3(KEYINPUT88), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  AND2_X1   g0464(.A1(new_n507), .A2(new_n493), .ZN(new_n665));
  AOI21_X1  g0465(.A(new_n654), .B1(new_n664), .B2(new_n665), .ZN(new_n666));
  AOI21_X1  g0466(.A(new_n511), .B1(new_n523), .B2(new_n530), .ZN(new_n667));
  INV_X1    g0467(.A(new_n513), .ZN(new_n668));
  NAND3_X1  g0468(.A1(new_n667), .A2(new_n541), .A3(new_n668), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n548), .A2(new_n550), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n669), .A2(new_n670), .ZN(new_n671));
  OAI21_X1  g0471(.A(KEYINPUT26), .B1(new_n671), .B2(new_n592), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n591), .A2(new_n587), .ZN(new_n673));
  NOR2_X1   g0473(.A1(new_n673), .A2(new_n593), .ZN(new_n674));
  INV_X1    g0474(.A(KEYINPUT26), .ZN(new_n675));
  NAND3_X1  g0475(.A1(new_n551), .A2(new_n674), .A3(new_n675), .ZN(new_n676));
  NAND3_X1  g0476(.A1(new_n672), .A2(new_n676), .A3(new_n670), .ZN(new_n677));
  OAI21_X1  g0477(.A(new_n458), .B1(new_n666), .B2(new_n677), .ZN(new_n678));
  INV_X1    g0478(.A(new_n305), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n299), .A2(KEYINPUT10), .ZN(new_n680));
  AND2_X1   g0480(.A1(new_n296), .A2(new_n298), .ZN(new_n681));
  NAND4_X1  g0481(.A1(new_n681), .A2(new_n300), .A3(new_n297), .A4(new_n270), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n680), .A2(new_n682), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n338), .A2(new_n320), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n684), .A2(new_n388), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n343), .A2(new_n352), .ZN(new_n686));
  AND4_X1   g0486(.A1(new_n454), .A2(new_n685), .A3(new_n456), .A4(new_n686), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n442), .A2(new_n447), .ZN(new_n688));
  OAI21_X1  g0488(.A(new_n683), .B1(new_n687), .B2(new_n688), .ZN(new_n689));
  NAND3_X1  g0489(.A1(new_n678), .A2(new_n679), .A3(new_n689), .ZN(G369));
  INV_X1    g0490(.A(new_n287), .ZN(new_n691));
  OR3_X1    g0491(.A1(new_n691), .A2(KEYINPUT27), .A3(G20), .ZN(new_n692));
  OAI21_X1  g0492(.A(KEYINPUT27), .B1(new_n691), .B2(G20), .ZN(new_n693));
  NAND3_X1  g0493(.A1(new_n692), .A2(G213), .A3(new_n693), .ZN(new_n694));
  INV_X1    g0494(.A(new_n694), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n695), .A2(G343), .ZN(new_n696));
  INV_X1    g0496(.A(new_n696), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n506), .A2(new_n697), .ZN(new_n698));
  INV_X1    g0498(.A(new_n698), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n665), .A2(new_n699), .ZN(new_n700));
  OAI211_X1 g0500(.A(new_n700), .B(G330), .C1(new_n509), .C2(new_n699), .ZN(new_n701));
  XNOR2_X1  g0501(.A(new_n701), .B(KEYINPUT89), .ZN(new_n702));
  NAND2_X1  g0502(.A1(new_n629), .A2(new_n697), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n652), .A2(new_n703), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n704), .A2(KEYINPUT90), .ZN(new_n705));
  INV_X1    g0505(.A(KEYINPUT90), .ZN(new_n706));
  NAND3_X1  g0506(.A1(new_n652), .A2(new_n706), .A3(new_n703), .ZN(new_n707));
  OAI211_X1 g0507(.A(new_n705), .B(new_n707), .C1(new_n643), .C2(new_n696), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n702), .A2(new_n708), .ZN(new_n709));
  NOR2_X1   g0509(.A1(new_n665), .A2(new_n697), .ZN(new_n710));
  INV_X1    g0510(.A(new_n710), .ZN(new_n711));
  AOI21_X1  g0511(.A(new_n711), .B1(new_n705), .B2(new_n707), .ZN(new_n712));
  NOR2_X1   g0512(.A1(new_n664), .A2(new_n697), .ZN(new_n713));
  NOR2_X1   g0513(.A1(new_n712), .A2(new_n713), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n709), .A2(new_n714), .ZN(G399));
  NAND2_X1  g0515(.A1(new_n209), .A2(new_n479), .ZN(new_n716));
  NOR4_X1   g0516(.A1(G87), .A2(G97), .A3(G107), .A4(G116), .ZN(new_n717));
  NAND3_X1  g0517(.A1(new_n716), .A2(G1), .A3(new_n717), .ZN(new_n718));
  OAI21_X1  g0518(.A(new_n718), .B1(new_n214), .B2(new_n716), .ZN(new_n719));
  XNOR2_X1  g0519(.A(new_n719), .B(KEYINPUT28), .ZN(new_n720));
  INV_X1    g0520(.A(new_n670), .ZN(new_n721));
  NAND2_X1  g0521(.A1(new_n551), .A2(new_n674), .ZN(new_n722));
  AOI21_X1  g0522(.A(new_n721), .B1(new_n722), .B2(KEYINPUT26), .ZN(new_n723));
  OR3_X1    g0523(.A1(new_n671), .A2(new_n592), .A3(KEYINPUT26), .ZN(new_n724));
  AND2_X1   g0524(.A1(new_n665), .A2(new_n643), .ZN(new_n725));
  OAI211_X1 g0525(.A(new_n723), .B(new_n724), .C1(new_n725), .C2(new_n654), .ZN(new_n726));
  AND3_X1   g0526(.A1(new_n726), .A2(KEYINPUT29), .A3(new_n696), .ZN(new_n727));
  OAI21_X1  g0527(.A(new_n696), .B1(new_n666), .B2(new_n677), .ZN(new_n728));
  INV_X1    g0528(.A(KEYINPUT93), .ZN(new_n729));
  NAND2_X1  g0529(.A1(new_n728), .A2(new_n729), .ZN(new_n730));
  OAI211_X1 g0530(.A(KEYINPUT93), .B(new_n696), .C1(new_n666), .C2(new_n677), .ZN(new_n731));
  XOR2_X1   g0531(.A(KEYINPUT94), .B(KEYINPUT29), .Z(new_n732));
  NAND3_X1  g0532(.A1(new_n730), .A2(new_n731), .A3(new_n732), .ZN(new_n733));
  INV_X1    g0533(.A(KEYINPUT95), .ZN(new_n734));
  NAND2_X1  g0534(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  NAND4_X1  g0535(.A1(new_n730), .A2(KEYINPUT95), .A3(new_n731), .A4(new_n732), .ZN(new_n736));
  AOI21_X1  g0536(.A(new_n727), .B1(new_n735), .B2(new_n736), .ZN(new_n737));
  NAND4_X1  g0537(.A1(new_n509), .A2(new_n600), .A3(new_n652), .A4(new_n696), .ZN(new_n738));
  INV_X1    g0538(.A(KEYINPUT91), .ZN(new_n739));
  AOI21_X1  g0539(.A(new_n739), .B1(new_n658), .B2(new_n539), .ZN(new_n740));
  INV_X1    g0540(.A(new_n740), .ZN(new_n741));
  NOR2_X1   g0541(.A1(new_n596), .A2(new_n504), .ZN(new_n742));
  NAND4_X1  g0542(.A1(new_n637), .A2(new_n539), .A3(new_n739), .A4(new_n639), .ZN(new_n743));
  NAND4_X1  g0543(.A1(new_n741), .A2(new_n742), .A3(KEYINPUT30), .A4(new_n743), .ZN(new_n744));
  AND2_X1   g0544(.A1(new_n538), .A2(new_n258), .ZN(new_n745));
  OAI211_X1 g0545(.A(new_n491), .B(new_n383), .C1(new_n745), .C2(new_n534), .ZN(new_n746));
  OR3_X1    g0546(.A1(new_n746), .A2(new_n649), .A3(new_n586), .ZN(new_n747));
  INV_X1    g0547(.A(KEYINPUT30), .ZN(new_n748));
  AND3_X1   g0548(.A1(new_n486), .A2(new_n490), .A3(G179), .ZN(new_n749));
  NAND3_X1  g0549(.A1(new_n743), .A2(new_n749), .A3(new_n586), .ZN(new_n750));
  OAI21_X1  g0550(.A(new_n748), .B1(new_n750), .B2(new_n740), .ZN(new_n751));
  NAND3_X1  g0551(.A1(new_n744), .A2(new_n747), .A3(new_n751), .ZN(new_n752));
  NAND2_X1  g0552(.A1(new_n752), .A2(new_n697), .ZN(new_n753));
  INV_X1    g0553(.A(KEYINPUT31), .ZN(new_n754));
  NAND2_X1  g0554(.A1(new_n753), .A2(new_n754), .ZN(new_n755));
  NOR3_X1   g0555(.A1(new_n746), .A2(new_n649), .A3(new_n586), .ZN(new_n756));
  NOR2_X1   g0556(.A1(new_n750), .A2(new_n740), .ZN(new_n757));
  AOI21_X1  g0557(.A(new_n756), .B1(new_n757), .B2(KEYINPUT30), .ZN(new_n758));
  AOI21_X1  g0558(.A(new_n696), .B1(new_n758), .B2(new_n751), .ZN(new_n759));
  NAND2_X1  g0559(.A1(new_n759), .A2(KEYINPUT31), .ZN(new_n760));
  NAND3_X1  g0560(.A1(new_n738), .A2(new_n755), .A3(new_n760), .ZN(new_n761));
  AND3_X1   g0561(.A1(new_n761), .A2(KEYINPUT92), .A3(G330), .ZN(new_n762));
  AOI21_X1  g0562(.A(KEYINPUT92), .B1(new_n761), .B2(G330), .ZN(new_n763));
  OR2_X1    g0563(.A1(new_n762), .A2(new_n763), .ZN(new_n764));
  NOR2_X1   g0564(.A1(new_n737), .A2(new_n764), .ZN(new_n765));
  OAI21_X1  g0565(.A(new_n720), .B1(new_n765), .B2(G1), .ZN(G364));
  NAND3_X1  g0566(.A1(new_n209), .A2(G355), .A3(new_n250), .ZN(new_n767));
  INV_X1    g0567(.A(new_n209), .ZN(new_n768));
  NOR2_X1   g0568(.A1(new_n768), .A2(new_n250), .ZN(new_n769));
  INV_X1    g0569(.A(new_n769), .ZN(new_n770));
  NOR2_X1   g0570(.A1(new_n215), .A2(G45), .ZN(new_n771));
  AOI21_X1  g0571(.A(new_n771), .B1(new_n243), .B2(G45), .ZN(new_n772));
  OAI221_X1 g0572(.A(new_n767), .B1(G116), .B2(new_n209), .C1(new_n770), .C2(new_n772), .ZN(new_n773));
  NOR2_X1   g0573(.A1(G13), .A2(G33), .ZN(new_n774));
  NAND2_X1  g0574(.A1(new_n774), .A2(new_n206), .ZN(new_n775));
  XOR2_X1   g0575(.A(new_n775), .B(KEYINPUT97), .Z(new_n776));
  AOI21_X1  g0576(.A(new_n212), .B1(G20), .B2(new_n381), .ZN(new_n777));
  INV_X1    g0577(.A(new_n777), .ZN(new_n778));
  NAND2_X1  g0578(.A1(new_n776), .A2(new_n778), .ZN(new_n779));
  XOR2_X1   g0579(.A(new_n779), .B(KEYINPUT98), .Z(new_n780));
  INV_X1    g0580(.A(new_n780), .ZN(new_n781));
  NAND2_X1  g0581(.A1(new_n773), .A2(new_n781), .ZN(new_n782));
  OR3_X1    g0582(.A1(new_n206), .A2(KEYINPUT100), .A3(G190), .ZN(new_n783));
  OAI21_X1  g0583(.A(KEYINPUT100), .B1(new_n206), .B2(G190), .ZN(new_n784));
  NOR2_X1   g0584(.A1(G179), .A2(G200), .ZN(new_n785));
  NAND3_X1  g0585(.A1(new_n783), .A2(new_n784), .A3(new_n785), .ZN(new_n786));
  INV_X1    g0586(.A(new_n786), .ZN(new_n787));
  NAND2_X1  g0587(.A1(new_n787), .A2(G159), .ZN(new_n788));
  XNOR2_X1  g0588(.A(new_n788), .B(KEYINPUT101), .ZN(new_n789));
  XNOR2_X1  g0589(.A(new_n789), .B(KEYINPUT32), .ZN(new_n790));
  NOR2_X1   g0590(.A1(new_n391), .A2(G179), .ZN(new_n791));
  NAND3_X1  g0591(.A1(new_n783), .A2(new_n791), .A3(new_n784), .ZN(new_n792));
  NOR2_X1   g0592(.A1(new_n792), .A2(new_n557), .ZN(new_n793));
  AOI21_X1  g0593(.A(new_n206), .B1(new_n785), .B2(G190), .ZN(new_n794));
  NOR2_X1   g0594(.A1(new_n794), .A2(new_n221), .ZN(new_n795));
  NOR2_X1   g0595(.A1(new_n383), .A2(new_n391), .ZN(new_n796));
  NOR2_X1   g0596(.A1(new_n206), .A2(G190), .ZN(new_n797));
  NAND2_X1  g0597(.A1(new_n796), .A2(new_n797), .ZN(new_n798));
  INV_X1    g0598(.A(new_n798), .ZN(new_n799));
  AOI211_X1 g0599(.A(new_n400), .B(new_n795), .C1(G68), .C2(new_n799), .ZN(new_n800));
  NOR2_X1   g0600(.A1(new_n206), .A2(new_n389), .ZN(new_n801));
  NAND2_X1  g0601(.A1(new_n801), .A2(new_n791), .ZN(new_n802));
  INV_X1    g0602(.A(new_n802), .ZN(new_n803));
  NOR2_X1   g0603(.A1(new_n383), .A2(G200), .ZN(new_n804));
  NAND2_X1  g0604(.A1(new_n804), .A2(new_n797), .ZN(new_n805));
  INV_X1    g0605(.A(new_n805), .ZN(new_n806));
  AOI22_X1  g0606(.A1(G87), .A2(new_n803), .B1(new_n806), .B2(G77), .ZN(new_n807));
  NAND2_X1  g0607(.A1(new_n801), .A2(new_n796), .ZN(new_n808));
  OAI211_X1 g0608(.A(new_n800), .B(new_n807), .C1(new_n285), .C2(new_n808), .ZN(new_n809));
  AND3_X1   g0609(.A1(new_n801), .A2(KEYINPUT99), .A3(new_n804), .ZN(new_n810));
  AOI21_X1  g0610(.A(KEYINPUT99), .B1(new_n801), .B2(new_n804), .ZN(new_n811));
  NOR2_X1   g0611(.A1(new_n810), .A2(new_n811), .ZN(new_n812));
  INV_X1    g0612(.A(new_n812), .ZN(new_n813));
  AOI211_X1 g0613(.A(new_n793), .B(new_n809), .C1(G58), .C2(new_n813), .ZN(new_n814));
  INV_X1    g0614(.A(G283), .ZN(new_n815));
  INV_X1    g0615(.A(G329), .ZN(new_n816));
  OAI22_X1  g0616(.A1(new_n815), .A2(new_n792), .B1(new_n786), .B2(new_n816), .ZN(new_n817));
  AOI21_X1  g0617(.A(new_n250), .B1(new_n806), .B2(G311), .ZN(new_n818));
  INV_X1    g0618(.A(G303), .ZN(new_n819));
  XOR2_X1   g0619(.A(KEYINPUT33), .B(G317), .Z(new_n820));
  OAI221_X1 g0620(.A(new_n818), .B1(new_n819), .B2(new_n802), .C1(new_n798), .C2(new_n820), .ZN(new_n821));
  AOI211_X1 g0621(.A(new_n817), .B(new_n821), .C1(G322), .C2(new_n813), .ZN(new_n822));
  INV_X1    g0622(.A(G326), .ZN(new_n823));
  INV_X1    g0623(.A(G294), .ZN(new_n824));
  OAI22_X1  g0624(.A1(new_n808), .A2(new_n823), .B1(new_n794), .B2(new_n824), .ZN(new_n825));
  XNOR2_X1  g0625(.A(new_n825), .B(KEYINPUT102), .ZN(new_n826));
  AOI22_X1  g0626(.A1(new_n790), .A2(new_n814), .B1(new_n822), .B2(new_n826), .ZN(new_n827));
  OAI21_X1  g0627(.A(new_n782), .B1(new_n827), .B2(new_n778), .ZN(new_n828));
  OAI21_X1  g0628(.A(new_n700), .B1(new_n509), .B2(new_n699), .ZN(new_n829));
  INV_X1    g0629(.A(new_n776), .ZN(new_n830));
  AOI21_X1  g0630(.A(new_n828), .B1(new_n829), .B2(new_n830), .ZN(new_n831));
  INV_X1    g0631(.A(G330), .ZN(new_n832));
  AND2_X1   g0632(.A1(new_n829), .A2(new_n832), .ZN(new_n833));
  NOR2_X1   g0633(.A1(new_n702), .A2(new_n833), .ZN(new_n834));
  NAND2_X1  g0634(.A1(new_n206), .A2(G13), .ZN(new_n835));
  NOR2_X1   g0635(.A1(new_n835), .A2(new_n481), .ZN(new_n836));
  XNOR2_X1  g0636(.A(new_n836), .B(KEYINPUT96), .ZN(new_n837));
  NAND3_X1  g0637(.A1(new_n716), .A2(G1), .A3(new_n837), .ZN(new_n838));
  MUX2_X1   g0638(.A(new_n831), .B(new_n834), .S(new_n838), .Z(G396));
  INV_X1    g0639(.A(new_n838), .ZN(new_n840));
  NOR2_X1   g0640(.A1(new_n777), .A2(new_n774), .ZN(new_n841));
  INV_X1    g0641(.A(new_n841), .ZN(new_n842));
  OAI22_X1  g0642(.A1(new_n808), .A2(new_n819), .B1(new_n805), .B2(new_n463), .ZN(new_n843));
  AOI21_X1  g0643(.A(new_n843), .B1(G283), .B2(new_n799), .ZN(new_n844));
  XNOR2_X1  g0644(.A(new_n844), .B(KEYINPUT103), .ZN(new_n845));
  AOI211_X1 g0645(.A(new_n250), .B(new_n795), .C1(G107), .C2(new_n803), .ZN(new_n846));
  OAI21_X1  g0646(.A(new_n846), .B1(new_n824), .B2(new_n812), .ZN(new_n847));
  INV_X1    g0647(.A(G311), .ZN(new_n848));
  OAI22_X1  g0648(.A1(new_n434), .A2(new_n792), .B1(new_n786), .B2(new_n848), .ZN(new_n849));
  NOR3_X1   g0649(.A1(new_n845), .A2(new_n847), .A3(new_n849), .ZN(new_n850));
  OAI22_X1  g0650(.A1(new_n802), .A2(new_n285), .B1(new_n794), .B2(new_n219), .ZN(new_n851));
  AOI21_X1  g0651(.A(new_n400), .B1(new_n787), .B2(G132), .ZN(new_n852));
  XOR2_X1   g0652(.A(new_n852), .B(KEYINPUT105), .Z(new_n853));
  INV_X1    g0653(.A(new_n792), .ZN(new_n854));
  AOI211_X1 g0654(.A(new_n851), .B(new_n853), .C1(G68), .C2(new_n854), .ZN(new_n855));
  INV_X1    g0655(.A(G137), .ZN(new_n856));
  OAI22_X1  g0656(.A1(new_n808), .A2(new_n856), .B1(new_n798), .B2(new_n271), .ZN(new_n857));
  XNOR2_X1  g0657(.A(new_n857), .B(KEYINPUT104), .ZN(new_n858));
  INV_X1    g0658(.A(G143), .ZN(new_n859));
  INV_X1    g0659(.A(G159), .ZN(new_n860));
  OAI221_X1 g0660(.A(new_n858), .B1(new_n859), .B2(new_n812), .C1(new_n860), .C2(new_n805), .ZN(new_n861));
  XNOR2_X1  g0661(.A(new_n861), .B(KEYINPUT34), .ZN(new_n862));
  AOI21_X1  g0662(.A(new_n850), .B1(new_n855), .B2(new_n862), .ZN(new_n863));
  OAI221_X1 g0663(.A(new_n840), .B1(G77), .B2(new_n842), .C1(new_n863), .C2(new_n778), .ZN(new_n864));
  XOR2_X1   g0664(.A(new_n864), .B(KEYINPUT106), .Z(new_n865));
  INV_X1    g0665(.A(new_n774), .ZN(new_n866));
  INV_X1    g0666(.A(new_n388), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n867), .A2(new_n697), .ZN(new_n868));
  NOR2_X1   g0668(.A1(new_n362), .A2(new_n696), .ZN(new_n869));
  INV_X1    g0669(.A(new_n869), .ZN(new_n870));
  AND4_X1   g0670(.A1(KEYINPUT107), .A2(new_n394), .A3(new_n388), .A4(new_n870), .ZN(new_n871));
  AOI21_X1  g0671(.A(new_n869), .B1(new_n393), .B2(new_n362), .ZN(new_n872));
  AOI21_X1  g0672(.A(KEYINPUT107), .B1(new_n872), .B2(new_n388), .ZN(new_n873));
  OAI21_X1  g0673(.A(new_n868), .B1(new_n871), .B2(new_n873), .ZN(new_n874));
  OAI21_X1  g0674(.A(new_n865), .B1(new_n866), .B2(new_n874), .ZN(new_n875));
  INV_X1    g0675(.A(new_n875), .ZN(new_n876));
  NAND3_X1  g0676(.A1(new_n394), .A2(new_n388), .A3(new_n870), .ZN(new_n877));
  INV_X1    g0677(.A(KEYINPUT107), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n877), .A2(new_n878), .ZN(new_n879));
  NAND3_X1  g0679(.A1(new_n872), .A2(KEYINPUT107), .A3(new_n388), .ZN(new_n880));
  AOI22_X1  g0680(.A1(new_n879), .A2(new_n880), .B1(new_n867), .B2(new_n697), .ZN(new_n881));
  NAND3_X1  g0681(.A1(new_n730), .A2(new_n731), .A3(new_n881), .ZN(new_n882));
  OAI21_X1  g0682(.A(new_n882), .B1(new_n728), .B2(new_n881), .ZN(new_n883));
  INV_X1    g0683(.A(new_n883), .ZN(new_n884));
  NOR2_X1   g0684(.A1(new_n884), .A2(new_n764), .ZN(new_n885));
  INV_X1    g0685(.A(new_n885), .ZN(new_n886));
  AOI21_X1  g0686(.A(new_n840), .B1(new_n884), .B2(new_n764), .ZN(new_n887));
  AOI21_X1  g0687(.A(new_n876), .B1(new_n886), .B2(new_n887), .ZN(new_n888));
  INV_X1    g0688(.A(new_n888), .ZN(G384));
  NAND2_X1  g0689(.A1(new_n560), .A2(new_n565), .ZN(new_n890));
  OAI211_X1 g0690(.A(G116), .B(new_n213), .C1(new_n890), .C2(KEYINPUT35), .ZN(new_n891));
  AOI21_X1  g0691(.A(new_n891), .B1(KEYINPUT35), .B2(new_n890), .ZN(new_n892));
  OAI21_X1  g0692(.A(G77), .B1(new_n219), .B2(new_n308), .ZN(new_n893));
  OAI22_X1  g0693(.A1(new_n893), .A2(new_n214), .B1(G50), .B2(new_n308), .ZN(new_n894));
  NOR2_X1   g0694(.A1(new_n205), .A2(G13), .ZN(new_n895));
  AOI22_X1  g0695(.A1(new_n892), .A2(KEYINPUT36), .B1(new_n894), .B2(new_n895), .ZN(new_n896));
  INV_X1    g0696(.A(KEYINPUT111), .ZN(new_n897));
  OAI21_X1  g0697(.A(new_n897), .B1(new_n759), .B2(KEYINPUT31), .ZN(new_n898));
  NAND3_X1  g0698(.A1(new_n753), .A2(KEYINPUT111), .A3(new_n754), .ZN(new_n899));
  NAND4_X1  g0699(.A1(new_n898), .A2(new_n738), .A3(new_n760), .A4(new_n899), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n332), .A2(new_n337), .ZN(new_n901));
  AOI21_X1  g0701(.A(new_n331), .B1(new_n350), .B2(G169), .ZN(new_n902));
  OAI211_X1 g0702(.A(new_n320), .B(new_n697), .C1(new_n901), .C2(new_n902), .ZN(new_n903));
  INV_X1    g0703(.A(new_n903), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n320), .A2(new_n697), .ZN(new_n905));
  AOI21_X1  g0705(.A(new_n904), .B1(new_n353), .B2(new_n905), .ZN(new_n906));
  INV_X1    g0706(.A(new_n906), .ZN(new_n907));
  AND4_X1   g0707(.A1(KEYINPUT40), .A2(new_n900), .A3(new_n874), .A4(new_n907), .ZN(new_n908));
  XOR2_X1   g0708(.A(KEYINPUT109), .B(KEYINPUT38), .Z(new_n909));
  AND3_X1   g0709(.A1(new_n457), .A2(new_n445), .A3(new_n695), .ZN(new_n910));
  OAI21_X1  g0710(.A(new_n694), .B1(new_n438), .B2(new_n439), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n445), .A2(new_n911), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n912), .A2(new_n452), .ZN(new_n913));
  AOI21_X1  g0713(.A(KEYINPUT110), .B1(new_n445), .B2(new_n911), .ZN(new_n914));
  INV_X1    g0714(.A(KEYINPUT37), .ZN(new_n915));
  OAI21_X1  g0715(.A(new_n913), .B1(new_n914), .B2(new_n915), .ZN(new_n916));
  NAND4_X1  g0716(.A1(new_n912), .A2(KEYINPUT110), .A3(KEYINPUT37), .A4(new_n452), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n916), .A2(new_n917), .ZN(new_n918));
  OAI21_X1  g0718(.A(new_n909), .B1(new_n910), .B2(new_n918), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n429), .A2(new_n284), .ZN(new_n920));
  AOI21_X1  g0720(.A(new_n409), .B1(new_n419), .B2(KEYINPUT77), .ZN(new_n921));
  AOI21_X1  g0721(.A(KEYINPUT16), .B1(new_n921), .B2(new_n428), .ZN(new_n922));
  OAI21_X1  g0722(.A(new_n397), .B1(new_n920), .B2(new_n922), .ZN(new_n923));
  AND2_X1   g0723(.A1(new_n923), .A2(new_n695), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n454), .A2(new_n456), .ZN(new_n925));
  OAI21_X1  g0725(.A(new_n924), .B1(new_n688), .B2(new_n925), .ZN(new_n926));
  NAND2_X1  g0726(.A1(new_n923), .A2(new_n911), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n452), .A2(new_n927), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n928), .A2(KEYINPUT37), .ZN(new_n929));
  INV_X1    g0729(.A(new_n911), .ZN(new_n930));
  OAI211_X1 g0730(.A(new_n452), .B(new_n915), .C1(new_n431), .C2(new_n930), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n929), .A2(new_n931), .ZN(new_n932));
  NAND3_X1  g0732(.A1(new_n926), .A2(KEYINPUT38), .A3(new_n932), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n919), .A2(new_n933), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n908), .A2(new_n934), .ZN(new_n935));
  INV_X1    g0735(.A(KEYINPUT40), .ZN(new_n936));
  INV_X1    g0736(.A(KEYINPUT38), .ZN(new_n937));
  AOI221_X4 g0737(.A(new_n937), .B1(new_n929), .B2(new_n931), .C1(new_n457), .C2(new_n924), .ZN(new_n938));
  AOI21_X1  g0738(.A(KEYINPUT38), .B1(new_n926), .B2(new_n932), .ZN(new_n939));
  NOR2_X1   g0739(.A1(new_n938), .A2(new_n939), .ZN(new_n940));
  NAND3_X1  g0740(.A1(new_n900), .A2(new_n874), .A3(new_n907), .ZN(new_n941));
  OAI21_X1  g0741(.A(new_n936), .B1(new_n940), .B2(new_n941), .ZN(new_n942));
  NAND3_X1  g0742(.A1(new_n935), .A2(new_n942), .A3(G330), .ZN(new_n943));
  AND3_X1   g0743(.A1(new_n458), .A2(G330), .A3(new_n900), .ZN(new_n944));
  INV_X1    g0744(.A(new_n944), .ZN(new_n945));
  AOI21_X1  g0745(.A(KEYINPUT112), .B1(new_n943), .B2(new_n945), .ZN(new_n946));
  AND3_X1   g0746(.A1(new_n943), .A2(KEYINPUT112), .A3(new_n945), .ZN(new_n947));
  AND2_X1   g0747(.A1(new_n458), .A2(new_n900), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n879), .A2(new_n880), .ZN(new_n949));
  AOI21_X1  g0749(.A(new_n906), .B1(new_n949), .B2(new_n868), .ZN(new_n950));
  OAI211_X1 g0750(.A(new_n950), .B(new_n900), .C1(new_n938), .C2(new_n939), .ZN(new_n951));
  AOI22_X1  g0751(.A1(new_n936), .A2(new_n951), .B1(new_n908), .B2(new_n934), .ZN(new_n952));
  AOI211_X1 g0752(.A(new_n946), .B(new_n947), .C1(new_n948), .C2(new_n952), .ZN(new_n953));
  NAND2_X1  g0753(.A1(new_n688), .A2(new_n694), .ZN(new_n954));
  NOR2_X1   g0754(.A1(new_n388), .A2(new_n697), .ZN(new_n955));
  INV_X1    g0755(.A(new_n955), .ZN(new_n956));
  OAI21_X1  g0756(.A(new_n956), .B1(new_n881), .B2(new_n728), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n957), .A2(new_n907), .ZN(new_n958));
  OAI21_X1  g0758(.A(new_n954), .B1(new_n958), .B2(new_n940), .ZN(new_n959));
  OAI21_X1  g0759(.A(KEYINPUT39), .B1(new_n938), .B2(new_n939), .ZN(new_n960));
  NAND2_X1  g0760(.A1(new_n960), .A2(KEYINPUT108), .ZN(new_n961));
  INV_X1    g0761(.A(KEYINPUT108), .ZN(new_n962));
  OAI211_X1 g0762(.A(new_n962), .B(KEYINPUT39), .C1(new_n938), .C2(new_n939), .ZN(new_n963));
  INV_X1    g0763(.A(KEYINPUT39), .ZN(new_n964));
  NAND3_X1  g0764(.A1(new_n919), .A2(new_n964), .A3(new_n933), .ZN(new_n965));
  NAND3_X1  g0765(.A1(new_n961), .A2(new_n963), .A3(new_n965), .ZN(new_n966));
  NAND3_X1  g0766(.A1(new_n338), .A2(new_n320), .A3(new_n696), .ZN(new_n967));
  INV_X1    g0767(.A(new_n967), .ZN(new_n968));
  AOI21_X1  g0768(.A(new_n959), .B1(new_n966), .B2(new_n968), .ZN(new_n969));
  NAND2_X1  g0769(.A1(new_n689), .A2(new_n679), .ZN(new_n970));
  AOI21_X1  g0770(.A(new_n970), .B1(new_n737), .B2(new_n458), .ZN(new_n971));
  XOR2_X1   g0771(.A(new_n969), .B(new_n971), .Z(new_n972));
  AOI22_X1  g0772(.A1(new_n953), .A2(new_n972), .B1(G1), .B2(new_n835), .ZN(new_n973));
  INV_X1    g0773(.A(KEYINPUT113), .ZN(new_n974));
  OAI22_X1  g0774(.A1(new_n973), .A2(new_n974), .B1(new_n953), .B2(new_n972), .ZN(new_n975));
  AND2_X1   g0775(.A1(new_n973), .A2(new_n974), .ZN(new_n976));
  OAI221_X1 g0776(.A(new_n896), .B1(KEYINPUT36), .B2(new_n892), .C1(new_n975), .C2(new_n976), .ZN(new_n977));
  XOR2_X1   g0777(.A(new_n977), .B(KEYINPUT114), .Z(G367));
  AOI22_X1  g0778(.A1(new_n769), .A2(new_n239), .B1(new_n768), .B2(new_n510), .ZN(new_n979));
  AOI21_X1  g0779(.A(new_n838), .B1(new_n781), .B2(new_n979), .ZN(new_n980));
  NOR2_X1   g0780(.A1(new_n802), .A2(new_n463), .ZN(new_n981));
  XNOR2_X1  g0781(.A(new_n981), .B(KEYINPUT46), .ZN(new_n982));
  INV_X1    g0782(.A(new_n794), .ZN(new_n983));
  AOI21_X1  g0783(.A(new_n982), .B1(G107), .B2(new_n983), .ZN(new_n984));
  NAND2_X1  g0784(.A1(new_n813), .A2(G303), .ZN(new_n985));
  OAI22_X1  g0785(.A1(new_n808), .A2(new_n848), .B1(new_n798), .B2(new_n824), .ZN(new_n986));
  AOI211_X1 g0786(.A(new_n250), .B(new_n986), .C1(G283), .C2(new_n806), .ZN(new_n987));
  AOI22_X1  g0787(.A1(G97), .A2(new_n854), .B1(new_n787), .B2(G317), .ZN(new_n988));
  NAND4_X1  g0788(.A1(new_n984), .A2(new_n985), .A3(new_n987), .A4(new_n988), .ZN(new_n989));
  NOR2_X1   g0789(.A1(new_n794), .A2(new_n308), .ZN(new_n990));
  INV_X1    g0790(.A(new_n808), .ZN(new_n991));
  AOI211_X1 g0791(.A(new_n400), .B(new_n990), .C1(G143), .C2(new_n991), .ZN(new_n992));
  AOI22_X1  g0792(.A1(G77), .A2(new_n854), .B1(new_n787), .B2(G137), .ZN(new_n993));
  NAND2_X1  g0793(.A1(new_n813), .A2(G150), .ZN(new_n994));
  OAI22_X1  g0794(.A1(new_n219), .A2(new_n802), .B1(new_n798), .B2(new_n860), .ZN(new_n995));
  AOI21_X1  g0795(.A(new_n995), .B1(G50), .B2(new_n806), .ZN(new_n996));
  NAND4_X1  g0796(.A1(new_n992), .A2(new_n993), .A3(new_n994), .A4(new_n996), .ZN(new_n997));
  NAND3_X1  g0797(.A1(new_n989), .A2(KEYINPUT47), .A3(new_n997), .ZN(new_n998));
  NAND2_X1  g0798(.A1(new_n998), .A2(new_n777), .ZN(new_n999));
  AOI21_X1  g0799(.A(KEYINPUT47), .B1(new_n989), .B2(new_n997), .ZN(new_n1000));
  OAI21_X1  g0800(.A(new_n980), .B1(new_n999), .B2(new_n1000), .ZN(new_n1001));
  XNOR2_X1  g0801(.A(new_n1001), .B(KEYINPUT118), .ZN(new_n1002));
  NOR2_X1   g0802(.A1(new_n531), .A2(new_n696), .ZN(new_n1003));
  XOR2_X1   g0803(.A(new_n1003), .B(KEYINPUT115), .Z(new_n1004));
  OR2_X1    g0804(.A1(new_n1004), .A2(new_n721), .ZN(new_n1005));
  NAND2_X1  g0805(.A1(new_n1004), .A2(new_n671), .ZN(new_n1006));
  NAND2_X1  g0806(.A1(new_n1005), .A2(new_n1006), .ZN(new_n1007));
  AOI21_X1  g0807(.A(new_n1002), .B1(new_n1007), .B2(new_n830), .ZN(new_n1008));
  XNOR2_X1  g0808(.A(new_n1008), .B(KEYINPUT119), .ZN(new_n1009));
  NAND2_X1  g0809(.A1(new_n837), .A2(G1), .ZN(new_n1010));
  NAND2_X1  g0810(.A1(new_n705), .A2(new_n707), .ZN(new_n1011));
  NAND2_X1  g0811(.A1(new_n1011), .A2(new_n710), .ZN(new_n1012));
  OAI21_X1  g0812(.A(new_n1012), .B1(new_n708), .B2(new_n710), .ZN(new_n1013));
  XNOR2_X1  g0813(.A(new_n1013), .B(new_n702), .ZN(new_n1014));
  AND2_X1   g0814(.A1(new_n765), .A2(new_n1014), .ZN(new_n1015));
  AOI21_X1  g0815(.A(KEYINPUT117), .B1(new_n702), .B2(new_n708), .ZN(new_n1016));
  OR2_X1    g0816(.A1(new_n712), .A2(new_n713), .ZN(new_n1017));
  INV_X1    g0817(.A(KEYINPUT44), .ZN(new_n1018));
  OAI211_X1 g0818(.A(new_n592), .B(new_n599), .C1(new_n593), .C2(new_n696), .ZN(new_n1019));
  NAND2_X1  g0819(.A1(new_n674), .A2(new_n697), .ZN(new_n1020));
  AND2_X1   g0820(.A1(new_n1019), .A2(new_n1020), .ZN(new_n1021));
  NAND3_X1  g0821(.A1(new_n1017), .A2(new_n1018), .A3(new_n1021), .ZN(new_n1022));
  OAI21_X1  g0822(.A(new_n1021), .B1(new_n712), .B2(new_n713), .ZN(new_n1023));
  NAND2_X1  g0823(.A1(new_n1023), .A2(KEYINPUT44), .ZN(new_n1024));
  NAND3_X1  g0824(.A1(new_n702), .A2(KEYINPUT117), .A3(new_n708), .ZN(new_n1025));
  NAND3_X1  g0825(.A1(new_n1022), .A2(new_n1024), .A3(new_n1025), .ZN(new_n1026));
  INV_X1    g0826(.A(new_n1021), .ZN(new_n1027));
  AOI21_X1  g0827(.A(KEYINPUT45), .B1(new_n714), .B2(new_n1027), .ZN(new_n1028));
  INV_X1    g0828(.A(KEYINPUT45), .ZN(new_n1029));
  NOR4_X1   g0829(.A1(new_n712), .A2(new_n1029), .A3(new_n713), .A4(new_n1021), .ZN(new_n1030));
  NOR2_X1   g0830(.A1(new_n1028), .A2(new_n1030), .ZN(new_n1031));
  OAI21_X1  g0831(.A(new_n1016), .B1(new_n1026), .B2(new_n1031), .ZN(new_n1032));
  OAI21_X1  g0832(.A(new_n1029), .B1(new_n1017), .B2(new_n1021), .ZN(new_n1033));
  INV_X1    g0833(.A(new_n1030), .ZN(new_n1034));
  NAND2_X1  g0834(.A1(new_n1033), .A2(new_n1034), .ZN(new_n1035));
  XNOR2_X1  g0835(.A(new_n1023), .B(new_n1018), .ZN(new_n1036));
  INV_X1    g0836(.A(new_n1016), .ZN(new_n1037));
  NAND4_X1  g0837(.A1(new_n1035), .A2(new_n1036), .A3(new_n1025), .A4(new_n1037), .ZN(new_n1038));
  NAND2_X1  g0838(.A1(new_n1032), .A2(new_n1038), .ZN(new_n1039));
  NAND2_X1  g0839(.A1(new_n1015), .A2(new_n1039), .ZN(new_n1040));
  NAND2_X1  g0840(.A1(new_n1040), .A2(new_n765), .ZN(new_n1041));
  XNOR2_X1  g0841(.A(new_n716), .B(KEYINPUT41), .ZN(new_n1042));
  INV_X1    g0842(.A(new_n1042), .ZN(new_n1043));
  AOI21_X1  g0843(.A(new_n1010), .B1(new_n1041), .B2(new_n1043), .ZN(new_n1044));
  NOR2_X1   g0844(.A1(new_n1012), .A2(new_n1021), .ZN(new_n1045));
  INV_X1    g0845(.A(KEYINPUT42), .ZN(new_n1046));
  NAND2_X1  g0846(.A1(new_n1045), .A2(new_n1046), .ZN(new_n1047));
  OAI21_X1  g0847(.A(new_n592), .B1(new_n1021), .B2(new_n643), .ZN(new_n1048));
  NAND2_X1  g0848(.A1(new_n1048), .A2(new_n696), .ZN(new_n1049));
  AND2_X1   g0849(.A1(new_n1047), .A2(new_n1049), .ZN(new_n1050));
  INV_X1    g0850(.A(KEYINPUT43), .ZN(new_n1051));
  NOR2_X1   g0851(.A1(new_n1045), .A2(new_n1046), .ZN(new_n1052));
  INV_X1    g0852(.A(new_n1052), .ZN(new_n1053));
  NAND4_X1  g0853(.A1(new_n1050), .A2(new_n1051), .A3(new_n1007), .A4(new_n1053), .ZN(new_n1054));
  NAND3_X1  g0854(.A1(new_n702), .A2(new_n708), .A3(new_n1027), .ZN(new_n1055));
  INV_X1    g0855(.A(new_n1055), .ZN(new_n1056));
  NAND2_X1  g0856(.A1(new_n1007), .A2(new_n1051), .ZN(new_n1057));
  INV_X1    g0857(.A(new_n1007), .ZN(new_n1058));
  NAND2_X1  g0858(.A1(new_n1058), .A2(KEYINPUT43), .ZN(new_n1059));
  NAND2_X1  g0859(.A1(new_n1047), .A2(new_n1049), .ZN(new_n1060));
  OAI211_X1 g0860(.A(new_n1057), .B(new_n1059), .C1(new_n1060), .C2(new_n1052), .ZN(new_n1061));
  NAND3_X1  g0861(.A1(new_n1054), .A2(new_n1056), .A3(new_n1061), .ZN(new_n1062));
  INV_X1    g0862(.A(KEYINPUT116), .ZN(new_n1063));
  NAND2_X1  g0863(.A1(new_n1062), .A2(new_n1063), .ZN(new_n1064));
  NAND4_X1  g0864(.A1(new_n1054), .A2(new_n1061), .A3(KEYINPUT116), .A4(new_n1056), .ZN(new_n1065));
  NAND2_X1  g0865(.A1(new_n1054), .A2(new_n1061), .ZN(new_n1066));
  NAND2_X1  g0866(.A1(new_n1066), .A2(new_n1055), .ZN(new_n1067));
  NAND3_X1  g0867(.A1(new_n1064), .A2(new_n1065), .A3(new_n1067), .ZN(new_n1068));
  OAI21_X1  g0868(.A(new_n1009), .B1(new_n1044), .B2(new_n1068), .ZN(G387));
  OR2_X1    g0869(.A1(new_n708), .A2(new_n776), .ZN(new_n1070));
  NAND3_X1  g0870(.A1(new_n236), .A2(G45), .A3(new_n400), .ZN(new_n1071));
  OAI21_X1  g0871(.A(new_n481), .B1(new_n308), .B2(new_n202), .ZN(new_n1072));
  INV_X1    g0872(.A(new_n275), .ZN(new_n1073));
  NAND3_X1  g0873(.A1(new_n1073), .A2(KEYINPUT50), .A3(new_n285), .ZN(new_n1074));
  INV_X1    g0874(.A(KEYINPUT50), .ZN(new_n1075));
  OAI21_X1  g0875(.A(new_n1075), .B1(new_n275), .B2(G50), .ZN(new_n1076));
  AOI21_X1  g0876(.A(new_n1072), .B1(new_n1074), .B2(new_n1076), .ZN(new_n1077));
  OAI21_X1  g0877(.A(new_n717), .B1(new_n1077), .B2(new_n250), .ZN(new_n1078));
  AOI21_X1  g0878(.A(new_n768), .B1(new_n1071), .B2(new_n1078), .ZN(new_n1079));
  OAI21_X1  g0879(.A(new_n781), .B1(new_n557), .B2(new_n209), .ZN(new_n1080));
  OAI21_X1  g0880(.A(new_n840), .B1(new_n1079), .B2(new_n1080), .ZN(new_n1081));
  AOI22_X1  g0881(.A1(new_n813), .A2(G50), .B1(G97), .B2(new_n854), .ZN(new_n1082));
  OAI22_X1  g0882(.A1(new_n202), .A2(new_n802), .B1(new_n798), .B2(new_n275), .ZN(new_n1083));
  AOI21_X1  g0883(.A(new_n1083), .B1(G68), .B2(new_n806), .ZN(new_n1084));
  NOR2_X1   g0884(.A1(new_n794), .A2(new_n355), .ZN(new_n1085));
  AOI211_X1 g0885(.A(new_n400), .B(new_n1085), .C1(G159), .C2(new_n991), .ZN(new_n1086));
  NAND2_X1  g0886(.A1(new_n787), .A2(G150), .ZN(new_n1087));
  NAND4_X1  g0887(.A1(new_n1082), .A2(new_n1084), .A3(new_n1086), .A4(new_n1087), .ZN(new_n1088));
  AOI22_X1  g0888(.A1(new_n803), .A2(G294), .B1(new_n983), .B2(G283), .ZN(new_n1089));
  AOI22_X1  g0889(.A1(G322), .A2(new_n991), .B1(new_n799), .B2(G311), .ZN(new_n1090));
  XNOR2_X1  g0890(.A(new_n1090), .B(KEYINPUT120), .ZN(new_n1091));
  INV_X1    g0891(.A(G317), .ZN(new_n1092));
  OAI221_X1 g0892(.A(new_n1091), .B1(new_n819), .B2(new_n805), .C1(new_n1092), .C2(new_n812), .ZN(new_n1093));
  INV_X1    g0893(.A(KEYINPUT48), .ZN(new_n1094));
  OAI21_X1  g0894(.A(new_n1089), .B1(new_n1093), .B2(new_n1094), .ZN(new_n1095));
  AOI21_X1  g0895(.A(new_n1095), .B1(new_n1094), .B2(new_n1093), .ZN(new_n1096));
  XNOR2_X1  g0896(.A(new_n1096), .B(KEYINPUT49), .ZN(new_n1097));
  OAI221_X1 g0897(.A(new_n400), .B1(new_n792), .B2(new_n463), .C1(new_n823), .C2(new_n786), .ZN(new_n1098));
  OAI21_X1  g0898(.A(new_n1088), .B1(new_n1097), .B2(new_n1098), .ZN(new_n1099));
  AOI21_X1  g0899(.A(new_n1081), .B1(new_n1099), .B2(new_n777), .ZN(new_n1100));
  AOI22_X1  g0900(.A1(new_n1014), .A2(new_n1010), .B1(new_n1070), .B2(new_n1100), .ZN(new_n1101));
  NAND2_X1  g0901(.A1(new_n765), .A2(new_n1014), .ZN(new_n1102));
  XOR2_X1   g0902(.A(new_n716), .B(KEYINPUT121), .Z(new_n1103));
  NAND2_X1  g0903(.A1(new_n1102), .A2(new_n1103), .ZN(new_n1104));
  NOR2_X1   g0904(.A1(new_n765), .A2(new_n1014), .ZN(new_n1105));
  OAI21_X1  g0905(.A(new_n1101), .B1(new_n1104), .B2(new_n1105), .ZN(G393));
  NAND2_X1  g0906(.A1(new_n1039), .A2(new_n1010), .ZN(new_n1107));
  OAI22_X1  g0907(.A1(new_n770), .A2(new_n246), .B1(new_n221), .B2(new_n209), .ZN(new_n1108));
  OAI21_X1  g0908(.A(new_n840), .B1(new_n1108), .B2(new_n780), .ZN(new_n1109));
  OAI22_X1  g0909(.A1(new_n812), .A2(new_n848), .B1(new_n1092), .B2(new_n808), .ZN(new_n1110));
  XNOR2_X1  g0910(.A(new_n1110), .B(KEYINPUT52), .ZN(new_n1111));
  OAI21_X1  g0911(.A(new_n400), .B1(new_n798), .B2(new_n819), .ZN(new_n1112));
  OAI22_X1  g0912(.A1(new_n802), .A2(new_n815), .B1(new_n805), .B2(new_n824), .ZN(new_n1113));
  AOI211_X1 g0913(.A(new_n1112), .B(new_n1113), .C1(G116), .C2(new_n983), .ZN(new_n1114));
  AOI21_X1  g0914(.A(new_n793), .B1(G322), .B2(new_n787), .ZN(new_n1115));
  NAND3_X1  g0915(.A1(new_n1111), .A2(new_n1114), .A3(new_n1115), .ZN(new_n1116));
  OAI22_X1  g0916(.A1(new_n812), .A2(new_n860), .B1(new_n271), .B2(new_n808), .ZN(new_n1117));
  XOR2_X1   g0917(.A(new_n1117), .B(KEYINPUT51), .Z(new_n1118));
  OAI22_X1  g0918(.A1(new_n285), .A2(new_n798), .B1(new_n802), .B2(new_n308), .ZN(new_n1119));
  OAI21_X1  g0919(.A(new_n250), .B1(new_n805), .B2(new_n275), .ZN(new_n1120));
  NOR2_X1   g0920(.A1(new_n794), .A2(new_n202), .ZN(new_n1121));
  NOR3_X1   g0921(.A1(new_n1119), .A2(new_n1120), .A3(new_n1121), .ZN(new_n1122));
  OAI221_X1 g0922(.A(new_n1122), .B1(new_n434), .B2(new_n792), .C1(new_n859), .C2(new_n786), .ZN(new_n1123));
  OAI21_X1  g0923(.A(new_n1116), .B1(new_n1118), .B2(new_n1123), .ZN(new_n1124));
  AOI21_X1  g0924(.A(new_n1109), .B1(new_n1124), .B2(new_n777), .ZN(new_n1125));
  OAI21_X1  g0925(.A(new_n1125), .B1(new_n1027), .B2(new_n776), .ZN(new_n1126));
  NAND2_X1  g0926(.A1(new_n1107), .A2(new_n1126), .ZN(new_n1127));
  NAND3_X1  g0927(.A1(new_n1102), .A2(new_n1032), .A3(new_n1038), .ZN(new_n1128));
  INV_X1    g0928(.A(new_n1103), .ZN(new_n1129));
  AOI21_X1  g0929(.A(new_n1129), .B1(new_n1015), .B2(new_n1039), .ZN(new_n1130));
  AOI21_X1  g0930(.A(new_n1127), .B1(new_n1128), .B2(new_n1130), .ZN(new_n1131));
  INV_X1    g0931(.A(new_n1131), .ZN(G390));
  NOR3_X1   g0932(.A1(new_n657), .A2(new_n661), .A3(new_n655), .ZN(new_n1133));
  AOI21_X1  g0933(.A(KEYINPUT88), .B1(new_n629), .B2(new_n642), .ZN(new_n1134));
  OAI21_X1  g0934(.A(new_n665), .B1(new_n1133), .B2(new_n1134), .ZN(new_n1135));
  INV_X1    g0935(.A(new_n654), .ZN(new_n1136));
  NAND2_X1  g0936(.A1(new_n1135), .A2(new_n1136), .ZN(new_n1137));
  AND3_X1   g0937(.A1(new_n672), .A2(new_n676), .A3(new_n670), .ZN(new_n1138));
  AOI21_X1  g0938(.A(new_n697), .B1(new_n1137), .B2(new_n1138), .ZN(new_n1139));
  AOI21_X1  g0939(.A(new_n955), .B1(new_n874), .B2(new_n1139), .ZN(new_n1140));
  OAI21_X1  g0940(.A(new_n967), .B1(new_n1140), .B2(new_n906), .ZN(new_n1141));
  NAND4_X1  g0941(.A1(new_n961), .A2(new_n1141), .A3(new_n963), .A4(new_n965), .ZN(new_n1142));
  NAND2_X1  g0942(.A1(new_n726), .A2(new_n696), .ZN(new_n1143));
  OAI21_X1  g0943(.A(new_n956), .B1(new_n1143), .B2(new_n949), .ZN(new_n1144));
  NAND2_X1  g0944(.A1(new_n1144), .A2(new_n907), .ZN(new_n1145));
  NAND3_X1  g0945(.A1(new_n1145), .A2(new_n934), .A3(new_n967), .ZN(new_n1146));
  NAND2_X1  g0946(.A1(new_n1142), .A2(new_n1146), .ZN(new_n1147));
  AND4_X1   g0947(.A1(G330), .A2(new_n900), .A3(new_n874), .A4(new_n907), .ZN(new_n1148));
  NAND2_X1  g0948(.A1(new_n1147), .A2(new_n1148), .ZN(new_n1149));
  OAI21_X1  g0949(.A(new_n950), .B1(new_n762), .B2(new_n763), .ZN(new_n1150));
  NAND3_X1  g0950(.A1(new_n1142), .A2(new_n1146), .A3(new_n1150), .ZN(new_n1151));
  NAND2_X1  g0951(.A1(new_n1149), .A2(new_n1151), .ZN(new_n1152));
  NOR2_X1   g0952(.A1(new_n881), .A2(new_n832), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n1153), .A2(new_n900), .ZN(new_n1154));
  AOI21_X1  g0954(.A(new_n1144), .B1(new_n1154), .B2(new_n906), .ZN(new_n1155));
  NAND2_X1  g0955(.A1(new_n1155), .A2(new_n1150), .ZN(new_n1156));
  OAI21_X1  g0956(.A(new_n874), .B1(new_n762), .B2(new_n763), .ZN(new_n1157));
  AOI21_X1  g0957(.A(new_n1148), .B1(new_n1157), .B2(new_n906), .ZN(new_n1158));
  OAI21_X1  g0958(.A(new_n1156), .B1(new_n1158), .B2(new_n1140), .ZN(new_n1159));
  NAND3_X1  g0959(.A1(new_n1159), .A2(new_n945), .A3(new_n971), .ZN(new_n1160));
  NAND2_X1  g0960(.A1(new_n1152), .A2(new_n1160), .ZN(new_n1161));
  AOI211_X1 g0961(.A(new_n970), .B(new_n944), .C1(new_n737), .C2(new_n458), .ZN(new_n1162));
  NAND4_X1  g0962(.A1(new_n1162), .A2(new_n1149), .A3(new_n1151), .A4(new_n1159), .ZN(new_n1163));
  NAND3_X1  g0963(.A1(new_n1161), .A2(new_n1103), .A3(new_n1163), .ZN(new_n1164));
  AND2_X1   g0964(.A1(new_n1149), .A2(new_n1151), .ZN(new_n1165));
  OR2_X1    g0965(.A1(new_n966), .A2(new_n866), .ZN(new_n1166));
  OAI21_X1  g0966(.A(new_n840), .B1(new_n1073), .B2(new_n842), .ZN(new_n1167));
  AOI211_X1 g0967(.A(new_n250), .B(new_n1121), .C1(G87), .C2(new_n803), .ZN(new_n1168));
  AOI22_X1  g0968(.A1(G68), .A2(new_n854), .B1(new_n787), .B2(G294), .ZN(new_n1169));
  NAND2_X1  g0969(.A1(new_n813), .A2(G116), .ZN(new_n1170));
  OAI22_X1  g0970(.A1(new_n808), .A2(new_n815), .B1(new_n798), .B2(new_n557), .ZN(new_n1171));
  AOI21_X1  g0971(.A(new_n1171), .B1(G97), .B2(new_n806), .ZN(new_n1172));
  NAND4_X1  g0972(.A1(new_n1168), .A2(new_n1169), .A3(new_n1170), .A4(new_n1172), .ZN(new_n1173));
  OAI21_X1  g0973(.A(new_n250), .B1(new_n792), .B2(new_n285), .ZN(new_n1174));
  XOR2_X1   g0974(.A(new_n1174), .B(KEYINPUT123), .Z(new_n1175));
  NAND2_X1  g0975(.A1(new_n813), .A2(G132), .ZN(new_n1176));
  INV_X1    g0976(.A(KEYINPUT53), .ZN(new_n1177));
  OAI21_X1  g0977(.A(new_n1177), .B1(new_n802), .B2(new_n271), .ZN(new_n1178));
  NAND3_X1  g0978(.A1(new_n803), .A2(KEYINPUT53), .A3(G150), .ZN(new_n1179));
  AOI22_X1  g0979(.A1(new_n1178), .A2(new_n1179), .B1(new_n787), .B2(G125), .ZN(new_n1180));
  XOR2_X1   g0980(.A(KEYINPUT54), .B(G143), .Z(new_n1181));
  XNOR2_X1  g0981(.A(new_n1181), .B(KEYINPUT122), .ZN(new_n1182));
  NAND2_X1  g0982(.A1(new_n1182), .A2(new_n806), .ZN(new_n1183));
  INV_X1    g0983(.A(G128), .ZN(new_n1184));
  OAI22_X1  g0984(.A1(new_n808), .A2(new_n1184), .B1(new_n798), .B2(new_n856), .ZN(new_n1185));
  AOI21_X1  g0985(.A(new_n1185), .B1(G159), .B2(new_n983), .ZN(new_n1186));
  NAND4_X1  g0986(.A1(new_n1176), .A2(new_n1180), .A3(new_n1183), .A4(new_n1186), .ZN(new_n1187));
  OAI21_X1  g0987(.A(new_n1173), .B1(new_n1175), .B2(new_n1187), .ZN(new_n1188));
  AOI21_X1  g0988(.A(new_n1167), .B1(new_n1188), .B2(new_n777), .ZN(new_n1189));
  XOR2_X1   g0989(.A(new_n1189), .B(KEYINPUT124), .Z(new_n1190));
  AOI22_X1  g0990(.A1(new_n1165), .A2(new_n1010), .B1(new_n1166), .B2(new_n1190), .ZN(new_n1191));
  NAND2_X1  g0991(.A1(new_n1164), .A2(new_n1191), .ZN(G378));
  AOI21_X1  g0992(.A(KEYINPUT125), .B1(new_n683), .B2(new_n679), .ZN(new_n1193));
  INV_X1    g0993(.A(KEYINPUT125), .ZN(new_n1194));
  AOI211_X1 g0994(.A(new_n1194), .B(new_n305), .C1(new_n680), .C2(new_n682), .ZN(new_n1195));
  OAI22_X1  g0995(.A1(new_n1193), .A2(new_n1195), .B1(new_n302), .B2(new_n694), .ZN(new_n1196));
  OAI21_X1  g0996(.A(new_n1194), .B1(new_n301), .B2(new_n305), .ZN(new_n1197));
  NOR2_X1   g0997(.A1(new_n302), .A2(new_n694), .ZN(new_n1198));
  NAND3_X1  g0998(.A1(new_n683), .A2(KEYINPUT125), .A3(new_n679), .ZN(new_n1199));
  NAND3_X1  g0999(.A1(new_n1197), .A2(new_n1198), .A3(new_n1199), .ZN(new_n1200));
  XOR2_X1   g1000(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1201));
  INV_X1    g1001(.A(new_n1201), .ZN(new_n1202));
  AND3_X1   g1002(.A1(new_n1196), .A2(new_n1200), .A3(new_n1202), .ZN(new_n1203));
  AOI21_X1  g1003(.A(new_n1202), .B1(new_n1196), .B2(new_n1200), .ZN(new_n1204));
  NOR2_X1   g1004(.A1(new_n1203), .A2(new_n1204), .ZN(new_n1205));
  NAND2_X1  g1005(.A1(new_n1205), .A2(new_n774), .ZN(new_n1206));
  NOR2_X1   g1006(.A1(new_n250), .A2(G41), .ZN(new_n1207));
  AOI211_X1 g1007(.A(G50), .B(new_n1207), .C1(new_n433), .C2(new_n479), .ZN(new_n1208));
  AOI22_X1  g1008(.A1(new_n813), .A2(G107), .B1(G58), .B2(new_n854), .ZN(new_n1209));
  OAI21_X1  g1009(.A(new_n1209), .B1(new_n815), .B2(new_n786), .ZN(new_n1210));
  OAI221_X1 g1010(.A(new_n1207), .B1(new_n221), .B2(new_n798), .C1(new_n463), .C2(new_n808), .ZN(new_n1211));
  OAI22_X1  g1011(.A1(new_n802), .A2(new_n202), .B1(new_n805), .B2(new_n355), .ZN(new_n1212));
  NOR4_X1   g1012(.A1(new_n1210), .A2(new_n990), .A3(new_n1211), .A4(new_n1212), .ZN(new_n1213));
  AOI21_X1  g1013(.A(new_n1208), .B1(new_n1213), .B2(KEYINPUT58), .ZN(new_n1214));
  AOI22_X1  g1014(.A1(G128), .A2(new_n813), .B1(new_n1182), .B2(new_n803), .ZN(new_n1215));
  NAND2_X1  g1015(.A1(new_n983), .A2(G150), .ZN(new_n1216));
  NAND2_X1  g1016(.A1(new_n806), .A2(G137), .ZN(new_n1217));
  AOI22_X1  g1017(.A1(G125), .A2(new_n991), .B1(new_n799), .B2(G132), .ZN(new_n1218));
  NAND4_X1  g1018(.A1(new_n1215), .A2(new_n1216), .A3(new_n1217), .A4(new_n1218), .ZN(new_n1219));
  NOR2_X1   g1019(.A1(new_n1219), .A2(KEYINPUT59), .ZN(new_n1220));
  NAND2_X1  g1020(.A1(new_n1219), .A2(KEYINPUT59), .ZN(new_n1221));
  OAI211_X1 g1021(.A(new_n433), .B(new_n479), .C1(new_n792), .C2(new_n860), .ZN(new_n1222));
  AOI21_X1  g1022(.A(new_n1222), .B1(G124), .B2(new_n787), .ZN(new_n1223));
  NAND2_X1  g1023(.A1(new_n1221), .A2(new_n1223), .ZN(new_n1224));
  OAI221_X1 g1024(.A(new_n1214), .B1(KEYINPUT58), .B2(new_n1213), .C1(new_n1220), .C2(new_n1224), .ZN(new_n1225));
  NAND2_X1  g1025(.A1(new_n1225), .A2(new_n777), .ZN(new_n1226));
  NAND2_X1  g1026(.A1(new_n841), .A2(new_n285), .ZN(new_n1227));
  NAND4_X1  g1027(.A1(new_n1206), .A2(new_n840), .A3(new_n1226), .A4(new_n1227), .ZN(new_n1228));
  INV_X1    g1028(.A(new_n1228), .ZN(new_n1229));
  OAI21_X1  g1029(.A(new_n943), .B1(new_n1203), .B2(new_n1204), .ZN(new_n1230));
  NAND3_X1  g1030(.A1(new_n952), .A2(G330), .A3(new_n1205), .ZN(new_n1231));
  AND2_X1   g1031(.A1(new_n966), .A2(new_n968), .ZN(new_n1232));
  OAI211_X1 g1032(.A(new_n1230), .B(new_n1231), .C1(new_n1232), .C2(new_n959), .ZN(new_n1233));
  AOI21_X1  g1033(.A(new_n1205), .B1(new_n952), .B2(G330), .ZN(new_n1234));
  AND4_X1   g1034(.A1(G330), .A2(new_n935), .A3(new_n1205), .A4(new_n942), .ZN(new_n1235));
  OAI21_X1  g1035(.A(new_n969), .B1(new_n1234), .B2(new_n1235), .ZN(new_n1236));
  NAND2_X1  g1036(.A1(new_n1233), .A2(new_n1236), .ZN(new_n1237));
  AOI21_X1  g1037(.A(new_n1229), .B1(new_n1237), .B2(new_n1010), .ZN(new_n1238));
  AOI22_X1  g1038(.A1(new_n1163), .A2(new_n1162), .B1(new_n1233), .B2(new_n1236), .ZN(new_n1239));
  OAI21_X1  g1039(.A(new_n1103), .B1(new_n1239), .B2(KEYINPUT57), .ZN(new_n1240));
  INV_X1    g1040(.A(KEYINPUT57), .ZN(new_n1241));
  AOI21_X1  g1041(.A(new_n1241), .B1(new_n1163), .B2(new_n1162), .ZN(new_n1242));
  NAND2_X1  g1042(.A1(new_n1236), .A2(KEYINPUT126), .ZN(new_n1243));
  INV_X1    g1043(.A(KEYINPUT126), .ZN(new_n1244));
  OAI211_X1 g1044(.A(new_n1244), .B(new_n969), .C1(new_n1234), .C2(new_n1235), .ZN(new_n1245));
  NAND3_X1  g1045(.A1(new_n1243), .A2(new_n1233), .A3(new_n1245), .ZN(new_n1246));
  AND2_X1   g1046(.A1(new_n1242), .A2(new_n1246), .ZN(new_n1247));
  OAI21_X1  g1047(.A(new_n1238), .B1(new_n1240), .B2(new_n1247), .ZN(G375));
  NAND2_X1  g1048(.A1(new_n906), .A2(new_n774), .ZN(new_n1249));
  NOR2_X1   g1049(.A1(new_n842), .A2(G68), .ZN(new_n1250));
  AOI22_X1  g1050(.A1(new_n1182), .A2(new_n799), .B1(new_n854), .B2(G58), .ZN(new_n1251));
  OAI221_X1 g1051(.A(new_n1251), .B1(new_n1184), .B2(new_n786), .C1(new_n856), .C2(new_n812), .ZN(new_n1252));
  AOI22_X1  g1052(.A1(G159), .A2(new_n803), .B1(new_n806), .B2(G150), .ZN(new_n1253));
  AOI21_X1  g1053(.A(new_n400), .B1(new_n991), .B2(G132), .ZN(new_n1254));
  OAI211_X1 g1054(.A(new_n1253), .B(new_n1254), .C1(new_n285), .C2(new_n794), .ZN(new_n1255));
  OAI21_X1  g1055(.A(new_n400), .B1(new_n798), .B2(new_n463), .ZN(new_n1256));
  NOR2_X1   g1056(.A1(new_n1256), .A2(new_n1085), .ZN(new_n1257));
  AOI22_X1  g1057(.A1(G294), .A2(new_n991), .B1(new_n806), .B2(G107), .ZN(new_n1258));
  OAI211_X1 g1058(.A(new_n1257), .B(new_n1258), .C1(new_n221), .C2(new_n802), .ZN(new_n1259));
  AOI22_X1  g1059(.A1(G77), .A2(new_n854), .B1(new_n787), .B2(G303), .ZN(new_n1260));
  OAI21_X1  g1060(.A(new_n1260), .B1(new_n815), .B2(new_n812), .ZN(new_n1261));
  OAI22_X1  g1061(.A1(new_n1252), .A2(new_n1255), .B1(new_n1259), .B2(new_n1261), .ZN(new_n1262));
  AOI211_X1 g1062(.A(new_n838), .B(new_n1250), .C1(new_n1262), .C2(new_n777), .ZN(new_n1263));
  AOI22_X1  g1063(.A1(new_n1159), .A2(new_n1010), .B1(new_n1249), .B2(new_n1263), .ZN(new_n1264));
  NAND2_X1  g1064(.A1(new_n1160), .A2(new_n1043), .ZN(new_n1265));
  NOR2_X1   g1065(.A1(new_n1162), .A2(new_n1159), .ZN(new_n1266));
  OAI21_X1  g1066(.A(new_n1264), .B1(new_n1265), .B2(new_n1266), .ZN(G381));
  INV_X1    g1067(.A(new_n1238), .ZN(new_n1268));
  OAI21_X1  g1068(.A(new_n1162), .B1(new_n1152), .B2(new_n1160), .ZN(new_n1269));
  NAND2_X1  g1069(.A1(new_n1269), .A2(new_n1237), .ZN(new_n1270));
  AOI21_X1  g1070(.A(new_n1129), .B1(new_n1270), .B2(new_n1241), .ZN(new_n1271));
  NAND2_X1  g1071(.A1(new_n1242), .A2(new_n1246), .ZN(new_n1272));
  AOI21_X1  g1072(.A(new_n1268), .B1(new_n1271), .B2(new_n1272), .ZN(new_n1273));
  AND3_X1   g1073(.A1(new_n1064), .A2(new_n1065), .A3(new_n1067), .ZN(new_n1274));
  AOI21_X1  g1074(.A(new_n1042), .B1(new_n1040), .B2(new_n765), .ZN(new_n1275));
  OAI21_X1  g1075(.A(new_n1274), .B1(new_n1275), .B2(new_n1010), .ZN(new_n1276));
  AND3_X1   g1076(.A1(new_n1276), .A2(new_n1009), .A3(new_n1131), .ZN(new_n1277));
  INV_X1    g1077(.A(G378), .ZN(new_n1278));
  OR2_X1    g1078(.A1(G393), .A2(G396), .ZN(new_n1279));
  NOR3_X1   g1079(.A1(new_n1279), .A2(G384), .A3(G381), .ZN(new_n1280));
  NAND4_X1  g1080(.A1(new_n1273), .A2(new_n1277), .A3(new_n1278), .A4(new_n1280), .ZN(new_n1281));
  XNOR2_X1  g1081(.A(new_n1281), .B(KEYINPUT127), .ZN(G407));
  NAND2_X1  g1082(.A1(new_n1273), .A2(new_n1278), .ZN(new_n1283));
  OAI211_X1 g1083(.A(G407), .B(G213), .C1(G343), .C2(new_n1283), .ZN(G409));
  XNOR2_X1  g1084(.A(G393), .B(G396), .ZN(new_n1285));
  INV_X1    g1085(.A(new_n1285), .ZN(new_n1286));
  AOI21_X1  g1086(.A(new_n1131), .B1(new_n1276), .B2(new_n1009), .ZN(new_n1287));
  OAI21_X1  g1087(.A(new_n1286), .B1(new_n1277), .B2(new_n1287), .ZN(new_n1288));
  NAND2_X1  g1088(.A1(G387), .A2(G390), .ZN(new_n1289));
  NAND3_X1  g1089(.A1(new_n1276), .A2(new_n1009), .A3(new_n1131), .ZN(new_n1290));
  NAND3_X1  g1090(.A1(new_n1289), .A2(new_n1290), .A3(new_n1285), .ZN(new_n1291));
  NAND2_X1  g1091(.A1(new_n1288), .A2(new_n1291), .ZN(new_n1292));
  NAND2_X1  g1092(.A1(new_n1160), .A2(new_n1103), .ZN(new_n1293));
  OAI21_X1  g1093(.A(KEYINPUT60), .B1(new_n1162), .B2(new_n1159), .ZN(new_n1294));
  INV_X1    g1094(.A(new_n1159), .ZN(new_n1295));
  NAND2_X1  g1095(.A1(new_n971), .A2(new_n945), .ZN(new_n1296));
  INV_X1    g1096(.A(KEYINPUT60), .ZN(new_n1297));
  NAND3_X1  g1097(.A1(new_n1295), .A2(new_n1296), .A3(new_n1297), .ZN(new_n1298));
  AOI21_X1  g1098(.A(new_n1293), .B1(new_n1294), .B2(new_n1298), .ZN(new_n1299));
  INV_X1    g1099(.A(new_n1264), .ZN(new_n1300));
  OAI21_X1  g1100(.A(new_n888), .B1(new_n1299), .B2(new_n1300), .ZN(new_n1301));
  AND2_X1   g1101(.A1(new_n1298), .A2(new_n1294), .ZN(new_n1302));
  OAI211_X1 g1102(.A(G384), .B(new_n1264), .C1(new_n1302), .C2(new_n1293), .ZN(new_n1303));
  INV_X1    g1103(.A(G213), .ZN(new_n1304));
  NOR2_X1   g1104(.A1(new_n1304), .A2(G343), .ZN(new_n1305));
  NAND2_X1  g1105(.A1(new_n1305), .A2(G2897), .ZN(new_n1306));
  AND3_X1   g1106(.A1(new_n1301), .A2(new_n1303), .A3(new_n1306), .ZN(new_n1307));
  AOI21_X1  g1107(.A(new_n1306), .B1(new_n1301), .B2(new_n1303), .ZN(new_n1308));
  NOR2_X1   g1108(.A1(new_n1307), .A2(new_n1308), .ZN(new_n1309));
  AOI21_X1  g1109(.A(new_n1229), .B1(new_n1246), .B2(new_n1010), .ZN(new_n1310));
  NAND2_X1  g1110(.A1(new_n1239), .A2(new_n1043), .ZN(new_n1311));
  AOI21_X1  g1111(.A(G378), .B1(new_n1310), .B2(new_n1311), .ZN(new_n1312));
  AOI21_X1  g1112(.A(new_n1312), .B1(new_n1273), .B2(G378), .ZN(new_n1313));
  OAI21_X1  g1113(.A(new_n1309), .B1(new_n1313), .B2(new_n1305), .ZN(new_n1314));
  INV_X1    g1114(.A(KEYINPUT61), .ZN(new_n1315));
  OAI211_X1 g1115(.A(G378), .B(new_n1238), .C1(new_n1240), .C2(new_n1247), .ZN(new_n1316));
  NAND2_X1  g1116(.A1(new_n1310), .A2(new_n1311), .ZN(new_n1317));
  NAND2_X1  g1117(.A1(new_n1317), .A2(new_n1278), .ZN(new_n1318));
  NAND2_X1  g1118(.A1(new_n1316), .A2(new_n1318), .ZN(new_n1319));
  INV_X1    g1119(.A(KEYINPUT62), .ZN(new_n1320));
  NAND2_X1  g1120(.A1(new_n1301), .A2(new_n1303), .ZN(new_n1321));
  INV_X1    g1121(.A(new_n1321), .ZN(new_n1322));
  INV_X1    g1122(.A(new_n1305), .ZN(new_n1323));
  NAND4_X1  g1123(.A1(new_n1319), .A2(new_n1320), .A3(new_n1322), .A4(new_n1323), .ZN(new_n1324));
  NAND3_X1  g1124(.A1(new_n1314), .A2(new_n1315), .A3(new_n1324), .ZN(new_n1325));
  AOI211_X1 g1125(.A(new_n1321), .B(new_n1305), .C1(new_n1316), .C2(new_n1318), .ZN(new_n1326));
  NOR2_X1   g1126(.A1(new_n1326), .A2(new_n1320), .ZN(new_n1327));
  OAI21_X1  g1127(.A(new_n1292), .B1(new_n1325), .B2(new_n1327), .ZN(new_n1328));
  AOI21_X1  g1128(.A(new_n1305), .B1(new_n1316), .B2(new_n1318), .ZN(new_n1329));
  NAND2_X1  g1129(.A1(new_n1329), .A2(new_n1322), .ZN(new_n1330));
  INV_X1    g1130(.A(new_n1306), .ZN(new_n1331));
  NAND2_X1  g1131(.A1(new_n1321), .A2(new_n1331), .ZN(new_n1332));
  NAND3_X1  g1132(.A1(new_n1301), .A2(new_n1303), .A3(new_n1306), .ZN(new_n1333));
  NAND2_X1  g1133(.A1(new_n1332), .A2(new_n1333), .ZN(new_n1334));
  NOR2_X1   g1134(.A1(new_n1329), .A2(new_n1334), .ZN(new_n1335));
  INV_X1    g1135(.A(KEYINPUT63), .ZN(new_n1336));
  OAI21_X1  g1136(.A(new_n1330), .B1(new_n1335), .B2(new_n1336), .ZN(new_n1337));
  NAND3_X1  g1137(.A1(new_n1288), .A2(new_n1315), .A3(new_n1291), .ZN(new_n1338));
  AOI21_X1  g1138(.A(new_n1338), .B1(KEYINPUT63), .B2(new_n1326), .ZN(new_n1339));
  NAND2_X1  g1139(.A1(new_n1337), .A2(new_n1339), .ZN(new_n1340));
  NAND2_X1  g1140(.A1(new_n1328), .A2(new_n1340), .ZN(G405));
  AND3_X1   g1141(.A1(new_n1288), .A2(new_n1291), .A3(new_n1322), .ZN(new_n1342));
  AOI21_X1  g1142(.A(new_n1322), .B1(new_n1288), .B2(new_n1291), .ZN(new_n1343));
  NAND2_X1  g1143(.A1(G375), .A2(G378), .ZN(new_n1344));
  NAND2_X1  g1144(.A1(new_n1344), .A2(new_n1283), .ZN(new_n1345));
  OR3_X1    g1145(.A1(new_n1342), .A2(new_n1343), .A3(new_n1345), .ZN(new_n1346));
  OAI21_X1  g1146(.A(new_n1345), .B1(new_n1342), .B2(new_n1343), .ZN(new_n1347));
  NAND2_X1  g1147(.A1(new_n1346), .A2(new_n1347), .ZN(G402));
endmodule


