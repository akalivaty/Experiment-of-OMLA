//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 1 0 0 0 0 0 0 1 1 0 1 0 1 0 1 1 1 1 1 0 1 1 0 0 1 1 1 0 1 1 1 1 1 1 0 0 0 0 1 1 0 1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 1 0 1 1 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:39:32 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n236, new_n237,
    new_n238, new_n240, new_n241, new_n242, new_n243, new_n244, new_n245,
    new_n246, new_n248, new_n249, new_n250, new_n251, new_n252, new_n253,
    new_n254, new_n255, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n993, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1025, new_n1026, new_n1027, new_n1028,
    new_n1029, new_n1030, new_n1031, new_n1032, new_n1033, new_n1034,
    new_n1035, new_n1036, new_n1037, new_n1038, new_n1039, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1050, new_n1051, new_n1052, new_n1053,
    new_n1054, new_n1055, new_n1056, new_n1057, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1106, new_n1107, new_n1108,
    new_n1109, new_n1110, new_n1111, new_n1112, new_n1113, new_n1114,
    new_n1115, new_n1116, new_n1117, new_n1118, new_n1119, new_n1120,
    new_n1121, new_n1122, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1160, new_n1161, new_n1162, new_n1163,
    new_n1164, new_n1165, new_n1166, new_n1167, new_n1168, new_n1169,
    new_n1170, new_n1171, new_n1172, new_n1173, new_n1174, new_n1175,
    new_n1176, new_n1177, new_n1178, new_n1179, new_n1180, new_n1181,
    new_n1182, new_n1184, new_n1185, new_n1186, new_n1187, new_n1190,
    new_n1191, new_n1192, new_n1193, new_n1194, new_n1195, new_n1196,
    new_n1197, new_n1198, new_n1199, new_n1200, new_n1201, new_n1202,
    new_n1203, new_n1204, new_n1205, new_n1206, new_n1207, new_n1208,
    new_n1209, new_n1210, new_n1211, new_n1212, new_n1213, new_n1214,
    new_n1215, new_n1216, new_n1217, new_n1218, new_n1219, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1232, new_n1233,
    new_n1234, new_n1235, new_n1236;
  NOR3_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .ZN(new_n201));
  XNOR2_X1  g0001(.A(new_n201), .B(KEYINPUT64), .ZN(new_n202));
  NOR2_X1   g0002(.A1(new_n202), .A2(G77), .ZN(G353));
  OAI21_X1  g0003(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  AOI22_X1  g0004(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n205));
  XOR2_X1   g0005(.A(new_n205), .B(KEYINPUT65), .Z(new_n206));
  INV_X1    g0006(.A(G87), .ZN(new_n207));
  INV_X1    g0007(.A(G250), .ZN(new_n208));
  INV_X1    g0008(.A(G97), .ZN(new_n209));
  INV_X1    g0009(.A(G257), .ZN(new_n210));
  OAI221_X1 g0010(.A(new_n206), .B1(new_n207), .B2(new_n208), .C1(new_n209), .C2(new_n210), .ZN(new_n211));
  INV_X1    g0011(.A(G50), .ZN(new_n212));
  INV_X1    g0012(.A(G226), .ZN(new_n213));
  OAI22_X1  g0013(.A1(new_n211), .A2(KEYINPUT66), .B1(new_n212), .B2(new_n213), .ZN(new_n214));
  AOI21_X1  g0014(.A(new_n214), .B1(KEYINPUT66), .B2(new_n211), .ZN(new_n215));
  INV_X1    g0015(.A(G68), .ZN(new_n216));
  INV_X1    g0016(.A(G238), .ZN(new_n217));
  INV_X1    g0017(.A(G116), .ZN(new_n218));
  INV_X1    g0018(.A(G270), .ZN(new_n219));
  OAI221_X1 g0019(.A(new_n215), .B1(new_n216), .B2(new_n217), .C1(new_n218), .C2(new_n219), .ZN(new_n220));
  AOI21_X1  g0020(.A(new_n220), .B1(G77), .B2(G244), .ZN(new_n221));
  INV_X1    g0021(.A(G1), .ZN(new_n222));
  INV_X1    g0022(.A(G20), .ZN(new_n223));
  NOR2_X1   g0023(.A1(new_n222), .A2(new_n223), .ZN(new_n224));
  INV_X1    g0024(.A(KEYINPUT67), .ZN(new_n225));
  OAI22_X1  g0025(.A1(new_n221), .A2(new_n224), .B1(new_n225), .B2(KEYINPUT1), .ZN(new_n226));
  NAND2_X1  g0026(.A1(new_n225), .A2(KEYINPUT1), .ZN(new_n227));
  XNOR2_X1  g0027(.A(new_n226), .B(new_n227), .ZN(new_n228));
  INV_X1    g0028(.A(G58), .ZN(new_n229));
  NAND2_X1  g0029(.A1(new_n229), .A2(new_n216), .ZN(new_n230));
  NAND2_X1  g0030(.A1(new_n230), .A2(G50), .ZN(new_n231));
  NAND2_X1  g0031(.A1(G1), .A2(G13), .ZN(new_n232));
  NOR3_X1   g0032(.A1(new_n231), .A2(new_n223), .A3(new_n232), .ZN(new_n233));
  INV_X1    g0033(.A(G13), .ZN(new_n234));
  NAND2_X1  g0034(.A1(new_n224), .A2(new_n234), .ZN(new_n235));
  INV_X1    g0035(.A(new_n235), .ZN(new_n236));
  OAI211_X1 g0036(.A(new_n236), .B(G250), .C1(G257), .C2(G264), .ZN(new_n237));
  XOR2_X1   g0037(.A(new_n237), .B(KEYINPUT0), .Z(new_n238));
  NOR3_X1   g0038(.A1(new_n228), .A2(new_n233), .A3(new_n238), .ZN(G361));
  XNOR2_X1  g0039(.A(KEYINPUT2), .B(G226), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n240), .B(G232), .ZN(new_n241));
  XNOR2_X1  g0041(.A(G238), .B(G244), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XNOR2_X1  g0043(.A(G250), .B(G257), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n244), .B(G264), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n245), .B(new_n219), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n243), .B(new_n246), .ZN(G358));
  XNOR2_X1  g0047(.A(G68), .B(G77), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n248), .B(KEYINPUT68), .ZN(new_n249));
  XNOR2_X1  g0049(.A(new_n249), .B(new_n212), .ZN(new_n250));
  XNOR2_X1  g0050(.A(new_n250), .B(new_n229), .ZN(new_n251));
  XNOR2_X1  g0051(.A(G87), .B(G97), .ZN(new_n252));
  XNOR2_X1  g0052(.A(G107), .B(G116), .ZN(new_n253));
  XNOR2_X1  g0053(.A(new_n252), .B(new_n253), .ZN(new_n254));
  INV_X1    g0054(.A(new_n254), .ZN(new_n255));
  XNOR2_X1  g0055(.A(new_n251), .B(new_n255), .ZN(G351));
  NOR2_X1   g0056(.A1(G20), .A2(G33), .ZN(new_n257));
  AOI22_X1  g0057(.A1(new_n202), .A2(G20), .B1(G150), .B2(new_n257), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n229), .A2(KEYINPUT70), .ZN(new_n259));
  OR2_X1    g0059(.A1(new_n229), .A2(KEYINPUT71), .ZN(new_n260));
  OAI211_X1 g0060(.A(KEYINPUT8), .B(new_n259), .C1(new_n260), .C2(KEYINPUT70), .ZN(new_n261));
  OR2_X1    g0061(.A1(new_n260), .A2(KEYINPUT8), .ZN(new_n262));
  NAND2_X1  g0062(.A1(new_n261), .A2(new_n262), .ZN(new_n263));
  INV_X1    g0063(.A(new_n263), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n223), .A2(G33), .ZN(new_n265));
  OAI21_X1  g0065(.A(new_n258), .B1(new_n264), .B2(new_n265), .ZN(new_n266));
  NAND3_X1  g0066(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n267), .A2(KEYINPUT69), .ZN(new_n268));
  INV_X1    g0068(.A(KEYINPUT69), .ZN(new_n269));
  NAND4_X1  g0069(.A1(new_n269), .A2(G1), .A3(G20), .A4(G33), .ZN(new_n270));
  NAND3_X1  g0070(.A1(new_n268), .A2(new_n232), .A3(new_n270), .ZN(new_n271));
  NOR2_X1   g0071(.A1(new_n223), .A2(G1), .ZN(new_n272));
  XOR2_X1   g0072(.A(new_n272), .B(KEYINPUT72), .Z(new_n273));
  NAND3_X1  g0073(.A1(new_n222), .A2(G13), .A3(G20), .ZN(new_n274));
  NAND4_X1  g0074(.A1(new_n268), .A2(new_n270), .A3(new_n232), .A4(new_n274), .ZN(new_n275));
  NOR2_X1   g0075(.A1(new_n273), .A2(new_n275), .ZN(new_n276));
  AOI22_X1  g0076(.A1(new_n266), .A2(new_n271), .B1(G50), .B2(new_n276), .ZN(new_n277));
  OAI21_X1  g0077(.A(new_n277), .B1(G50), .B2(new_n274), .ZN(new_n278));
  INV_X1    g0078(.A(KEYINPUT3), .ZN(new_n279));
  INV_X1    g0079(.A(G33), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n279), .A2(new_n280), .ZN(new_n281));
  NAND2_X1  g0081(.A1(KEYINPUT3), .A2(G33), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n281), .A2(new_n282), .ZN(new_n283));
  INV_X1    g0083(.A(G1698), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n284), .A2(G222), .ZN(new_n285));
  NAND2_X1  g0085(.A1(G223), .A2(G1698), .ZN(new_n286));
  NAND3_X1  g0086(.A1(new_n283), .A2(new_n285), .A3(new_n286), .ZN(new_n287));
  INV_X1    g0087(.A(G41), .ZN(new_n288));
  OAI211_X1 g0088(.A(G1), .B(G13), .C1(new_n280), .C2(new_n288), .ZN(new_n289));
  INV_X1    g0089(.A(new_n289), .ZN(new_n290));
  OAI211_X1 g0090(.A(new_n287), .B(new_n290), .C1(G77), .C2(new_n283), .ZN(new_n291));
  OAI21_X1  g0091(.A(new_n222), .B1(G41), .B2(G45), .ZN(new_n292));
  INV_X1    g0092(.A(G274), .ZN(new_n293));
  NOR2_X1   g0093(.A1(new_n292), .A2(new_n293), .ZN(new_n294));
  INV_X1    g0094(.A(new_n294), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n289), .A2(new_n292), .ZN(new_n296));
  OAI211_X1 g0096(.A(new_n291), .B(new_n295), .C1(new_n213), .C2(new_n296), .ZN(new_n297));
  INV_X1    g0097(.A(G169), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n297), .A2(new_n298), .ZN(new_n299));
  OAI211_X1 g0099(.A(new_n278), .B(new_n299), .C1(G179), .C2(new_n297), .ZN(new_n300));
  XNOR2_X1  g0100(.A(KEYINPUT8), .B(G58), .ZN(new_n301));
  INV_X1    g0101(.A(new_n301), .ZN(new_n302));
  AOI22_X1  g0102(.A1(new_n302), .A2(new_n257), .B1(G20), .B2(G77), .ZN(new_n303));
  XOR2_X1   g0103(.A(KEYINPUT15), .B(G87), .Z(new_n304));
  INV_X1    g0104(.A(new_n304), .ZN(new_n305));
  OAI21_X1  g0105(.A(new_n303), .B1(new_n265), .B2(new_n305), .ZN(new_n306));
  AOI22_X1  g0106(.A1(new_n271), .A2(new_n306), .B1(new_n276), .B2(G77), .ZN(new_n307));
  INV_X1    g0107(.A(new_n274), .ZN(new_n308));
  INV_X1    g0108(.A(G77), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n308), .A2(new_n309), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n307), .A2(new_n310), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n284), .A2(G232), .ZN(new_n312));
  OAI211_X1 g0112(.A(new_n283), .B(new_n312), .C1(new_n217), .C2(new_n284), .ZN(new_n313));
  OAI211_X1 g0113(.A(new_n313), .B(new_n290), .C1(G107), .C2(new_n283), .ZN(new_n314));
  INV_X1    g0114(.A(new_n296), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n315), .A2(G244), .ZN(new_n316));
  NAND3_X1  g0116(.A1(new_n314), .A2(new_n295), .A3(new_n316), .ZN(new_n317));
  INV_X1    g0117(.A(new_n317), .ZN(new_n318));
  INV_X1    g0118(.A(G179), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n318), .A2(new_n319), .ZN(new_n320));
  OAI211_X1 g0120(.A(new_n311), .B(new_n320), .C1(G169), .C2(new_n318), .ZN(new_n321));
  INV_X1    g0121(.A(KEYINPUT73), .ZN(new_n322));
  INV_X1    g0122(.A(KEYINPUT9), .ZN(new_n323));
  AOI21_X1  g0123(.A(new_n278), .B1(new_n322), .B2(new_n323), .ZN(new_n324));
  NAND2_X1  g0124(.A1(KEYINPUT73), .A2(KEYINPUT9), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n324), .A2(new_n325), .ZN(new_n326));
  NAND3_X1  g0126(.A1(new_n278), .A2(KEYINPUT73), .A3(KEYINPUT9), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n326), .A2(new_n327), .ZN(new_n328));
  INV_X1    g0128(.A(KEYINPUT10), .ZN(new_n329));
  INV_X1    g0129(.A(G190), .ZN(new_n330));
  NOR2_X1   g0130(.A1(new_n297), .A2(new_n330), .ZN(new_n331));
  AOI21_X1  g0131(.A(new_n331), .B1(G200), .B2(new_n297), .ZN(new_n332));
  AND3_X1   g0132(.A1(new_n328), .A2(new_n329), .A3(new_n332), .ZN(new_n333));
  AOI21_X1  g0133(.A(new_n329), .B1(new_n328), .B2(new_n332), .ZN(new_n334));
  OAI211_X1 g0134(.A(new_n300), .B(new_n321), .C1(new_n333), .C2(new_n334), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n213), .A2(new_n284), .ZN(new_n336));
  OAI211_X1 g0136(.A(new_n283), .B(new_n336), .C1(G232), .C2(new_n284), .ZN(new_n337));
  NAND2_X1  g0137(.A1(G33), .A2(G97), .ZN(new_n338));
  AOI21_X1  g0138(.A(new_n289), .B1(new_n337), .B2(new_n338), .ZN(new_n339));
  AOI211_X1 g0139(.A(new_n294), .B(new_n339), .C1(G238), .C2(new_n315), .ZN(new_n340));
  XNOR2_X1  g0140(.A(KEYINPUT74), .B(KEYINPUT13), .ZN(new_n341));
  INV_X1    g0141(.A(new_n341), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n340), .A2(new_n342), .ZN(new_n343));
  NOR2_X1   g0143(.A1(new_n339), .A2(new_n294), .ZN(new_n344));
  OAI21_X1  g0144(.A(new_n344), .B1(new_n217), .B2(new_n296), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n345), .A2(new_n341), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n343), .A2(new_n346), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n347), .A2(G169), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n348), .A2(KEYINPUT14), .ZN(new_n349));
  INV_X1    g0149(.A(KEYINPUT75), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n340), .A2(new_n350), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n345), .A2(KEYINPUT75), .ZN(new_n352));
  NAND3_X1  g0152(.A1(new_n351), .A2(KEYINPUT13), .A3(new_n352), .ZN(new_n353));
  NAND3_X1  g0153(.A1(new_n353), .A2(G179), .A3(new_n343), .ZN(new_n354));
  INV_X1    g0154(.A(KEYINPUT14), .ZN(new_n355));
  NAND3_X1  g0155(.A1(new_n347), .A2(new_n355), .A3(G169), .ZN(new_n356));
  NAND3_X1  g0156(.A1(new_n349), .A2(new_n354), .A3(new_n356), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n276), .A2(G68), .ZN(new_n358));
  XOR2_X1   g0158(.A(new_n358), .B(KEYINPUT76), .Z(new_n359));
  AOI22_X1  g0159(.A1(new_n257), .A2(G50), .B1(G20), .B2(new_n216), .ZN(new_n360));
  OAI21_X1  g0160(.A(new_n360), .B1(new_n309), .B2(new_n265), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n361), .A2(new_n271), .ZN(new_n362));
  XNOR2_X1  g0162(.A(new_n362), .B(KEYINPUT11), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n222), .A2(G13), .ZN(new_n364));
  INV_X1    g0164(.A(new_n364), .ZN(new_n365));
  NAND3_X1  g0165(.A1(new_n365), .A2(G20), .A3(new_n216), .ZN(new_n366));
  XNOR2_X1  g0166(.A(new_n366), .B(KEYINPUT12), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n363), .A2(new_n367), .ZN(new_n368));
  NOR2_X1   g0168(.A1(new_n359), .A2(new_n368), .ZN(new_n369));
  INV_X1    g0169(.A(new_n369), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n357), .A2(new_n370), .ZN(new_n371));
  INV_X1    g0171(.A(KEYINPUT18), .ZN(new_n372));
  OR2_X1    g0172(.A1(G223), .A2(G1698), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n213), .A2(G1698), .ZN(new_n374));
  AND2_X1   g0174(.A1(KEYINPUT3), .A2(G33), .ZN(new_n375));
  NOR2_X1   g0175(.A1(KEYINPUT3), .A2(G33), .ZN(new_n376));
  OAI211_X1 g0176(.A(new_n373), .B(new_n374), .C1(new_n375), .C2(new_n376), .ZN(new_n377));
  NAND2_X1  g0177(.A1(G33), .A2(G87), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n377), .A2(new_n378), .ZN(new_n379));
  INV_X1    g0179(.A(KEYINPUT78), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n379), .A2(new_n380), .ZN(new_n381));
  NAND3_X1  g0181(.A1(new_n377), .A2(KEYINPUT78), .A3(new_n378), .ZN(new_n382));
  NAND3_X1  g0182(.A1(new_n381), .A2(new_n290), .A3(new_n382), .ZN(new_n383));
  AOI21_X1  g0183(.A(new_n294), .B1(new_n315), .B2(G232), .ZN(new_n384));
  NAND2_X1  g0184(.A1(new_n383), .A2(new_n384), .ZN(new_n385));
  NAND2_X1  g0185(.A1(new_n385), .A2(G169), .ZN(new_n386));
  NAND3_X1  g0186(.A1(new_n383), .A2(G179), .A3(new_n384), .ZN(new_n387));
  XNOR2_X1  g0187(.A(KEYINPUT70), .B(G58), .ZN(new_n388));
  OAI21_X1  g0188(.A(new_n230), .B1(new_n388), .B2(new_n216), .ZN(new_n389));
  AOI22_X1  g0189(.A1(new_n389), .A2(G20), .B1(G159), .B2(new_n257), .ZN(new_n390));
  NAND3_X1  g0190(.A1(new_n281), .A2(new_n223), .A3(new_n282), .ZN(new_n391));
  INV_X1    g0191(.A(KEYINPUT7), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n391), .A2(new_n392), .ZN(new_n393));
  NAND4_X1  g0193(.A1(new_n281), .A2(KEYINPUT7), .A3(new_n223), .A4(new_n282), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n393), .A2(new_n394), .ZN(new_n395));
  AOI21_X1  g0195(.A(KEYINPUT77), .B1(new_n395), .B2(G68), .ZN(new_n396));
  INV_X1    g0196(.A(KEYINPUT77), .ZN(new_n397));
  AOI211_X1 g0197(.A(new_n397), .B(new_n216), .C1(new_n393), .C2(new_n394), .ZN(new_n398));
  OAI211_X1 g0198(.A(KEYINPUT16), .B(new_n390), .C1(new_n396), .C2(new_n398), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n395), .A2(G68), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n400), .A2(new_n390), .ZN(new_n401));
  INV_X1    g0201(.A(KEYINPUT16), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n401), .A2(new_n402), .ZN(new_n403));
  NAND3_X1  g0203(.A1(new_n399), .A2(new_n403), .A3(new_n271), .ZN(new_n404));
  NOR2_X1   g0204(.A1(new_n263), .A2(new_n274), .ZN(new_n405));
  AOI21_X1  g0205(.A(new_n405), .B1(new_n276), .B2(new_n263), .ZN(new_n406));
  AOI221_X4 g0206(.A(new_n372), .B1(new_n386), .B2(new_n387), .C1(new_n404), .C2(new_n406), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n404), .A2(new_n406), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n386), .A2(new_n387), .ZN(new_n409));
  AOI21_X1  g0209(.A(KEYINPUT18), .B1(new_n408), .B2(new_n409), .ZN(new_n410));
  NOR2_X1   g0210(.A1(new_n407), .A2(new_n410), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n385), .A2(G200), .ZN(new_n412));
  NAND3_X1  g0212(.A1(new_n383), .A2(G190), .A3(new_n384), .ZN(new_n413));
  NAND4_X1  g0213(.A1(new_n404), .A2(new_n406), .A3(new_n412), .A4(new_n413), .ZN(new_n414));
  NOR2_X1   g0214(.A1(KEYINPUT79), .A2(KEYINPUT17), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n414), .A2(new_n415), .ZN(new_n416));
  AND2_X1   g0216(.A1(new_n412), .A2(new_n413), .ZN(new_n417));
  XOR2_X1   g0217(.A(KEYINPUT79), .B(KEYINPUT17), .Z(new_n418));
  NAND4_X1  g0218(.A1(new_n417), .A2(new_n404), .A3(new_n406), .A4(new_n418), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n416), .A2(new_n419), .ZN(new_n420));
  NOR2_X1   g0220(.A1(new_n411), .A2(new_n420), .ZN(new_n421));
  NAND3_X1  g0221(.A1(new_n353), .A2(G190), .A3(new_n343), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n347), .A2(G200), .ZN(new_n423));
  NAND3_X1  g0223(.A1(new_n422), .A2(new_n369), .A3(new_n423), .ZN(new_n424));
  AOI21_X1  g0224(.A(new_n311), .B1(G190), .B2(new_n318), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n317), .A2(G200), .ZN(new_n426));
  AND2_X1   g0226(.A1(new_n425), .A2(new_n426), .ZN(new_n427));
  INV_X1    g0227(.A(new_n427), .ZN(new_n428));
  NAND4_X1  g0228(.A1(new_n371), .A2(new_n421), .A3(new_n424), .A4(new_n428), .ZN(new_n429));
  NOR2_X1   g0229(.A1(new_n335), .A2(new_n429), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n218), .A2(G20), .ZN(new_n431));
  NAND2_X1  g0231(.A1(G33), .A2(G283), .ZN(new_n432));
  OAI211_X1 g0232(.A(new_n432), .B(new_n223), .C1(G33), .C2(new_n209), .ZN(new_n433));
  NAND3_X1  g0233(.A1(new_n271), .A2(new_n431), .A3(new_n433), .ZN(new_n434));
  XNOR2_X1  g0234(.A(KEYINPUT92), .B(KEYINPUT20), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n434), .A2(new_n435), .ZN(new_n436));
  AND3_X1   g0236(.A1(new_n268), .A2(new_n232), .A3(new_n270), .ZN(new_n437));
  NOR2_X1   g0237(.A1(new_n280), .A2(G1), .ZN(new_n438));
  INV_X1    g0238(.A(new_n438), .ZN(new_n439));
  NAND4_X1  g0239(.A1(new_n437), .A2(G116), .A3(new_n274), .A4(new_n439), .ZN(new_n440));
  INV_X1    g0240(.A(KEYINPUT92), .ZN(new_n441));
  NOR2_X1   g0241(.A1(new_n441), .A2(KEYINPUT20), .ZN(new_n442));
  NAND4_X1  g0242(.A1(new_n271), .A2(new_n442), .A3(new_n431), .A4(new_n433), .ZN(new_n443));
  OR2_X1    g0243(.A1(new_n364), .A2(new_n431), .ZN(new_n444));
  NAND4_X1  g0244(.A1(new_n436), .A2(new_n440), .A3(new_n443), .A4(new_n444), .ZN(new_n445));
  NAND2_X1  g0245(.A1(G264), .A2(G1698), .ZN(new_n446));
  OAI221_X1 g0246(.A(new_n446), .B1(new_n210), .B2(G1698), .C1(new_n375), .C2(new_n376), .ZN(new_n447));
  NOR2_X1   g0247(.A1(new_n375), .A2(new_n376), .ZN(new_n448));
  INV_X1    g0248(.A(G303), .ZN(new_n449));
  NAND2_X1  g0249(.A1(new_n448), .A2(new_n449), .ZN(new_n450));
  NAND3_X1  g0250(.A1(new_n447), .A2(new_n450), .A3(new_n290), .ZN(new_n451));
  INV_X1    g0251(.A(KEYINPUT83), .ZN(new_n452));
  INV_X1    g0252(.A(KEYINPUT5), .ZN(new_n453));
  OAI21_X1  g0253(.A(new_n452), .B1(new_n453), .B2(G41), .ZN(new_n454));
  NAND3_X1  g0254(.A1(new_n288), .A2(KEYINPUT83), .A3(KEYINPUT5), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n454), .A2(new_n455), .ZN(new_n456));
  OAI211_X1 g0256(.A(new_n222), .B(G45), .C1(new_n288), .C2(KEYINPUT5), .ZN(new_n457));
  OAI211_X1 g0257(.A(G270), .B(new_n289), .C1(new_n456), .C2(new_n457), .ZN(new_n458));
  AND3_X1   g0258(.A1(new_n454), .A2(KEYINPUT84), .A3(new_n455), .ZN(new_n459));
  AOI21_X1  g0259(.A(KEYINPUT84), .B1(new_n454), .B2(new_n455), .ZN(new_n460));
  NOR2_X1   g0260(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  NAND2_X1  g0261(.A1(new_n457), .A2(KEYINPUT82), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n453), .A2(G41), .ZN(new_n463));
  INV_X1    g0263(.A(KEYINPUT82), .ZN(new_n464));
  NAND4_X1  g0264(.A1(new_n463), .A2(new_n464), .A3(new_n222), .A4(G45), .ZN(new_n465));
  NAND4_X1  g0265(.A1(new_n462), .A2(new_n465), .A3(new_n289), .A4(G274), .ZN(new_n466));
  OAI211_X1 g0266(.A(new_n451), .B(new_n458), .C1(new_n461), .C2(new_n466), .ZN(new_n467));
  NAND3_X1  g0267(.A1(new_n445), .A2(G169), .A3(new_n467), .ZN(new_n468));
  INV_X1    g0268(.A(KEYINPUT21), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n470), .A2(KEYINPUT93), .ZN(new_n471));
  NAND3_X1  g0271(.A1(new_n467), .A2(KEYINPUT21), .A3(G169), .ZN(new_n472));
  AND2_X1   g0272(.A1(new_n465), .A2(new_n289), .ZN(new_n473));
  AOI21_X1  g0273(.A(new_n293), .B1(new_n457), .B2(KEYINPUT82), .ZN(new_n474));
  OAI211_X1 g0274(.A(new_n473), .B(new_n474), .C1(new_n460), .C2(new_n459), .ZN(new_n475));
  NAND4_X1  g0275(.A1(new_n475), .A2(G179), .A3(new_n451), .A4(new_n458), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n472), .A2(new_n476), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n477), .A2(new_n445), .ZN(new_n478));
  INV_X1    g0278(.A(KEYINPUT93), .ZN(new_n479));
  NAND3_X1  g0279(.A1(new_n468), .A2(new_n479), .A3(new_n469), .ZN(new_n480));
  NAND3_X1  g0280(.A1(new_n471), .A2(new_n478), .A3(new_n480), .ZN(new_n481));
  INV_X1    g0281(.A(new_n481), .ZN(new_n482));
  NOR2_X1   g0282(.A1(new_n223), .A2(G107), .ZN(new_n483));
  XNOR2_X1  g0283(.A(new_n483), .B(KEYINPUT23), .ZN(new_n484));
  NAND2_X1  g0284(.A1(G33), .A2(G116), .ZN(new_n485));
  NOR2_X1   g0285(.A1(new_n485), .A2(G20), .ZN(new_n486));
  INV_X1    g0286(.A(new_n486), .ZN(new_n487));
  INV_X1    g0287(.A(KEYINPUT22), .ZN(new_n488));
  AOI21_X1  g0288(.A(G20), .B1(new_n281), .B2(new_n282), .ZN(new_n489));
  AOI21_X1  g0289(.A(new_n488), .B1(new_n489), .B2(G87), .ZN(new_n490));
  OAI211_X1 g0290(.A(new_n223), .B(G87), .C1(new_n375), .C2(new_n376), .ZN(new_n491));
  NOR2_X1   g0291(.A1(new_n491), .A2(KEYINPUT22), .ZN(new_n492));
  OAI211_X1 g0292(.A(new_n484), .B(new_n487), .C1(new_n490), .C2(new_n492), .ZN(new_n493));
  INV_X1    g0293(.A(KEYINPUT24), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n491), .A2(KEYINPUT22), .ZN(new_n496));
  NAND4_X1  g0296(.A1(new_n283), .A2(new_n488), .A3(new_n223), .A4(G87), .ZN(new_n497));
  AOI21_X1  g0297(.A(new_n486), .B1(new_n496), .B2(new_n497), .ZN(new_n498));
  NAND3_X1  g0298(.A1(new_n498), .A2(KEYINPUT24), .A3(new_n484), .ZN(new_n499));
  NAND3_X1  g0299(.A1(new_n495), .A2(new_n271), .A3(new_n499), .ZN(new_n500));
  NOR2_X1   g0300(.A1(new_n275), .A2(new_n438), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n501), .A2(G107), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n365), .A2(new_n483), .ZN(new_n503));
  XOR2_X1   g0303(.A(new_n503), .B(KEYINPUT25), .Z(new_n504));
  NAND3_X1  g0304(.A1(new_n500), .A2(new_n502), .A3(new_n504), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n210), .A2(G1698), .ZN(new_n506));
  OAI221_X1 g0306(.A(new_n506), .B1(G250), .B2(G1698), .C1(new_n375), .C2(new_n376), .ZN(new_n507));
  NAND2_X1  g0307(.A1(G33), .A2(G294), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n509), .A2(new_n290), .ZN(new_n510));
  OAI211_X1 g0310(.A(G264), .B(new_n289), .C1(new_n456), .C2(new_n457), .ZN(new_n511));
  OAI211_X1 g0311(.A(new_n510), .B(new_n511), .C1(new_n461), .C2(new_n466), .ZN(new_n512));
  NOR2_X1   g0312(.A1(new_n512), .A2(G179), .ZN(new_n513));
  INV_X1    g0313(.A(new_n456), .ZN(new_n514));
  INV_X1    g0314(.A(new_n457), .ZN(new_n515));
  AOI21_X1  g0315(.A(new_n290), .B1(new_n514), .B2(new_n515), .ZN(new_n516));
  AOI22_X1  g0316(.A1(new_n516), .A2(G264), .B1(new_n509), .B2(new_n290), .ZN(new_n517));
  AOI21_X1  g0317(.A(G169), .B1(new_n517), .B2(new_n475), .ZN(new_n518));
  NOR2_X1   g0318(.A1(new_n513), .A2(new_n518), .ZN(new_n519));
  AND2_X1   g0319(.A1(new_n505), .A2(new_n519), .ZN(new_n520));
  INV_X1    g0320(.A(new_n520), .ZN(new_n521));
  INV_X1    g0321(.A(new_n445), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n467), .A2(G200), .ZN(new_n523));
  OAI211_X1 g0323(.A(new_n522), .B(new_n523), .C1(new_n330), .C2(new_n467), .ZN(new_n524));
  AND2_X1   g0324(.A1(new_n500), .A2(new_n504), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n512), .A2(G200), .ZN(new_n526));
  NAND3_X1  g0326(.A1(new_n517), .A2(G190), .A3(new_n475), .ZN(new_n527));
  NAND4_X1  g0327(.A1(new_n525), .A2(new_n502), .A3(new_n526), .A4(new_n527), .ZN(new_n528));
  NAND4_X1  g0328(.A1(new_n482), .A2(new_n521), .A3(new_n524), .A4(new_n528), .ZN(new_n529));
  INV_X1    g0329(.A(KEYINPUT81), .ZN(new_n530));
  NAND2_X1  g0330(.A1(KEYINPUT80), .A2(KEYINPUT4), .ZN(new_n531));
  OAI211_X1 g0331(.A(new_n284), .B(G244), .C1(KEYINPUT80), .C2(KEYINPUT4), .ZN(new_n532));
  OAI21_X1  g0332(.A(new_n531), .B1(new_n448), .B2(new_n532), .ZN(new_n533));
  INV_X1    g0333(.A(G244), .ZN(new_n534));
  NOR2_X1   g0334(.A1(new_n534), .A2(G1698), .ZN(new_n535));
  NAND4_X1  g0335(.A1(new_n283), .A2(KEYINPUT80), .A3(KEYINPUT4), .A4(new_n535), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n533), .A2(new_n536), .ZN(new_n537));
  NAND3_X1  g0337(.A1(new_n283), .A2(G250), .A3(G1698), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n538), .A2(new_n432), .ZN(new_n539));
  OAI21_X1  g0339(.A(new_n530), .B1(new_n537), .B2(new_n539), .ZN(new_n540));
  AOI21_X1  g0340(.A(new_n208), .B1(new_n281), .B2(new_n282), .ZN(new_n541));
  AOI22_X1  g0341(.A1(new_n541), .A2(G1698), .B1(G33), .B2(G283), .ZN(new_n542));
  NAND4_X1  g0342(.A1(new_n542), .A2(KEYINPUT81), .A3(new_n533), .A4(new_n536), .ZN(new_n543));
  NAND3_X1  g0343(.A1(new_n540), .A2(new_n290), .A3(new_n543), .ZN(new_n544));
  INV_X1    g0344(.A(KEYINPUT85), .ZN(new_n545));
  OAI211_X1 g0345(.A(G257), .B(new_n289), .C1(new_n456), .C2(new_n457), .ZN(new_n546));
  AOI21_X1  g0346(.A(new_n545), .B1(new_n475), .B2(new_n546), .ZN(new_n547));
  OAI211_X1 g0347(.A(new_n545), .B(new_n546), .C1(new_n461), .C2(new_n466), .ZN(new_n548));
  INV_X1    g0348(.A(new_n548), .ZN(new_n549));
  OAI21_X1  g0349(.A(new_n544), .B1(new_n547), .B2(new_n549), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n550), .A2(new_n298), .ZN(new_n551));
  NOR3_X1   g0351(.A1(new_n275), .A2(new_n209), .A3(new_n438), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n395), .A2(G107), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n257), .A2(G77), .ZN(new_n554));
  INV_X1    g0354(.A(G107), .ZN(new_n555));
  NOR2_X1   g0355(.A1(new_n209), .A2(new_n555), .ZN(new_n556));
  NOR2_X1   g0356(.A1(G97), .A2(G107), .ZN(new_n557));
  NOR2_X1   g0357(.A1(new_n556), .A2(new_n557), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n555), .A2(G97), .ZN(new_n559));
  MUX2_X1   g0359(.A(new_n558), .B(new_n559), .S(KEYINPUT6), .Z(new_n560));
  OAI211_X1 g0360(.A(new_n553), .B(new_n554), .C1(new_n560), .C2(new_n223), .ZN(new_n561));
  AOI21_X1  g0361(.A(new_n552), .B1(new_n561), .B2(new_n271), .ZN(new_n562));
  NOR2_X1   g0362(.A1(new_n274), .A2(G97), .ZN(new_n563));
  INV_X1    g0363(.A(new_n563), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n562), .A2(new_n564), .ZN(new_n565));
  OAI21_X1  g0365(.A(new_n546), .B1(new_n461), .B2(new_n466), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n566), .A2(KEYINPUT85), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n567), .A2(new_n548), .ZN(new_n568));
  NAND3_X1  g0368(.A1(new_n568), .A2(new_n319), .A3(new_n544), .ZN(new_n569));
  NAND3_X1  g0369(.A1(new_n551), .A2(new_n565), .A3(new_n569), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n550), .A2(G200), .ZN(new_n571));
  AOI211_X1 g0371(.A(new_n563), .B(new_n552), .C1(new_n561), .C2(new_n271), .ZN(new_n572));
  NAND3_X1  g0372(.A1(new_n568), .A2(G190), .A3(new_n544), .ZN(new_n573));
  NAND3_X1  g0373(.A1(new_n571), .A2(new_n572), .A3(new_n573), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n570), .A2(new_n574), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n575), .A2(KEYINPUT86), .ZN(new_n576));
  INV_X1    g0376(.A(KEYINPUT90), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n217), .A2(new_n284), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n534), .A2(G1698), .ZN(new_n579));
  OAI211_X1 g0379(.A(new_n578), .B(new_n579), .C1(new_n375), .C2(new_n376), .ZN(new_n580));
  AOI21_X1  g0380(.A(new_n289), .B1(new_n580), .B2(new_n485), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n222), .A2(G45), .ZN(new_n582));
  AND2_X1   g0382(.A1(G33), .A2(G41), .ZN(new_n583));
  OAI211_X1 g0383(.A(new_n582), .B(G250), .C1(new_n583), .C2(new_n232), .ZN(new_n584));
  INV_X1    g0384(.A(new_n584), .ZN(new_n585));
  NOR2_X1   g0385(.A1(new_n581), .A2(new_n585), .ZN(new_n586));
  NAND3_X1  g0386(.A1(new_n222), .A2(G45), .A3(G274), .ZN(new_n587));
  INV_X1    g0387(.A(KEYINPUT87), .ZN(new_n588));
  XNOR2_X1  g0388(.A(new_n587), .B(new_n588), .ZN(new_n589));
  INV_X1    g0389(.A(new_n589), .ZN(new_n590));
  AND4_X1   g0390(.A1(KEYINPUT89), .A2(new_n586), .A3(G190), .A4(new_n590), .ZN(new_n591));
  NOR3_X1   g0391(.A1(new_n581), .A2(new_n589), .A3(new_n585), .ZN(new_n592));
  AOI21_X1  g0392(.A(KEYINPUT89), .B1(new_n592), .B2(G190), .ZN(new_n593));
  OAI21_X1  g0393(.A(new_n577), .B1(new_n591), .B2(new_n593), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n489), .A2(G68), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n557), .A2(new_n207), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n338), .A2(new_n223), .ZN(new_n597));
  NAND3_X1  g0397(.A1(new_n596), .A2(KEYINPUT19), .A3(new_n597), .ZN(new_n598));
  INV_X1    g0398(.A(KEYINPUT19), .ZN(new_n599));
  OAI21_X1  g0399(.A(new_n599), .B1(new_n338), .B2(G20), .ZN(new_n600));
  NAND3_X1  g0400(.A1(new_n595), .A2(new_n598), .A3(new_n600), .ZN(new_n601));
  AOI22_X1  g0401(.A1(new_n601), .A2(new_n271), .B1(new_n308), .B2(new_n305), .ZN(new_n602));
  AOI21_X1  g0402(.A(KEYINPUT88), .B1(new_n501), .B2(G87), .ZN(new_n603));
  INV_X1    g0403(.A(KEYINPUT88), .ZN(new_n604));
  NOR4_X1   g0404(.A1(new_n275), .A2(new_n604), .A3(new_n207), .A4(new_n438), .ZN(new_n605));
  OAI21_X1  g0405(.A(new_n602), .B1(new_n603), .B2(new_n605), .ZN(new_n606));
  INV_X1    g0406(.A(G200), .ZN(new_n607));
  NOR2_X1   g0407(.A1(new_n592), .A2(new_n607), .ZN(new_n608));
  NOR2_X1   g0408(.A1(new_n606), .A2(new_n608), .ZN(new_n609));
  NAND3_X1  g0409(.A1(new_n586), .A2(G190), .A3(new_n590), .ZN(new_n610));
  INV_X1    g0410(.A(KEYINPUT89), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  NAND3_X1  g0412(.A1(new_n592), .A2(KEYINPUT89), .A3(G190), .ZN(new_n613));
  NAND3_X1  g0413(.A1(new_n612), .A2(KEYINPUT90), .A3(new_n613), .ZN(new_n614));
  NAND3_X1  g0414(.A1(new_n594), .A2(new_n609), .A3(new_n614), .ZN(new_n615));
  INV_X1    g0415(.A(new_n592), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n501), .A2(new_n304), .ZN(new_n617));
  AOI22_X1  g0417(.A1(new_n298), .A2(new_n616), .B1(new_n602), .B2(new_n617), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n592), .A2(new_n319), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  AND2_X1   g0420(.A1(new_n615), .A2(new_n620), .ZN(new_n621));
  INV_X1    g0421(.A(KEYINPUT86), .ZN(new_n622));
  NAND3_X1  g0422(.A1(new_n570), .A2(new_n574), .A3(new_n622), .ZN(new_n623));
  NAND3_X1  g0423(.A1(new_n576), .A2(new_n621), .A3(new_n623), .ZN(new_n624));
  INV_X1    g0424(.A(KEYINPUT91), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  NAND4_X1  g0426(.A1(new_n576), .A2(KEYINPUT91), .A3(new_n621), .A4(new_n623), .ZN(new_n627));
  AOI21_X1  g0427(.A(new_n529), .B1(new_n626), .B2(new_n627), .ZN(new_n628));
  AND2_X1   g0428(.A1(new_n430), .A2(new_n628), .ZN(G372));
  INV_X1    g0429(.A(new_n424), .ZN(new_n630));
  AOI21_X1  g0430(.A(new_n630), .B1(new_n371), .B2(new_n321), .ZN(new_n631));
  INV_X1    g0431(.A(new_n420), .ZN(new_n632));
  AND2_X1   g0432(.A1(new_n631), .A2(new_n632), .ZN(new_n633));
  OAI22_X1  g0433(.A1(new_n633), .A2(new_n411), .B1(new_n334), .B2(new_n333), .ZN(new_n634));
  AND2_X1   g0434(.A1(new_n634), .A2(new_n300), .ZN(new_n635));
  INV_X1    g0435(.A(new_n430), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n615), .A2(new_n620), .ZN(new_n637));
  OAI21_X1  g0437(.A(KEYINPUT26), .B1(new_n637), .B2(new_n570), .ZN(new_n638));
  INV_X1    g0438(.A(new_n569), .ZN(new_n639));
  AOI21_X1  g0439(.A(G169), .B1(new_n568), .B2(new_n544), .ZN(new_n640));
  NOR2_X1   g0440(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  INV_X1    g0441(.A(KEYINPUT26), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n612), .A2(new_n613), .ZN(new_n643));
  AOI22_X1  g0443(.A1(new_n609), .A2(new_n643), .B1(new_n618), .B2(new_n619), .ZN(new_n644));
  NAND4_X1  g0444(.A1(new_n641), .A2(new_n642), .A3(new_n565), .A4(new_n644), .ZN(new_n645));
  NAND3_X1  g0445(.A1(new_n638), .A2(new_n620), .A3(new_n645), .ZN(new_n646));
  OAI21_X1  g0446(.A(new_n644), .B1(new_n481), .B2(new_n520), .ZN(new_n647));
  NAND3_X1  g0447(.A1(new_n528), .A2(new_n570), .A3(new_n574), .ZN(new_n648));
  NOR2_X1   g0448(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  NOR2_X1   g0449(.A1(new_n646), .A2(new_n649), .ZN(new_n650));
  OAI21_X1  g0450(.A(new_n635), .B1(new_n636), .B2(new_n650), .ZN(G369));
  OR3_X1    g0451(.A1(new_n364), .A2(KEYINPUT27), .A3(G20), .ZN(new_n652));
  OAI21_X1  g0452(.A(KEYINPUT27), .B1(new_n364), .B2(G20), .ZN(new_n653));
  AND3_X1   g0453(.A1(new_n652), .A2(G213), .A3(new_n653), .ZN(new_n654));
  INV_X1    g0454(.A(new_n654), .ZN(new_n655));
  INV_X1    g0455(.A(G343), .ZN(new_n656));
  NOR2_X1   g0456(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  INV_X1    g0457(.A(new_n657), .ZN(new_n658));
  NOR2_X1   g0458(.A1(new_n658), .A2(new_n522), .ZN(new_n659));
  XNOR2_X1  g0459(.A(new_n481), .B(new_n659), .ZN(new_n660));
  NAND3_X1  g0460(.A1(new_n660), .A2(G330), .A3(new_n524), .ZN(new_n661));
  NOR2_X1   g0461(.A1(new_n521), .A2(new_n657), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n505), .A2(new_n657), .ZN(new_n663));
  AOI21_X1  g0463(.A(new_n520), .B1(new_n528), .B2(new_n663), .ZN(new_n664));
  NOR2_X1   g0464(.A1(new_n662), .A2(new_n664), .ZN(new_n665));
  INV_X1    g0465(.A(new_n665), .ZN(new_n666));
  NOR2_X1   g0466(.A1(new_n661), .A2(new_n666), .ZN(new_n667));
  INV_X1    g0467(.A(new_n667), .ZN(new_n668));
  NOR2_X1   g0468(.A1(new_n482), .A2(new_n657), .ZN(new_n669));
  AOI21_X1  g0469(.A(new_n662), .B1(new_n665), .B2(new_n669), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n668), .A2(new_n670), .ZN(new_n671));
  XNOR2_X1  g0471(.A(new_n671), .B(KEYINPUT94), .ZN(G399));
  NOR2_X1   g0472(.A1(new_n235), .A2(G41), .ZN(new_n673));
  INV_X1    g0473(.A(new_n673), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n674), .A2(G1), .ZN(new_n675));
  NAND3_X1  g0475(.A1(new_n557), .A2(new_n207), .A3(new_n218), .ZN(new_n676));
  OAI22_X1  g0476(.A1(new_n675), .A2(new_n676), .B1(new_n231), .B2(new_n674), .ZN(new_n677));
  XNOR2_X1  g0477(.A(new_n677), .B(KEYINPUT28), .ZN(new_n678));
  INV_X1    g0478(.A(new_n570), .ZN(new_n679));
  NAND3_X1  g0479(.A1(new_n621), .A2(new_n642), .A3(new_n679), .ZN(new_n680));
  INV_X1    g0480(.A(new_n644), .ZN(new_n681));
  OAI21_X1  g0481(.A(KEYINPUT26), .B1(new_n681), .B2(new_n570), .ZN(new_n682));
  OAI211_X1 g0482(.A(new_n680), .B(new_n682), .C1(new_n648), .C2(new_n647), .ZN(new_n683));
  XOR2_X1   g0483(.A(new_n620), .B(KEYINPUT98), .Z(new_n684));
  OAI21_X1  g0484(.A(new_n658), .B1(new_n683), .B2(new_n684), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n685), .A2(KEYINPUT29), .ZN(new_n686));
  NOR2_X1   g0486(.A1(new_n650), .A2(new_n657), .ZN(new_n687));
  INV_X1    g0487(.A(new_n687), .ZN(new_n688));
  OAI21_X1  g0488(.A(new_n686), .B1(new_n688), .B2(KEYINPUT29), .ZN(new_n689));
  INV_X1    g0489(.A(new_n529), .ZN(new_n690));
  AND3_X1   g0490(.A1(new_n570), .A2(new_n574), .A3(new_n622), .ZN(new_n691));
  AOI21_X1  g0491(.A(new_n622), .B1(new_n570), .B2(new_n574), .ZN(new_n692));
  NOR2_X1   g0492(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  AOI21_X1  g0493(.A(KEYINPUT91), .B1(new_n693), .B2(new_n621), .ZN(new_n694));
  INV_X1    g0494(.A(new_n627), .ZN(new_n695));
  OAI211_X1 g0495(.A(new_n690), .B(new_n658), .C1(new_n694), .C2(new_n695), .ZN(new_n696));
  NOR2_X1   g0496(.A1(new_n550), .A2(new_n476), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n697), .A2(new_n517), .ZN(new_n698));
  OAI21_X1  g0498(.A(KEYINPUT96), .B1(new_n698), .B2(new_n616), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n699), .A2(KEYINPUT30), .ZN(new_n700));
  NAND3_X1  g0500(.A1(new_n616), .A2(new_n467), .A3(new_n319), .ZN(new_n701));
  OR2_X1    g0501(.A1(new_n701), .A2(KEYINPUT97), .ZN(new_n702));
  NAND2_X1  g0502(.A1(new_n701), .A2(KEYINPUT97), .ZN(new_n703));
  NAND4_X1  g0503(.A1(new_n702), .A2(new_n550), .A3(new_n512), .A4(new_n703), .ZN(new_n704));
  INV_X1    g0504(.A(KEYINPUT30), .ZN(new_n705));
  OAI211_X1 g0505(.A(KEYINPUT96), .B(new_n705), .C1(new_n698), .C2(new_n616), .ZN(new_n706));
  NAND3_X1  g0506(.A1(new_n700), .A2(new_n704), .A3(new_n706), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n707), .A2(new_n657), .ZN(new_n708));
  INV_X1    g0508(.A(KEYINPUT31), .ZN(new_n709));
  NAND2_X1  g0509(.A1(new_n708), .A2(new_n709), .ZN(new_n710));
  XNOR2_X1  g0510(.A(KEYINPUT95), .B(KEYINPUT31), .ZN(new_n711));
  NAND3_X1  g0511(.A1(new_n707), .A2(new_n657), .A3(new_n711), .ZN(new_n712));
  NAND3_X1  g0512(.A1(new_n696), .A2(new_n710), .A3(new_n712), .ZN(new_n713));
  AOI21_X1  g0513(.A(new_n689), .B1(G330), .B2(new_n713), .ZN(new_n714));
  OAI21_X1  g0514(.A(new_n678), .B1(new_n714), .B2(G1), .ZN(G364));
  NAND3_X1  g0515(.A1(new_n236), .A2(G355), .A3(new_n283), .ZN(new_n716));
  INV_X1    g0516(.A(G45), .ZN(new_n717));
  NOR2_X1   g0517(.A1(new_n251), .A2(new_n717), .ZN(new_n718));
  NOR2_X1   g0518(.A1(new_n235), .A2(new_n283), .ZN(new_n719));
  OAI21_X1  g0519(.A(new_n719), .B1(G45), .B2(new_n231), .ZN(new_n720));
  OAI221_X1 g0520(.A(new_n716), .B1(G116), .B2(new_n236), .C1(new_n718), .C2(new_n720), .ZN(new_n721));
  NOR2_X1   g0521(.A1(G13), .A2(G33), .ZN(new_n722));
  INV_X1    g0522(.A(new_n722), .ZN(new_n723));
  NOR2_X1   g0523(.A1(new_n723), .A2(G20), .ZN(new_n724));
  AOI21_X1  g0524(.A(new_n232), .B1(G20), .B2(new_n298), .ZN(new_n725));
  NOR2_X1   g0525(.A1(new_n724), .A2(new_n725), .ZN(new_n726));
  NAND2_X1  g0526(.A1(new_n721), .A2(new_n726), .ZN(new_n727));
  NOR2_X1   g0527(.A1(new_n234), .A2(G20), .ZN(new_n728));
  NAND2_X1  g0528(.A1(new_n728), .A2(G45), .ZN(new_n729));
  NAND3_X1  g0529(.A1(new_n674), .A2(G1), .A3(new_n729), .ZN(new_n730));
  INV_X1    g0530(.A(new_n730), .ZN(new_n731));
  NOR2_X1   g0531(.A1(new_n223), .A2(new_n319), .ZN(new_n732));
  OR2_X1    g0532(.A1(new_n732), .A2(KEYINPUT100), .ZN(new_n733));
  NAND2_X1  g0533(.A1(new_n732), .A2(KEYINPUT100), .ZN(new_n734));
  NOR2_X1   g0534(.A1(new_n330), .A2(G200), .ZN(new_n735));
  NAND3_X1  g0535(.A1(new_n733), .A2(new_n734), .A3(new_n735), .ZN(new_n736));
  INV_X1    g0536(.A(new_n736), .ZN(new_n737));
  INV_X1    g0537(.A(new_n388), .ZN(new_n738));
  NAND2_X1  g0538(.A1(new_n732), .A2(G200), .ZN(new_n739));
  NOR2_X1   g0539(.A1(new_n739), .A2(G190), .ZN(new_n740));
  AOI22_X1  g0540(.A1(new_n737), .A2(new_n738), .B1(G68), .B2(new_n740), .ZN(new_n741));
  NOR2_X1   g0541(.A1(G190), .A2(G200), .ZN(new_n742));
  NAND3_X1  g0542(.A1(new_n733), .A2(new_n742), .A3(new_n734), .ZN(new_n743));
  OAI21_X1  g0543(.A(new_n741), .B1(new_n309), .B2(new_n743), .ZN(new_n744));
  INV_X1    g0544(.A(new_n744), .ZN(new_n745));
  NOR2_X1   g0545(.A1(new_n223), .A2(G179), .ZN(new_n746));
  NAND3_X1  g0546(.A1(new_n746), .A2(G190), .A3(G200), .ZN(new_n747));
  INV_X1    g0547(.A(new_n747), .ZN(new_n748));
  AOI21_X1  g0548(.A(new_n448), .B1(new_n748), .B2(G87), .ZN(new_n749));
  NAND3_X1  g0549(.A1(new_n746), .A2(new_n330), .A3(G200), .ZN(new_n750));
  NOR2_X1   g0550(.A1(new_n750), .A2(new_n555), .ZN(new_n751));
  NAND2_X1  g0551(.A1(new_n735), .A2(new_n319), .ZN(new_n752));
  NAND2_X1  g0552(.A1(new_n752), .A2(G20), .ZN(new_n753));
  INV_X1    g0553(.A(new_n753), .ZN(new_n754));
  NOR2_X1   g0554(.A1(new_n754), .A2(new_n209), .ZN(new_n755));
  NOR2_X1   g0555(.A1(new_n739), .A2(new_n330), .ZN(new_n756));
  AOI211_X1 g0556(.A(new_n751), .B(new_n755), .C1(G50), .C2(new_n756), .ZN(new_n757));
  NAND2_X1  g0557(.A1(new_n746), .A2(new_n742), .ZN(new_n758));
  INV_X1    g0558(.A(G159), .ZN(new_n759));
  NOR2_X1   g0559(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  XNOR2_X1  g0560(.A(new_n760), .B(KEYINPUT32), .ZN(new_n761));
  NAND4_X1  g0561(.A1(new_n745), .A2(new_n749), .A3(new_n757), .A4(new_n761), .ZN(new_n762));
  XOR2_X1   g0562(.A(new_n758), .B(KEYINPUT101), .Z(new_n763));
  INV_X1    g0563(.A(G329), .ZN(new_n764));
  INV_X1    g0564(.A(G326), .ZN(new_n765));
  INV_X1    g0565(.A(new_n756), .ZN(new_n766));
  OAI22_X1  g0566(.A1(new_n763), .A2(new_n764), .B1(new_n765), .B2(new_n766), .ZN(new_n767));
  AOI21_X1  g0567(.A(new_n767), .B1(G294), .B2(new_n753), .ZN(new_n768));
  INV_X1    g0568(.A(G283), .ZN(new_n769));
  OAI221_X1 g0569(.A(new_n448), .B1(new_n747), .B2(new_n449), .C1(new_n769), .C2(new_n750), .ZN(new_n770));
  XNOR2_X1  g0570(.A(KEYINPUT33), .B(G317), .ZN(new_n771));
  AOI21_X1  g0571(.A(new_n770), .B1(new_n740), .B2(new_n771), .ZN(new_n772));
  INV_X1    g0572(.A(G322), .ZN(new_n773));
  OAI211_X1 g0573(.A(new_n768), .B(new_n772), .C1(new_n773), .C2(new_n736), .ZN(new_n774));
  INV_X1    g0574(.A(G311), .ZN(new_n775));
  NOR2_X1   g0575(.A1(new_n743), .A2(new_n775), .ZN(new_n776));
  OAI21_X1  g0576(.A(new_n762), .B1(new_n774), .B2(new_n776), .ZN(new_n777));
  NAND2_X1  g0577(.A1(new_n777), .A2(new_n725), .ZN(new_n778));
  NAND3_X1  g0578(.A1(new_n727), .A2(new_n731), .A3(new_n778), .ZN(new_n779));
  XOR2_X1   g0579(.A(new_n779), .B(KEYINPUT102), .Z(new_n780));
  NAND2_X1  g0580(.A1(new_n660), .A2(new_n524), .ZN(new_n781));
  AOI21_X1  g0581(.A(new_n780), .B1(new_n781), .B2(new_n724), .ZN(new_n782));
  INV_X1    g0582(.A(G330), .ZN(new_n783));
  NAND2_X1  g0583(.A1(new_n781), .A2(new_n783), .ZN(new_n784));
  INV_X1    g0584(.A(KEYINPUT99), .ZN(new_n785));
  XNOR2_X1  g0585(.A(new_n661), .B(new_n785), .ZN(new_n786));
  NOR2_X1   g0586(.A1(new_n786), .A2(new_n731), .ZN(new_n787));
  AOI21_X1  g0587(.A(new_n782), .B1(new_n784), .B2(new_n787), .ZN(new_n788));
  INV_X1    g0588(.A(new_n788), .ZN(G396));
  AOI22_X1  g0589(.A1(new_n740), .A2(G150), .B1(new_n756), .B2(G137), .ZN(new_n790));
  XOR2_X1   g0590(.A(new_n790), .B(KEYINPUT106), .Z(new_n791));
  INV_X1    g0591(.A(G143), .ZN(new_n792));
  OAI221_X1 g0592(.A(new_n791), .B1(new_n792), .B2(new_n736), .C1(new_n759), .C2(new_n743), .ZN(new_n793));
  XOR2_X1   g0593(.A(new_n793), .B(KEYINPUT34), .Z(new_n794));
  AOI21_X1  g0594(.A(new_n794), .B1(G50), .B2(new_n748), .ZN(new_n795));
  AOI21_X1  g0595(.A(new_n448), .B1(new_n753), .B2(new_n738), .ZN(new_n796));
  INV_X1    g0596(.A(new_n763), .ZN(new_n797));
  NAND2_X1  g0597(.A1(new_n797), .A2(G132), .ZN(new_n798));
  NOR2_X1   g0598(.A1(new_n750), .A2(new_n216), .ZN(new_n799));
  INV_X1    g0599(.A(new_n799), .ZN(new_n800));
  NAND4_X1  g0600(.A1(new_n795), .A2(new_n796), .A3(new_n798), .A4(new_n800), .ZN(new_n801));
  INV_X1    g0601(.A(new_n740), .ZN(new_n802));
  OAI22_X1  g0602(.A1(new_n802), .A2(new_n769), .B1(new_n750), .B2(new_n207), .ZN(new_n803));
  AOI21_X1  g0603(.A(new_n755), .B1(G294), .B2(new_n737), .ZN(new_n804));
  XOR2_X1   g0604(.A(new_n804), .B(KEYINPUT105), .Z(new_n805));
  AOI211_X1 g0605(.A(new_n803), .B(new_n805), .C1(G303), .C2(new_n756), .ZN(new_n806));
  INV_X1    g0606(.A(new_n743), .ZN(new_n807));
  NAND2_X1  g0607(.A1(new_n807), .A2(G116), .ZN(new_n808));
  NAND2_X1  g0608(.A1(new_n797), .A2(G311), .ZN(new_n809));
  OAI21_X1  g0609(.A(new_n448), .B1(new_n747), .B2(new_n555), .ZN(new_n810));
  XOR2_X1   g0610(.A(new_n810), .B(KEYINPUT104), .Z(new_n811));
  NAND4_X1  g0611(.A1(new_n806), .A2(new_n808), .A3(new_n809), .A4(new_n811), .ZN(new_n812));
  AND2_X1   g0612(.A1(new_n801), .A2(new_n812), .ZN(new_n813));
  INV_X1    g0613(.A(new_n725), .ZN(new_n814));
  OAI21_X1  g0614(.A(new_n731), .B1(new_n813), .B2(new_n814), .ZN(new_n815));
  NOR2_X1   g0615(.A1(new_n725), .A2(new_n722), .ZN(new_n816));
  XOR2_X1   g0616(.A(new_n816), .B(KEYINPUT103), .Z(new_n817));
  AOI21_X1  g0617(.A(new_n815), .B1(new_n309), .B2(new_n817), .ZN(new_n818));
  XNOR2_X1  g0618(.A(new_n818), .B(KEYINPUT107), .ZN(new_n819));
  XNOR2_X1  g0619(.A(new_n321), .B(KEYINPUT108), .ZN(new_n820));
  NOR2_X1   g0620(.A1(new_n820), .A2(new_n427), .ZN(new_n821));
  INV_X1    g0621(.A(new_n311), .ZN(new_n822));
  OAI21_X1  g0622(.A(new_n821), .B1(new_n822), .B2(new_n658), .ZN(new_n823));
  OR2_X1    g0623(.A1(new_n321), .A2(new_n658), .ZN(new_n824));
  NAND2_X1  g0624(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  OAI21_X1  g0625(.A(new_n819), .B1(new_n723), .B2(new_n825), .ZN(new_n826));
  NAND2_X1  g0626(.A1(new_n713), .A2(G330), .ZN(new_n827));
  OAI211_X1 g0627(.A(new_n658), .B(new_n821), .C1(new_n646), .C2(new_n649), .ZN(new_n828));
  OAI21_X1  g0628(.A(new_n828), .B1(new_n687), .B2(new_n825), .ZN(new_n829));
  XOR2_X1   g0629(.A(new_n827), .B(new_n829), .Z(new_n830));
  NAND2_X1  g0630(.A1(new_n830), .A2(new_n730), .ZN(new_n831));
  AND2_X1   g0631(.A1(new_n826), .A2(new_n831), .ZN(new_n832));
  INV_X1    g0632(.A(new_n832), .ZN(G384));
  INV_X1    g0633(.A(KEYINPUT39), .ZN(new_n834));
  OAI21_X1  g0634(.A(new_n390), .B1(new_n396), .B2(new_n398), .ZN(new_n835));
  NAND2_X1  g0635(.A1(new_n835), .A2(new_n402), .ZN(new_n836));
  NAND3_X1  g0636(.A1(new_n836), .A2(new_n399), .A3(new_n271), .ZN(new_n837));
  AOI21_X1  g0637(.A(new_n655), .B1(new_n837), .B2(new_n406), .ZN(new_n838));
  OAI21_X1  g0638(.A(new_n838), .B1(new_n411), .B2(new_n420), .ZN(new_n839));
  AND3_X1   g0639(.A1(new_n383), .A2(G179), .A3(new_n384), .ZN(new_n840));
  AOI21_X1  g0640(.A(new_n298), .B1(new_n383), .B2(new_n384), .ZN(new_n841));
  NOR3_X1   g0641(.A1(new_n840), .A2(new_n841), .A3(new_n654), .ZN(new_n842));
  AOI21_X1  g0642(.A(new_n842), .B1(new_n837), .B2(new_n406), .ZN(new_n843));
  AND4_X1   g0643(.A1(new_n404), .A2(new_n406), .A3(new_n412), .A4(new_n413), .ZN(new_n844));
  OAI21_X1  g0644(.A(KEYINPUT37), .B1(new_n843), .B2(new_n844), .ZN(new_n845));
  NAND2_X1  g0645(.A1(new_n408), .A2(new_n654), .ZN(new_n846));
  INV_X1    g0646(.A(KEYINPUT109), .ZN(new_n847));
  AOI22_X1  g0647(.A1(new_n404), .A2(new_n406), .B1(new_n386), .B2(new_n387), .ZN(new_n848));
  OAI211_X1 g0648(.A(new_n846), .B(new_n414), .C1(new_n847), .C2(new_n848), .ZN(new_n849));
  INV_X1    g0649(.A(KEYINPUT37), .ZN(new_n850));
  NAND2_X1  g0650(.A1(new_n408), .A2(new_n409), .ZN(new_n851));
  OAI21_X1  g0651(.A(new_n850), .B1(new_n851), .B2(KEYINPUT109), .ZN(new_n852));
  OAI21_X1  g0652(.A(new_n845), .B1(new_n849), .B2(new_n852), .ZN(new_n853));
  AND3_X1   g0653(.A1(new_n839), .A2(KEYINPUT38), .A3(new_n853), .ZN(new_n854));
  INV_X1    g0654(.A(new_n854), .ZN(new_n855));
  AOI21_X1  g0655(.A(new_n655), .B1(new_n404), .B2(new_n406), .ZN(new_n856));
  NOR2_X1   g0656(.A1(new_n844), .A2(new_n856), .ZN(new_n857));
  AOI21_X1  g0657(.A(KEYINPUT37), .B1(new_n848), .B2(new_n847), .ZN(new_n858));
  NAND2_X1  g0658(.A1(new_n851), .A2(KEYINPUT109), .ZN(new_n859));
  NAND3_X1  g0659(.A1(new_n857), .A2(new_n858), .A3(new_n859), .ZN(new_n860));
  NAND3_X1  g0660(.A1(new_n851), .A2(new_n846), .A3(new_n414), .ZN(new_n861));
  NAND2_X1  g0661(.A1(new_n861), .A2(KEYINPUT37), .ZN(new_n862));
  INV_X1    g0662(.A(KEYINPUT112), .ZN(new_n863));
  AND3_X1   g0663(.A1(new_n860), .A2(new_n862), .A3(new_n863), .ZN(new_n864));
  AOI21_X1  g0664(.A(new_n863), .B1(new_n860), .B2(new_n862), .ZN(new_n865));
  OR2_X1    g0665(.A1(new_n407), .A2(new_n410), .ZN(new_n866));
  AOI21_X1  g0666(.A(new_n846), .B1(new_n866), .B2(new_n632), .ZN(new_n867));
  NOR3_X1   g0667(.A1(new_n864), .A2(new_n865), .A3(new_n867), .ZN(new_n868));
  XOR2_X1   g0668(.A(KEYINPUT111), .B(KEYINPUT38), .Z(new_n869));
  INV_X1    g0669(.A(new_n869), .ZN(new_n870));
  OAI211_X1 g0670(.A(new_n834), .B(new_n855), .C1(new_n868), .C2(new_n870), .ZN(new_n871));
  AOI21_X1  g0671(.A(KEYINPUT38), .B1(new_n839), .B2(new_n853), .ZN(new_n872));
  OAI21_X1  g0672(.A(KEYINPUT39), .B1(new_n854), .B2(new_n872), .ZN(new_n873));
  NAND2_X1  g0673(.A1(new_n873), .A2(KEYINPUT110), .ZN(new_n874));
  INV_X1    g0674(.A(KEYINPUT110), .ZN(new_n875));
  OAI211_X1 g0675(.A(new_n875), .B(KEYINPUT39), .C1(new_n854), .C2(new_n872), .ZN(new_n876));
  NAND3_X1  g0676(.A1(new_n871), .A2(new_n874), .A3(new_n876), .ZN(new_n877));
  NAND3_X1  g0677(.A1(new_n357), .A2(new_n370), .A3(new_n658), .ZN(new_n878));
  INV_X1    g0678(.A(new_n878), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n877), .A2(new_n879), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n820), .A2(new_n658), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n828), .A2(new_n881), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n370), .A2(new_n657), .ZN(new_n883));
  NAND3_X1  g0683(.A1(new_n371), .A2(new_n424), .A3(new_n883), .ZN(new_n884));
  OAI211_X1 g0684(.A(new_n370), .B(new_n657), .C1(new_n630), .C2(new_n357), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n884), .A2(new_n885), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n882), .A2(new_n886), .ZN(new_n887));
  INV_X1    g0687(.A(new_n887), .ZN(new_n888));
  OR2_X1    g0688(.A1(new_n854), .A2(new_n872), .ZN(new_n889));
  AOI22_X1  g0689(.A1(new_n888), .A2(new_n889), .B1(new_n411), .B2(new_n655), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n880), .A2(new_n890), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n891), .A2(KEYINPUT113), .ZN(new_n892));
  INV_X1    g0692(.A(KEYINPUT113), .ZN(new_n893));
  NAND3_X1  g0693(.A1(new_n880), .A2(new_n893), .A3(new_n890), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n892), .A2(new_n894), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n689), .A2(new_n430), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n635), .A2(new_n896), .ZN(new_n897));
  XNOR2_X1  g0697(.A(new_n895), .B(new_n897), .ZN(new_n898));
  INV_X1    g0698(.A(KEYINPUT40), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n886), .A2(new_n825), .ZN(new_n900));
  INV_X1    g0700(.A(new_n711), .ZN(new_n901));
  AOI22_X1  g0701(.A1(new_n628), .A2(new_n658), .B1(new_n708), .B2(new_n901), .ZN(new_n902));
  NAND3_X1  g0702(.A1(new_n707), .A2(KEYINPUT31), .A3(new_n657), .ZN(new_n903));
  AOI21_X1  g0703(.A(new_n900), .B1(new_n902), .B2(new_n903), .ZN(new_n904));
  OAI21_X1  g0704(.A(new_n855), .B1(new_n868), .B2(new_n870), .ZN(new_n905));
  AOI21_X1  g0705(.A(new_n899), .B1(new_n904), .B2(new_n905), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n708), .A2(new_n901), .ZN(new_n907));
  NAND3_X1  g0707(.A1(new_n696), .A2(new_n903), .A3(new_n907), .ZN(new_n908));
  INV_X1    g0708(.A(new_n900), .ZN(new_n909));
  AND4_X1   g0709(.A1(new_n899), .A2(new_n908), .A3(new_n909), .A4(new_n889), .ZN(new_n910));
  NOR2_X1   g0710(.A1(new_n906), .A2(new_n910), .ZN(new_n911));
  AND2_X1   g0711(.A1(new_n908), .A2(new_n430), .ZN(new_n912));
  XNOR2_X1  g0712(.A(new_n911), .B(new_n912), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n913), .A2(G330), .ZN(new_n914));
  XNOR2_X1  g0714(.A(new_n898), .B(new_n914), .ZN(new_n915));
  OAI21_X1  g0715(.A(new_n915), .B1(new_n222), .B2(new_n728), .ZN(new_n916));
  INV_X1    g0716(.A(KEYINPUT35), .ZN(new_n917));
  AOI211_X1 g0717(.A(new_n223), .B(new_n232), .C1(new_n560), .C2(new_n917), .ZN(new_n918));
  OAI211_X1 g0718(.A(new_n918), .B(G116), .C1(new_n917), .C2(new_n560), .ZN(new_n919));
  XNOR2_X1  g0719(.A(new_n919), .B(KEYINPUT36), .ZN(new_n920));
  AOI211_X1 g0720(.A(new_n309), .B(new_n231), .C1(new_n738), .C2(G68), .ZN(new_n921));
  NOR2_X1   g0721(.A1(new_n216), .A2(G50), .ZN(new_n922));
  OAI211_X1 g0722(.A(G1), .B(new_n234), .C1(new_n921), .C2(new_n922), .ZN(new_n923));
  NAND3_X1  g0723(.A1(new_n916), .A2(new_n920), .A3(new_n923), .ZN(G367));
  AOI21_X1  g0724(.A(KEYINPUT116), .B1(new_n748), .B2(G116), .ZN(new_n925));
  XOR2_X1   g0725(.A(new_n925), .B(KEYINPUT46), .Z(new_n926));
  INV_X1    g0726(.A(new_n758), .ZN(new_n927));
  AOI22_X1  g0727(.A1(new_n756), .A2(G311), .B1(G317), .B2(new_n927), .ZN(new_n928));
  OAI221_X1 g0728(.A(new_n928), .B1(new_n209), .B2(new_n750), .C1(new_n555), .C2(new_n754), .ZN(new_n929));
  INV_X1    g0729(.A(G294), .ZN(new_n930));
  OAI221_X1 g0730(.A(new_n448), .B1(new_n802), .B2(new_n930), .C1(new_n449), .C2(new_n736), .ZN(new_n931));
  NOR2_X1   g0731(.A1(new_n743), .A2(new_n769), .ZN(new_n932));
  NOR4_X1   g0732(.A1(new_n926), .A2(new_n929), .A3(new_n931), .A4(new_n932), .ZN(new_n933));
  NOR2_X1   g0733(.A1(new_n754), .A2(new_n216), .ZN(new_n934));
  INV_X1    g0734(.A(new_n934), .ZN(new_n935));
  INV_X1    g0735(.A(G150), .ZN(new_n936));
  OAI221_X1 g0736(.A(new_n935), .B1(new_n792), .B2(new_n766), .C1(new_n936), .C2(new_n736), .ZN(new_n937));
  OR2_X1    g0737(.A1(new_n937), .A2(KEYINPUT117), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n927), .A2(G137), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n937), .A2(KEYINPUT117), .ZN(new_n940));
  NOR2_X1   g0740(.A1(new_n750), .A2(new_n309), .ZN(new_n941));
  AOI211_X1 g0741(.A(new_n448), .B(new_n941), .C1(G159), .C2(new_n740), .ZN(new_n942));
  NAND4_X1  g0742(.A1(new_n938), .A2(new_n939), .A3(new_n940), .A4(new_n942), .ZN(new_n943));
  AOI21_X1  g0743(.A(new_n943), .B1(G50), .B2(new_n807), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n748), .A2(new_n738), .ZN(new_n945));
  AOI21_X1  g0745(.A(new_n933), .B1(new_n944), .B2(new_n945), .ZN(new_n946));
  XOR2_X1   g0746(.A(new_n946), .B(KEYINPUT47), .Z(new_n947));
  NAND2_X1  g0747(.A1(new_n947), .A2(new_n725), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n606), .A2(new_n657), .ZN(new_n949));
  NOR2_X1   g0749(.A1(new_n620), .A2(new_n949), .ZN(new_n950));
  AOI21_X1  g0750(.A(new_n950), .B1(new_n644), .B2(new_n949), .ZN(new_n951));
  INV_X1    g0751(.A(KEYINPUT114), .ZN(new_n952));
  NOR2_X1   g0752(.A1(new_n951), .A2(new_n952), .ZN(new_n953));
  NOR2_X1   g0753(.A1(new_n950), .A2(KEYINPUT114), .ZN(new_n954));
  NOR2_X1   g0754(.A1(new_n953), .A2(new_n954), .ZN(new_n955));
  NAND2_X1  g0755(.A1(new_n955), .A2(new_n724), .ZN(new_n956));
  INV_X1    g0756(.A(new_n719), .ZN(new_n957));
  OAI221_X1 g0757(.A(new_n726), .B1(new_n236), .B2(new_n305), .C1(new_n246), .C2(new_n957), .ZN(new_n958));
  NAND4_X1  g0758(.A1(new_n948), .A2(new_n731), .A3(new_n956), .A4(new_n958), .ZN(new_n959));
  NAND2_X1  g0759(.A1(new_n729), .A2(G1), .ZN(new_n960));
  NAND2_X1  g0760(.A1(new_n679), .A2(new_n657), .ZN(new_n961));
  OAI211_X1 g0761(.A(new_n570), .B(new_n574), .C1(new_n572), .C2(new_n658), .ZN(new_n962));
  NAND2_X1  g0762(.A1(new_n961), .A2(new_n962), .ZN(new_n963));
  NOR2_X1   g0763(.A1(new_n670), .A2(new_n963), .ZN(new_n964));
  XOR2_X1   g0764(.A(new_n964), .B(KEYINPUT44), .Z(new_n965));
  NAND2_X1  g0765(.A1(new_n670), .A2(new_n963), .ZN(new_n966));
  XNOR2_X1  g0766(.A(new_n966), .B(KEYINPUT45), .ZN(new_n967));
  NOR2_X1   g0767(.A1(new_n965), .A2(new_n967), .ZN(new_n968));
  XNOR2_X1  g0768(.A(new_n968), .B(new_n668), .ZN(new_n969));
  XOR2_X1   g0769(.A(new_n665), .B(new_n669), .Z(new_n970));
  INV_X1    g0770(.A(KEYINPUT115), .ZN(new_n971));
  OAI211_X1 g0771(.A(new_n970), .B(new_n661), .C1(new_n785), .C2(new_n971), .ZN(new_n972));
  NOR2_X1   g0772(.A1(new_n786), .A2(KEYINPUT115), .ZN(new_n973));
  OAI21_X1  g0773(.A(new_n972), .B1(new_n973), .B2(new_n970), .ZN(new_n974));
  NAND2_X1  g0774(.A1(new_n714), .A2(new_n974), .ZN(new_n975));
  OR2_X1    g0775(.A1(new_n969), .A2(new_n975), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n976), .A2(new_n714), .ZN(new_n977));
  XNOR2_X1  g0777(.A(new_n673), .B(KEYINPUT41), .ZN(new_n978));
  AOI21_X1  g0778(.A(new_n960), .B1(new_n977), .B2(new_n978), .ZN(new_n979));
  INV_X1    g0779(.A(new_n955), .ZN(new_n980));
  NAND2_X1  g0780(.A1(new_n980), .A2(KEYINPUT43), .ZN(new_n981));
  NAND3_X1  g0781(.A1(new_n665), .A2(new_n669), .A3(new_n963), .ZN(new_n982));
  XNOR2_X1  g0782(.A(new_n982), .B(KEYINPUT42), .ZN(new_n983));
  OAI21_X1  g0783(.A(new_n570), .B1(new_n962), .B2(new_n521), .ZN(new_n984));
  AND2_X1   g0784(.A1(new_n984), .A2(new_n658), .ZN(new_n985));
  OAI21_X1  g0785(.A(new_n981), .B1(new_n983), .B2(new_n985), .ZN(new_n986));
  INV_X1    g0786(.A(new_n963), .ZN(new_n987));
  NOR2_X1   g0787(.A1(new_n668), .A2(new_n987), .ZN(new_n988));
  XNOR2_X1  g0788(.A(new_n986), .B(new_n988), .ZN(new_n989));
  NOR2_X1   g0789(.A1(new_n980), .A2(KEYINPUT43), .ZN(new_n990));
  XOR2_X1   g0790(.A(new_n989), .B(new_n990), .Z(new_n991));
  OAI21_X1  g0791(.A(new_n959), .B1(new_n979), .B2(new_n991), .ZN(G387));
  NAND2_X1  g0792(.A1(new_n975), .A2(new_n673), .ZN(new_n993));
  XOR2_X1   g0793(.A(new_n993), .B(KEYINPUT119), .Z(new_n994));
  OAI21_X1  g0794(.A(new_n994), .B1(new_n714), .B2(new_n974), .ZN(new_n995));
  OAI21_X1  g0795(.A(new_n448), .B1(new_n758), .B2(new_n765), .ZN(new_n996));
  AOI22_X1  g0796(.A1(new_n737), .A2(G317), .B1(G311), .B2(new_n740), .ZN(new_n997));
  OAI221_X1 g0797(.A(new_n997), .B1(new_n449), .B2(new_n743), .C1(new_n773), .C2(new_n766), .ZN(new_n998));
  XNOR2_X1  g0798(.A(new_n998), .B(KEYINPUT48), .ZN(new_n999));
  OAI221_X1 g0799(.A(new_n999), .B1(new_n769), .B2(new_n754), .C1(new_n930), .C2(new_n747), .ZN(new_n1000));
  XOR2_X1   g0800(.A(new_n1000), .B(KEYINPUT49), .Z(new_n1001));
  INV_X1    g0801(.A(new_n750), .ZN(new_n1002));
  AOI211_X1 g0802(.A(new_n996), .B(new_n1001), .C1(G116), .C2(new_n1002), .ZN(new_n1003));
  NOR2_X1   g0803(.A1(new_n736), .A2(new_n212), .ZN(new_n1004));
  NAND2_X1  g0804(.A1(new_n753), .A2(new_n304), .ZN(new_n1005));
  OAI221_X1 g0805(.A(new_n1005), .B1(new_n766), .B2(new_n759), .C1(new_n216), .C2(new_n743), .ZN(new_n1006));
  AOI211_X1 g0806(.A(new_n1004), .B(new_n1006), .C1(G150), .C2(new_n927), .ZN(new_n1007));
  OAI221_X1 g0807(.A(new_n1007), .B1(new_n309), .B2(new_n747), .C1(new_n264), .C2(new_n802), .ZN(new_n1008));
  AOI211_X1 g0808(.A(new_n448), .B(new_n1008), .C1(G97), .C2(new_n1002), .ZN(new_n1009));
  OAI21_X1  g0809(.A(new_n725), .B1(new_n1003), .B2(new_n1009), .ZN(new_n1010));
  NAND2_X1  g0810(.A1(new_n302), .A2(new_n212), .ZN(new_n1011));
  XNOR2_X1  g0811(.A(new_n1011), .B(KEYINPUT50), .ZN(new_n1012));
  NOR2_X1   g0812(.A1(new_n216), .A2(new_n309), .ZN(new_n1013));
  NOR4_X1   g0813(.A1(new_n1012), .A2(G45), .A3(new_n1013), .A4(new_n676), .ZN(new_n1014));
  OAI21_X1  g0814(.A(new_n719), .B1(new_n243), .B2(new_n717), .ZN(new_n1015));
  NAND3_X1  g0815(.A1(new_n236), .A2(new_n283), .A3(new_n676), .ZN(new_n1016));
  AOI21_X1  g0816(.A(new_n1014), .B1(new_n1015), .B2(new_n1016), .ZN(new_n1017));
  NOR2_X1   g0817(.A1(new_n236), .A2(G107), .ZN(new_n1018));
  OAI21_X1  g0818(.A(new_n726), .B1(new_n1017), .B2(new_n1018), .ZN(new_n1019));
  AOI21_X1  g0819(.A(new_n730), .B1(new_n666), .B2(new_n724), .ZN(new_n1020));
  NAND3_X1  g0820(.A1(new_n1010), .A2(new_n1019), .A3(new_n1020), .ZN(new_n1021));
  XNOR2_X1  g0821(.A(new_n1021), .B(KEYINPUT118), .ZN(new_n1022));
  NAND2_X1  g0822(.A1(new_n974), .A2(new_n960), .ZN(new_n1023));
  NAND3_X1  g0823(.A1(new_n995), .A2(new_n1022), .A3(new_n1023), .ZN(G393));
  AOI21_X1  g0824(.A(new_n674), .B1(new_n969), .B2(new_n975), .ZN(new_n1025));
  NAND2_X1  g0825(.A1(new_n976), .A2(new_n1025), .ZN(new_n1026));
  AOI22_X1  g0826(.A1(new_n737), .A2(G311), .B1(G317), .B2(new_n756), .ZN(new_n1027));
  XNOR2_X1  g0827(.A(new_n1027), .B(KEYINPUT121), .ZN(new_n1028));
  XOR2_X1   g0828(.A(new_n1028), .B(KEYINPUT52), .Z(new_n1029));
  OAI21_X1  g0829(.A(new_n448), .B1(new_n743), .B2(new_n930), .ZN(new_n1030));
  NOR2_X1   g0830(.A1(new_n747), .A2(new_n769), .ZN(new_n1031));
  NOR4_X1   g0831(.A1(new_n1029), .A2(new_n751), .A3(new_n1030), .A4(new_n1031), .ZN(new_n1032));
  OAI221_X1 g0832(.A(new_n1032), .B1(new_n218), .B2(new_n754), .C1(new_n773), .C2(new_n758), .ZN(new_n1033));
  AOI21_X1  g0833(.A(new_n1033), .B1(G303), .B2(new_n740), .ZN(new_n1034));
  OAI221_X1 g0834(.A(new_n283), .B1(new_n802), .B2(new_n212), .C1(new_n301), .C2(new_n743), .ZN(new_n1035));
  INV_X1    g0835(.A(new_n1035), .ZN(new_n1036));
  NAND2_X1  g0836(.A1(new_n753), .A2(G77), .ZN(new_n1037));
  OAI211_X1 g0837(.A(new_n1036), .B(new_n1037), .C1(new_n216), .C2(new_n747), .ZN(new_n1038));
  OAI22_X1  g0838(.A1(new_n759), .A2(new_n736), .B1(new_n766), .B2(new_n936), .ZN(new_n1039));
  XNOR2_X1  g0839(.A(new_n1039), .B(KEYINPUT51), .ZN(new_n1040));
  OAI21_X1  g0840(.A(new_n1040), .B1(new_n207), .B2(new_n750), .ZN(new_n1041));
  AOI211_X1 g0841(.A(new_n1038), .B(new_n1041), .C1(G143), .C2(new_n927), .ZN(new_n1042));
  XNOR2_X1  g0842(.A(new_n1042), .B(KEYINPUT120), .ZN(new_n1043));
  OAI21_X1  g0843(.A(new_n725), .B1(new_n1034), .B2(new_n1043), .ZN(new_n1044));
  OAI221_X1 g0844(.A(new_n726), .B1(new_n209), .B2(new_n236), .C1(new_n255), .C2(new_n957), .ZN(new_n1045));
  AOI21_X1  g0845(.A(new_n730), .B1(new_n987), .B2(new_n724), .ZN(new_n1046));
  NAND3_X1  g0846(.A1(new_n1044), .A2(new_n1045), .A3(new_n1046), .ZN(new_n1047));
  INV_X1    g0847(.A(new_n960), .ZN(new_n1048));
  OAI211_X1 g0848(.A(new_n1026), .B(new_n1047), .C1(new_n1048), .C2(new_n969), .ZN(G390));
  OR2_X1    g0849(.A1(new_n877), .A2(new_n723), .ZN(new_n1050));
  NAND2_X1  g0850(.A1(new_n817), .A2(new_n264), .ZN(new_n1051));
  OAI21_X1  g0851(.A(new_n283), .B1(new_n750), .B2(new_n212), .ZN(new_n1052));
  XNOR2_X1  g0852(.A(new_n1052), .B(KEYINPUT123), .ZN(new_n1053));
  AOI22_X1  g0853(.A1(new_n740), .A2(G137), .B1(new_n756), .B2(G128), .ZN(new_n1054));
  AND2_X1   g0854(.A1(new_n1053), .A2(new_n1054), .ZN(new_n1055));
  XOR2_X1   g0855(.A(KEYINPUT54), .B(G143), .Z(new_n1056));
  NAND2_X1  g0856(.A1(new_n807), .A2(new_n1056), .ZN(new_n1057));
  INV_X1    g0857(.A(G132), .ZN(new_n1058));
  OAI22_X1  g0858(.A1(new_n736), .A2(new_n1058), .B1(new_n754), .B2(new_n759), .ZN(new_n1059));
  AOI21_X1  g0859(.A(new_n1059), .B1(G125), .B2(new_n797), .ZN(new_n1060));
  NOR2_X1   g0860(.A1(new_n747), .A2(new_n936), .ZN(new_n1061));
  XNOR2_X1  g0861(.A(new_n1061), .B(KEYINPUT53), .ZN(new_n1062));
  NAND4_X1  g0862(.A1(new_n1055), .A2(new_n1057), .A3(new_n1060), .A4(new_n1062), .ZN(new_n1063));
  OAI22_X1  g0863(.A1(new_n763), .A2(new_n930), .B1(new_n769), .B2(new_n766), .ZN(new_n1064));
  AOI211_X1 g0864(.A(new_n799), .B(new_n1064), .C1(G97), .C2(new_n807), .ZN(new_n1065));
  AND2_X1   g0865(.A1(new_n1065), .A2(new_n1037), .ZN(new_n1066));
  OAI221_X1 g0866(.A(new_n1066), .B1(new_n207), .B2(new_n747), .C1(new_n218), .C2(new_n736), .ZN(new_n1067));
  OAI21_X1  g0867(.A(new_n448), .B1(new_n802), .B2(new_n555), .ZN(new_n1068));
  OAI21_X1  g0868(.A(new_n1063), .B1(new_n1067), .B2(new_n1068), .ZN(new_n1069));
  NAND2_X1  g0869(.A1(new_n1069), .A2(new_n725), .ZN(new_n1070));
  NAND4_X1  g0870(.A1(new_n1050), .A2(new_n731), .A3(new_n1051), .A4(new_n1070), .ZN(new_n1071));
  NAND2_X1  g0871(.A1(new_n887), .A2(new_n878), .ZN(new_n1072));
  NAND4_X1  g0872(.A1(new_n1072), .A2(new_n871), .A3(new_n874), .A4(new_n876), .ZN(new_n1073));
  INV_X1    g0873(.A(new_n821), .ZN(new_n1074));
  OAI21_X1  g0874(.A(new_n881), .B1(new_n685), .B2(new_n1074), .ZN(new_n1075));
  NAND2_X1  g0875(.A1(new_n1075), .A2(new_n886), .ZN(new_n1076));
  NAND3_X1  g0876(.A1(new_n1076), .A2(new_n905), .A3(new_n878), .ZN(new_n1077));
  NAND2_X1  g0877(.A1(new_n1073), .A2(new_n1077), .ZN(new_n1078));
  AND3_X1   g0878(.A1(new_n908), .A2(new_n909), .A3(G330), .ZN(new_n1079));
  INV_X1    g0879(.A(new_n1079), .ZN(new_n1080));
  NAND2_X1  g0880(.A1(new_n1078), .A2(new_n1080), .ZN(new_n1081));
  NAND2_X1  g0881(.A1(new_n825), .A2(G330), .ZN(new_n1082));
  INV_X1    g0882(.A(new_n1082), .ZN(new_n1083));
  NAND3_X1  g0883(.A1(new_n713), .A2(new_n886), .A3(new_n1083), .ZN(new_n1084));
  INV_X1    g0884(.A(new_n1084), .ZN(new_n1085));
  NAND3_X1  g0885(.A1(new_n1085), .A2(new_n1073), .A3(new_n1077), .ZN(new_n1086));
  NAND2_X1  g0886(.A1(new_n1081), .A2(new_n1086), .ZN(new_n1087));
  INV_X1    g0887(.A(new_n1087), .ZN(new_n1088));
  OAI21_X1  g0888(.A(new_n1071), .B1(new_n1088), .B2(new_n1048), .ZN(new_n1089));
  NAND3_X1  g0889(.A1(new_n908), .A2(new_n430), .A3(G330), .ZN(new_n1090));
  NAND4_X1  g0890(.A1(new_n1090), .A2(new_n896), .A3(new_n300), .A4(new_n634), .ZN(new_n1091));
  AOI21_X1  g0891(.A(new_n886), .B1(new_n713), .B2(new_n1083), .ZN(new_n1092));
  OAI21_X1  g0892(.A(new_n882), .B1(new_n1079), .B2(new_n1092), .ZN(new_n1093));
  INV_X1    g0893(.A(new_n1075), .ZN(new_n1094));
  AOI21_X1  g0894(.A(new_n1082), .B1(new_n902), .B2(new_n903), .ZN(new_n1095));
  OAI211_X1 g0895(.A(new_n1094), .B(new_n1084), .C1(new_n1095), .C2(new_n886), .ZN(new_n1096));
  AOI21_X1  g0896(.A(new_n1091), .B1(new_n1093), .B2(new_n1096), .ZN(new_n1097));
  INV_X1    g0897(.A(KEYINPUT122), .ZN(new_n1098));
  AND3_X1   g0898(.A1(new_n1097), .A2(new_n1087), .A3(new_n1098), .ZN(new_n1099));
  AOI21_X1  g0899(.A(new_n1098), .B1(new_n1097), .B2(new_n1087), .ZN(new_n1100));
  NOR2_X1   g0900(.A1(new_n1099), .A2(new_n1100), .ZN(new_n1101));
  INV_X1    g0901(.A(new_n1097), .ZN(new_n1102));
  AOI21_X1  g0902(.A(new_n1101), .B1(new_n1088), .B2(new_n1102), .ZN(new_n1103));
  AOI21_X1  g0903(.A(new_n1089), .B1(new_n1103), .B2(new_n673), .ZN(new_n1104));
  INV_X1    g0904(.A(new_n1104), .ZN(G378));
  INV_X1    g0905(.A(new_n1091), .ZN(new_n1106));
  OAI21_X1  g0906(.A(new_n1106), .B1(new_n1099), .B2(new_n1100), .ZN(new_n1107));
  INV_X1    g0907(.A(KEYINPUT125), .ZN(new_n1108));
  NAND2_X1  g0908(.A1(new_n1107), .A2(new_n1108), .ZN(new_n1109));
  OAI21_X1  g0909(.A(new_n300), .B1(new_n333), .B2(new_n334), .ZN(new_n1110));
  XNOR2_X1  g0910(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1111));
  XNOR2_X1  g0911(.A(new_n1110), .B(new_n1111), .ZN(new_n1112));
  NAND2_X1  g0912(.A1(new_n278), .A2(new_n654), .ZN(new_n1113));
  XNOR2_X1  g0913(.A(new_n1112), .B(new_n1113), .ZN(new_n1114));
  INV_X1    g0914(.A(new_n1114), .ZN(new_n1115));
  OAI21_X1  g0915(.A(G330), .B1(new_n906), .B2(new_n910), .ZN(new_n1116));
  AND3_X1   g0916(.A1(new_n892), .A2(new_n1116), .A3(new_n894), .ZN(new_n1117));
  AOI21_X1  g0917(.A(new_n1116), .B1(new_n892), .B2(new_n894), .ZN(new_n1118));
  OAI21_X1  g0918(.A(new_n1115), .B1(new_n1117), .B2(new_n1118), .ZN(new_n1119));
  INV_X1    g0919(.A(new_n1116), .ZN(new_n1120));
  NAND2_X1  g0920(.A1(new_n895), .A2(new_n1120), .ZN(new_n1121));
  NAND3_X1  g0921(.A1(new_n892), .A2(new_n1116), .A3(new_n894), .ZN(new_n1122));
  NAND3_X1  g0922(.A1(new_n1121), .A2(new_n1114), .A3(new_n1122), .ZN(new_n1123));
  NAND2_X1  g0923(.A1(new_n1119), .A2(new_n1123), .ZN(new_n1124));
  OAI211_X1 g0924(.A(KEYINPUT125), .B(new_n1106), .C1(new_n1099), .C2(new_n1100), .ZN(new_n1125));
  NAND3_X1  g0925(.A1(new_n1109), .A2(new_n1124), .A3(new_n1125), .ZN(new_n1126));
  INV_X1    g0926(.A(KEYINPUT57), .ZN(new_n1127));
  NAND2_X1  g0927(.A1(new_n1126), .A2(new_n1127), .ZN(new_n1128));
  NAND4_X1  g0928(.A1(new_n1109), .A2(new_n1124), .A3(KEYINPUT57), .A4(new_n1125), .ZN(new_n1129));
  NAND3_X1  g0929(.A1(new_n1128), .A2(new_n673), .A3(new_n1129), .ZN(new_n1130));
  AOI21_X1  g0930(.A(new_n1048), .B1(new_n1119), .B2(new_n1123), .ZN(new_n1131));
  NAND2_X1  g0931(.A1(new_n816), .A2(new_n212), .ZN(new_n1132));
  OAI21_X1  g0932(.A(new_n1132), .B1(new_n1114), .B2(new_n723), .ZN(new_n1133));
  AOI22_X1  g0933(.A1(new_n797), .A2(G283), .B1(new_n737), .B2(G107), .ZN(new_n1134));
  OAI221_X1 g0934(.A(new_n1134), .B1(new_n218), .B2(new_n766), .C1(new_n388), .C2(new_n750), .ZN(new_n1135));
  AOI211_X1 g0935(.A(new_n934), .B(new_n1135), .C1(new_n304), .C2(new_n807), .ZN(new_n1136));
  AOI211_X1 g0936(.A(G41), .B(new_n283), .C1(new_n740), .C2(G97), .ZN(new_n1137));
  OAI211_X1 g0937(.A(new_n1136), .B(new_n1137), .C1(new_n309), .C2(new_n747), .ZN(new_n1138));
  XNOR2_X1  g0938(.A(new_n1138), .B(KEYINPUT58), .ZN(new_n1139));
  INV_X1    g0939(.A(G124), .ZN(new_n1140));
  OAI21_X1  g0940(.A(new_n280), .B1(new_n758), .B2(new_n1140), .ZN(new_n1141));
  AOI22_X1  g0941(.A1(new_n737), .A2(G128), .B1(G125), .B2(new_n756), .ZN(new_n1142));
  AOI22_X1  g0942(.A1(new_n807), .A2(G137), .B1(G150), .B2(new_n753), .ZN(new_n1143));
  NAND2_X1  g0943(.A1(new_n740), .A2(G132), .ZN(new_n1144));
  NAND2_X1  g0944(.A1(new_n748), .A2(new_n1056), .ZN(new_n1145));
  NAND4_X1  g0945(.A1(new_n1142), .A2(new_n1143), .A3(new_n1144), .A4(new_n1145), .ZN(new_n1146));
  AOI211_X1 g0946(.A(G41), .B(new_n1141), .C1(new_n1146), .C2(KEYINPUT59), .ZN(new_n1147));
  OAI221_X1 g0947(.A(new_n1147), .B1(KEYINPUT59), .B2(new_n1146), .C1(new_n759), .C2(new_n750), .ZN(new_n1148));
  OAI21_X1  g0948(.A(new_n212), .B1(new_n375), .B2(G41), .ZN(new_n1149));
  NAND2_X1  g0949(.A1(new_n1148), .A2(new_n1149), .ZN(new_n1150));
  INV_X1    g0950(.A(new_n1150), .ZN(new_n1151));
  AOI21_X1  g0951(.A(new_n814), .B1(new_n1139), .B2(new_n1151), .ZN(new_n1152));
  NOR3_X1   g0952(.A1(new_n1133), .A2(new_n730), .A3(new_n1152), .ZN(new_n1153));
  NOR2_X1   g0953(.A1(new_n1131), .A2(new_n1153), .ZN(new_n1154));
  NAND2_X1  g0954(.A1(new_n1154), .A2(KEYINPUT124), .ZN(new_n1155));
  INV_X1    g0955(.A(KEYINPUT124), .ZN(new_n1156));
  OAI21_X1  g0956(.A(new_n1156), .B1(new_n1131), .B2(new_n1153), .ZN(new_n1157));
  NAND2_X1  g0957(.A1(new_n1155), .A2(new_n1157), .ZN(new_n1158));
  NAND2_X1  g0958(.A1(new_n1130), .A2(new_n1158), .ZN(G375));
  AOI22_X1  g0959(.A1(new_n807), .A2(G107), .B1(G116), .B2(new_n740), .ZN(new_n1160));
  INV_X1    g0960(.A(KEYINPUT126), .ZN(new_n1161));
  NAND2_X1  g0961(.A1(new_n1160), .A2(new_n1161), .ZN(new_n1162));
  AOI21_X1  g0962(.A(new_n283), .B1(new_n737), .B2(G283), .ZN(new_n1163));
  OAI211_X1 g0963(.A(new_n1162), .B(new_n1163), .C1(new_n449), .C2(new_n763), .ZN(new_n1164));
  OAI221_X1 g0964(.A(new_n1005), .B1(new_n930), .B2(new_n766), .C1(new_n1160), .C2(new_n1161), .ZN(new_n1165));
  NOR2_X1   g0965(.A1(new_n747), .A2(new_n209), .ZN(new_n1166));
  NOR4_X1   g0966(.A1(new_n1164), .A2(new_n1165), .A3(new_n941), .A4(new_n1166), .ZN(new_n1167));
  NOR2_X1   g0967(.A1(new_n743), .A2(new_n936), .ZN(new_n1168));
  OAI22_X1  g0968(.A1(new_n754), .A2(new_n212), .B1(new_n750), .B2(new_n388), .ZN(new_n1169));
  AOI21_X1  g0969(.A(new_n1169), .B1(G159), .B2(new_n748), .ZN(new_n1170));
  NAND2_X1  g0970(.A1(new_n797), .A2(G128), .ZN(new_n1171));
  NAND2_X1  g0971(.A1(new_n740), .A2(new_n1056), .ZN(new_n1172));
  AOI21_X1  g0972(.A(new_n448), .B1(new_n737), .B2(G137), .ZN(new_n1173));
  NAND4_X1  g0973(.A1(new_n1170), .A2(new_n1171), .A3(new_n1172), .A4(new_n1173), .ZN(new_n1174));
  AOI211_X1 g0974(.A(new_n1168), .B(new_n1174), .C1(G132), .C2(new_n756), .ZN(new_n1175));
  OAI21_X1  g0975(.A(new_n725), .B1(new_n1167), .B2(new_n1175), .ZN(new_n1176));
  OAI211_X1 g0976(.A(new_n731), .B(new_n1176), .C1(new_n886), .C2(new_n723), .ZN(new_n1177));
  AOI21_X1  g0977(.A(new_n1177), .B1(new_n216), .B2(new_n817), .ZN(new_n1178));
  NAND2_X1  g0978(.A1(new_n1093), .A2(new_n1096), .ZN(new_n1179));
  AOI21_X1  g0979(.A(new_n1178), .B1(new_n1179), .B2(new_n960), .ZN(new_n1180));
  NAND3_X1  g0980(.A1(new_n1093), .A2(new_n1091), .A3(new_n1096), .ZN(new_n1181));
  NAND2_X1  g0981(.A1(new_n1181), .A2(new_n978), .ZN(new_n1182));
  OAI21_X1  g0982(.A(new_n1180), .B1(new_n1182), .B2(new_n1097), .ZN(G381));
  NAND3_X1  g0983(.A1(new_n1130), .A2(new_n1158), .A3(new_n1104), .ZN(new_n1184));
  NOR3_X1   g0984(.A1(new_n1184), .A2(G384), .A3(G381), .ZN(new_n1185));
  NOR2_X1   g0985(.A1(G387), .A2(G390), .ZN(new_n1186));
  NOR2_X1   g0986(.A1(G393), .A2(G396), .ZN(new_n1187));
  NAND3_X1  g0987(.A1(new_n1185), .A2(new_n1186), .A3(new_n1187), .ZN(G407));
  OAI211_X1 g0988(.A(G407), .B(G213), .C1(G343), .C2(new_n1184), .ZN(G409));
  NAND2_X1  g0989(.A1(G375), .A2(G378), .ZN(new_n1190));
  INV_X1    g0990(.A(KEYINPUT60), .ZN(new_n1191));
  OR2_X1    g0991(.A1(new_n1181), .A2(new_n1191), .ZN(new_n1192));
  NAND2_X1  g0992(.A1(new_n1181), .A2(new_n1191), .ZN(new_n1193));
  NAND4_X1  g0993(.A1(new_n1192), .A2(new_n673), .A3(new_n1102), .A4(new_n1193), .ZN(new_n1194));
  NAND2_X1  g0994(.A1(new_n1194), .A2(new_n1180), .ZN(new_n1195));
  OR2_X1    g0995(.A1(new_n1195), .A2(new_n832), .ZN(new_n1196));
  NAND2_X1  g0996(.A1(new_n832), .A2(new_n1195), .ZN(new_n1197));
  NAND2_X1  g0997(.A1(new_n1196), .A2(new_n1197), .ZN(new_n1198));
  INV_X1    g0998(.A(new_n1198), .ZN(new_n1199));
  INV_X1    g0999(.A(G213), .ZN(new_n1200));
  NOR2_X1   g1000(.A1(new_n1200), .A2(G343), .ZN(new_n1201));
  INV_X1    g1001(.A(new_n1201), .ZN(new_n1202));
  NAND4_X1  g1002(.A1(new_n1109), .A2(new_n1124), .A3(new_n978), .A4(new_n1125), .ZN(new_n1203));
  NAND3_X1  g1003(.A1(new_n1104), .A2(new_n1154), .A3(new_n1203), .ZN(new_n1204));
  NAND4_X1  g1004(.A1(new_n1190), .A2(new_n1199), .A3(new_n1202), .A4(new_n1204), .ZN(new_n1205));
  NAND2_X1  g1005(.A1(new_n1205), .A2(KEYINPUT62), .ZN(new_n1206));
  NAND3_X1  g1006(.A1(new_n1190), .A2(new_n1202), .A3(new_n1204), .ZN(new_n1207));
  NAND2_X1  g1007(.A1(new_n1201), .A2(G2897), .ZN(new_n1208));
  XNOR2_X1  g1008(.A(new_n1198), .B(new_n1208), .ZN(new_n1209));
  NAND2_X1  g1009(.A1(new_n1207), .A2(new_n1209), .ZN(new_n1210));
  INV_X1    g1010(.A(KEYINPUT61), .ZN(new_n1211));
  AOI21_X1  g1011(.A(new_n1201), .B1(G375), .B2(G378), .ZN(new_n1212));
  INV_X1    g1012(.A(KEYINPUT62), .ZN(new_n1213));
  NAND4_X1  g1013(.A1(new_n1212), .A2(new_n1213), .A3(new_n1199), .A4(new_n1204), .ZN(new_n1214));
  NAND4_X1  g1014(.A1(new_n1206), .A2(new_n1210), .A3(new_n1211), .A4(new_n1214), .ZN(new_n1215));
  XNOR2_X1  g1015(.A(G387), .B(G390), .ZN(new_n1216));
  XNOR2_X1  g1016(.A(G393), .B(new_n788), .ZN(new_n1217));
  XNOR2_X1  g1017(.A(new_n1216), .B(new_n1217), .ZN(new_n1218));
  NAND2_X1  g1018(.A1(new_n1215), .A2(new_n1218), .ZN(new_n1219));
  NAND2_X1  g1019(.A1(new_n1207), .A2(KEYINPUT127), .ZN(new_n1220));
  INV_X1    g1020(.A(KEYINPUT127), .ZN(new_n1221));
  NAND3_X1  g1021(.A1(new_n1212), .A2(new_n1221), .A3(new_n1204), .ZN(new_n1222));
  NAND3_X1  g1022(.A1(new_n1220), .A2(new_n1209), .A3(new_n1222), .ZN(new_n1223));
  INV_X1    g1023(.A(KEYINPUT63), .ZN(new_n1224));
  AOI21_X1  g1024(.A(new_n1218), .B1(new_n1205), .B2(new_n1224), .ZN(new_n1225));
  AOI21_X1  g1025(.A(new_n1104), .B1(new_n1130), .B2(new_n1158), .ZN(new_n1226));
  INV_X1    g1026(.A(new_n1204), .ZN(new_n1227));
  NOR4_X1   g1027(.A1(new_n1226), .A2(new_n1198), .A3(new_n1201), .A4(new_n1227), .ZN(new_n1228));
  AOI21_X1  g1028(.A(KEYINPUT61), .B1(new_n1228), .B2(KEYINPUT63), .ZN(new_n1229));
  NAND3_X1  g1029(.A1(new_n1223), .A2(new_n1225), .A3(new_n1229), .ZN(new_n1230));
  NAND2_X1  g1030(.A1(new_n1219), .A2(new_n1230), .ZN(G405));
  NAND2_X1  g1031(.A1(new_n1190), .A2(new_n1184), .ZN(new_n1232));
  NAND2_X1  g1032(.A1(new_n1232), .A2(new_n1199), .ZN(new_n1233));
  NAND3_X1  g1033(.A1(new_n1190), .A2(new_n1184), .A3(new_n1198), .ZN(new_n1234));
  NAND2_X1  g1034(.A1(new_n1233), .A2(new_n1234), .ZN(new_n1235));
  INV_X1    g1035(.A(new_n1218), .ZN(new_n1236));
  XNOR2_X1  g1036(.A(new_n1235), .B(new_n1236), .ZN(G402));
endmodule


