//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 1 1 0 1 0 1 0 0 1 1 0 1 1 0 1 0 0 1 1 0 0 0 0 1 1 1 0 0 1 1 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 0 1 1 1 1 0 0 0 1 1 1 0 0 1 0 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:34:43 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n445, new_n447, new_n451, new_n452, new_n453, new_n454, new_n455,
    new_n458, new_n459, new_n460, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n483, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n532, new_n533, new_n534, new_n535, new_n536, new_n537, new_n538,
    new_n541, new_n542, new_n543, new_n544, new_n545, new_n546, new_n547,
    new_n548, new_n549, new_n550, new_n551, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n570, new_n572, new_n573,
    new_n575, new_n576, new_n577, new_n578, new_n579, new_n580, new_n581,
    new_n582, new_n583, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n592, new_n593, new_n594, new_n595, new_n596, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n619, new_n622, new_n624, new_n625, new_n626,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1151, new_n1152, new_n1153, new_n1154,
    new_n1156;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  NAND2_X1  g019(.A1(G94), .A2(G452), .ZN(new_n445));
  XNOR2_X1  g020(.A(new_n445), .B(KEYINPUT64), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g025(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n451));
  XOR2_X1   g026(.A(KEYINPUT65), .B(KEYINPUT2), .Z(new_n452));
  XNOR2_X1  g027(.A(new_n451), .B(new_n452), .ZN(new_n453));
  NOR4_X1   g028(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(new_n455));
  NOR2_X1   g030(.A1(new_n453), .A2(new_n455), .ZN(G325));
  INV_X1    g031(.A(G325), .ZN(G261));
  NAND2_X1  g032(.A1(new_n453), .A2(G2106), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n455), .A2(G567), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  INV_X1    g035(.A(new_n460), .ZN(G319));
  INV_X1    g036(.A(KEYINPUT67), .ZN(new_n462));
  INV_X1    g037(.A(G2104), .ZN(new_n463));
  AOI21_X1  g038(.A(new_n462), .B1(KEYINPUT3), .B2(new_n463), .ZN(new_n464));
  XNOR2_X1  g039(.A(KEYINPUT66), .B(KEYINPUT3), .ZN(new_n465));
  OAI21_X1  g040(.A(new_n464), .B1(new_n465), .B2(new_n463), .ZN(new_n466));
  INV_X1    g041(.A(KEYINPUT66), .ZN(new_n467));
  NOR2_X1   g042(.A1(new_n467), .A2(KEYINPUT3), .ZN(new_n468));
  INV_X1    g043(.A(KEYINPUT3), .ZN(new_n469));
  NOR2_X1   g044(.A1(new_n469), .A2(KEYINPUT66), .ZN(new_n470));
  OAI211_X1 g045(.A(new_n462), .B(G2104), .C1(new_n468), .C2(new_n470), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n466), .A2(new_n471), .ZN(new_n472));
  INV_X1    g047(.A(G2105), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n472), .A2(new_n473), .ZN(new_n474));
  INV_X1    g049(.A(new_n474), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n475), .A2(G137), .ZN(new_n476));
  XNOR2_X1  g051(.A(KEYINPUT3), .B(G2104), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n477), .A2(G125), .ZN(new_n478));
  INV_X1    g053(.A(G113), .ZN(new_n479));
  OAI21_X1  g054(.A(new_n478), .B1(new_n479), .B2(new_n463), .ZN(new_n480));
  NOR2_X1   g055(.A1(new_n463), .A2(G2105), .ZN(new_n481));
  AOI22_X1  g056(.A1(new_n480), .A2(G2105), .B1(G101), .B2(new_n481), .ZN(new_n482));
  NAND2_X1  g057(.A1(new_n476), .A2(new_n482), .ZN(new_n483));
  INV_X1    g058(.A(new_n483), .ZN(G160));
  NAND2_X1  g059(.A1(new_n475), .A2(G136), .ZN(new_n485));
  NAND2_X1  g060(.A1(new_n472), .A2(G2105), .ZN(new_n486));
  INV_X1    g061(.A(new_n486), .ZN(new_n487));
  NAND2_X1  g062(.A1(new_n487), .A2(G124), .ZN(new_n488));
  OR2_X1    g063(.A1(G100), .A2(G2105), .ZN(new_n489));
  OAI211_X1 g064(.A(new_n489), .B(G2104), .C1(G112), .C2(new_n473), .ZN(new_n490));
  NAND3_X1  g065(.A1(new_n485), .A2(new_n488), .A3(new_n490), .ZN(new_n491));
  INV_X1    g066(.A(new_n491), .ZN(G162));
  NAND3_X1  g067(.A1(new_n477), .A2(G138), .A3(new_n473), .ZN(new_n493));
  INV_X1    g068(.A(KEYINPUT4), .ZN(new_n494));
  NAND2_X1  g069(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  NAND2_X1  g070(.A1(KEYINPUT4), .A2(G138), .ZN(new_n496));
  OAI21_X1  g071(.A(new_n495), .B1(new_n474), .B2(new_n496), .ZN(new_n497));
  OAI21_X1  g072(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n498));
  INV_X1    g073(.A(G114), .ZN(new_n499));
  AOI21_X1  g074(.A(new_n498), .B1(new_n499), .B2(G2105), .ZN(new_n500));
  INV_X1    g075(.A(new_n500), .ZN(new_n501));
  NAND2_X1  g076(.A1(G126), .A2(G2105), .ZN(new_n502));
  INV_X1    g077(.A(new_n502), .ZN(new_n503));
  AOI21_X1  g078(.A(KEYINPUT68), .B1(new_n472), .B2(new_n503), .ZN(new_n504));
  INV_X1    g079(.A(KEYINPUT68), .ZN(new_n505));
  AOI211_X1 g080(.A(new_n505), .B(new_n502), .C1(new_n466), .C2(new_n471), .ZN(new_n506));
  OAI21_X1  g081(.A(new_n501), .B1(new_n504), .B2(new_n506), .ZN(new_n507));
  INV_X1    g082(.A(KEYINPUT69), .ZN(new_n508));
  NAND2_X1  g083(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  OAI211_X1 g084(.A(KEYINPUT69), .B(new_n501), .C1(new_n504), .C2(new_n506), .ZN(new_n510));
  AOI21_X1  g085(.A(new_n497), .B1(new_n509), .B2(new_n510), .ZN(G164));
  INV_X1    g086(.A(G651), .ZN(new_n512));
  OR2_X1    g087(.A1(KEYINPUT70), .A2(KEYINPUT6), .ZN(new_n513));
  NAND2_X1  g088(.A1(KEYINPUT70), .A2(KEYINPUT6), .ZN(new_n514));
  AOI21_X1  g089(.A(new_n512), .B1(new_n513), .B2(new_n514), .ZN(new_n515));
  INV_X1    g090(.A(KEYINPUT71), .ZN(new_n516));
  NAND2_X1  g091(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  INV_X1    g092(.A(KEYINPUT6), .ZN(new_n518));
  OAI21_X1  g093(.A(KEYINPUT71), .B1(new_n518), .B2(G651), .ZN(new_n519));
  OAI21_X1  g094(.A(new_n517), .B1(new_n515), .B2(new_n519), .ZN(new_n520));
  AND2_X1   g095(.A1(new_n520), .A2(G543), .ZN(new_n521));
  NAND2_X1  g096(.A1(G75), .A2(G543), .ZN(new_n522));
  INV_X1    g097(.A(KEYINPUT72), .ZN(new_n523));
  INV_X1    g098(.A(G543), .ZN(new_n524));
  OAI21_X1  g099(.A(new_n523), .B1(new_n524), .B2(KEYINPUT5), .ZN(new_n525));
  INV_X1    g100(.A(KEYINPUT5), .ZN(new_n526));
  NAND3_X1  g101(.A1(new_n526), .A2(KEYINPUT72), .A3(G543), .ZN(new_n527));
  AOI22_X1  g102(.A1(new_n525), .A2(new_n527), .B1(KEYINPUT5), .B2(new_n524), .ZN(new_n528));
  INV_X1    g103(.A(new_n528), .ZN(new_n529));
  INV_X1    g104(.A(G62), .ZN(new_n530));
  OAI21_X1  g105(.A(new_n522), .B1(new_n529), .B2(new_n530), .ZN(new_n531));
  AOI22_X1  g106(.A1(new_n521), .A2(G50), .B1(G651), .B2(new_n531), .ZN(new_n532));
  NAND2_X1  g107(.A1(new_n520), .A2(new_n528), .ZN(new_n533));
  INV_X1    g108(.A(KEYINPUT73), .ZN(new_n534));
  NAND2_X1  g109(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  NAND3_X1  g110(.A1(new_n520), .A2(KEYINPUT73), .A3(new_n528), .ZN(new_n536));
  NAND2_X1  g111(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  INV_X1    g112(.A(G88), .ZN(new_n538));
  OAI21_X1  g113(.A(new_n532), .B1(new_n537), .B2(new_n538), .ZN(G303));
  INV_X1    g114(.A(G303), .ZN(G166));
  NAND2_X1  g115(.A1(new_n521), .A2(G51), .ZN(new_n541));
  INV_X1    g116(.A(KEYINPUT74), .ZN(new_n542));
  XNOR2_X1  g117(.A(new_n528), .B(new_n542), .ZN(new_n543));
  NAND2_X1  g118(.A1(G63), .A2(G651), .ZN(new_n544));
  OR2_X1    g119(.A1(new_n543), .A2(new_n544), .ZN(new_n545));
  NAND3_X1  g120(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n546));
  XNOR2_X1  g121(.A(new_n546), .B(KEYINPUT7), .ZN(new_n547));
  AND3_X1   g122(.A1(new_n541), .A2(new_n545), .A3(new_n547), .ZN(new_n548));
  INV_X1    g123(.A(G89), .ZN(new_n549));
  OAI21_X1  g124(.A(new_n548), .B1(new_n549), .B2(new_n537), .ZN(new_n550));
  INV_X1    g125(.A(KEYINPUT75), .ZN(new_n551));
  XNOR2_X1  g126(.A(new_n550), .B(new_n551), .ZN(G168));
  AND2_X1   g127(.A1(new_n535), .A2(new_n536), .ZN(new_n553));
  XOR2_X1   g128(.A(KEYINPUT76), .B(G90), .Z(new_n554));
  NAND2_X1  g129(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  NAND2_X1  g130(.A1(G77), .A2(G543), .ZN(new_n556));
  INV_X1    g131(.A(G64), .ZN(new_n557));
  OAI21_X1  g132(.A(new_n556), .B1(new_n543), .B2(new_n557), .ZN(new_n558));
  AOI22_X1  g133(.A1(new_n558), .A2(G651), .B1(G52), .B2(new_n521), .ZN(new_n559));
  NAND2_X1  g134(.A1(new_n555), .A2(new_n559), .ZN(G301));
  INV_X1    g135(.A(G301), .ZN(G171));
  NAND2_X1  g136(.A1(new_n553), .A2(G81), .ZN(new_n562));
  NAND2_X1  g137(.A1(G68), .A2(G543), .ZN(new_n563));
  INV_X1    g138(.A(G56), .ZN(new_n564));
  OAI21_X1  g139(.A(new_n563), .B1(new_n543), .B2(new_n564), .ZN(new_n565));
  AOI22_X1  g140(.A1(new_n565), .A2(G651), .B1(G43), .B2(new_n521), .ZN(new_n566));
  AND2_X1   g141(.A1(new_n562), .A2(new_n566), .ZN(new_n567));
  NAND2_X1  g142(.A1(new_n567), .A2(G860), .ZN(new_n568));
  XNOR2_X1  g143(.A(new_n568), .B(KEYINPUT77), .ZN(G153));
  AND3_X1   g144(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n570));
  NAND2_X1  g145(.A1(new_n570), .A2(G36), .ZN(G176));
  NAND2_X1  g146(.A1(G1), .A2(G3), .ZN(new_n572));
  XNOR2_X1  g147(.A(new_n572), .B(KEYINPUT8), .ZN(new_n573));
  NAND2_X1  g148(.A1(new_n570), .A2(new_n573), .ZN(G188));
  NAND2_X1  g149(.A1(new_n520), .A2(G543), .ZN(new_n575));
  INV_X1    g150(.A(G53), .ZN(new_n576));
  OAI21_X1  g151(.A(KEYINPUT9), .B1(new_n575), .B2(new_n576), .ZN(new_n577));
  INV_X1    g152(.A(KEYINPUT9), .ZN(new_n578));
  NAND4_X1  g153(.A1(new_n520), .A2(new_n578), .A3(G53), .A4(G543), .ZN(new_n579));
  NAND2_X1  g154(.A1(new_n577), .A2(new_n579), .ZN(new_n580));
  NAND3_X1  g155(.A1(new_n535), .A2(G91), .A3(new_n536), .ZN(new_n581));
  AOI22_X1  g156(.A1(new_n528), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n582));
  OR2_X1    g157(.A1(new_n582), .A2(new_n512), .ZN(new_n583));
  NAND3_X1  g158(.A1(new_n580), .A2(new_n581), .A3(new_n583), .ZN(G299));
  XNOR2_X1  g159(.A(new_n550), .B(KEYINPUT75), .ZN(G286));
  AOI22_X1  g160(.A1(new_n553), .A2(G87), .B1(G49), .B2(new_n521), .ZN(new_n586));
  INV_X1    g161(.A(G74), .ZN(new_n587));
  AOI21_X1  g162(.A(new_n512), .B1(new_n543), .B2(new_n587), .ZN(new_n588));
  INV_X1    g163(.A(KEYINPUT78), .ZN(new_n589));
  XNOR2_X1  g164(.A(new_n588), .B(new_n589), .ZN(new_n590));
  NAND2_X1  g165(.A1(new_n586), .A2(new_n590), .ZN(G288));
  NAND2_X1  g166(.A1(G73), .A2(G543), .ZN(new_n592));
  INV_X1    g167(.A(G61), .ZN(new_n593));
  OAI21_X1  g168(.A(new_n592), .B1(new_n529), .B2(new_n593), .ZN(new_n594));
  AOI22_X1  g169(.A1(new_n521), .A2(G48), .B1(G651), .B2(new_n594), .ZN(new_n595));
  INV_X1    g170(.A(G86), .ZN(new_n596));
  OAI21_X1  g171(.A(new_n595), .B1(new_n537), .B2(new_n596), .ZN(G305));
  NAND2_X1  g172(.A1(G72), .A2(G543), .ZN(new_n598));
  INV_X1    g173(.A(G60), .ZN(new_n599));
  OAI21_X1  g174(.A(new_n598), .B1(new_n543), .B2(new_n599), .ZN(new_n600));
  AOI22_X1  g175(.A1(new_n600), .A2(G651), .B1(G47), .B2(new_n521), .ZN(new_n601));
  INV_X1    g176(.A(G85), .ZN(new_n602));
  OAI21_X1  g177(.A(new_n601), .B1(new_n602), .B2(new_n537), .ZN(G290));
  NAND2_X1  g178(.A1(G301), .A2(G868), .ZN(new_n604));
  AOI22_X1  g179(.A1(new_n528), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n605));
  AOI21_X1  g180(.A(new_n512), .B1(new_n605), .B2(KEYINPUT80), .ZN(new_n606));
  OAI21_X1  g181(.A(new_n606), .B1(KEYINPUT80), .B2(new_n605), .ZN(new_n607));
  OAI21_X1  g182(.A(G54), .B1(new_n521), .B2(KEYINPUT79), .ZN(new_n608));
  AND3_X1   g183(.A1(new_n520), .A2(KEYINPUT79), .A3(G543), .ZN(new_n609));
  OAI21_X1  g184(.A(new_n607), .B1(new_n608), .B2(new_n609), .ZN(new_n610));
  AND2_X1   g185(.A1(new_n610), .A2(KEYINPUT81), .ZN(new_n611));
  NOR2_X1   g186(.A1(new_n610), .A2(KEYINPUT81), .ZN(new_n612));
  NOR2_X1   g187(.A1(new_n611), .A2(new_n612), .ZN(new_n613));
  NAND2_X1  g188(.A1(new_n553), .A2(G92), .ZN(new_n614));
  XNOR2_X1  g189(.A(new_n614), .B(KEYINPUT10), .ZN(new_n615));
  NOR2_X1   g190(.A1(new_n613), .A2(new_n615), .ZN(new_n616));
  OAI21_X1  g191(.A(new_n604), .B1(new_n616), .B2(G868), .ZN(G284));
  OAI21_X1  g192(.A(new_n604), .B1(new_n616), .B2(G868), .ZN(G321));
  XOR2_X1   g193(.A(G299), .B(KEYINPUT82), .Z(new_n619));
  MUX2_X1   g194(.A(new_n619), .B(G286), .S(G868), .Z(G280));
  XNOR2_X1  g195(.A(G280), .B(KEYINPUT83), .ZN(G297));
  XOR2_X1   g196(.A(KEYINPUT84), .B(G559), .Z(new_n622));
  OAI21_X1  g197(.A(new_n616), .B1(G860), .B2(new_n622), .ZN(G148));
  NOR2_X1   g198(.A1(new_n567), .A2(G868), .ZN(new_n624));
  NAND2_X1  g199(.A1(new_n616), .A2(new_n622), .ZN(new_n625));
  AOI21_X1  g200(.A(new_n624), .B1(new_n625), .B2(G868), .ZN(new_n626));
  XNOR2_X1  g201(.A(new_n626), .B(KEYINPUT85), .ZN(G323));
  XNOR2_X1  g202(.A(G323), .B(KEYINPUT11), .ZN(G282));
  OR2_X1    g203(.A1(G99), .A2(G2105), .ZN(new_n629));
  OAI211_X1 g204(.A(new_n629), .B(G2104), .C1(G111), .C2(new_n473), .ZN(new_n630));
  INV_X1    g205(.A(G135), .ZN(new_n631));
  INV_X1    g206(.A(G123), .ZN(new_n632));
  OAI221_X1 g207(.A(new_n630), .B1(new_n474), .B2(new_n631), .C1(new_n632), .C2(new_n486), .ZN(new_n633));
  OR2_X1    g208(.A1(new_n633), .A2(G2096), .ZN(new_n634));
  NAND2_X1  g209(.A1(new_n633), .A2(G2096), .ZN(new_n635));
  NAND3_X1  g210(.A1(new_n473), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n636));
  XNOR2_X1  g211(.A(new_n636), .B(KEYINPUT12), .ZN(new_n637));
  XNOR2_X1  g212(.A(new_n637), .B(KEYINPUT13), .ZN(new_n638));
  XNOR2_X1  g213(.A(new_n638), .B(G2100), .ZN(new_n639));
  NAND3_X1  g214(.A1(new_n634), .A2(new_n635), .A3(new_n639), .ZN(new_n640));
  XOR2_X1   g215(.A(new_n640), .B(KEYINPUT86), .Z(G156));
  XNOR2_X1  g216(.A(G2427), .B(G2438), .ZN(new_n642));
  XNOR2_X1  g217(.A(new_n642), .B(G2430), .ZN(new_n643));
  XNOR2_X1  g218(.A(KEYINPUT15), .B(G2435), .ZN(new_n644));
  OR2_X1    g219(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  NAND2_X1  g220(.A1(new_n643), .A2(new_n644), .ZN(new_n646));
  NAND3_X1  g221(.A1(new_n645), .A2(KEYINPUT14), .A3(new_n646), .ZN(new_n647));
  XNOR2_X1  g222(.A(G1341), .B(G1348), .ZN(new_n648));
  XNOR2_X1  g223(.A(KEYINPUT87), .B(KEYINPUT16), .ZN(new_n649));
  XNOR2_X1  g224(.A(new_n648), .B(new_n649), .ZN(new_n650));
  XNOR2_X1  g225(.A(new_n647), .B(new_n650), .ZN(new_n651));
  XOR2_X1   g226(.A(G2451), .B(G2454), .Z(new_n652));
  XNOR2_X1  g227(.A(G2443), .B(G2446), .ZN(new_n653));
  XNOR2_X1  g228(.A(new_n652), .B(new_n653), .ZN(new_n654));
  OR2_X1    g229(.A1(new_n651), .A2(new_n654), .ZN(new_n655));
  NAND2_X1  g230(.A1(new_n651), .A2(new_n654), .ZN(new_n656));
  NAND3_X1  g231(.A1(new_n655), .A2(G14), .A3(new_n656), .ZN(new_n657));
  XNOR2_X1  g232(.A(new_n657), .B(KEYINPUT88), .ZN(G401));
  XOR2_X1   g233(.A(G2084), .B(G2090), .Z(new_n659));
  XNOR2_X1  g234(.A(G2067), .B(G2678), .ZN(new_n660));
  NAND2_X1  g235(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  AND2_X1   g236(.A1(new_n661), .A2(KEYINPUT17), .ZN(new_n662));
  OR2_X1    g237(.A1(new_n659), .A2(new_n660), .ZN(new_n663));
  AOI21_X1  g238(.A(KEYINPUT18), .B1(new_n662), .B2(new_n663), .ZN(new_n664));
  XOR2_X1   g239(.A(G2072), .B(G2078), .Z(new_n665));
  AOI21_X1  g240(.A(new_n665), .B1(new_n661), .B2(KEYINPUT18), .ZN(new_n666));
  XNOR2_X1  g241(.A(new_n664), .B(new_n666), .ZN(new_n667));
  XOR2_X1   g242(.A(G2096), .B(G2100), .Z(new_n668));
  XNOR2_X1  g243(.A(new_n667), .B(new_n668), .ZN(G227));
  XOR2_X1   g244(.A(G1971), .B(G1976), .Z(new_n670));
  XNOR2_X1  g245(.A(new_n670), .B(KEYINPUT19), .ZN(new_n671));
  XOR2_X1   g246(.A(G1956), .B(G2474), .Z(new_n672));
  XOR2_X1   g247(.A(G1961), .B(G1966), .Z(new_n673));
  NOR2_X1   g248(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  AND2_X1   g249(.A1(new_n671), .A2(new_n674), .ZN(new_n675));
  AND2_X1   g250(.A1(new_n672), .A2(new_n673), .ZN(new_n676));
  NOR3_X1   g251(.A1(new_n671), .A2(new_n676), .A3(new_n674), .ZN(new_n677));
  NAND2_X1  g252(.A1(new_n671), .A2(new_n676), .ZN(new_n678));
  XOR2_X1   g253(.A(KEYINPUT89), .B(KEYINPUT20), .Z(new_n679));
  AOI211_X1 g254(.A(new_n675), .B(new_n677), .C1(new_n678), .C2(new_n679), .ZN(new_n680));
  OAI21_X1  g255(.A(new_n680), .B1(new_n678), .B2(new_n679), .ZN(new_n681));
  INV_X1    g256(.A(KEYINPUT90), .ZN(new_n682));
  XNOR2_X1  g257(.A(new_n681), .B(new_n682), .ZN(new_n683));
  XNOR2_X1  g258(.A(new_n683), .B(KEYINPUT91), .ZN(new_n684));
  XOR2_X1   g259(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n685));
  XNOR2_X1  g260(.A(new_n684), .B(new_n685), .ZN(new_n686));
  XNOR2_X1  g261(.A(G1991), .B(G1996), .ZN(new_n687));
  XNOR2_X1  g262(.A(new_n686), .B(new_n687), .ZN(new_n688));
  XNOR2_X1  g263(.A(G1981), .B(G1986), .ZN(new_n689));
  INV_X1    g264(.A(new_n689), .ZN(new_n690));
  XNOR2_X1  g265(.A(new_n688), .B(new_n690), .ZN(new_n691));
  INV_X1    g266(.A(new_n691), .ZN(G229));
  INV_X1    g267(.A(G29), .ZN(new_n693));
  NAND2_X1  g268(.A1(new_n693), .A2(G35), .ZN(new_n694));
  OAI21_X1  g269(.A(new_n694), .B1(G162), .B2(new_n693), .ZN(new_n695));
  XOR2_X1   g270(.A(new_n695), .B(KEYINPUT29), .Z(new_n696));
  INV_X1    g271(.A(G2090), .ZN(new_n697));
  NOR2_X1   g272(.A1(new_n696), .A2(new_n697), .ZN(new_n698));
  AND2_X1   g273(.A1(new_n698), .A2(KEYINPUT103), .ZN(new_n699));
  NOR2_X1   g274(.A1(new_n698), .A2(KEYINPUT103), .ZN(new_n700));
  INV_X1    g275(.A(G16), .ZN(new_n701));
  NAND2_X1  g276(.A1(new_n701), .A2(G20), .ZN(new_n702));
  XOR2_X1   g277(.A(new_n702), .B(KEYINPUT23), .Z(new_n703));
  AOI21_X1  g278(.A(new_n703), .B1(G299), .B2(G16), .ZN(new_n704));
  XOR2_X1   g279(.A(new_n704), .B(G1956), .Z(new_n705));
  OR3_X1    g280(.A1(new_n699), .A2(new_n700), .A3(new_n705), .ZN(new_n706));
  OR2_X1    g281(.A1(new_n706), .A2(KEYINPUT104), .ZN(new_n707));
  NOR2_X1   g282(.A1(G4), .A2(G16), .ZN(new_n708));
  AOI21_X1  g283(.A(new_n708), .B1(new_n616), .B2(G16), .ZN(new_n709));
  XNOR2_X1  g284(.A(new_n709), .B(KEYINPUT95), .ZN(new_n710));
  XNOR2_X1  g285(.A(KEYINPUT96), .B(G1348), .ZN(new_n711));
  XNOR2_X1  g286(.A(new_n710), .B(new_n711), .ZN(new_n712));
  NAND2_X1  g287(.A1(new_n693), .A2(G26), .ZN(new_n713));
  XOR2_X1   g288(.A(new_n713), .B(KEYINPUT28), .Z(new_n714));
  NAND2_X1  g289(.A1(new_n475), .A2(G140), .ZN(new_n715));
  NAND2_X1  g290(.A1(new_n487), .A2(G128), .ZN(new_n716));
  NOR2_X1   g291(.A1(new_n473), .A2(G116), .ZN(new_n717));
  OAI21_X1  g292(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n718));
  OAI211_X1 g293(.A(new_n715), .B(new_n716), .C1(new_n717), .C2(new_n718), .ZN(new_n719));
  AOI21_X1  g294(.A(new_n714), .B1(new_n719), .B2(G29), .ZN(new_n720));
  XOR2_X1   g295(.A(KEYINPUT97), .B(G2067), .Z(new_n721));
  XNOR2_X1  g296(.A(new_n720), .B(new_n721), .ZN(new_n722));
  XOR2_X1   g297(.A(KEYINPUT31), .B(G11), .Z(new_n723));
  NOR2_X1   g298(.A1(new_n633), .A2(new_n693), .ZN(new_n724));
  XNOR2_X1  g299(.A(KEYINPUT30), .B(G28), .ZN(new_n725));
  AOI211_X1 g300(.A(new_n723), .B(new_n724), .C1(new_n693), .C2(new_n725), .ZN(new_n726));
  AND2_X1   g301(.A1(new_n693), .A2(G32), .ZN(new_n727));
  NAND3_X1  g302(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n728));
  INV_X1    g303(.A(KEYINPUT26), .ZN(new_n729));
  OR2_X1    g304(.A1(new_n728), .A2(new_n729), .ZN(new_n730));
  NAND2_X1  g305(.A1(new_n728), .A2(new_n729), .ZN(new_n731));
  AOI22_X1  g306(.A1(new_n730), .A2(new_n731), .B1(G105), .B2(new_n481), .ZN(new_n732));
  INV_X1    g307(.A(G141), .ZN(new_n733));
  INV_X1    g308(.A(G129), .ZN(new_n734));
  OAI221_X1 g309(.A(new_n732), .B1(new_n474), .B2(new_n733), .C1(new_n734), .C2(new_n486), .ZN(new_n735));
  AOI21_X1  g310(.A(new_n727), .B1(new_n735), .B2(G29), .ZN(new_n736));
  XNOR2_X1  g311(.A(KEYINPUT27), .B(G1996), .ZN(new_n737));
  OR2_X1    g312(.A1(new_n736), .A2(new_n737), .ZN(new_n738));
  INV_X1    g313(.A(G34), .ZN(new_n739));
  AOI21_X1  g314(.A(G29), .B1(new_n739), .B2(KEYINPUT24), .ZN(new_n740));
  OAI21_X1  g315(.A(new_n740), .B1(KEYINPUT24), .B2(new_n739), .ZN(new_n741));
  OAI21_X1  g316(.A(new_n741), .B1(new_n483), .B2(new_n693), .ZN(new_n742));
  INV_X1    g317(.A(G2084), .ZN(new_n743));
  NAND2_X1  g318(.A1(new_n742), .A2(new_n743), .ZN(new_n744));
  OR2_X1    g319(.A1(new_n742), .A2(new_n743), .ZN(new_n745));
  NAND4_X1  g320(.A1(new_n726), .A2(new_n738), .A3(new_n744), .A4(new_n745), .ZN(new_n746));
  INV_X1    g321(.A(G2072), .ZN(new_n747));
  NAND2_X1  g322(.A1(new_n693), .A2(G33), .ZN(new_n748));
  NAND3_X1  g323(.A1(new_n473), .A2(G103), .A3(G2104), .ZN(new_n749));
  INV_X1    g324(.A(KEYINPUT25), .ZN(new_n750));
  XNOR2_X1  g325(.A(new_n749), .B(new_n750), .ZN(new_n751));
  AOI22_X1  g326(.A1(new_n477), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n752));
  OAI21_X1  g327(.A(new_n751), .B1(new_n752), .B2(new_n473), .ZN(new_n753));
  AOI21_X1  g328(.A(new_n753), .B1(new_n475), .B2(G139), .ZN(new_n754));
  OAI21_X1  g329(.A(new_n748), .B1(new_n754), .B2(new_n693), .ZN(new_n755));
  XOR2_X1   g330(.A(new_n755), .B(KEYINPUT98), .Z(new_n756));
  AOI211_X1 g331(.A(new_n722), .B(new_n746), .C1(new_n747), .C2(new_n756), .ZN(new_n757));
  NAND2_X1  g332(.A1(new_n693), .A2(G27), .ZN(new_n758));
  XNOR2_X1  g333(.A(new_n758), .B(KEYINPUT101), .ZN(new_n759));
  OAI21_X1  g334(.A(new_n759), .B1(G164), .B2(new_n693), .ZN(new_n760));
  XOR2_X1   g335(.A(KEYINPUT102), .B(G2078), .Z(new_n761));
  OR2_X1    g336(.A1(new_n760), .A2(new_n761), .ZN(new_n762));
  NAND2_X1  g337(.A1(new_n760), .A2(new_n761), .ZN(new_n763));
  NAND3_X1  g338(.A1(new_n757), .A2(new_n762), .A3(new_n763), .ZN(new_n764));
  NOR2_X1   g339(.A1(G16), .A2(G21), .ZN(new_n765));
  AOI21_X1  g340(.A(new_n765), .B1(G168), .B2(G16), .ZN(new_n766));
  XNOR2_X1  g341(.A(new_n766), .B(G1966), .ZN(new_n767));
  NOR2_X1   g342(.A1(G16), .A2(G19), .ZN(new_n768));
  AOI21_X1  g343(.A(new_n768), .B1(new_n567), .B2(G16), .ZN(new_n769));
  NOR2_X1   g344(.A1(new_n769), .A2(G1341), .ZN(new_n770));
  NAND2_X1  g345(.A1(new_n701), .A2(G5), .ZN(new_n771));
  OAI21_X1  g346(.A(new_n771), .B1(G171), .B2(new_n701), .ZN(new_n772));
  AOI21_X1  g347(.A(new_n770), .B1(G1961), .B2(new_n772), .ZN(new_n773));
  NAND2_X1  g348(.A1(new_n696), .A2(new_n697), .ZN(new_n774));
  OAI211_X1 g349(.A(new_n773), .B(new_n774), .C1(G1961), .C2(new_n772), .ZN(new_n775));
  NOR2_X1   g350(.A1(new_n756), .A2(new_n747), .ZN(new_n776));
  INV_X1    g351(.A(KEYINPUT99), .ZN(new_n777));
  AOI22_X1  g352(.A1(new_n776), .A2(new_n777), .B1(G1341), .B2(new_n769), .ZN(new_n778));
  NAND2_X1  g353(.A1(new_n736), .A2(new_n737), .ZN(new_n779));
  XNOR2_X1  g354(.A(new_n779), .B(KEYINPUT100), .ZN(new_n780));
  OAI211_X1 g355(.A(new_n778), .B(new_n780), .C1(new_n777), .C2(new_n776), .ZN(new_n781));
  NOR4_X1   g356(.A1(new_n764), .A2(new_n767), .A3(new_n775), .A4(new_n781), .ZN(new_n782));
  NAND2_X1  g357(.A1(new_n706), .A2(KEYINPUT104), .ZN(new_n783));
  NAND4_X1  g358(.A1(new_n707), .A2(new_n712), .A3(new_n782), .A4(new_n783), .ZN(new_n784));
  NAND2_X1  g359(.A1(new_n693), .A2(G25), .ZN(new_n785));
  NAND2_X1  g360(.A1(new_n475), .A2(G131), .ZN(new_n786));
  NAND2_X1  g361(.A1(new_n487), .A2(G119), .ZN(new_n787));
  OR2_X1    g362(.A1(G95), .A2(G2105), .ZN(new_n788));
  OAI211_X1 g363(.A(new_n788), .B(G2104), .C1(G107), .C2(new_n473), .ZN(new_n789));
  NAND3_X1  g364(.A1(new_n786), .A2(new_n787), .A3(new_n789), .ZN(new_n790));
  INV_X1    g365(.A(new_n790), .ZN(new_n791));
  OAI21_X1  g366(.A(new_n785), .B1(new_n791), .B2(new_n693), .ZN(new_n792));
  XOR2_X1   g367(.A(KEYINPUT35), .B(G1991), .Z(new_n793));
  XNOR2_X1  g368(.A(new_n792), .B(new_n793), .ZN(new_n794));
  AND2_X1   g369(.A1(new_n701), .A2(G24), .ZN(new_n795));
  AOI21_X1  g370(.A(new_n795), .B1(G290), .B2(G16), .ZN(new_n796));
  XNOR2_X1  g371(.A(KEYINPUT92), .B(G1986), .ZN(new_n797));
  OR2_X1    g372(.A1(new_n796), .A2(new_n797), .ZN(new_n798));
  NAND2_X1  g373(.A1(new_n796), .A2(new_n797), .ZN(new_n799));
  NAND3_X1  g374(.A1(new_n794), .A2(new_n798), .A3(new_n799), .ZN(new_n800));
  NOR2_X1   g375(.A1(G16), .A2(G23), .ZN(new_n801));
  XOR2_X1   g376(.A(new_n801), .B(KEYINPUT94), .Z(new_n802));
  OAI21_X1  g377(.A(new_n802), .B1(G288), .B2(new_n701), .ZN(new_n803));
  XNOR2_X1  g378(.A(new_n803), .B(KEYINPUT33), .ZN(new_n804));
  XNOR2_X1  g379(.A(new_n804), .B(G1976), .ZN(new_n805));
  MUX2_X1   g380(.A(G6), .B(G305), .S(G16), .Z(new_n806));
  XNOR2_X1  g381(.A(KEYINPUT32), .B(G1981), .ZN(new_n807));
  XNOR2_X1  g382(.A(new_n806), .B(new_n807), .ZN(new_n808));
  NAND2_X1  g383(.A1(new_n701), .A2(G22), .ZN(new_n809));
  OAI21_X1  g384(.A(new_n809), .B1(G166), .B2(new_n701), .ZN(new_n810));
  XNOR2_X1  g385(.A(new_n810), .B(G1971), .ZN(new_n811));
  OR2_X1    g386(.A1(new_n808), .A2(new_n811), .ZN(new_n812));
  NOR2_X1   g387(.A1(new_n805), .A2(new_n812), .ZN(new_n813));
  XNOR2_X1  g388(.A(KEYINPUT93), .B(KEYINPUT34), .ZN(new_n814));
  AOI21_X1  g389(.A(new_n800), .B1(new_n813), .B2(new_n814), .ZN(new_n815));
  OAI21_X1  g390(.A(new_n815), .B1(new_n814), .B2(new_n813), .ZN(new_n816));
  NAND2_X1  g391(.A1(new_n816), .A2(KEYINPUT36), .ZN(new_n817));
  INV_X1    g392(.A(KEYINPUT36), .ZN(new_n818));
  OAI211_X1 g393(.A(new_n815), .B(new_n818), .C1(new_n814), .C2(new_n813), .ZN(new_n819));
  AOI21_X1  g394(.A(new_n784), .B1(new_n817), .B2(new_n819), .ZN(G311));
  XNOR2_X1  g395(.A(G311), .B(KEYINPUT105), .ZN(G150));
  NAND2_X1  g396(.A1(new_n616), .A2(G559), .ZN(new_n822));
  XOR2_X1   g397(.A(new_n822), .B(KEYINPUT38), .Z(new_n823));
  NAND2_X1  g398(.A1(new_n562), .A2(new_n566), .ZN(new_n824));
  NAND2_X1  g399(.A1(G80), .A2(G543), .ZN(new_n825));
  INV_X1    g400(.A(G67), .ZN(new_n826));
  OAI21_X1  g401(.A(new_n825), .B1(new_n543), .B2(new_n826), .ZN(new_n827));
  AOI22_X1  g402(.A1(new_n827), .A2(G651), .B1(G55), .B2(new_n521), .ZN(new_n828));
  XNOR2_X1  g403(.A(KEYINPUT106), .B(G93), .ZN(new_n829));
  OAI21_X1  g404(.A(new_n828), .B1(new_n537), .B2(new_n829), .ZN(new_n830));
  XNOR2_X1  g405(.A(new_n824), .B(new_n830), .ZN(new_n831));
  XNOR2_X1  g406(.A(new_n823), .B(new_n831), .ZN(new_n832));
  AND2_X1   g407(.A1(new_n832), .A2(KEYINPUT39), .ZN(new_n833));
  NOR2_X1   g408(.A1(new_n832), .A2(KEYINPUT39), .ZN(new_n834));
  NOR3_X1   g409(.A1(new_n833), .A2(new_n834), .A3(G860), .ZN(new_n835));
  NAND2_X1  g410(.A1(new_n830), .A2(G860), .ZN(new_n836));
  XNOR2_X1  g411(.A(new_n836), .B(KEYINPUT37), .ZN(new_n837));
  OR2_X1    g412(.A1(new_n835), .A2(new_n837), .ZN(G145));
  XNOR2_X1  g413(.A(new_n719), .B(new_n735), .ZN(new_n839));
  XNOR2_X1  g414(.A(new_n637), .B(KEYINPUT107), .ZN(new_n840));
  XNOR2_X1  g415(.A(new_n839), .B(new_n840), .ZN(new_n841));
  NAND2_X1  g416(.A1(new_n475), .A2(G142), .ZN(new_n842));
  NAND2_X1  g417(.A1(new_n487), .A2(G130), .ZN(new_n843));
  NOR2_X1   g418(.A1(new_n473), .A2(G118), .ZN(new_n844));
  OAI21_X1  g419(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n845));
  OAI211_X1 g420(.A(new_n842), .B(new_n843), .C1(new_n844), .C2(new_n845), .ZN(new_n846));
  XNOR2_X1  g421(.A(new_n846), .B(KEYINPUT108), .ZN(new_n847));
  XNOR2_X1  g422(.A(new_n847), .B(new_n790), .ZN(new_n848));
  XNOR2_X1  g423(.A(new_n841), .B(new_n848), .ZN(new_n849));
  OAI21_X1  g424(.A(KEYINPUT67), .B1(new_n469), .B2(G2104), .ZN(new_n850));
  NAND2_X1  g425(.A1(new_n469), .A2(KEYINPUT66), .ZN(new_n851));
  NAND2_X1  g426(.A1(new_n467), .A2(KEYINPUT3), .ZN(new_n852));
  NAND2_X1  g427(.A1(new_n851), .A2(new_n852), .ZN(new_n853));
  AOI21_X1  g428(.A(new_n850), .B1(new_n853), .B2(G2104), .ZN(new_n854));
  AOI211_X1 g429(.A(KEYINPUT67), .B(new_n463), .C1(new_n851), .C2(new_n852), .ZN(new_n855));
  OAI21_X1  g430(.A(new_n503), .B1(new_n854), .B2(new_n855), .ZN(new_n856));
  NAND2_X1  g431(.A1(new_n856), .A2(new_n505), .ZN(new_n857));
  NAND3_X1  g432(.A1(new_n472), .A2(KEYINPUT68), .A3(new_n503), .ZN(new_n858));
  AOI21_X1  g433(.A(new_n500), .B1(new_n857), .B2(new_n858), .ZN(new_n859));
  INV_X1    g434(.A(new_n497), .ZN(new_n860));
  NAND2_X1  g435(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  INV_X1    g436(.A(new_n861), .ZN(new_n862));
  NOR2_X1   g437(.A1(new_n849), .A2(new_n862), .ZN(new_n863));
  INV_X1    g438(.A(new_n863), .ZN(new_n864));
  NAND2_X1  g439(.A1(new_n849), .A2(new_n862), .ZN(new_n865));
  AND3_X1   g440(.A1(new_n864), .A2(new_n754), .A3(new_n865), .ZN(new_n866));
  AOI21_X1  g441(.A(new_n754), .B1(new_n864), .B2(new_n865), .ZN(new_n867));
  XNOR2_X1  g442(.A(new_n633), .B(new_n483), .ZN(new_n868));
  XNOR2_X1  g443(.A(new_n868), .B(new_n491), .ZN(new_n869));
  INV_X1    g444(.A(new_n869), .ZN(new_n870));
  OR3_X1    g445(.A1(new_n866), .A2(new_n867), .A3(new_n870), .ZN(new_n871));
  INV_X1    g446(.A(G37), .ZN(new_n872));
  OAI21_X1  g447(.A(new_n870), .B1(new_n866), .B2(new_n867), .ZN(new_n873));
  NAND3_X1  g448(.A1(new_n871), .A2(new_n872), .A3(new_n873), .ZN(new_n874));
  XNOR2_X1  g449(.A(new_n874), .B(KEYINPUT40), .ZN(G395));
  NOR2_X1   g450(.A1(new_n830), .A2(G868), .ZN(new_n876));
  XNOR2_X1  g451(.A(new_n567), .B(new_n830), .ZN(new_n877));
  XNOR2_X1  g452(.A(new_n625), .B(new_n877), .ZN(new_n878));
  NAND2_X1  g453(.A1(new_n616), .A2(G299), .ZN(new_n879));
  INV_X1    g454(.A(G299), .ZN(new_n880));
  OAI21_X1  g455(.A(new_n880), .B1(new_n613), .B2(new_n615), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n879), .A2(new_n881), .ZN(new_n882));
  INV_X1    g457(.A(new_n882), .ZN(new_n883));
  NOR2_X1   g458(.A1(new_n878), .A2(new_n883), .ZN(new_n884));
  XNOR2_X1  g459(.A(new_n884), .B(KEYINPUT109), .ZN(new_n885));
  NAND3_X1  g460(.A1(new_n879), .A2(KEYINPUT110), .A3(new_n881), .ZN(new_n886));
  INV_X1    g461(.A(KEYINPUT41), .ZN(new_n887));
  OR2_X1    g462(.A1(new_n881), .A2(KEYINPUT110), .ZN(new_n888));
  NAND3_X1  g463(.A1(new_n886), .A2(new_n887), .A3(new_n888), .ZN(new_n889));
  OAI21_X1  g464(.A(KEYINPUT111), .B1(new_n882), .B2(new_n887), .ZN(new_n890));
  INV_X1    g465(.A(KEYINPUT111), .ZN(new_n891));
  NAND4_X1  g466(.A1(new_n879), .A2(new_n891), .A3(KEYINPUT41), .A4(new_n881), .ZN(new_n892));
  NAND3_X1  g467(.A1(new_n889), .A2(new_n890), .A3(new_n892), .ZN(new_n893));
  NAND2_X1  g468(.A1(new_n893), .A2(new_n878), .ZN(new_n894));
  XNOR2_X1  g469(.A(G288), .B(G305), .ZN(new_n895));
  XNOR2_X1  g470(.A(G166), .B(G290), .ZN(new_n896));
  XNOR2_X1  g471(.A(new_n895), .B(new_n896), .ZN(new_n897));
  XOR2_X1   g472(.A(new_n897), .B(KEYINPUT42), .Z(new_n898));
  NAND3_X1  g473(.A1(new_n885), .A2(new_n894), .A3(new_n898), .ZN(new_n899));
  NAND2_X1  g474(.A1(new_n899), .A2(KEYINPUT112), .ZN(new_n900));
  AOI21_X1  g475(.A(new_n898), .B1(new_n885), .B2(new_n894), .ZN(new_n901));
  XNOR2_X1  g476(.A(new_n900), .B(new_n901), .ZN(new_n902));
  AOI21_X1  g477(.A(new_n876), .B1(new_n902), .B2(G868), .ZN(G295));
  AOI21_X1  g478(.A(new_n876), .B1(new_n902), .B2(G868), .ZN(G331));
  NAND2_X1  g479(.A1(new_n877), .A2(G168), .ZN(new_n905));
  NAND2_X1  g480(.A1(G286), .A2(new_n831), .ZN(new_n906));
  AND3_X1   g481(.A1(new_n905), .A2(G171), .A3(new_n906), .ZN(new_n907));
  AOI21_X1  g482(.A(G171), .B1(new_n905), .B2(new_n906), .ZN(new_n908));
  OR2_X1    g483(.A1(new_n907), .A2(new_n908), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n893), .A2(new_n909), .ZN(new_n910));
  INV_X1    g485(.A(KEYINPUT113), .ZN(new_n911));
  NOR2_X1   g486(.A1(new_n907), .A2(new_n908), .ZN(new_n912));
  AOI21_X1  g487(.A(new_n911), .B1(new_n912), .B2(new_n882), .ZN(new_n913));
  NAND2_X1  g488(.A1(new_n910), .A2(new_n913), .ZN(new_n914));
  NAND3_X1  g489(.A1(new_n893), .A2(new_n909), .A3(new_n911), .ZN(new_n915));
  AOI21_X1  g490(.A(new_n897), .B1(new_n914), .B2(new_n915), .ZN(new_n916));
  NOR2_X1   g491(.A1(new_n916), .A2(G37), .ZN(new_n917));
  NAND3_X1  g492(.A1(new_n914), .A2(new_n897), .A3(new_n915), .ZN(new_n918));
  AOI21_X1  g493(.A(KEYINPUT43), .B1(new_n917), .B2(new_n918), .ZN(new_n919));
  OAI21_X1  g494(.A(KEYINPUT41), .B1(new_n907), .B2(new_n908), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n886), .A2(new_n888), .ZN(new_n921));
  OAI21_X1  g496(.A(new_n897), .B1(new_n920), .B2(new_n921), .ZN(new_n922));
  AOI21_X1  g497(.A(new_n922), .B1(new_n883), .B2(new_n920), .ZN(new_n923));
  INV_X1    g498(.A(KEYINPUT43), .ZN(new_n924));
  NOR4_X1   g499(.A1(new_n916), .A2(new_n923), .A3(new_n924), .A4(G37), .ZN(new_n925));
  OAI21_X1  g500(.A(KEYINPUT44), .B1(new_n919), .B2(new_n925), .ZN(new_n926));
  INV_X1    g501(.A(KEYINPUT44), .ZN(new_n927));
  AOI21_X1  g502(.A(new_n924), .B1(new_n917), .B2(new_n918), .ZN(new_n928));
  NOR4_X1   g503(.A1(new_n916), .A2(new_n923), .A3(KEYINPUT43), .A4(G37), .ZN(new_n929));
  OAI21_X1  g504(.A(new_n927), .B1(new_n928), .B2(new_n929), .ZN(new_n930));
  NAND2_X1  g505(.A1(new_n926), .A2(new_n930), .ZN(G397));
  INV_X1    g506(.A(KEYINPUT124), .ZN(new_n932));
  XNOR2_X1  g507(.A(KEYINPUT116), .B(G8), .ZN(new_n933));
  INV_X1    g508(.A(new_n933), .ZN(new_n934));
  NAND2_X1  g509(.A1(G286), .A2(new_n934), .ZN(new_n935));
  INV_X1    g510(.A(KEYINPUT51), .ZN(new_n936));
  NAND2_X1  g511(.A1(new_n935), .A2(new_n936), .ZN(new_n937));
  INV_X1    g512(.A(new_n937), .ZN(new_n938));
  NAND3_X1  g513(.A1(new_n476), .A2(G40), .A3(new_n482), .ZN(new_n939));
  INV_X1    g514(.A(new_n939), .ZN(new_n940));
  AOI21_X1  g515(.A(G1384), .B1(new_n859), .B2(new_n860), .ZN(new_n941));
  OAI21_X1  g516(.A(new_n940), .B1(new_n941), .B2(KEYINPUT45), .ZN(new_n942));
  NAND2_X1  g517(.A1(new_n857), .A2(new_n858), .ZN(new_n943));
  AOI21_X1  g518(.A(KEYINPUT69), .B1(new_n943), .B2(new_n501), .ZN(new_n944));
  INV_X1    g519(.A(new_n510), .ZN(new_n945));
  OAI21_X1  g520(.A(new_n860), .B1(new_n944), .B2(new_n945), .ZN(new_n946));
  INV_X1    g521(.A(G1384), .ZN(new_n947));
  NAND3_X1  g522(.A1(new_n946), .A2(KEYINPUT45), .A3(new_n947), .ZN(new_n948));
  AOI21_X1  g523(.A(new_n942), .B1(new_n948), .B2(KEYINPUT118), .ZN(new_n949));
  NAND2_X1  g524(.A1(new_n509), .A2(new_n510), .ZN(new_n950));
  AOI21_X1  g525(.A(G1384), .B1(new_n950), .B2(new_n860), .ZN(new_n951));
  INV_X1    g526(.A(KEYINPUT118), .ZN(new_n952));
  NAND3_X1  g527(.A1(new_n951), .A2(new_n952), .A3(KEYINPUT45), .ZN(new_n953));
  AOI21_X1  g528(.A(G1966), .B1(new_n949), .B2(new_n953), .ZN(new_n954));
  INV_X1    g529(.A(KEYINPUT50), .ZN(new_n955));
  NAND2_X1  g530(.A1(new_n941), .A2(new_n955), .ZN(new_n956));
  OAI211_X1 g531(.A(new_n956), .B(new_n940), .C1(new_n951), .C2(new_n955), .ZN(new_n957));
  NOR2_X1   g532(.A1(new_n957), .A2(G2084), .ZN(new_n958));
  NOR2_X1   g533(.A1(new_n954), .A2(new_n958), .ZN(new_n959));
  OAI21_X1  g534(.A(new_n938), .B1(new_n959), .B2(new_n933), .ZN(new_n960));
  NOR2_X1   g535(.A1(G168), .A2(new_n933), .ZN(new_n961));
  NAND2_X1  g536(.A1(new_n956), .A2(new_n940), .ZN(new_n962));
  NAND2_X1  g537(.A1(new_n946), .A2(new_n947), .ZN(new_n963));
  AOI21_X1  g538(.A(new_n962), .B1(new_n963), .B2(KEYINPUT50), .ZN(new_n964));
  NAND2_X1  g539(.A1(new_n964), .A2(new_n743), .ZN(new_n965));
  AOI21_X1  g540(.A(new_n952), .B1(new_n951), .B2(KEYINPUT45), .ZN(new_n966));
  INV_X1    g541(.A(KEYINPUT45), .ZN(new_n967));
  NOR4_X1   g542(.A1(G164), .A2(KEYINPUT118), .A3(new_n967), .A4(G1384), .ZN(new_n968));
  NOR3_X1   g543(.A1(new_n966), .A2(new_n968), .A3(new_n942), .ZN(new_n969));
  OAI21_X1  g544(.A(new_n965), .B1(new_n969), .B2(G1966), .ZN(new_n970));
  AOI21_X1  g545(.A(new_n961), .B1(new_n970), .B2(G8), .ZN(new_n971));
  OAI21_X1  g546(.A(new_n960), .B1(new_n971), .B2(new_n936), .ZN(new_n972));
  NAND2_X1  g547(.A1(new_n970), .A2(new_n961), .ZN(new_n973));
  AOI21_X1  g548(.A(new_n932), .B1(new_n972), .B2(new_n973), .ZN(new_n974));
  OAI21_X1  g549(.A(G8), .B1(new_n954), .B2(new_n958), .ZN(new_n975));
  AOI21_X1  g550(.A(new_n936), .B1(new_n975), .B2(new_n935), .ZN(new_n976));
  AOI21_X1  g551(.A(new_n937), .B1(new_n970), .B2(new_n934), .ZN(new_n977));
  OAI211_X1 g552(.A(new_n932), .B(new_n973), .C1(new_n976), .C2(new_n977), .ZN(new_n978));
  INV_X1    g553(.A(new_n978), .ZN(new_n979));
  OAI21_X1  g554(.A(KEYINPUT62), .B1(new_n974), .B2(new_n979), .ZN(new_n980));
  NOR2_X1   g555(.A1(new_n976), .A2(new_n977), .ZN(new_n981));
  INV_X1    g556(.A(new_n973), .ZN(new_n982));
  OAI21_X1  g557(.A(KEYINPUT124), .B1(new_n981), .B2(new_n982), .ZN(new_n983));
  INV_X1    g558(.A(KEYINPUT62), .ZN(new_n984));
  NAND3_X1  g559(.A1(new_n983), .A2(new_n984), .A3(new_n978), .ZN(new_n985));
  INV_X1    g560(.A(G8), .ZN(new_n986));
  NAND2_X1  g561(.A1(new_n963), .A2(new_n967), .ZN(new_n987));
  XNOR2_X1  g562(.A(KEYINPUT114), .B(G1384), .ZN(new_n988));
  AOI21_X1  g563(.A(new_n988), .B1(new_n859), .B2(new_n860), .ZN(new_n989));
  AOI21_X1  g564(.A(new_n939), .B1(new_n989), .B2(KEYINPUT45), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n987), .A2(new_n990), .ZN(new_n991));
  INV_X1    g566(.A(G1971), .ZN(new_n992));
  NAND2_X1  g567(.A1(new_n991), .A2(new_n992), .ZN(new_n993));
  XOR2_X1   g568(.A(KEYINPUT115), .B(G2090), .Z(new_n994));
  NAND2_X1  g569(.A1(new_n964), .A2(new_n994), .ZN(new_n995));
  AOI21_X1  g570(.A(new_n986), .B1(new_n993), .B2(new_n995), .ZN(new_n996));
  NAND2_X1  g571(.A1(G303), .A2(G8), .ZN(new_n997));
  XOR2_X1   g572(.A(new_n997), .B(KEYINPUT55), .Z(new_n998));
  NAND2_X1  g573(.A1(new_n996), .A2(new_n998), .ZN(new_n999));
  NAND2_X1  g574(.A1(new_n941), .A2(new_n940), .ZN(new_n1000));
  NAND2_X1  g575(.A1(new_n1000), .A2(new_n934), .ZN(new_n1001));
  AND2_X1   g576(.A1(new_n586), .A2(new_n590), .ZN(new_n1002));
  AOI21_X1  g577(.A(new_n1001), .B1(new_n1002), .B2(G1976), .ZN(new_n1003));
  INV_X1    g578(.A(KEYINPUT52), .ZN(new_n1004));
  OR2_X1    g579(.A1(new_n1003), .A2(new_n1004), .ZN(new_n1005));
  OAI211_X1 g580(.A(new_n1003), .B(new_n1004), .C1(G1976), .C2(new_n1002), .ZN(new_n1006));
  INV_X1    g581(.A(G1981), .ZN(new_n1007));
  XOR2_X1   g582(.A(KEYINPUT117), .B(G86), .Z(new_n1008));
  NAND2_X1  g583(.A1(new_n553), .A2(new_n1008), .ZN(new_n1009));
  AOI21_X1  g584(.A(new_n1007), .B1(new_n1009), .B2(new_n595), .ZN(new_n1010));
  NOR2_X1   g585(.A1(G305), .A2(G1981), .ZN(new_n1011));
  INV_X1    g586(.A(KEYINPUT49), .ZN(new_n1012));
  OR3_X1    g587(.A1(new_n1010), .A2(new_n1011), .A3(new_n1012), .ZN(new_n1013));
  OAI21_X1  g588(.A(new_n1012), .B1(new_n1010), .B2(new_n1011), .ZN(new_n1014));
  NAND4_X1  g589(.A1(new_n1013), .A2(new_n934), .A3(new_n1000), .A4(new_n1014), .ZN(new_n1015));
  AND3_X1   g590(.A1(new_n1005), .A2(new_n1006), .A3(new_n1015), .ZN(new_n1016));
  OAI21_X1  g591(.A(new_n940), .B1(new_n941), .B2(new_n955), .ZN(new_n1017));
  AOI21_X1  g592(.A(new_n1017), .B1(new_n951), .B2(new_n955), .ZN(new_n1018));
  NAND2_X1  g593(.A1(new_n1018), .A2(new_n994), .ZN(new_n1019));
  AOI21_X1  g594(.A(new_n933), .B1(new_n993), .B2(new_n1019), .ZN(new_n1020));
  OAI211_X1 g595(.A(new_n999), .B(new_n1016), .C1(new_n998), .C2(new_n1020), .ZN(new_n1021));
  INV_X1    g596(.A(G2078), .ZN(new_n1022));
  NAND3_X1  g597(.A1(new_n987), .A2(new_n1022), .A3(new_n990), .ZN(new_n1023));
  INV_X1    g598(.A(KEYINPUT53), .ZN(new_n1024));
  NAND2_X1  g599(.A1(new_n1023), .A2(new_n1024), .ZN(new_n1025));
  INV_X1    g600(.A(G1961), .ZN(new_n1026));
  NAND2_X1  g601(.A1(new_n957), .A2(new_n1026), .ZN(new_n1027));
  NAND2_X1  g602(.A1(new_n1025), .A2(new_n1027), .ZN(new_n1028));
  NAND3_X1  g603(.A1(new_n949), .A2(new_n1022), .A3(new_n953), .ZN(new_n1029));
  INV_X1    g604(.A(KEYINPUT125), .ZN(new_n1030));
  AOI21_X1  g605(.A(new_n1024), .B1(new_n1029), .B2(new_n1030), .ZN(new_n1031));
  NAND3_X1  g606(.A1(new_n969), .A2(KEYINPUT125), .A3(new_n1022), .ZN(new_n1032));
  AOI21_X1  g607(.A(new_n1028), .B1(new_n1031), .B2(new_n1032), .ZN(new_n1033));
  NOR3_X1   g608(.A1(new_n1021), .A2(G301), .A3(new_n1033), .ZN(new_n1034));
  NAND3_X1  g609(.A1(new_n980), .A2(new_n985), .A3(new_n1034), .ZN(new_n1035));
  NAND2_X1  g610(.A1(new_n1035), .A2(KEYINPUT127), .ZN(new_n1036));
  INV_X1    g611(.A(KEYINPUT127), .ZN(new_n1037));
  NAND4_X1  g612(.A1(new_n980), .A2(new_n985), .A3(new_n1037), .A4(new_n1034), .ZN(new_n1038));
  INV_X1    g613(.A(KEYINPUT63), .ZN(new_n1039));
  NOR3_X1   g614(.A1(new_n959), .A2(G286), .A3(new_n933), .ZN(new_n1040));
  INV_X1    g615(.A(new_n1040), .ZN(new_n1041));
  OAI21_X1  g616(.A(new_n1039), .B1(new_n1021), .B2(new_n1041), .ZN(new_n1042));
  NOR2_X1   g617(.A1(new_n996), .A2(new_n998), .ZN(new_n1043));
  NOR2_X1   g618(.A1(new_n1043), .A2(new_n1039), .ZN(new_n1044));
  NAND4_X1  g619(.A1(new_n1044), .A2(new_n999), .A3(new_n1016), .A4(new_n1040), .ZN(new_n1045));
  NAND2_X1  g620(.A1(new_n1042), .A2(new_n1045), .ZN(new_n1046));
  INV_X1    g621(.A(G1976), .ZN(new_n1047));
  NAND3_X1  g622(.A1(new_n1015), .A2(new_n1047), .A3(new_n1002), .ZN(new_n1048));
  INV_X1    g623(.A(new_n1011), .ZN(new_n1049));
  AOI21_X1  g624(.A(new_n1001), .B1(new_n1048), .B2(new_n1049), .ZN(new_n1050));
  INV_X1    g625(.A(new_n999), .ZN(new_n1051));
  AOI21_X1  g626(.A(new_n1050), .B1(new_n1051), .B2(new_n1016), .ZN(new_n1052));
  NAND2_X1  g627(.A1(new_n1046), .A2(new_n1052), .ZN(new_n1053));
  INV_X1    g628(.A(KEYINPUT119), .ZN(new_n1054));
  NAND2_X1  g629(.A1(new_n1054), .A2(KEYINPUT57), .ZN(new_n1055));
  NOR2_X1   g630(.A1(new_n1054), .A2(KEYINPUT57), .ZN(new_n1056));
  INV_X1    g631(.A(new_n1056), .ZN(new_n1057));
  NAND3_X1  g632(.A1(G299), .A2(new_n1055), .A3(new_n1057), .ZN(new_n1058));
  INV_X1    g633(.A(new_n1058), .ZN(new_n1059));
  AOI21_X1  g634(.A(new_n1057), .B1(G299), .B2(new_n1055), .ZN(new_n1060));
  NOR2_X1   g635(.A1(new_n1059), .A2(new_n1060), .ZN(new_n1061));
  XNOR2_X1  g636(.A(KEYINPUT56), .B(G2072), .ZN(new_n1062));
  OAI211_X1 g637(.A(new_n990), .B(new_n1062), .C1(new_n951), .C2(KEYINPUT45), .ZN(new_n1063));
  OAI211_X1 g638(.A(new_n1061), .B(new_n1063), .C1(new_n1018), .C2(G1956), .ZN(new_n1064));
  OAI21_X1  g639(.A(KEYINPUT120), .B1(new_n1059), .B2(new_n1060), .ZN(new_n1065));
  OR3_X1    g640(.A1(G299), .A2(new_n1054), .A3(KEYINPUT57), .ZN(new_n1066));
  INV_X1    g641(.A(KEYINPUT120), .ZN(new_n1067));
  NAND3_X1  g642(.A1(new_n1066), .A2(new_n1067), .A3(new_n1058), .ZN(new_n1068));
  NAND2_X1  g643(.A1(new_n1065), .A2(new_n1068), .ZN(new_n1069));
  OAI21_X1  g644(.A(new_n1063), .B1(new_n1018), .B2(G1956), .ZN(new_n1070));
  AND2_X1   g645(.A1(new_n1069), .A2(new_n1070), .ZN(new_n1071));
  NOR2_X1   g646(.A1(new_n1000), .A2(G2067), .ZN(new_n1072));
  AOI21_X1  g647(.A(new_n1072), .B1(new_n957), .B2(new_n711), .ZN(new_n1073));
  OR2_X1    g648(.A1(new_n613), .A2(new_n615), .ZN(new_n1074));
  NOR2_X1   g649(.A1(new_n1073), .A2(new_n1074), .ZN(new_n1075));
  OAI21_X1  g650(.A(new_n1064), .B1(new_n1071), .B2(new_n1075), .ZN(new_n1076));
  NAND2_X1  g651(.A1(new_n1076), .A2(KEYINPUT121), .ZN(new_n1077));
  INV_X1    g652(.A(KEYINPUT121), .ZN(new_n1078));
  OAI211_X1 g653(.A(new_n1078), .B(new_n1064), .C1(new_n1071), .C2(new_n1075), .ZN(new_n1079));
  NAND2_X1  g654(.A1(new_n1077), .A2(new_n1079), .ZN(new_n1080));
  INV_X1    g655(.A(new_n1061), .ZN(new_n1081));
  NAND2_X1  g656(.A1(new_n1070), .A2(new_n1081), .ZN(new_n1082));
  NAND2_X1  g657(.A1(new_n1082), .A2(new_n1064), .ZN(new_n1083));
  INV_X1    g658(.A(KEYINPUT61), .ZN(new_n1084));
  NOR2_X1   g659(.A1(new_n1074), .A2(KEYINPUT60), .ZN(new_n1085));
  AOI22_X1  g660(.A1(new_n1083), .A2(new_n1084), .B1(new_n1073), .B2(new_n1085), .ZN(new_n1086));
  AND2_X1   g661(.A1(new_n1073), .A2(new_n1074), .ZN(new_n1087));
  OAI21_X1  g662(.A(KEYINPUT60), .B1(new_n1087), .B2(new_n1075), .ZN(new_n1088));
  INV_X1    g663(.A(KEYINPUT122), .ZN(new_n1089));
  INV_X1    g664(.A(G1996), .ZN(new_n1090));
  NAND4_X1  g665(.A1(new_n987), .A2(new_n1089), .A3(new_n1090), .A4(new_n990), .ZN(new_n1091));
  OAI211_X1 g666(.A(new_n1090), .B(new_n990), .C1(new_n951), .C2(KEYINPUT45), .ZN(new_n1092));
  NAND2_X1  g667(.A1(new_n1092), .A2(KEYINPUT122), .ZN(new_n1093));
  XOR2_X1   g668(.A(KEYINPUT58), .B(G1341), .Z(new_n1094));
  NAND2_X1  g669(.A1(new_n1000), .A2(new_n1094), .ZN(new_n1095));
  NAND3_X1  g670(.A1(new_n1091), .A2(new_n1093), .A3(new_n1095), .ZN(new_n1096));
  NAND2_X1  g671(.A1(new_n1096), .A2(new_n567), .ZN(new_n1097));
  INV_X1    g672(.A(KEYINPUT59), .ZN(new_n1098));
  NAND2_X1  g673(.A1(new_n1097), .A2(new_n1098), .ZN(new_n1099));
  NAND3_X1  g674(.A1(new_n1096), .A2(KEYINPUT59), .A3(new_n567), .ZN(new_n1100));
  NAND4_X1  g675(.A1(new_n1086), .A2(new_n1088), .A3(new_n1099), .A4(new_n1100), .ZN(new_n1101));
  AOI21_X1  g676(.A(new_n1084), .B1(new_n1069), .B2(new_n1070), .ZN(new_n1102));
  AND3_X1   g677(.A1(new_n1102), .A2(KEYINPUT123), .A3(new_n1064), .ZN(new_n1103));
  AOI21_X1  g678(.A(KEYINPUT123), .B1(new_n1102), .B2(new_n1064), .ZN(new_n1104));
  NOR2_X1   g679(.A1(new_n1103), .A2(new_n1104), .ZN(new_n1105));
  OAI21_X1  g680(.A(new_n1080), .B1(new_n1101), .B2(new_n1105), .ZN(new_n1106));
  OAI21_X1  g681(.A(new_n967), .B1(new_n862), .B2(new_n988), .ZN(new_n1107));
  NAND4_X1  g682(.A1(new_n1107), .A2(new_n990), .A3(KEYINPUT53), .A4(new_n1022), .ZN(new_n1108));
  NAND3_X1  g683(.A1(new_n1025), .A2(new_n1027), .A3(new_n1108), .ZN(new_n1109));
  OR2_X1    g684(.A1(new_n1109), .A2(G171), .ZN(new_n1110));
  OAI21_X1  g685(.A(new_n1110), .B1(new_n1033), .B2(G301), .ZN(new_n1111));
  INV_X1    g686(.A(KEYINPUT54), .ZN(new_n1112));
  AOI21_X1  g687(.A(new_n1021), .B1(new_n1111), .B2(new_n1112), .ZN(new_n1113));
  AND2_X1   g688(.A1(new_n1106), .A2(new_n1113), .ZN(new_n1114));
  NAND2_X1  g689(.A1(new_n1033), .A2(G301), .ZN(new_n1115));
  OR2_X1    g690(.A1(new_n1115), .A2(KEYINPUT126), .ZN(new_n1116));
  NAND2_X1  g691(.A1(new_n1109), .A2(G171), .ZN(new_n1117));
  NAND2_X1  g692(.A1(new_n1117), .A2(KEYINPUT54), .ZN(new_n1118));
  AOI21_X1  g693(.A(new_n1118), .B1(new_n1115), .B2(KEYINPUT126), .ZN(new_n1119));
  AOI22_X1  g694(.A1(new_n983), .A2(new_n978), .B1(new_n1116), .B2(new_n1119), .ZN(new_n1120));
  AOI21_X1  g695(.A(new_n1053), .B1(new_n1114), .B2(new_n1120), .ZN(new_n1121));
  NAND3_X1  g696(.A1(new_n1036), .A2(new_n1038), .A3(new_n1121), .ZN(new_n1122));
  NOR2_X1   g697(.A1(new_n1107), .A2(new_n939), .ZN(new_n1123));
  XOR2_X1   g698(.A(new_n719), .B(G2067), .Z(new_n1124));
  XNOR2_X1  g699(.A(new_n735), .B(new_n1090), .ZN(new_n1125));
  NAND2_X1  g700(.A1(new_n1124), .A2(new_n1125), .ZN(new_n1126));
  XOR2_X1   g701(.A(new_n790), .B(new_n793), .Z(new_n1127));
  NOR2_X1   g702(.A1(new_n1126), .A2(new_n1127), .ZN(new_n1128));
  INV_X1    g703(.A(new_n1128), .ZN(new_n1129));
  XNOR2_X1  g704(.A(G290), .B(G1986), .ZN(new_n1130));
  OAI21_X1  g705(.A(new_n1123), .B1(new_n1129), .B2(new_n1130), .ZN(new_n1131));
  NAND2_X1  g706(.A1(new_n1122), .A2(new_n1131), .ZN(new_n1132));
  INV_X1    g707(.A(new_n1123), .ZN(new_n1133));
  OR3_X1    g708(.A1(new_n1133), .A2(G1986), .A3(G290), .ZN(new_n1134));
  INV_X1    g709(.A(new_n1134), .ZN(new_n1135));
  AOI22_X1  g710(.A1(new_n1135), .A2(KEYINPUT48), .B1(new_n1129), .B2(new_n1123), .ZN(new_n1136));
  OAI21_X1  g711(.A(new_n1136), .B1(KEYINPUT48), .B2(new_n1135), .ZN(new_n1137));
  INV_X1    g712(.A(KEYINPUT46), .ZN(new_n1138));
  OAI21_X1  g713(.A(new_n1138), .B1(new_n1133), .B2(G1996), .ZN(new_n1139));
  NAND3_X1  g714(.A1(new_n1123), .A2(KEYINPUT46), .A3(new_n1090), .ZN(new_n1140));
  INV_X1    g715(.A(new_n1124), .ZN(new_n1141));
  OAI21_X1  g716(.A(new_n1123), .B1(new_n1141), .B2(new_n735), .ZN(new_n1142));
  NAND3_X1  g717(.A1(new_n1139), .A2(new_n1140), .A3(new_n1142), .ZN(new_n1143));
  XNOR2_X1  g718(.A(new_n1143), .B(KEYINPUT47), .ZN(new_n1144));
  NAND2_X1  g719(.A1(new_n791), .A2(new_n793), .ZN(new_n1145));
  OAI22_X1  g720(.A1(new_n1126), .A2(new_n1145), .B1(G2067), .B2(new_n719), .ZN(new_n1146));
  NAND2_X1  g721(.A1(new_n1146), .A2(new_n1123), .ZN(new_n1147));
  AND3_X1   g722(.A1(new_n1137), .A2(new_n1144), .A3(new_n1147), .ZN(new_n1148));
  NAND2_X1  g723(.A1(new_n1132), .A2(new_n1148), .ZN(G329));
  assign    G231 = 1'b0;
  NOR2_X1   g724(.A1(new_n928), .A2(new_n929), .ZN(new_n1151));
  INV_X1    g725(.A(new_n657), .ZN(new_n1152));
  NOR3_X1   g726(.A1(new_n1152), .A2(new_n460), .A3(G227), .ZN(new_n1153));
  NAND3_X1  g727(.A1(new_n874), .A2(new_n691), .A3(new_n1153), .ZN(new_n1154));
  NOR2_X1   g728(.A1(new_n1151), .A2(new_n1154), .ZN(G308));
  AND2_X1   g729(.A1(new_n691), .A2(new_n1153), .ZN(new_n1156));
  OAI211_X1 g730(.A(new_n1156), .B(new_n874), .C1(new_n928), .C2(new_n929), .ZN(G225));
endmodule


