//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 1 0 1 1 1 0 1 0 0 0 1 1 1 1 0 0 1 1 1 0 0 1 0 0 1 0 1 0 0 1 1 0 1 0 0 0 1 0 1 0 0 0 0 0 1 1 1 1 0 1 0 0 1 0 1 1 1 1 1 0 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:28:43 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n455, new_n456, new_n457,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n498, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n517, new_n518,
    new_n519, new_n520, new_n521, new_n522, new_n523, new_n524, new_n525,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n535,
    new_n536, new_n537, new_n538, new_n539, new_n540, new_n541, new_n542,
    new_n543, new_n545, new_n546, new_n548, new_n549, new_n551, new_n552,
    new_n553, new_n554, new_n555, new_n556, new_n557, new_n558, new_n559,
    new_n560, new_n561, new_n562, new_n563, new_n564, new_n568, new_n569,
    new_n571, new_n572, new_n573, new_n574, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n596, new_n598,
    new_n599, new_n600, new_n602, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n619, new_n620, new_n621, new_n622,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n638, new_n639, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n806, new_n807, new_n808, new_n809, new_n810,
    new_n811, new_n812, new_n813, new_n814, new_n815, new_n816, new_n817,
    new_n818, new_n819, new_n820, new_n821, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n890, new_n891,
    new_n892, new_n893, new_n894, new_n895, new_n896, new_n897, new_n898,
    new_n899, new_n900, new_n901, new_n902, new_n903, new_n904, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n450));
  XNOR2_X1  g025(.A(new_n450), .B(KEYINPUT2), .ZN(new_n451));
  NOR4_X1   g026(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n452));
  NAND2_X1  g027(.A1(new_n451), .A2(new_n452), .ZN(G261));
  INV_X1    g028(.A(G261), .ZN(G325));
  INV_X1    g029(.A(G2106), .ZN(new_n455));
  INV_X1    g030(.A(G567), .ZN(new_n456));
  OAI22_X1  g031(.A1(new_n451), .A2(new_n455), .B1(new_n456), .B2(new_n452), .ZN(new_n457));
  XNOR2_X1  g032(.A(new_n457), .B(KEYINPUT64), .ZN(G319));
  INV_X1    g033(.A(KEYINPUT65), .ZN(new_n459));
  AND2_X1   g034(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n460));
  NOR2_X1   g035(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n461));
  OAI211_X1 g036(.A(new_n459), .B(G125), .C1(new_n460), .C2(new_n461), .ZN(new_n462));
  NAND2_X1  g037(.A1(G113), .A2(G2104), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  XNOR2_X1  g039(.A(KEYINPUT3), .B(G2104), .ZN(new_n465));
  AOI21_X1  g040(.A(new_n459), .B1(new_n465), .B2(G125), .ZN(new_n466));
  OAI21_X1  g041(.A(G2105), .B1(new_n464), .B2(new_n466), .ZN(new_n467));
  NOR2_X1   g042(.A1(new_n460), .A2(new_n461), .ZN(new_n468));
  NOR2_X1   g043(.A1(new_n468), .A2(G2105), .ZN(new_n469));
  INV_X1    g044(.A(G2104), .ZN(new_n470));
  NOR2_X1   g045(.A1(new_n470), .A2(G2105), .ZN(new_n471));
  AOI22_X1  g046(.A1(new_n469), .A2(G137), .B1(G101), .B2(new_n471), .ZN(new_n472));
  AND2_X1   g047(.A1(new_n467), .A2(new_n472), .ZN(G160));
  XNOR2_X1  g048(.A(new_n469), .B(KEYINPUT66), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n474), .A2(G136), .ZN(new_n475));
  INV_X1    g050(.A(G2105), .ZN(new_n476));
  NOR2_X1   g051(.A1(new_n468), .A2(new_n476), .ZN(new_n477));
  MUX2_X1   g052(.A(G100), .B(G112), .S(G2105), .Z(new_n478));
  AOI22_X1  g053(.A1(new_n477), .A2(G124), .B1(G2104), .B2(new_n478), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n475), .A2(new_n479), .ZN(new_n480));
  INV_X1    g055(.A(new_n480), .ZN(G162));
  INV_X1    g056(.A(G126), .ZN(new_n482));
  OR2_X1    g057(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n483));
  NAND2_X1  g058(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n484));
  AOI21_X1  g059(.A(new_n482), .B1(new_n483), .B2(new_n484), .ZN(new_n485));
  AND2_X1   g060(.A1(G114), .A2(G2104), .ZN(new_n486));
  OAI21_X1  g061(.A(G2105), .B1(new_n485), .B2(new_n486), .ZN(new_n487));
  NAND2_X1  g062(.A1(KEYINPUT4), .A2(G138), .ZN(new_n488));
  AOI21_X1  g063(.A(new_n488), .B1(new_n483), .B2(new_n484), .ZN(new_n489));
  NAND2_X1  g064(.A1(G102), .A2(G2104), .ZN(new_n490));
  INV_X1    g065(.A(new_n490), .ZN(new_n491));
  OAI21_X1  g066(.A(new_n476), .B1(new_n489), .B2(new_n491), .ZN(new_n492));
  OAI211_X1 g067(.A(G138), .B(new_n476), .C1(new_n460), .C2(new_n461), .ZN(new_n493));
  INV_X1    g068(.A(KEYINPUT4), .ZN(new_n494));
  NAND2_X1  g069(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  NAND3_X1  g070(.A1(new_n487), .A2(new_n492), .A3(new_n495), .ZN(new_n496));
  INV_X1    g071(.A(new_n496), .ZN(G164));
  INV_X1    g072(.A(KEYINPUT5), .ZN(new_n498));
  INV_X1    g073(.A(G543), .ZN(new_n499));
  OAI21_X1  g074(.A(new_n498), .B1(new_n499), .B2(KEYINPUT67), .ZN(new_n500));
  INV_X1    g075(.A(KEYINPUT67), .ZN(new_n501));
  NAND3_X1  g076(.A1(new_n501), .A2(KEYINPUT5), .A3(G543), .ZN(new_n502));
  NAND2_X1  g077(.A1(new_n500), .A2(new_n502), .ZN(new_n503));
  XNOR2_X1  g078(.A(KEYINPUT6), .B(G651), .ZN(new_n504));
  NAND2_X1  g079(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  XOR2_X1   g080(.A(KEYINPUT68), .B(G88), .Z(new_n506));
  NAND2_X1  g081(.A1(new_n504), .A2(G543), .ZN(new_n507));
  INV_X1    g082(.A(G50), .ZN(new_n508));
  OAI22_X1  g083(.A1(new_n505), .A2(new_n506), .B1(new_n507), .B2(new_n508), .ZN(new_n509));
  XNOR2_X1  g084(.A(new_n509), .B(KEYINPUT69), .ZN(new_n510));
  INV_X1    g085(.A(G651), .ZN(new_n511));
  AND2_X1   g086(.A1(new_n503), .A2(G62), .ZN(new_n512));
  OR2_X1    g087(.A1(new_n512), .A2(KEYINPUT70), .ZN(new_n513));
  AOI22_X1  g088(.A1(new_n512), .A2(KEYINPUT70), .B1(G75), .B2(G543), .ZN(new_n514));
  AOI21_X1  g089(.A(new_n511), .B1(new_n513), .B2(new_n514), .ZN(new_n515));
  NOR2_X1   g090(.A1(new_n510), .A2(new_n515), .ZN(G166));
  XNOR2_X1  g091(.A(new_n503), .B(KEYINPUT71), .ZN(new_n517));
  INV_X1    g092(.A(new_n517), .ZN(new_n518));
  NAND3_X1  g093(.A1(new_n518), .A2(G63), .A3(G651), .ZN(new_n519));
  INV_X1    g094(.A(new_n505), .ZN(new_n520));
  NAND2_X1  g095(.A1(new_n520), .A2(G89), .ZN(new_n521));
  NAND3_X1  g096(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n522));
  XOR2_X1   g097(.A(new_n522), .B(KEYINPUT7), .Z(new_n523));
  INV_X1    g098(.A(new_n507), .ZN(new_n524));
  AOI21_X1  g099(.A(new_n523), .B1(G51), .B2(new_n524), .ZN(new_n525));
  NAND3_X1  g100(.A1(new_n519), .A2(new_n521), .A3(new_n525), .ZN(G286));
  INV_X1    g101(.A(G286), .ZN(G168));
  INV_X1    g102(.A(G90), .ZN(new_n528));
  INV_X1    g103(.A(G52), .ZN(new_n529));
  OAI22_X1  g104(.A1(new_n505), .A2(new_n528), .B1(new_n507), .B2(new_n529), .ZN(new_n530));
  NAND2_X1  g105(.A1(G77), .A2(G543), .ZN(new_n531));
  INV_X1    g106(.A(G64), .ZN(new_n532));
  OAI21_X1  g107(.A(new_n531), .B1(new_n517), .B2(new_n532), .ZN(new_n533));
  AOI21_X1  g108(.A(new_n530), .B1(new_n533), .B2(G651), .ZN(G171));
  NAND2_X1  g109(.A1(G68), .A2(G543), .ZN(new_n535));
  INV_X1    g110(.A(G56), .ZN(new_n536));
  OAI21_X1  g111(.A(new_n535), .B1(new_n517), .B2(new_n536), .ZN(new_n537));
  INV_X1    g112(.A(KEYINPUT72), .ZN(new_n538));
  AOI21_X1  g113(.A(new_n511), .B1(new_n537), .B2(new_n538), .ZN(new_n539));
  OAI21_X1  g114(.A(new_n539), .B1(new_n538), .B2(new_n537), .ZN(new_n540));
  AOI22_X1  g115(.A1(new_n520), .A2(G81), .B1(new_n524), .B2(G43), .ZN(new_n541));
  NAND2_X1  g116(.A1(new_n540), .A2(new_n541), .ZN(new_n542));
  INV_X1    g117(.A(new_n542), .ZN(new_n543));
  NAND2_X1  g118(.A1(new_n543), .A2(G860), .ZN(G153));
  AND3_X1   g119(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n545));
  NAND2_X1  g120(.A1(new_n545), .A2(G36), .ZN(new_n546));
  XOR2_X1   g121(.A(new_n546), .B(KEYINPUT73), .Z(G176));
  NAND2_X1  g122(.A1(G1), .A2(G3), .ZN(new_n548));
  XNOR2_X1  g123(.A(new_n548), .B(KEYINPUT8), .ZN(new_n549));
  NAND2_X1  g124(.A1(new_n545), .A2(new_n549), .ZN(G188));
  INV_X1    g125(.A(KEYINPUT74), .ZN(new_n551));
  NAND4_X1  g126(.A1(new_n524), .A2(new_n551), .A3(KEYINPUT9), .A4(G53), .ZN(new_n552));
  NAND2_X1  g127(.A1(new_n520), .A2(G91), .ZN(new_n553));
  XNOR2_X1  g128(.A(KEYINPUT74), .B(KEYINPUT9), .ZN(new_n554));
  INV_X1    g129(.A(G53), .ZN(new_n555));
  OAI21_X1  g130(.A(new_n554), .B1(new_n507), .B2(new_n555), .ZN(new_n556));
  NAND3_X1  g131(.A1(new_n552), .A2(new_n553), .A3(new_n556), .ZN(new_n557));
  INV_X1    g132(.A(G65), .ZN(new_n558));
  AND2_X1   g133(.A1(new_n558), .A2(KEYINPUT75), .ZN(new_n559));
  NOR2_X1   g134(.A1(new_n558), .A2(KEYINPUT75), .ZN(new_n560));
  OAI21_X1  g135(.A(new_n503), .B1(new_n559), .B2(new_n560), .ZN(new_n561));
  NAND2_X1  g136(.A1(G78), .A2(G543), .ZN(new_n562));
  AOI21_X1  g137(.A(new_n511), .B1(new_n561), .B2(new_n562), .ZN(new_n563));
  NOR2_X1   g138(.A1(new_n557), .A2(new_n563), .ZN(new_n564));
  INV_X1    g139(.A(new_n564), .ZN(G299));
  INV_X1    g140(.A(G171), .ZN(G301));
  INV_X1    g141(.A(G166), .ZN(G303));
  OAI21_X1  g142(.A(G651), .B1(new_n518), .B2(G74), .ZN(new_n568));
  AOI22_X1  g143(.A1(new_n520), .A2(G87), .B1(new_n524), .B2(G49), .ZN(new_n569));
  NAND2_X1  g144(.A1(new_n568), .A2(new_n569), .ZN(G288));
  AOI22_X1  g145(.A1(new_n503), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n571));
  OR2_X1    g146(.A1(new_n571), .A2(new_n511), .ZN(new_n572));
  NAND2_X1  g147(.A1(new_n520), .A2(G86), .ZN(new_n573));
  NAND2_X1  g148(.A1(new_n524), .A2(G48), .ZN(new_n574));
  NAND3_X1  g149(.A1(new_n572), .A2(new_n573), .A3(new_n574), .ZN(G305));
  AND2_X1   g150(.A1(new_n518), .A2(G60), .ZN(new_n576));
  AND2_X1   g151(.A1(G72), .A2(G543), .ZN(new_n577));
  OAI21_X1  g152(.A(G651), .B1(new_n576), .B2(new_n577), .ZN(new_n578));
  XNOR2_X1  g153(.A(KEYINPUT76), .B(G47), .ZN(new_n579));
  AOI22_X1  g154(.A1(new_n520), .A2(G85), .B1(new_n524), .B2(new_n579), .ZN(new_n580));
  NAND2_X1  g155(.A1(new_n578), .A2(new_n580), .ZN(G290));
  INV_X1    g156(.A(G868), .ZN(new_n582));
  NOR2_X1   g157(.A1(G301), .A2(new_n582), .ZN(new_n583));
  NAND2_X1  g158(.A1(new_n520), .A2(G92), .ZN(new_n584));
  XNOR2_X1  g159(.A(new_n584), .B(KEYINPUT10), .ZN(new_n585));
  AOI21_X1  g160(.A(new_n585), .B1(G54), .B2(new_n524), .ZN(new_n586));
  AOI22_X1  g161(.A1(new_n503), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n587));
  AOI21_X1  g162(.A(new_n511), .B1(new_n587), .B2(KEYINPUT77), .ZN(new_n588));
  OAI21_X1  g163(.A(new_n588), .B1(KEYINPUT77), .B2(new_n587), .ZN(new_n589));
  NAND2_X1  g164(.A1(new_n586), .A2(new_n589), .ZN(new_n590));
  INV_X1    g165(.A(new_n590), .ZN(new_n591));
  AOI21_X1  g166(.A(new_n583), .B1(new_n591), .B2(new_n582), .ZN(G284));
  AOI21_X1  g167(.A(new_n583), .B1(new_n591), .B2(new_n582), .ZN(G321));
  MUX2_X1   g168(.A(G286), .B(G299), .S(new_n582), .Z(G297));
  XNOR2_X1  g169(.A(G297), .B(KEYINPUT78), .ZN(G280));
  INV_X1    g170(.A(G559), .ZN(new_n596));
  OAI21_X1  g171(.A(new_n591), .B1(new_n596), .B2(G860), .ZN(G148));
  NOR2_X1   g172(.A1(new_n542), .A2(G868), .ZN(new_n598));
  NOR2_X1   g173(.A1(new_n590), .A2(G559), .ZN(new_n599));
  AOI21_X1  g174(.A(new_n598), .B1(new_n599), .B2(G868), .ZN(new_n600));
  XNOR2_X1  g175(.A(new_n600), .B(KEYINPUT79), .ZN(G323));
  XOR2_X1   g176(.A(KEYINPUT80), .B(KEYINPUT11), .Z(new_n602));
  XNOR2_X1  g177(.A(G323), .B(new_n602), .ZN(G282));
  NAND2_X1  g178(.A1(new_n469), .A2(G2104), .ZN(new_n604));
  XOR2_X1   g179(.A(new_n604), .B(KEYINPUT12), .Z(new_n605));
  INV_X1    g180(.A(new_n605), .ZN(new_n606));
  INV_X1    g181(.A(G2100), .ZN(new_n607));
  AOI22_X1  g182(.A1(new_n606), .A2(KEYINPUT13), .B1(KEYINPUT81), .B2(new_n607), .ZN(new_n608));
  OAI21_X1  g183(.A(new_n608), .B1(KEYINPUT13), .B2(new_n606), .ZN(new_n609));
  OR3_X1    g184(.A1(new_n609), .A2(KEYINPUT81), .A3(new_n607), .ZN(new_n610));
  OAI21_X1  g185(.A(new_n609), .B1(KEYINPUT81), .B2(new_n607), .ZN(new_n611));
  MUX2_X1   g186(.A(G99), .B(G111), .S(G2105), .Z(new_n612));
  AOI22_X1  g187(.A1(new_n477), .A2(G123), .B1(G2104), .B2(new_n612), .ZN(new_n613));
  INV_X1    g188(.A(new_n474), .ZN(new_n614));
  INV_X1    g189(.A(G135), .ZN(new_n615));
  OAI21_X1  g190(.A(new_n613), .B1(new_n614), .B2(new_n615), .ZN(new_n616));
  XOR2_X1   g191(.A(new_n616), .B(G2096), .Z(new_n617));
  NAND3_X1  g192(.A1(new_n610), .A2(new_n611), .A3(new_n617), .ZN(G156));
  XNOR2_X1  g193(.A(KEYINPUT15), .B(G2435), .ZN(new_n619));
  XNOR2_X1  g194(.A(new_n619), .B(G2438), .ZN(new_n620));
  XNOR2_X1  g195(.A(G2427), .B(G2430), .ZN(new_n621));
  NAND2_X1  g196(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  AND3_X1   g197(.A1(new_n622), .A2(KEYINPUT83), .A3(KEYINPUT14), .ZN(new_n623));
  AOI21_X1  g198(.A(KEYINPUT83), .B1(new_n622), .B2(KEYINPUT14), .ZN(new_n624));
  OAI22_X1  g199(.A1(new_n623), .A2(new_n624), .B1(new_n620), .B2(new_n621), .ZN(new_n625));
  XOR2_X1   g200(.A(KEYINPUT82), .B(KEYINPUT16), .Z(new_n626));
  XNOR2_X1  g201(.A(new_n625), .B(new_n626), .ZN(new_n627));
  XOR2_X1   g202(.A(G1341), .B(G1348), .Z(new_n628));
  XNOR2_X1  g203(.A(new_n627), .B(new_n628), .ZN(new_n629));
  XNOR2_X1  g204(.A(G2451), .B(G2454), .ZN(new_n630));
  XNOR2_X1  g205(.A(G2443), .B(G2446), .ZN(new_n631));
  XOR2_X1   g206(.A(new_n630), .B(new_n631), .Z(new_n632));
  INV_X1    g207(.A(new_n632), .ZN(new_n633));
  OR2_X1    g208(.A1(new_n629), .A2(new_n633), .ZN(new_n634));
  INV_X1    g209(.A(G14), .ZN(new_n635));
  AOI21_X1  g210(.A(new_n635), .B1(new_n629), .B2(new_n633), .ZN(new_n636));
  AND2_X1   g211(.A1(new_n634), .A2(new_n636), .ZN(G401));
  XNOR2_X1  g212(.A(G2067), .B(G2678), .ZN(new_n638));
  XNOR2_X1  g213(.A(new_n638), .B(KEYINPUT84), .ZN(new_n639));
  XNOR2_X1  g214(.A(G2072), .B(G2078), .ZN(new_n640));
  XOR2_X1   g215(.A(G2084), .B(G2090), .Z(new_n641));
  NAND3_X1  g216(.A1(new_n639), .A2(new_n640), .A3(new_n641), .ZN(new_n642));
  INV_X1    g217(.A(KEYINPUT18), .ZN(new_n643));
  XNOR2_X1  g218(.A(new_n642), .B(new_n643), .ZN(new_n644));
  OR2_X1    g219(.A1(new_n639), .A2(new_n641), .ZN(new_n645));
  AOI21_X1  g220(.A(new_n640), .B1(new_n645), .B2(KEYINPUT17), .ZN(new_n646));
  INV_X1    g221(.A(new_n641), .ZN(new_n647));
  NAND2_X1  g222(.A1(new_n640), .A2(KEYINPUT17), .ZN(new_n648));
  NAND2_X1  g223(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  NAND2_X1  g224(.A1(new_n639), .A2(new_n649), .ZN(new_n650));
  OAI21_X1  g225(.A(new_n650), .B1(new_n647), .B2(new_n648), .ZN(new_n651));
  OAI21_X1  g226(.A(new_n644), .B1(new_n646), .B2(new_n651), .ZN(new_n652));
  XNOR2_X1  g227(.A(new_n652), .B(G2096), .ZN(new_n653));
  XNOR2_X1  g228(.A(KEYINPUT85), .B(G2100), .ZN(new_n654));
  XNOR2_X1  g229(.A(new_n653), .B(new_n654), .ZN(G227));
  XOR2_X1   g230(.A(G1971), .B(G1976), .Z(new_n656));
  XNOR2_X1  g231(.A(new_n656), .B(KEYINPUT19), .ZN(new_n657));
  XNOR2_X1  g232(.A(G1956), .B(G2474), .ZN(new_n658));
  XNOR2_X1  g233(.A(G1961), .B(G1966), .ZN(new_n659));
  NOR2_X1   g234(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  AND2_X1   g235(.A1(new_n658), .A2(new_n659), .ZN(new_n661));
  NOR3_X1   g236(.A1(new_n657), .A2(new_n660), .A3(new_n661), .ZN(new_n662));
  NAND2_X1  g237(.A1(new_n657), .A2(new_n660), .ZN(new_n663));
  XOR2_X1   g238(.A(new_n663), .B(KEYINPUT20), .Z(new_n664));
  AOI211_X1 g239(.A(new_n662), .B(new_n664), .C1(new_n657), .C2(new_n661), .ZN(new_n665));
  XOR2_X1   g240(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n666));
  XOR2_X1   g241(.A(new_n665), .B(new_n666), .Z(new_n667));
  XNOR2_X1  g242(.A(G1991), .B(G1996), .ZN(new_n668));
  XNOR2_X1  g243(.A(G1981), .B(G1986), .ZN(new_n669));
  XNOR2_X1  g244(.A(new_n668), .B(new_n669), .ZN(new_n670));
  XNOR2_X1  g245(.A(new_n667), .B(new_n670), .ZN(new_n671));
  INV_X1    g246(.A(new_n671), .ZN(G229));
  NOR2_X1   g247(.A1(G25), .A2(G29), .ZN(new_n673));
  NAND2_X1  g248(.A1(new_n474), .A2(G131), .ZN(new_n674));
  MUX2_X1   g249(.A(G95), .B(G107), .S(G2105), .Z(new_n675));
  AOI22_X1  g250(.A1(new_n477), .A2(G119), .B1(G2104), .B2(new_n675), .ZN(new_n676));
  NAND2_X1  g251(.A1(new_n674), .A2(new_n676), .ZN(new_n677));
  INV_X1    g252(.A(new_n677), .ZN(new_n678));
  AOI21_X1  g253(.A(new_n673), .B1(new_n678), .B2(G29), .ZN(new_n679));
  XOR2_X1   g254(.A(KEYINPUT35), .B(G1991), .Z(new_n680));
  XNOR2_X1  g255(.A(new_n679), .B(new_n680), .ZN(new_n681));
  MUX2_X1   g256(.A(G24), .B(G290), .S(G16), .Z(new_n682));
  OAI21_X1  g257(.A(new_n681), .B1(G1986), .B2(new_n682), .ZN(new_n683));
  AOI21_X1  g258(.A(new_n683), .B1(G1986), .B2(new_n682), .ZN(new_n684));
  NOR2_X1   g259(.A1(G16), .A2(G23), .ZN(new_n685));
  XNOR2_X1  g260(.A(new_n685), .B(KEYINPUT86), .ZN(new_n686));
  INV_X1    g261(.A(G16), .ZN(new_n687));
  OAI21_X1  g262(.A(new_n686), .B1(G288), .B2(new_n687), .ZN(new_n688));
  XNOR2_X1  g263(.A(KEYINPUT33), .B(G1976), .ZN(new_n689));
  XNOR2_X1  g264(.A(new_n688), .B(new_n689), .ZN(new_n690));
  NAND2_X1  g265(.A1(G166), .A2(G16), .ZN(new_n691));
  OAI21_X1  g266(.A(new_n691), .B1(G16), .B2(G22), .ZN(new_n692));
  INV_X1    g267(.A(G1971), .ZN(new_n693));
  AOI21_X1  g268(.A(new_n690), .B1(new_n692), .B2(new_n693), .ZN(new_n694));
  NOR2_X1   g269(.A1(G6), .A2(G16), .ZN(new_n695));
  INV_X1    g270(.A(G305), .ZN(new_n696));
  AOI21_X1  g271(.A(new_n695), .B1(new_n696), .B2(G16), .ZN(new_n697));
  XOR2_X1   g272(.A(KEYINPUT32), .B(G1981), .Z(new_n698));
  XNOR2_X1  g273(.A(new_n697), .B(new_n698), .ZN(new_n699));
  OAI211_X1 g274(.A(new_n694), .B(new_n699), .C1(new_n693), .C2(new_n692), .ZN(new_n700));
  OAI21_X1  g275(.A(new_n684), .B1(new_n700), .B2(KEYINPUT34), .ZN(new_n701));
  AOI21_X1  g276(.A(new_n701), .B1(KEYINPUT34), .B2(new_n700), .ZN(new_n702));
  XOR2_X1   g277(.A(new_n702), .B(KEYINPUT36), .Z(new_n703));
  NAND2_X1  g278(.A1(new_n687), .A2(G20), .ZN(new_n704));
  XNOR2_X1  g279(.A(new_n704), .B(KEYINPUT23), .ZN(new_n705));
  OAI21_X1  g280(.A(new_n705), .B1(new_n564), .B2(new_n687), .ZN(new_n706));
  XNOR2_X1  g281(.A(new_n706), .B(G1956), .ZN(new_n707));
  NAND2_X1  g282(.A1(new_n687), .A2(G21), .ZN(new_n708));
  OAI21_X1  g283(.A(new_n708), .B1(G168), .B2(new_n687), .ZN(new_n709));
  INV_X1    g284(.A(G1966), .ZN(new_n710));
  XNOR2_X1  g285(.A(new_n709), .B(new_n710), .ZN(new_n711));
  INV_X1    g286(.A(G29), .ZN(new_n712));
  OR3_X1    g287(.A1(new_n616), .A2(KEYINPUT92), .A3(new_n712), .ZN(new_n713));
  OAI21_X1  g288(.A(KEYINPUT92), .B1(new_n616), .B2(new_n712), .ZN(new_n714));
  NAND2_X1  g289(.A1(G164), .A2(G29), .ZN(new_n715));
  OAI21_X1  g290(.A(new_n715), .B1(G27), .B2(G29), .ZN(new_n716));
  INV_X1    g291(.A(G2078), .ZN(new_n717));
  AOI22_X1  g292(.A1(new_n713), .A2(new_n714), .B1(new_n716), .B2(new_n717), .ZN(new_n718));
  NOR2_X1   g293(.A1(G29), .A2(G35), .ZN(new_n719));
  AOI21_X1  g294(.A(new_n719), .B1(G162), .B2(G29), .ZN(new_n720));
  XOR2_X1   g295(.A(new_n720), .B(KEYINPUT29), .Z(new_n721));
  INV_X1    g296(.A(G2090), .ZN(new_n722));
  OAI211_X1 g297(.A(new_n711), .B(new_n718), .C1(new_n721), .C2(new_n722), .ZN(new_n723));
  AOI211_X1 g298(.A(new_n707), .B(new_n723), .C1(new_n722), .C2(new_n721), .ZN(new_n724));
  NAND2_X1  g299(.A1(new_n474), .A2(G141), .ZN(new_n725));
  AND2_X1   g300(.A1(new_n471), .A2(G105), .ZN(new_n726));
  NAND3_X1  g301(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n727));
  XNOR2_X1  g302(.A(new_n727), .B(KEYINPUT26), .ZN(new_n728));
  AOI211_X1 g303(.A(new_n726), .B(new_n728), .C1(G129), .C2(new_n477), .ZN(new_n729));
  NAND2_X1  g304(.A1(new_n725), .A2(new_n729), .ZN(new_n730));
  INV_X1    g305(.A(new_n730), .ZN(new_n731));
  NAND2_X1  g306(.A1(new_n731), .A2(G29), .ZN(new_n732));
  NOR2_X1   g307(.A1(G29), .A2(G32), .ZN(new_n733));
  OAI21_X1  g308(.A(new_n732), .B1(KEYINPUT91), .B2(new_n733), .ZN(new_n734));
  OAI21_X1  g309(.A(new_n734), .B1(KEYINPUT91), .B2(new_n732), .ZN(new_n735));
  XNOR2_X1  g310(.A(KEYINPUT27), .B(G1996), .ZN(new_n736));
  OR2_X1    g311(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  NAND2_X1  g312(.A1(new_n735), .A2(new_n736), .ZN(new_n738));
  OR2_X1    g313(.A1(KEYINPUT24), .A2(G34), .ZN(new_n739));
  NAND2_X1  g314(.A1(KEYINPUT24), .A2(G34), .ZN(new_n740));
  AOI21_X1  g315(.A(G29), .B1(new_n739), .B2(new_n740), .ZN(new_n741));
  AOI21_X1  g316(.A(new_n741), .B1(G160), .B2(G29), .ZN(new_n742));
  NAND2_X1  g317(.A1(new_n742), .A2(G2084), .ZN(new_n743));
  NAND3_X1  g318(.A1(new_n737), .A2(new_n738), .A3(new_n743), .ZN(new_n744));
  NOR2_X1   g319(.A1(G29), .A2(G33), .ZN(new_n745));
  XNOR2_X1  g320(.A(new_n745), .B(KEYINPUT89), .ZN(new_n746));
  NAND2_X1  g321(.A1(new_n474), .A2(G139), .ZN(new_n747));
  XOR2_X1   g322(.A(KEYINPUT90), .B(KEYINPUT25), .Z(new_n748));
  NAND2_X1  g323(.A1(new_n471), .A2(G103), .ZN(new_n749));
  XNOR2_X1  g324(.A(new_n748), .B(new_n749), .ZN(new_n750));
  AOI22_X1  g325(.A1(new_n465), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n751));
  OAI211_X1 g326(.A(new_n747), .B(new_n750), .C1(new_n476), .C2(new_n751), .ZN(new_n752));
  OAI21_X1  g327(.A(new_n746), .B1(new_n752), .B2(new_n712), .ZN(new_n753));
  XNOR2_X1  g328(.A(new_n753), .B(G2072), .ZN(new_n754));
  XOR2_X1   g329(.A(KEYINPUT31), .B(G11), .Z(new_n755));
  XNOR2_X1  g330(.A(KEYINPUT30), .B(G28), .ZN(new_n756));
  AOI21_X1  g331(.A(new_n755), .B1(new_n712), .B2(new_n756), .ZN(new_n757));
  OAI211_X1 g332(.A(new_n754), .B(new_n757), .C1(new_n717), .C2(new_n716), .ZN(new_n758));
  NAND2_X1  g333(.A1(new_n712), .A2(G26), .ZN(new_n759));
  XOR2_X1   g334(.A(new_n759), .B(KEYINPUT28), .Z(new_n760));
  NAND2_X1  g335(.A1(new_n474), .A2(G140), .ZN(new_n761));
  NOR2_X1   g336(.A1(G104), .A2(G2105), .ZN(new_n762));
  XNOR2_X1  g337(.A(new_n762), .B(KEYINPUT88), .ZN(new_n763));
  INV_X1    g338(.A(G116), .ZN(new_n764));
  AOI21_X1  g339(.A(new_n470), .B1(new_n764), .B2(G2105), .ZN(new_n765));
  AOI22_X1  g340(.A1(G128), .A2(new_n477), .B1(new_n763), .B2(new_n765), .ZN(new_n766));
  NAND2_X1  g341(.A1(new_n761), .A2(new_n766), .ZN(new_n767));
  AOI21_X1  g342(.A(new_n760), .B1(new_n767), .B2(G29), .ZN(new_n768));
  XNOR2_X1  g343(.A(new_n768), .B(G2067), .ZN(new_n769));
  OAI21_X1  g344(.A(new_n769), .B1(G2084), .B2(new_n742), .ZN(new_n770));
  NOR3_X1   g345(.A1(new_n744), .A2(new_n758), .A3(new_n770), .ZN(new_n771));
  NAND2_X1  g346(.A1(new_n724), .A2(new_n771), .ZN(new_n772));
  NOR2_X1   g347(.A1(G16), .A2(G19), .ZN(new_n773));
  AOI21_X1  g348(.A(new_n773), .B1(new_n543), .B2(G16), .ZN(new_n774));
  XNOR2_X1  g349(.A(KEYINPUT87), .B(G1341), .ZN(new_n775));
  XNOR2_X1  g350(.A(new_n774), .B(new_n775), .ZN(new_n776));
  NOR2_X1   g351(.A1(G4), .A2(G16), .ZN(new_n777));
  AOI21_X1  g352(.A(new_n777), .B1(new_n591), .B2(G16), .ZN(new_n778));
  INV_X1    g353(.A(G1348), .ZN(new_n779));
  XNOR2_X1  g354(.A(new_n778), .B(new_n779), .ZN(new_n780));
  NAND2_X1  g355(.A1(new_n687), .A2(G5), .ZN(new_n781));
  OAI21_X1  g356(.A(new_n781), .B1(G171), .B2(new_n687), .ZN(new_n782));
  NAND2_X1  g357(.A1(new_n782), .A2(G1961), .ZN(new_n783));
  XOR2_X1   g358(.A(new_n783), .B(KEYINPUT93), .Z(new_n784));
  OAI211_X1 g359(.A(new_n780), .B(new_n784), .C1(G1961), .C2(new_n782), .ZN(new_n785));
  NOR3_X1   g360(.A1(new_n772), .A2(new_n776), .A3(new_n785), .ZN(new_n786));
  NAND2_X1  g361(.A1(new_n703), .A2(new_n786), .ZN(G150));
  INV_X1    g362(.A(G150), .ZN(G311));
  AOI22_X1  g363(.A1(new_n520), .A2(G93), .B1(new_n524), .B2(G55), .ZN(new_n789));
  XNOR2_X1  g364(.A(new_n789), .B(KEYINPUT94), .ZN(new_n790));
  NAND2_X1  g365(.A1(G80), .A2(G543), .ZN(new_n791));
  INV_X1    g366(.A(G67), .ZN(new_n792));
  OAI21_X1  g367(.A(new_n791), .B1(new_n517), .B2(new_n792), .ZN(new_n793));
  AOI21_X1  g368(.A(new_n790), .B1(G651), .B2(new_n793), .ZN(new_n794));
  INV_X1    g369(.A(G860), .ZN(new_n795));
  NOR2_X1   g370(.A1(new_n794), .A2(new_n795), .ZN(new_n796));
  XNOR2_X1  g371(.A(new_n796), .B(KEYINPUT37), .ZN(new_n797));
  XNOR2_X1  g372(.A(new_n542), .B(new_n794), .ZN(new_n798));
  XNOR2_X1  g373(.A(new_n798), .B(KEYINPUT38), .ZN(new_n799));
  NOR2_X1   g374(.A1(new_n590), .A2(new_n596), .ZN(new_n800));
  XNOR2_X1  g375(.A(new_n799), .B(new_n800), .ZN(new_n801));
  INV_X1    g376(.A(new_n801), .ZN(new_n802));
  AND2_X1   g377(.A1(new_n802), .A2(KEYINPUT39), .ZN(new_n803));
  OAI21_X1  g378(.A(new_n795), .B1(new_n802), .B2(KEYINPUT39), .ZN(new_n804));
  OAI21_X1  g379(.A(new_n797), .B1(new_n803), .B2(new_n804), .ZN(G145));
  XNOR2_X1  g380(.A(new_n677), .B(new_n605), .ZN(new_n806));
  MUX2_X1   g381(.A(G106), .B(G118), .S(G2105), .Z(new_n807));
  AOI22_X1  g382(.A1(new_n477), .A2(G130), .B1(G2104), .B2(new_n807), .ZN(new_n808));
  INV_X1    g383(.A(G142), .ZN(new_n809));
  OAI21_X1  g384(.A(new_n808), .B1(new_n614), .B2(new_n809), .ZN(new_n810));
  XNOR2_X1  g385(.A(new_n806), .B(new_n810), .ZN(new_n811));
  XNOR2_X1  g386(.A(new_n767), .B(G164), .ZN(new_n812));
  XNOR2_X1  g387(.A(new_n811), .B(new_n812), .ZN(new_n813));
  XNOR2_X1  g388(.A(new_n752), .B(new_n730), .ZN(new_n814));
  XNOR2_X1  g389(.A(new_n813), .B(new_n814), .ZN(new_n815));
  XNOR2_X1  g390(.A(new_n480), .B(G160), .ZN(new_n816));
  XOR2_X1   g391(.A(new_n816), .B(new_n616), .Z(new_n817));
  OR2_X1    g392(.A1(new_n815), .A2(new_n817), .ZN(new_n818));
  NAND2_X1  g393(.A1(new_n815), .A2(new_n817), .ZN(new_n819));
  XOR2_X1   g394(.A(KEYINPUT95), .B(G37), .Z(new_n820));
  NAND3_X1  g395(.A1(new_n818), .A2(new_n819), .A3(new_n820), .ZN(new_n821));
  XNOR2_X1  g396(.A(new_n821), .B(KEYINPUT40), .ZN(G395));
  XNOR2_X1  g397(.A(new_n798), .B(new_n599), .ZN(new_n823));
  OAI21_X1  g398(.A(KEYINPUT96), .B1(new_n590), .B2(new_n564), .ZN(new_n824));
  INV_X1    g399(.A(KEYINPUT96), .ZN(new_n825));
  NAND4_X1  g400(.A1(new_n586), .A2(G299), .A3(new_n825), .A4(new_n589), .ZN(new_n826));
  NAND2_X1  g401(.A1(new_n824), .A2(new_n826), .ZN(new_n827));
  NAND2_X1  g402(.A1(new_n590), .A2(new_n564), .ZN(new_n828));
  NAND3_X1  g403(.A1(new_n823), .A2(new_n827), .A3(new_n828), .ZN(new_n829));
  NAND2_X1  g404(.A1(new_n827), .A2(new_n828), .ZN(new_n830));
  INV_X1    g405(.A(KEYINPUT41), .ZN(new_n831));
  NAND2_X1  g406(.A1(new_n830), .A2(new_n831), .ZN(new_n832));
  NAND3_X1  g407(.A1(new_n827), .A2(KEYINPUT41), .A3(new_n828), .ZN(new_n833));
  NAND2_X1  g408(.A1(new_n832), .A2(new_n833), .ZN(new_n834));
  OAI21_X1  g409(.A(new_n829), .B1(new_n823), .B2(new_n834), .ZN(new_n835));
  XNOR2_X1  g410(.A(G166), .B(KEYINPUT97), .ZN(new_n836));
  XNOR2_X1  g411(.A(new_n836), .B(new_n696), .ZN(new_n837));
  INV_X1    g412(.A(KEYINPUT98), .ZN(new_n838));
  XOR2_X1   g413(.A(G290), .B(G288), .Z(new_n839));
  AND3_X1   g414(.A1(new_n837), .A2(new_n838), .A3(new_n839), .ZN(new_n840));
  AOI21_X1  g415(.A(new_n838), .B1(new_n837), .B2(new_n839), .ZN(new_n841));
  OAI22_X1  g416(.A1(new_n840), .A2(new_n841), .B1(new_n837), .B2(new_n839), .ZN(new_n842));
  INV_X1    g417(.A(KEYINPUT42), .ZN(new_n843));
  OR2_X1    g418(.A1(new_n842), .A2(new_n843), .ZN(new_n844));
  NAND2_X1  g419(.A1(new_n842), .A2(new_n843), .ZN(new_n845));
  AOI21_X1  g420(.A(new_n835), .B1(new_n844), .B2(new_n845), .ZN(new_n846));
  INV_X1    g421(.A(KEYINPUT99), .ZN(new_n847));
  AND2_X1   g422(.A1(new_n846), .A2(new_n847), .ZN(new_n848));
  NAND3_X1  g423(.A1(new_n844), .A2(new_n835), .A3(new_n845), .ZN(new_n849));
  OAI21_X1  g424(.A(new_n849), .B1(new_n846), .B2(new_n847), .ZN(new_n850));
  OAI21_X1  g425(.A(G868), .B1(new_n848), .B2(new_n850), .ZN(new_n851));
  OAI21_X1  g426(.A(new_n851), .B1(G868), .B2(new_n794), .ZN(G295));
  OAI21_X1  g427(.A(new_n851), .B1(G868), .B2(new_n794), .ZN(G331));
  INV_X1    g428(.A(KEYINPUT44), .ZN(new_n854));
  AOI21_X1  g429(.A(G286), .B1(G171), .B2(KEYINPUT100), .ZN(new_n855));
  OAI21_X1  g430(.A(new_n855), .B1(KEYINPUT100), .B2(G171), .ZN(new_n856));
  OR3_X1    g431(.A1(G168), .A2(KEYINPUT100), .A3(G171), .ZN(new_n857));
  AND2_X1   g432(.A1(new_n856), .A2(new_n857), .ZN(new_n858));
  OR2_X1    g433(.A1(new_n858), .A2(new_n798), .ZN(new_n859));
  NAND2_X1  g434(.A1(new_n858), .A2(new_n798), .ZN(new_n860));
  NAND3_X1  g435(.A1(new_n859), .A2(new_n830), .A3(new_n860), .ZN(new_n861));
  NAND2_X1  g436(.A1(new_n859), .A2(new_n860), .ZN(new_n862));
  AND3_X1   g437(.A1(new_n834), .A2(new_n862), .A3(KEYINPUT101), .ZN(new_n863));
  AOI21_X1  g438(.A(KEYINPUT101), .B1(new_n834), .B2(new_n862), .ZN(new_n864));
  OAI211_X1 g439(.A(new_n842), .B(new_n861), .C1(new_n863), .C2(new_n864), .ZN(new_n865));
  INV_X1    g440(.A(new_n865), .ZN(new_n866));
  NAND2_X1  g441(.A1(new_n861), .A2(KEYINPUT104), .ZN(new_n867));
  INV_X1    g442(.A(KEYINPUT104), .ZN(new_n868));
  NAND4_X1  g443(.A1(new_n859), .A2(new_n868), .A3(new_n830), .A4(new_n860), .ZN(new_n869));
  AOI21_X1  g444(.A(KEYINPUT41), .B1(new_n827), .B2(new_n828), .ZN(new_n870));
  AOI22_X1  g445(.A1(new_n859), .A2(new_n860), .B1(new_n870), .B2(KEYINPUT103), .ZN(new_n871));
  INV_X1    g446(.A(KEYINPUT103), .ZN(new_n872));
  NAND3_X1  g447(.A1(new_n832), .A2(new_n872), .A3(new_n833), .ZN(new_n873));
  AOI22_X1  g448(.A1(new_n867), .A2(new_n869), .B1(new_n871), .B2(new_n873), .ZN(new_n874));
  OAI21_X1  g449(.A(new_n820), .B1(new_n874), .B2(new_n842), .ZN(new_n875));
  OAI21_X1  g450(.A(KEYINPUT43), .B1(new_n866), .B2(new_n875), .ZN(new_n876));
  OAI21_X1  g451(.A(new_n861), .B1(new_n863), .B2(new_n864), .ZN(new_n877));
  INV_X1    g452(.A(KEYINPUT102), .ZN(new_n878));
  NOR2_X1   g453(.A1(new_n842), .A2(new_n878), .ZN(new_n879));
  NAND2_X1  g454(.A1(new_n877), .A2(new_n879), .ZN(new_n880));
  OAI221_X1 g455(.A(new_n861), .B1(new_n842), .B2(new_n878), .C1(new_n863), .C2(new_n864), .ZN(new_n881));
  INV_X1    g456(.A(KEYINPUT43), .ZN(new_n882));
  INV_X1    g457(.A(G37), .ZN(new_n883));
  NAND4_X1  g458(.A1(new_n880), .A2(new_n881), .A3(new_n882), .A4(new_n883), .ZN(new_n884));
  AOI21_X1  g459(.A(new_n854), .B1(new_n876), .B2(new_n884), .ZN(new_n885));
  OAI21_X1  g460(.A(new_n882), .B1(new_n866), .B2(new_n875), .ZN(new_n886));
  NAND4_X1  g461(.A1(new_n880), .A2(new_n881), .A3(KEYINPUT43), .A4(new_n883), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n886), .A2(new_n887), .ZN(new_n888));
  AOI21_X1  g463(.A(new_n885), .B1(new_n854), .B2(new_n888), .ZN(G397));
  NAND2_X1  g464(.A1(KEYINPUT124), .A2(KEYINPUT46), .ZN(new_n890));
  NAND3_X1  g465(.A1(new_n467), .A2(G40), .A3(new_n472), .ZN(new_n891));
  INV_X1    g466(.A(new_n891), .ZN(new_n892));
  INV_X1    g467(.A(G1384), .ZN(new_n893));
  AOI21_X1  g468(.A(KEYINPUT45), .B1(new_n496), .B2(new_n893), .ZN(new_n894));
  NAND2_X1  g469(.A1(new_n892), .A2(new_n894), .ZN(new_n895));
  NOR2_X1   g470(.A1(new_n895), .A2(G1996), .ZN(new_n896));
  INV_X1    g471(.A(new_n896), .ZN(new_n897));
  NOR2_X1   g472(.A1(KEYINPUT124), .A2(KEYINPUT46), .ZN(new_n898));
  OAI21_X1  g473(.A(new_n890), .B1(new_n897), .B2(new_n898), .ZN(new_n899));
  INV_X1    g474(.A(new_n895), .ZN(new_n900));
  NAND2_X1  g475(.A1(new_n767), .A2(G2067), .ZN(new_n901));
  INV_X1    g476(.A(G2067), .ZN(new_n902));
  NAND3_X1  g477(.A1(new_n761), .A2(new_n902), .A3(new_n766), .ZN(new_n903));
  NAND2_X1  g478(.A1(new_n901), .A2(new_n903), .ZN(new_n904));
  OAI21_X1  g479(.A(new_n900), .B1(new_n904), .B2(new_n730), .ZN(new_n905));
  OAI211_X1 g480(.A(new_n899), .B(new_n905), .C1(new_n897), .C2(new_n890), .ZN(new_n906));
  XOR2_X1   g481(.A(new_n906), .B(KEYINPUT47), .Z(new_n907));
  NAND3_X1  g482(.A1(new_n900), .A2(G1996), .A3(new_n730), .ZN(new_n908));
  XNOR2_X1  g483(.A(new_n908), .B(KEYINPUT106), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n896), .A2(new_n731), .ZN(new_n910));
  XNOR2_X1  g485(.A(new_n910), .B(KEYINPUT105), .ZN(new_n911));
  AOI211_X1 g486(.A(new_n909), .B(new_n911), .C1(new_n900), .C2(new_n904), .ZN(new_n912));
  AND2_X1   g487(.A1(new_n678), .A2(new_n680), .ZN(new_n913));
  NAND2_X1  g488(.A1(new_n912), .A2(new_n913), .ZN(new_n914));
  AOI21_X1  g489(.A(new_n895), .B1(new_n914), .B2(new_n903), .ZN(new_n915));
  NOR2_X1   g490(.A1(new_n678), .A2(new_n680), .ZN(new_n916));
  OAI21_X1  g491(.A(new_n900), .B1(new_n913), .B2(new_n916), .ZN(new_n917));
  AND2_X1   g492(.A1(new_n912), .A2(new_n917), .ZN(new_n918));
  NOR3_X1   g493(.A1(G290), .A2(new_n895), .A3(G1986), .ZN(new_n919));
  XOR2_X1   g494(.A(new_n919), .B(KEYINPUT48), .Z(new_n920));
  AOI211_X1 g495(.A(new_n907), .B(new_n915), .C1(new_n918), .C2(new_n920), .ZN(new_n921));
  INV_X1    g496(.A(G1981), .ZN(new_n922));
  AOI21_X1  g497(.A(new_n922), .B1(new_n572), .B2(KEYINPUT109), .ZN(new_n923));
  XNOR2_X1  g498(.A(new_n923), .B(G305), .ZN(new_n924));
  INV_X1    g499(.A(KEYINPUT49), .ZN(new_n925));
  NAND2_X1  g500(.A1(new_n924), .A2(new_n925), .ZN(new_n926));
  XOR2_X1   g501(.A(new_n926), .B(KEYINPUT110), .Z(new_n927));
  NAND2_X1  g502(.A1(new_n496), .A2(new_n893), .ZN(new_n928));
  NOR2_X1   g503(.A1(new_n928), .A2(new_n891), .ZN(new_n929));
  INV_X1    g504(.A(G8), .ZN(new_n930));
  NOR2_X1   g505(.A1(new_n929), .A2(new_n930), .ZN(new_n931));
  OAI21_X1  g506(.A(new_n931), .B1(new_n924), .B2(new_n925), .ZN(new_n932));
  NOR2_X1   g507(.A1(new_n927), .A2(new_n932), .ZN(new_n933));
  AOI21_X1  g508(.A(KEYINPUT108), .B1(new_n928), .B2(KEYINPUT50), .ZN(new_n934));
  INV_X1    g509(.A(KEYINPUT108), .ZN(new_n935));
  INV_X1    g510(.A(KEYINPUT50), .ZN(new_n936));
  AOI211_X1 g511(.A(new_n935), .B(new_n936), .C1(new_n496), .C2(new_n893), .ZN(new_n937));
  OR2_X1    g512(.A1(new_n934), .A2(new_n937), .ZN(new_n938));
  INV_X1    g513(.A(new_n488), .ZN(new_n939));
  OAI21_X1  g514(.A(new_n939), .B1(new_n460), .B2(new_n461), .ZN(new_n940));
  NAND2_X1  g515(.A1(new_n940), .A2(new_n490), .ZN(new_n941));
  AOI22_X1  g516(.A1(new_n941), .A2(new_n476), .B1(new_n494), .B2(new_n493), .ZN(new_n942));
  AOI21_X1  g517(.A(G1384), .B1(new_n942), .B2(new_n487), .ZN(new_n943));
  XNOR2_X1  g518(.A(KEYINPUT107), .B(KEYINPUT50), .ZN(new_n944));
  AOI21_X1  g519(.A(new_n891), .B1(new_n943), .B2(new_n944), .ZN(new_n945));
  NAND3_X1  g520(.A1(new_n938), .A2(new_n722), .A3(new_n945), .ZN(new_n946));
  NOR2_X1   g521(.A1(new_n894), .A2(new_n891), .ZN(new_n947));
  NAND3_X1  g522(.A1(new_n496), .A2(KEYINPUT45), .A3(new_n893), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n947), .A2(new_n948), .ZN(new_n949));
  NAND2_X1  g524(.A1(new_n949), .A2(new_n693), .ZN(new_n950));
  AOI21_X1  g525(.A(new_n930), .B1(new_n946), .B2(new_n950), .ZN(new_n951));
  INV_X1    g526(.A(new_n951), .ZN(new_n952));
  NAND2_X1  g527(.A1(G303), .A2(G8), .ZN(new_n953));
  XNOR2_X1  g528(.A(new_n953), .B(KEYINPUT55), .ZN(new_n954));
  OR2_X1    g529(.A1(new_n952), .A2(new_n954), .ZN(new_n955));
  INV_X1    g530(.A(G1976), .ZN(new_n956));
  AOI21_X1  g531(.A(KEYINPUT52), .B1(G288), .B2(new_n956), .ZN(new_n957));
  OAI21_X1  g532(.A(new_n931), .B1(new_n956), .B2(G288), .ZN(new_n958));
  MUX2_X1   g533(.A(new_n957), .B(KEYINPUT52), .S(new_n958), .Z(new_n959));
  NOR3_X1   g534(.A1(new_n933), .A2(new_n955), .A3(new_n959), .ZN(new_n960));
  NAND3_X1  g535(.A1(new_n568), .A2(new_n956), .A3(new_n569), .ZN(new_n961));
  OAI22_X1  g536(.A1(new_n933), .A2(new_n961), .B1(G1981), .B2(G305), .ZN(new_n962));
  INV_X1    g537(.A(KEYINPUT111), .ZN(new_n963));
  AOI211_X1 g538(.A(new_n930), .B(new_n929), .C1(new_n962), .C2(new_n963), .ZN(new_n964));
  OR2_X1    g539(.A1(new_n962), .A2(new_n963), .ZN(new_n965));
  AOI21_X1  g540(.A(new_n960), .B1(new_n964), .B2(new_n965), .ZN(new_n966));
  OR3_X1    g541(.A1(new_n933), .A2(KEYINPUT112), .A3(new_n959), .ZN(new_n967));
  NOR2_X1   g542(.A1(new_n943), .A2(new_n944), .ZN(new_n968));
  AOI211_X1 g543(.A(new_n891), .B(new_n968), .C1(new_n936), .C2(new_n943), .ZN(new_n969));
  AOI22_X1  g544(.A1(new_n969), .A2(new_n722), .B1(new_n693), .B2(new_n949), .ZN(new_n970));
  OAI21_X1  g545(.A(new_n954), .B1(new_n930), .B2(new_n970), .ZN(new_n971));
  OAI21_X1  g546(.A(KEYINPUT112), .B1(new_n933), .B2(new_n959), .ZN(new_n972));
  NAND4_X1  g547(.A1(new_n967), .A2(new_n955), .A3(new_n971), .A4(new_n972), .ZN(new_n973));
  INV_X1    g548(.A(new_n973), .ZN(new_n974));
  INV_X1    g549(.A(KEYINPUT113), .ZN(new_n975));
  AOI21_X1  g550(.A(new_n975), .B1(new_n943), .B2(KEYINPUT45), .ZN(new_n976));
  NAND4_X1  g551(.A1(new_n496), .A2(new_n975), .A3(KEYINPUT45), .A4(new_n893), .ZN(new_n977));
  INV_X1    g552(.A(new_n977), .ZN(new_n978));
  OAI21_X1  g553(.A(new_n947), .B1(new_n976), .B2(new_n978), .ZN(new_n979));
  NAND2_X1  g554(.A1(new_n979), .A2(new_n710), .ZN(new_n980));
  INV_X1    g555(.A(G2084), .ZN(new_n981));
  OAI211_X1 g556(.A(new_n945), .B(new_n981), .C1(new_n934), .C2(new_n937), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n980), .A2(new_n982), .ZN(new_n983));
  NAND2_X1  g558(.A1(new_n983), .A2(G8), .ZN(new_n984));
  NOR2_X1   g559(.A1(new_n984), .A2(G286), .ZN(new_n985));
  AOI21_X1  g560(.A(KEYINPUT63), .B1(new_n974), .B2(new_n985), .ZN(new_n986));
  NOR2_X1   g561(.A1(new_n933), .A2(new_n959), .ZN(new_n987));
  AOI211_X1 g562(.A(G286), .B(new_n984), .C1(new_n952), .C2(new_n954), .ZN(new_n988));
  AND4_X1   g563(.A1(KEYINPUT63), .A2(new_n987), .A3(new_n955), .A4(new_n988), .ZN(new_n989));
  OAI21_X1  g564(.A(new_n966), .B1(new_n986), .B2(new_n989), .ZN(new_n990));
  INV_X1    g565(.A(new_n949), .ZN(new_n991));
  AOI21_X1  g566(.A(KEYINPUT53), .B1(new_n991), .B2(new_n717), .ZN(new_n992));
  INV_X1    g567(.A(G1961), .ZN(new_n993));
  NAND2_X1  g568(.A1(new_n938), .A2(new_n945), .ZN(new_n994));
  AOI21_X1  g569(.A(new_n992), .B1(new_n993), .B2(new_n994), .ZN(new_n995));
  NAND2_X1  g570(.A1(new_n717), .A2(KEYINPUT53), .ZN(new_n996));
  OAI21_X1  g571(.A(new_n995), .B1(new_n979), .B2(new_n996), .ZN(new_n997));
  INV_X1    g572(.A(new_n997), .ZN(new_n998));
  NOR2_X1   g573(.A1(new_n998), .A2(G301), .ZN(new_n999));
  NOR2_X1   g574(.A1(G168), .A2(new_n930), .ZN(new_n1000));
  AOI211_X1 g575(.A(KEYINPUT51), .B(new_n1000), .C1(new_n983), .C2(G8), .ZN(new_n1001));
  INV_X1    g576(.A(new_n982), .ZN(new_n1002));
  NAND2_X1  g577(.A1(new_n948), .A2(KEYINPUT113), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n1003), .A2(new_n977), .ZN(new_n1004));
  AOI21_X1  g579(.A(G1966), .B1(new_n1004), .B2(new_n947), .ZN(new_n1005));
  NOR3_X1   g580(.A1(new_n1002), .A2(new_n1005), .A3(KEYINPUT118), .ZN(new_n1006));
  INV_X1    g581(.A(KEYINPUT118), .ZN(new_n1007));
  AOI21_X1  g582(.A(new_n1007), .B1(new_n980), .B2(new_n982), .ZN(new_n1008));
  OAI21_X1  g583(.A(G8), .B1(new_n1006), .B2(new_n1008), .ZN(new_n1009));
  INV_X1    g584(.A(KEYINPUT120), .ZN(new_n1010));
  NAND2_X1  g585(.A1(new_n1009), .A2(new_n1010), .ZN(new_n1011));
  OAI21_X1  g586(.A(KEYINPUT118), .B1(new_n1002), .B2(new_n1005), .ZN(new_n1012));
  NAND3_X1  g587(.A1(new_n980), .A2(new_n1007), .A3(new_n982), .ZN(new_n1013));
  AOI21_X1  g588(.A(new_n930), .B1(new_n1012), .B2(new_n1013), .ZN(new_n1014));
  NAND2_X1  g589(.A1(new_n1014), .A2(KEYINPUT120), .ZN(new_n1015));
  INV_X1    g590(.A(new_n1000), .ZN(new_n1016));
  NAND3_X1  g591(.A1(new_n1011), .A2(new_n1015), .A3(new_n1016), .ZN(new_n1017));
  XOR2_X1   g592(.A(KEYINPUT119), .B(KEYINPUT51), .Z(new_n1018));
  AOI21_X1  g593(.A(new_n1001), .B1(new_n1017), .B2(new_n1018), .ZN(new_n1019));
  AOI21_X1  g594(.A(new_n1016), .B1(new_n1012), .B2(new_n1013), .ZN(new_n1020));
  OAI21_X1  g595(.A(KEYINPUT121), .B1(new_n1019), .B2(new_n1020), .ZN(new_n1021));
  INV_X1    g596(.A(new_n1020), .ZN(new_n1022));
  INV_X1    g597(.A(KEYINPUT121), .ZN(new_n1023));
  INV_X1    g598(.A(new_n1018), .ZN(new_n1024));
  AOI21_X1  g599(.A(new_n1000), .B1(new_n1014), .B2(KEYINPUT120), .ZN(new_n1025));
  AOI21_X1  g600(.A(new_n1024), .B1(new_n1025), .B2(new_n1011), .ZN(new_n1026));
  OAI211_X1 g601(.A(new_n1022), .B(new_n1023), .C1(new_n1026), .C2(new_n1001), .ZN(new_n1027));
  AND3_X1   g602(.A1(new_n1021), .A2(KEYINPUT62), .A3(new_n1027), .ZN(new_n1028));
  AOI21_X1  g603(.A(KEYINPUT62), .B1(new_n1021), .B2(new_n1027), .ZN(new_n1029));
  OAI21_X1  g604(.A(new_n999), .B1(new_n1028), .B2(new_n1029), .ZN(new_n1030));
  XNOR2_X1  g605(.A(G171), .B(KEYINPUT54), .ZN(new_n1031));
  NAND2_X1  g606(.A1(new_n472), .A2(G40), .ZN(new_n1032));
  NOR2_X1   g607(.A1(new_n464), .A2(new_n466), .ZN(new_n1033));
  XOR2_X1   g608(.A(new_n1033), .B(KEYINPUT122), .Z(new_n1034));
  AOI21_X1  g609(.A(new_n1032), .B1(new_n1034), .B2(G2105), .ZN(new_n1035));
  INV_X1    g610(.A(KEYINPUT123), .ZN(new_n1036));
  OR2_X1    g611(.A1(new_n1035), .A2(new_n1036), .ZN(new_n1037));
  NAND2_X1  g612(.A1(new_n1035), .A2(new_n1036), .ZN(new_n1038));
  NOR2_X1   g613(.A1(new_n894), .A2(new_n996), .ZN(new_n1039));
  NAND4_X1  g614(.A1(new_n1037), .A2(new_n948), .A3(new_n1038), .A4(new_n1039), .ZN(new_n1040));
  NAND3_X1  g615(.A1(new_n995), .A2(new_n1031), .A3(new_n1040), .ZN(new_n1041));
  OAI21_X1  g616(.A(new_n1041), .B1(new_n998), .B2(new_n1031), .ZN(new_n1042));
  OR2_X1    g617(.A1(new_n949), .A2(G1996), .ZN(new_n1043));
  XOR2_X1   g618(.A(KEYINPUT58), .B(G1341), .Z(new_n1044));
  OAI21_X1  g619(.A(new_n1044), .B1(new_n928), .B2(new_n891), .ZN(new_n1045));
  AOI21_X1  g620(.A(new_n542), .B1(new_n1043), .B2(new_n1045), .ZN(new_n1046));
  XOR2_X1   g621(.A(new_n1046), .B(KEYINPUT59), .Z(new_n1047));
  INV_X1    g622(.A(KEYINPUT115), .ZN(new_n1048));
  INV_X1    g623(.A(KEYINPUT114), .ZN(new_n1049));
  AOI21_X1  g624(.A(new_n1048), .B1(G299), .B2(new_n1049), .ZN(new_n1050));
  INV_X1    g625(.A(KEYINPUT57), .ZN(new_n1051));
  NAND2_X1  g626(.A1(new_n1050), .A2(new_n1051), .ZN(new_n1052));
  OAI21_X1  g627(.A(KEYINPUT57), .B1(new_n564), .B2(KEYINPUT115), .ZN(new_n1053));
  OAI21_X1  g628(.A(new_n1052), .B1(new_n1050), .B2(new_n1053), .ZN(new_n1054));
  XOR2_X1   g629(.A(KEYINPUT56), .B(G2072), .Z(new_n1055));
  OAI22_X1  g630(.A1(new_n969), .A2(G1956), .B1(new_n949), .B2(new_n1055), .ZN(new_n1056));
  OR2_X1    g631(.A1(new_n1054), .A2(new_n1056), .ZN(new_n1057));
  NAND2_X1  g632(.A1(new_n1054), .A2(new_n1056), .ZN(new_n1058));
  NAND3_X1  g633(.A1(new_n1057), .A2(KEYINPUT61), .A3(new_n1058), .ZN(new_n1059));
  NAND2_X1  g634(.A1(new_n929), .A2(new_n902), .ZN(new_n1060));
  XNOR2_X1  g635(.A(new_n1060), .B(KEYINPUT116), .ZN(new_n1061));
  AOI21_X1  g636(.A(new_n1061), .B1(new_n779), .B2(new_n994), .ZN(new_n1062));
  INV_X1    g637(.A(KEYINPUT60), .ZN(new_n1063));
  NAND3_X1  g638(.A1(new_n1062), .A2(new_n1063), .A3(new_n591), .ZN(new_n1064));
  AND3_X1   g639(.A1(new_n1047), .A2(new_n1059), .A3(new_n1064), .ZN(new_n1065));
  AND2_X1   g640(.A1(new_n1062), .A2(new_n590), .ZN(new_n1066));
  NOR2_X1   g641(.A1(new_n1062), .A2(new_n590), .ZN(new_n1067));
  OAI21_X1  g642(.A(KEYINPUT60), .B1(new_n1066), .B2(new_n1067), .ZN(new_n1068));
  NAND2_X1  g643(.A1(new_n1057), .A2(new_n1058), .ZN(new_n1069));
  INV_X1    g644(.A(KEYINPUT61), .ZN(new_n1070));
  AND3_X1   g645(.A1(new_n1069), .A2(KEYINPUT117), .A3(new_n1070), .ZN(new_n1071));
  AOI21_X1  g646(.A(KEYINPUT117), .B1(new_n1069), .B2(new_n1070), .ZN(new_n1072));
  OAI211_X1 g647(.A(new_n1065), .B(new_n1068), .C1(new_n1071), .C2(new_n1072), .ZN(new_n1073));
  INV_X1    g648(.A(new_n1058), .ZN(new_n1074));
  AOI21_X1  g649(.A(new_n1074), .B1(new_n1067), .B2(new_n1057), .ZN(new_n1075));
  AOI21_X1  g650(.A(new_n1042), .B1(new_n1073), .B2(new_n1075), .ZN(new_n1076));
  NAND2_X1  g651(.A1(new_n1021), .A2(new_n1027), .ZN(new_n1077));
  NAND2_X1  g652(.A1(new_n1076), .A2(new_n1077), .ZN(new_n1078));
  NAND2_X1  g653(.A1(new_n1030), .A2(new_n1078), .ZN(new_n1079));
  AOI21_X1  g654(.A(new_n990), .B1(new_n1079), .B2(new_n974), .ZN(new_n1080));
  XOR2_X1   g655(.A(G290), .B(G1986), .Z(new_n1081));
  OAI21_X1  g656(.A(new_n918), .B1(new_n895), .B2(new_n1081), .ZN(new_n1082));
  OAI21_X1  g657(.A(new_n921), .B1(new_n1080), .B2(new_n1082), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g658(.A(KEYINPUT126), .ZN(new_n1085));
  INV_X1    g659(.A(KEYINPUT125), .ZN(new_n1086));
  OR2_X1    g660(.A1(G227), .A2(new_n457), .ZN(new_n1087));
  OAI21_X1  g661(.A(new_n1086), .B1(G401), .B2(new_n1087), .ZN(new_n1088));
  NAND2_X1  g662(.A1(new_n1088), .A2(new_n671), .ZN(new_n1089));
  NOR3_X1   g663(.A1(G401), .A2(new_n1086), .A3(new_n1087), .ZN(new_n1090));
  OAI21_X1  g664(.A(new_n1085), .B1(new_n1089), .B2(new_n1090), .ZN(new_n1091));
  AOI21_X1  g665(.A(new_n1087), .B1(new_n636), .B2(new_n634), .ZN(new_n1092));
  NAND2_X1  g666(.A1(new_n1092), .A2(KEYINPUT125), .ZN(new_n1093));
  NAND4_X1  g667(.A1(new_n1093), .A2(KEYINPUT126), .A3(new_n671), .A4(new_n1088), .ZN(new_n1094));
  AND3_X1   g668(.A1(new_n1091), .A2(new_n821), .A3(new_n1094), .ZN(new_n1095));
  INV_X1    g669(.A(KEYINPUT127), .ZN(new_n1096));
  NAND4_X1  g670(.A1(new_n1095), .A2(new_n1096), .A3(new_n886), .A4(new_n887), .ZN(new_n1097));
  NAND3_X1  g671(.A1(new_n1091), .A2(new_n1094), .A3(new_n821), .ZN(new_n1098));
  OAI21_X1  g672(.A(KEYINPUT127), .B1(new_n888), .B2(new_n1098), .ZN(new_n1099));
  AND2_X1   g673(.A1(new_n1097), .A2(new_n1099), .ZN(G308));
  NAND2_X1  g674(.A1(new_n1097), .A2(new_n1099), .ZN(G225));
endmodule


