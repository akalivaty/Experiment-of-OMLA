//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 0 0 1 1 0 0 0 0 1 1 1 0 1 1 0 0 0 0 0 0 0 1 0 0 1 0 0 0 0 0 1 0 1 0 0 1 0 1 1 0 0 1 1 1 0 1 1 0 1 0 1 1 1 1 0 1 1 1 1 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:20:12 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n750, new_n751, new_n752, new_n753, new_n754, new_n755, new_n757,
    new_n758, new_n759, new_n760, new_n761, new_n762, new_n763, new_n764,
    new_n765, new_n766, new_n767, new_n768, new_n769, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n798, new_n799, new_n800, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n809, new_n810,
    new_n811, new_n812, new_n813, new_n814, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n848, new_n850,
    new_n851, new_n852, new_n853, new_n854, new_n855, new_n856, new_n857,
    new_n858, new_n859, new_n860, new_n861, new_n862, new_n863, new_n864,
    new_n865, new_n866, new_n867, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n885, new_n886, new_n887,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n906, new_n907, new_n908, new_n909, new_n910,
    new_n911, new_n912, new_n913, new_n914, new_n915, new_n916, new_n917,
    new_n918, new_n919, new_n920, new_n921, new_n922, new_n923, new_n924,
    new_n925, new_n926, new_n927, new_n928, new_n929, new_n930, new_n931,
    new_n932, new_n934, new_n935, new_n937, new_n938, new_n940, new_n941,
    new_n942, new_n943, new_n944, new_n945, new_n946, new_n948, new_n949,
    new_n950, new_n951, new_n952, new_n953, new_n954, new_n955, new_n956,
    new_n957, new_n958, new_n959, new_n960, new_n961, new_n962, new_n963,
    new_n964, new_n965, new_n966, new_n968, new_n969, new_n970, new_n971,
    new_n972, new_n973, new_n974, new_n975, new_n976, new_n978, new_n979,
    new_n981, new_n982, new_n983, new_n984, new_n985, new_n986, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n999, new_n1000, new_n1001, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1017, new_n1018, new_n1019, new_n1020, new_n1021, new_n1022,
    new_n1023, new_n1024, new_n1026, new_n1027, new_n1028, new_n1029,
    new_n1030, new_n1031, new_n1032, new_n1033, new_n1035, new_n1036,
    new_n1037, new_n1038, new_n1040, new_n1041, new_n1042, new_n1043,
    new_n1044, new_n1045, new_n1046, new_n1047, new_n1049, new_n1050,
    new_n1051, new_n1052;
  NAND3_X1  g000(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n202));
  NAND2_X1  g001(.A1(G85gat), .A2(G92gat), .ZN(new_n203));
  XNOR2_X1  g002(.A(new_n203), .B(KEYINPUT7), .ZN(new_n204));
  NAND2_X1  g003(.A1(G99gat), .A2(G106gat), .ZN(new_n205));
  INV_X1    g004(.A(G85gat), .ZN(new_n206));
  INV_X1    g005(.A(G92gat), .ZN(new_n207));
  AOI22_X1  g006(.A1(KEYINPUT8), .A2(new_n205), .B1(new_n206), .B2(new_n207), .ZN(new_n208));
  NAND2_X1  g007(.A1(new_n204), .A2(new_n208), .ZN(new_n209));
  XNOR2_X1  g008(.A(G99gat), .B(G106gat), .ZN(new_n210));
  XOR2_X1   g009(.A(new_n209), .B(new_n210), .Z(new_n211));
  INV_X1    g010(.A(new_n211), .ZN(new_n212));
  XOR2_X1   g011(.A(G43gat), .B(G50gat), .Z(new_n213));
  INV_X1    g012(.A(KEYINPUT93), .ZN(new_n214));
  NAND2_X1  g013(.A1(new_n213), .A2(new_n214), .ZN(new_n215));
  XNOR2_X1  g014(.A(G43gat), .B(G50gat), .ZN(new_n216));
  NAND2_X1  g015(.A1(new_n216), .A2(KEYINPUT93), .ZN(new_n217));
  NAND3_X1  g016(.A1(new_n215), .A2(KEYINPUT15), .A3(new_n217), .ZN(new_n218));
  NOR2_X1   g017(.A1(G29gat), .A2(G36gat), .ZN(new_n219));
  NAND2_X1  g018(.A1(new_n219), .A2(KEYINPUT14), .ZN(new_n220));
  INV_X1    g019(.A(KEYINPUT14), .ZN(new_n221));
  AOI21_X1  g020(.A(new_n221), .B1(G29gat), .B2(G36gat), .ZN(new_n222));
  OAI21_X1  g021(.A(new_n220), .B1(new_n222), .B2(new_n219), .ZN(new_n223));
  INV_X1    g022(.A(new_n223), .ZN(new_n224));
  OAI211_X1 g023(.A(new_n218), .B(new_n224), .C1(KEYINPUT15), .C2(new_n216), .ZN(new_n225));
  AND3_X1   g024(.A1(new_n215), .A2(KEYINPUT15), .A3(new_n217), .ZN(new_n226));
  AOI21_X1  g025(.A(KEYINPUT94), .B1(new_n226), .B2(new_n223), .ZN(new_n227));
  INV_X1    g026(.A(KEYINPUT94), .ZN(new_n228));
  NOR3_X1   g027(.A1(new_n218), .A2(new_n228), .A3(new_n224), .ZN(new_n229));
  OAI21_X1  g028(.A(new_n225), .B1(new_n227), .B2(new_n229), .ZN(new_n230));
  INV_X1    g029(.A(KEYINPUT95), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n230), .A2(new_n231), .ZN(new_n232));
  INV_X1    g031(.A(KEYINPUT17), .ZN(new_n233));
  OAI211_X1 g032(.A(KEYINPUT95), .B(new_n225), .C1(new_n227), .C2(new_n229), .ZN(new_n234));
  NAND3_X1  g033(.A1(new_n232), .A2(new_n233), .A3(new_n234), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n230), .A2(KEYINPUT17), .ZN(new_n236));
  AOI21_X1  g035(.A(new_n212), .B1(new_n235), .B2(new_n236), .ZN(new_n237));
  OAI21_X1  g036(.A(new_n202), .B1(new_n237), .B2(KEYINPUT103), .ZN(new_n238));
  NAND2_X1  g037(.A1(new_n232), .A2(new_n234), .ZN(new_n239));
  INV_X1    g038(.A(new_n239), .ZN(new_n240));
  NOR2_X1   g039(.A1(new_n240), .A2(new_n211), .ZN(new_n241));
  INV_X1    g040(.A(KEYINPUT103), .ZN(new_n242));
  AOI211_X1 g041(.A(new_n242), .B(new_n212), .C1(new_n235), .C2(new_n236), .ZN(new_n243));
  NOR3_X1   g042(.A1(new_n238), .A2(new_n241), .A3(new_n243), .ZN(new_n244));
  XOR2_X1   g043(.A(G190gat), .B(G218gat), .Z(new_n245));
  NOR3_X1   g044(.A1(new_n244), .A2(KEYINPUT105), .A3(new_n245), .ZN(new_n246));
  INV_X1    g045(.A(KEYINPUT105), .ZN(new_n247));
  NAND2_X1  g046(.A1(new_n235), .A2(new_n236), .ZN(new_n248));
  NAND2_X1  g047(.A1(new_n248), .A2(new_n211), .ZN(new_n249));
  NAND2_X1  g048(.A1(new_n249), .A2(new_n242), .ZN(new_n250));
  INV_X1    g049(.A(new_n241), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n237), .A2(KEYINPUT103), .ZN(new_n252));
  NAND4_X1  g051(.A1(new_n250), .A2(new_n251), .A3(new_n252), .A4(new_n202), .ZN(new_n253));
  INV_X1    g052(.A(new_n245), .ZN(new_n254));
  AOI21_X1  g053(.A(new_n247), .B1(new_n253), .B2(new_n254), .ZN(new_n255));
  NOR2_X1   g054(.A1(new_n246), .A2(new_n255), .ZN(new_n256));
  NAND2_X1  g055(.A1(new_n244), .A2(new_n245), .ZN(new_n257));
  INV_X1    g056(.A(KEYINPUT104), .ZN(new_n258));
  AOI21_X1  g057(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n259));
  XNOR2_X1  g058(.A(new_n259), .B(G134gat), .ZN(new_n260));
  INV_X1    g059(.A(G162gat), .ZN(new_n261));
  XNOR2_X1  g060(.A(new_n260), .B(new_n261), .ZN(new_n262));
  INV_X1    g061(.A(new_n262), .ZN(new_n263));
  OAI211_X1 g062(.A(new_n256), .B(new_n257), .C1(new_n258), .C2(new_n263), .ZN(new_n264));
  OAI21_X1  g063(.A(KEYINPUT105), .B1(new_n244), .B2(new_n245), .ZN(new_n265));
  NAND3_X1  g064(.A1(new_n253), .A2(new_n247), .A3(new_n254), .ZN(new_n266));
  NAND3_X1  g065(.A1(new_n265), .A2(new_n257), .A3(new_n266), .ZN(new_n267));
  NAND3_X1  g066(.A1(new_n265), .A2(new_n258), .A3(new_n266), .ZN(new_n268));
  NAND3_X1  g067(.A1(new_n267), .A2(new_n268), .A3(new_n262), .ZN(new_n269));
  INV_X1    g068(.A(G57gat), .ZN(new_n270));
  INV_X1    g069(.A(G64gat), .ZN(new_n271));
  NAND2_X1  g070(.A1(new_n270), .A2(new_n271), .ZN(new_n272));
  NAND2_X1  g071(.A1(G57gat), .A2(G64gat), .ZN(new_n273));
  NAND2_X1  g072(.A1(G71gat), .A2(G78gat), .ZN(new_n274));
  INV_X1    g073(.A(new_n274), .ZN(new_n275));
  OAI211_X1 g074(.A(new_n272), .B(new_n273), .C1(new_n275), .C2(KEYINPUT9), .ZN(new_n276));
  OAI21_X1  g075(.A(KEYINPUT96), .B1(G71gat), .B2(G78gat), .ZN(new_n277));
  INV_X1    g076(.A(new_n277), .ZN(new_n278));
  NOR3_X1   g077(.A1(KEYINPUT96), .A2(G71gat), .A3(G78gat), .ZN(new_n279));
  OAI21_X1  g078(.A(new_n274), .B1(new_n278), .B2(new_n279), .ZN(new_n280));
  NOR2_X1   g079(.A1(new_n280), .A2(KEYINPUT97), .ZN(new_n281));
  INV_X1    g080(.A(KEYINPUT97), .ZN(new_n282));
  NOR2_X1   g081(.A1(G71gat), .A2(G78gat), .ZN(new_n283));
  INV_X1    g082(.A(KEYINPUT96), .ZN(new_n284));
  NAND2_X1  g083(.A1(new_n283), .A2(new_n284), .ZN(new_n285));
  NAND2_X1  g084(.A1(new_n285), .A2(new_n277), .ZN(new_n286));
  AOI21_X1  g085(.A(new_n282), .B1(new_n286), .B2(new_n274), .ZN(new_n287));
  OAI21_X1  g086(.A(new_n276), .B1(new_n281), .B2(new_n287), .ZN(new_n288));
  NAND2_X1  g087(.A1(new_n288), .A2(KEYINPUT98), .ZN(new_n289));
  INV_X1    g088(.A(KEYINPUT98), .ZN(new_n290));
  OAI211_X1 g089(.A(new_n290), .B(new_n276), .C1(new_n281), .C2(new_n287), .ZN(new_n291));
  NAND2_X1  g090(.A1(new_n289), .A2(new_n291), .ZN(new_n292));
  INV_X1    g091(.A(KEYINPUT99), .ZN(new_n293));
  NAND2_X1  g092(.A1(new_n293), .A2(G57gat), .ZN(new_n294));
  XNOR2_X1  g093(.A(new_n294), .B(new_n271), .ZN(new_n295));
  AOI21_X1  g094(.A(new_n275), .B1(KEYINPUT9), .B2(new_n283), .ZN(new_n296));
  NOR2_X1   g095(.A1(new_n295), .A2(new_n296), .ZN(new_n297));
  INV_X1    g096(.A(new_n297), .ZN(new_n298));
  AOI21_X1  g097(.A(KEYINPUT100), .B1(new_n292), .B2(new_n298), .ZN(new_n299));
  INV_X1    g098(.A(KEYINPUT100), .ZN(new_n300));
  AOI211_X1 g099(.A(new_n300), .B(new_n297), .C1(new_n289), .C2(new_n291), .ZN(new_n301));
  INV_X1    g100(.A(KEYINPUT21), .ZN(new_n302));
  NOR3_X1   g101(.A1(new_n299), .A2(new_n301), .A3(new_n302), .ZN(new_n303));
  XNOR2_X1  g102(.A(G15gat), .B(G22gat), .ZN(new_n304));
  INV_X1    g103(.A(KEYINPUT16), .ZN(new_n305));
  OAI21_X1  g104(.A(new_n304), .B1(new_n305), .B2(G1gat), .ZN(new_n306));
  OAI21_X1  g105(.A(new_n306), .B1(G1gat), .B2(new_n304), .ZN(new_n307));
  INV_X1    g106(.A(G8gat), .ZN(new_n308));
  XNOR2_X1  g107(.A(new_n307), .B(new_n308), .ZN(new_n309));
  INV_X1    g108(.A(new_n309), .ZN(new_n310));
  OAI21_X1  g109(.A(KEYINPUT102), .B1(new_n303), .B2(new_n310), .ZN(new_n311));
  INV_X1    g110(.A(KEYINPUT101), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n292), .A2(new_n298), .ZN(new_n313));
  NAND2_X1  g112(.A1(new_n313), .A2(new_n300), .ZN(new_n314));
  NAND3_X1  g113(.A1(new_n292), .A2(KEYINPUT100), .A3(new_n298), .ZN(new_n315));
  NAND3_X1  g114(.A1(new_n314), .A2(KEYINPUT21), .A3(new_n315), .ZN(new_n316));
  INV_X1    g115(.A(KEYINPUT102), .ZN(new_n317));
  NAND3_X1  g116(.A1(new_n316), .A2(new_n317), .A3(new_n309), .ZN(new_n318));
  NAND3_X1  g117(.A1(new_n311), .A2(new_n312), .A3(new_n318), .ZN(new_n319));
  INV_X1    g118(.A(new_n319), .ZN(new_n320));
  AOI21_X1  g119(.A(new_n312), .B1(new_n311), .B2(new_n318), .ZN(new_n321));
  INV_X1    g120(.A(KEYINPUT19), .ZN(new_n322));
  NOR3_X1   g121(.A1(new_n320), .A2(new_n321), .A3(new_n322), .ZN(new_n323));
  INV_X1    g122(.A(new_n318), .ZN(new_n324));
  AOI21_X1  g123(.A(new_n317), .B1(new_n316), .B2(new_n309), .ZN(new_n325));
  OAI21_X1  g124(.A(KEYINPUT101), .B1(new_n324), .B2(new_n325), .ZN(new_n326));
  AOI21_X1  g125(.A(KEYINPUT19), .B1(new_n326), .B2(new_n319), .ZN(new_n327));
  XNOR2_X1  g126(.A(G127gat), .B(G155gat), .ZN(new_n328));
  XOR2_X1   g127(.A(new_n328), .B(KEYINPUT20), .Z(new_n329));
  NOR3_X1   g128(.A1(new_n323), .A2(new_n327), .A3(new_n329), .ZN(new_n330));
  INV_X1    g129(.A(new_n329), .ZN(new_n331));
  OAI21_X1  g130(.A(new_n322), .B1(new_n320), .B2(new_n321), .ZN(new_n332));
  NAND3_X1  g131(.A1(new_n326), .A2(KEYINPUT19), .A3(new_n319), .ZN(new_n333));
  AOI21_X1  g132(.A(new_n331), .B1(new_n332), .B2(new_n333), .ZN(new_n334));
  OAI21_X1  g133(.A(new_n302), .B1(new_n299), .B2(new_n301), .ZN(new_n335));
  XOR2_X1   g134(.A(G183gat), .B(G211gat), .Z(new_n336));
  NAND2_X1  g135(.A1(G231gat), .A2(G233gat), .ZN(new_n337));
  XNOR2_X1  g136(.A(new_n336), .B(new_n337), .ZN(new_n338));
  XNOR2_X1  g137(.A(new_n335), .B(new_n338), .ZN(new_n339));
  INV_X1    g138(.A(new_n339), .ZN(new_n340));
  NOR3_X1   g139(.A1(new_n330), .A2(new_n334), .A3(new_n340), .ZN(new_n341));
  OAI21_X1  g140(.A(new_n329), .B1(new_n323), .B2(new_n327), .ZN(new_n342));
  NAND3_X1  g141(.A1(new_n332), .A2(new_n331), .A3(new_n333), .ZN(new_n343));
  AOI21_X1  g142(.A(new_n339), .B1(new_n342), .B2(new_n343), .ZN(new_n344));
  OAI211_X1 g143(.A(new_n264), .B(new_n269), .C1(new_n341), .C2(new_n344), .ZN(new_n345));
  INV_X1    g144(.A(G127gat), .ZN(new_n346));
  INV_X1    g145(.A(G134gat), .ZN(new_n347));
  NAND2_X1  g146(.A1(new_n346), .A2(new_n347), .ZN(new_n348));
  NAND2_X1  g147(.A1(G127gat), .A2(G134gat), .ZN(new_n349));
  AOI21_X1  g148(.A(KEYINPUT1), .B1(new_n348), .B2(new_n349), .ZN(new_n350));
  INV_X1    g149(.A(KEYINPUT69), .ZN(new_n351));
  INV_X1    g150(.A(G113gat), .ZN(new_n352));
  OAI21_X1  g151(.A(new_n351), .B1(new_n352), .B2(G120gat), .ZN(new_n353));
  INV_X1    g152(.A(G120gat), .ZN(new_n354));
  NAND3_X1  g153(.A1(new_n354), .A2(KEYINPUT69), .A3(G113gat), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n353), .A2(new_n355), .ZN(new_n356));
  NOR2_X1   g155(.A1(new_n354), .A2(G113gat), .ZN(new_n357));
  OAI21_X1  g156(.A(new_n350), .B1(new_n356), .B2(new_n357), .ZN(new_n358));
  INV_X1    g157(.A(KEYINPUT1), .ZN(new_n359));
  NOR2_X1   g158(.A1(new_n352), .A2(G120gat), .ZN(new_n360));
  OAI21_X1  g159(.A(new_n359), .B1(new_n357), .B2(new_n360), .ZN(new_n361));
  AND2_X1   g160(.A1(new_n348), .A2(new_n349), .ZN(new_n362));
  NAND2_X1  g161(.A1(new_n361), .A2(new_n362), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n358), .A2(new_n363), .ZN(new_n364));
  INV_X1    g163(.A(new_n364), .ZN(new_n365));
  NAND2_X1  g164(.A1(G183gat), .A2(G190gat), .ZN(new_n366));
  NAND2_X1  g165(.A1(G169gat), .A2(G176gat), .ZN(new_n367));
  INV_X1    g166(.A(KEYINPUT66), .ZN(new_n368));
  NAND2_X1  g167(.A1(new_n367), .A2(new_n368), .ZN(new_n369));
  NAND3_X1  g168(.A1(KEYINPUT66), .A2(G169gat), .A3(G176gat), .ZN(new_n370));
  NAND2_X1  g169(.A1(new_n369), .A2(new_n370), .ZN(new_n371));
  OAI21_X1  g170(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n372));
  NOR2_X1   g171(.A1(G169gat), .A2(G176gat), .ZN(new_n373));
  INV_X1    g172(.A(KEYINPUT26), .ZN(new_n374));
  NAND2_X1  g173(.A1(new_n373), .A2(new_n374), .ZN(new_n375));
  NAND3_X1  g174(.A1(new_n371), .A2(new_n372), .A3(new_n375), .ZN(new_n376));
  INV_X1    g175(.A(KEYINPUT28), .ZN(new_n377));
  NOR2_X1   g176(.A1(new_n377), .A2(G190gat), .ZN(new_n378));
  INV_X1    g177(.A(new_n378), .ZN(new_n379));
  AND2_X1   g178(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n380));
  NOR2_X1   g179(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n381));
  OAI21_X1  g180(.A(KEYINPUT68), .B1(new_n380), .B2(new_n381), .ZN(new_n382));
  INV_X1    g181(.A(KEYINPUT27), .ZN(new_n383));
  INV_X1    g182(.A(G183gat), .ZN(new_n384));
  NAND2_X1  g183(.A1(new_n383), .A2(new_n384), .ZN(new_n385));
  INV_X1    g184(.A(KEYINPUT68), .ZN(new_n386));
  NAND2_X1  g185(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n387));
  NAND3_X1  g186(.A1(new_n385), .A2(new_n386), .A3(new_n387), .ZN(new_n388));
  AOI21_X1  g187(.A(new_n379), .B1(new_n382), .B2(new_n388), .ZN(new_n389));
  NAND2_X1  g188(.A1(new_n385), .A2(new_n387), .ZN(new_n390));
  INV_X1    g189(.A(G190gat), .ZN(new_n391));
  AOI21_X1  g190(.A(KEYINPUT28), .B1(new_n390), .B2(new_n391), .ZN(new_n392));
  OAI211_X1 g191(.A(new_n366), .B(new_n376), .C1(new_n389), .C2(new_n392), .ZN(new_n393));
  INV_X1    g192(.A(G169gat), .ZN(new_n394));
  INV_X1    g193(.A(G176gat), .ZN(new_n395));
  NAND3_X1  g194(.A1(new_n394), .A2(new_n395), .A3(KEYINPUT23), .ZN(new_n396));
  NAND2_X1  g195(.A1(new_n396), .A2(KEYINPUT65), .ZN(new_n397));
  INV_X1    g196(.A(KEYINPUT65), .ZN(new_n398));
  NAND3_X1  g197(.A1(new_n373), .A2(new_n398), .A3(KEYINPUT23), .ZN(new_n399));
  AND2_X1   g198(.A1(new_n397), .A2(new_n399), .ZN(new_n400));
  AOI21_X1  g199(.A(KEYINPUT25), .B1(new_n369), .B2(new_n370), .ZN(new_n401));
  INV_X1    g200(.A(KEYINPUT64), .ZN(new_n402));
  NAND3_X1  g201(.A1(new_n402), .A2(new_n384), .A3(new_n391), .ZN(new_n403));
  OAI21_X1  g202(.A(KEYINPUT64), .B1(G183gat), .B2(G190gat), .ZN(new_n404));
  NAND2_X1  g203(.A1(new_n403), .A2(new_n404), .ZN(new_n405));
  NAND2_X1  g204(.A1(new_n366), .A2(KEYINPUT24), .ZN(new_n406));
  INV_X1    g205(.A(KEYINPUT24), .ZN(new_n407));
  NAND3_X1  g206(.A1(new_n407), .A2(G183gat), .A3(G190gat), .ZN(new_n408));
  NAND2_X1  g207(.A1(new_n406), .A2(new_n408), .ZN(new_n409));
  NAND2_X1  g208(.A1(new_n405), .A2(new_n409), .ZN(new_n410));
  INV_X1    g209(.A(KEYINPUT23), .ZN(new_n411));
  OAI21_X1  g210(.A(new_n411), .B1(G169gat), .B2(G176gat), .ZN(new_n412));
  NAND4_X1  g211(.A1(new_n400), .A2(new_n401), .A3(new_n410), .A4(new_n412), .ZN(new_n413));
  NAND2_X1  g212(.A1(new_n393), .A2(new_n413), .ZN(new_n414));
  INV_X1    g213(.A(KEYINPUT25), .ZN(new_n415));
  NAND2_X1  g214(.A1(new_n396), .A2(new_n412), .ZN(new_n416));
  AOI21_X1  g215(.A(KEYINPUT67), .B1(G183gat), .B2(G190gat), .ZN(new_n417));
  XNOR2_X1  g216(.A(new_n417), .B(KEYINPUT24), .ZN(new_n418));
  NAND2_X1  g217(.A1(new_n384), .A2(new_n391), .ZN(new_n419));
  AOI21_X1  g218(.A(new_n416), .B1(new_n418), .B2(new_n419), .ZN(new_n420));
  AOI21_X1  g219(.A(new_n415), .B1(new_n420), .B2(new_n371), .ZN(new_n421));
  OAI21_X1  g220(.A(new_n365), .B1(new_n414), .B2(new_n421), .ZN(new_n422));
  INV_X1    g221(.A(KEYINPUT67), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n366), .A2(new_n423), .ZN(new_n424));
  NAND2_X1  g223(.A1(new_n424), .A2(KEYINPUT24), .ZN(new_n425));
  NAND2_X1  g224(.A1(new_n417), .A2(new_n407), .ZN(new_n426));
  NAND3_X1  g225(.A1(new_n425), .A2(new_n419), .A3(new_n426), .ZN(new_n427));
  NAND4_X1  g226(.A1(new_n427), .A2(new_n371), .A3(new_n412), .A4(new_n396), .ZN(new_n428));
  NAND2_X1  g227(.A1(new_n428), .A2(KEYINPUT25), .ZN(new_n429));
  NAND4_X1  g228(.A1(new_n429), .A2(new_n364), .A3(new_n393), .A4(new_n413), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n422), .A2(new_n430), .ZN(new_n431));
  INV_X1    g230(.A(G227gat), .ZN(new_n432));
  INV_X1    g231(.A(G233gat), .ZN(new_n433));
  NOR2_X1   g232(.A1(new_n432), .A2(new_n433), .ZN(new_n434));
  INV_X1    g233(.A(new_n434), .ZN(new_n435));
  NAND2_X1  g234(.A1(new_n431), .A2(new_n435), .ZN(new_n436));
  AND2_X1   g235(.A1(new_n436), .A2(KEYINPUT34), .ZN(new_n437));
  NOR2_X1   g236(.A1(new_n436), .A2(KEYINPUT34), .ZN(new_n438));
  NOR2_X1   g237(.A1(new_n437), .A2(new_n438), .ZN(new_n439));
  INV_X1    g238(.A(new_n439), .ZN(new_n440));
  INV_X1    g239(.A(KEYINPUT32), .ZN(new_n441));
  NAND3_X1  g240(.A1(new_n422), .A2(new_n434), .A3(new_n430), .ZN(new_n442));
  INV_X1    g241(.A(KEYINPUT70), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  NAND4_X1  g243(.A1(new_n422), .A2(KEYINPUT70), .A3(new_n434), .A4(new_n430), .ZN(new_n445));
  AOI21_X1  g244(.A(new_n441), .B1(new_n444), .B2(new_n445), .ZN(new_n446));
  AOI21_X1  g245(.A(KEYINPUT33), .B1(new_n444), .B2(new_n445), .ZN(new_n447));
  XNOR2_X1  g246(.A(G15gat), .B(G43gat), .ZN(new_n448));
  XNOR2_X1  g247(.A(G71gat), .B(G99gat), .ZN(new_n449));
  XOR2_X1   g248(.A(new_n448), .B(new_n449), .Z(new_n450));
  INV_X1    g249(.A(new_n450), .ZN(new_n451));
  NOR3_X1   g250(.A1(new_n446), .A2(new_n447), .A3(new_n451), .ZN(new_n452));
  AOI221_X4 g251(.A(new_n441), .B1(KEYINPUT33), .B2(new_n450), .C1(new_n444), .C2(new_n445), .ZN(new_n453));
  OAI21_X1  g252(.A(new_n440), .B1(new_n452), .B2(new_n453), .ZN(new_n454));
  INV_X1    g253(.A(KEYINPUT71), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n444), .A2(new_n445), .ZN(new_n456));
  INV_X1    g255(.A(KEYINPUT33), .ZN(new_n457));
  AOI21_X1  g256(.A(new_n451), .B1(new_n456), .B2(new_n457), .ZN(new_n458));
  INV_X1    g257(.A(new_n446), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  INV_X1    g259(.A(new_n453), .ZN(new_n461));
  NAND3_X1  g260(.A1(new_n460), .A2(new_n461), .A3(new_n439), .ZN(new_n462));
  NAND3_X1  g261(.A1(new_n454), .A2(new_n455), .A3(new_n462), .ZN(new_n463));
  AOI21_X1  g262(.A(new_n439), .B1(new_n460), .B2(new_n461), .ZN(new_n464));
  NAND2_X1  g263(.A1(new_n464), .A2(KEYINPUT71), .ZN(new_n465));
  NAND2_X1  g264(.A1(new_n463), .A2(new_n465), .ZN(new_n466));
  XOR2_X1   g265(.A(G78gat), .B(G106gat), .Z(new_n467));
  XNOR2_X1  g266(.A(new_n467), .B(G50gat), .ZN(new_n468));
  XNOR2_X1  g267(.A(new_n468), .B(KEYINPUT83), .ZN(new_n469));
  XOR2_X1   g268(.A(new_n469), .B(KEYINPUT31), .Z(new_n470));
  INV_X1    g269(.A(G22gat), .ZN(new_n471));
  NAND2_X1  g270(.A1(G211gat), .A2(G218gat), .ZN(new_n472));
  INV_X1    g271(.A(KEYINPUT22), .ZN(new_n473));
  NAND2_X1  g272(.A1(new_n472), .A2(new_n473), .ZN(new_n474));
  NAND2_X1  g273(.A1(new_n474), .A2(KEYINPUT73), .ZN(new_n475));
  XNOR2_X1  g274(.A(G197gat), .B(G204gat), .ZN(new_n476));
  INV_X1    g275(.A(KEYINPUT73), .ZN(new_n477));
  NAND3_X1  g276(.A1(new_n472), .A2(new_n477), .A3(new_n473), .ZN(new_n478));
  NAND3_X1  g277(.A1(new_n475), .A2(new_n476), .A3(new_n478), .ZN(new_n479));
  XOR2_X1   g278(.A(G211gat), .B(G218gat), .Z(new_n480));
  INV_X1    g279(.A(new_n480), .ZN(new_n481));
  AND3_X1   g280(.A1(new_n479), .A2(KEYINPUT74), .A3(new_n481), .ZN(new_n482));
  AOI21_X1  g281(.A(new_n481), .B1(new_n479), .B2(KEYINPUT74), .ZN(new_n483));
  NOR2_X1   g282(.A1(new_n482), .A2(new_n483), .ZN(new_n484));
  INV_X1    g283(.A(KEYINPUT2), .ZN(new_n485));
  INV_X1    g284(.A(G141gat), .ZN(new_n486));
  NAND2_X1  g285(.A1(new_n486), .A2(G148gat), .ZN(new_n487));
  INV_X1    g286(.A(new_n487), .ZN(new_n488));
  NOR2_X1   g287(.A1(new_n486), .A2(G148gat), .ZN(new_n489));
  OAI21_X1  g288(.A(new_n485), .B1(new_n488), .B2(new_n489), .ZN(new_n490));
  INV_X1    g289(.A(G155gat), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n491), .A2(new_n261), .ZN(new_n492));
  NAND2_X1  g291(.A1(G155gat), .A2(G162gat), .ZN(new_n493));
  AND2_X1   g292(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  INV_X1    g293(.A(KEYINPUT78), .ZN(new_n495));
  OAI21_X1  g294(.A(new_n495), .B1(new_n486), .B2(G148gat), .ZN(new_n496));
  INV_X1    g295(.A(G148gat), .ZN(new_n497));
  NAND3_X1  g296(.A1(new_n497), .A2(KEYINPUT78), .A3(G141gat), .ZN(new_n498));
  NAND3_X1  g297(.A1(new_n496), .A2(new_n487), .A3(new_n498), .ZN(new_n499));
  OAI21_X1  g298(.A(new_n493), .B1(new_n492), .B2(KEYINPUT2), .ZN(new_n500));
  AOI22_X1  g299(.A1(new_n490), .A2(new_n494), .B1(new_n499), .B2(new_n500), .ZN(new_n501));
  XOR2_X1   g300(.A(KEYINPUT79), .B(KEYINPUT3), .Z(new_n502));
  AOI21_X1  g301(.A(KEYINPUT29), .B1(new_n501), .B2(new_n502), .ZN(new_n503));
  OAI21_X1  g302(.A(KEYINPUT84), .B1(new_n484), .B2(new_n503), .ZN(new_n504));
  NAND2_X1  g303(.A1(new_n479), .A2(new_n481), .ZN(new_n505));
  INV_X1    g304(.A(KEYINPUT29), .ZN(new_n506));
  NAND4_X1  g305(.A1(new_n480), .A2(new_n475), .A3(new_n476), .A4(new_n478), .ZN(new_n507));
  NAND3_X1  g306(.A1(new_n505), .A2(new_n506), .A3(new_n507), .ZN(new_n508));
  NAND2_X1  g307(.A1(new_n508), .A2(new_n502), .ZN(new_n509));
  XNOR2_X1  g308(.A(G141gat), .B(G148gat), .ZN(new_n510));
  OAI211_X1 g309(.A(new_n493), .B(new_n492), .C1(new_n510), .C2(KEYINPUT2), .ZN(new_n511));
  NAND2_X1  g310(.A1(new_n499), .A2(new_n500), .ZN(new_n512));
  NAND2_X1  g311(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  NAND2_X1  g312(.A1(new_n509), .A2(new_n513), .ZN(new_n514));
  NAND2_X1  g313(.A1(new_n479), .A2(KEYINPUT74), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n515), .A2(new_n480), .ZN(new_n516));
  NAND3_X1  g315(.A1(new_n479), .A2(KEYINPUT74), .A3(new_n481), .ZN(new_n517));
  NAND2_X1  g316(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  INV_X1    g317(.A(KEYINPUT84), .ZN(new_n519));
  NAND3_X1  g318(.A1(new_n511), .A2(new_n512), .A3(new_n502), .ZN(new_n520));
  NAND2_X1  g319(.A1(new_n520), .A2(new_n506), .ZN(new_n521));
  NAND3_X1  g320(.A1(new_n518), .A2(new_n519), .A3(new_n521), .ZN(new_n522));
  NAND3_X1  g321(.A1(new_n504), .A2(new_n514), .A3(new_n522), .ZN(new_n523));
  NAND2_X1  g322(.A1(G228gat), .A2(G233gat), .ZN(new_n524));
  NAND2_X1  g323(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  NOR3_X1   g324(.A1(new_n482), .A2(new_n483), .A3(KEYINPUT29), .ZN(new_n526));
  OAI21_X1  g325(.A(new_n513), .B1(new_n526), .B2(KEYINPUT3), .ZN(new_n527));
  AOI22_X1  g326(.A1(new_n516), .A2(new_n517), .B1(new_n520), .B2(new_n506), .ZN(new_n528));
  INV_X1    g327(.A(new_n528), .ZN(new_n529));
  NAND4_X1  g328(.A1(new_n527), .A2(G228gat), .A3(G233gat), .A4(new_n529), .ZN(new_n530));
  AOI21_X1  g329(.A(new_n471), .B1(new_n525), .B2(new_n530), .ZN(new_n531));
  INV_X1    g330(.A(KEYINPUT85), .ZN(new_n532));
  AOI21_X1  g331(.A(new_n470), .B1(new_n531), .B2(new_n532), .ZN(new_n533));
  NAND3_X1  g332(.A1(new_n516), .A2(new_n506), .A3(new_n517), .ZN(new_n534));
  INV_X1    g333(.A(KEYINPUT3), .ZN(new_n535));
  AOI21_X1  g334(.A(new_n501), .B1(new_n534), .B2(new_n535), .ZN(new_n536));
  NOR3_X1   g335(.A1(new_n536), .A2(new_n524), .A3(new_n528), .ZN(new_n537));
  AOI21_X1  g336(.A(new_n537), .B1(new_n524), .B2(new_n523), .ZN(new_n538));
  OAI21_X1  g337(.A(KEYINPUT85), .B1(new_n538), .B2(new_n471), .ZN(new_n539));
  NAND3_X1  g338(.A1(new_n525), .A2(new_n530), .A3(new_n471), .ZN(new_n540));
  NAND2_X1  g339(.A1(new_n540), .A2(KEYINPUT86), .ZN(new_n541));
  INV_X1    g340(.A(KEYINPUT86), .ZN(new_n542));
  NAND3_X1  g341(.A1(new_n538), .A2(new_n542), .A3(new_n471), .ZN(new_n543));
  NAND4_X1  g342(.A1(new_n533), .A2(new_n539), .A3(new_n541), .A4(new_n543), .ZN(new_n544));
  INV_X1    g343(.A(new_n540), .ZN(new_n545));
  OAI21_X1  g344(.A(new_n470), .B1(new_n545), .B2(new_n531), .ZN(new_n546));
  NAND2_X1  g345(.A1(new_n544), .A2(new_n546), .ZN(new_n547));
  NAND2_X1  g346(.A1(new_n466), .A2(new_n547), .ZN(new_n548));
  INV_X1    g347(.A(KEYINPUT77), .ZN(new_n549));
  XNOR2_X1  g348(.A(G8gat), .B(G36gat), .ZN(new_n550));
  XNOR2_X1  g349(.A(new_n550), .B(KEYINPUT76), .ZN(new_n551));
  XNOR2_X1  g350(.A(new_n551), .B(new_n271), .ZN(new_n552));
  XNOR2_X1  g351(.A(new_n552), .B(new_n207), .ZN(new_n553));
  INV_X1    g352(.A(new_n553), .ZN(new_n554));
  NAND2_X1  g353(.A1(G226gat), .A2(G233gat), .ZN(new_n555));
  INV_X1    g354(.A(new_n555), .ZN(new_n556));
  NAND3_X1  g355(.A1(new_n429), .A2(new_n393), .A3(new_n413), .ZN(new_n557));
  AOI21_X1  g356(.A(new_n556), .B1(new_n557), .B2(new_n506), .ZN(new_n558));
  NOR3_X1   g357(.A1(new_n380), .A2(new_n381), .A3(KEYINPUT68), .ZN(new_n559));
  AOI21_X1  g358(.A(new_n386), .B1(new_n385), .B2(new_n387), .ZN(new_n560));
  OAI21_X1  g359(.A(new_n378), .B1(new_n559), .B2(new_n560), .ZN(new_n561));
  NAND2_X1  g360(.A1(new_n390), .A2(new_n391), .ZN(new_n562));
  NAND2_X1  g361(.A1(new_n562), .A2(new_n377), .ZN(new_n563));
  NAND2_X1  g362(.A1(new_n561), .A2(new_n563), .ZN(new_n564));
  AND2_X1   g363(.A1(new_n376), .A2(new_n366), .ZN(new_n565));
  NAND3_X1  g364(.A1(new_n397), .A2(new_n412), .A3(new_n399), .ZN(new_n566));
  AOI22_X1  g365(.A1(new_n404), .A2(new_n403), .B1(new_n406), .B2(new_n408), .ZN(new_n567));
  NOR2_X1   g366(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  AOI22_X1  g367(.A1(new_n564), .A2(new_n565), .B1(new_n568), .B2(new_n401), .ZN(new_n569));
  AOI21_X1  g368(.A(new_n555), .B1(new_n569), .B2(new_n429), .ZN(new_n570));
  OAI21_X1  g369(.A(new_n484), .B1(new_n558), .B2(new_n570), .ZN(new_n571));
  NAND2_X1  g370(.A1(new_n557), .A2(new_n556), .ZN(new_n572));
  AOI21_X1  g371(.A(KEYINPUT29), .B1(new_n569), .B2(new_n429), .ZN(new_n573));
  OAI211_X1 g372(.A(new_n572), .B(new_n518), .C1(new_n573), .C2(new_n556), .ZN(new_n574));
  NAND2_X1  g373(.A1(new_n571), .A2(new_n574), .ZN(new_n575));
  INV_X1    g374(.A(KEYINPUT75), .ZN(new_n576));
  NAND2_X1  g375(.A1(new_n575), .A2(new_n576), .ZN(new_n577));
  NAND3_X1  g376(.A1(new_n571), .A2(new_n574), .A3(KEYINPUT75), .ZN(new_n578));
  AOI21_X1  g377(.A(new_n554), .B1(new_n577), .B2(new_n578), .ZN(new_n579));
  NAND3_X1  g378(.A1(new_n575), .A2(KEYINPUT30), .A3(new_n554), .ZN(new_n580));
  INV_X1    g379(.A(new_n580), .ZN(new_n581));
  OAI21_X1  g380(.A(new_n549), .B1(new_n579), .B2(new_n581), .ZN(new_n582));
  XNOR2_X1  g381(.A(G1gat), .B(G29gat), .ZN(new_n583));
  XNOR2_X1  g382(.A(new_n583), .B(KEYINPUT0), .ZN(new_n584));
  XNOR2_X1  g383(.A(new_n584), .B(G57gat), .ZN(new_n585));
  XNOR2_X1  g384(.A(new_n585), .B(new_n206), .ZN(new_n586));
  INV_X1    g385(.A(new_n586), .ZN(new_n587));
  NAND2_X1  g386(.A1(G225gat), .A2(G233gat), .ZN(new_n588));
  XNOR2_X1  g387(.A(new_n588), .B(KEYINPUT80), .ZN(new_n589));
  NAND4_X1  g388(.A1(new_n358), .A2(new_n363), .A3(new_n512), .A4(new_n511), .ZN(new_n590));
  INV_X1    g389(.A(new_n590), .ZN(new_n591));
  AOI22_X1  g390(.A1(new_n363), .A2(new_n358), .B1(new_n511), .B2(new_n512), .ZN(new_n592));
  OAI21_X1  g391(.A(new_n589), .B1(new_n591), .B2(new_n592), .ZN(new_n593));
  NAND2_X1  g392(.A1(new_n593), .A2(KEYINPUT5), .ZN(new_n594));
  INV_X1    g393(.A(KEYINPUT82), .ZN(new_n595));
  XOR2_X1   g394(.A(KEYINPUT81), .B(KEYINPUT4), .Z(new_n596));
  AOI21_X1  g395(.A(new_n595), .B1(new_n590), .B2(new_n596), .ZN(new_n597));
  INV_X1    g396(.A(new_n597), .ZN(new_n598));
  NOR2_X1   g397(.A1(new_n590), .A2(KEYINPUT4), .ZN(new_n599));
  INV_X1    g398(.A(new_n599), .ZN(new_n600));
  NAND3_X1  g399(.A1(new_n590), .A2(new_n595), .A3(new_n596), .ZN(new_n601));
  NAND3_X1  g400(.A1(new_n598), .A2(new_n600), .A3(new_n601), .ZN(new_n602));
  OAI211_X1 g401(.A(new_n520), .B(new_n364), .C1(new_n501), .C2(new_n535), .ZN(new_n603));
  INV_X1    g402(.A(new_n589), .ZN(new_n604));
  NAND2_X1  g403(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  INV_X1    g404(.A(new_n605), .ZN(new_n606));
  AOI21_X1  g405(.A(new_n594), .B1(new_n602), .B2(new_n606), .ZN(new_n607));
  OR2_X1    g406(.A1(new_n591), .A2(KEYINPUT4), .ZN(new_n608));
  NAND2_X1  g407(.A1(new_n591), .A2(new_n596), .ZN(new_n609));
  NOR2_X1   g408(.A1(new_n589), .A2(KEYINPUT5), .ZN(new_n610));
  NAND4_X1  g409(.A1(new_n608), .A2(new_n603), .A3(new_n609), .A4(new_n610), .ZN(new_n611));
  INV_X1    g410(.A(new_n611), .ZN(new_n612));
  OAI21_X1  g411(.A(new_n587), .B1(new_n607), .B2(new_n612), .ZN(new_n613));
  INV_X1    g412(.A(KEYINPUT5), .ZN(new_n614));
  INV_X1    g413(.A(new_n592), .ZN(new_n615));
  NAND2_X1  g414(.A1(new_n615), .A2(new_n590), .ZN(new_n616));
  AOI21_X1  g415(.A(new_n614), .B1(new_n616), .B2(new_n589), .ZN(new_n617));
  AND3_X1   g416(.A1(new_n590), .A2(new_n595), .A3(new_n596), .ZN(new_n618));
  NOR3_X1   g417(.A1(new_n618), .A2(new_n597), .A3(new_n599), .ZN(new_n619));
  OAI21_X1  g418(.A(new_n617), .B1(new_n619), .B2(new_n605), .ZN(new_n620));
  NAND3_X1  g419(.A1(new_n620), .A2(new_n586), .A3(new_n611), .ZN(new_n621));
  INV_X1    g420(.A(KEYINPUT6), .ZN(new_n622));
  NAND3_X1  g421(.A1(new_n613), .A2(new_n621), .A3(new_n622), .ZN(new_n623));
  AOI21_X1  g422(.A(new_n586), .B1(new_n620), .B2(new_n611), .ZN(new_n624));
  NAND2_X1  g423(.A1(new_n624), .A2(KEYINPUT6), .ZN(new_n625));
  NAND2_X1  g424(.A1(new_n623), .A2(new_n625), .ZN(new_n626));
  AND3_X1   g425(.A1(new_n571), .A2(new_n574), .A3(KEYINPUT75), .ZN(new_n627));
  AOI21_X1  g426(.A(KEYINPUT75), .B1(new_n571), .B2(new_n574), .ZN(new_n628));
  OAI21_X1  g427(.A(new_n553), .B1(new_n627), .B2(new_n628), .ZN(new_n629));
  NAND3_X1  g428(.A1(new_n629), .A2(KEYINPUT77), .A3(new_n580), .ZN(new_n630));
  NAND2_X1  g429(.A1(new_n575), .A2(new_n554), .ZN(new_n631));
  INV_X1    g430(.A(KEYINPUT30), .ZN(new_n632));
  NAND2_X1  g431(.A1(new_n631), .A2(new_n632), .ZN(new_n633));
  NAND4_X1  g432(.A1(new_n582), .A2(new_n626), .A3(new_n630), .A4(new_n633), .ZN(new_n634));
  OR2_X1    g433(.A1(new_n548), .A2(new_n634), .ZN(new_n635));
  INV_X1    g434(.A(new_n547), .ZN(new_n636));
  NAND3_X1  g435(.A1(new_n629), .A2(new_n580), .A3(new_n633), .ZN(new_n637));
  NOR2_X1   g436(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  INV_X1    g437(.A(new_n462), .ZN(new_n639));
  NOR3_X1   g438(.A1(new_n639), .A2(new_n464), .A3(KEYINPUT35), .ZN(new_n640));
  NAND2_X1  g439(.A1(new_n626), .A2(KEYINPUT90), .ZN(new_n641));
  INV_X1    g440(.A(KEYINPUT90), .ZN(new_n642));
  NAND2_X1  g441(.A1(new_n625), .A2(new_n642), .ZN(new_n643));
  NAND2_X1  g442(.A1(new_n641), .A2(new_n643), .ZN(new_n644));
  NAND3_X1  g443(.A1(new_n638), .A2(new_n640), .A3(new_n644), .ZN(new_n645));
  INV_X1    g444(.A(KEYINPUT91), .ZN(new_n646));
  NAND2_X1  g445(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  NAND4_X1  g446(.A1(new_n638), .A2(new_n640), .A3(KEYINPUT91), .A4(new_n644), .ZN(new_n648));
  AOI22_X1  g447(.A1(new_n635), .A2(KEYINPUT35), .B1(new_n647), .B2(new_n648), .ZN(new_n649));
  INV_X1    g448(.A(new_n649), .ZN(new_n650));
  NAND2_X1  g449(.A1(new_n466), .A2(KEYINPUT36), .ZN(new_n651));
  NAND2_X1  g450(.A1(new_n651), .A2(KEYINPUT72), .ZN(new_n652));
  NOR2_X1   g451(.A1(new_n639), .A2(new_n464), .ZN(new_n653));
  NOR2_X1   g452(.A1(new_n653), .A2(KEYINPUT36), .ZN(new_n654));
  INV_X1    g453(.A(new_n654), .ZN(new_n655));
  INV_X1    g454(.A(KEYINPUT72), .ZN(new_n656));
  NAND3_X1  g455(.A1(new_n466), .A2(new_n656), .A3(KEYINPUT36), .ZN(new_n657));
  NAND3_X1  g456(.A1(new_n652), .A2(new_n655), .A3(new_n657), .ZN(new_n658));
  INV_X1    g457(.A(KEYINPUT37), .ZN(new_n659));
  NAND2_X1  g458(.A1(new_n575), .A2(new_n659), .ZN(new_n660));
  XOR2_X1   g459(.A(KEYINPUT89), .B(KEYINPUT38), .Z(new_n661));
  INV_X1    g460(.A(new_n661), .ZN(new_n662));
  NAND3_X1  g461(.A1(new_n571), .A2(new_n574), .A3(KEYINPUT37), .ZN(new_n663));
  NAND4_X1  g462(.A1(new_n660), .A2(new_n553), .A3(new_n662), .A4(new_n663), .ZN(new_n664));
  NAND3_X1  g463(.A1(new_n641), .A2(new_n643), .A3(new_n664), .ZN(new_n665));
  AOI21_X1  g464(.A(new_n659), .B1(new_n577), .B2(new_n578), .ZN(new_n666));
  NAND2_X1  g465(.A1(new_n660), .A2(new_n553), .ZN(new_n667));
  OAI21_X1  g466(.A(new_n661), .B1(new_n666), .B2(new_n667), .ZN(new_n668));
  NAND2_X1  g467(.A1(new_n668), .A2(new_n631), .ZN(new_n669));
  NOR2_X1   g468(.A1(new_n665), .A2(new_n669), .ZN(new_n670));
  OAI211_X1 g469(.A(new_n609), .B(new_n603), .C1(KEYINPUT4), .C2(new_n591), .ZN(new_n671));
  NAND2_X1  g470(.A1(new_n671), .A2(new_n589), .ZN(new_n672));
  NOR2_X1   g471(.A1(new_n616), .A2(new_n589), .ZN(new_n673));
  INV_X1    g472(.A(KEYINPUT88), .ZN(new_n674));
  NAND2_X1  g473(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  NAND2_X1  g474(.A1(new_n672), .A2(new_n675), .ZN(new_n676));
  OAI21_X1  g475(.A(KEYINPUT39), .B1(new_n673), .B2(new_n674), .ZN(new_n677));
  OAI221_X1 g476(.A(new_n586), .B1(KEYINPUT39), .B2(new_n672), .C1(new_n676), .C2(new_n677), .ZN(new_n678));
  INV_X1    g477(.A(KEYINPUT40), .ZN(new_n679));
  AOI21_X1  g478(.A(new_n624), .B1(new_n678), .B2(new_n679), .ZN(new_n680));
  OAI211_X1 g479(.A(new_n637), .B(new_n680), .C1(new_n679), .C2(new_n678), .ZN(new_n681));
  NAND2_X1  g480(.A1(new_n681), .A2(new_n547), .ZN(new_n682));
  OR2_X1    g481(.A1(new_n670), .A2(new_n682), .ZN(new_n683));
  AND3_X1   g482(.A1(new_n544), .A2(KEYINPUT87), .A3(new_n546), .ZN(new_n684));
  AOI21_X1  g483(.A(KEYINPUT87), .B1(new_n544), .B2(new_n546), .ZN(new_n685));
  OAI21_X1  g484(.A(new_n634), .B1(new_n684), .B2(new_n685), .ZN(new_n686));
  NAND3_X1  g485(.A1(new_n658), .A2(new_n683), .A3(new_n686), .ZN(new_n687));
  AOI21_X1  g486(.A(new_n345), .B1(new_n650), .B2(new_n687), .ZN(new_n688));
  XNOR2_X1  g487(.A(G169gat), .B(G197gat), .ZN(new_n689));
  XNOR2_X1  g488(.A(G113gat), .B(G141gat), .ZN(new_n690));
  XNOR2_X1  g489(.A(new_n689), .B(new_n690), .ZN(new_n691));
  XNOR2_X1  g490(.A(KEYINPUT92), .B(KEYINPUT11), .ZN(new_n692));
  XNOR2_X1  g491(.A(new_n691), .B(new_n692), .ZN(new_n693));
  XOR2_X1   g492(.A(new_n693), .B(KEYINPUT12), .Z(new_n694));
  INV_X1    g493(.A(new_n694), .ZN(new_n695));
  AOI21_X1  g494(.A(new_n310), .B1(new_n235), .B2(new_n236), .ZN(new_n696));
  AOI21_X1  g495(.A(new_n309), .B1(new_n232), .B2(new_n234), .ZN(new_n697));
  NOR2_X1   g496(.A1(new_n696), .A2(new_n697), .ZN(new_n698));
  NAND2_X1  g497(.A1(G229gat), .A2(G233gat), .ZN(new_n699));
  AOI21_X1  g498(.A(KEYINPUT18), .B1(new_n698), .B2(new_n699), .ZN(new_n700));
  INV_X1    g499(.A(KEYINPUT18), .ZN(new_n701));
  INV_X1    g500(.A(new_n699), .ZN(new_n702));
  NOR4_X1   g501(.A1(new_n696), .A2(new_n701), .A3(new_n697), .A4(new_n702), .ZN(new_n703));
  NOR2_X1   g502(.A1(new_n700), .A2(new_n703), .ZN(new_n704));
  XNOR2_X1  g503(.A(new_n699), .B(KEYINPUT13), .ZN(new_n705));
  NAND2_X1  g504(.A1(new_n240), .A2(new_n309), .ZN(new_n706));
  INV_X1    g505(.A(new_n697), .ZN(new_n707));
  AOI21_X1  g506(.A(new_n705), .B1(new_n706), .B2(new_n707), .ZN(new_n708));
  INV_X1    g507(.A(new_n708), .ZN(new_n709));
  AOI21_X1  g508(.A(new_n695), .B1(new_n704), .B2(new_n709), .ZN(new_n710));
  INV_X1    g509(.A(new_n710), .ZN(new_n711));
  NOR4_X1   g510(.A1(new_n700), .A2(new_n703), .A3(new_n694), .A4(new_n708), .ZN(new_n712));
  INV_X1    g511(.A(new_n712), .ZN(new_n713));
  NAND2_X1  g512(.A1(new_n711), .A2(new_n713), .ZN(new_n714));
  INV_X1    g513(.A(new_n714), .ZN(new_n715));
  INV_X1    g514(.A(G230gat), .ZN(new_n716));
  NOR2_X1   g515(.A1(new_n716), .A2(new_n433), .ZN(new_n717));
  OAI21_X1  g516(.A(new_n211), .B1(new_n299), .B2(new_n301), .ZN(new_n718));
  INV_X1    g517(.A(KEYINPUT10), .ZN(new_n719));
  NAND3_X1  g518(.A1(new_n292), .A2(new_n212), .A3(new_n298), .ZN(new_n720));
  NAND3_X1  g519(.A1(new_n718), .A2(new_n719), .A3(new_n720), .ZN(new_n721));
  NAND4_X1  g520(.A1(new_n314), .A2(KEYINPUT10), .A3(new_n212), .A4(new_n315), .ZN(new_n722));
  AOI21_X1  g521(.A(new_n717), .B1(new_n721), .B2(new_n722), .ZN(new_n723));
  INV_X1    g522(.A(new_n723), .ZN(new_n724));
  NAND2_X1  g523(.A1(new_n718), .A2(new_n720), .ZN(new_n725));
  NAND2_X1  g524(.A1(new_n725), .A2(new_n717), .ZN(new_n726));
  NAND2_X1  g525(.A1(new_n724), .A2(new_n726), .ZN(new_n727));
  XNOR2_X1  g526(.A(G120gat), .B(G148gat), .ZN(new_n728));
  XNOR2_X1  g527(.A(new_n728), .B(KEYINPUT106), .ZN(new_n729));
  XNOR2_X1  g528(.A(new_n729), .B(new_n395), .ZN(new_n730));
  INV_X1    g529(.A(G204gat), .ZN(new_n731));
  XNOR2_X1  g530(.A(new_n730), .B(new_n731), .ZN(new_n732));
  INV_X1    g531(.A(new_n732), .ZN(new_n733));
  NAND2_X1  g532(.A1(new_n727), .A2(new_n733), .ZN(new_n734));
  NAND3_X1  g533(.A1(new_n724), .A2(new_n726), .A3(new_n732), .ZN(new_n735));
  NAND2_X1  g534(.A1(new_n734), .A2(new_n735), .ZN(new_n736));
  NOR2_X1   g535(.A1(new_n715), .A2(new_n736), .ZN(new_n737));
  NAND2_X1  g536(.A1(new_n688), .A2(new_n737), .ZN(new_n738));
  INV_X1    g537(.A(new_n738), .ZN(new_n739));
  INV_X1    g538(.A(new_n626), .ZN(new_n740));
  NAND2_X1  g539(.A1(new_n739), .A2(new_n740), .ZN(new_n741));
  XNOR2_X1  g540(.A(new_n741), .B(G1gat), .ZN(G1324gat));
  INV_X1    g541(.A(new_n637), .ZN(new_n743));
  OAI21_X1  g542(.A(G8gat), .B1(new_n738), .B2(new_n743), .ZN(new_n744));
  NAND2_X1  g543(.A1(new_n744), .A2(KEYINPUT42), .ZN(new_n745));
  XNOR2_X1  g544(.A(KEYINPUT107), .B(G8gat), .ZN(new_n746));
  XNOR2_X1  g545(.A(new_n746), .B(new_n305), .ZN(new_n747));
  NAND3_X1  g546(.A1(new_n739), .A2(new_n637), .A3(new_n747), .ZN(new_n748));
  MUX2_X1   g547(.A(KEYINPUT42), .B(new_n745), .S(new_n748), .Z(G1325gat));
  AOI21_X1  g548(.A(new_n656), .B1(new_n466), .B2(KEYINPUT36), .ZN(new_n750));
  INV_X1    g549(.A(KEYINPUT36), .ZN(new_n751));
  AOI211_X1 g550(.A(KEYINPUT72), .B(new_n751), .C1(new_n463), .C2(new_n465), .ZN(new_n752));
  NOR3_X1   g551(.A1(new_n750), .A2(new_n752), .A3(new_n654), .ZN(new_n753));
  AND3_X1   g552(.A1(new_n739), .A2(G15gat), .A3(new_n753), .ZN(new_n754));
  AOI21_X1  g553(.A(G15gat), .B1(new_n739), .B2(new_n653), .ZN(new_n755));
  NOR2_X1   g554(.A1(new_n754), .A2(new_n755), .ZN(G1326gat));
  INV_X1    g555(.A(KEYINPUT87), .ZN(new_n757));
  NAND2_X1  g556(.A1(new_n547), .A2(new_n757), .ZN(new_n758));
  NAND3_X1  g557(.A1(new_n544), .A2(KEYINPUT87), .A3(new_n546), .ZN(new_n759));
  NAND2_X1  g558(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  INV_X1    g559(.A(new_n760), .ZN(new_n761));
  OAI21_X1  g560(.A(KEYINPUT108), .B1(new_n738), .B2(new_n761), .ZN(new_n762));
  INV_X1    g561(.A(new_n762), .ZN(new_n763));
  NOR3_X1   g562(.A1(new_n738), .A2(KEYINPUT108), .A3(new_n761), .ZN(new_n764));
  OAI21_X1  g563(.A(KEYINPUT43), .B1(new_n763), .B2(new_n764), .ZN(new_n765));
  INV_X1    g564(.A(new_n764), .ZN(new_n766));
  INV_X1    g565(.A(KEYINPUT43), .ZN(new_n767));
  NAND3_X1  g566(.A1(new_n766), .A2(new_n767), .A3(new_n762), .ZN(new_n768));
  NAND2_X1  g567(.A1(new_n765), .A2(new_n768), .ZN(new_n769));
  XNOR2_X1  g568(.A(new_n769), .B(G22gat), .ZN(G1327gat));
  NAND2_X1  g569(.A1(new_n264), .A2(new_n269), .ZN(new_n771));
  INV_X1    g570(.A(new_n771), .ZN(new_n772));
  AOI21_X1  g571(.A(new_n772), .B1(new_n650), .B2(new_n687), .ZN(new_n773));
  NOR2_X1   g572(.A1(new_n341), .A2(new_n344), .ZN(new_n774));
  AND2_X1   g573(.A1(new_n774), .A2(new_n737), .ZN(new_n775));
  NAND2_X1  g574(.A1(new_n773), .A2(new_n775), .ZN(new_n776));
  NOR3_X1   g575(.A1(new_n776), .A2(G29gat), .A3(new_n626), .ZN(new_n777));
  XOR2_X1   g576(.A(new_n777), .B(KEYINPUT45), .Z(new_n778));
  INV_X1    g577(.A(KEYINPUT44), .ZN(new_n779));
  INV_X1    g578(.A(KEYINPUT110), .ZN(new_n780));
  INV_X1    g579(.A(KEYINPUT109), .ZN(new_n781));
  AOI21_X1  g580(.A(new_n781), .B1(new_n760), .B2(new_n634), .ZN(new_n782));
  OAI211_X1 g581(.A(new_n781), .B(new_n634), .C1(new_n684), .C2(new_n685), .ZN(new_n783));
  INV_X1    g582(.A(new_n783), .ZN(new_n784));
  OAI21_X1  g583(.A(new_n683), .B1(new_n782), .B2(new_n784), .ZN(new_n785));
  OAI21_X1  g584(.A(new_n780), .B1(new_n753), .B2(new_n785), .ZN(new_n786));
  NOR2_X1   g585(.A1(new_n670), .A2(new_n682), .ZN(new_n787));
  NAND2_X1  g586(.A1(new_n686), .A2(KEYINPUT109), .ZN(new_n788));
  AOI21_X1  g587(.A(new_n787), .B1(new_n788), .B2(new_n783), .ZN(new_n789));
  NAND3_X1  g588(.A1(new_n658), .A2(new_n789), .A3(KEYINPUT110), .ZN(new_n790));
  AOI21_X1  g589(.A(new_n649), .B1(new_n786), .B2(new_n790), .ZN(new_n791));
  OAI21_X1  g590(.A(new_n779), .B1(new_n791), .B2(new_n772), .ZN(new_n792));
  NAND2_X1  g591(.A1(new_n773), .A2(KEYINPUT44), .ZN(new_n793));
  AND2_X1   g592(.A1(new_n792), .A2(new_n793), .ZN(new_n794));
  NAND2_X1  g593(.A1(new_n794), .A2(new_n775), .ZN(new_n795));
  OAI21_X1  g594(.A(G29gat), .B1(new_n795), .B2(new_n626), .ZN(new_n796));
  NAND2_X1  g595(.A1(new_n778), .A2(new_n796), .ZN(G1328gat));
  OAI21_X1  g596(.A(G36gat), .B1(new_n795), .B2(new_n743), .ZN(new_n798));
  NOR3_X1   g597(.A1(new_n776), .A2(G36gat), .A3(new_n743), .ZN(new_n799));
  XNOR2_X1  g598(.A(new_n799), .B(KEYINPUT46), .ZN(new_n800));
  NAND2_X1  g599(.A1(new_n798), .A2(new_n800), .ZN(G1329gat));
  OAI21_X1  g600(.A(G43gat), .B1(new_n795), .B2(new_n658), .ZN(new_n802));
  OR4_X1    g601(.A1(G43gat), .A2(new_n776), .A3(new_n464), .A4(new_n639), .ZN(new_n803));
  NAND2_X1  g602(.A1(new_n802), .A2(new_n803), .ZN(new_n804));
  INV_X1    g603(.A(KEYINPUT47), .ZN(new_n805));
  NAND2_X1  g604(.A1(new_n804), .A2(new_n805), .ZN(new_n806));
  NAND3_X1  g605(.A1(new_n802), .A2(KEYINPUT47), .A3(new_n803), .ZN(new_n807));
  NAND2_X1  g606(.A1(new_n806), .A2(new_n807), .ZN(G1330gat));
  OAI21_X1  g607(.A(G50gat), .B1(new_n795), .B2(new_n547), .ZN(new_n809));
  NOR3_X1   g608(.A1(new_n776), .A2(G50gat), .A3(new_n761), .ZN(new_n810));
  INV_X1    g609(.A(new_n810), .ZN(new_n811));
  NAND3_X1  g610(.A1(new_n809), .A2(KEYINPUT48), .A3(new_n811), .ZN(new_n812));
  NAND3_X1  g611(.A1(new_n794), .A2(new_n760), .A3(new_n775), .ZN(new_n813));
  AOI21_X1  g612(.A(new_n810), .B1(new_n813), .B2(G50gat), .ZN(new_n814));
  OAI21_X1  g613(.A(new_n812), .B1(new_n814), .B2(KEYINPUT48), .ZN(G1331gat));
  AND3_X1   g614(.A1(new_n658), .A2(KEYINPUT110), .A3(new_n789), .ZN(new_n816));
  AOI21_X1  g615(.A(KEYINPUT110), .B1(new_n658), .B2(new_n789), .ZN(new_n817));
  OAI21_X1  g616(.A(new_n650), .B1(new_n816), .B2(new_n817), .ZN(new_n818));
  NOR2_X1   g617(.A1(new_n345), .A2(new_n714), .ZN(new_n819));
  NAND3_X1  g618(.A1(new_n818), .A2(new_n736), .A3(new_n819), .ZN(new_n820));
  NAND2_X1  g619(.A1(new_n820), .A2(KEYINPUT111), .ZN(new_n821));
  INV_X1    g620(.A(KEYINPUT111), .ZN(new_n822));
  NAND4_X1  g621(.A1(new_n818), .A2(new_n822), .A3(new_n736), .A4(new_n819), .ZN(new_n823));
  NAND2_X1  g622(.A1(new_n821), .A2(new_n823), .ZN(new_n824));
  NOR2_X1   g623(.A1(new_n824), .A2(new_n626), .ZN(new_n825));
  XNOR2_X1  g624(.A(new_n825), .B(new_n270), .ZN(G1332gat));
  XNOR2_X1  g625(.A(new_n637), .B(KEYINPUT112), .ZN(new_n827));
  INV_X1    g626(.A(new_n827), .ZN(new_n828));
  NOR2_X1   g627(.A1(new_n824), .A2(new_n828), .ZN(new_n829));
  XNOR2_X1  g628(.A(KEYINPUT49), .B(G64gat), .ZN(new_n830));
  NAND2_X1  g629(.A1(new_n829), .A2(new_n830), .ZN(new_n831));
  NOR2_X1   g630(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n832));
  OAI21_X1  g631(.A(new_n831), .B1(new_n829), .B2(new_n832), .ZN(G1333gat));
  INV_X1    g632(.A(KEYINPUT50), .ZN(new_n834));
  NAND3_X1  g633(.A1(new_n821), .A2(new_n653), .A3(new_n823), .ZN(new_n835));
  INV_X1    g634(.A(G71gat), .ZN(new_n836));
  NAND2_X1  g635(.A1(new_n835), .A2(new_n836), .ZN(new_n837));
  INV_X1    g636(.A(KEYINPUT113), .ZN(new_n838));
  NAND4_X1  g637(.A1(new_n821), .A2(G71gat), .A3(new_n753), .A4(new_n823), .ZN(new_n839));
  AND3_X1   g638(.A1(new_n837), .A2(new_n838), .A3(new_n839), .ZN(new_n840));
  AOI21_X1  g639(.A(new_n838), .B1(new_n837), .B2(new_n839), .ZN(new_n841));
  OAI21_X1  g640(.A(new_n834), .B1(new_n840), .B2(new_n841), .ZN(new_n842));
  NAND2_X1  g641(.A1(new_n837), .A2(new_n839), .ZN(new_n843));
  NAND2_X1  g642(.A1(new_n843), .A2(KEYINPUT113), .ZN(new_n844));
  NAND3_X1  g643(.A1(new_n837), .A2(new_n838), .A3(new_n839), .ZN(new_n845));
  NAND3_X1  g644(.A1(new_n844), .A2(KEYINPUT50), .A3(new_n845), .ZN(new_n846));
  NAND2_X1  g645(.A1(new_n842), .A2(new_n846), .ZN(G1334gat));
  NOR2_X1   g646(.A1(new_n824), .A2(new_n761), .ZN(new_n848));
  XOR2_X1   g647(.A(new_n848), .B(G78gat), .Z(G1335gat));
  NAND2_X1  g648(.A1(new_n774), .A2(new_n715), .ZN(new_n850));
  INV_X1    g649(.A(new_n736), .ZN(new_n851));
  NOR2_X1   g650(.A1(new_n850), .A2(new_n851), .ZN(new_n852));
  NAND2_X1  g651(.A1(new_n794), .A2(new_n852), .ZN(new_n853));
  OAI21_X1  g652(.A(G85gat), .B1(new_n853), .B2(new_n626), .ZN(new_n854));
  NAND2_X1  g653(.A1(new_n786), .A2(new_n790), .ZN(new_n855));
  AOI21_X1  g654(.A(new_n772), .B1(new_n855), .B2(new_n650), .ZN(new_n856));
  INV_X1    g655(.A(new_n850), .ZN(new_n857));
  AOI21_X1  g656(.A(KEYINPUT51), .B1(new_n856), .B2(new_n857), .ZN(new_n858));
  INV_X1    g657(.A(KEYINPUT51), .ZN(new_n859));
  NOR4_X1   g658(.A1(new_n791), .A2(new_n859), .A3(new_n772), .A4(new_n850), .ZN(new_n860));
  OAI21_X1  g659(.A(KEYINPUT114), .B1(new_n858), .B2(new_n860), .ZN(new_n861));
  NAND3_X1  g660(.A1(new_n818), .A2(new_n771), .A3(new_n857), .ZN(new_n862));
  NAND2_X1  g661(.A1(new_n862), .A2(new_n859), .ZN(new_n863));
  INV_X1    g662(.A(KEYINPUT114), .ZN(new_n864));
  NAND2_X1  g663(.A1(new_n863), .A2(new_n864), .ZN(new_n865));
  NAND2_X1  g664(.A1(new_n861), .A2(new_n865), .ZN(new_n866));
  NAND3_X1  g665(.A1(new_n866), .A2(new_n206), .A3(new_n736), .ZN(new_n867));
  OAI21_X1  g666(.A(new_n854), .B1(new_n867), .B2(new_n626), .ZN(G1336gat));
  NAND3_X1  g667(.A1(new_n736), .A2(new_n827), .A3(new_n207), .ZN(new_n869));
  AOI21_X1  g668(.A(new_n869), .B1(new_n861), .B2(new_n865), .ZN(new_n870));
  NAND4_X1  g669(.A1(new_n792), .A2(new_n793), .A3(new_n827), .A4(new_n852), .ZN(new_n871));
  NAND2_X1  g670(.A1(new_n871), .A2(G92gat), .ZN(new_n872));
  INV_X1    g671(.A(KEYINPUT52), .ZN(new_n873));
  NAND2_X1  g672(.A1(new_n872), .A2(new_n873), .ZN(new_n874));
  NAND3_X1  g673(.A1(new_n856), .A2(KEYINPUT51), .A3(new_n857), .ZN(new_n875));
  NAND2_X1  g674(.A1(new_n863), .A2(new_n875), .ZN(new_n876));
  XNOR2_X1  g675(.A(new_n869), .B(KEYINPUT115), .ZN(new_n877));
  NAND4_X1  g676(.A1(new_n792), .A2(new_n793), .A3(new_n637), .A4(new_n852), .ZN(new_n878));
  AOI22_X1  g677(.A1(new_n876), .A2(new_n877), .B1(new_n878), .B2(G92gat), .ZN(new_n879));
  OAI22_X1  g678(.A1(new_n870), .A2(new_n874), .B1(new_n879), .B2(new_n873), .ZN(new_n880));
  NAND2_X1  g679(.A1(new_n880), .A2(KEYINPUT116), .ZN(new_n881));
  INV_X1    g680(.A(KEYINPUT116), .ZN(new_n882));
  OAI221_X1 g681(.A(new_n882), .B1(new_n879), .B2(new_n873), .C1(new_n870), .C2(new_n874), .ZN(new_n883));
  NAND2_X1  g682(.A1(new_n881), .A2(new_n883), .ZN(G1337gat));
  NOR2_X1   g683(.A1(new_n851), .A2(G99gat), .ZN(new_n885));
  NAND3_X1  g684(.A1(new_n866), .A2(new_n653), .A3(new_n885), .ZN(new_n886));
  OAI21_X1  g685(.A(G99gat), .B1(new_n853), .B2(new_n658), .ZN(new_n887));
  NAND2_X1  g686(.A1(new_n886), .A2(new_n887), .ZN(G1338gat));
  NOR2_X1   g687(.A1(new_n853), .A2(new_n761), .ZN(new_n889));
  INV_X1    g688(.A(G106gat), .ZN(new_n890));
  NOR2_X1   g689(.A1(new_n889), .A2(new_n890), .ZN(new_n891));
  NAND3_X1  g690(.A1(new_n736), .A2(new_n890), .A3(new_n636), .ZN(new_n892));
  XNOR2_X1  g691(.A(new_n892), .B(KEYINPUT117), .ZN(new_n893));
  AOI21_X1  g692(.A(new_n893), .B1(new_n863), .B2(new_n875), .ZN(new_n894));
  OAI21_X1  g693(.A(KEYINPUT53), .B1(new_n891), .B2(new_n894), .ZN(new_n895));
  OAI21_X1  g694(.A(G106gat), .B1(new_n853), .B2(new_n547), .ZN(new_n896));
  INV_X1    g695(.A(KEYINPUT53), .ZN(new_n897));
  INV_X1    g696(.A(new_n866), .ZN(new_n898));
  OAI211_X1 g697(.A(new_n896), .B(new_n897), .C1(new_n898), .C2(new_n892), .ZN(new_n899));
  NAND2_X1  g698(.A1(new_n895), .A2(new_n899), .ZN(G1339gat));
  OR2_X1    g699(.A1(new_n341), .A2(new_n344), .ZN(new_n901));
  NOR2_X1   g700(.A1(new_n698), .A2(new_n699), .ZN(new_n902));
  AND3_X1   g701(.A1(new_n706), .A2(new_n707), .A3(new_n705), .ZN(new_n903));
  OAI21_X1  g702(.A(new_n693), .B1(new_n902), .B2(new_n903), .ZN(new_n904));
  AND2_X1   g703(.A1(new_n713), .A2(new_n904), .ZN(new_n905));
  INV_X1    g704(.A(KEYINPUT54), .ZN(new_n906));
  AOI21_X1  g705(.A(new_n732), .B1(new_n723), .B2(new_n906), .ZN(new_n907));
  NAND3_X1  g706(.A1(new_n721), .A2(new_n717), .A3(new_n722), .ZN(new_n908));
  NAND2_X1  g707(.A1(new_n908), .A2(KEYINPUT54), .ZN(new_n909));
  OAI21_X1  g708(.A(new_n907), .B1(new_n723), .B2(new_n909), .ZN(new_n910));
  INV_X1    g709(.A(KEYINPUT55), .ZN(new_n911));
  OAI21_X1  g710(.A(new_n735), .B1(new_n910), .B2(new_n911), .ZN(new_n912));
  AOI21_X1  g711(.A(new_n912), .B1(new_n911), .B2(new_n910), .ZN(new_n913));
  NAND3_X1  g712(.A1(new_n771), .A2(new_n905), .A3(new_n913), .ZN(new_n914));
  NAND3_X1  g713(.A1(new_n713), .A2(new_n736), .A3(new_n904), .ZN(new_n915));
  NAND2_X1  g714(.A1(new_n910), .A2(new_n911), .ZN(new_n916));
  OAI21_X1  g715(.A(new_n916), .B1(new_n710), .B2(new_n712), .ZN(new_n917));
  OAI21_X1  g716(.A(new_n915), .B1(new_n917), .B2(new_n912), .ZN(new_n918));
  NAND3_X1  g717(.A1(new_n918), .A2(new_n264), .A3(new_n269), .ZN(new_n919));
  AOI21_X1  g718(.A(new_n901), .B1(new_n914), .B2(new_n919), .ZN(new_n920));
  NOR3_X1   g719(.A1(new_n345), .A2(new_n714), .A3(new_n736), .ZN(new_n921));
  NOR2_X1   g720(.A1(new_n920), .A2(new_n921), .ZN(new_n922));
  NOR2_X1   g721(.A1(new_n922), .A2(new_n626), .ZN(new_n923));
  NAND2_X1  g722(.A1(new_n923), .A2(new_n828), .ZN(new_n924));
  NAND2_X1  g723(.A1(new_n761), .A2(new_n653), .ZN(new_n925));
  NOR2_X1   g724(.A1(new_n924), .A2(new_n925), .ZN(new_n926));
  INV_X1    g725(.A(new_n926), .ZN(new_n927));
  OAI21_X1  g726(.A(G113gat), .B1(new_n927), .B2(new_n715), .ZN(new_n928));
  NOR2_X1   g727(.A1(new_n924), .A2(new_n548), .ZN(new_n929));
  NAND2_X1  g728(.A1(new_n714), .A2(new_n352), .ZN(new_n930));
  XOR2_X1   g729(.A(new_n930), .B(KEYINPUT118), .Z(new_n931));
  NAND2_X1  g730(.A1(new_n929), .A2(new_n931), .ZN(new_n932));
  NAND2_X1  g731(.A1(new_n928), .A2(new_n932), .ZN(G1340gat));
  OAI21_X1  g732(.A(G120gat), .B1(new_n927), .B2(new_n851), .ZN(new_n934));
  NAND3_X1  g733(.A1(new_n929), .A2(new_n354), .A3(new_n736), .ZN(new_n935));
  NAND2_X1  g734(.A1(new_n934), .A2(new_n935), .ZN(G1341gat));
  AOI21_X1  g735(.A(G127gat), .B1(new_n929), .B2(new_n901), .ZN(new_n937));
  NOR2_X1   g736(.A1(new_n774), .A2(new_n346), .ZN(new_n938));
  AOI21_X1  g737(.A(new_n937), .B1(new_n926), .B2(new_n938), .ZN(G1342gat));
  INV_X1    g738(.A(new_n548), .ZN(new_n940));
  NAND2_X1  g739(.A1(new_n771), .A2(new_n743), .ZN(new_n941));
  XNOR2_X1  g740(.A(new_n941), .B(KEYINPUT119), .ZN(new_n942));
  INV_X1    g741(.A(new_n942), .ZN(new_n943));
  NAND4_X1  g742(.A1(new_n923), .A2(new_n347), .A3(new_n940), .A4(new_n943), .ZN(new_n944));
  XOR2_X1   g743(.A(new_n944), .B(KEYINPUT56), .Z(new_n945));
  OAI21_X1  g744(.A(G134gat), .B1(new_n927), .B2(new_n772), .ZN(new_n946));
  NAND2_X1  g745(.A1(new_n945), .A2(new_n946), .ZN(G1343gat));
  NOR2_X1   g746(.A1(new_n922), .A2(new_n547), .ZN(new_n948));
  NAND2_X1  g747(.A1(new_n658), .A2(new_n740), .ZN(new_n949));
  NOR2_X1   g748(.A1(new_n949), .A2(new_n827), .ZN(new_n950));
  NAND2_X1  g749(.A1(new_n948), .A2(new_n950), .ZN(new_n951));
  INV_X1    g750(.A(new_n951), .ZN(new_n952));
  NAND3_X1  g751(.A1(new_n952), .A2(new_n486), .A3(new_n714), .ZN(new_n953));
  INV_X1    g752(.A(KEYINPUT120), .ZN(new_n954));
  NAND3_X1  g753(.A1(new_n772), .A2(new_n954), .A3(new_n918), .ZN(new_n955));
  NAND2_X1  g754(.A1(new_n919), .A2(KEYINPUT120), .ZN(new_n956));
  NAND3_X1  g755(.A1(new_n955), .A2(new_n956), .A3(new_n914), .ZN(new_n957));
  AOI21_X1  g756(.A(new_n921), .B1(new_n957), .B2(new_n774), .ZN(new_n958));
  OAI21_X1  g757(.A(KEYINPUT57), .B1(new_n958), .B2(new_n761), .ZN(new_n959));
  OR3_X1    g758(.A1(new_n922), .A2(KEYINPUT57), .A3(new_n547), .ZN(new_n960));
  NAND3_X1  g759(.A1(new_n959), .A2(new_n960), .A3(new_n950), .ZN(new_n961));
  NOR2_X1   g760(.A1(new_n961), .A2(new_n715), .ZN(new_n962));
  OAI21_X1  g761(.A(new_n953), .B1(new_n962), .B2(new_n486), .ZN(new_n963));
  NAND2_X1  g762(.A1(new_n963), .A2(KEYINPUT58), .ZN(new_n964));
  INV_X1    g763(.A(KEYINPUT58), .ZN(new_n965));
  OAI211_X1 g764(.A(new_n965), .B(new_n953), .C1(new_n962), .C2(new_n486), .ZN(new_n966));
  NAND2_X1  g765(.A1(new_n964), .A2(new_n966), .ZN(G1344gat));
  NAND3_X1  g766(.A1(new_n952), .A2(new_n497), .A3(new_n736), .ZN(new_n968));
  INV_X1    g767(.A(KEYINPUT59), .ZN(new_n969));
  OAI21_X1  g768(.A(new_n969), .B1(new_n961), .B2(new_n851), .ZN(new_n970));
  NOR2_X1   g769(.A1(new_n970), .A2(new_n497), .ZN(new_n971));
  INV_X1    g770(.A(new_n948), .ZN(new_n972));
  NAND2_X1  g771(.A1(new_n972), .A2(KEYINPUT57), .ZN(new_n973));
  OR3_X1    g772(.A1(new_n922), .A2(KEYINPUT57), .A3(new_n761), .ZN(new_n974));
  NAND4_X1  g773(.A1(new_n973), .A2(new_n736), .A3(new_n974), .A4(new_n950), .ZN(new_n975));
  AOI21_X1  g774(.A(new_n969), .B1(new_n975), .B2(G148gat), .ZN(new_n976));
  OAI21_X1  g775(.A(new_n968), .B1(new_n971), .B2(new_n976), .ZN(G1345gat));
  NOR3_X1   g776(.A1(new_n961), .A2(new_n491), .A3(new_n774), .ZN(new_n978));
  AOI21_X1  g777(.A(G155gat), .B1(new_n952), .B2(new_n901), .ZN(new_n979));
  NOR2_X1   g778(.A1(new_n978), .A2(new_n979), .ZN(G1346gat));
  OR4_X1    g779(.A1(G162gat), .A2(new_n972), .A3(new_n942), .A4(new_n949), .ZN(new_n981));
  NOR2_X1   g780(.A1(new_n961), .A2(new_n772), .ZN(new_n982));
  OAI21_X1  g781(.A(new_n981), .B1(new_n982), .B2(new_n261), .ZN(new_n983));
  NAND2_X1  g782(.A1(new_n983), .A2(KEYINPUT121), .ZN(new_n984));
  INV_X1    g783(.A(KEYINPUT121), .ZN(new_n985));
  OAI211_X1 g784(.A(new_n981), .B(new_n985), .C1(new_n982), .C2(new_n261), .ZN(new_n986));
  NAND2_X1  g785(.A1(new_n984), .A2(new_n986), .ZN(G1347gat));
  NOR2_X1   g786(.A1(new_n922), .A2(new_n925), .ZN(new_n988));
  NOR2_X1   g787(.A1(new_n743), .A2(new_n740), .ZN(new_n989));
  NAND2_X1  g788(.A1(new_n988), .A2(new_n989), .ZN(new_n990));
  OAI21_X1  g789(.A(G169gat), .B1(new_n990), .B2(new_n715), .ZN(new_n991));
  OAI21_X1  g790(.A(new_n626), .B1(new_n920), .B2(new_n921), .ZN(new_n992));
  NAND2_X1  g791(.A1(new_n992), .A2(KEYINPUT122), .ZN(new_n993));
  INV_X1    g792(.A(KEYINPUT122), .ZN(new_n994));
  OAI211_X1 g793(.A(new_n994), .B(new_n626), .C1(new_n920), .C2(new_n921), .ZN(new_n995));
  NAND4_X1  g794(.A1(new_n993), .A2(new_n940), .A3(new_n827), .A4(new_n995), .ZN(new_n996));
  NAND2_X1  g795(.A1(new_n714), .A2(new_n394), .ZN(new_n997));
  OAI21_X1  g796(.A(new_n991), .B1(new_n996), .B2(new_n997), .ZN(G1348gat));
  NOR3_X1   g797(.A1(new_n990), .A2(new_n395), .A3(new_n851), .ZN(new_n999));
  INV_X1    g798(.A(new_n996), .ZN(new_n1000));
  NAND2_X1  g799(.A1(new_n1000), .A2(new_n736), .ZN(new_n1001));
  AOI21_X1  g800(.A(new_n999), .B1(new_n1001), .B2(new_n395), .ZN(G1349gat));
  INV_X1    g801(.A(KEYINPUT124), .ZN(new_n1003));
  OAI21_X1  g802(.A(new_n1003), .B1(new_n990), .B2(new_n774), .ZN(new_n1004));
  NAND4_X1  g803(.A1(new_n988), .A2(KEYINPUT124), .A3(new_n901), .A4(new_n989), .ZN(new_n1005));
  NAND3_X1  g804(.A1(new_n1004), .A2(new_n1005), .A3(G183gat), .ZN(new_n1006));
  INV_X1    g805(.A(KEYINPUT123), .ZN(new_n1007));
  AOI21_X1  g806(.A(new_n774), .B1(new_n382), .B2(new_n388), .ZN(new_n1008));
  AOI21_X1  g807(.A(new_n1007), .B1(new_n1000), .B2(new_n1008), .ZN(new_n1009));
  INV_X1    g808(.A(new_n1008), .ZN(new_n1010));
  NOR3_X1   g809(.A1(new_n996), .A2(KEYINPUT123), .A3(new_n1010), .ZN(new_n1011));
  OAI21_X1  g810(.A(new_n1006), .B1(new_n1009), .B2(new_n1011), .ZN(new_n1012));
  NAND2_X1  g811(.A1(new_n1012), .A2(KEYINPUT60), .ZN(new_n1013));
  INV_X1    g812(.A(KEYINPUT60), .ZN(new_n1014));
  OAI211_X1 g813(.A(new_n1014), .B(new_n1006), .C1(new_n1009), .C2(new_n1011), .ZN(new_n1015));
  NAND2_X1  g814(.A1(new_n1013), .A2(new_n1015), .ZN(G1350gat));
  NAND3_X1  g815(.A1(new_n1000), .A2(new_n391), .A3(new_n771), .ZN(new_n1017));
  OAI21_X1  g816(.A(G190gat), .B1(new_n990), .B2(new_n772), .ZN(new_n1018));
  NAND2_X1  g817(.A1(new_n1018), .A2(KEYINPUT125), .ZN(new_n1019));
  INV_X1    g818(.A(KEYINPUT61), .ZN(new_n1020));
  INV_X1    g819(.A(KEYINPUT125), .ZN(new_n1021));
  OAI211_X1 g820(.A(new_n1021), .B(G190gat), .C1(new_n990), .C2(new_n772), .ZN(new_n1022));
  AND3_X1   g821(.A1(new_n1019), .A2(new_n1020), .A3(new_n1022), .ZN(new_n1023));
  AOI21_X1  g822(.A(new_n1020), .B1(new_n1019), .B2(new_n1022), .ZN(new_n1024));
  OAI21_X1  g823(.A(new_n1017), .B1(new_n1023), .B2(new_n1024), .ZN(G1351gat));
  AND2_X1   g824(.A1(new_n973), .A2(new_n974), .ZN(new_n1026));
  AND2_X1   g825(.A1(new_n658), .A2(new_n989), .ZN(new_n1027));
  NAND2_X1  g826(.A1(new_n1026), .A2(new_n1027), .ZN(new_n1028));
  OAI21_X1  g827(.A(G197gat), .B1(new_n1028), .B2(new_n715), .ZN(new_n1029));
  AND4_X1   g828(.A1(new_n636), .A2(new_n993), .A3(new_n827), .A4(new_n995), .ZN(new_n1030));
  AND2_X1   g829(.A1(new_n1030), .A2(new_n658), .ZN(new_n1031));
  INV_X1    g830(.A(G197gat), .ZN(new_n1032));
  NAND3_X1  g831(.A1(new_n1031), .A2(new_n1032), .A3(new_n714), .ZN(new_n1033));
  NAND2_X1  g832(.A1(new_n1029), .A2(new_n1033), .ZN(G1352gat));
  NAND4_X1  g833(.A1(new_n1030), .A2(new_n731), .A3(new_n736), .A4(new_n658), .ZN(new_n1035));
  OR2_X1    g834(.A1(new_n1035), .A2(KEYINPUT62), .ZN(new_n1036));
  NAND2_X1  g835(.A1(new_n1035), .A2(KEYINPUT62), .ZN(new_n1037));
  AND3_X1   g836(.A1(new_n1026), .A2(new_n736), .A3(new_n1027), .ZN(new_n1038));
  OAI211_X1 g837(.A(new_n1036), .B(new_n1037), .C1(new_n731), .C2(new_n1038), .ZN(G1353gat));
  NAND4_X1  g838(.A1(new_n973), .A2(new_n901), .A3(new_n974), .A4(new_n1027), .ZN(new_n1040));
  NAND2_X1  g839(.A1(new_n1040), .A2(G211gat), .ZN(new_n1041));
  NAND3_X1  g840(.A1(new_n1041), .A2(KEYINPUT126), .A3(KEYINPUT63), .ZN(new_n1042));
  INV_X1    g841(.A(G211gat), .ZN(new_n1043));
  NAND3_X1  g842(.A1(new_n1031), .A2(new_n1043), .A3(new_n901), .ZN(new_n1044));
  OR2_X1    g843(.A1(KEYINPUT126), .A2(KEYINPUT63), .ZN(new_n1045));
  NAND2_X1  g844(.A1(KEYINPUT126), .A2(KEYINPUT63), .ZN(new_n1046));
  NAND4_X1  g845(.A1(new_n1040), .A2(G211gat), .A3(new_n1045), .A4(new_n1046), .ZN(new_n1047));
  NAND3_X1  g846(.A1(new_n1042), .A2(new_n1044), .A3(new_n1047), .ZN(G1354gat));
  AOI21_X1  g847(.A(G218gat), .B1(new_n1031), .B2(new_n771), .ZN(new_n1049));
  INV_X1    g848(.A(new_n1028), .ZN(new_n1050));
  NAND2_X1  g849(.A1(new_n771), .A2(G218gat), .ZN(new_n1051));
  XNOR2_X1  g850(.A(new_n1051), .B(KEYINPUT127), .ZN(new_n1052));
  AOI21_X1  g851(.A(new_n1049), .B1(new_n1050), .B2(new_n1052), .ZN(G1355gat));
endmodule


