//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 1 0 0 1 0 1 1 1 0 0 1 0 1 1 1 1 1 1 0 1 0 1 0 1 0 0 0 0 1 1 0 1 1 1 0 0 1 1 0 1 1 1 1 1 1 1 1 0 0 1 0 0 1 1 0 0 0 0 0 1 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:40:00 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1233, new_n1234, new_n1235, new_n1237,
    new_n1238, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1296, new_n1297, new_n1298, new_n1299,
    new_n1300, new_n1301;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0005(.A(G250), .ZN(new_n206));
  NAND2_X1  g0006(.A1(G1), .A2(G20), .ZN(new_n207));
  NOR2_X1   g0007(.A1(new_n207), .A2(G13), .ZN(new_n208));
  INV_X1    g0008(.A(new_n208), .ZN(new_n209));
  INV_X1    g0009(.A(G257), .ZN(new_n210));
  INV_X1    g0010(.A(G264), .ZN(new_n211));
  AOI211_X1 g0011(.A(new_n206), .B(new_n209), .C1(new_n210), .C2(new_n211), .ZN(new_n212));
  NAND2_X1  g0012(.A1(G1), .A2(G13), .ZN(new_n213));
  INV_X1    g0013(.A(G20), .ZN(new_n214));
  NOR2_X1   g0014(.A1(new_n213), .A2(new_n214), .ZN(new_n215));
  INV_X1    g0015(.A(new_n215), .ZN(new_n216));
  OAI21_X1  g0016(.A(G50), .B1(G58), .B2(G68), .ZN(new_n217));
  OAI22_X1  g0017(.A1(new_n212), .A2(KEYINPUT0), .B1(new_n216), .B2(new_n217), .ZN(new_n218));
  AOI22_X1  g0018(.A1(G77), .A2(G244), .B1(G97), .B2(G257), .ZN(new_n219));
  INV_X1    g0019(.A(G226), .ZN(new_n220));
  INV_X1    g0020(.A(G87), .ZN(new_n221));
  OAI221_X1 g0021(.A(new_n219), .B1(new_n202), .B2(new_n220), .C1(new_n221), .C2(new_n206), .ZN(new_n222));
  AOI22_X1  g0022(.A1(G107), .A2(G264), .B1(G116), .B2(G270), .ZN(new_n223));
  INV_X1    g0023(.A(G58), .ZN(new_n224));
  INV_X1    g0024(.A(G232), .ZN(new_n225));
  INV_X1    g0025(.A(G68), .ZN(new_n226));
  INV_X1    g0026(.A(G238), .ZN(new_n227));
  OAI221_X1 g0027(.A(new_n223), .B1(new_n224), .B2(new_n225), .C1(new_n226), .C2(new_n227), .ZN(new_n228));
  OAI21_X1  g0028(.A(new_n207), .B1(new_n222), .B2(new_n228), .ZN(new_n229));
  XNOR2_X1  g0029(.A(new_n229), .B(KEYINPUT1), .ZN(new_n230));
  AOI211_X1 g0030(.A(new_n218), .B(new_n230), .C1(KEYINPUT0), .C2(new_n212), .ZN(G361));
  XNOR2_X1  g0031(.A(G238), .B(G244), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n232), .B(G232), .ZN(new_n233));
  XNOR2_X1  g0033(.A(KEYINPUT2), .B(G226), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n233), .B(new_n234), .ZN(new_n235));
  XOR2_X1   g0035(.A(G250), .B(G257), .Z(new_n236));
  XNOR2_X1  g0036(.A(G264), .B(G270), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n235), .B(new_n238), .ZN(G358));
  XNOR2_X1  g0039(.A(G87), .B(G97), .ZN(new_n240));
  INV_X1    g0040(.A(G116), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XNOR2_X1  g0042(.A(KEYINPUT64), .B(G107), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XOR2_X1   g0044(.A(G50), .B(G68), .Z(new_n245));
  XNOR2_X1  g0045(.A(G58), .B(G77), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n245), .B(new_n246), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n244), .B(new_n247), .ZN(G351));
  NAND2_X1  g0048(.A1(new_n203), .A2(G20), .ZN(new_n249));
  INV_X1    g0049(.A(G33), .ZN(new_n250));
  NAND2_X1  g0050(.A1(new_n214), .A2(new_n250), .ZN(new_n251));
  INV_X1    g0051(.A(new_n251), .ZN(new_n252));
  AOI22_X1  g0052(.A1(new_n249), .A2(KEYINPUT68), .B1(G150), .B2(new_n252), .ZN(new_n253));
  INV_X1    g0053(.A(KEYINPUT8), .ZN(new_n254));
  NAND2_X1  g0054(.A1(new_n254), .A2(G58), .ZN(new_n255));
  OR2_X1    g0055(.A1(new_n255), .A2(KEYINPUT67), .ZN(new_n256));
  NOR2_X1   g0056(.A1(new_n254), .A2(G58), .ZN(new_n257));
  OAI21_X1  g0057(.A(new_n255), .B1(new_n257), .B2(KEYINPUT67), .ZN(new_n258));
  AND2_X1   g0058(.A1(new_n256), .A2(new_n258), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n214), .A2(G33), .ZN(new_n260));
  OAI221_X1 g0060(.A(new_n253), .B1(KEYINPUT68), .B2(new_n249), .C1(new_n259), .C2(new_n260), .ZN(new_n261));
  NAND3_X1  g0061(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n262));
  NAND2_X1  g0062(.A1(new_n262), .A2(new_n213), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n261), .A2(new_n263), .ZN(new_n264));
  INV_X1    g0064(.A(G1), .ZN(new_n265));
  NAND3_X1  g0065(.A1(new_n265), .A2(G13), .A3(G20), .ZN(new_n266));
  AND2_X1   g0066(.A1(new_n262), .A2(new_n213), .ZN(new_n267));
  OAI21_X1  g0067(.A(new_n267), .B1(G1), .B2(new_n214), .ZN(new_n268));
  MUX2_X1   g0068(.A(new_n266), .B(new_n268), .S(G50), .Z(new_n269));
  NAND2_X1  g0069(.A1(new_n264), .A2(new_n269), .ZN(new_n270));
  AOI21_X1  g0070(.A(new_n270), .B1(KEYINPUT72), .B2(KEYINPUT9), .ZN(new_n271));
  NAND2_X1  g0071(.A1(KEYINPUT72), .A2(KEYINPUT9), .ZN(new_n272));
  AOI21_X1  g0072(.A(new_n272), .B1(new_n264), .B2(new_n269), .ZN(new_n273));
  NOR2_X1   g0073(.A1(new_n271), .A2(new_n273), .ZN(new_n274));
  NOR2_X1   g0074(.A1(KEYINPUT72), .A2(KEYINPUT9), .ZN(new_n275));
  NOR2_X1   g0075(.A1(new_n274), .A2(new_n275), .ZN(new_n276));
  INV_X1    g0076(.A(G41), .ZN(new_n277));
  INV_X1    g0077(.A(G45), .ZN(new_n278));
  AOI21_X1  g0078(.A(G1), .B1(new_n277), .B2(new_n278), .ZN(new_n279));
  INV_X1    g0079(.A(new_n279), .ZN(new_n280));
  OAI211_X1 g0080(.A(G1), .B(G13), .C1(new_n250), .C2(new_n277), .ZN(new_n281));
  NAND2_X1  g0081(.A1(new_n280), .A2(new_n281), .ZN(new_n282));
  INV_X1    g0082(.A(KEYINPUT65), .ZN(new_n283));
  OAI211_X1 g0083(.A(new_n283), .B(new_n265), .C1(G41), .C2(G45), .ZN(new_n284));
  NAND3_X1  g0084(.A1(new_n281), .A2(G274), .A3(new_n284), .ZN(new_n285));
  NOR2_X1   g0085(.A1(new_n279), .A2(new_n283), .ZN(new_n286));
  OAI22_X1  g0086(.A1(new_n282), .A2(new_n220), .B1(new_n285), .B2(new_n286), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n250), .A2(KEYINPUT3), .ZN(new_n288));
  INV_X1    g0088(.A(KEYINPUT3), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n289), .A2(G33), .ZN(new_n290));
  NAND2_X1  g0090(.A1(new_n288), .A2(new_n290), .ZN(new_n291));
  NOR2_X1   g0091(.A1(new_n291), .A2(G1698), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n292), .A2(G222), .ZN(new_n293));
  INV_X1    g0093(.A(G77), .ZN(new_n294));
  NOR2_X1   g0094(.A1(new_n289), .A2(G33), .ZN(new_n295));
  NOR2_X1   g0095(.A1(new_n250), .A2(KEYINPUT3), .ZN(new_n296));
  NOR2_X1   g0096(.A1(new_n295), .A2(new_n296), .ZN(new_n297));
  INV_X1    g0097(.A(G223), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n297), .A2(G1698), .ZN(new_n299));
  OAI221_X1 g0099(.A(new_n293), .B1(new_n294), .B2(new_n297), .C1(new_n298), .C2(new_n299), .ZN(new_n300));
  INV_X1    g0100(.A(KEYINPUT66), .ZN(new_n301));
  AOI21_X1  g0101(.A(new_n281), .B1(new_n300), .B2(new_n301), .ZN(new_n302));
  NOR2_X1   g0102(.A1(new_n299), .A2(new_n298), .ZN(new_n303));
  AOI21_X1  g0103(.A(new_n303), .B1(G77), .B2(new_n291), .ZN(new_n304));
  NAND3_X1  g0104(.A1(new_n304), .A2(KEYINPUT66), .A3(new_n293), .ZN(new_n305));
  AOI21_X1  g0105(.A(new_n287), .B1(new_n302), .B2(new_n305), .ZN(new_n306));
  INV_X1    g0106(.A(G200), .ZN(new_n307));
  NOR2_X1   g0107(.A1(new_n306), .A2(new_n307), .ZN(new_n308));
  INV_X1    g0108(.A(KEYINPUT73), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n302), .A2(new_n305), .ZN(new_n310));
  INV_X1    g0110(.A(new_n287), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n310), .A2(new_n311), .ZN(new_n312));
  INV_X1    g0112(.A(G190), .ZN(new_n313));
  OAI22_X1  g0113(.A1(new_n308), .A2(new_n309), .B1(new_n312), .B2(new_n313), .ZN(new_n314));
  INV_X1    g0114(.A(KEYINPUT10), .ZN(new_n315));
  NAND3_X1  g0115(.A1(new_n306), .A2(KEYINPUT73), .A3(G190), .ZN(new_n316));
  NAND4_X1  g0116(.A1(new_n276), .A2(new_n314), .A3(new_n315), .A4(new_n316), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n312), .A2(G200), .ZN(new_n318));
  AOI22_X1  g0118(.A1(new_n318), .A2(KEYINPUT73), .B1(G190), .B2(new_n306), .ZN(new_n319));
  INV_X1    g0119(.A(new_n275), .ZN(new_n320));
  OAI211_X1 g0120(.A(new_n316), .B(new_n320), .C1(new_n273), .C2(new_n271), .ZN(new_n321));
  OAI21_X1  g0121(.A(KEYINPUT10), .B1(new_n319), .B2(new_n321), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n317), .A2(new_n322), .ZN(new_n323));
  OAI21_X1  g0123(.A(new_n270), .B1(new_n306), .B2(G169), .ZN(new_n324));
  NOR2_X1   g0124(.A1(new_n324), .A2(KEYINPUT69), .ZN(new_n325));
  INV_X1    g0125(.A(KEYINPUT70), .ZN(new_n326));
  INV_X1    g0126(.A(G179), .ZN(new_n327));
  AOI21_X1  g0127(.A(new_n326), .B1(new_n306), .B2(new_n327), .ZN(new_n328));
  NOR3_X1   g0128(.A1(new_n312), .A2(KEYINPUT70), .A3(G179), .ZN(new_n329));
  NOR3_X1   g0129(.A1(new_n325), .A2(new_n328), .A3(new_n329), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n324), .A2(KEYINPUT69), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n330), .A2(new_n331), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n323), .A2(new_n332), .ZN(new_n333));
  INV_X1    g0133(.A(new_n285), .ZN(new_n334));
  INV_X1    g0134(.A(new_n286), .ZN(new_n335));
  AOI21_X1  g0135(.A(new_n213), .B1(G33), .B2(G41), .ZN(new_n336));
  NOR2_X1   g0136(.A1(new_n336), .A2(new_n279), .ZN(new_n337));
  AOI22_X1  g0137(.A1(new_n334), .A2(new_n335), .B1(new_n337), .B2(G232), .ZN(new_n338));
  NOR2_X1   g0138(.A1(G223), .A2(G1698), .ZN(new_n339));
  AOI21_X1  g0139(.A(new_n339), .B1(new_n220), .B2(G1698), .ZN(new_n340));
  AND2_X1   g0140(.A1(KEYINPUT77), .A2(KEYINPUT3), .ZN(new_n341));
  NOR2_X1   g0141(.A1(KEYINPUT77), .A2(KEYINPUT3), .ZN(new_n342));
  OAI21_X1  g0142(.A(G33), .B1(new_n341), .B2(new_n342), .ZN(new_n343));
  NAND3_X1  g0143(.A1(new_n340), .A2(new_n343), .A3(new_n288), .ZN(new_n344));
  NAND2_X1  g0144(.A1(G33), .A2(G87), .ZN(new_n345));
  AND2_X1   g0145(.A1(new_n344), .A2(new_n345), .ZN(new_n346));
  OAI211_X1 g0146(.A(new_n338), .B(G190), .C1(new_n346), .C2(new_n281), .ZN(new_n347));
  AOI21_X1  g0147(.A(new_n281), .B1(new_n344), .B2(new_n345), .ZN(new_n348));
  OAI22_X1  g0148(.A1(new_n282), .A2(new_n225), .B1(new_n285), .B2(new_n286), .ZN(new_n349));
  OAI21_X1  g0149(.A(G200), .B1(new_n348), .B2(new_n349), .ZN(new_n350));
  AND2_X1   g0150(.A1(new_n347), .A2(new_n350), .ZN(new_n351));
  INV_X1    g0151(.A(KEYINPUT16), .ZN(new_n352));
  INV_X1    g0152(.A(KEYINPUT7), .ZN(new_n353));
  NOR2_X1   g0153(.A1(new_n353), .A2(G20), .ZN(new_n354));
  NOR3_X1   g0154(.A1(new_n341), .A2(new_n342), .A3(G33), .ZN(new_n355));
  OAI21_X1  g0155(.A(new_n354), .B1(new_n355), .B2(new_n296), .ZN(new_n356));
  OAI21_X1  g0156(.A(new_n353), .B1(new_n297), .B2(G20), .ZN(new_n357));
  AOI21_X1  g0157(.A(new_n226), .B1(new_n356), .B2(new_n357), .ZN(new_n358));
  NOR2_X1   g0158(.A1(new_n224), .A2(new_n226), .ZN(new_n359));
  OAI21_X1  g0159(.A(G20), .B1(new_n359), .B2(new_n201), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n252), .A2(G159), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n360), .A2(new_n361), .ZN(new_n362));
  OAI21_X1  g0162(.A(new_n352), .B1(new_n358), .B2(new_n362), .ZN(new_n363));
  INV_X1    g0163(.A(new_n362), .ZN(new_n364));
  AOI21_X1  g0164(.A(G20), .B1(new_n343), .B2(new_n288), .ZN(new_n365));
  OAI21_X1  g0165(.A(G68), .B1(new_n365), .B2(new_n353), .ZN(new_n366));
  XNOR2_X1  g0166(.A(KEYINPUT77), .B(KEYINPUT3), .ZN(new_n367));
  AOI21_X1  g0167(.A(new_n295), .B1(new_n367), .B2(G33), .ZN(new_n368));
  NOR3_X1   g0168(.A1(new_n368), .A2(KEYINPUT7), .A3(G20), .ZN(new_n369));
  OAI211_X1 g0169(.A(KEYINPUT16), .B(new_n364), .C1(new_n366), .C2(new_n369), .ZN(new_n370));
  NAND3_X1  g0170(.A1(new_n363), .A2(new_n370), .A3(new_n263), .ZN(new_n371));
  INV_X1    g0171(.A(new_n259), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n372), .A2(new_n268), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n259), .A2(new_n266), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n373), .A2(new_n374), .ZN(new_n375));
  NAND3_X1  g0175(.A1(new_n351), .A2(new_n371), .A3(new_n375), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n376), .A2(KEYINPUT17), .ZN(new_n377));
  INV_X1    g0177(.A(KEYINPUT17), .ZN(new_n378));
  NAND4_X1  g0178(.A1(new_n351), .A2(new_n371), .A3(new_n378), .A4(new_n375), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n371), .A2(new_n375), .ZN(new_n380));
  OAI21_X1  g0180(.A(new_n338), .B1(new_n346), .B2(new_n281), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n381), .A2(G169), .ZN(new_n382));
  OAI21_X1  g0182(.A(new_n382), .B1(new_n381), .B2(new_n327), .ZN(new_n383));
  AOI21_X1  g0183(.A(KEYINPUT18), .B1(new_n380), .B2(new_n383), .ZN(new_n384));
  INV_X1    g0184(.A(KEYINPUT78), .ZN(new_n385));
  AOI22_X1  g0185(.A1(new_n377), .A2(new_n379), .B1(new_n384), .B2(new_n385), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n380), .A2(new_n383), .ZN(new_n387));
  INV_X1    g0187(.A(KEYINPUT18), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n387), .A2(new_n388), .ZN(new_n389));
  NAND3_X1  g0189(.A1(new_n380), .A2(KEYINPUT18), .A3(new_n383), .ZN(new_n390));
  NAND3_X1  g0190(.A1(new_n389), .A2(KEYINPUT78), .A3(new_n390), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n386), .A2(new_n391), .ZN(new_n392));
  NAND3_X1  g0192(.A1(new_n297), .A2(G232), .A3(G1698), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n393), .A2(KEYINPUT74), .ZN(new_n394));
  INV_X1    g0194(.A(KEYINPUT74), .ZN(new_n395));
  NAND4_X1  g0195(.A1(new_n297), .A2(new_n395), .A3(G232), .A4(G1698), .ZN(new_n396));
  NAND2_X1  g0196(.A1(G33), .A2(G97), .ZN(new_n397));
  NAND2_X1  g0197(.A1(new_n292), .A2(G226), .ZN(new_n398));
  NAND4_X1  g0198(.A1(new_n394), .A2(new_n396), .A3(new_n397), .A4(new_n398), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n399), .A2(new_n336), .ZN(new_n400));
  OAI22_X1  g0200(.A1(new_n282), .A2(new_n227), .B1(new_n285), .B2(new_n286), .ZN(new_n401));
  INV_X1    g0201(.A(new_n401), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n400), .A2(new_n402), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n403), .A2(KEYINPUT13), .ZN(new_n404));
  INV_X1    g0204(.A(KEYINPUT13), .ZN(new_n405));
  NAND3_X1  g0205(.A1(new_n400), .A2(new_n402), .A3(new_n405), .ZN(new_n406));
  NAND3_X1  g0206(.A1(new_n404), .A2(G190), .A3(new_n406), .ZN(new_n407));
  AOI21_X1  g0207(.A(new_n405), .B1(new_n400), .B2(new_n402), .ZN(new_n408));
  AOI211_X1 g0208(.A(KEYINPUT13), .B(new_n401), .C1(new_n399), .C2(new_n336), .ZN(new_n409));
  OAI21_X1  g0209(.A(G200), .B1(new_n408), .B2(new_n409), .ZN(new_n410));
  OAI211_X1 g0210(.A(new_n267), .B(KEYINPUT71), .C1(G1), .C2(new_n214), .ZN(new_n411));
  NOR2_X1   g0211(.A1(new_n411), .A2(new_n226), .ZN(new_n412));
  XOR2_X1   g0212(.A(new_n412), .B(KEYINPUT75), .Z(new_n413));
  NAND3_X1  g0213(.A1(new_n214), .A2(G33), .A3(G77), .ZN(new_n414));
  OAI221_X1 g0214(.A(new_n414), .B1(new_n214), .B2(G68), .C1(new_n251), .C2(new_n202), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n415), .A2(new_n263), .ZN(new_n416));
  XNOR2_X1  g0216(.A(new_n416), .B(KEYINPUT11), .ZN(new_n417));
  INV_X1    g0217(.A(new_n266), .ZN(new_n418));
  AOI21_X1  g0218(.A(KEYINPUT12), .B1(new_n418), .B2(new_n226), .ZN(new_n419));
  INV_X1    g0219(.A(KEYINPUT71), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n266), .A2(new_n420), .ZN(new_n421));
  NAND4_X1  g0221(.A1(new_n265), .A2(KEYINPUT71), .A3(G13), .A4(G20), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n421), .A2(new_n422), .ZN(new_n423));
  AND2_X1   g0223(.A1(new_n226), .A2(KEYINPUT12), .ZN(new_n424));
  AOI21_X1  g0224(.A(new_n419), .B1(new_n423), .B2(new_n424), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n417), .A2(new_n425), .ZN(new_n426));
  NOR2_X1   g0226(.A1(new_n413), .A2(new_n426), .ZN(new_n427));
  NAND3_X1  g0227(.A1(new_n407), .A2(new_n410), .A3(new_n427), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n428), .A2(KEYINPUT76), .ZN(new_n429));
  INV_X1    g0229(.A(KEYINPUT76), .ZN(new_n430));
  NAND4_X1  g0230(.A1(new_n407), .A2(new_n410), .A3(new_n430), .A4(new_n427), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n429), .A2(new_n431), .ZN(new_n432));
  OAI21_X1  g0232(.A(G169), .B1(new_n408), .B2(new_n409), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n433), .A2(KEYINPUT14), .ZN(new_n434));
  INV_X1    g0234(.A(KEYINPUT14), .ZN(new_n435));
  OAI211_X1 g0235(.A(new_n435), .B(G169), .C1(new_n408), .C2(new_n409), .ZN(new_n436));
  NAND3_X1  g0236(.A1(new_n404), .A2(G179), .A3(new_n406), .ZN(new_n437));
  NAND3_X1  g0237(.A1(new_n434), .A2(new_n436), .A3(new_n437), .ZN(new_n438));
  OR2_X1    g0238(.A1(new_n413), .A2(new_n426), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n438), .A2(new_n439), .ZN(new_n440));
  NAND2_X1  g0240(.A1(new_n432), .A2(new_n440), .ZN(new_n441));
  INV_X1    g0241(.A(new_n255), .ZN(new_n442));
  OR2_X1    g0242(.A1(new_n442), .A2(new_n257), .ZN(new_n443));
  AOI22_X1  g0243(.A1(new_n443), .A2(new_n252), .B1(G20), .B2(G77), .ZN(new_n444));
  XNOR2_X1  g0244(.A(KEYINPUT15), .B(G87), .ZN(new_n445));
  OR2_X1    g0245(.A1(new_n445), .A2(new_n260), .ZN(new_n446));
  AOI21_X1  g0246(.A(new_n267), .B1(new_n444), .B2(new_n446), .ZN(new_n447));
  NAND2_X1  g0247(.A1(new_n423), .A2(new_n294), .ZN(new_n448));
  OAI21_X1  g0248(.A(new_n448), .B1(new_n411), .B2(new_n294), .ZN(new_n449));
  OR2_X1    g0249(.A1(new_n447), .A2(new_n449), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n292), .A2(G232), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n291), .A2(G107), .ZN(new_n452));
  OAI211_X1 g0252(.A(new_n451), .B(new_n452), .C1(new_n227), .C2(new_n299), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n453), .A2(new_n336), .ZN(new_n454));
  AND2_X1   g0254(.A1(new_n337), .A2(G244), .ZN(new_n455));
  NOR2_X1   g0255(.A1(new_n285), .A2(new_n286), .ZN(new_n456));
  NOR2_X1   g0256(.A1(new_n455), .A2(new_n456), .ZN(new_n457));
  NAND3_X1  g0257(.A1(new_n454), .A2(new_n457), .A3(new_n327), .ZN(new_n458));
  AOI211_X1 g0258(.A(new_n456), .B(new_n455), .C1(new_n453), .C2(new_n336), .ZN(new_n459));
  OAI211_X1 g0259(.A(new_n450), .B(new_n458), .C1(new_n459), .C2(G169), .ZN(new_n460));
  NAND3_X1  g0260(.A1(new_n454), .A2(new_n457), .A3(G190), .ZN(new_n461));
  NOR2_X1   g0261(.A1(new_n447), .A2(new_n449), .ZN(new_n462));
  OAI211_X1 g0262(.A(new_n461), .B(new_n462), .C1(new_n459), .C2(new_n307), .ZN(new_n463));
  AND2_X1   g0263(.A1(new_n460), .A2(new_n463), .ZN(new_n464));
  INV_X1    g0264(.A(new_n464), .ZN(new_n465));
  NOR4_X1   g0265(.A1(new_n333), .A2(new_n392), .A3(new_n441), .A4(new_n465), .ZN(new_n466));
  INV_X1    g0266(.A(new_n466), .ZN(new_n467));
  INV_X1    g0267(.A(G1698), .ZN(new_n468));
  NAND4_X1  g0268(.A1(new_n343), .A2(G244), .A3(new_n468), .A4(new_n288), .ZN(new_n469));
  INV_X1    g0269(.A(KEYINPUT4), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n469), .A2(new_n470), .ZN(new_n471));
  AND2_X1   g0271(.A1(KEYINPUT4), .A2(G244), .ZN(new_n472));
  NAND4_X1  g0272(.A1(new_n288), .A2(new_n290), .A3(new_n472), .A4(new_n468), .ZN(new_n473));
  NAND4_X1  g0273(.A1(new_n288), .A2(new_n290), .A3(G250), .A4(G1698), .ZN(new_n474));
  NAND2_X1  g0274(.A1(G33), .A2(G283), .ZN(new_n475));
  AND3_X1   g0275(.A1(new_n473), .A2(new_n474), .A3(new_n475), .ZN(new_n476));
  AOI21_X1  g0276(.A(new_n281), .B1(new_n471), .B2(new_n476), .ZN(new_n477));
  INV_X1    g0277(.A(new_n477), .ZN(new_n478));
  INV_X1    g0278(.A(KEYINPUT5), .ZN(new_n479));
  OAI21_X1  g0279(.A(KEYINPUT81), .B1(new_n479), .B2(G41), .ZN(new_n480));
  INV_X1    g0280(.A(KEYINPUT81), .ZN(new_n481));
  NAND3_X1  g0281(.A1(new_n481), .A2(new_n277), .A3(KEYINPUT5), .ZN(new_n482));
  AND2_X1   g0282(.A1(new_n480), .A2(new_n482), .ZN(new_n483));
  OAI211_X1 g0283(.A(new_n265), .B(G45), .C1(new_n277), .C2(KEYINPUT5), .ZN(new_n484));
  OAI211_X1 g0284(.A(G257), .B(new_n281), .C1(new_n483), .C2(new_n484), .ZN(new_n485));
  AOI21_X1  g0285(.A(new_n484), .B1(new_n480), .B2(new_n482), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n486), .A2(G274), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n485), .A2(new_n487), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n488), .A2(KEYINPUT82), .ZN(new_n489));
  INV_X1    g0289(.A(KEYINPUT82), .ZN(new_n490));
  NAND3_X1  g0290(.A1(new_n485), .A2(new_n490), .A3(new_n487), .ZN(new_n491));
  NAND3_X1  g0291(.A1(new_n478), .A2(new_n489), .A3(new_n491), .ZN(new_n492));
  INV_X1    g0292(.A(G169), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  NAND4_X1  g0294(.A1(new_n478), .A2(new_n489), .A3(new_n327), .A4(new_n491), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  NOR2_X1   g0296(.A1(new_n250), .A2(G1), .ZN(new_n497));
  NOR2_X1   g0297(.A1(new_n263), .A2(new_n497), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n498), .A2(new_n266), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n499), .A2(G97), .ZN(new_n500));
  INV_X1    g0300(.A(KEYINPUT80), .ZN(new_n501));
  INV_X1    g0301(.A(G97), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n266), .A2(new_n502), .ZN(new_n503));
  AND3_X1   g0303(.A1(new_n500), .A2(new_n501), .A3(new_n503), .ZN(new_n504));
  AOI21_X1  g0304(.A(new_n501), .B1(new_n500), .B2(new_n503), .ZN(new_n505));
  NOR2_X1   g0305(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  INV_X1    g0306(.A(G107), .ZN(new_n507));
  AOI21_X1  g0307(.A(new_n507), .B1(new_n356), .B2(new_n357), .ZN(new_n508));
  INV_X1    g0308(.A(KEYINPUT6), .ZN(new_n509));
  NOR3_X1   g0309(.A1(new_n509), .A2(new_n502), .A3(G107), .ZN(new_n510));
  XNOR2_X1  g0310(.A(G97), .B(G107), .ZN(new_n511));
  AOI21_X1  g0311(.A(new_n510), .B1(new_n509), .B2(new_n511), .ZN(new_n512));
  OAI22_X1  g0312(.A1(new_n512), .A2(new_n214), .B1(new_n294), .B2(new_n251), .ZN(new_n513));
  OAI21_X1  g0313(.A(new_n263), .B1(new_n508), .B2(new_n513), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n514), .A2(KEYINPUT79), .ZN(new_n515));
  INV_X1    g0315(.A(KEYINPUT79), .ZN(new_n516));
  OAI211_X1 g0316(.A(new_n516), .B(new_n263), .C1(new_n508), .C2(new_n513), .ZN(new_n517));
  AOI21_X1  g0317(.A(new_n506), .B1(new_n515), .B2(new_n517), .ZN(new_n518));
  NOR2_X1   g0318(.A1(new_n496), .A2(new_n518), .ZN(new_n519));
  NAND4_X1  g0319(.A1(new_n478), .A2(new_n489), .A3(new_n313), .A4(new_n491), .ZN(new_n520));
  AND3_X1   g0320(.A1(new_n485), .A2(new_n490), .A3(new_n487), .ZN(new_n521));
  AOI21_X1  g0321(.A(new_n490), .B1(new_n485), .B2(new_n487), .ZN(new_n522));
  NOR3_X1   g0322(.A1(new_n521), .A2(new_n477), .A3(new_n522), .ZN(new_n523));
  OAI21_X1  g0323(.A(new_n520), .B1(new_n523), .B2(G200), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n524), .A2(new_n518), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n525), .A2(KEYINPUT83), .ZN(new_n526));
  INV_X1    g0326(.A(KEYINPUT83), .ZN(new_n527));
  NAND3_X1  g0327(.A1(new_n524), .A2(new_n518), .A3(new_n527), .ZN(new_n528));
  AOI21_X1  g0328(.A(new_n519), .B1(new_n526), .B2(new_n528), .ZN(new_n529));
  INV_X1    g0329(.A(KEYINPUT24), .ZN(new_n530));
  NOR4_X1   g0330(.A1(new_n291), .A2(KEYINPUT22), .A3(G20), .A4(new_n221), .ZN(new_n531));
  NOR2_X1   g0331(.A1(new_n221), .A2(G20), .ZN(new_n532));
  NAND3_X1  g0332(.A1(new_n343), .A2(new_n288), .A3(new_n532), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n533), .A2(KEYINPUT86), .ZN(new_n534));
  INV_X1    g0334(.A(KEYINPUT86), .ZN(new_n535));
  NAND4_X1  g0335(.A1(new_n343), .A2(new_n535), .A3(new_n288), .A4(new_n532), .ZN(new_n536));
  NAND3_X1  g0336(.A1(new_n534), .A2(KEYINPUT22), .A3(new_n536), .ZN(new_n537));
  INV_X1    g0337(.A(KEYINPUT87), .ZN(new_n538));
  AOI21_X1  g0338(.A(new_n531), .B1(new_n537), .B2(new_n538), .ZN(new_n539));
  NAND4_X1  g0339(.A1(new_n534), .A2(KEYINPUT87), .A3(KEYINPUT22), .A4(new_n536), .ZN(new_n540));
  AND2_X1   g0340(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  NAND3_X1  g0341(.A1(new_n214), .A2(G33), .A3(G116), .ZN(new_n542));
  INV_X1    g0342(.A(KEYINPUT88), .ZN(new_n543));
  INV_X1    g0343(.A(KEYINPUT23), .ZN(new_n544));
  OAI211_X1 g0344(.A(G20), .B(new_n507), .C1(new_n543), .C2(new_n544), .ZN(new_n545));
  AOI21_X1  g0345(.A(new_n545), .B1(new_n543), .B2(new_n544), .ZN(new_n546));
  AOI211_X1 g0346(.A(KEYINPUT88), .B(KEYINPUT23), .C1(new_n507), .C2(G20), .ZN(new_n547));
  OAI21_X1  g0347(.A(new_n542), .B1(new_n546), .B2(new_n547), .ZN(new_n548));
  OAI21_X1  g0348(.A(new_n530), .B1(new_n541), .B2(new_n548), .ZN(new_n549));
  AOI21_X1  g0349(.A(new_n548), .B1(new_n539), .B2(new_n540), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n550), .A2(KEYINPUT24), .ZN(new_n551));
  NAND3_X1  g0351(.A1(new_n549), .A2(new_n263), .A3(new_n551), .ZN(new_n552));
  OAI21_X1  g0352(.A(KEYINPUT25), .B1(new_n266), .B2(G107), .ZN(new_n553));
  OR3_X1    g0353(.A1(new_n266), .A2(KEYINPUT25), .A3(G107), .ZN(new_n554));
  OAI211_X1 g0354(.A(new_n553), .B(new_n554), .C1(new_n499), .C2(new_n507), .ZN(new_n555));
  XOR2_X1   g0355(.A(new_n555), .B(KEYINPUT89), .Z(new_n556));
  NAND3_X1  g0356(.A1(new_n368), .A2(G250), .A3(new_n468), .ZN(new_n557));
  INV_X1    g0357(.A(KEYINPUT90), .ZN(new_n558));
  NOR2_X1   g0358(.A1(new_n210), .A2(new_n468), .ZN(new_n559));
  NAND3_X1  g0359(.A1(new_n368), .A2(new_n558), .A3(new_n559), .ZN(new_n560));
  NAND3_X1  g0360(.A1(new_n343), .A2(new_n288), .A3(new_n559), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n561), .A2(KEYINPUT90), .ZN(new_n562));
  NAND2_X1  g0362(.A1(G33), .A2(G294), .ZN(new_n563));
  NAND4_X1  g0363(.A1(new_n557), .A2(new_n560), .A3(new_n562), .A4(new_n563), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n480), .A2(new_n482), .ZN(new_n565));
  INV_X1    g0365(.A(new_n484), .ZN(new_n566));
  AOI21_X1  g0366(.A(new_n336), .B1(new_n565), .B2(new_n566), .ZN(new_n567));
  AOI22_X1  g0367(.A1(new_n564), .A2(new_n336), .B1(G264), .B2(new_n567), .ZN(new_n568));
  AOI21_X1  g0368(.A(new_n307), .B1(new_n568), .B2(new_n487), .ZN(new_n569));
  AND2_X1   g0369(.A1(new_n568), .A2(new_n487), .ZN(new_n570));
  AOI21_X1  g0370(.A(new_n569), .B1(G190), .B2(new_n570), .ZN(new_n571));
  NAND3_X1  g0371(.A1(new_n552), .A2(new_n556), .A3(new_n571), .ZN(new_n572));
  OAI21_X1  g0372(.A(new_n263), .B1(new_n550), .B2(KEYINPUT24), .ZN(new_n573));
  AOI211_X1 g0373(.A(new_n530), .B(new_n548), .C1(new_n539), .C2(new_n540), .ZN(new_n574));
  OAI21_X1  g0374(.A(new_n556), .B1(new_n573), .B2(new_n574), .ZN(new_n575));
  AOI21_X1  g0375(.A(G169), .B1(new_n568), .B2(new_n487), .ZN(new_n576));
  AOI21_X1  g0376(.A(new_n576), .B1(new_n327), .B2(new_n570), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n575), .A2(new_n577), .ZN(new_n578));
  NAND4_X1  g0378(.A1(new_n343), .A2(G238), .A3(new_n468), .A4(new_n288), .ZN(new_n579));
  NAND4_X1  g0379(.A1(new_n343), .A2(G244), .A3(G1698), .A4(new_n288), .ZN(new_n580));
  OAI211_X1 g0380(.A(new_n579), .B(new_n580), .C1(new_n250), .C2(new_n241), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n581), .A2(new_n336), .ZN(new_n582));
  NOR2_X1   g0382(.A1(new_n278), .A2(G1), .ZN(new_n583));
  NOR2_X1   g0383(.A1(new_n583), .A2(new_n206), .ZN(new_n584));
  AOI22_X1  g0384(.A1(new_n584), .A2(new_n281), .B1(G274), .B2(new_n583), .ZN(new_n585));
  NAND3_X1  g0385(.A1(new_n582), .A2(new_n327), .A3(new_n585), .ZN(new_n586));
  NAND4_X1  g0386(.A1(new_n343), .A2(new_n214), .A3(G68), .A4(new_n288), .ZN(new_n587));
  INV_X1    g0387(.A(KEYINPUT19), .ZN(new_n588));
  OAI21_X1  g0388(.A(new_n214), .B1(new_n397), .B2(new_n588), .ZN(new_n589));
  NAND3_X1  g0389(.A1(new_n221), .A2(new_n502), .A3(new_n507), .ZN(new_n590));
  NAND3_X1  g0390(.A1(new_n214), .A2(G33), .A3(G97), .ZN(new_n591));
  AOI22_X1  g0391(.A1(new_n589), .A2(new_n590), .B1(new_n588), .B2(new_n591), .ZN(new_n592));
  AOI21_X1  g0392(.A(new_n267), .B1(new_n587), .B2(new_n592), .ZN(new_n593));
  AND2_X1   g0393(.A1(new_n423), .A2(new_n445), .ZN(new_n594));
  NOR2_X1   g0394(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  XNOR2_X1  g0395(.A(new_n445), .B(KEYINPUT84), .ZN(new_n596));
  NAND3_X1  g0396(.A1(new_n596), .A2(new_n266), .A3(new_n498), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n595), .A2(new_n597), .ZN(new_n598));
  INV_X1    g0398(.A(new_n585), .ZN(new_n599));
  AOI21_X1  g0399(.A(new_n599), .B1(new_n581), .B2(new_n336), .ZN(new_n600));
  OAI211_X1 g0400(.A(new_n586), .B(new_n598), .C1(G169), .C2(new_n600), .ZN(new_n601));
  NAND3_X1  g0401(.A1(new_n582), .A2(G190), .A3(new_n585), .ZN(new_n602));
  NOR2_X1   g0402(.A1(new_n499), .A2(new_n221), .ZN(new_n603));
  NOR3_X1   g0403(.A1(new_n593), .A2(new_n603), .A3(new_n594), .ZN(new_n604));
  OAI211_X1 g0404(.A(new_n602), .B(new_n604), .C1(new_n307), .C2(new_n600), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n601), .A2(new_n605), .ZN(new_n606));
  INV_X1    g0406(.A(KEYINPUT85), .ZN(new_n607));
  NOR2_X1   g0407(.A1(new_n607), .A2(KEYINPUT21), .ZN(new_n608));
  NAND4_X1  g0408(.A1(new_n498), .A2(G116), .A3(new_n421), .A4(new_n422), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n423), .A2(new_n241), .ZN(new_n610));
  AOI22_X1  g0410(.A1(new_n262), .A2(new_n213), .B1(G20), .B2(new_n241), .ZN(new_n611));
  OAI211_X1 g0411(.A(new_n475), .B(new_n214), .C1(G33), .C2(new_n502), .ZN(new_n612));
  AND3_X1   g0412(.A1(new_n611), .A2(KEYINPUT20), .A3(new_n612), .ZN(new_n613));
  AOI21_X1  g0413(.A(KEYINPUT20), .B1(new_n611), .B2(new_n612), .ZN(new_n614));
  OAI211_X1 g0414(.A(new_n609), .B(new_n610), .C1(new_n613), .C2(new_n614), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n615), .A2(G169), .ZN(new_n616));
  OAI211_X1 g0416(.A(G270), .B(new_n281), .C1(new_n483), .C2(new_n484), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n617), .A2(new_n487), .ZN(new_n618));
  NOR2_X1   g0418(.A1(G257), .A2(G1698), .ZN(new_n619));
  AOI21_X1  g0419(.A(new_n619), .B1(new_n211), .B2(G1698), .ZN(new_n620));
  NAND3_X1  g0420(.A1(new_n620), .A2(new_n343), .A3(new_n288), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n291), .A2(G303), .ZN(new_n622));
  AOI21_X1  g0422(.A(new_n281), .B1(new_n621), .B2(new_n622), .ZN(new_n623));
  NOR2_X1   g0423(.A1(new_n618), .A2(new_n623), .ZN(new_n624));
  OAI21_X1  g0424(.A(new_n608), .B1(new_n616), .B2(new_n624), .ZN(new_n625));
  INV_X1    g0425(.A(new_n623), .ZN(new_n626));
  AOI22_X1  g0426(.A1(new_n567), .A2(G270), .B1(G274), .B2(new_n486), .ZN(new_n627));
  NAND3_X1  g0427(.A1(new_n626), .A2(new_n627), .A3(G190), .ZN(new_n628));
  OAI21_X1  g0428(.A(G200), .B1(new_n618), .B2(new_n623), .ZN(new_n629));
  INV_X1    g0429(.A(new_n615), .ZN(new_n630));
  NAND3_X1  g0430(.A1(new_n628), .A2(new_n629), .A3(new_n630), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n626), .A2(new_n627), .ZN(new_n632));
  INV_X1    g0432(.A(new_n608), .ZN(new_n633));
  NAND4_X1  g0433(.A1(new_n632), .A2(G169), .A3(new_n633), .A4(new_n615), .ZN(new_n634));
  NAND3_X1  g0434(.A1(new_n624), .A2(G179), .A3(new_n615), .ZN(new_n635));
  NAND4_X1  g0435(.A1(new_n625), .A2(new_n631), .A3(new_n634), .A4(new_n635), .ZN(new_n636));
  NOR2_X1   g0436(.A1(new_n606), .A2(new_n636), .ZN(new_n637));
  NAND4_X1  g0437(.A1(new_n529), .A2(new_n572), .A3(new_n578), .A4(new_n637), .ZN(new_n638));
  NOR2_X1   g0438(.A1(new_n467), .A2(new_n638), .ZN(G372));
  NAND2_X1  g0439(.A1(new_n377), .A2(new_n379), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n460), .A2(KEYINPUT92), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n454), .A2(new_n457), .ZN(new_n642));
  AOI21_X1  g0442(.A(new_n462), .B1(new_n642), .B2(new_n493), .ZN(new_n643));
  INV_X1    g0443(.A(KEYINPUT92), .ZN(new_n644));
  NAND3_X1  g0444(.A1(new_n643), .A2(new_n644), .A3(new_n458), .ZN(new_n645));
  AOI22_X1  g0445(.A1(new_n429), .A2(new_n431), .B1(new_n641), .B2(new_n645), .ZN(new_n646));
  INV_X1    g0446(.A(new_n440), .ZN(new_n647));
  OAI21_X1  g0447(.A(new_n640), .B1(new_n646), .B2(new_n647), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n389), .A2(new_n390), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n648), .A2(new_n649), .ZN(new_n650));
  AOI22_X1  g0450(.A1(new_n650), .A2(new_n323), .B1(new_n331), .B2(new_n330), .ZN(new_n651));
  NAND3_X1  g0451(.A1(new_n625), .A2(new_n634), .A3(new_n635), .ZN(new_n652));
  INV_X1    g0452(.A(new_n652), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n578), .A2(new_n653), .ZN(new_n654));
  AND2_X1   g0454(.A1(new_n586), .A2(new_n598), .ZN(new_n655));
  XOR2_X1   g0455(.A(new_n585), .B(KEYINPUT91), .Z(new_n656));
  NAND2_X1  g0456(.A1(new_n656), .A2(new_n582), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n657), .A2(new_n493), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n655), .A2(new_n658), .ZN(new_n659));
  AND2_X1   g0459(.A1(new_n602), .A2(new_n604), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n657), .A2(G200), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  AND2_X1   g0462(.A1(new_n659), .A2(new_n662), .ZN(new_n663));
  NAND4_X1  g0463(.A1(new_n654), .A2(new_n572), .A3(new_n529), .A4(new_n663), .ZN(new_n664));
  INV_X1    g0464(.A(KEYINPUT26), .ZN(new_n665));
  NAND3_X1  g0465(.A1(new_n663), .A2(new_n519), .A3(new_n665), .ZN(new_n666));
  INV_X1    g0466(.A(new_n518), .ZN(new_n667));
  NAND3_X1  g0467(.A1(new_n667), .A2(new_n494), .A3(new_n495), .ZN(new_n668));
  OAI21_X1  g0468(.A(KEYINPUT26), .B1(new_n668), .B2(new_n606), .ZN(new_n669));
  AND3_X1   g0469(.A1(new_n666), .A2(new_n669), .A3(new_n659), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n664), .A2(new_n670), .ZN(new_n671));
  INV_X1    g0471(.A(new_n671), .ZN(new_n672));
  OAI21_X1  g0472(.A(new_n651), .B1(new_n467), .B2(new_n672), .ZN(G369));
  INV_X1    g0473(.A(new_n572), .ZN(new_n674));
  INV_X1    g0474(.A(G13), .ZN(new_n675));
  NOR2_X1   g0475(.A1(new_n675), .A2(G20), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n676), .A2(new_n265), .ZN(new_n677));
  OR2_X1    g0477(.A1(new_n677), .A2(KEYINPUT27), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n677), .A2(KEYINPUT27), .ZN(new_n679));
  NAND3_X1  g0479(.A1(new_n678), .A2(G213), .A3(new_n679), .ZN(new_n680));
  INV_X1    g0480(.A(G343), .ZN(new_n681));
  NOR2_X1   g0481(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  INV_X1    g0482(.A(new_n682), .ZN(new_n683));
  AOI21_X1  g0483(.A(new_n683), .B1(new_n552), .B2(new_n556), .ZN(new_n684));
  OAI21_X1  g0484(.A(new_n578), .B1(new_n674), .B2(new_n684), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n568), .A2(new_n487), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n686), .A2(new_n493), .ZN(new_n687));
  OAI21_X1  g0487(.A(new_n687), .B1(G179), .B2(new_n686), .ZN(new_n688));
  AOI21_X1  g0488(.A(new_n688), .B1(new_n552), .B2(new_n556), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n689), .A2(new_n683), .ZN(new_n690));
  AND2_X1   g0490(.A1(new_n685), .A2(new_n690), .ZN(new_n691));
  NOR2_X1   g0491(.A1(new_n653), .A2(new_n682), .ZN(new_n692));
  NOR2_X1   g0492(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  NOR2_X1   g0493(.A1(new_n683), .A2(new_n630), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n652), .A2(new_n694), .ZN(new_n695));
  OAI21_X1  g0495(.A(new_n695), .B1(new_n636), .B2(new_n694), .ZN(new_n696));
  NAND2_X1  g0496(.A1(new_n696), .A2(G330), .ZN(new_n697));
  NOR2_X1   g0497(.A1(new_n693), .A2(new_n697), .ZN(new_n698));
  INV_X1    g0498(.A(new_n698), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n691), .A2(new_n692), .ZN(new_n700));
  AND2_X1   g0500(.A1(new_n700), .A2(new_n690), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n699), .A2(new_n701), .ZN(G399));
  NOR2_X1   g0502(.A1(new_n209), .A2(G41), .ZN(new_n703));
  INV_X1    g0503(.A(new_n703), .ZN(new_n704));
  NOR2_X1   g0504(.A1(new_n590), .A2(G116), .ZN(new_n705));
  NAND3_X1  g0505(.A1(new_n704), .A2(G1), .A3(new_n705), .ZN(new_n706));
  OAI21_X1  g0506(.A(new_n706), .B1(new_n217), .B2(new_n704), .ZN(new_n707));
  XNOR2_X1  g0507(.A(new_n707), .B(KEYINPUT28), .ZN(new_n708));
  AOI21_X1  g0508(.A(new_n682), .B1(new_n664), .B2(new_n670), .ZN(new_n709));
  INV_X1    g0509(.A(KEYINPUT95), .ZN(new_n710));
  OR3_X1    g0510(.A1(new_n709), .A2(new_n710), .A3(KEYINPUT29), .ZN(new_n711));
  OAI21_X1  g0511(.A(new_n710), .B1(new_n709), .B2(KEYINPUT29), .ZN(new_n712));
  AND3_X1   g0512(.A1(new_n524), .A2(new_n527), .A3(new_n518), .ZN(new_n713));
  AOI21_X1  g0513(.A(new_n527), .B1(new_n524), .B2(new_n518), .ZN(new_n714));
  OAI211_X1 g0514(.A(new_n663), .B(new_n668), .C1(new_n713), .C2(new_n714), .ZN(new_n715));
  AOI21_X1  g0515(.A(new_n652), .B1(new_n575), .B2(new_n577), .ZN(new_n716));
  NOR3_X1   g0516(.A1(new_n674), .A2(new_n715), .A3(new_n716), .ZN(new_n717));
  NAND2_X1  g0517(.A1(new_n662), .A2(new_n659), .ZN(new_n718));
  OAI21_X1  g0518(.A(KEYINPUT26), .B1(new_n668), .B2(new_n718), .ZN(new_n719));
  NAND4_X1  g0519(.A1(new_n519), .A2(new_n665), .A3(new_n601), .A4(new_n605), .ZN(new_n720));
  NAND3_X1  g0520(.A1(new_n719), .A2(new_n720), .A3(new_n659), .ZN(new_n721));
  OAI211_X1 g0521(.A(KEYINPUT29), .B(new_n683), .C1(new_n717), .C2(new_n721), .ZN(new_n722));
  NAND3_X1  g0522(.A1(new_n711), .A2(new_n712), .A3(new_n722), .ZN(new_n723));
  INV_X1    g0523(.A(KEYINPUT94), .ZN(new_n724));
  OAI21_X1  g0524(.A(new_n724), .B1(new_n638), .B2(new_n682), .ZN(new_n725));
  OAI211_X1 g0525(.A(new_n637), .B(new_n668), .C1(new_n713), .C2(new_n714), .ZN(new_n726));
  NOR2_X1   g0526(.A1(new_n726), .A2(new_n689), .ZN(new_n727));
  NAND4_X1  g0527(.A1(new_n727), .A2(KEYINPUT94), .A3(new_n572), .A4(new_n683), .ZN(new_n728));
  AND4_X1   g0528(.A1(new_n478), .A2(new_n600), .A3(new_n489), .A4(new_n491), .ZN(new_n729));
  INV_X1    g0529(.A(KEYINPUT30), .ZN(new_n730));
  NAND2_X1  g0530(.A1(new_n730), .A2(KEYINPUT93), .ZN(new_n731));
  AND3_X1   g0531(.A1(new_n624), .A2(G179), .A3(new_n731), .ZN(new_n732));
  NAND3_X1  g0532(.A1(new_n729), .A2(new_n568), .A3(new_n732), .ZN(new_n733));
  OAI21_X1  g0533(.A(new_n733), .B1(KEYINPUT93), .B2(new_n730), .ZN(new_n734));
  NOR2_X1   g0534(.A1(new_n730), .A2(KEYINPUT93), .ZN(new_n735));
  NAND4_X1  g0535(.A1(new_n729), .A2(new_n568), .A3(new_n735), .A4(new_n732), .ZN(new_n736));
  NOR2_X1   g0536(.A1(new_n624), .A2(G179), .ZN(new_n737));
  NAND4_X1  g0537(.A1(new_n686), .A2(new_n492), .A3(new_n657), .A4(new_n737), .ZN(new_n738));
  NAND3_X1  g0538(.A1(new_n734), .A2(new_n736), .A3(new_n738), .ZN(new_n739));
  AND3_X1   g0539(.A1(new_n739), .A2(KEYINPUT31), .A3(new_n682), .ZN(new_n740));
  AOI21_X1  g0540(.A(KEYINPUT31), .B1(new_n739), .B2(new_n682), .ZN(new_n741));
  NOR2_X1   g0541(.A1(new_n740), .A2(new_n741), .ZN(new_n742));
  NAND3_X1  g0542(.A1(new_n725), .A2(new_n728), .A3(new_n742), .ZN(new_n743));
  NAND2_X1  g0543(.A1(new_n743), .A2(G330), .ZN(new_n744));
  NAND2_X1  g0544(.A1(new_n723), .A2(new_n744), .ZN(new_n745));
  XNOR2_X1  g0545(.A(new_n745), .B(KEYINPUT96), .ZN(new_n746));
  OAI21_X1  g0546(.A(new_n708), .B1(new_n746), .B2(G1), .ZN(G364));
  NOR2_X1   g0547(.A1(new_n209), .A2(new_n291), .ZN(new_n748));
  AOI22_X1  g0548(.A1(new_n748), .A2(G355), .B1(new_n241), .B2(new_n209), .ZN(new_n749));
  NOR2_X1   g0549(.A1(new_n247), .A2(new_n278), .ZN(new_n750));
  NOR2_X1   g0550(.A1(new_n368), .A2(new_n209), .ZN(new_n751));
  OAI21_X1  g0551(.A(new_n751), .B1(G45), .B2(new_n217), .ZN(new_n752));
  OAI21_X1  g0552(.A(new_n749), .B1(new_n750), .B2(new_n752), .ZN(new_n753));
  INV_X1    g0553(.A(KEYINPUT98), .ZN(new_n754));
  OR2_X1    g0554(.A1(new_n753), .A2(new_n754), .ZN(new_n755));
  NAND2_X1  g0555(.A1(new_n753), .A2(new_n754), .ZN(new_n756));
  NOR2_X1   g0556(.A1(G13), .A2(G33), .ZN(new_n757));
  INV_X1    g0557(.A(new_n757), .ZN(new_n758));
  NOR2_X1   g0558(.A1(new_n758), .A2(G20), .ZN(new_n759));
  AOI21_X1  g0559(.A(new_n213), .B1(G20), .B2(new_n493), .ZN(new_n760));
  NOR2_X1   g0560(.A1(new_n759), .A2(new_n760), .ZN(new_n761));
  NAND3_X1  g0561(.A1(new_n755), .A2(new_n756), .A3(new_n761), .ZN(new_n762));
  AOI21_X1  g0562(.A(new_n265), .B1(new_n676), .B2(G45), .ZN(new_n763));
  INV_X1    g0563(.A(new_n763), .ZN(new_n764));
  NOR2_X1   g0564(.A1(new_n703), .A2(new_n764), .ZN(new_n765));
  INV_X1    g0565(.A(new_n765), .ZN(new_n766));
  NOR2_X1   g0566(.A1(new_n214), .A2(G190), .ZN(new_n767));
  INV_X1    g0567(.A(new_n767), .ZN(new_n768));
  NOR3_X1   g0568(.A1(new_n768), .A2(G179), .A3(new_n307), .ZN(new_n769));
  INV_X1    g0569(.A(new_n769), .ZN(new_n770));
  NOR2_X1   g0570(.A1(new_n770), .A2(new_n507), .ZN(new_n771));
  NOR2_X1   g0571(.A1(new_n327), .A2(new_n307), .ZN(new_n772));
  NAND2_X1  g0572(.A1(new_n772), .A2(new_n767), .ZN(new_n773));
  INV_X1    g0573(.A(new_n773), .ZN(new_n774));
  AOI21_X1  g0574(.A(new_n771), .B1(G68), .B2(new_n774), .ZN(new_n775));
  NOR2_X1   g0575(.A1(G179), .A2(G200), .ZN(new_n776));
  NAND2_X1  g0576(.A1(new_n767), .A2(new_n776), .ZN(new_n777));
  INV_X1    g0577(.A(G159), .ZN(new_n778));
  NOR2_X1   g0578(.A1(new_n777), .A2(new_n778), .ZN(new_n779));
  XNOR2_X1  g0579(.A(new_n779), .B(KEYINPUT32), .ZN(new_n780));
  NOR2_X1   g0580(.A1(new_n327), .A2(G200), .ZN(new_n781));
  NAND2_X1  g0581(.A1(new_n781), .A2(new_n767), .ZN(new_n782));
  OAI211_X1 g0582(.A(new_n775), .B(new_n780), .C1(new_n294), .C2(new_n782), .ZN(new_n783));
  NOR2_X1   g0583(.A1(new_n214), .A2(new_n313), .ZN(new_n784));
  NAND2_X1  g0584(.A1(new_n784), .A2(new_n772), .ZN(new_n785));
  INV_X1    g0585(.A(new_n785), .ZN(new_n786));
  AOI21_X1  g0586(.A(new_n291), .B1(new_n786), .B2(G50), .ZN(new_n787));
  NAND2_X1  g0587(.A1(new_n776), .A2(G190), .ZN(new_n788));
  NAND2_X1  g0588(.A1(new_n788), .A2(G20), .ZN(new_n789));
  NAND2_X1  g0589(.A1(new_n789), .A2(G97), .ZN(new_n790));
  NAND2_X1  g0590(.A1(new_n784), .A2(new_n781), .ZN(new_n791));
  INV_X1    g0591(.A(new_n791), .ZN(new_n792));
  NAND2_X1  g0592(.A1(new_n792), .A2(G58), .ZN(new_n793));
  NAND3_X1  g0593(.A1(new_n784), .A2(new_n327), .A3(G200), .ZN(new_n794));
  INV_X1    g0594(.A(new_n794), .ZN(new_n795));
  NAND2_X1  g0595(.A1(new_n795), .A2(G87), .ZN(new_n796));
  NAND4_X1  g0596(.A1(new_n787), .A2(new_n790), .A3(new_n793), .A4(new_n796), .ZN(new_n797));
  INV_X1    g0597(.A(new_n777), .ZN(new_n798));
  AOI22_X1  g0598(.A1(G322), .A2(new_n792), .B1(new_n798), .B2(G329), .ZN(new_n799));
  NAND2_X1  g0599(.A1(new_n786), .A2(G326), .ZN(new_n800));
  XOR2_X1   g0600(.A(KEYINPUT33), .B(G317), .Z(new_n801));
  OAI211_X1 g0601(.A(new_n799), .B(new_n800), .C1(new_n773), .C2(new_n801), .ZN(new_n802));
  INV_X1    g0602(.A(new_n782), .ZN(new_n803));
  AOI22_X1  g0603(.A1(new_n769), .A2(G283), .B1(new_n803), .B2(G311), .ZN(new_n804));
  AOI21_X1  g0604(.A(new_n297), .B1(new_n795), .B2(G303), .ZN(new_n805));
  INV_X1    g0605(.A(G294), .ZN(new_n806));
  INV_X1    g0606(.A(new_n789), .ZN(new_n807));
  OAI211_X1 g0607(.A(new_n804), .B(new_n805), .C1(new_n806), .C2(new_n807), .ZN(new_n808));
  OAI22_X1  g0608(.A1(new_n783), .A2(new_n797), .B1(new_n802), .B2(new_n808), .ZN(new_n809));
  AOI21_X1  g0609(.A(new_n766), .B1(new_n809), .B2(new_n760), .ZN(new_n810));
  INV_X1    g0610(.A(new_n759), .ZN(new_n811));
  OAI211_X1 g0611(.A(new_n762), .B(new_n810), .C1(new_n696), .C2(new_n811), .ZN(new_n812));
  OR2_X1    g0612(.A1(new_n696), .A2(G330), .ZN(new_n813));
  INV_X1    g0613(.A(KEYINPUT97), .ZN(new_n814));
  NAND2_X1  g0614(.A1(new_n813), .A2(new_n814), .ZN(new_n815));
  NAND3_X1  g0615(.A1(new_n815), .A2(new_n697), .A3(new_n766), .ZN(new_n816));
  NOR2_X1   g0616(.A1(new_n813), .A2(new_n814), .ZN(new_n817));
  OAI21_X1  g0617(.A(new_n812), .B1(new_n816), .B2(new_n817), .ZN(G396));
  NAND2_X1  g0618(.A1(new_n450), .A2(new_n682), .ZN(new_n819));
  NAND3_X1  g0619(.A1(new_n460), .A2(new_n463), .A3(new_n819), .ZN(new_n820));
  AND2_X1   g0620(.A1(new_n820), .A2(KEYINPUT101), .ZN(new_n821));
  NOR2_X1   g0621(.A1(new_n820), .A2(KEYINPUT101), .ZN(new_n822));
  AOI21_X1  g0622(.A(new_n819), .B1(new_n641), .B2(new_n645), .ZN(new_n823));
  NOR3_X1   g0623(.A1(new_n821), .A2(new_n822), .A3(new_n823), .ZN(new_n824));
  INV_X1    g0624(.A(new_n824), .ZN(new_n825));
  XNOR2_X1  g0625(.A(new_n709), .B(new_n825), .ZN(new_n826));
  OAI21_X1  g0626(.A(new_n766), .B1(new_n826), .B2(new_n744), .ZN(new_n827));
  AOI21_X1  g0627(.A(KEYINPUT102), .B1(new_n826), .B2(new_n744), .ZN(new_n828));
  NOR2_X1   g0628(.A1(new_n827), .A2(new_n828), .ZN(new_n829));
  NAND3_X1  g0629(.A1(new_n826), .A2(KEYINPUT102), .A3(new_n744), .ZN(new_n830));
  NAND2_X1  g0630(.A1(new_n829), .A2(new_n830), .ZN(new_n831));
  NOR2_X1   g0631(.A1(new_n760), .A2(new_n757), .ZN(new_n832));
  XOR2_X1   g0632(.A(new_n832), .B(KEYINPUT99), .Z(new_n833));
  OAI21_X1  g0633(.A(new_n765), .B1(new_n833), .B2(G77), .ZN(new_n834));
  AOI22_X1  g0634(.A1(new_n786), .A2(G137), .B1(new_n803), .B2(G159), .ZN(new_n835));
  INV_X1    g0635(.A(new_n835), .ZN(new_n836));
  INV_X1    g0636(.A(G143), .ZN(new_n837));
  INV_X1    g0637(.A(G150), .ZN(new_n838));
  OAI22_X1  g0638(.A1(new_n837), .A2(new_n791), .B1(new_n773), .B2(new_n838), .ZN(new_n839));
  XNOR2_X1  g0639(.A(KEYINPUT100), .B(KEYINPUT34), .ZN(new_n840));
  OR3_X1    g0640(.A1(new_n836), .A2(new_n839), .A3(new_n840), .ZN(new_n841));
  OAI21_X1  g0641(.A(new_n840), .B1(new_n836), .B2(new_n839), .ZN(new_n842));
  NAND2_X1  g0642(.A1(new_n769), .A2(G68), .ZN(new_n843));
  OAI21_X1  g0643(.A(new_n843), .B1(new_n202), .B2(new_n794), .ZN(new_n844));
  AOI21_X1  g0644(.A(new_n844), .B1(G132), .B2(new_n798), .ZN(new_n845));
  INV_X1    g0645(.A(new_n368), .ZN(new_n846));
  AOI21_X1  g0646(.A(new_n846), .B1(G58), .B2(new_n789), .ZN(new_n847));
  NAND4_X1  g0647(.A1(new_n841), .A2(new_n842), .A3(new_n845), .A4(new_n847), .ZN(new_n848));
  NOR2_X1   g0648(.A1(new_n770), .A2(new_n221), .ZN(new_n849));
  AOI21_X1  g0649(.A(new_n849), .B1(G311), .B2(new_n798), .ZN(new_n850));
  INV_X1    g0650(.A(G283), .ZN(new_n851));
  OAI22_X1  g0651(.A1(new_n794), .A2(new_n507), .B1(new_n773), .B2(new_n851), .ZN(new_n852));
  AOI211_X1 g0652(.A(new_n297), .B(new_n852), .C1(G294), .C2(new_n792), .ZN(new_n853));
  AOI22_X1  g0653(.A1(new_n786), .A2(G303), .B1(new_n803), .B2(G116), .ZN(new_n854));
  NAND4_X1  g0654(.A1(new_n850), .A2(new_n853), .A3(new_n790), .A4(new_n854), .ZN(new_n855));
  NAND2_X1  g0655(.A1(new_n848), .A2(new_n855), .ZN(new_n856));
  AOI21_X1  g0656(.A(new_n834), .B1(new_n856), .B2(new_n760), .ZN(new_n857));
  OAI21_X1  g0657(.A(new_n857), .B1(new_n825), .B2(new_n758), .ZN(new_n858));
  AND2_X1   g0658(.A1(new_n831), .A2(new_n858), .ZN(new_n859));
  INV_X1    g0659(.A(new_n859), .ZN(G384));
  OAI21_X1  g0660(.A(G77), .B1(new_n224), .B2(new_n226), .ZN(new_n861));
  OAI22_X1  g0661(.A1(new_n861), .A2(new_n217), .B1(G50), .B2(new_n226), .ZN(new_n862));
  NAND3_X1  g0662(.A1(new_n862), .A2(G1), .A3(new_n675), .ZN(new_n863));
  XNOR2_X1  g0663(.A(new_n512), .B(KEYINPUT103), .ZN(new_n864));
  INV_X1    g0664(.A(new_n864), .ZN(new_n865));
  OR2_X1    g0665(.A1(new_n865), .A2(KEYINPUT35), .ZN(new_n866));
  NAND3_X1  g0666(.A1(new_n866), .A2(G116), .A3(new_n215), .ZN(new_n867));
  AOI21_X1  g0667(.A(new_n867), .B1(KEYINPUT35), .B2(new_n865), .ZN(new_n868));
  OAI21_X1  g0668(.A(new_n863), .B1(new_n868), .B2(KEYINPUT36), .ZN(new_n869));
  AOI21_X1  g0669(.A(new_n869), .B1(KEYINPUT36), .B2(new_n868), .ZN(new_n870));
  NOR2_X1   g0670(.A1(new_n460), .A2(new_n682), .ZN(new_n871));
  XNOR2_X1  g0671(.A(new_n871), .B(KEYINPUT104), .ZN(new_n872));
  INV_X1    g0672(.A(new_n872), .ZN(new_n873));
  AOI21_X1  g0673(.A(new_n873), .B1(new_n709), .B2(new_n825), .ZN(new_n874));
  INV_X1    g0674(.A(new_n874), .ZN(new_n875));
  INV_X1    g0675(.A(KEYINPUT38), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n387), .A2(new_n376), .ZN(new_n877));
  INV_X1    g0677(.A(KEYINPUT107), .ZN(new_n878));
  INV_X1    g0678(.A(new_n680), .ZN(new_n879));
  NAND3_X1  g0679(.A1(new_n380), .A2(new_n878), .A3(new_n879), .ZN(new_n880));
  INV_X1    g0680(.A(new_n375), .ZN(new_n881));
  INV_X1    g0681(.A(KEYINPUT77), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n882), .A2(new_n289), .ZN(new_n883));
  NAND2_X1  g0683(.A1(KEYINPUT77), .A2(KEYINPUT3), .ZN(new_n884));
  AOI21_X1  g0684(.A(new_n250), .B1(new_n883), .B2(new_n884), .ZN(new_n885));
  OAI21_X1  g0685(.A(new_n214), .B1(new_n885), .B2(new_n295), .ZN(new_n886));
  AOI21_X1  g0686(.A(new_n226), .B1(new_n886), .B2(KEYINPUT7), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n365), .A2(new_n353), .ZN(new_n888));
  AOI21_X1  g0688(.A(new_n362), .B1(new_n887), .B2(new_n888), .ZN(new_n889));
  AOI21_X1  g0689(.A(new_n267), .B1(new_n889), .B2(KEYINPUT16), .ZN(new_n890));
  AOI21_X1  g0690(.A(new_n881), .B1(new_n890), .B2(new_n363), .ZN(new_n891));
  OAI21_X1  g0691(.A(KEYINPUT107), .B1(new_n891), .B2(new_n680), .ZN(new_n892));
  AOI21_X1  g0692(.A(new_n877), .B1(new_n880), .B2(new_n892), .ZN(new_n893));
  XNOR2_X1  g0693(.A(KEYINPUT108), .B(KEYINPUT37), .ZN(new_n894));
  INV_X1    g0694(.A(new_n894), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n370), .A2(new_n263), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n886), .A2(KEYINPUT7), .ZN(new_n897));
  NAND3_X1  g0697(.A1(new_n897), .A2(new_n888), .A3(G68), .ZN(new_n898));
  AOI21_X1  g0698(.A(KEYINPUT16), .B1(new_n898), .B2(new_n364), .ZN(new_n899));
  OAI21_X1  g0699(.A(new_n375), .B1(new_n896), .B2(new_n899), .ZN(new_n900));
  AOI22_X1  g0700(.A1(new_n891), .A2(new_n351), .B1(new_n900), .B2(new_n383), .ZN(new_n901));
  INV_X1    g0701(.A(KEYINPUT106), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n898), .A2(new_n364), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n903), .A2(new_n352), .ZN(new_n904));
  AOI21_X1  g0704(.A(new_n881), .B1(new_n890), .B2(new_n904), .ZN(new_n905));
  OAI21_X1  g0705(.A(new_n902), .B1(new_n905), .B2(new_n680), .ZN(new_n906));
  NAND3_X1  g0706(.A1(new_n900), .A2(KEYINPUT106), .A3(new_n879), .ZN(new_n907));
  NAND3_X1  g0707(.A1(new_n901), .A2(new_n906), .A3(new_n907), .ZN(new_n908));
  AOI22_X1  g0708(.A1(new_n893), .A2(new_n895), .B1(new_n908), .B2(KEYINPUT37), .ZN(new_n909));
  AOI22_X1  g0709(.A1(new_n386), .A2(new_n391), .B1(new_n906), .B2(new_n907), .ZN(new_n910));
  OAI21_X1  g0710(.A(new_n876), .B1(new_n909), .B2(new_n910), .ZN(new_n911));
  INV_X1    g0711(.A(new_n877), .ZN(new_n912));
  INV_X1    g0712(.A(new_n880), .ZN(new_n913));
  AOI21_X1  g0713(.A(new_n878), .B1(new_n380), .B2(new_n879), .ZN(new_n914));
  OAI211_X1 g0714(.A(new_n912), .B(new_n895), .C1(new_n913), .C2(new_n914), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n908), .A2(KEYINPUT37), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n915), .A2(new_n916), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n906), .A2(new_n907), .ZN(new_n918));
  AND3_X1   g0718(.A1(new_n389), .A2(KEYINPUT78), .A3(new_n390), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n384), .A2(new_n385), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n640), .A2(new_n920), .ZN(new_n921));
  OAI21_X1  g0721(.A(new_n918), .B1(new_n919), .B2(new_n921), .ZN(new_n922));
  NAND3_X1  g0722(.A1(new_n917), .A2(new_n922), .A3(KEYINPUT38), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n911), .A2(new_n923), .ZN(new_n924));
  NOR2_X1   g0724(.A1(new_n427), .A2(new_n683), .ZN(new_n925));
  XNOR2_X1  g0725(.A(new_n925), .B(KEYINPUT105), .ZN(new_n926));
  AND3_X1   g0726(.A1(new_n432), .A2(new_n440), .A3(new_n926), .ZN(new_n927));
  AOI21_X1  g0727(.A(new_n926), .B1(new_n432), .B2(new_n440), .ZN(new_n928));
  NOR2_X1   g0728(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  NAND3_X1  g0729(.A1(new_n875), .A2(new_n924), .A3(new_n929), .ZN(new_n930));
  OAI21_X1  g0730(.A(new_n930), .B1(new_n649), .B2(new_n879), .ZN(new_n931));
  NOR2_X1   g0731(.A1(new_n913), .A2(new_n914), .ZN(new_n932));
  OAI21_X1  g0732(.A(new_n894), .B1(new_n932), .B2(new_n877), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n649), .A2(new_n640), .ZN(new_n934));
  AOI22_X1  g0734(.A1(new_n933), .A2(new_n915), .B1(new_n934), .B2(new_n932), .ZN(new_n935));
  OAI21_X1  g0735(.A(new_n923), .B1(new_n935), .B2(KEYINPUT38), .ZN(new_n936));
  NOR2_X1   g0736(.A1(new_n936), .A2(KEYINPUT39), .ZN(new_n937));
  INV_X1    g0737(.A(KEYINPUT39), .ZN(new_n938));
  AOI21_X1  g0738(.A(new_n938), .B1(new_n911), .B2(new_n923), .ZN(new_n939));
  NOR2_X1   g0739(.A1(new_n937), .A2(new_n939), .ZN(new_n940));
  NOR2_X1   g0740(.A1(new_n440), .A2(new_n682), .ZN(new_n941));
  INV_X1    g0741(.A(new_n941), .ZN(new_n942));
  NOR2_X1   g0742(.A1(new_n940), .A2(new_n942), .ZN(new_n943));
  NOR2_X1   g0743(.A1(new_n931), .A2(new_n943), .ZN(new_n944));
  NAND4_X1  g0744(.A1(new_n711), .A2(new_n466), .A3(new_n712), .A4(new_n722), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n945), .A2(new_n651), .ZN(new_n946));
  XNOR2_X1  g0746(.A(new_n944), .B(new_n946), .ZN(new_n947));
  NOR3_X1   g0747(.A1(new_n927), .A2(new_n928), .A3(new_n824), .ZN(new_n948));
  NAND4_X1  g0748(.A1(new_n936), .A2(new_n743), .A3(KEYINPUT40), .A4(new_n948), .ZN(new_n949));
  NAND3_X1  g0749(.A1(new_n743), .A2(new_n924), .A3(new_n948), .ZN(new_n950));
  INV_X1    g0750(.A(KEYINPUT109), .ZN(new_n951));
  INV_X1    g0751(.A(KEYINPUT40), .ZN(new_n952));
  AND3_X1   g0752(.A1(new_n950), .A2(new_n951), .A3(new_n952), .ZN(new_n953));
  AOI21_X1  g0753(.A(new_n951), .B1(new_n950), .B2(new_n952), .ZN(new_n954));
  OAI211_X1 g0754(.A(G330), .B(new_n949), .C1(new_n953), .C2(new_n954), .ZN(new_n955));
  INV_X1    g0755(.A(new_n744), .ZN(new_n956));
  NAND2_X1  g0756(.A1(new_n956), .A2(new_n466), .ZN(new_n957));
  INV_X1    g0757(.A(new_n949), .ZN(new_n958));
  NAND2_X1  g0758(.A1(new_n950), .A2(new_n952), .ZN(new_n959));
  NAND2_X1  g0759(.A1(new_n959), .A2(KEYINPUT109), .ZN(new_n960));
  NAND3_X1  g0760(.A1(new_n950), .A2(new_n951), .A3(new_n952), .ZN(new_n961));
  AOI21_X1  g0761(.A(new_n958), .B1(new_n960), .B2(new_n961), .ZN(new_n962));
  AND2_X1   g0762(.A1(new_n466), .A2(new_n743), .ZN(new_n963));
  AOI22_X1  g0763(.A1(new_n955), .A2(new_n957), .B1(new_n962), .B2(new_n963), .ZN(new_n964));
  NAND2_X1  g0764(.A1(new_n947), .A2(new_n964), .ZN(new_n965));
  OAI21_X1  g0765(.A(new_n965), .B1(new_n265), .B2(new_n676), .ZN(new_n966));
  OAI22_X1  g0766(.A1(new_n966), .A2(KEYINPUT110), .B1(new_n947), .B2(new_n964), .ZN(new_n967));
  AND2_X1   g0767(.A1(new_n966), .A2(KEYINPUT110), .ZN(new_n968));
  OAI21_X1  g0768(.A(new_n870), .B1(new_n967), .B2(new_n968), .ZN(G367));
  OR2_X1    g0769(.A1(new_n683), .A2(new_n604), .ZN(new_n970));
  NAND2_X1  g0770(.A1(new_n663), .A2(new_n970), .ZN(new_n971));
  OR2_X1    g0771(.A1(new_n659), .A2(new_n970), .ZN(new_n972));
  NAND2_X1  g0772(.A1(new_n971), .A2(new_n972), .ZN(new_n973));
  INV_X1    g0773(.A(new_n973), .ZN(new_n974));
  NAND2_X1  g0774(.A1(new_n974), .A2(new_n759), .ZN(new_n975));
  INV_X1    g0775(.A(new_n751), .ZN(new_n976));
  OAI221_X1 g0776(.A(new_n761), .B1(new_n208), .B2(new_n445), .C1(new_n976), .C2(new_n238), .ZN(new_n977));
  NAND2_X1  g0777(.A1(new_n977), .A2(new_n765), .ZN(new_n978));
  INV_X1    g0778(.A(G317), .ZN(new_n979));
  OAI22_X1  g0779(.A1(new_n782), .A2(new_n851), .B1(new_n777), .B2(new_n979), .ZN(new_n980));
  NOR2_X1   g0780(.A1(new_n770), .A2(new_n502), .ZN(new_n981));
  AOI211_X1 g0781(.A(new_n980), .B(new_n981), .C1(G294), .C2(new_n774), .ZN(new_n982));
  NOR2_X1   g0782(.A1(new_n794), .A2(new_n241), .ZN(new_n983));
  XNOR2_X1  g0783(.A(new_n983), .B(KEYINPUT46), .ZN(new_n984));
  AOI21_X1  g0784(.A(new_n984), .B1(G107), .B2(new_n789), .ZN(new_n985));
  AOI22_X1  g0785(.A1(G311), .A2(new_n786), .B1(new_n792), .B2(G303), .ZN(new_n986));
  NAND4_X1  g0786(.A1(new_n982), .A2(new_n846), .A3(new_n985), .A4(new_n986), .ZN(new_n987));
  INV_X1    g0787(.A(G137), .ZN(new_n988));
  OAI22_X1  g0788(.A1(new_n794), .A2(new_n224), .B1(new_n777), .B2(new_n988), .ZN(new_n989));
  AOI211_X1 g0789(.A(new_n291), .B(new_n989), .C1(G77), .C2(new_n769), .ZN(new_n990));
  AOI22_X1  g0790(.A1(G150), .A2(new_n792), .B1(new_n803), .B2(G50), .ZN(new_n991));
  AOI22_X1  g0791(.A1(G143), .A2(new_n786), .B1(new_n774), .B2(G159), .ZN(new_n992));
  NAND2_X1  g0792(.A1(new_n789), .A2(G68), .ZN(new_n993));
  NAND4_X1  g0793(.A1(new_n990), .A2(new_n991), .A3(new_n992), .A4(new_n993), .ZN(new_n994));
  AOI21_X1  g0794(.A(KEYINPUT47), .B1(new_n987), .B2(new_n994), .ZN(new_n995));
  INV_X1    g0795(.A(new_n760), .ZN(new_n996));
  NOR2_X1   g0796(.A1(new_n995), .A2(new_n996), .ZN(new_n997));
  NAND3_X1  g0797(.A1(new_n987), .A2(KEYINPUT47), .A3(new_n994), .ZN(new_n998));
  AOI21_X1  g0798(.A(new_n978), .B1(new_n997), .B2(new_n998), .ZN(new_n999));
  NAND2_X1  g0799(.A1(new_n975), .A2(new_n999), .ZN(new_n1000));
  NAND2_X1  g0800(.A1(new_n699), .A2(new_n700), .ZN(new_n1001));
  AOI21_X1  g0801(.A(new_n1001), .B1(new_n697), .B2(new_n693), .ZN(new_n1002));
  OAI21_X1  g0802(.A(new_n529), .B1(new_n518), .B2(new_n683), .ZN(new_n1003));
  NAND2_X1  g0803(.A1(new_n519), .A2(new_n682), .ZN(new_n1004));
  NAND2_X1  g0804(.A1(new_n1003), .A2(new_n1004), .ZN(new_n1005));
  NOR2_X1   g0805(.A1(new_n701), .A2(new_n1005), .ZN(new_n1006));
  XNOR2_X1  g0806(.A(new_n1006), .B(KEYINPUT44), .ZN(new_n1007));
  NAND2_X1  g0807(.A1(new_n701), .A2(new_n1005), .ZN(new_n1008));
  INV_X1    g0808(.A(KEYINPUT45), .ZN(new_n1009));
  XNOR2_X1  g0809(.A(new_n1008), .B(new_n1009), .ZN(new_n1010));
  NAND2_X1  g0810(.A1(new_n1007), .A2(new_n1010), .ZN(new_n1011));
  OAI211_X1 g0811(.A(new_n746), .B(new_n1002), .C1(new_n1011), .C2(new_n698), .ZN(new_n1012));
  NAND2_X1  g0812(.A1(new_n1012), .A2(new_n746), .ZN(new_n1013));
  XNOR2_X1  g0813(.A(new_n703), .B(KEYINPUT41), .ZN(new_n1014));
  AOI21_X1  g0814(.A(new_n764), .B1(new_n1013), .B2(new_n1014), .ZN(new_n1015));
  NAND3_X1  g0815(.A1(new_n691), .A2(new_n692), .A3(new_n1005), .ZN(new_n1016));
  OAI21_X1  g0816(.A(new_n668), .B1(new_n1003), .B2(new_n578), .ZN(new_n1017));
  AOI22_X1  g0817(.A1(new_n1016), .A2(KEYINPUT42), .B1(new_n683), .B2(new_n1017), .ZN(new_n1018));
  OAI21_X1  g0818(.A(new_n1018), .B1(KEYINPUT42), .B2(new_n1016), .ZN(new_n1019));
  INV_X1    g0819(.A(KEYINPUT43), .ZN(new_n1020));
  OAI21_X1  g0820(.A(new_n1019), .B1(new_n1020), .B2(new_n974), .ZN(new_n1021));
  NAND2_X1  g0821(.A1(new_n974), .A2(new_n1020), .ZN(new_n1022));
  XNOR2_X1  g0822(.A(new_n1021), .B(new_n1022), .ZN(new_n1023));
  INV_X1    g0823(.A(new_n1005), .ZN(new_n1024));
  NOR2_X1   g0824(.A1(new_n699), .A2(new_n1024), .ZN(new_n1025));
  XNOR2_X1  g0825(.A(new_n1023), .B(new_n1025), .ZN(new_n1026));
  OAI21_X1  g0826(.A(new_n1000), .B1(new_n1015), .B2(new_n1026), .ZN(G387));
  NAND2_X1  g0827(.A1(new_n1002), .A2(new_n764), .ZN(new_n1028));
  OAI211_X1 g0828(.A(new_n705), .B(new_n278), .C1(new_n226), .C2(new_n294), .ZN(new_n1029));
  NAND2_X1  g0829(.A1(new_n443), .A2(new_n202), .ZN(new_n1030));
  AOI21_X1  g0830(.A(new_n1029), .B1(new_n1030), .B2(KEYINPUT50), .ZN(new_n1031));
  OAI21_X1  g0831(.A(new_n1031), .B1(KEYINPUT50), .B2(new_n1030), .ZN(new_n1032));
  OAI211_X1 g0832(.A(new_n1032), .B(new_n751), .C1(new_n235), .C2(new_n278), .ZN(new_n1033));
  INV_X1    g0833(.A(new_n748), .ZN(new_n1034));
  OAI22_X1  g0834(.A1(new_n1034), .A2(new_n705), .B1(G107), .B2(new_n208), .ZN(new_n1035));
  XOR2_X1   g0835(.A(new_n1035), .B(KEYINPUT111), .Z(new_n1036));
  NAND3_X1  g0836(.A1(new_n1033), .A2(new_n1036), .A3(KEYINPUT112), .ZN(new_n1037));
  NAND2_X1  g0837(.A1(new_n1037), .A2(new_n761), .ZN(new_n1038));
  AOI21_X1  g0838(.A(KEYINPUT112), .B1(new_n1033), .B2(new_n1036), .ZN(new_n1039));
  OAI21_X1  g0839(.A(new_n765), .B1(new_n1038), .B2(new_n1039), .ZN(new_n1040));
  INV_X1    g0840(.A(new_n596), .ZN(new_n1041));
  NOR2_X1   g0841(.A1(new_n1041), .A2(new_n807), .ZN(new_n1042));
  AOI21_X1  g0842(.A(new_n1042), .B1(new_n372), .B2(new_n774), .ZN(new_n1043));
  OAI22_X1  g0843(.A1(new_n785), .A2(new_n778), .B1(new_n791), .B2(new_n202), .ZN(new_n1044));
  OAI22_X1  g0844(.A1(new_n782), .A2(new_n226), .B1(new_n777), .B2(new_n838), .ZN(new_n1045));
  NOR2_X1   g0845(.A1(new_n1044), .A2(new_n1045), .ZN(new_n1046));
  AOI21_X1  g0846(.A(new_n981), .B1(G77), .B2(new_n795), .ZN(new_n1047));
  NAND4_X1  g0847(.A1(new_n1043), .A2(new_n368), .A3(new_n1046), .A4(new_n1047), .ZN(new_n1048));
  AOI22_X1  g0848(.A1(new_n786), .A2(G322), .B1(new_n803), .B2(G303), .ZN(new_n1049));
  INV_X1    g0849(.A(G311), .ZN(new_n1050));
  OAI221_X1 g0850(.A(new_n1049), .B1(new_n1050), .B2(new_n773), .C1(new_n979), .C2(new_n791), .ZN(new_n1051));
  XNOR2_X1  g0851(.A(new_n1051), .B(KEYINPUT48), .ZN(new_n1052));
  OAI221_X1 g0852(.A(new_n1052), .B1(new_n851), .B2(new_n807), .C1(new_n806), .C2(new_n794), .ZN(new_n1053));
  XOR2_X1   g0853(.A(new_n1053), .B(KEYINPUT49), .Z(new_n1054));
  AOI22_X1  g0854(.A1(new_n769), .A2(G116), .B1(G326), .B2(new_n798), .ZN(new_n1055));
  NAND2_X1  g0855(.A1(new_n1055), .A2(new_n846), .ZN(new_n1056));
  OAI21_X1  g0856(.A(new_n1048), .B1(new_n1054), .B2(new_n1056), .ZN(new_n1057));
  AOI21_X1  g0857(.A(new_n1040), .B1(new_n1057), .B2(new_n760), .ZN(new_n1058));
  OAI21_X1  g0858(.A(new_n1058), .B1(new_n691), .B2(new_n811), .ZN(new_n1059));
  NAND2_X1  g0859(.A1(new_n746), .A2(new_n1002), .ZN(new_n1060));
  NAND2_X1  g0860(.A1(new_n1060), .A2(new_n703), .ZN(new_n1061));
  NOR2_X1   g0861(.A1(new_n746), .A2(new_n1002), .ZN(new_n1062));
  OAI211_X1 g0862(.A(new_n1028), .B(new_n1059), .C1(new_n1061), .C2(new_n1062), .ZN(G393));
  XNOR2_X1  g0863(.A(new_n1011), .B(new_n698), .ZN(new_n1064));
  NAND2_X1  g0864(.A1(new_n1064), .A2(new_n1060), .ZN(new_n1065));
  NAND2_X1  g0865(.A1(new_n1065), .A2(KEYINPUT113), .ZN(new_n1066));
  INV_X1    g0866(.A(KEYINPUT113), .ZN(new_n1067));
  NAND3_X1  g0867(.A1(new_n1064), .A2(new_n1067), .A3(new_n1060), .ZN(new_n1068));
  NAND4_X1  g0868(.A1(new_n1066), .A2(new_n703), .A3(new_n1012), .A4(new_n1068), .ZN(new_n1069));
  NOR2_X1   g0869(.A1(new_n1064), .A2(new_n763), .ZN(new_n1070));
  AOI211_X1 g0870(.A(new_n297), .B(new_n771), .C1(G116), .C2(new_n789), .ZN(new_n1071));
  OAI22_X1  g0871(.A1(new_n785), .A2(new_n979), .B1(new_n791), .B2(new_n1050), .ZN(new_n1072));
  XNOR2_X1  g0872(.A(new_n1072), .B(KEYINPUT52), .ZN(new_n1073));
  AOI22_X1  g0873(.A1(G294), .A2(new_n803), .B1(new_n798), .B2(G322), .ZN(new_n1074));
  AOI22_X1  g0874(.A1(new_n795), .A2(G283), .B1(new_n774), .B2(G303), .ZN(new_n1075));
  NAND4_X1  g0875(.A1(new_n1071), .A2(new_n1073), .A3(new_n1074), .A4(new_n1075), .ZN(new_n1076));
  AOI211_X1 g0876(.A(new_n846), .B(new_n849), .C1(G68), .C2(new_n795), .ZN(new_n1077));
  OAI22_X1  g0877(.A1(new_n785), .A2(new_n838), .B1(new_n791), .B2(new_n778), .ZN(new_n1078));
  XNOR2_X1  g0878(.A(new_n1078), .B(KEYINPUT51), .ZN(new_n1079));
  NAND2_X1  g0879(.A1(new_n443), .A2(new_n803), .ZN(new_n1080));
  OAI21_X1  g0880(.A(new_n1080), .B1(new_n837), .B2(new_n777), .ZN(new_n1081));
  AOI21_X1  g0881(.A(new_n1081), .B1(G50), .B2(new_n774), .ZN(new_n1082));
  NAND2_X1  g0882(.A1(new_n789), .A2(G77), .ZN(new_n1083));
  NAND4_X1  g0883(.A1(new_n1077), .A2(new_n1079), .A3(new_n1082), .A4(new_n1083), .ZN(new_n1084));
  AOI21_X1  g0884(.A(new_n996), .B1(new_n1076), .B2(new_n1084), .ZN(new_n1085));
  OAI221_X1 g0885(.A(new_n761), .B1(new_n502), .B2(new_n208), .C1(new_n244), .C2(new_n976), .ZN(new_n1086));
  NAND2_X1  g0886(.A1(new_n1086), .A2(new_n765), .ZN(new_n1087));
  AOI211_X1 g0887(.A(new_n1085), .B(new_n1087), .C1(new_n1024), .C2(new_n759), .ZN(new_n1088));
  NOR2_X1   g0888(.A1(new_n1070), .A2(new_n1088), .ZN(new_n1089));
  NAND2_X1  g0889(.A1(new_n1069), .A2(new_n1089), .ZN(G390));
  NAND2_X1  g0890(.A1(new_n940), .A2(new_n757), .ZN(new_n1091));
  OAI21_X1  g0891(.A(new_n765), .B1(new_n833), .B2(new_n372), .ZN(new_n1092));
  NOR2_X1   g0892(.A1(new_n794), .A2(new_n838), .ZN(new_n1093));
  XNOR2_X1  g0893(.A(KEYINPUT118), .B(KEYINPUT53), .ZN(new_n1094));
  XNOR2_X1  g0894(.A(new_n1093), .B(new_n1094), .ZN(new_n1095));
  XOR2_X1   g0895(.A(KEYINPUT54), .B(G143), .Z(new_n1096));
  XNOR2_X1  g0896(.A(new_n1096), .B(KEYINPUT117), .ZN(new_n1097));
  OAI21_X1  g0897(.A(new_n1095), .B1(new_n782), .B2(new_n1097), .ZN(new_n1098));
  AOI22_X1  g0898(.A1(new_n769), .A2(G50), .B1(new_n792), .B2(G132), .ZN(new_n1099));
  AOI22_X1  g0899(.A1(G128), .A2(new_n786), .B1(new_n774), .B2(G137), .ZN(new_n1100));
  NAND2_X1  g0900(.A1(new_n789), .A2(G159), .ZN(new_n1101));
  AOI21_X1  g0901(.A(new_n291), .B1(new_n798), .B2(G125), .ZN(new_n1102));
  NAND4_X1  g0902(.A1(new_n1099), .A2(new_n1100), .A3(new_n1101), .A4(new_n1102), .ZN(new_n1103));
  AOI22_X1  g0903(.A1(new_n786), .A2(G283), .B1(new_n798), .B2(G294), .ZN(new_n1104));
  OAI221_X1 g0904(.A(new_n1104), .B1(new_n502), .B2(new_n782), .C1(new_n507), .C2(new_n773), .ZN(new_n1105));
  AOI21_X1  g0905(.A(new_n297), .B1(new_n795), .B2(G87), .ZN(new_n1106));
  NAND2_X1  g0906(.A1(new_n792), .A2(G116), .ZN(new_n1107));
  NAND4_X1  g0907(.A1(new_n1106), .A2(new_n843), .A3(new_n1083), .A4(new_n1107), .ZN(new_n1108));
  OAI22_X1  g0908(.A1(new_n1098), .A2(new_n1103), .B1(new_n1105), .B2(new_n1108), .ZN(new_n1109));
  AOI21_X1  g0909(.A(new_n1092), .B1(new_n1109), .B2(new_n760), .ZN(new_n1110));
  NAND2_X1  g0910(.A1(new_n1091), .A2(new_n1110), .ZN(new_n1111));
  AND3_X1   g0911(.A1(new_n719), .A2(new_n659), .A3(new_n720), .ZN(new_n1112));
  AOI211_X1 g0912(.A(new_n682), .B(new_n824), .C1(new_n664), .C2(new_n1112), .ZN(new_n1113));
  OAI21_X1  g0913(.A(KEYINPUT114), .B1(new_n1113), .B2(new_n873), .ZN(new_n1114));
  INV_X1    g0914(.A(KEYINPUT114), .ZN(new_n1115));
  OAI21_X1  g0915(.A(new_n683), .B1(new_n717), .B2(new_n721), .ZN(new_n1116));
  OAI211_X1 g0916(.A(new_n1115), .B(new_n872), .C1(new_n1116), .C2(new_n824), .ZN(new_n1117));
  NAND3_X1  g0917(.A1(new_n1114), .A2(new_n929), .A3(new_n1117), .ZN(new_n1118));
  AND2_X1   g0918(.A1(new_n936), .A2(new_n942), .ZN(new_n1119));
  INV_X1    g0919(.A(new_n929), .ZN(new_n1120));
  OAI21_X1  g0920(.A(new_n942), .B1(new_n874), .B2(new_n1120), .ZN(new_n1121));
  AOI22_X1  g0921(.A1(new_n1118), .A2(new_n1119), .B1(new_n940), .B2(new_n1121), .ZN(new_n1122));
  NOR3_X1   g0922(.A1(new_n744), .A2(new_n824), .A3(new_n1120), .ZN(new_n1123));
  AND2_X1   g0923(.A1(new_n1123), .A2(KEYINPUT115), .ZN(new_n1124));
  NOR2_X1   g0924(.A1(new_n1123), .A2(KEYINPUT115), .ZN(new_n1125));
  NOR3_X1   g0925(.A1(new_n1122), .A2(new_n1124), .A3(new_n1125), .ZN(new_n1126));
  NAND2_X1  g0926(.A1(new_n1118), .A2(new_n1119), .ZN(new_n1127));
  NAND2_X1  g0927(.A1(new_n940), .A2(new_n1121), .ZN(new_n1128));
  AND4_X1   g0928(.A1(KEYINPUT115), .A2(new_n1127), .A3(new_n1123), .A4(new_n1128), .ZN(new_n1129));
  NOR2_X1   g0929(.A1(new_n1126), .A2(new_n1129), .ZN(new_n1130));
  OAI21_X1  g0930(.A(new_n1111), .B1(new_n1130), .B2(new_n763), .ZN(new_n1131));
  NAND3_X1  g0931(.A1(new_n945), .A2(new_n957), .A3(new_n651), .ZN(new_n1132));
  AOI21_X1  g0932(.A(new_n929), .B1(new_n956), .B2(new_n825), .ZN(new_n1133));
  OAI21_X1  g0933(.A(new_n875), .B1(new_n1133), .B2(new_n1123), .ZN(new_n1134));
  NAND3_X1  g0934(.A1(new_n956), .A2(new_n825), .A3(new_n929), .ZN(new_n1135));
  NAND2_X1  g0935(.A1(new_n1114), .A2(new_n1117), .ZN(new_n1136));
  OAI21_X1  g0936(.A(new_n1120), .B1(new_n744), .B2(new_n824), .ZN(new_n1137));
  NAND3_X1  g0937(.A1(new_n1135), .A2(new_n1136), .A3(new_n1137), .ZN(new_n1138));
  AOI21_X1  g0938(.A(new_n1132), .B1(new_n1134), .B2(new_n1138), .ZN(new_n1139));
  XNOR2_X1  g0939(.A(new_n1139), .B(KEYINPUT116), .ZN(new_n1140));
  NAND2_X1  g0940(.A1(new_n1140), .A2(new_n1130), .ZN(new_n1141));
  OAI21_X1  g0941(.A(new_n1139), .B1(new_n1126), .B2(new_n1129), .ZN(new_n1142));
  AND2_X1   g0942(.A1(new_n1142), .A2(new_n703), .ZN(new_n1143));
  AOI21_X1  g0943(.A(new_n1131), .B1(new_n1141), .B2(new_n1143), .ZN(new_n1144));
  INV_X1    g0944(.A(new_n1144), .ZN(G378));
  INV_X1    g0945(.A(new_n944), .ZN(new_n1146));
  XNOR2_X1  g0946(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1147));
  INV_X1    g0947(.A(new_n1147), .ZN(new_n1148));
  INV_X1    g0948(.A(KEYINPUT120), .ZN(new_n1149));
  NAND2_X1  g0949(.A1(new_n333), .A2(new_n1149), .ZN(new_n1150));
  NAND2_X1  g0950(.A1(new_n270), .A2(new_n879), .ZN(new_n1151));
  AOI22_X1  g0951(.A1(new_n317), .A2(new_n322), .B1(new_n330), .B2(new_n331), .ZN(new_n1152));
  NAND2_X1  g0952(.A1(new_n1152), .A2(KEYINPUT120), .ZN(new_n1153));
  NAND3_X1  g0953(.A1(new_n1150), .A2(new_n1151), .A3(new_n1153), .ZN(new_n1154));
  INV_X1    g0954(.A(new_n1154), .ZN(new_n1155));
  AOI21_X1  g0955(.A(new_n1151), .B1(new_n1150), .B2(new_n1153), .ZN(new_n1156));
  OAI21_X1  g0956(.A(new_n1148), .B1(new_n1155), .B2(new_n1156), .ZN(new_n1157));
  INV_X1    g0957(.A(new_n1151), .ZN(new_n1158));
  NOR2_X1   g0958(.A1(new_n333), .A2(new_n1149), .ZN(new_n1159));
  NOR2_X1   g0959(.A1(new_n1152), .A2(KEYINPUT120), .ZN(new_n1160));
  OAI21_X1  g0960(.A(new_n1158), .B1(new_n1159), .B2(new_n1160), .ZN(new_n1161));
  NAND3_X1  g0961(.A1(new_n1161), .A2(new_n1147), .A3(new_n1154), .ZN(new_n1162));
  NAND2_X1  g0962(.A1(new_n1157), .A2(new_n1162), .ZN(new_n1163));
  AOI21_X1  g0963(.A(new_n1163), .B1(new_n962), .B2(G330), .ZN(new_n1164));
  NOR3_X1   g0964(.A1(new_n1155), .A2(new_n1156), .A3(new_n1148), .ZN(new_n1165));
  AOI21_X1  g0965(.A(new_n1147), .B1(new_n1161), .B2(new_n1154), .ZN(new_n1166));
  NOR2_X1   g0966(.A1(new_n1165), .A2(new_n1166), .ZN(new_n1167));
  NOR2_X1   g0967(.A1(new_n955), .A2(new_n1167), .ZN(new_n1168));
  OAI21_X1  g0968(.A(new_n1146), .B1(new_n1164), .B2(new_n1168), .ZN(new_n1169));
  INV_X1    g0969(.A(KEYINPUT121), .ZN(new_n1170));
  NAND3_X1  g0970(.A1(new_n962), .A2(G330), .A3(new_n1163), .ZN(new_n1171));
  NAND2_X1  g0971(.A1(new_n955), .A2(new_n1167), .ZN(new_n1172));
  NAND3_X1  g0972(.A1(new_n1171), .A2(new_n1172), .A3(new_n944), .ZN(new_n1173));
  NAND3_X1  g0973(.A1(new_n1169), .A2(new_n1170), .A3(new_n1173), .ZN(new_n1174));
  NAND4_X1  g0974(.A1(new_n1171), .A2(new_n1172), .A3(KEYINPUT121), .A4(new_n944), .ZN(new_n1175));
  INV_X1    g0975(.A(new_n1132), .ZN(new_n1176));
  NAND2_X1  g0976(.A1(new_n1142), .A2(new_n1176), .ZN(new_n1177));
  NAND3_X1  g0977(.A1(new_n1174), .A2(new_n1175), .A3(new_n1177), .ZN(new_n1178));
  INV_X1    g0978(.A(KEYINPUT57), .ZN(new_n1179));
  NAND2_X1  g0979(.A1(new_n1178), .A2(new_n1179), .ZN(new_n1180));
  AOI21_X1  g0980(.A(new_n1179), .B1(new_n1142), .B2(new_n1176), .ZN(new_n1181));
  NAND2_X1  g0981(.A1(new_n1169), .A2(new_n1173), .ZN(new_n1182));
  AOI21_X1  g0982(.A(new_n704), .B1(new_n1181), .B2(new_n1182), .ZN(new_n1183));
  NAND2_X1  g0983(.A1(new_n1180), .A2(new_n1183), .ZN(new_n1184));
  NAND3_X1  g0984(.A1(new_n1174), .A2(new_n764), .A3(new_n1175), .ZN(new_n1185));
  NOR2_X1   g0985(.A1(new_n1163), .A2(new_n758), .ZN(new_n1186));
  AOI22_X1  g0986(.A1(G125), .A2(new_n786), .B1(new_n774), .B2(G132), .ZN(new_n1187));
  AOI22_X1  g0987(.A1(G128), .A2(new_n792), .B1(new_n803), .B2(G137), .ZN(new_n1188));
  AND2_X1   g0988(.A1(new_n1187), .A2(new_n1188), .ZN(new_n1189));
  OAI221_X1 g0989(.A(new_n1189), .B1(new_n838), .B2(new_n807), .C1(new_n794), .C2(new_n1097), .ZN(new_n1190));
  NAND2_X1  g0990(.A1(new_n1190), .A2(KEYINPUT59), .ZN(new_n1191));
  NAND2_X1  g0991(.A1(new_n769), .A2(G159), .ZN(new_n1192));
  AOI211_X1 g0992(.A(G33), .B(G41), .C1(new_n798), .C2(G124), .ZN(new_n1193));
  NAND3_X1  g0993(.A1(new_n1191), .A2(new_n1192), .A3(new_n1193), .ZN(new_n1194));
  NOR2_X1   g0994(.A1(new_n1190), .A2(KEYINPUT59), .ZN(new_n1195));
  NOR2_X1   g0995(.A1(new_n1194), .A2(new_n1195), .ZN(new_n1196));
  NOR2_X1   g0996(.A1(new_n368), .A2(G41), .ZN(new_n1197));
  AOI211_X1 g0997(.A(G50), .B(new_n1197), .C1(new_n250), .C2(new_n277), .ZN(new_n1198));
  OAI22_X1  g0998(.A1(new_n770), .A2(new_n224), .B1(new_n777), .B2(new_n851), .ZN(new_n1199));
  OAI221_X1 g0999(.A(new_n993), .B1(new_n294), .B2(new_n794), .C1(new_n507), .C2(new_n791), .ZN(new_n1200));
  OAI22_X1  g1000(.A1(new_n785), .A2(new_n241), .B1(new_n773), .B2(new_n502), .ZN(new_n1201));
  NOR3_X1   g1001(.A1(new_n1199), .A2(new_n1200), .A3(new_n1201), .ZN(new_n1202));
  OAI211_X1 g1002(.A(new_n1202), .B(new_n1197), .C1(new_n1041), .C2(new_n782), .ZN(new_n1203));
  INV_X1    g1003(.A(KEYINPUT58), .ZN(new_n1204));
  AOI21_X1  g1004(.A(new_n1198), .B1(new_n1203), .B2(new_n1204), .ZN(new_n1205));
  OAI21_X1  g1005(.A(new_n1205), .B1(new_n1204), .B2(new_n1203), .ZN(new_n1206));
  OAI21_X1  g1006(.A(new_n760), .B1(new_n1196), .B2(new_n1206), .ZN(new_n1207));
  XNOR2_X1  g1007(.A(new_n1207), .B(KEYINPUT119), .ZN(new_n1208));
  NAND2_X1  g1008(.A1(new_n832), .A2(new_n202), .ZN(new_n1209));
  NAND3_X1  g1009(.A1(new_n1208), .A2(new_n765), .A3(new_n1209), .ZN(new_n1210));
  NOR2_X1   g1010(.A1(new_n1186), .A2(new_n1210), .ZN(new_n1211));
  INV_X1    g1011(.A(new_n1211), .ZN(new_n1212));
  AND2_X1   g1012(.A1(new_n1185), .A2(new_n1212), .ZN(new_n1213));
  NAND2_X1  g1013(.A1(new_n1184), .A2(new_n1213), .ZN(G375));
  NAND3_X1  g1014(.A1(new_n1134), .A2(new_n1132), .A3(new_n1138), .ZN(new_n1215));
  NAND3_X1  g1015(.A1(new_n1140), .A2(new_n1014), .A3(new_n1215), .ZN(new_n1216));
  OAI221_X1 g1016(.A(new_n368), .B1(new_n988), .B2(new_n791), .C1(new_n770), .C2(new_n224), .ZN(new_n1217));
  AOI22_X1  g1017(.A1(new_n795), .A2(G159), .B1(new_n786), .B2(G132), .ZN(new_n1218));
  AOI22_X1  g1018(.A1(G150), .A2(new_n803), .B1(new_n798), .B2(G128), .ZN(new_n1219));
  OAI211_X1 g1019(.A(new_n1218), .B(new_n1219), .C1(new_n1097), .C2(new_n773), .ZN(new_n1220));
  AOI211_X1 g1020(.A(new_n1217), .B(new_n1220), .C1(G50), .C2(new_n789), .ZN(new_n1221));
  AOI22_X1  g1021(.A1(new_n786), .A2(G294), .B1(new_n798), .B2(G303), .ZN(new_n1222));
  OAI221_X1 g1022(.A(new_n1222), .B1(new_n502), .B2(new_n794), .C1(new_n241), .C2(new_n773), .ZN(new_n1223));
  AOI22_X1  g1023(.A1(G283), .A2(new_n792), .B1(new_n803), .B2(G107), .ZN(new_n1224));
  OAI211_X1 g1024(.A(new_n1224), .B(new_n291), .C1(new_n294), .C2(new_n770), .ZN(new_n1225));
  NOR3_X1   g1025(.A1(new_n1223), .A2(new_n1225), .A3(new_n1042), .ZN(new_n1226));
  OAI21_X1  g1026(.A(new_n760), .B1(new_n1221), .B2(new_n1226), .ZN(new_n1227));
  OAI211_X1 g1027(.A(new_n1227), .B(new_n765), .C1(G68), .C2(new_n833), .ZN(new_n1228));
  AOI21_X1  g1028(.A(new_n1228), .B1(new_n1120), .B2(new_n757), .ZN(new_n1229));
  NAND2_X1  g1029(.A1(new_n1134), .A2(new_n1138), .ZN(new_n1230));
  AOI21_X1  g1030(.A(new_n1229), .B1(new_n1230), .B2(new_n764), .ZN(new_n1231));
  NAND2_X1  g1031(.A1(new_n1216), .A2(new_n1231), .ZN(G381));
  OR4_X1    g1032(.A1(G396), .A2(G390), .A3(G384), .A4(G393), .ZN(new_n1233));
  NOR2_X1   g1033(.A1(G375), .A2(G378), .ZN(new_n1234));
  INV_X1    g1034(.A(new_n1234), .ZN(new_n1235));
  OR4_X1    g1035(.A1(G387), .A2(new_n1233), .A3(G381), .A4(new_n1235), .ZN(G407));
  NAND2_X1  g1036(.A1(new_n681), .A2(G213), .ZN(new_n1237));
  XOR2_X1   g1037(.A(new_n1237), .B(KEYINPUT122), .Z(new_n1238));
  OAI211_X1 g1038(.A(G407), .B(G213), .C1(new_n1235), .C2(new_n1238), .ZN(G409));
  NAND3_X1  g1039(.A1(new_n1184), .A2(G378), .A3(new_n1213), .ZN(new_n1240));
  NAND4_X1  g1040(.A1(new_n1174), .A2(new_n1177), .A3(new_n1014), .A4(new_n1175), .ZN(new_n1241));
  AOI21_X1  g1041(.A(new_n1211), .B1(new_n1182), .B2(new_n764), .ZN(new_n1242));
  NAND2_X1  g1042(.A1(new_n1241), .A2(new_n1242), .ZN(new_n1243));
  AND3_X1   g1043(.A1(new_n1243), .A2(new_n1144), .A3(KEYINPUT123), .ZN(new_n1244));
  AOI21_X1  g1044(.A(KEYINPUT123), .B1(new_n1243), .B2(new_n1144), .ZN(new_n1245));
  OAI21_X1  g1045(.A(new_n1240), .B1(new_n1244), .B2(new_n1245), .ZN(new_n1246));
  AND2_X1   g1046(.A1(new_n1246), .A2(new_n1238), .ZN(new_n1247));
  INV_X1    g1047(.A(KEYINPUT60), .ZN(new_n1248));
  OR2_X1    g1048(.A1(new_n1215), .A2(new_n1248), .ZN(new_n1249));
  NAND2_X1  g1049(.A1(new_n1215), .A2(new_n1248), .ZN(new_n1250));
  NOR2_X1   g1050(.A1(new_n1139), .A2(new_n704), .ZN(new_n1251));
  NAND3_X1  g1051(.A1(new_n1249), .A2(new_n1250), .A3(new_n1251), .ZN(new_n1252));
  AND3_X1   g1052(.A1(new_n1252), .A2(G384), .A3(new_n1231), .ZN(new_n1253));
  AOI21_X1  g1053(.A(G384), .B1(new_n1252), .B2(new_n1231), .ZN(new_n1254));
  NOR2_X1   g1054(.A1(new_n1253), .A2(new_n1254), .ZN(new_n1255));
  NAND3_X1  g1055(.A1(new_n1247), .A2(KEYINPUT63), .A3(new_n1255), .ZN(new_n1256));
  XOR2_X1   g1056(.A(G393), .B(G396), .Z(new_n1257));
  INV_X1    g1057(.A(new_n1257), .ZN(new_n1258));
  NAND3_X1  g1058(.A1(new_n1069), .A2(G387), .A3(new_n1089), .ZN(new_n1259));
  INV_X1    g1059(.A(new_n1259), .ZN(new_n1260));
  AOI21_X1  g1060(.A(G387), .B1(new_n1069), .B2(new_n1089), .ZN(new_n1261));
  OAI21_X1  g1061(.A(new_n1258), .B1(new_n1260), .B2(new_n1261), .ZN(new_n1262));
  INV_X1    g1062(.A(new_n1261), .ZN(new_n1263));
  NAND3_X1  g1063(.A1(new_n1263), .A2(new_n1257), .A3(new_n1259), .ZN(new_n1264));
  NAND2_X1  g1064(.A1(new_n1262), .A2(new_n1264), .ZN(new_n1265));
  NOR2_X1   g1065(.A1(new_n1265), .A2(KEYINPUT61), .ZN(new_n1266));
  INV_X1    g1066(.A(KEYINPUT63), .ZN(new_n1267));
  INV_X1    g1067(.A(G2897), .ZN(new_n1268));
  OR2_X1    g1068(.A1(new_n1238), .A2(new_n1268), .ZN(new_n1269));
  NOR2_X1   g1069(.A1(new_n1255), .A2(new_n1269), .ZN(new_n1270));
  INV_X1    g1070(.A(KEYINPUT124), .ZN(new_n1271));
  NOR2_X1   g1071(.A1(new_n1237), .A2(new_n1268), .ZN(new_n1272));
  NOR3_X1   g1072(.A1(new_n1253), .A2(new_n1254), .A3(new_n1272), .ZN(new_n1273));
  OR3_X1    g1073(.A1(new_n1270), .A2(new_n1271), .A3(new_n1273), .ZN(new_n1274));
  OAI21_X1  g1074(.A(new_n1271), .B1(new_n1270), .B2(new_n1273), .ZN(new_n1275));
  AND2_X1   g1075(.A1(new_n1274), .A2(new_n1275), .ZN(new_n1276));
  NAND2_X1  g1076(.A1(new_n1246), .A2(new_n1237), .ZN(new_n1277));
  AOI21_X1  g1077(.A(new_n1267), .B1(new_n1276), .B2(new_n1277), .ZN(new_n1278));
  NAND3_X1  g1078(.A1(new_n1246), .A2(new_n1237), .A3(new_n1255), .ZN(new_n1279));
  INV_X1    g1079(.A(new_n1279), .ZN(new_n1280));
  OAI211_X1 g1080(.A(new_n1256), .B(new_n1266), .C1(new_n1278), .C2(new_n1280), .ZN(new_n1281));
  XOR2_X1   g1081(.A(KEYINPUT125), .B(KEYINPUT61), .Z(new_n1282));
  NAND2_X1  g1082(.A1(new_n1274), .A2(new_n1275), .ZN(new_n1283));
  OAI21_X1  g1083(.A(new_n1282), .B1(new_n1283), .B2(new_n1247), .ZN(new_n1284));
  INV_X1    g1084(.A(new_n1255), .ZN(new_n1285));
  INV_X1    g1085(.A(KEYINPUT62), .ZN(new_n1286));
  NOR2_X1   g1086(.A1(new_n1285), .A2(new_n1286), .ZN(new_n1287));
  AND3_X1   g1087(.A1(new_n1246), .A2(new_n1238), .A3(new_n1287), .ZN(new_n1288));
  NAND2_X1  g1088(.A1(new_n1279), .A2(new_n1286), .ZN(new_n1289));
  AOI21_X1  g1089(.A(new_n1288), .B1(new_n1289), .B2(KEYINPUT126), .ZN(new_n1290));
  INV_X1    g1090(.A(KEYINPUT126), .ZN(new_n1291));
  NAND3_X1  g1091(.A1(new_n1279), .A2(new_n1291), .A3(new_n1286), .ZN(new_n1292));
  AOI21_X1  g1092(.A(new_n1284), .B1(new_n1290), .B2(new_n1292), .ZN(new_n1293));
  INV_X1    g1093(.A(new_n1265), .ZN(new_n1294));
  OAI21_X1  g1094(.A(new_n1281), .B1(new_n1293), .B2(new_n1294), .ZN(G405));
  OR2_X1    g1095(.A1(new_n1265), .A2(KEYINPUT127), .ZN(new_n1296));
  NAND2_X1  g1096(.A1(G375), .A2(new_n1144), .ZN(new_n1297));
  NAND2_X1  g1097(.A1(new_n1297), .A2(new_n1240), .ZN(new_n1298));
  XNOR2_X1  g1098(.A(new_n1298), .B(new_n1285), .ZN(new_n1299));
  NAND2_X1  g1099(.A1(new_n1265), .A2(KEYINPUT127), .ZN(new_n1300));
  NAND3_X1  g1100(.A1(new_n1296), .A2(new_n1299), .A3(new_n1300), .ZN(new_n1301));
  OAI21_X1  g1101(.A(new_n1301), .B1(new_n1299), .B2(new_n1300), .ZN(G402));
endmodule


