

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300,
         n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311,
         n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322,
         n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333,
         n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344,
         n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355,
         n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
         n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
         n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
         n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
         n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410,
         n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421,
         n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432,
         n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443,
         n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454,
         n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465,
         n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
         n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487,
         n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
         n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
         n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586;

  XNOR2_X1 U322 ( .A(G99GAT), .B(G106GAT), .ZN(n343) );
  XNOR2_X1 U323 ( .A(n367), .B(n366), .ZN(n368) );
  XNOR2_X1 U324 ( .A(n449), .B(KEYINPUT116), .ZN(n562) );
  XNOR2_X1 U325 ( .A(n359), .B(n358), .ZN(n556) );
  XNOR2_X1 U326 ( .A(n355), .B(n354), .ZN(n359) );
  XOR2_X1 U327 ( .A(n292), .B(n447), .Z(n530) );
  XNOR2_X2 U328 ( .A(n339), .B(n338), .ZN(n574) );
  XNOR2_X1 U329 ( .A(G176GAT), .B(KEYINPUT117), .ZN(n290) );
  AND2_X1 U330 ( .A1(G227GAT), .A2(G233GAT), .ZN(n291) );
  XNOR2_X1 U331 ( .A(n446), .B(n445), .ZN(n292) );
  INV_X1 U332 ( .A(KEYINPUT107), .ZN(n366) );
  XNOR2_X1 U333 ( .A(n440), .B(n291), .ZN(n441) );
  INV_X1 U334 ( .A(KEYINPUT93), .ZN(n474) );
  XNOR2_X1 U335 ( .A(n442), .B(n441), .ZN(n444) );
  XNOR2_X1 U336 ( .A(n475), .B(n474), .ZN(n476) );
  XNOR2_X1 U337 ( .A(n390), .B(KEYINPUT115), .ZN(n391) );
  NAND2_X1 U338 ( .A1(n477), .A2(n476), .ZN(n490) );
  XOR2_X1 U339 ( .A(G120GAT), .B(G71GAT), .Z(n434) );
  XNOR2_X1 U340 ( .A(n357), .B(n356), .ZN(n358) );
  NOR2_X1 U341 ( .A1(n583), .A2(n491), .ZN(n492) );
  XOR2_X1 U342 ( .A(KEYINPUT36), .B(n541), .Z(n583) );
  XOR2_X1 U343 ( .A(n469), .B(KEYINPUT26), .Z(n570) );
  XNOR2_X1 U344 ( .A(KEYINPUT38), .B(n494), .ZN(n502) );
  XNOR2_X1 U345 ( .A(n450), .B(G190GAT), .ZN(n451) );
  XNOR2_X1 U346 ( .A(n452), .B(n451), .ZN(G1351GAT) );
  XOR2_X1 U347 ( .A(G78GAT), .B(G71GAT), .Z(n294) );
  XNOR2_X1 U348 ( .A(G22GAT), .B(G127GAT), .ZN(n293) );
  XNOR2_X1 U349 ( .A(n294), .B(n293), .ZN(n308) );
  XOR2_X1 U350 ( .A(KEYINPUT13), .B(G57GAT), .Z(n328) );
  XOR2_X1 U351 ( .A(n328), .B(G211GAT), .Z(n297) );
  XNOR2_X1 U352 ( .A(G15GAT), .B(G1GAT), .ZN(n295) );
  XNOR2_X1 U353 ( .A(n295), .B(KEYINPUT70), .ZN(n318) );
  XNOR2_X1 U354 ( .A(n318), .B(G155GAT), .ZN(n296) );
  XNOR2_X1 U355 ( .A(n297), .B(n296), .ZN(n301) );
  XOR2_X1 U356 ( .A(KEYINPUT12), .B(G64GAT), .Z(n299) );
  NAND2_X1 U357 ( .A1(G231GAT), .A2(G233GAT), .ZN(n298) );
  XNOR2_X1 U358 ( .A(n299), .B(n298), .ZN(n300) );
  XOR2_X1 U359 ( .A(n301), .B(n300), .Z(n306) );
  XOR2_X1 U360 ( .A(KEYINPUT15), .B(KEYINPUT14), .Z(n303) );
  XNOR2_X1 U361 ( .A(G8GAT), .B(G183GAT), .ZN(n302) );
  XNOR2_X1 U362 ( .A(n303), .B(n302), .ZN(n304) );
  XNOR2_X1 U363 ( .A(n304), .B(KEYINPUT77), .ZN(n305) );
  XNOR2_X1 U364 ( .A(n306), .B(n305), .ZN(n307) );
  XOR2_X1 U365 ( .A(n308), .B(n307), .Z(n579) );
  INV_X1 U366 ( .A(n579), .ZN(n561) );
  XOR2_X1 U367 ( .A(KEYINPUT29), .B(KEYINPUT30), .Z(n310) );
  XNOR2_X1 U368 ( .A(KEYINPUT69), .B(KEYINPUT67), .ZN(n309) );
  XNOR2_X1 U369 ( .A(n310), .B(n309), .ZN(n314) );
  XOR2_X1 U370 ( .A(G113GAT), .B(G197GAT), .Z(n312) );
  XOR2_X1 U371 ( .A(G141GAT), .B(G22GAT), .Z(n405) );
  XOR2_X1 U372 ( .A(G169GAT), .B(G8GAT), .Z(n375) );
  XNOR2_X1 U373 ( .A(n405), .B(n375), .ZN(n311) );
  XNOR2_X1 U374 ( .A(n312), .B(n311), .ZN(n313) );
  XOR2_X1 U375 ( .A(n314), .B(n313), .Z(n316) );
  NAND2_X1 U376 ( .A1(G229GAT), .A2(G233GAT), .ZN(n315) );
  XNOR2_X1 U377 ( .A(n316), .B(n315), .ZN(n317) );
  XOR2_X1 U378 ( .A(n317), .B(KEYINPUT66), .Z(n320) );
  XNOR2_X1 U379 ( .A(n318), .B(KEYINPUT68), .ZN(n319) );
  XNOR2_X1 U380 ( .A(n320), .B(n319), .ZN(n325) );
  XOR2_X1 U381 ( .A(G29GAT), .B(KEYINPUT8), .Z(n322) );
  XNOR2_X1 U382 ( .A(G43GAT), .B(G36GAT), .ZN(n321) );
  XNOR2_X1 U383 ( .A(n322), .B(n321), .ZN(n324) );
  XOR2_X1 U384 ( .A(G50GAT), .B(KEYINPUT7), .Z(n323) );
  XNOR2_X1 U385 ( .A(n324), .B(n323), .ZN(n357) );
  XNOR2_X1 U386 ( .A(n325), .B(n357), .ZN(n571) );
  XOR2_X1 U387 ( .A(G85GAT), .B(G92GAT), .Z(n344) );
  XNOR2_X1 U388 ( .A(n344), .B(n343), .ZN(n326) );
  XNOR2_X1 U389 ( .A(n326), .B(KEYINPUT31), .ZN(n327) );
  XNOR2_X1 U390 ( .A(n327), .B(KEYINPUT73), .ZN(n331) );
  XNOR2_X1 U391 ( .A(n328), .B(KEYINPUT33), .ZN(n329) );
  XNOR2_X1 U392 ( .A(n329), .B(KEYINPUT32), .ZN(n330) );
  XNOR2_X1 U393 ( .A(n331), .B(n330), .ZN(n336) );
  XOR2_X1 U394 ( .A(G78GAT), .B(G148GAT), .Z(n333) );
  XNOR2_X1 U395 ( .A(KEYINPUT72), .B(G204GAT), .ZN(n332) );
  XNOR2_X1 U396 ( .A(n333), .B(n332), .ZN(n402) );
  XNOR2_X1 U397 ( .A(G176GAT), .B(G64GAT), .ZN(n334) );
  XNOR2_X1 U398 ( .A(n334), .B(KEYINPUT74), .ZN(n376) );
  XNOR2_X1 U399 ( .A(n402), .B(n376), .ZN(n335) );
  XNOR2_X1 U400 ( .A(n336), .B(n335), .ZN(n337) );
  XNOR2_X1 U401 ( .A(n434), .B(n337), .ZN(n339) );
  NAND2_X1 U402 ( .A1(G230GAT), .A2(G233GAT), .ZN(n338) );
  INV_X1 U403 ( .A(KEYINPUT41), .ZN(n340) );
  XNOR2_X1 U404 ( .A(n574), .B(n340), .ZN(n550) );
  NOR2_X1 U405 ( .A1(n571), .A2(n550), .ZN(n341) );
  XNOR2_X1 U406 ( .A(n341), .B(KEYINPUT46), .ZN(n342) );
  NOR2_X1 U407 ( .A1(n561), .A2(n342), .ZN(n360) );
  XNOR2_X1 U408 ( .A(n343), .B(KEYINPUT64), .ZN(n345) );
  XNOR2_X1 U409 ( .A(n345), .B(n344), .ZN(n349) );
  INV_X1 U410 ( .A(n349), .ZN(n347) );
  AND2_X1 U411 ( .A1(G232GAT), .A2(G233GAT), .ZN(n348) );
  INV_X1 U412 ( .A(n348), .ZN(n346) );
  NAND2_X1 U413 ( .A1(n347), .A2(n346), .ZN(n351) );
  NAND2_X1 U414 ( .A1(n349), .A2(n348), .ZN(n350) );
  NAND2_X1 U415 ( .A1(n351), .A2(n350), .ZN(n355) );
  XOR2_X1 U416 ( .A(KEYINPUT10), .B(KEYINPUT11), .Z(n353) );
  XNOR2_X1 U417 ( .A(KEYINPUT9), .B(KEYINPUT75), .ZN(n352) );
  XOR2_X1 U418 ( .A(n353), .B(n352), .Z(n354) );
  XOR2_X1 U419 ( .A(G190GAT), .B(G134GAT), .Z(n435) );
  XOR2_X1 U420 ( .A(G218GAT), .B(G162GAT), .Z(n404) );
  XNOR2_X1 U421 ( .A(n435), .B(n404), .ZN(n356) );
  NAND2_X1 U422 ( .A1(n360), .A2(n556), .ZN(n361) );
  XNOR2_X1 U423 ( .A(n361), .B(KEYINPUT106), .ZN(n362) );
  XNOR2_X1 U424 ( .A(KEYINPUT47), .B(n362), .ZN(n371) );
  XNOR2_X1 U425 ( .A(KEYINPUT71), .B(n571), .ZN(n559) );
  INV_X1 U426 ( .A(KEYINPUT76), .ZN(n363) );
  XNOR2_X1 U427 ( .A(n556), .B(n363), .ZN(n541) );
  NOR2_X1 U428 ( .A1(n579), .A2(n583), .ZN(n364) );
  XNOR2_X1 U429 ( .A(n364), .B(KEYINPUT45), .ZN(n365) );
  NAND2_X1 U430 ( .A1(n365), .A2(n574), .ZN(n367) );
  NOR2_X1 U431 ( .A1(n559), .A2(n368), .ZN(n369) );
  XNOR2_X1 U432 ( .A(n369), .B(KEYINPUT108), .ZN(n370) );
  NOR2_X1 U433 ( .A1(n371), .A2(n370), .ZN(n372) );
  XNOR2_X1 U434 ( .A(n372), .B(KEYINPUT48), .ZN(n528) );
  XOR2_X1 U435 ( .A(G92GAT), .B(G218GAT), .Z(n374) );
  XNOR2_X1 U436 ( .A(G36GAT), .B(G190GAT), .ZN(n373) );
  XNOR2_X1 U437 ( .A(n374), .B(n373), .ZN(n385) );
  XOR2_X1 U438 ( .A(n376), .B(n375), .Z(n378) );
  NAND2_X1 U439 ( .A1(G226GAT), .A2(G233GAT), .ZN(n377) );
  XNOR2_X1 U440 ( .A(n378), .B(n377), .ZN(n379) );
  XOR2_X1 U441 ( .A(n379), .B(KEYINPUT90), .Z(n383) );
  XOR2_X1 U442 ( .A(G211GAT), .B(KEYINPUT84), .Z(n381) );
  XNOR2_X1 U443 ( .A(G197GAT), .B(KEYINPUT21), .ZN(n380) );
  XNOR2_X1 U444 ( .A(n381), .B(n380), .ZN(n399) );
  XNOR2_X1 U445 ( .A(n399), .B(G204GAT), .ZN(n382) );
  XNOR2_X1 U446 ( .A(n383), .B(n382), .ZN(n384) );
  XNOR2_X1 U447 ( .A(n385), .B(n384), .ZN(n389) );
  XOR2_X1 U448 ( .A(KEYINPUT19), .B(KEYINPUT18), .Z(n387) );
  XNOR2_X1 U449 ( .A(KEYINPUT81), .B(G183GAT), .ZN(n386) );
  XNOR2_X1 U450 ( .A(n387), .B(n386), .ZN(n388) );
  XNOR2_X1 U451 ( .A(KEYINPUT17), .B(n388), .ZN(n447) );
  XOR2_X1 U452 ( .A(n389), .B(n447), .Z(n521) );
  INV_X1 U453 ( .A(n521), .ZN(n463) );
  NOR2_X1 U454 ( .A1(n528), .A2(n463), .ZN(n392) );
  INV_X1 U455 ( .A(KEYINPUT54), .ZN(n390) );
  XNOR2_X1 U456 ( .A(n392), .B(n391), .ZN(n568) );
  XOR2_X1 U457 ( .A(KEYINPUT24), .B(KEYINPUT22), .Z(n394) );
  XNOR2_X1 U458 ( .A(G50GAT), .B(G106GAT), .ZN(n393) );
  XNOR2_X1 U459 ( .A(n394), .B(n393), .ZN(n409) );
  XOR2_X1 U460 ( .A(KEYINPUT83), .B(KEYINPUT23), .Z(n396) );
  NAND2_X1 U461 ( .A1(G228GAT), .A2(G233GAT), .ZN(n395) );
  XNOR2_X1 U462 ( .A(n396), .B(n395), .ZN(n397) );
  XOR2_X1 U463 ( .A(n397), .B(KEYINPUT85), .Z(n401) );
  XNOR2_X1 U464 ( .A(G155GAT), .B(KEYINPUT2), .ZN(n398) );
  XNOR2_X1 U465 ( .A(n398), .B(KEYINPUT3), .ZN(n425) );
  XNOR2_X1 U466 ( .A(n425), .B(n399), .ZN(n400) );
  XNOR2_X1 U467 ( .A(n401), .B(n400), .ZN(n403) );
  XOR2_X1 U468 ( .A(n403), .B(n402), .Z(n407) );
  XNOR2_X1 U469 ( .A(n405), .B(n404), .ZN(n406) );
  XNOR2_X1 U470 ( .A(n407), .B(n406), .ZN(n408) );
  XNOR2_X1 U471 ( .A(n409), .B(n408), .ZN(n468) );
  XOR2_X1 U472 ( .A(G148GAT), .B(G120GAT), .Z(n411) );
  XNOR2_X1 U473 ( .A(G1GAT), .B(G141GAT), .ZN(n410) );
  XNOR2_X1 U474 ( .A(n411), .B(n410), .ZN(n415) );
  XOR2_X1 U475 ( .A(KEYINPUT1), .B(KEYINPUT6), .Z(n413) );
  XNOR2_X1 U476 ( .A(G57GAT), .B(KEYINPUT86), .ZN(n412) );
  XNOR2_X1 U477 ( .A(n413), .B(n412), .ZN(n414) );
  XOR2_X1 U478 ( .A(n415), .B(n414), .Z(n422) );
  XOR2_X1 U479 ( .A(G127GAT), .B(KEYINPUT0), .Z(n417) );
  XNOR2_X1 U480 ( .A(G113GAT), .B(KEYINPUT79), .ZN(n416) );
  XNOR2_X1 U481 ( .A(n417), .B(n416), .ZN(n443) );
  XOR2_X1 U482 ( .A(G85GAT), .B(G162GAT), .Z(n419) );
  XNOR2_X1 U483 ( .A(G29GAT), .B(G134GAT), .ZN(n418) );
  XNOR2_X1 U484 ( .A(n419), .B(n418), .ZN(n420) );
  XNOR2_X1 U485 ( .A(n443), .B(n420), .ZN(n421) );
  XNOR2_X1 U486 ( .A(n422), .B(n421), .ZN(n431) );
  XOR2_X1 U487 ( .A(KEYINPUT89), .B(KEYINPUT4), .Z(n424) );
  XNOR2_X1 U488 ( .A(KEYINPUT87), .B(KEYINPUT5), .ZN(n423) );
  XNOR2_X1 U489 ( .A(n424), .B(n423), .ZN(n429) );
  XOR2_X1 U490 ( .A(n425), .B(KEYINPUT88), .Z(n427) );
  NAND2_X1 U491 ( .A1(G225GAT), .A2(G233GAT), .ZN(n426) );
  XNOR2_X1 U492 ( .A(n427), .B(n426), .ZN(n428) );
  XOR2_X1 U493 ( .A(n429), .B(n428), .Z(n430) );
  XOR2_X1 U494 ( .A(n431), .B(n430), .Z(n519) );
  NOR2_X1 U495 ( .A1(n468), .A2(n519), .ZN(n432) );
  AND2_X1 U496 ( .A1(n568), .A2(n432), .ZN(n433) );
  XNOR2_X1 U497 ( .A(n433), .B(KEYINPUT55), .ZN(n448) );
  XOR2_X1 U498 ( .A(G99GAT), .B(n434), .Z(n437) );
  XNOR2_X1 U499 ( .A(G43GAT), .B(n435), .ZN(n436) );
  XNOR2_X1 U500 ( .A(n437), .B(n436), .ZN(n442) );
  XOR2_X1 U501 ( .A(KEYINPUT20), .B(KEYINPUT80), .Z(n439) );
  XNOR2_X1 U502 ( .A(G176GAT), .B(KEYINPUT82), .ZN(n438) );
  XNOR2_X1 U503 ( .A(n439), .B(n438), .ZN(n440) );
  XOR2_X1 U504 ( .A(n444), .B(n443), .Z(n446) );
  XNOR2_X1 U505 ( .A(G169GAT), .B(G15GAT), .ZN(n445) );
  INV_X1 U506 ( .A(n530), .ZN(n467) );
  NOR2_X1 U507 ( .A1(n448), .A2(n467), .ZN(n449) );
  NAND2_X1 U508 ( .A1(n562), .A2(n541), .ZN(n452) );
  XOR2_X1 U509 ( .A(KEYINPUT58), .B(KEYINPUT121), .Z(n450) );
  INV_X1 U510 ( .A(n550), .ZN(n535) );
  NAND2_X1 U511 ( .A1(n562), .A2(n535), .ZN(n457) );
  XOR2_X1 U512 ( .A(KEYINPUT119), .B(KEYINPUT118), .Z(n454) );
  XNOR2_X1 U513 ( .A(KEYINPUT56), .B(KEYINPUT57), .ZN(n453) );
  XNOR2_X1 U514 ( .A(n454), .B(n453), .ZN(n455) );
  XNOR2_X1 U515 ( .A(n455), .B(n290), .ZN(n456) );
  XNOR2_X1 U516 ( .A(n457), .B(n456), .ZN(G1349GAT) );
  XOR2_X1 U517 ( .A(KEYINPUT78), .B(KEYINPUT16), .Z(n459) );
  OR2_X1 U518 ( .A1(n541), .A2(n579), .ZN(n458) );
  XNOR2_X1 U519 ( .A(n459), .B(n458), .ZN(n478) );
  XOR2_X1 U520 ( .A(KEYINPUT65), .B(KEYINPUT28), .Z(n460) );
  XNOR2_X1 U521 ( .A(n468), .B(n460), .ZN(n533) );
  XNOR2_X1 U522 ( .A(KEYINPUT27), .B(n521), .ZN(n470) );
  NAND2_X1 U523 ( .A1(n519), .A2(n470), .ZN(n529) );
  NOR2_X1 U524 ( .A1(n533), .A2(n529), .ZN(n461) );
  NAND2_X1 U525 ( .A1(n467), .A2(n461), .ZN(n462) );
  XOR2_X1 U526 ( .A(KEYINPUT91), .B(n462), .Z(n477) );
  INV_X1 U527 ( .A(n519), .ZN(n567) );
  XNOR2_X1 U528 ( .A(KEYINPUT92), .B(KEYINPUT25), .ZN(n466) );
  NOR2_X1 U529 ( .A1(n467), .A2(n463), .ZN(n464) );
  NOR2_X1 U530 ( .A1(n468), .A2(n464), .ZN(n465) );
  XNOR2_X1 U531 ( .A(n466), .B(n465), .ZN(n472) );
  NAND2_X1 U532 ( .A1(n468), .A2(n467), .ZN(n469) );
  NAND2_X1 U533 ( .A1(n570), .A2(n470), .ZN(n471) );
  NAND2_X1 U534 ( .A1(n472), .A2(n471), .ZN(n473) );
  NAND2_X1 U535 ( .A1(n567), .A2(n473), .ZN(n475) );
  NAND2_X1 U536 ( .A1(n478), .A2(n490), .ZN(n505) );
  NAND2_X1 U537 ( .A1(n574), .A2(n559), .ZN(n493) );
  NOR2_X1 U538 ( .A1(n505), .A2(n493), .ZN(n479) );
  XNOR2_X1 U539 ( .A(n479), .B(KEYINPUT94), .ZN(n488) );
  NAND2_X1 U540 ( .A1(n488), .A2(n519), .ZN(n483) );
  XOR2_X1 U541 ( .A(KEYINPUT34), .B(KEYINPUT95), .Z(n481) );
  XNOR2_X1 U542 ( .A(G1GAT), .B(KEYINPUT96), .ZN(n480) );
  XNOR2_X1 U543 ( .A(n481), .B(n480), .ZN(n482) );
  XNOR2_X1 U544 ( .A(n483), .B(n482), .ZN(G1324GAT) );
  XOR2_X1 U545 ( .A(G8GAT), .B(KEYINPUT97), .Z(n485) );
  NAND2_X1 U546 ( .A1(n521), .A2(n488), .ZN(n484) );
  XNOR2_X1 U547 ( .A(n485), .B(n484), .ZN(G1325GAT) );
  XOR2_X1 U548 ( .A(G15GAT), .B(KEYINPUT35), .Z(n487) );
  NAND2_X1 U549 ( .A1(n488), .A2(n530), .ZN(n486) );
  XNOR2_X1 U550 ( .A(n487), .B(n486), .ZN(G1326GAT) );
  NAND2_X1 U551 ( .A1(n488), .A2(n533), .ZN(n489) );
  XNOR2_X1 U552 ( .A(n489), .B(G22GAT), .ZN(G1327GAT) );
  XOR2_X1 U553 ( .A(KEYINPUT98), .B(KEYINPUT39), .Z(n496) );
  NAND2_X1 U554 ( .A1(n579), .A2(n490), .ZN(n491) );
  XNOR2_X1 U555 ( .A(KEYINPUT37), .B(n492), .ZN(n518) );
  NOR2_X1 U556 ( .A1(n518), .A2(n493), .ZN(n494) );
  NAND2_X1 U557 ( .A1(n519), .A2(n502), .ZN(n495) );
  XNOR2_X1 U558 ( .A(n496), .B(n495), .ZN(n497) );
  XNOR2_X1 U559 ( .A(G29GAT), .B(n497), .ZN(G1328GAT) );
  NAND2_X1 U560 ( .A1(n521), .A2(n502), .ZN(n498) );
  XNOR2_X1 U561 ( .A(G36GAT), .B(n498), .ZN(G1329GAT) );
  XOR2_X1 U562 ( .A(KEYINPUT40), .B(KEYINPUT99), .Z(n500) );
  NAND2_X1 U563 ( .A1(n502), .A2(n530), .ZN(n499) );
  XNOR2_X1 U564 ( .A(n500), .B(n499), .ZN(n501) );
  XNOR2_X1 U565 ( .A(G43GAT), .B(n501), .ZN(G1330GAT) );
  NAND2_X1 U566 ( .A1(n502), .A2(n533), .ZN(n503) );
  XNOR2_X1 U567 ( .A(n503), .B(KEYINPUT100), .ZN(n504) );
  XNOR2_X1 U568 ( .A(G50GAT), .B(n504), .ZN(G1331GAT) );
  XNOR2_X1 U569 ( .A(G57GAT), .B(KEYINPUT42), .ZN(n508) );
  NAND2_X1 U570 ( .A1(n571), .A2(n535), .ZN(n517) );
  NOR2_X1 U571 ( .A1(n505), .A2(n517), .ZN(n506) );
  XOR2_X1 U572 ( .A(KEYINPUT101), .B(n506), .Z(n512) );
  NAND2_X1 U573 ( .A1(n519), .A2(n512), .ZN(n507) );
  XNOR2_X1 U574 ( .A(n508), .B(n507), .ZN(G1332GAT) );
  NAND2_X1 U575 ( .A1(n512), .A2(n521), .ZN(n509) );
  XNOR2_X1 U576 ( .A(n509), .B(G64GAT), .ZN(G1333GAT) );
  NAND2_X1 U577 ( .A1(n530), .A2(n512), .ZN(n510) );
  XNOR2_X1 U578 ( .A(n510), .B(KEYINPUT102), .ZN(n511) );
  XNOR2_X1 U579 ( .A(G71GAT), .B(n511), .ZN(G1334GAT) );
  XOR2_X1 U580 ( .A(KEYINPUT104), .B(KEYINPUT43), .Z(n514) );
  NAND2_X1 U581 ( .A1(n512), .A2(n533), .ZN(n513) );
  XNOR2_X1 U582 ( .A(n514), .B(n513), .ZN(n516) );
  XOR2_X1 U583 ( .A(G78GAT), .B(KEYINPUT103), .Z(n515) );
  XNOR2_X1 U584 ( .A(n516), .B(n515), .ZN(G1335GAT) );
  NOR2_X1 U585 ( .A1(n518), .A2(n517), .ZN(n524) );
  NAND2_X1 U586 ( .A1(n519), .A2(n524), .ZN(n520) );
  XNOR2_X1 U587 ( .A(G85GAT), .B(n520), .ZN(G1336GAT) );
  NAND2_X1 U588 ( .A1(n524), .A2(n521), .ZN(n522) );
  XNOR2_X1 U589 ( .A(n522), .B(G92GAT), .ZN(G1337GAT) );
  NAND2_X1 U590 ( .A1(n530), .A2(n524), .ZN(n523) );
  XNOR2_X1 U591 ( .A(n523), .B(G99GAT), .ZN(G1338GAT) );
  XOR2_X1 U592 ( .A(KEYINPUT105), .B(KEYINPUT44), .Z(n526) );
  NAND2_X1 U593 ( .A1(n524), .A2(n533), .ZN(n525) );
  XNOR2_X1 U594 ( .A(n526), .B(n525), .ZN(n527) );
  XNOR2_X1 U595 ( .A(G106GAT), .B(n527), .ZN(G1339GAT) );
  NOR2_X1 U596 ( .A1(n528), .A2(n529), .ZN(n546) );
  NAND2_X1 U597 ( .A1(n546), .A2(n530), .ZN(n531) );
  XOR2_X1 U598 ( .A(KEYINPUT109), .B(n531), .Z(n532) );
  NOR2_X1 U599 ( .A1(n533), .A2(n532), .ZN(n542) );
  NAND2_X1 U600 ( .A1(n559), .A2(n542), .ZN(n534) );
  XNOR2_X1 U601 ( .A(n534), .B(G113GAT), .ZN(G1340GAT) );
  XOR2_X1 U602 ( .A(G120GAT), .B(KEYINPUT49), .Z(n537) );
  NAND2_X1 U603 ( .A1(n542), .A2(n535), .ZN(n536) );
  XNOR2_X1 U604 ( .A(n537), .B(n536), .ZN(G1341GAT) );
  XOR2_X1 U605 ( .A(KEYINPUT50), .B(KEYINPUT110), .Z(n539) );
  NAND2_X1 U606 ( .A1(n542), .A2(n561), .ZN(n538) );
  XNOR2_X1 U607 ( .A(n539), .B(n538), .ZN(n540) );
  XOR2_X1 U608 ( .A(G127GAT), .B(n540), .Z(G1342GAT) );
  XOR2_X1 U609 ( .A(KEYINPUT51), .B(KEYINPUT111), .Z(n544) );
  NAND2_X1 U610 ( .A1(n542), .A2(n541), .ZN(n543) );
  XNOR2_X1 U611 ( .A(n544), .B(n543), .ZN(n545) );
  XOR2_X1 U612 ( .A(G134GAT), .B(n545), .Z(G1343GAT) );
  NAND2_X1 U613 ( .A1(n546), .A2(n570), .ZN(n555) );
  NOR2_X1 U614 ( .A1(n571), .A2(n555), .ZN(n547) );
  XOR2_X1 U615 ( .A(G141GAT), .B(n547), .Z(G1344GAT) );
  XOR2_X1 U616 ( .A(KEYINPUT53), .B(KEYINPUT52), .Z(n549) );
  XNOR2_X1 U617 ( .A(G148GAT), .B(KEYINPUT112), .ZN(n548) );
  XNOR2_X1 U618 ( .A(n549), .B(n548), .ZN(n552) );
  NOR2_X1 U619 ( .A1(n550), .A2(n555), .ZN(n551) );
  XOR2_X1 U620 ( .A(n552), .B(n551), .Z(G1345GAT) );
  NOR2_X1 U621 ( .A1(n579), .A2(n555), .ZN(n554) );
  XNOR2_X1 U622 ( .A(G155GAT), .B(KEYINPUT113), .ZN(n553) );
  XNOR2_X1 U623 ( .A(n554), .B(n553), .ZN(G1346GAT) );
  NOR2_X1 U624 ( .A1(n556), .A2(n555), .ZN(n557) );
  XOR2_X1 U625 ( .A(KEYINPUT114), .B(n557), .Z(n558) );
  XNOR2_X1 U626 ( .A(G162GAT), .B(n558), .ZN(G1347GAT) );
  NAND2_X1 U627 ( .A1(n559), .A2(n562), .ZN(n560) );
  XNOR2_X1 U628 ( .A(G169GAT), .B(n560), .ZN(G1348GAT) );
  NAND2_X1 U629 ( .A1(n562), .A2(n561), .ZN(n563) );
  XNOR2_X1 U630 ( .A(n563), .B(KEYINPUT120), .ZN(n564) );
  XNOR2_X1 U631 ( .A(G183GAT), .B(n564), .ZN(G1350GAT) );
  XOR2_X1 U632 ( .A(KEYINPUT60), .B(KEYINPUT59), .Z(n566) );
  XNOR2_X1 U633 ( .A(G197GAT), .B(KEYINPUT122), .ZN(n565) );
  XNOR2_X1 U634 ( .A(n566), .B(n565), .ZN(n573) );
  AND2_X1 U635 ( .A1(n568), .A2(n567), .ZN(n569) );
  NAND2_X1 U636 ( .A1(n570), .A2(n569), .ZN(n582) );
  NOR2_X1 U637 ( .A1(n571), .A2(n582), .ZN(n572) );
  XOR2_X1 U638 ( .A(n573), .B(n572), .Z(G1352GAT) );
  NOR2_X1 U639 ( .A1(n582), .A2(n574), .ZN(n578) );
  XOR2_X1 U640 ( .A(KEYINPUT123), .B(KEYINPUT124), .Z(n576) );
  XNOR2_X1 U641 ( .A(G204GAT), .B(KEYINPUT61), .ZN(n575) );
  XNOR2_X1 U642 ( .A(n576), .B(n575), .ZN(n577) );
  XNOR2_X1 U643 ( .A(n578), .B(n577), .ZN(G1353GAT) );
  NOR2_X1 U644 ( .A1(n579), .A2(n582), .ZN(n581) );
  XNOR2_X1 U645 ( .A(G211GAT), .B(KEYINPUT125), .ZN(n580) );
  XNOR2_X1 U646 ( .A(n581), .B(n580), .ZN(G1354GAT) );
  NOR2_X1 U647 ( .A1(n583), .A2(n582), .ZN(n585) );
  XNOR2_X1 U648 ( .A(KEYINPUT62), .B(KEYINPUT126), .ZN(n584) );
  XNOR2_X1 U649 ( .A(n585), .B(n584), .ZN(n586) );
  XOR2_X1 U650 ( .A(G218GAT), .B(n586), .Z(G1355GAT) );
endmodule

