//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 1 1 1 0 0 0 1 0 0 1 0 1 1 0 1 1 1 0 1 1 0 1 0 0 1 0 1 0 0 0 0 0 0 1 1 0 0 0 0 1 0 0 0 1 0 1 0 0 0 0 0 1 0 0 1 0 1 0 0 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:36:03 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1186, new_n1187, new_n1188, new_n1189, new_n1190, new_n1191,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1251, new_n1252,
    new_n1253, new_n1254, new_n1255, new_n1256, new_n1257, new_n1258,
    new_n1259, new_n1260, new_n1262, new_n1263, new_n1264, new_n1265,
    new_n1266, new_n1267, new_n1268, new_n1269, new_n1270, new_n1271,
    new_n1272, new_n1273, new_n1274, new_n1275, new_n1276, new_n1277,
    new_n1278, new_n1279, new_n1280, new_n1281, new_n1282, new_n1283,
    new_n1285, new_n1286, new_n1287, new_n1288, new_n1289, new_n1290,
    new_n1291, new_n1292, new_n1293, new_n1295, new_n1296, new_n1297,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1346,
    new_n1347, new_n1348, new_n1349, new_n1350, new_n1351, new_n1353,
    new_n1354, new_n1355, new_n1356, new_n1357, new_n1358, new_n1359,
    new_n1360, new_n1361;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(new_n201), .ZN(new_n202));
  NOR3_X1   g0002(.A1(new_n202), .A2(G50), .A3(G77), .ZN(G353));
  OAI21_X1  g0003(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0004(.A1(G1), .A2(G20), .ZN(new_n205));
  AOI22_X1  g0005(.A1(G68), .A2(G238), .B1(G87), .B2(G250), .ZN(new_n206));
  INV_X1    g0006(.A(G50), .ZN(new_n207));
  INV_X1    g0007(.A(G226), .ZN(new_n208));
  INV_X1    g0008(.A(G116), .ZN(new_n209));
  INV_X1    g0009(.A(G270), .ZN(new_n210));
  OAI221_X1 g0010(.A(new_n206), .B1(new_n207), .B2(new_n208), .C1(new_n209), .C2(new_n210), .ZN(new_n211));
  AOI22_X1  g0011(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n212));
  INV_X1    g0012(.A(G58), .ZN(new_n213));
  INV_X1    g0013(.A(G232), .ZN(new_n214));
  INV_X1    g0014(.A(G97), .ZN(new_n215));
  INV_X1    g0015(.A(G257), .ZN(new_n216));
  OAI221_X1 g0016(.A(new_n212), .B1(new_n213), .B2(new_n214), .C1(new_n215), .C2(new_n216), .ZN(new_n217));
  OAI21_X1  g0017(.A(new_n205), .B1(new_n211), .B2(new_n217), .ZN(new_n218));
  XNOR2_X1  g0018(.A(new_n218), .B(KEYINPUT1), .ZN(new_n219));
  OR3_X1    g0019(.A1(new_n205), .A2(KEYINPUT64), .A3(G13), .ZN(new_n220));
  OAI21_X1  g0020(.A(KEYINPUT64), .B1(new_n205), .B2(G13), .ZN(new_n221));
  NAND2_X1  g0021(.A1(new_n220), .A2(new_n221), .ZN(new_n222));
  OAI211_X1 g0022(.A(new_n222), .B(G250), .C1(G257), .C2(G264), .ZN(new_n223));
  XOR2_X1   g0023(.A(new_n223), .B(KEYINPUT0), .Z(new_n224));
  NAND2_X1  g0024(.A1(G1), .A2(G13), .ZN(new_n225));
  INV_X1    g0025(.A(G20), .ZN(new_n226));
  NOR2_X1   g0026(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  NAND2_X1  g0027(.A1(new_n202), .A2(G50), .ZN(new_n228));
  INV_X1    g0028(.A(new_n228), .ZN(new_n229));
  AOI211_X1 g0029(.A(new_n219), .B(new_n224), .C1(new_n227), .C2(new_n229), .ZN(G361));
  XNOR2_X1  g0030(.A(G238), .B(G244), .ZN(new_n231));
  XNOR2_X1  g0031(.A(new_n231), .B(G232), .ZN(new_n232));
  XNOR2_X1  g0032(.A(KEYINPUT2), .B(G226), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n232), .B(new_n233), .ZN(new_n234));
  XOR2_X1   g0034(.A(G264), .B(G270), .Z(new_n235));
  XNOR2_X1  g0035(.A(G250), .B(G257), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n234), .B(new_n237), .ZN(G358));
  XOR2_X1   g0038(.A(G87), .B(G97), .Z(new_n239));
  XNOR2_X1  g0039(.A(G107), .B(G116), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  NAND2_X1  g0041(.A1(new_n207), .A2(G68), .ZN(new_n242));
  INV_X1    g0042(.A(G68), .ZN(new_n243));
  NAND2_X1  g0043(.A1(new_n243), .A2(G50), .ZN(new_n244));
  NAND2_X1  g0044(.A1(new_n242), .A2(new_n244), .ZN(new_n245));
  XNOR2_X1  g0045(.A(G58), .B(G77), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n245), .B(new_n246), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n241), .B(new_n247), .ZN(G351));
  INV_X1    g0048(.A(G1), .ZN(new_n249));
  NAND3_X1  g0049(.A1(new_n249), .A2(G13), .A3(G20), .ZN(new_n250));
  INV_X1    g0050(.A(new_n250), .ZN(new_n251));
  NAND2_X1  g0051(.A1(new_n251), .A2(new_n207), .ZN(new_n252));
  NAND3_X1  g0052(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n253));
  NAND3_X1  g0053(.A1(new_n250), .A2(new_n225), .A3(new_n253), .ZN(new_n254));
  NAND2_X1  g0054(.A1(new_n249), .A2(G20), .ZN(new_n255));
  NAND2_X1  g0055(.A1(new_n255), .A2(G50), .ZN(new_n256));
  AOI21_X1  g0056(.A(new_n226), .B1(new_n201), .B2(new_n207), .ZN(new_n257));
  NOR2_X1   g0057(.A1(G20), .A2(G33), .ZN(new_n258));
  INV_X1    g0058(.A(new_n258), .ZN(new_n259));
  INV_X1    g0059(.A(G150), .ZN(new_n260));
  NOR2_X1   g0060(.A1(new_n259), .A2(new_n260), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n213), .A2(KEYINPUT8), .ZN(new_n262));
  INV_X1    g0062(.A(KEYINPUT8), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n263), .A2(G58), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n262), .A2(new_n264), .ZN(new_n265));
  INV_X1    g0065(.A(G33), .ZN(new_n266));
  NOR2_X1   g0066(.A1(new_n266), .A2(G20), .ZN(new_n267));
  AOI211_X1 g0067(.A(new_n257), .B(new_n261), .C1(new_n265), .C2(new_n267), .ZN(new_n268));
  AND2_X1   g0068(.A1(new_n253), .A2(new_n225), .ZN(new_n269));
  OAI221_X1 g0069(.A(new_n252), .B1(new_n254), .B2(new_n256), .C1(new_n268), .C2(new_n269), .ZN(new_n270));
  XNOR2_X1  g0070(.A(new_n270), .B(KEYINPUT9), .ZN(new_n271));
  OAI21_X1  g0071(.A(new_n249), .B1(G41), .B2(G45), .ZN(new_n272));
  INV_X1    g0072(.A(new_n272), .ZN(new_n273));
  NAND2_X1  g0073(.A1(G33), .A2(G41), .ZN(new_n274));
  NAND3_X1  g0074(.A1(new_n274), .A2(G1), .A3(G13), .ZN(new_n275));
  NAND3_X1  g0075(.A1(new_n273), .A2(new_n275), .A3(G274), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n275), .A2(new_n272), .ZN(new_n277));
  OAI21_X1  g0077(.A(new_n276), .B1(new_n208), .B2(new_n277), .ZN(new_n278));
  XOR2_X1   g0078(.A(new_n278), .B(KEYINPUT65), .Z(new_n279));
  INV_X1    g0079(.A(KEYINPUT3), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n280), .A2(new_n266), .ZN(new_n281));
  NAND2_X1  g0081(.A1(KEYINPUT3), .A2(G33), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n281), .A2(new_n282), .ZN(new_n283));
  AND2_X1   g0083(.A1(KEYINPUT66), .A2(G1698), .ZN(new_n284));
  NOR2_X1   g0084(.A1(KEYINPUT66), .A2(G1698), .ZN(new_n285));
  NOR2_X1   g0085(.A1(new_n284), .A2(new_n285), .ZN(new_n286));
  NAND3_X1  g0086(.A1(new_n283), .A2(new_n286), .A3(G222), .ZN(new_n287));
  NAND3_X1  g0087(.A1(new_n283), .A2(G223), .A3(G1698), .ZN(new_n288));
  INV_X1    g0088(.A(G77), .ZN(new_n289));
  OAI211_X1 g0089(.A(new_n287), .B(new_n288), .C1(new_n289), .C2(new_n283), .ZN(new_n290));
  INV_X1    g0090(.A(new_n290), .ZN(new_n291));
  OAI21_X1  g0091(.A(new_n279), .B1(new_n275), .B2(new_n291), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n292), .A2(G200), .ZN(new_n293));
  INV_X1    g0093(.A(G190), .ZN(new_n294));
  OAI211_X1 g0094(.A(new_n271), .B(new_n293), .C1(new_n294), .C2(new_n292), .ZN(new_n295));
  XNOR2_X1  g0095(.A(new_n295), .B(KEYINPUT10), .ZN(new_n296));
  OR2_X1    g0096(.A1(new_n292), .A2(G179), .ZN(new_n297));
  INV_X1    g0097(.A(G169), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n292), .A2(new_n298), .ZN(new_n299));
  NAND3_X1  g0099(.A1(new_n297), .A2(new_n270), .A3(new_n299), .ZN(new_n300));
  XNOR2_X1  g0100(.A(KEYINPUT15), .B(G87), .ZN(new_n301));
  INV_X1    g0101(.A(new_n301), .ZN(new_n302));
  AOI22_X1  g0102(.A1(new_n302), .A2(new_n267), .B1(G20), .B2(G77), .ZN(new_n303));
  NOR2_X1   g0103(.A1(new_n259), .A2(KEYINPUT67), .ZN(new_n304));
  INV_X1    g0104(.A(KEYINPUT67), .ZN(new_n305));
  OAI21_X1  g0105(.A(new_n265), .B1(new_n305), .B2(new_n258), .ZN(new_n306));
  OAI21_X1  g0106(.A(new_n303), .B1(new_n304), .B2(new_n306), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n253), .A2(new_n225), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n307), .A2(new_n308), .ZN(new_n309));
  INV_X1    g0109(.A(new_n254), .ZN(new_n310));
  AOI21_X1  g0110(.A(new_n289), .B1(new_n249), .B2(G20), .ZN(new_n311));
  AOI22_X1  g0111(.A1(new_n310), .A2(new_n311), .B1(new_n289), .B2(new_n251), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n309), .A2(new_n312), .ZN(new_n313));
  INV_X1    g0113(.A(G238), .ZN(new_n314));
  INV_X1    g0114(.A(G1698), .ZN(new_n315));
  INV_X1    g0115(.A(KEYINPUT66), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n316), .A2(new_n315), .ZN(new_n317));
  NAND2_X1  g0117(.A1(KEYINPUT66), .A2(G1698), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n317), .A2(new_n318), .ZN(new_n319));
  OAI221_X1 g0119(.A(new_n283), .B1(new_n314), .B2(new_n315), .C1(new_n319), .C2(new_n214), .ZN(new_n320));
  AOI21_X1  g0120(.A(new_n225), .B1(G33), .B2(G41), .ZN(new_n321));
  OAI211_X1 g0121(.A(new_n320), .B(new_n321), .C1(G107), .C2(new_n283), .ZN(new_n322));
  INV_X1    g0122(.A(G244), .ZN(new_n323));
  NOR2_X1   g0123(.A1(new_n277), .A2(new_n323), .ZN(new_n324));
  INV_X1    g0124(.A(G274), .ZN(new_n325));
  NOR3_X1   g0125(.A1(new_n321), .A2(new_n325), .A3(new_n272), .ZN(new_n326));
  NOR2_X1   g0126(.A1(new_n324), .A2(new_n326), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n322), .A2(new_n327), .ZN(new_n328));
  INV_X1    g0128(.A(new_n328), .ZN(new_n329));
  AOI21_X1  g0129(.A(new_n313), .B1(new_n329), .B2(G190), .ZN(new_n330));
  INV_X1    g0130(.A(G200), .ZN(new_n331));
  OAI21_X1  g0131(.A(new_n330), .B1(new_n331), .B2(new_n329), .ZN(new_n332));
  INV_X1    g0132(.A(G179), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n329), .A2(new_n333), .ZN(new_n334));
  AOI22_X1  g0134(.A1(new_n328), .A2(new_n298), .B1(new_n309), .B2(new_n312), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n334), .A2(new_n335), .ZN(new_n336));
  AND4_X1   g0136(.A1(new_n296), .A2(new_n300), .A3(new_n332), .A4(new_n336), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n258), .A2(G159), .ZN(new_n338));
  AND2_X1   g0138(.A1(G58), .A2(G68), .ZN(new_n339));
  OAI21_X1  g0139(.A(G20), .B1(new_n339), .B2(new_n201), .ZN(new_n340));
  OAI21_X1  g0140(.A(new_n338), .B1(new_n340), .B2(KEYINPUT69), .ZN(new_n341));
  INV_X1    g0141(.A(KEYINPUT69), .ZN(new_n342));
  XNOR2_X1  g0142(.A(G58), .B(G68), .ZN(new_n343));
  AOI21_X1  g0143(.A(new_n342), .B1(new_n343), .B2(G20), .ZN(new_n344));
  NOR2_X1   g0144(.A1(new_n341), .A2(new_n344), .ZN(new_n345));
  INV_X1    g0145(.A(KEYINPUT7), .ZN(new_n346));
  NOR2_X1   g0146(.A1(KEYINPUT3), .A2(G33), .ZN(new_n347));
  XNOR2_X1  g0147(.A(KEYINPUT68), .B(G33), .ZN(new_n348));
  AOI21_X1  g0148(.A(new_n347), .B1(new_n348), .B2(KEYINPUT3), .ZN(new_n349));
  AOI21_X1  g0149(.A(new_n346), .B1(new_n349), .B2(new_n226), .ZN(new_n350));
  AND2_X1   g0150(.A1(KEYINPUT68), .A2(G33), .ZN(new_n351));
  NOR2_X1   g0151(.A1(KEYINPUT68), .A2(G33), .ZN(new_n352));
  OAI21_X1  g0152(.A(KEYINPUT3), .B1(new_n351), .B2(new_n352), .ZN(new_n353));
  NAND4_X1  g0153(.A1(new_n353), .A2(new_n346), .A3(new_n226), .A4(new_n281), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n354), .A2(G68), .ZN(new_n355));
  OAI211_X1 g0155(.A(KEYINPUT16), .B(new_n345), .C1(new_n350), .C2(new_n355), .ZN(new_n356));
  XNOR2_X1  g0156(.A(KEYINPUT70), .B(KEYINPUT16), .ZN(new_n357));
  INV_X1    g0157(.A(KEYINPUT68), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n358), .A2(new_n266), .ZN(new_n359));
  NAND2_X1  g0159(.A1(KEYINPUT68), .A2(G33), .ZN(new_n360));
  NAND3_X1  g0160(.A1(new_n359), .A2(new_n280), .A3(new_n360), .ZN(new_n361));
  AND3_X1   g0161(.A1(new_n282), .A2(KEYINPUT7), .A3(new_n226), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n361), .A2(new_n362), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n282), .A2(new_n226), .ZN(new_n364));
  OAI21_X1  g0164(.A(new_n346), .B1(new_n364), .B2(new_n347), .ZN(new_n365));
  AOI21_X1  g0165(.A(new_n243), .B1(new_n363), .B2(new_n365), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n340), .A2(KEYINPUT69), .ZN(new_n367));
  NAND3_X1  g0167(.A1(new_n343), .A2(new_n342), .A3(G20), .ZN(new_n368));
  NAND3_X1  g0168(.A1(new_n367), .A2(new_n368), .A3(new_n338), .ZN(new_n369));
  OAI21_X1  g0169(.A(new_n357), .B1(new_n366), .B2(new_n369), .ZN(new_n370));
  NAND3_X1  g0170(.A1(new_n356), .A2(new_n370), .A3(new_n308), .ZN(new_n371));
  INV_X1    g0171(.A(KEYINPUT72), .ZN(new_n372));
  INV_X1    g0172(.A(G13), .ZN(new_n373));
  NOR2_X1   g0173(.A1(new_n373), .A2(G1), .ZN(new_n374));
  NAND4_X1  g0174(.A1(new_n374), .A2(new_n262), .A3(new_n264), .A4(G20), .ZN(new_n375));
  NOR2_X1   g0175(.A1(new_n263), .A2(G58), .ZN(new_n376));
  NOR2_X1   g0176(.A1(new_n213), .A2(KEYINPUT8), .ZN(new_n377));
  OAI21_X1  g0177(.A(new_n255), .B1(new_n376), .B2(new_n377), .ZN(new_n378));
  OAI211_X1 g0178(.A(KEYINPUT71), .B(new_n375), .C1(new_n378), .C2(new_n254), .ZN(new_n379));
  INV_X1    g0179(.A(new_n379), .ZN(new_n380));
  NAND4_X1  g0180(.A1(new_n269), .A2(new_n265), .A3(new_n250), .A4(new_n255), .ZN(new_n381));
  AOI21_X1  g0181(.A(KEYINPUT71), .B1(new_n381), .B2(new_n375), .ZN(new_n382));
  OAI21_X1  g0182(.A(new_n372), .B1(new_n380), .B2(new_n382), .ZN(new_n383));
  OAI21_X1  g0183(.A(new_n375), .B1(new_n378), .B2(new_n254), .ZN(new_n384));
  INV_X1    g0184(.A(KEYINPUT71), .ZN(new_n385));
  NAND2_X1  g0185(.A1(new_n384), .A2(new_n385), .ZN(new_n386));
  NAND3_X1  g0186(.A1(new_n386), .A2(KEYINPUT72), .A3(new_n379), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n383), .A2(new_n387), .ZN(new_n388));
  NOR2_X1   g0188(.A1(new_n277), .A2(new_n214), .ZN(new_n389));
  NOR2_X1   g0189(.A1(new_n389), .A2(new_n326), .ZN(new_n390));
  NAND2_X1  g0190(.A1(new_n353), .A2(new_n281), .ZN(new_n391));
  NAND3_X1  g0191(.A1(new_n317), .A2(G223), .A3(new_n318), .ZN(new_n392));
  NAND2_X1  g0192(.A1(G226), .A2(G1698), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n392), .A2(new_n393), .ZN(new_n394));
  AOI22_X1  g0194(.A1(new_n391), .A2(new_n394), .B1(G33), .B2(G87), .ZN(new_n395));
  OAI21_X1  g0195(.A(new_n390), .B1(new_n395), .B2(new_n275), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n396), .A2(G169), .ZN(new_n397));
  OAI211_X1 g0197(.A(new_n390), .B(G179), .C1(new_n395), .C2(new_n275), .ZN(new_n398));
  AOI22_X1  g0198(.A1(new_n371), .A2(new_n388), .B1(new_n397), .B2(new_n398), .ZN(new_n399));
  INV_X1    g0199(.A(KEYINPUT18), .ZN(new_n400));
  XNOR2_X1  g0200(.A(new_n399), .B(new_n400), .ZN(new_n401));
  OAI211_X1 g0201(.A(new_n390), .B(new_n294), .C1(new_n395), .C2(new_n275), .ZN(new_n402));
  OAI21_X1  g0202(.A(new_n276), .B1(new_n277), .B2(new_n214), .ZN(new_n403));
  NAND2_X1  g0203(.A1(G33), .A2(G87), .ZN(new_n404));
  AOI22_X1  g0204(.A1(new_n286), .A2(G223), .B1(G226), .B2(G1698), .ZN(new_n405));
  OAI21_X1  g0205(.A(new_n404), .B1(new_n405), .B2(new_n349), .ZN(new_n406));
  AOI21_X1  g0206(.A(new_n403), .B1(new_n406), .B2(new_n321), .ZN(new_n407));
  OAI21_X1  g0207(.A(new_n402), .B1(new_n407), .B2(G200), .ZN(new_n408));
  NAND3_X1  g0208(.A1(new_n408), .A2(new_n371), .A3(new_n388), .ZN(new_n409));
  INV_X1    g0209(.A(KEYINPUT17), .ZN(new_n410));
  XNOR2_X1  g0210(.A(new_n409), .B(new_n410), .ZN(new_n411));
  NOR2_X1   g0211(.A1(new_n401), .A2(new_n411), .ZN(new_n412));
  OAI22_X1  g0212(.A1(new_n319), .A2(new_n208), .B1(new_n214), .B2(new_n315), .ZN(new_n413));
  AOI22_X1  g0213(.A1(new_n413), .A2(new_n283), .B1(G33), .B2(G97), .ZN(new_n414));
  NOR2_X1   g0214(.A1(new_n414), .A2(new_n275), .ZN(new_n415));
  OAI21_X1  g0215(.A(new_n276), .B1(new_n277), .B2(new_n314), .ZN(new_n416));
  OR3_X1    g0216(.A1(new_n415), .A2(KEYINPUT13), .A3(new_n416), .ZN(new_n417));
  OAI21_X1  g0217(.A(KEYINPUT13), .B1(new_n415), .B2(new_n416), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n417), .A2(new_n418), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n419), .A2(G200), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n251), .A2(new_n243), .ZN(new_n421));
  XNOR2_X1  g0221(.A(new_n421), .B(KEYINPUT12), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n267), .A2(G77), .ZN(new_n423));
  OAI221_X1 g0223(.A(new_n423), .B1(new_n226), .B2(G68), .C1(new_n207), .C2(new_n259), .ZN(new_n424));
  NAND3_X1  g0224(.A1(new_n424), .A2(KEYINPUT11), .A3(new_n308), .ZN(new_n425));
  NAND3_X1  g0225(.A1(new_n310), .A2(G68), .A3(new_n255), .ZN(new_n426));
  NAND3_X1  g0226(.A1(new_n422), .A2(new_n425), .A3(new_n426), .ZN(new_n427));
  AOI21_X1  g0227(.A(KEYINPUT11), .B1(new_n424), .B2(new_n308), .ZN(new_n428));
  NOR2_X1   g0228(.A1(new_n427), .A2(new_n428), .ZN(new_n429));
  NAND3_X1  g0229(.A1(new_n417), .A2(G190), .A3(new_n418), .ZN(new_n430));
  NAND3_X1  g0230(.A1(new_n420), .A2(new_n429), .A3(new_n430), .ZN(new_n431));
  INV_X1    g0231(.A(new_n431), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n419), .A2(G169), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n433), .A2(KEYINPUT14), .ZN(new_n434));
  NAND3_X1  g0234(.A1(new_n417), .A2(G179), .A3(new_n418), .ZN(new_n435));
  INV_X1    g0235(.A(KEYINPUT14), .ZN(new_n436));
  NAND3_X1  g0236(.A1(new_n419), .A2(new_n436), .A3(G169), .ZN(new_n437));
  NAND3_X1  g0237(.A1(new_n434), .A2(new_n435), .A3(new_n437), .ZN(new_n438));
  INV_X1    g0238(.A(new_n429), .ZN(new_n439));
  AOI21_X1  g0239(.A(new_n432), .B1(new_n438), .B2(new_n439), .ZN(new_n440));
  NAND3_X1  g0240(.A1(new_n337), .A2(new_n412), .A3(new_n440), .ZN(new_n441));
  NAND2_X1  g0241(.A1(G33), .A2(G283), .ZN(new_n442));
  OAI211_X1 g0242(.A(new_n442), .B(new_n226), .C1(G33), .C2(new_n215), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n209), .A2(G20), .ZN(new_n444));
  NAND3_X1  g0244(.A1(new_n443), .A2(new_n308), .A3(new_n444), .ZN(new_n445));
  INV_X1    g0245(.A(KEYINPUT20), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n445), .A2(new_n446), .ZN(new_n447));
  NAND4_X1  g0247(.A1(new_n443), .A2(KEYINPUT20), .A3(new_n308), .A4(new_n444), .ZN(new_n448));
  NAND3_X1  g0248(.A1(new_n447), .A2(KEYINPUT77), .A3(new_n448), .ZN(new_n449));
  NAND2_X1  g0249(.A1(new_n249), .A2(G33), .ZN(new_n450));
  NAND3_X1  g0250(.A1(new_n269), .A2(new_n250), .A3(new_n450), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n451), .A2(G116), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n250), .A2(new_n209), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n452), .A2(new_n453), .ZN(new_n454));
  INV_X1    g0254(.A(KEYINPUT77), .ZN(new_n455));
  NAND3_X1  g0255(.A1(new_n445), .A2(new_n455), .A3(new_n446), .ZN(new_n456));
  NAND3_X1  g0256(.A1(new_n449), .A2(new_n454), .A3(new_n456), .ZN(new_n457));
  NAND3_X1  g0257(.A1(new_n391), .A2(G264), .A3(G1698), .ZN(new_n458));
  NAND3_X1  g0258(.A1(new_n391), .A2(G257), .A3(new_n286), .ZN(new_n459));
  INV_X1    g0259(.A(new_n283), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n460), .A2(G303), .ZN(new_n461));
  NAND3_X1  g0261(.A1(new_n458), .A2(new_n459), .A3(new_n461), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n462), .A2(new_n321), .ZN(new_n463));
  XNOR2_X1  g0263(.A(KEYINPUT5), .B(G41), .ZN(new_n464));
  INV_X1    g0264(.A(G45), .ZN(new_n465));
  NOR2_X1   g0265(.A1(new_n465), .A2(G1), .ZN(new_n466));
  NAND4_X1  g0266(.A1(new_n464), .A2(new_n275), .A3(G274), .A4(new_n466), .ZN(new_n467));
  INV_X1    g0267(.A(new_n467), .ZN(new_n468));
  AOI21_X1  g0268(.A(new_n321), .B1(new_n466), .B2(new_n464), .ZN(new_n469));
  AOI21_X1  g0269(.A(new_n468), .B1(G270), .B2(new_n469), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n463), .A2(new_n470), .ZN(new_n471));
  AOI21_X1  g0271(.A(new_n457), .B1(new_n471), .B2(G200), .ZN(new_n472));
  AOI21_X1  g0272(.A(new_n319), .B1(new_n353), .B2(new_n281), .ZN(new_n473));
  AOI22_X1  g0273(.A1(new_n473), .A2(G257), .B1(G303), .B2(new_n460), .ZN(new_n474));
  AOI21_X1  g0274(.A(new_n275), .B1(new_n474), .B2(new_n458), .ZN(new_n475));
  INV_X1    g0275(.A(new_n470), .ZN(new_n476));
  NOR2_X1   g0276(.A1(new_n475), .A2(new_n476), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n477), .A2(G190), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n472), .A2(new_n478), .ZN(new_n479));
  OAI211_X1 g0279(.A(G169), .B(new_n457), .C1(new_n475), .C2(new_n476), .ZN(new_n480));
  INV_X1    g0280(.A(KEYINPUT21), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n480), .A2(new_n481), .ZN(new_n482));
  NAND3_X1  g0282(.A1(new_n477), .A2(G179), .A3(new_n457), .ZN(new_n483));
  NAND4_X1  g0283(.A1(new_n471), .A2(KEYINPUT21), .A3(G169), .A4(new_n457), .ZN(new_n484));
  NAND4_X1  g0284(.A1(new_n479), .A2(new_n482), .A3(new_n483), .A4(new_n484), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n469), .A2(G264), .ZN(new_n486));
  NAND3_X1  g0286(.A1(new_n317), .A2(G250), .A3(new_n318), .ZN(new_n487));
  NAND2_X1  g0287(.A1(G257), .A2(G1698), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n487), .A2(new_n488), .ZN(new_n489));
  AOI22_X1  g0289(.A1(new_n391), .A2(new_n489), .B1(G294), .B2(new_n348), .ZN(new_n490));
  OAI211_X1 g0290(.A(new_n467), .B(new_n486), .C1(new_n490), .C2(new_n275), .ZN(new_n491));
  NAND3_X1  g0291(.A1(new_n491), .A2(KEYINPUT78), .A3(G169), .ZN(new_n492));
  AND2_X1   g0292(.A1(new_n391), .A2(new_n489), .ZN(new_n493));
  INV_X1    g0293(.A(G294), .ZN(new_n494));
  AOI21_X1  g0294(.A(new_n494), .B1(new_n359), .B2(new_n360), .ZN(new_n495));
  OAI21_X1  g0295(.A(new_n321), .B1(new_n493), .B2(new_n495), .ZN(new_n496));
  NAND4_X1  g0296(.A1(new_n496), .A2(G179), .A3(new_n467), .A4(new_n486), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n492), .A2(new_n497), .ZN(new_n498));
  AOI21_X1  g0298(.A(KEYINPUT78), .B1(new_n491), .B2(G169), .ZN(new_n499));
  NAND2_X1  g0299(.A1(KEYINPUT22), .A2(G87), .ZN(new_n500));
  NOR3_X1   g0300(.A1(new_n349), .A2(G20), .A3(new_n500), .ZN(new_n501));
  OAI211_X1 g0301(.A(new_n226), .B(G116), .C1(new_n351), .C2(new_n352), .ZN(new_n502));
  INV_X1    g0302(.A(KEYINPUT23), .ZN(new_n503));
  OAI21_X1  g0303(.A(new_n503), .B1(new_n226), .B2(G107), .ZN(new_n504));
  INV_X1    g0304(.A(G107), .ZN(new_n505));
  NAND3_X1  g0305(.A1(new_n505), .A2(KEYINPUT23), .A3(G20), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n504), .A2(new_n506), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n226), .A2(G87), .ZN(new_n508));
  AOI21_X1  g0308(.A(new_n508), .B1(new_n281), .B2(new_n282), .ZN(new_n509));
  OAI211_X1 g0309(.A(new_n502), .B(new_n507), .C1(new_n509), .C2(KEYINPUT22), .ZN(new_n510));
  OAI21_X1  g0310(.A(KEYINPUT24), .B1(new_n501), .B2(new_n510), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n502), .A2(new_n507), .ZN(new_n512));
  INV_X1    g0312(.A(new_n508), .ZN(new_n513));
  AOI21_X1  g0313(.A(KEYINPUT22), .B1(new_n283), .B2(new_n513), .ZN(new_n514));
  NOR2_X1   g0314(.A1(new_n512), .A2(new_n514), .ZN(new_n515));
  NAND4_X1  g0315(.A1(new_n391), .A2(KEYINPUT22), .A3(new_n226), .A4(G87), .ZN(new_n516));
  INV_X1    g0316(.A(KEYINPUT24), .ZN(new_n517));
  NAND3_X1  g0317(.A1(new_n515), .A2(new_n516), .A3(new_n517), .ZN(new_n518));
  AOI21_X1  g0318(.A(new_n269), .B1(new_n511), .B2(new_n518), .ZN(new_n519));
  INV_X1    g0319(.A(new_n451), .ZN(new_n520));
  INV_X1    g0320(.A(KEYINPUT25), .ZN(new_n521));
  OAI21_X1  g0321(.A(new_n521), .B1(new_n250), .B2(G107), .ZN(new_n522));
  NOR3_X1   g0322(.A1(new_n250), .A2(new_n521), .A3(G107), .ZN(new_n523));
  INV_X1    g0323(.A(new_n523), .ZN(new_n524));
  AOI22_X1  g0324(.A1(new_n520), .A2(G107), .B1(new_n522), .B2(new_n524), .ZN(new_n525));
  INV_X1    g0325(.A(new_n525), .ZN(new_n526));
  OAI22_X1  g0326(.A1(new_n498), .A2(new_n499), .B1(new_n519), .B2(new_n526), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n511), .A2(new_n518), .ZN(new_n528));
  AOI21_X1  g0328(.A(new_n526), .B1(new_n528), .B2(new_n308), .ZN(new_n529));
  OR2_X1    g0329(.A1(new_n491), .A2(new_n294), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n491), .A2(G200), .ZN(new_n531));
  NAND3_X1  g0331(.A1(new_n529), .A2(new_n530), .A3(new_n531), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n527), .A2(new_n532), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n520), .A2(new_n302), .ZN(new_n534));
  INV_X1    g0334(.A(KEYINPUT76), .ZN(new_n535));
  AOI211_X1 g0335(.A(G20), .B(new_n243), .C1(new_n353), .C2(new_n281), .ZN(new_n536));
  NOR3_X1   g0336(.A1(G87), .A2(G97), .A3(G107), .ZN(new_n537));
  AOI21_X1  g0337(.A(G20), .B1(G33), .B2(G97), .ZN(new_n538));
  OAI21_X1  g0338(.A(KEYINPUT19), .B1(new_n537), .B2(new_n538), .ZN(new_n539));
  INV_X1    g0339(.A(KEYINPUT19), .ZN(new_n540));
  NAND3_X1  g0340(.A1(new_n267), .A2(new_n540), .A3(G97), .ZN(new_n541));
  AND2_X1   g0341(.A1(new_n539), .A2(new_n541), .ZN(new_n542));
  OAI21_X1  g0342(.A(new_n308), .B1(new_n536), .B2(new_n542), .ZN(new_n543));
  NOR2_X1   g0343(.A1(new_n302), .A2(new_n250), .ZN(new_n544));
  INV_X1    g0344(.A(new_n544), .ZN(new_n545));
  AOI21_X1  g0345(.A(new_n535), .B1(new_n543), .B2(new_n545), .ZN(new_n546));
  AOI21_X1  g0346(.A(new_n280), .B1(new_n359), .B2(new_n360), .ZN(new_n547));
  OAI211_X1 g0347(.A(new_n226), .B(G68), .C1(new_n547), .C2(new_n347), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n539), .A2(new_n541), .ZN(new_n549));
  AOI21_X1  g0349(.A(new_n269), .B1(new_n548), .B2(new_n549), .ZN(new_n550));
  NOR3_X1   g0350(.A1(new_n550), .A2(KEYINPUT76), .A3(new_n544), .ZN(new_n551));
  OAI21_X1  g0351(.A(new_n534), .B1(new_n546), .B2(new_n551), .ZN(new_n552));
  AOI22_X1  g0352(.A1(new_n473), .A2(G238), .B1(G116), .B2(new_n348), .ZN(new_n553));
  OAI211_X1 g0353(.A(G244), .B(G1698), .C1(new_n547), .C2(new_n347), .ZN(new_n554));
  INV_X1    g0354(.A(KEYINPUT75), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  NAND4_X1  g0356(.A1(new_n391), .A2(KEYINPUT75), .A3(G244), .A4(G1698), .ZN(new_n557));
  NAND3_X1  g0357(.A1(new_n553), .A2(new_n556), .A3(new_n557), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n558), .A2(new_n321), .ZN(new_n559));
  OAI21_X1  g0359(.A(KEYINPUT74), .B1(new_n465), .B2(G1), .ZN(new_n560));
  INV_X1    g0360(.A(KEYINPUT74), .ZN(new_n561));
  NAND3_X1  g0361(.A1(new_n561), .A2(new_n249), .A3(G45), .ZN(new_n562));
  NAND4_X1  g0362(.A1(new_n275), .A2(new_n560), .A3(new_n562), .A4(G250), .ZN(new_n563));
  NAND3_X1  g0363(.A1(new_n275), .A2(G274), .A3(new_n466), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n563), .A2(new_n564), .ZN(new_n565));
  INV_X1    g0365(.A(new_n565), .ZN(new_n566));
  NAND3_X1  g0366(.A1(new_n559), .A2(new_n333), .A3(new_n566), .ZN(new_n567));
  AOI21_X1  g0367(.A(new_n565), .B1(new_n558), .B2(new_n321), .ZN(new_n568));
  OAI211_X1 g0368(.A(new_n552), .B(new_n567), .C1(G169), .C2(new_n568), .ZN(new_n569));
  NAND3_X1  g0369(.A1(new_n559), .A2(G190), .A3(new_n566), .ZN(new_n570));
  INV_X1    g0370(.A(G87), .ZN(new_n571));
  NOR2_X1   g0371(.A1(new_n451), .A2(new_n571), .ZN(new_n572));
  OAI21_X1  g0372(.A(KEYINPUT76), .B1(new_n550), .B2(new_n544), .ZN(new_n573));
  AOI21_X1  g0373(.A(G20), .B1(new_n353), .B2(new_n281), .ZN(new_n574));
  AOI22_X1  g0374(.A1(new_n574), .A2(G68), .B1(new_n539), .B2(new_n541), .ZN(new_n575));
  OAI211_X1 g0375(.A(new_n535), .B(new_n545), .C1(new_n575), .C2(new_n269), .ZN(new_n576));
  AOI21_X1  g0376(.A(new_n572), .B1(new_n573), .B2(new_n576), .ZN(new_n577));
  OAI211_X1 g0377(.A(new_n570), .B(new_n577), .C1(new_n331), .C2(new_n568), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n258), .A2(G77), .ZN(new_n579));
  AND3_X1   g0379(.A1(new_n505), .A2(KEYINPUT6), .A3(G97), .ZN(new_n580));
  XNOR2_X1  g0380(.A(G97), .B(G107), .ZN(new_n581));
  INV_X1    g0381(.A(KEYINPUT6), .ZN(new_n582));
  AOI21_X1  g0382(.A(new_n580), .B1(new_n581), .B2(new_n582), .ZN(new_n583));
  OAI21_X1  g0383(.A(new_n579), .B1(new_n583), .B2(new_n226), .ZN(new_n584));
  AOI21_X1  g0384(.A(new_n505), .B1(new_n363), .B2(new_n365), .ZN(new_n585));
  OAI21_X1  g0385(.A(new_n308), .B1(new_n584), .B2(new_n585), .ZN(new_n586));
  NOR2_X1   g0386(.A1(new_n250), .A2(G97), .ZN(new_n587));
  AOI21_X1  g0387(.A(new_n587), .B1(new_n520), .B2(G97), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n586), .A2(new_n588), .ZN(new_n589));
  NOR3_X1   g0389(.A1(new_n284), .A2(new_n285), .A3(new_n323), .ZN(new_n590));
  INV_X1    g0390(.A(KEYINPUT4), .ZN(new_n591));
  AOI21_X1  g0391(.A(new_n591), .B1(new_n281), .B2(new_n282), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n590), .A2(new_n592), .ZN(new_n593));
  NAND3_X1  g0393(.A1(new_n283), .A2(G250), .A3(G1698), .ZN(new_n594));
  NAND3_X1  g0394(.A1(new_n593), .A2(new_n442), .A3(new_n594), .ZN(new_n595));
  AOI21_X1  g0395(.A(KEYINPUT4), .B1(new_n391), .B2(new_n590), .ZN(new_n596));
  OAI21_X1  g0396(.A(new_n321), .B1(new_n595), .B2(new_n596), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n464), .A2(new_n466), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n598), .A2(new_n275), .ZN(new_n599));
  OAI21_X1  g0399(.A(new_n467), .B1(new_n599), .B2(new_n216), .ZN(new_n600));
  INV_X1    g0400(.A(new_n600), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n597), .A2(new_n601), .ZN(new_n602));
  AOI21_X1  g0402(.A(new_n589), .B1(G200), .B2(new_n602), .ZN(new_n603));
  OAI21_X1  g0403(.A(new_n603), .B1(new_n294), .B2(new_n602), .ZN(new_n604));
  AOI22_X1  g0404(.A1(new_n602), .A2(new_n298), .B1(new_n586), .B2(new_n588), .ZN(new_n605));
  INV_X1    g0405(.A(new_n442), .ZN(new_n606));
  AOI21_X1  g0406(.A(new_n606), .B1(new_n590), .B2(new_n592), .ZN(new_n607));
  NAND3_X1  g0407(.A1(new_n317), .A2(G244), .A3(new_n318), .ZN(new_n608));
  AOI21_X1  g0408(.A(new_n608), .B1(new_n281), .B2(new_n353), .ZN(new_n609));
  OAI211_X1 g0409(.A(new_n607), .B(new_n594), .C1(new_n609), .C2(KEYINPUT4), .ZN(new_n610));
  AOI21_X1  g0410(.A(new_n600), .B1(new_n610), .B2(new_n321), .ZN(new_n611));
  AOI21_X1  g0411(.A(KEYINPUT73), .B1(new_n611), .B2(new_n333), .ZN(new_n612));
  AND4_X1   g0412(.A1(KEYINPUT73), .A2(new_n597), .A3(new_n333), .A4(new_n601), .ZN(new_n613));
  OAI21_X1  g0413(.A(new_n605), .B1(new_n612), .B2(new_n613), .ZN(new_n614));
  NAND4_X1  g0414(.A1(new_n569), .A2(new_n578), .A3(new_n604), .A4(new_n614), .ZN(new_n615));
  NOR4_X1   g0415(.A1(new_n441), .A2(new_n485), .A3(new_n533), .A4(new_n615), .ZN(G372));
  INV_X1    g0416(.A(new_n441), .ZN(new_n617));
  AND2_X1   g0417(.A1(new_n492), .A2(new_n497), .ZN(new_n618));
  INV_X1    g0418(.A(new_n499), .ZN(new_n619));
  AOI21_X1  g0419(.A(new_n529), .B1(new_n618), .B2(new_n619), .ZN(new_n620));
  NAND3_X1  g0420(.A1(new_n482), .A2(new_n484), .A3(new_n483), .ZN(new_n621));
  NOR2_X1   g0421(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  INV_X1    g0422(.A(KEYINPUT79), .ZN(new_n623));
  XNOR2_X1  g0423(.A(new_n565), .B(new_n623), .ZN(new_n624));
  AOI21_X1  g0424(.A(new_n624), .B1(new_n558), .B2(new_n321), .ZN(new_n625));
  OAI211_X1 g0425(.A(new_n552), .B(new_n567), .C1(G169), .C2(new_n625), .ZN(new_n626));
  OAI211_X1 g0426(.A(new_n570), .B(new_n577), .C1(new_n331), .C2(new_n625), .ZN(new_n627));
  NAND3_X1  g0427(.A1(new_n626), .A2(new_n532), .A3(new_n627), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n604), .A2(new_n614), .ZN(new_n629));
  NOR3_X1   g0429(.A1(new_n622), .A2(new_n628), .A3(new_n629), .ZN(new_n630));
  OAI21_X1  g0430(.A(new_n589), .B1(new_n611), .B2(G169), .ZN(new_n631));
  INV_X1    g0431(.A(KEYINPUT73), .ZN(new_n632));
  OAI21_X1  g0432(.A(new_n632), .B1(new_n602), .B2(G179), .ZN(new_n633));
  NAND3_X1  g0433(.A1(new_n611), .A2(KEYINPUT73), .A3(new_n333), .ZN(new_n634));
  AOI21_X1  g0434(.A(new_n631), .B1(new_n633), .B2(new_n634), .ZN(new_n635));
  NAND3_X1  g0435(.A1(new_n569), .A2(new_n578), .A3(new_n635), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n636), .A2(KEYINPUT26), .ZN(new_n637));
  INV_X1    g0437(.A(KEYINPUT26), .ZN(new_n638));
  NAND4_X1  g0438(.A1(new_n626), .A2(new_n627), .A3(new_n635), .A4(new_n638), .ZN(new_n639));
  NAND3_X1  g0439(.A1(new_n637), .A2(new_n626), .A3(new_n639), .ZN(new_n640));
  OAI21_X1  g0440(.A(new_n617), .B1(new_n630), .B2(new_n640), .ZN(new_n641));
  XNOR2_X1  g0441(.A(new_n641), .B(KEYINPUT80), .ZN(new_n642));
  INV_X1    g0442(.A(new_n300), .ZN(new_n643));
  XNOR2_X1  g0443(.A(new_n399), .B(KEYINPUT18), .ZN(new_n644));
  INV_X1    g0444(.A(new_n336), .ZN(new_n645));
  AOI22_X1  g0445(.A1(new_n438), .A2(new_n439), .B1(new_n431), .B2(new_n645), .ZN(new_n646));
  AND2_X1   g0446(.A1(new_n646), .A2(KEYINPUT81), .ZN(new_n647));
  XNOR2_X1  g0447(.A(new_n409), .B(KEYINPUT17), .ZN(new_n648));
  OAI21_X1  g0448(.A(new_n648), .B1(new_n646), .B2(KEYINPUT81), .ZN(new_n649));
  OAI21_X1  g0449(.A(new_n644), .B1(new_n647), .B2(new_n649), .ZN(new_n650));
  AOI21_X1  g0450(.A(new_n643), .B1(new_n650), .B2(new_n296), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n642), .A2(new_n651), .ZN(G369));
  NAND2_X1  g0452(.A1(new_n374), .A2(new_n226), .ZN(new_n653));
  OR2_X1    g0453(.A1(new_n653), .A2(KEYINPUT27), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n653), .A2(KEYINPUT27), .ZN(new_n655));
  NAND3_X1  g0455(.A1(new_n654), .A2(new_n655), .A3(G213), .ZN(new_n656));
  INV_X1    g0456(.A(G343), .ZN(new_n657));
  NOR2_X1   g0457(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  AND2_X1   g0458(.A1(new_n457), .A2(new_n658), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n621), .A2(new_n659), .ZN(new_n660));
  OAI21_X1  g0460(.A(new_n660), .B1(new_n485), .B2(new_n659), .ZN(new_n661));
  XNOR2_X1  g0461(.A(new_n661), .B(KEYINPUT82), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n662), .A2(G330), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n620), .A2(new_n658), .ZN(new_n664));
  INV_X1    g0464(.A(KEYINPUT83), .ZN(new_n665));
  XNOR2_X1  g0465(.A(new_n664), .B(new_n665), .ZN(new_n666));
  INV_X1    g0466(.A(new_n533), .ZN(new_n667));
  INV_X1    g0467(.A(new_n658), .ZN(new_n668));
  OAI21_X1  g0468(.A(new_n667), .B1(new_n529), .B2(new_n668), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n666), .A2(new_n669), .ZN(new_n670));
  INV_X1    g0470(.A(new_n670), .ZN(new_n671));
  NOR2_X1   g0471(.A1(new_n663), .A2(new_n671), .ZN(new_n672));
  INV_X1    g0472(.A(new_n672), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n621), .A2(new_n668), .ZN(new_n674));
  INV_X1    g0474(.A(new_n674), .ZN(new_n675));
  AOI22_X1  g0475(.A1(new_n670), .A2(new_n675), .B1(new_n620), .B2(new_n668), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n673), .A2(new_n676), .ZN(G399));
  INV_X1    g0477(.A(new_n222), .ZN(new_n678));
  NOR2_X1   g0478(.A1(new_n678), .A2(G41), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n537), .A2(new_n209), .ZN(new_n680));
  NOR3_X1   g0480(.A1(new_n679), .A2(new_n249), .A3(new_n680), .ZN(new_n681));
  AOI21_X1  g0481(.A(new_n681), .B1(new_n229), .B2(new_n679), .ZN(new_n682));
  XOR2_X1   g0482(.A(new_n682), .B(KEYINPUT28), .Z(new_n683));
  OAI21_X1  g0483(.A(new_n668), .B1(new_n640), .B2(new_n630), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n684), .A2(KEYINPUT86), .ZN(new_n685));
  INV_X1    g0485(.A(KEYINPUT29), .ZN(new_n686));
  INV_X1    g0486(.A(KEYINPUT86), .ZN(new_n687));
  OAI211_X1 g0487(.A(new_n687), .B(new_n668), .C1(new_n640), .C2(new_n630), .ZN(new_n688));
  NAND3_X1  g0488(.A1(new_n685), .A2(new_n686), .A3(new_n688), .ZN(new_n689));
  INV_X1    g0489(.A(KEYINPUT87), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  NAND3_X1  g0491(.A1(new_n626), .A2(new_n635), .A3(new_n627), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n692), .A2(KEYINPUT26), .ZN(new_n693));
  NAND4_X1  g0493(.A1(new_n569), .A2(new_n578), .A3(new_n635), .A4(new_n638), .ZN(new_n694));
  AND3_X1   g0494(.A1(new_n693), .A2(new_n626), .A3(new_n694), .ZN(new_n695));
  AND3_X1   g0495(.A1(new_n626), .A2(new_n532), .A3(new_n627), .ZN(new_n696));
  NAND4_X1  g0496(.A1(new_n527), .A2(new_n482), .A3(new_n483), .A4(new_n484), .ZN(new_n697));
  INV_X1    g0497(.A(KEYINPUT88), .ZN(new_n698));
  NOR2_X1   g0498(.A1(new_n602), .A2(new_n294), .ZN(new_n699));
  NOR2_X1   g0499(.A1(new_n611), .A2(new_n331), .ZN(new_n700));
  NOR3_X1   g0500(.A1(new_n699), .A2(new_n700), .A3(new_n589), .ZN(new_n701));
  OAI21_X1  g0501(.A(new_n698), .B1(new_n635), .B2(new_n701), .ZN(new_n702));
  NAND3_X1  g0502(.A1(new_n604), .A2(new_n614), .A3(KEYINPUT88), .ZN(new_n703));
  NAND4_X1  g0503(.A1(new_n696), .A2(new_n697), .A3(new_n702), .A4(new_n703), .ZN(new_n704));
  AOI21_X1  g0504(.A(new_n658), .B1(new_n695), .B2(new_n704), .ZN(new_n705));
  NAND2_X1  g0505(.A1(new_n705), .A2(KEYINPUT29), .ZN(new_n706));
  NAND4_X1  g0506(.A1(new_n685), .A2(KEYINPUT87), .A3(new_n686), .A4(new_n688), .ZN(new_n707));
  NAND3_X1  g0507(.A1(new_n691), .A2(new_n706), .A3(new_n707), .ZN(new_n708));
  AND4_X1   g0508(.A1(new_n569), .A2(new_n578), .A3(new_n604), .A4(new_n614), .ZN(new_n709));
  INV_X1    g0509(.A(new_n485), .ZN(new_n710));
  NAND4_X1  g0510(.A1(new_n709), .A2(new_n710), .A3(new_n667), .A4(new_n668), .ZN(new_n711));
  NAND4_X1  g0511(.A1(new_n568), .A2(new_n496), .A3(new_n486), .A4(new_n611), .ZN(new_n712));
  INV_X1    g0512(.A(KEYINPUT30), .ZN(new_n713));
  NAND2_X1  g0513(.A1(new_n477), .A2(G179), .ZN(new_n714));
  OR3_X1    g0514(.A1(new_n712), .A2(new_n713), .A3(new_n714), .ZN(new_n715));
  NOR2_X1   g0515(.A1(new_n477), .A2(G179), .ZN(new_n716));
  INV_X1    g0516(.A(new_n625), .ZN(new_n717));
  INV_X1    g0517(.A(new_n491), .ZN(new_n718));
  OAI21_X1  g0518(.A(KEYINPUT84), .B1(new_n718), .B2(new_n611), .ZN(new_n719));
  INV_X1    g0519(.A(KEYINPUT84), .ZN(new_n720));
  NAND3_X1  g0520(.A1(new_n602), .A2(new_n720), .A3(new_n491), .ZN(new_n721));
  NAND4_X1  g0521(.A1(new_n716), .A2(new_n717), .A3(new_n719), .A4(new_n721), .ZN(new_n722));
  INV_X1    g0522(.A(KEYINPUT85), .ZN(new_n723));
  NAND2_X1  g0523(.A1(new_n722), .A2(new_n723), .ZN(new_n724));
  OAI21_X1  g0524(.A(new_n713), .B1(new_n712), .B2(new_n714), .ZN(new_n725));
  NOR3_X1   g0525(.A1(new_n625), .A2(new_n477), .A3(G179), .ZN(new_n726));
  NAND4_X1  g0526(.A1(new_n726), .A2(KEYINPUT85), .A3(new_n719), .A4(new_n721), .ZN(new_n727));
  NAND4_X1  g0527(.A1(new_n715), .A2(new_n724), .A3(new_n725), .A4(new_n727), .ZN(new_n728));
  AOI22_X1  g0528(.A1(new_n711), .A2(KEYINPUT31), .B1(new_n658), .B2(new_n728), .ZN(new_n729));
  NAND3_X1  g0529(.A1(new_n715), .A2(new_n725), .A3(new_n722), .ZN(new_n730));
  AND3_X1   g0530(.A1(new_n730), .A2(KEYINPUT31), .A3(new_n658), .ZN(new_n731));
  OAI21_X1  g0531(.A(G330), .B1(new_n729), .B2(new_n731), .ZN(new_n732));
  NAND2_X1  g0532(.A1(new_n708), .A2(new_n732), .ZN(new_n733));
  INV_X1    g0533(.A(new_n733), .ZN(new_n734));
  OAI21_X1  g0534(.A(new_n683), .B1(new_n734), .B2(G1), .ZN(G364));
  AND2_X1   g0535(.A1(new_n662), .A2(G330), .ZN(new_n736));
  NOR2_X1   g0536(.A1(new_n662), .A2(G330), .ZN(new_n737));
  NOR2_X1   g0537(.A1(new_n373), .A2(G20), .ZN(new_n738));
  NAND2_X1  g0538(.A1(new_n738), .A2(G45), .ZN(new_n739));
  OR2_X1    g0539(.A1(new_n739), .A2(KEYINPUT89), .ZN(new_n740));
  NAND2_X1  g0540(.A1(new_n739), .A2(KEYINPUT89), .ZN(new_n741));
  NAND3_X1  g0541(.A1(new_n740), .A2(G1), .A3(new_n741), .ZN(new_n742));
  NOR2_X1   g0542(.A1(new_n679), .A2(new_n742), .ZN(new_n743));
  NOR3_X1   g0543(.A1(new_n736), .A2(new_n737), .A3(new_n743), .ZN(new_n744));
  XOR2_X1   g0544(.A(new_n744), .B(KEYINPUT90), .Z(new_n745));
  AOI21_X1  g0545(.A(new_n225), .B1(G20), .B2(new_n298), .ZN(new_n746));
  NOR2_X1   g0546(.A1(new_n226), .A2(new_n333), .ZN(new_n747));
  NOR2_X1   g0547(.A1(G190), .A2(G200), .ZN(new_n748));
  NAND2_X1  g0548(.A1(new_n747), .A2(new_n748), .ZN(new_n749));
  INV_X1    g0549(.A(new_n749), .ZN(new_n750));
  NAND3_X1  g0550(.A1(new_n333), .A2(new_n331), .A3(G190), .ZN(new_n751));
  NAND2_X1  g0551(.A1(new_n751), .A2(G20), .ZN(new_n752));
  AOI22_X1  g0552(.A1(new_n750), .A2(G311), .B1(G294), .B2(new_n752), .ZN(new_n753));
  INV_X1    g0553(.A(G326), .ZN(new_n754));
  NAND2_X1  g0554(.A1(new_n747), .A2(G200), .ZN(new_n755));
  NOR2_X1   g0555(.A1(new_n755), .A2(new_n294), .ZN(new_n756));
  INV_X1    g0556(.A(new_n756), .ZN(new_n757));
  OAI21_X1  g0557(.A(new_n753), .B1(new_n754), .B2(new_n757), .ZN(new_n758));
  XNOR2_X1  g0558(.A(new_n758), .B(KEYINPUT92), .ZN(new_n759));
  NOR2_X1   g0559(.A1(new_n226), .A2(G179), .ZN(new_n760));
  NAND2_X1  g0560(.A1(new_n760), .A2(new_n748), .ZN(new_n761));
  INV_X1    g0561(.A(G329), .ZN(new_n762));
  NAND3_X1  g0562(.A1(new_n747), .A2(G190), .A3(new_n331), .ZN(new_n763));
  INV_X1    g0563(.A(G322), .ZN(new_n764));
  OAI221_X1 g0564(.A(new_n460), .B1(new_n761), .B2(new_n762), .C1(new_n763), .C2(new_n764), .ZN(new_n765));
  NOR2_X1   g0565(.A1(new_n755), .A2(G190), .ZN(new_n766));
  INV_X1    g0566(.A(G317), .ZN(new_n767));
  NAND2_X1  g0567(.A1(new_n767), .A2(KEYINPUT33), .ZN(new_n768));
  OR2_X1    g0568(.A1(new_n767), .A2(KEYINPUT33), .ZN(new_n769));
  NAND3_X1  g0569(.A1(new_n766), .A2(new_n768), .A3(new_n769), .ZN(new_n770));
  INV_X1    g0570(.A(G283), .ZN(new_n771));
  NAND3_X1  g0571(.A1(new_n760), .A2(new_n294), .A3(G200), .ZN(new_n772));
  INV_X1    g0572(.A(G303), .ZN(new_n773));
  NAND3_X1  g0573(.A1(new_n760), .A2(G190), .A3(G200), .ZN(new_n774));
  OAI221_X1 g0574(.A(new_n770), .B1(new_n771), .B2(new_n772), .C1(new_n773), .C2(new_n774), .ZN(new_n775));
  NOR3_X1   g0575(.A1(new_n759), .A2(new_n765), .A3(new_n775), .ZN(new_n776));
  XOR2_X1   g0576(.A(new_n752), .B(KEYINPUT91), .Z(new_n777));
  NAND2_X1  g0577(.A1(new_n777), .A2(G97), .ZN(new_n778));
  OAI22_X1  g0578(.A1(new_n757), .A2(new_n207), .B1(new_n772), .B2(new_n505), .ZN(new_n779));
  INV_X1    g0579(.A(new_n766), .ZN(new_n780));
  OAI22_X1  g0580(.A1(new_n780), .A2(new_n243), .B1(new_n774), .B2(new_n571), .ZN(new_n781));
  NOR2_X1   g0581(.A1(new_n779), .A2(new_n781), .ZN(new_n782));
  INV_X1    g0582(.A(G159), .ZN(new_n783));
  NOR2_X1   g0583(.A1(new_n761), .A2(new_n783), .ZN(new_n784));
  XNOR2_X1  g0584(.A(new_n784), .B(KEYINPUT32), .ZN(new_n785));
  OAI21_X1  g0585(.A(new_n283), .B1(new_n763), .B2(new_n213), .ZN(new_n786));
  AOI21_X1  g0586(.A(new_n786), .B1(G77), .B2(new_n750), .ZN(new_n787));
  AND4_X1   g0587(.A1(new_n778), .A2(new_n782), .A3(new_n785), .A4(new_n787), .ZN(new_n788));
  OAI21_X1  g0588(.A(new_n746), .B1(new_n776), .B2(new_n788), .ZN(new_n789));
  INV_X1    g0589(.A(new_n743), .ZN(new_n790));
  NAND3_X1  g0590(.A1(new_n222), .A2(G355), .A3(new_n283), .ZN(new_n791));
  NOR2_X1   g0591(.A1(new_n678), .A2(new_n391), .ZN(new_n792));
  OAI21_X1  g0592(.A(new_n792), .B1(G45), .B2(new_n228), .ZN(new_n793));
  NOR2_X1   g0593(.A1(new_n247), .A2(new_n465), .ZN(new_n794));
  OAI221_X1 g0594(.A(new_n791), .B1(G116), .B2(new_n222), .C1(new_n793), .C2(new_n794), .ZN(new_n795));
  NOR2_X1   g0595(.A1(G13), .A2(G33), .ZN(new_n796));
  INV_X1    g0596(.A(new_n796), .ZN(new_n797));
  NOR2_X1   g0597(.A1(new_n797), .A2(G20), .ZN(new_n798));
  NOR2_X1   g0598(.A1(new_n798), .A2(new_n746), .ZN(new_n799));
  AOI21_X1  g0599(.A(new_n790), .B1(new_n795), .B2(new_n799), .ZN(new_n800));
  INV_X1    g0600(.A(new_n798), .ZN(new_n801));
  OAI211_X1 g0601(.A(new_n789), .B(new_n800), .C1(new_n662), .C2(new_n801), .ZN(new_n802));
  NAND2_X1  g0602(.A1(new_n745), .A2(new_n802), .ZN(G396));
  NAND2_X1  g0603(.A1(new_n645), .A2(new_n668), .ZN(new_n804));
  INV_X1    g0604(.A(new_n804), .ZN(new_n805));
  NAND2_X1  g0605(.A1(new_n313), .A2(new_n658), .ZN(new_n806));
  NAND2_X1  g0606(.A1(new_n332), .A2(new_n806), .ZN(new_n807));
  AOI21_X1  g0607(.A(new_n805), .B1(new_n336), .B2(new_n807), .ZN(new_n808));
  INV_X1    g0608(.A(new_n808), .ZN(new_n809));
  NAND3_X1  g0609(.A1(new_n685), .A2(new_n688), .A3(new_n809), .ZN(new_n810));
  OAI211_X1 g0610(.A(new_n668), .B(new_n808), .C1(new_n640), .C2(new_n630), .ZN(new_n811));
  NAND2_X1  g0611(.A1(new_n810), .A2(new_n811), .ZN(new_n812));
  AOI21_X1  g0612(.A(new_n743), .B1(new_n812), .B2(new_n732), .ZN(new_n813));
  OAI21_X1  g0613(.A(new_n813), .B1(new_n732), .B2(new_n812), .ZN(new_n814));
  INV_X1    g0614(.A(new_n746), .ZN(new_n815));
  NAND2_X1  g0615(.A1(new_n815), .A2(new_n797), .ZN(new_n816));
  OAI21_X1  g0616(.A(new_n743), .B1(G77), .B2(new_n816), .ZN(new_n817));
  XNOR2_X1  g0617(.A(new_n817), .B(KEYINPUT93), .ZN(new_n818));
  INV_X1    g0618(.A(new_n763), .ZN(new_n819));
  AOI22_X1  g0619(.A1(new_n819), .A2(G143), .B1(new_n750), .B2(G159), .ZN(new_n820));
  INV_X1    g0620(.A(G137), .ZN(new_n821));
  OAI221_X1 g0621(.A(new_n820), .B1(new_n757), .B2(new_n821), .C1(new_n260), .C2(new_n780), .ZN(new_n822));
  XNOR2_X1  g0622(.A(KEYINPUT94), .B(KEYINPUT34), .ZN(new_n823));
  OR2_X1    g0623(.A1(new_n822), .A2(new_n823), .ZN(new_n824));
  NAND2_X1  g0624(.A1(new_n822), .A2(new_n823), .ZN(new_n825));
  INV_X1    g0625(.A(new_n761), .ZN(new_n826));
  AOI21_X1  g0626(.A(new_n349), .B1(G132), .B2(new_n826), .ZN(new_n827));
  NOR2_X1   g0627(.A1(new_n774), .A2(new_n207), .ZN(new_n828));
  NOR2_X1   g0628(.A1(new_n772), .A2(new_n243), .ZN(new_n829));
  AOI211_X1 g0629(.A(new_n828), .B(new_n829), .C1(G58), .C2(new_n752), .ZN(new_n830));
  NAND4_X1  g0630(.A1(new_n824), .A2(new_n825), .A3(new_n827), .A4(new_n830), .ZN(new_n831));
  INV_X1    g0631(.A(G311), .ZN(new_n832));
  OAI22_X1  g0632(.A1(new_n763), .A2(new_n494), .B1(new_n761), .B2(new_n832), .ZN(new_n833));
  AOI211_X1 g0633(.A(new_n283), .B(new_n833), .C1(G116), .C2(new_n750), .ZN(new_n834));
  INV_X1    g0634(.A(new_n774), .ZN(new_n835));
  AOI22_X1  g0635(.A1(new_n756), .A2(G303), .B1(new_n835), .B2(G107), .ZN(new_n836));
  INV_X1    g0636(.A(new_n772), .ZN(new_n837));
  AOI22_X1  g0637(.A1(new_n766), .A2(G283), .B1(new_n837), .B2(G87), .ZN(new_n838));
  NAND4_X1  g0638(.A1(new_n834), .A2(new_n778), .A3(new_n836), .A4(new_n838), .ZN(new_n839));
  AND2_X1   g0639(.A1(new_n831), .A2(new_n839), .ZN(new_n840));
  OAI221_X1 g0640(.A(new_n818), .B1(new_n815), .B2(new_n840), .C1(new_n808), .C2(new_n797), .ZN(new_n841));
  NAND2_X1  g0641(.A1(new_n814), .A2(new_n841), .ZN(G384));
  INV_X1    g0642(.A(new_n583), .ZN(new_n843));
  OR2_X1    g0643(.A1(new_n843), .A2(KEYINPUT35), .ZN(new_n844));
  NAND2_X1  g0644(.A1(new_n843), .A2(KEYINPUT35), .ZN(new_n845));
  NAND4_X1  g0645(.A1(new_n844), .A2(G116), .A3(new_n227), .A4(new_n845), .ZN(new_n846));
  XNOR2_X1  g0646(.A(KEYINPUT95), .B(KEYINPUT36), .ZN(new_n847));
  XNOR2_X1  g0647(.A(new_n846), .B(new_n847), .ZN(new_n848));
  OR3_X1    g0648(.A1(new_n228), .A2(new_n289), .A3(new_n339), .ZN(new_n849));
  AOI211_X1 g0649(.A(new_n249), .B(G13), .C1(new_n849), .C2(new_n242), .ZN(new_n850));
  NOR2_X1   g0650(.A1(new_n848), .A2(new_n850), .ZN(new_n851));
  NAND2_X1  g0651(.A1(new_n811), .A2(new_n804), .ZN(new_n852));
  OAI211_X1 g0652(.A(new_n439), .B(new_n658), .C1(new_n438), .C2(new_n432), .ZN(new_n853));
  NAND2_X1  g0653(.A1(new_n437), .A2(new_n435), .ZN(new_n854));
  AOI21_X1  g0654(.A(new_n436), .B1(new_n419), .B2(G169), .ZN(new_n855));
  OAI21_X1  g0655(.A(new_n439), .B1(new_n854), .B2(new_n855), .ZN(new_n856));
  NOR2_X1   g0656(.A1(new_n429), .A2(new_n668), .ZN(new_n857));
  INV_X1    g0657(.A(new_n857), .ZN(new_n858));
  NAND3_X1  g0658(.A1(new_n856), .A2(new_n431), .A3(new_n858), .ZN(new_n859));
  NAND2_X1  g0659(.A1(new_n853), .A2(new_n859), .ZN(new_n860));
  NAND2_X1  g0660(.A1(new_n852), .A2(new_n860), .ZN(new_n861));
  INV_X1    g0661(.A(KEYINPUT96), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n861), .A2(new_n862), .ZN(new_n863));
  NAND3_X1  g0663(.A1(new_n852), .A2(KEYINPUT96), .A3(new_n860), .ZN(new_n864));
  INV_X1    g0664(.A(KEYINPUT38), .ZN(new_n865));
  NAND2_X1  g0665(.A1(new_n371), .A2(new_n388), .ZN(new_n866));
  NAND2_X1  g0666(.A1(new_n397), .A2(new_n398), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n866), .A2(new_n867), .ZN(new_n868));
  INV_X1    g0668(.A(KEYINPUT97), .ZN(new_n869));
  XNOR2_X1  g0669(.A(new_n656), .B(new_n869), .ZN(new_n870));
  INV_X1    g0670(.A(new_n870), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n866), .A2(new_n871), .ZN(new_n872));
  INV_X1    g0672(.A(KEYINPUT37), .ZN(new_n873));
  NAND4_X1  g0673(.A1(new_n868), .A2(new_n872), .A3(new_n873), .A4(new_n409), .ZN(new_n874));
  INV_X1    g0674(.A(KEYINPUT98), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n874), .A2(new_n875), .ZN(new_n876));
  AND3_X1   g0676(.A1(new_n408), .A2(new_n371), .A3(new_n388), .ZN(new_n877));
  NOR2_X1   g0677(.A1(new_n877), .A2(new_n399), .ZN(new_n878));
  AOI21_X1  g0678(.A(new_n870), .B1(new_n371), .B2(new_n388), .ZN(new_n879));
  NOR2_X1   g0679(.A1(new_n879), .A2(KEYINPUT37), .ZN(new_n880));
  NAND3_X1  g0680(.A1(new_n878), .A2(KEYINPUT98), .A3(new_n880), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n356), .A2(new_n308), .ZN(new_n882));
  INV_X1    g0682(.A(new_n357), .ZN(new_n883));
  OAI21_X1  g0683(.A(KEYINPUT7), .B1(new_n391), .B2(G20), .ZN(new_n884));
  NAND3_X1  g0684(.A1(new_n884), .A2(G68), .A3(new_n354), .ZN(new_n885));
  AOI21_X1  g0685(.A(new_n883), .B1(new_n885), .B2(new_n345), .ZN(new_n886));
  OAI211_X1 g0686(.A(new_n386), .B(new_n379), .C1(new_n882), .C2(new_n886), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n887), .A2(new_n867), .ZN(new_n888));
  INV_X1    g0688(.A(new_n656), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n887), .A2(new_n889), .ZN(new_n890));
  NAND3_X1  g0690(.A1(new_n888), .A2(new_n890), .A3(new_n409), .ZN(new_n891));
  AOI22_X1  g0691(.A1(new_n876), .A2(new_n881), .B1(KEYINPUT37), .B2(new_n891), .ZN(new_n892));
  AOI21_X1  g0692(.A(new_n890), .B1(new_n644), .B2(new_n648), .ZN(new_n893));
  OAI21_X1  g0693(.A(new_n865), .B1(new_n892), .B2(new_n893), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n891), .A2(KEYINPUT37), .ZN(new_n895));
  NOR2_X1   g0695(.A1(new_n874), .A2(new_n875), .ZN(new_n896));
  AOI21_X1  g0696(.A(KEYINPUT98), .B1(new_n878), .B2(new_n880), .ZN(new_n897));
  OAI21_X1  g0697(.A(new_n895), .B1(new_n896), .B2(new_n897), .ZN(new_n898));
  OAI211_X1 g0698(.A(new_n889), .B(new_n887), .C1(new_n401), .C2(new_n411), .ZN(new_n899));
  NAND3_X1  g0699(.A1(new_n898), .A2(KEYINPUT38), .A3(new_n899), .ZN(new_n900));
  NAND3_X1  g0700(.A1(new_n894), .A2(new_n900), .A3(KEYINPUT99), .ZN(new_n901));
  INV_X1    g0701(.A(KEYINPUT99), .ZN(new_n902));
  OAI211_X1 g0702(.A(new_n902), .B(new_n865), .C1(new_n892), .C2(new_n893), .ZN(new_n903));
  AND3_X1   g0703(.A1(new_n901), .A2(KEYINPUT100), .A3(new_n903), .ZN(new_n904));
  AOI21_X1  g0704(.A(KEYINPUT100), .B1(new_n901), .B2(new_n903), .ZN(new_n905));
  OAI211_X1 g0705(.A(new_n863), .B(new_n864), .C1(new_n904), .C2(new_n905), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n401), .A2(new_n870), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  INV_X1    g0708(.A(KEYINPUT101), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  NAND3_X1  g0710(.A1(new_n438), .A2(new_n439), .A3(new_n668), .ZN(new_n911));
  INV_X1    g0711(.A(new_n911), .ZN(new_n912));
  OAI21_X1  g0712(.A(KEYINPUT103), .B1(new_n896), .B2(new_n897), .ZN(new_n913));
  INV_X1    g0713(.A(KEYINPUT103), .ZN(new_n914));
  NAND3_X1  g0714(.A1(new_n876), .A2(new_n914), .A3(new_n881), .ZN(new_n915));
  NAND3_X1  g0715(.A1(new_n868), .A2(new_n872), .A3(new_n409), .ZN(new_n916));
  INV_X1    g0716(.A(KEYINPUT102), .ZN(new_n917));
  NAND3_X1  g0717(.A1(new_n916), .A2(new_n917), .A3(KEYINPUT37), .ZN(new_n918));
  NOR3_X1   g0718(.A1(new_n877), .A2(new_n399), .A3(new_n879), .ZN(new_n919));
  OAI21_X1  g0719(.A(KEYINPUT102), .B1(new_n919), .B2(new_n873), .ZN(new_n920));
  NAND4_X1  g0720(.A1(new_n913), .A2(new_n915), .A3(new_n918), .A4(new_n920), .ZN(new_n921));
  NOR2_X1   g0721(.A1(new_n412), .A2(new_n872), .ZN(new_n922));
  INV_X1    g0722(.A(new_n922), .ZN(new_n923));
  AOI21_X1  g0723(.A(KEYINPUT38), .B1(new_n921), .B2(new_n923), .ZN(new_n924));
  INV_X1    g0724(.A(new_n900), .ZN(new_n925));
  NOR3_X1   g0725(.A1(new_n924), .A2(KEYINPUT39), .A3(new_n925), .ZN(new_n926));
  AND3_X1   g0726(.A1(new_n901), .A2(KEYINPUT39), .A3(new_n903), .ZN(new_n927));
  OAI21_X1  g0727(.A(new_n912), .B1(new_n926), .B2(new_n927), .ZN(new_n928));
  NAND3_X1  g0728(.A1(new_n906), .A2(KEYINPUT101), .A3(new_n907), .ZN(new_n929));
  NAND3_X1  g0729(.A1(new_n910), .A2(new_n928), .A3(new_n929), .ZN(new_n930));
  NAND4_X1  g0730(.A1(new_n691), .A2(new_n617), .A3(new_n706), .A4(new_n707), .ZN(new_n931));
  AND2_X1   g0731(.A1(new_n931), .A2(new_n651), .ZN(new_n932));
  XOR2_X1   g0732(.A(new_n930), .B(new_n932), .Z(new_n933));
  INV_X1    g0733(.A(G330), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n921), .A2(new_n923), .ZN(new_n935));
  AOI21_X1  g0735(.A(new_n925), .B1(new_n935), .B2(new_n865), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n728), .A2(new_n658), .ZN(new_n937));
  NOR4_X1   g0737(.A1(new_n615), .A2(new_n485), .A3(new_n533), .A4(new_n658), .ZN(new_n938));
  INV_X1    g0738(.A(KEYINPUT31), .ZN(new_n939));
  OAI21_X1  g0739(.A(new_n937), .B1(new_n938), .B2(new_n939), .ZN(new_n940));
  NAND3_X1  g0740(.A1(new_n728), .A2(KEYINPUT31), .A3(new_n658), .ZN(new_n941));
  NAND2_X1  g0741(.A1(new_n940), .A2(new_n941), .ZN(new_n942));
  AOI21_X1  g0742(.A(new_n809), .B1(new_n859), .B2(new_n853), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n942), .A2(new_n943), .ZN(new_n944));
  INV_X1    g0744(.A(KEYINPUT40), .ZN(new_n945));
  NOR3_X1   g0745(.A1(new_n936), .A2(new_n944), .A3(new_n945), .ZN(new_n946));
  INV_X1    g0746(.A(new_n944), .ZN(new_n947));
  OAI21_X1  g0747(.A(new_n947), .B1(new_n904), .B2(new_n905), .ZN(new_n948));
  AOI21_X1  g0748(.A(new_n946), .B1(new_n948), .B2(new_n945), .ZN(new_n949));
  AOI21_X1  g0749(.A(new_n441), .B1(new_n940), .B2(new_n941), .ZN(new_n950));
  AOI21_X1  g0750(.A(new_n934), .B1(new_n949), .B2(new_n950), .ZN(new_n951));
  OAI21_X1  g0751(.A(new_n951), .B1(new_n950), .B2(new_n949), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n933), .A2(new_n952), .ZN(new_n953));
  OAI21_X1  g0753(.A(new_n953), .B1(new_n249), .B2(new_n738), .ZN(new_n954));
  NOR2_X1   g0754(.A1(new_n933), .A2(new_n952), .ZN(new_n955));
  OAI21_X1  g0755(.A(new_n851), .B1(new_n954), .B2(new_n955), .ZN(G367));
  INV_X1    g0756(.A(new_n792), .ZN(new_n957));
  NOR2_X1   g0757(.A1(new_n957), .A2(new_n237), .ZN(new_n958));
  OAI21_X1  g0758(.A(new_n799), .B1(new_n222), .B2(new_n301), .ZN(new_n959));
  OAI21_X1  g0759(.A(new_n743), .B1(new_n958), .B2(new_n959), .ZN(new_n960));
  OAI22_X1  g0760(.A1(new_n763), .A2(new_n260), .B1(new_n749), .B2(new_n207), .ZN(new_n961));
  AOI211_X1 g0761(.A(new_n460), .B(new_n961), .C1(G137), .C2(new_n826), .ZN(new_n962));
  NAND2_X1  g0762(.A1(new_n777), .A2(G68), .ZN(new_n963));
  AOI22_X1  g0763(.A1(new_n766), .A2(G159), .B1(new_n756), .B2(G143), .ZN(new_n964));
  NOR2_X1   g0764(.A1(new_n772), .A2(new_n289), .ZN(new_n965));
  AOI21_X1  g0765(.A(new_n965), .B1(G58), .B2(new_n835), .ZN(new_n966));
  NAND4_X1  g0766(.A1(new_n962), .A2(new_n963), .A3(new_n964), .A4(new_n966), .ZN(new_n967));
  OAI22_X1  g0767(.A1(new_n757), .A2(new_n832), .B1(new_n772), .B2(new_n215), .ZN(new_n968));
  AOI21_X1  g0768(.A(new_n968), .B1(G294), .B2(new_n766), .ZN(new_n969));
  OAI22_X1  g0769(.A1(new_n763), .A2(new_n773), .B1(new_n749), .B2(new_n771), .ZN(new_n970));
  AOI21_X1  g0770(.A(new_n970), .B1(G317), .B2(new_n826), .ZN(new_n971));
  AOI21_X1  g0771(.A(new_n391), .B1(G107), .B2(new_n752), .ZN(new_n972));
  NAND3_X1  g0772(.A1(new_n969), .A2(new_n971), .A3(new_n972), .ZN(new_n973));
  NOR2_X1   g0773(.A1(new_n774), .A2(new_n209), .ZN(new_n974));
  XNOR2_X1  g0774(.A(new_n974), .B(KEYINPUT46), .ZN(new_n975));
  OAI21_X1  g0775(.A(new_n967), .B1(new_n973), .B2(new_n975), .ZN(new_n976));
  XOR2_X1   g0776(.A(KEYINPUT107), .B(KEYINPUT47), .Z(new_n977));
  XNOR2_X1  g0777(.A(new_n976), .B(new_n977), .ZN(new_n978));
  AOI21_X1  g0778(.A(new_n960), .B1(new_n978), .B2(new_n746), .ZN(new_n979));
  OR3_X1    g0779(.A1(new_n626), .A2(new_n577), .A3(new_n668), .ZN(new_n980));
  OAI211_X1 g0780(.A(new_n626), .B(new_n627), .C1(new_n577), .C2(new_n668), .ZN(new_n981));
  NAND2_X1  g0781(.A1(new_n980), .A2(new_n981), .ZN(new_n982));
  OAI21_X1  g0782(.A(new_n979), .B1(new_n982), .B2(new_n801), .ZN(new_n983));
  NAND2_X1  g0783(.A1(new_n589), .A2(new_n658), .ZN(new_n984));
  NAND3_X1  g0784(.A1(new_n702), .A2(new_n703), .A3(new_n984), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n635), .A2(new_n658), .ZN(new_n986));
  NAND2_X1  g0786(.A1(new_n985), .A2(new_n986), .ZN(new_n987));
  NAND3_X1  g0787(.A1(new_n670), .A2(new_n675), .A3(new_n987), .ZN(new_n988));
  AND2_X1   g0788(.A1(new_n988), .A2(KEYINPUT42), .ZN(new_n989));
  OR2_X1    g0789(.A1(new_n985), .A2(new_n527), .ZN(new_n990));
  AOI21_X1  g0790(.A(new_n658), .B1(new_n990), .B2(new_n614), .ZN(new_n991));
  NOR3_X1   g0791(.A1(new_n989), .A2(KEYINPUT105), .A3(new_n991), .ZN(new_n992));
  NOR2_X1   g0792(.A1(new_n988), .A2(KEYINPUT42), .ZN(new_n993));
  NOR2_X1   g0793(.A1(new_n992), .A2(new_n993), .ZN(new_n994));
  OAI21_X1  g0794(.A(KEYINPUT105), .B1(new_n989), .B2(new_n991), .ZN(new_n995));
  NAND2_X1  g0795(.A1(new_n994), .A2(new_n995), .ZN(new_n996));
  INV_X1    g0796(.A(new_n982), .ZN(new_n997));
  NAND2_X1  g0797(.A1(new_n997), .A2(KEYINPUT104), .ZN(new_n998));
  INV_X1    g0798(.A(KEYINPUT104), .ZN(new_n999));
  AOI21_X1  g0799(.A(KEYINPUT43), .B1(new_n982), .B2(new_n999), .ZN(new_n1000));
  NAND2_X1  g0800(.A1(new_n998), .A2(new_n1000), .ZN(new_n1001));
  INV_X1    g0801(.A(KEYINPUT43), .ZN(new_n1002));
  OAI21_X1  g0802(.A(new_n1001), .B1(new_n1002), .B2(new_n997), .ZN(new_n1003));
  INV_X1    g0803(.A(new_n1003), .ZN(new_n1004));
  NAND2_X1  g0804(.A1(new_n996), .A2(new_n1004), .ZN(new_n1005));
  NAND4_X1  g0805(.A1(new_n994), .A2(new_n995), .A3(new_n998), .A4(new_n1000), .ZN(new_n1006));
  NAND2_X1  g0806(.A1(new_n1005), .A2(new_n1006), .ZN(new_n1007));
  INV_X1    g0807(.A(new_n987), .ZN(new_n1008));
  NOR2_X1   g0808(.A1(new_n673), .A2(new_n1008), .ZN(new_n1009));
  INV_X1    g0809(.A(new_n1009), .ZN(new_n1010));
  NAND2_X1  g0810(.A1(new_n1007), .A2(new_n1010), .ZN(new_n1011));
  NAND3_X1  g0811(.A1(new_n1005), .A2(new_n1009), .A3(new_n1006), .ZN(new_n1012));
  NAND2_X1  g0812(.A1(new_n1011), .A2(new_n1012), .ZN(new_n1013));
  INV_X1    g0813(.A(KEYINPUT45), .ZN(new_n1014));
  NAND2_X1  g0814(.A1(new_n670), .A2(new_n675), .ZN(new_n1015));
  NAND2_X1  g0815(.A1(new_n620), .A2(new_n668), .ZN(new_n1016));
  NAND2_X1  g0816(.A1(new_n1015), .A2(new_n1016), .ZN(new_n1017));
  OAI21_X1  g0817(.A(new_n1014), .B1(new_n1017), .B2(new_n1008), .ZN(new_n1018));
  NAND3_X1  g0818(.A1(new_n676), .A2(KEYINPUT45), .A3(new_n987), .ZN(new_n1019));
  NAND2_X1  g0819(.A1(new_n1018), .A2(new_n1019), .ZN(new_n1020));
  NAND3_X1  g0820(.A1(new_n1017), .A2(KEYINPUT44), .A3(new_n1008), .ZN(new_n1021));
  INV_X1    g0821(.A(KEYINPUT44), .ZN(new_n1022));
  OAI21_X1  g0822(.A(new_n1022), .B1(new_n676), .B2(new_n987), .ZN(new_n1023));
  NAND2_X1  g0823(.A1(new_n1021), .A2(new_n1023), .ZN(new_n1024));
  NAND2_X1  g0824(.A1(new_n1020), .A2(new_n1024), .ZN(new_n1025));
  NAND2_X1  g0825(.A1(new_n1025), .A2(new_n672), .ZN(new_n1026));
  NAND3_X1  g0826(.A1(new_n1020), .A2(new_n673), .A3(new_n1024), .ZN(new_n1027));
  NAND2_X1  g0827(.A1(new_n1026), .A2(new_n1027), .ZN(new_n1028));
  INV_X1    g0828(.A(KEYINPUT106), .ZN(new_n1029));
  NAND2_X1  g0829(.A1(new_n1015), .A2(new_n1029), .ZN(new_n1030));
  XNOR2_X1  g0830(.A(new_n1030), .B(new_n663), .ZN(new_n1031));
  NOR2_X1   g0831(.A1(new_n670), .A2(new_n675), .ZN(new_n1032));
  INV_X1    g0832(.A(new_n1032), .ZN(new_n1033));
  XNOR2_X1  g0833(.A(new_n1031), .B(new_n1033), .ZN(new_n1034));
  OAI21_X1  g0834(.A(new_n734), .B1(new_n1028), .B2(new_n1034), .ZN(new_n1035));
  XOR2_X1   g0835(.A(new_n679), .B(KEYINPUT41), .Z(new_n1036));
  INV_X1    g0836(.A(new_n1036), .ZN(new_n1037));
  AOI21_X1  g0837(.A(new_n742), .B1(new_n1035), .B2(new_n1037), .ZN(new_n1038));
  OAI21_X1  g0838(.A(new_n983), .B1(new_n1013), .B2(new_n1038), .ZN(G387));
  NAND2_X1  g0839(.A1(new_n265), .A2(new_n207), .ZN(new_n1040));
  XNOR2_X1  g0840(.A(new_n1040), .B(KEYINPUT50), .ZN(new_n1041));
  INV_X1    g0841(.A(new_n1041), .ZN(new_n1042));
  AOI211_X1 g0842(.A(G45), .B(new_n680), .C1(G68), .C2(G77), .ZN(new_n1043));
  AOI21_X1  g0843(.A(new_n957), .B1(new_n1042), .B2(new_n1043), .ZN(new_n1044));
  OR2_X1    g0844(.A1(new_n1044), .A2(KEYINPUT108), .ZN(new_n1045));
  NAND2_X1  g0845(.A1(new_n1044), .A2(KEYINPUT108), .ZN(new_n1046));
  OAI211_X1 g0846(.A(new_n1045), .B(new_n1046), .C1(new_n465), .C2(new_n234), .ZN(new_n1047));
  NAND3_X1  g0847(.A1(new_n222), .A2(new_n283), .A3(new_n680), .ZN(new_n1048));
  OAI211_X1 g0848(.A(new_n1047), .B(new_n1048), .C1(G107), .C2(new_n222), .ZN(new_n1049));
  AOI21_X1  g0849(.A(new_n790), .B1(new_n1049), .B2(new_n799), .ZN(new_n1050));
  NAND2_X1  g0850(.A1(new_n777), .A2(new_n302), .ZN(new_n1051));
  OAI22_X1  g0851(.A1(new_n757), .A2(new_n783), .B1(new_n774), .B2(new_n289), .ZN(new_n1052));
  AOI21_X1  g0852(.A(new_n1052), .B1(new_n265), .B2(new_n766), .ZN(new_n1053));
  OAI22_X1  g0853(.A1(new_n749), .A2(new_n243), .B1(new_n761), .B2(new_n260), .ZN(new_n1054));
  AOI21_X1  g0854(.A(new_n1054), .B1(G50), .B2(new_n819), .ZN(new_n1055));
  AOI21_X1  g0855(.A(new_n349), .B1(G97), .B2(new_n837), .ZN(new_n1056));
  AND4_X1   g0856(.A1(new_n1051), .A2(new_n1053), .A3(new_n1055), .A4(new_n1056), .ZN(new_n1057));
  AOI22_X1  g0857(.A1(new_n819), .A2(G317), .B1(new_n750), .B2(G303), .ZN(new_n1058));
  OAI221_X1 g0858(.A(new_n1058), .B1(new_n757), .B2(new_n764), .C1(new_n832), .C2(new_n780), .ZN(new_n1059));
  INV_X1    g0859(.A(KEYINPUT48), .ZN(new_n1060));
  OR2_X1    g0860(.A1(new_n1059), .A2(new_n1060), .ZN(new_n1061));
  NAND2_X1  g0861(.A1(new_n1059), .A2(new_n1060), .ZN(new_n1062));
  AOI22_X1  g0862(.A1(new_n835), .A2(G294), .B1(new_n752), .B2(G283), .ZN(new_n1063));
  NAND3_X1  g0863(.A1(new_n1061), .A2(new_n1062), .A3(new_n1063), .ZN(new_n1064));
  XOR2_X1   g0864(.A(new_n1064), .B(KEYINPUT49), .Z(new_n1065));
  OR2_X1    g0865(.A1(new_n1065), .A2(KEYINPUT109), .ZN(new_n1066));
  OAI221_X1 g0866(.A(new_n349), .B1(new_n209), .B2(new_n772), .C1(new_n754), .C2(new_n761), .ZN(new_n1067));
  AOI21_X1  g0867(.A(new_n1067), .B1(new_n1065), .B2(KEYINPUT109), .ZN(new_n1068));
  AOI21_X1  g0868(.A(new_n1057), .B1(new_n1066), .B2(new_n1068), .ZN(new_n1069));
  OAI21_X1  g0869(.A(new_n1050), .B1(new_n1069), .B2(new_n815), .ZN(new_n1070));
  AOI21_X1  g0870(.A(new_n1070), .B1(new_n671), .B2(new_n798), .ZN(new_n1071));
  XNOR2_X1  g0871(.A(new_n1031), .B(new_n1032), .ZN(new_n1072));
  AOI21_X1  g0872(.A(new_n1071), .B1(new_n1072), .B2(new_n742), .ZN(new_n1073));
  OAI21_X1  g0873(.A(KEYINPUT110), .B1(new_n1072), .B2(new_n734), .ZN(new_n1074));
  NAND2_X1  g0874(.A1(new_n1072), .A2(new_n734), .ZN(new_n1075));
  NAND3_X1  g0875(.A1(new_n1074), .A2(new_n679), .A3(new_n1075), .ZN(new_n1076));
  NOR3_X1   g0876(.A1(new_n1072), .A2(KEYINPUT110), .A3(new_n734), .ZN(new_n1077));
  OAI21_X1  g0877(.A(new_n1073), .B1(new_n1076), .B2(new_n1077), .ZN(G393));
  NAND3_X1  g0878(.A1(new_n1026), .A2(new_n742), .A3(new_n1027), .ZN(new_n1079));
  NOR2_X1   g0879(.A1(new_n957), .A2(new_n241), .ZN(new_n1080));
  OAI21_X1  g0880(.A(new_n799), .B1(new_n222), .B2(new_n215), .ZN(new_n1081));
  OAI21_X1  g0881(.A(new_n743), .B1(new_n1080), .B2(new_n1081), .ZN(new_n1082));
  OAI22_X1  g0882(.A1(new_n757), .A2(new_n767), .B1(new_n832), .B2(new_n763), .ZN(new_n1083));
  XNOR2_X1  g0883(.A(new_n1083), .B(KEYINPUT52), .ZN(new_n1084));
  OAI221_X1 g0884(.A(new_n460), .B1(new_n749), .B2(new_n494), .C1(new_n505), .C2(new_n772), .ZN(new_n1085));
  NOR2_X1   g0885(.A1(new_n780), .A2(new_n773), .ZN(new_n1086));
  AOI211_X1 g0886(.A(new_n1085), .B(new_n1086), .C1(G116), .C2(new_n752), .ZN(new_n1087));
  AOI22_X1  g0887(.A1(new_n835), .A2(G283), .B1(new_n826), .B2(G322), .ZN(new_n1088));
  OR2_X1    g0888(.A1(new_n1088), .A2(KEYINPUT112), .ZN(new_n1089));
  NAND2_X1  g0889(.A1(new_n1088), .A2(KEYINPUT112), .ZN(new_n1090));
  NAND4_X1  g0890(.A1(new_n1084), .A2(new_n1087), .A3(new_n1089), .A4(new_n1090), .ZN(new_n1091));
  AOI22_X1  g0891(.A1(G150), .A2(new_n756), .B1(new_n819), .B2(G159), .ZN(new_n1092));
  XNOR2_X1  g0892(.A(new_n1092), .B(KEYINPUT111), .ZN(new_n1093));
  NAND2_X1  g0893(.A1(new_n1093), .A2(KEYINPUT51), .ZN(new_n1094));
  NAND2_X1  g0894(.A1(new_n777), .A2(G77), .ZN(new_n1095));
  AOI22_X1  g0895(.A1(new_n265), .A2(new_n750), .B1(new_n826), .B2(G143), .ZN(new_n1096));
  AND2_X1   g0896(.A1(new_n1096), .A2(new_n391), .ZN(new_n1097));
  OAI22_X1  g0897(.A1(new_n780), .A2(new_n207), .B1(new_n772), .B2(new_n571), .ZN(new_n1098));
  AOI21_X1  g0898(.A(new_n1098), .B1(G68), .B2(new_n835), .ZN(new_n1099));
  NAND4_X1  g0899(.A1(new_n1094), .A2(new_n1095), .A3(new_n1097), .A4(new_n1099), .ZN(new_n1100));
  NOR2_X1   g0900(.A1(new_n1093), .A2(KEYINPUT51), .ZN(new_n1101));
  OAI21_X1  g0901(.A(new_n1091), .B1(new_n1100), .B2(new_n1101), .ZN(new_n1102));
  AOI21_X1  g0902(.A(new_n1082), .B1(new_n1102), .B2(new_n746), .ZN(new_n1103));
  OAI21_X1  g0903(.A(new_n1103), .B1(new_n987), .B2(new_n801), .ZN(new_n1104));
  NAND2_X1  g0904(.A1(new_n1075), .A2(new_n1028), .ZN(new_n1105));
  INV_X1    g0905(.A(new_n1105), .ZN(new_n1106));
  OAI21_X1  g0906(.A(new_n679), .B1(new_n1075), .B2(new_n1028), .ZN(new_n1107));
  OAI211_X1 g0907(.A(new_n1079), .B(new_n1104), .C1(new_n1106), .C2(new_n1107), .ZN(G390));
  NAND2_X1  g0908(.A1(new_n861), .A2(new_n911), .ZN(new_n1109));
  NAND3_X1  g0909(.A1(new_n901), .A2(KEYINPUT39), .A3(new_n903), .ZN(new_n1110));
  INV_X1    g0910(.A(KEYINPUT39), .ZN(new_n1111));
  NAND2_X1  g0911(.A1(new_n920), .A2(new_n918), .ZN(new_n1112));
  AOI21_X1  g0912(.A(new_n914), .B1(new_n876), .B2(new_n881), .ZN(new_n1113));
  NOR2_X1   g0913(.A1(new_n1112), .A2(new_n1113), .ZN(new_n1114));
  AOI21_X1  g0914(.A(new_n922), .B1(new_n1114), .B2(new_n915), .ZN(new_n1115));
  OAI211_X1 g0915(.A(new_n1111), .B(new_n900), .C1(new_n1115), .C2(KEYINPUT38), .ZN(new_n1116));
  NAND3_X1  g0916(.A1(new_n1109), .A2(new_n1110), .A3(new_n1116), .ZN(new_n1117));
  OAI211_X1 g0917(.A(G330), .B(new_n808), .C1(new_n729), .C2(new_n731), .ZN(new_n1118));
  AND2_X1   g0918(.A1(new_n853), .A2(new_n859), .ZN(new_n1119));
  NOR2_X1   g0919(.A1(new_n1118), .A2(new_n1119), .ZN(new_n1120));
  AOI21_X1  g0920(.A(new_n934), .B1(new_n940), .B2(new_n941), .ZN(new_n1121));
  NAND3_X1  g0921(.A1(new_n1121), .A2(KEYINPUT113), .A3(new_n943), .ZN(new_n1122));
  NAND2_X1  g0922(.A1(new_n1120), .A2(new_n1122), .ZN(new_n1123));
  OAI21_X1  g0923(.A(new_n900), .B1(new_n1115), .B2(KEYINPUT38), .ZN(new_n1124));
  NAND2_X1  g0924(.A1(new_n807), .A2(new_n336), .ZN(new_n1125));
  AND4_X1   g0925(.A1(new_n697), .A2(new_n696), .A3(new_n702), .A4(new_n703), .ZN(new_n1126));
  NAND3_X1  g0926(.A1(new_n693), .A2(new_n626), .A3(new_n694), .ZN(new_n1127));
  OAI211_X1 g0927(.A(new_n668), .B(new_n1125), .C1(new_n1126), .C2(new_n1127), .ZN(new_n1128));
  NAND2_X1  g0928(.A1(new_n1128), .A2(new_n804), .ZN(new_n1129));
  NAND2_X1  g0929(.A1(new_n1129), .A2(new_n860), .ZN(new_n1130));
  NAND3_X1  g0930(.A1(new_n1124), .A2(new_n1130), .A3(new_n911), .ZN(new_n1131));
  AND3_X1   g0931(.A1(new_n1117), .A2(new_n1123), .A3(new_n1131), .ZN(new_n1132));
  INV_X1    g0932(.A(KEYINPUT113), .ZN(new_n1133));
  NAND3_X1  g0933(.A1(new_n1121), .A2(new_n1133), .A3(new_n943), .ZN(new_n1134));
  AOI21_X1  g0934(.A(new_n1134), .B1(new_n1117), .B2(new_n1131), .ZN(new_n1135));
  NOR2_X1   g0935(.A1(new_n1132), .A2(new_n1135), .ZN(new_n1136));
  AND2_X1   g0936(.A1(new_n1136), .A2(new_n742), .ZN(new_n1137));
  XOR2_X1   g0937(.A(KEYINPUT54), .B(G143), .Z(new_n1138));
  AOI22_X1  g0938(.A1(new_n819), .A2(G132), .B1(new_n750), .B2(new_n1138), .ZN(new_n1139));
  INV_X1    g0939(.A(G128), .ZN(new_n1140));
  OAI21_X1  g0940(.A(new_n1139), .B1(new_n1140), .B2(new_n757), .ZN(new_n1141));
  AOI21_X1  g0941(.A(new_n1141), .B1(G137), .B2(new_n766), .ZN(new_n1142));
  NAND2_X1  g0942(.A1(new_n835), .A2(G150), .ZN(new_n1143));
  XOR2_X1   g0943(.A(new_n1143), .B(KEYINPUT53), .Z(new_n1144));
  INV_X1    g0944(.A(new_n777), .ZN(new_n1145));
  OAI211_X1 g0945(.A(new_n1142), .B(new_n1144), .C1(new_n783), .C2(new_n1145), .ZN(new_n1146));
  AOI21_X1  g0946(.A(new_n460), .B1(new_n826), .B2(G125), .ZN(new_n1147));
  OAI21_X1  g0947(.A(new_n1147), .B1(new_n207), .B2(new_n772), .ZN(new_n1148));
  XOR2_X1   g0948(.A(new_n1148), .B(KEYINPUT116), .Z(new_n1149));
  AOI22_X1  g0949(.A1(new_n756), .A2(G283), .B1(new_n750), .B2(G97), .ZN(new_n1150));
  OAI21_X1  g0950(.A(new_n1150), .B1(new_n505), .B2(new_n780), .ZN(new_n1151));
  XNOR2_X1  g0951(.A(new_n1151), .B(KEYINPUT117), .ZN(new_n1152));
  OAI21_X1  g0952(.A(new_n460), .B1(new_n774), .B2(new_n571), .ZN(new_n1153));
  XNOR2_X1  g0953(.A(new_n1153), .B(KEYINPUT118), .ZN(new_n1154));
  OAI22_X1  g0954(.A1(new_n763), .A2(new_n209), .B1(new_n761), .B2(new_n494), .ZN(new_n1155));
  NOR2_X1   g0955(.A1(new_n1155), .A2(new_n829), .ZN(new_n1156));
  NAND3_X1  g0956(.A1(new_n1154), .A2(new_n1095), .A3(new_n1156), .ZN(new_n1157));
  OAI22_X1  g0957(.A1(new_n1146), .A2(new_n1149), .B1(new_n1152), .B2(new_n1157), .ZN(new_n1158));
  AND2_X1   g0958(.A1(new_n1158), .A2(new_n746), .ZN(new_n1159));
  OAI21_X1  g0959(.A(new_n743), .B1(new_n265), .B2(new_n816), .ZN(new_n1160));
  NOR2_X1   g0960(.A1(new_n926), .A2(new_n927), .ZN(new_n1161));
  AOI211_X1 g0961(.A(new_n1159), .B(new_n1160), .C1(new_n1161), .C2(new_n796), .ZN(new_n1162));
  NOR2_X1   g0962(.A1(new_n1137), .A2(new_n1162), .ZN(new_n1163));
  OAI21_X1  g0963(.A(KEYINPUT115), .B1(new_n1132), .B2(new_n1135), .ZN(new_n1164));
  INV_X1    g0964(.A(KEYINPUT115), .ZN(new_n1165));
  NAND3_X1  g0965(.A1(new_n1117), .A2(new_n1123), .A3(new_n1131), .ZN(new_n1166));
  AOI21_X1  g0966(.A(new_n1119), .B1(new_n1128), .B2(new_n804), .ZN(new_n1167));
  NOR3_X1   g0967(.A1(new_n936), .A2(new_n1167), .A3(new_n912), .ZN(new_n1168));
  AOI21_X1  g0968(.A(new_n1168), .B1(new_n1161), .B2(new_n1109), .ZN(new_n1169));
  OAI211_X1 g0969(.A(new_n1165), .B(new_n1166), .C1(new_n1169), .C2(new_n1134), .ZN(new_n1170));
  NAND2_X1  g0970(.A1(new_n1118), .A2(new_n1119), .ZN(new_n1171));
  NAND2_X1  g0971(.A1(new_n1121), .A2(new_n943), .ZN(new_n1172));
  AND2_X1   g0972(.A1(new_n1171), .A2(new_n1172), .ZN(new_n1173));
  INV_X1    g0973(.A(new_n852), .ZN(new_n1174));
  AOI21_X1  g0974(.A(new_n860), .B1(new_n1121), .B2(new_n808), .ZN(new_n1175));
  AOI21_X1  g0975(.A(new_n805), .B1(new_n705), .B2(new_n1125), .ZN(new_n1176));
  OAI21_X1  g0976(.A(new_n1176), .B1(new_n1118), .B2(new_n1119), .ZN(new_n1177));
  OAI22_X1  g0977(.A1(new_n1173), .A2(new_n1174), .B1(new_n1175), .B2(new_n1177), .ZN(new_n1178));
  NAND2_X1  g0978(.A1(new_n617), .A2(new_n1121), .ZN(new_n1179));
  NAND3_X1  g0979(.A1(new_n932), .A2(new_n1178), .A3(new_n1179), .ZN(new_n1180));
  NAND3_X1  g0980(.A1(new_n1164), .A2(new_n1170), .A3(new_n1180), .ZN(new_n1181));
  INV_X1    g0981(.A(new_n679), .ZN(new_n1182));
  NAND3_X1  g0982(.A1(new_n931), .A2(new_n651), .A3(new_n1179), .ZN(new_n1183));
  NOR2_X1   g0983(.A1(new_n1177), .A2(new_n1175), .ZN(new_n1184));
  AOI21_X1  g0984(.A(new_n1174), .B1(new_n1171), .B2(new_n1172), .ZN(new_n1185));
  NOR2_X1   g0985(.A1(new_n1184), .A2(new_n1185), .ZN(new_n1186));
  NOR2_X1   g0986(.A1(new_n1183), .A2(new_n1186), .ZN(new_n1187));
  AOI21_X1  g0987(.A(new_n1182), .B1(new_n1136), .B2(new_n1187), .ZN(new_n1188));
  OAI21_X1  g0988(.A(new_n1181), .B1(new_n1188), .B2(KEYINPUT114), .ZN(new_n1189));
  INV_X1    g0989(.A(KEYINPUT114), .ZN(new_n1190));
  AOI211_X1 g0990(.A(new_n1190), .B(new_n1182), .C1(new_n1136), .C2(new_n1187), .ZN(new_n1191));
  OAI21_X1  g0991(.A(new_n1163), .B1(new_n1189), .B2(new_n1191), .ZN(G378));
  NAND2_X1  g0992(.A1(new_n929), .A2(new_n928), .ZN(new_n1193));
  AOI21_X1  g0993(.A(KEYINPUT101), .B1(new_n906), .B2(new_n907), .ZN(new_n1194));
  OAI21_X1  g0994(.A(KEYINPUT120), .B1(new_n1193), .B2(new_n1194), .ZN(new_n1195));
  NAND3_X1  g0995(.A1(new_n947), .A2(new_n1124), .A3(KEYINPUT40), .ZN(new_n1196));
  NAND2_X1  g0996(.A1(new_n901), .A2(new_n903), .ZN(new_n1197));
  INV_X1    g0997(.A(KEYINPUT100), .ZN(new_n1198));
  NAND2_X1  g0998(.A1(new_n1197), .A2(new_n1198), .ZN(new_n1199));
  NAND3_X1  g0999(.A1(new_n901), .A2(KEYINPUT100), .A3(new_n903), .ZN(new_n1200));
  AOI21_X1  g1000(.A(new_n944), .B1(new_n1199), .B2(new_n1200), .ZN(new_n1201));
  OAI211_X1 g1001(.A(G330), .B(new_n1196), .C1(new_n1201), .C2(KEYINPUT40), .ZN(new_n1202));
  NAND2_X1  g1002(.A1(new_n296), .A2(new_n300), .ZN(new_n1203));
  NAND2_X1  g1003(.A1(new_n270), .A2(new_n889), .ZN(new_n1204));
  XNOR2_X1  g1004(.A(new_n1203), .B(new_n1204), .ZN(new_n1205));
  XNOR2_X1  g1005(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1206));
  XNOR2_X1  g1006(.A(new_n1205), .B(new_n1206), .ZN(new_n1207));
  INV_X1    g1007(.A(new_n1207), .ZN(new_n1208));
  NAND2_X1  g1008(.A1(new_n1202), .A2(new_n1208), .ZN(new_n1209));
  NAND3_X1  g1009(.A1(new_n949), .A2(G330), .A3(new_n1207), .ZN(new_n1210));
  NAND2_X1  g1010(.A1(new_n1209), .A2(new_n1210), .ZN(new_n1211));
  NAND2_X1  g1011(.A1(new_n1195), .A2(new_n1211), .ZN(new_n1212));
  NAND4_X1  g1012(.A1(new_n930), .A2(KEYINPUT120), .A3(new_n1210), .A4(new_n1209), .ZN(new_n1213));
  INV_X1    g1013(.A(KEYINPUT121), .ZN(new_n1214));
  NAND2_X1  g1014(.A1(new_n1183), .A2(new_n1214), .ZN(new_n1215));
  NAND3_X1  g1015(.A1(new_n932), .A2(KEYINPUT121), .A3(new_n1179), .ZN(new_n1216));
  OAI21_X1  g1016(.A(new_n1166), .B1(new_n1169), .B2(new_n1134), .ZN(new_n1217));
  OAI211_X1 g1017(.A(new_n1215), .B(new_n1216), .C1(new_n1180), .C2(new_n1217), .ZN(new_n1218));
  NAND3_X1  g1018(.A1(new_n1212), .A2(new_n1213), .A3(new_n1218), .ZN(new_n1219));
  INV_X1    g1019(.A(KEYINPUT57), .ZN(new_n1220));
  NAND2_X1  g1020(.A1(new_n1219), .A2(new_n1220), .ZN(new_n1221));
  NOR2_X1   g1021(.A1(new_n1202), .A2(new_n1208), .ZN(new_n1222));
  AOI21_X1  g1022(.A(new_n1207), .B1(new_n949), .B2(G330), .ZN(new_n1223));
  OAI22_X1  g1023(.A1(new_n1222), .A2(new_n1223), .B1(new_n1194), .B2(new_n1193), .ZN(new_n1224));
  AND2_X1   g1024(.A1(new_n929), .A2(new_n928), .ZN(new_n1225));
  NAND4_X1  g1025(.A1(new_n1225), .A2(new_n1209), .A3(new_n1210), .A4(new_n910), .ZN(new_n1226));
  NAND2_X1  g1026(.A1(new_n1224), .A2(new_n1226), .ZN(new_n1227));
  XNOR2_X1  g1027(.A(new_n1183), .B(KEYINPUT121), .ZN(new_n1228));
  NAND2_X1  g1028(.A1(new_n1136), .A2(new_n1187), .ZN(new_n1229));
  AOI21_X1  g1029(.A(new_n1220), .B1(new_n1228), .B2(new_n1229), .ZN(new_n1230));
  AOI21_X1  g1030(.A(new_n1182), .B1(new_n1227), .B2(new_n1230), .ZN(new_n1231));
  NAND2_X1  g1031(.A1(new_n1221), .A2(new_n1231), .ZN(new_n1232));
  NAND3_X1  g1032(.A1(new_n1212), .A2(new_n1213), .A3(new_n742), .ZN(new_n1233));
  NAND2_X1  g1033(.A1(new_n1208), .A2(new_n796), .ZN(new_n1234));
  OAI21_X1  g1034(.A(new_n743), .B1(G50), .B2(new_n816), .ZN(new_n1235));
  AOI22_X1  g1035(.A1(new_n819), .A2(G107), .B1(new_n750), .B2(new_n302), .ZN(new_n1236));
  OAI21_X1  g1036(.A(new_n1236), .B1(new_n771), .B2(new_n761), .ZN(new_n1237));
  NOR3_X1   g1037(.A1(new_n1237), .A2(G41), .A3(new_n391), .ZN(new_n1238));
  AOI22_X1  g1038(.A1(new_n835), .A2(G77), .B1(new_n837), .B2(G58), .ZN(new_n1239));
  AOI22_X1  g1039(.A1(new_n766), .A2(G97), .B1(new_n756), .B2(G116), .ZN(new_n1240));
  NAND4_X1  g1040(.A1(new_n1238), .A2(new_n963), .A3(new_n1239), .A4(new_n1240), .ZN(new_n1241));
  INV_X1    g1041(.A(KEYINPUT58), .ZN(new_n1242));
  NAND2_X1  g1042(.A1(new_n1241), .A2(new_n1242), .ZN(new_n1243));
  NOR2_X1   g1043(.A1(G33), .A2(G41), .ZN(new_n1244));
  XNOR2_X1  g1044(.A(new_n1244), .B(KEYINPUT119), .ZN(new_n1245));
  OAI211_X1 g1045(.A(new_n207), .B(new_n1245), .C1(new_n391), .C2(G41), .ZN(new_n1246));
  AND2_X1   g1046(.A1(new_n1243), .A2(new_n1246), .ZN(new_n1247));
  OAI22_X1  g1047(.A1(new_n763), .A2(new_n1140), .B1(new_n749), .B2(new_n821), .ZN(new_n1248));
  AOI21_X1  g1048(.A(new_n1248), .B1(G132), .B2(new_n766), .ZN(new_n1249));
  AOI22_X1  g1049(.A1(new_n756), .A2(G125), .B1(new_n835), .B2(new_n1138), .ZN(new_n1250));
  OAI211_X1 g1050(.A(new_n1249), .B(new_n1250), .C1(new_n1145), .C2(new_n260), .ZN(new_n1251));
  NOR2_X1   g1051(.A1(new_n1251), .A2(KEYINPUT59), .ZN(new_n1252));
  NAND2_X1  g1052(.A1(new_n1251), .A2(KEYINPUT59), .ZN(new_n1253));
  AOI21_X1  g1053(.A(new_n1245), .B1(G124), .B2(new_n826), .ZN(new_n1254));
  OAI211_X1 g1054(.A(new_n1253), .B(new_n1254), .C1(new_n783), .C2(new_n772), .ZN(new_n1255));
  OAI221_X1 g1055(.A(new_n1247), .B1(new_n1242), .B2(new_n1241), .C1(new_n1252), .C2(new_n1255), .ZN(new_n1256));
  AOI21_X1  g1056(.A(new_n1235), .B1(new_n1256), .B2(new_n746), .ZN(new_n1257));
  NAND2_X1  g1057(.A1(new_n1234), .A2(new_n1257), .ZN(new_n1258));
  NAND2_X1  g1058(.A1(new_n1233), .A2(new_n1258), .ZN(new_n1259));
  INV_X1    g1059(.A(new_n1259), .ZN(new_n1260));
  NAND2_X1  g1060(.A1(new_n1232), .A2(new_n1260), .ZN(G375));
  NAND2_X1  g1061(.A1(new_n1183), .A2(new_n1186), .ZN(new_n1262));
  NAND3_X1  g1062(.A1(new_n1180), .A2(new_n1037), .A3(new_n1262), .ZN(new_n1263));
  OAI21_X1  g1063(.A(new_n743), .B1(G68), .B2(new_n816), .ZN(new_n1264));
  OAI22_X1  g1064(.A1(new_n763), .A2(new_n771), .B1(new_n749), .B2(new_n505), .ZN(new_n1265));
  AOI211_X1 g1065(.A(new_n283), .B(new_n1265), .C1(G303), .C2(new_n826), .ZN(new_n1266));
  AOI21_X1  g1066(.A(new_n965), .B1(G116), .B2(new_n766), .ZN(new_n1267));
  AOI22_X1  g1067(.A1(new_n756), .A2(G294), .B1(new_n835), .B2(G97), .ZN(new_n1268));
  NAND4_X1  g1068(.A1(new_n1266), .A2(new_n1051), .A3(new_n1267), .A4(new_n1268), .ZN(new_n1269));
  OAI21_X1  g1069(.A(new_n391), .B1(new_n213), .B2(new_n772), .ZN(new_n1270));
  XNOR2_X1  g1070(.A(new_n1270), .B(KEYINPUT122), .ZN(new_n1271));
  NAND2_X1  g1071(.A1(new_n777), .A2(G50), .ZN(new_n1272));
  OAI22_X1  g1072(.A1(new_n763), .A2(new_n821), .B1(new_n749), .B2(new_n260), .ZN(new_n1273));
  AOI21_X1  g1073(.A(new_n1273), .B1(G128), .B2(new_n826), .ZN(new_n1274));
  NAND2_X1  g1074(.A1(new_n756), .A2(G132), .ZN(new_n1275));
  AOI22_X1  g1075(.A1(new_n766), .A2(new_n1138), .B1(new_n835), .B2(G159), .ZN(new_n1276));
  NAND4_X1  g1076(.A1(new_n1272), .A2(new_n1274), .A3(new_n1275), .A4(new_n1276), .ZN(new_n1277));
  OAI21_X1  g1077(.A(new_n1269), .B1(new_n1271), .B2(new_n1277), .ZN(new_n1278));
  AOI21_X1  g1078(.A(new_n1264), .B1(new_n1278), .B2(new_n746), .ZN(new_n1279));
  OAI21_X1  g1079(.A(new_n1279), .B1(new_n860), .B2(new_n797), .ZN(new_n1280));
  INV_X1    g1080(.A(new_n742), .ZN(new_n1281));
  OAI21_X1  g1081(.A(new_n1280), .B1(new_n1186), .B2(new_n1281), .ZN(new_n1282));
  INV_X1    g1082(.A(new_n1282), .ZN(new_n1283));
  NAND2_X1  g1083(.A1(new_n1263), .A2(new_n1283), .ZN(G381));
  OR2_X1    g1084(.A1(G393), .A2(G396), .ZN(new_n1285));
  NAND2_X1  g1085(.A1(new_n1079), .A2(new_n1104), .ZN(new_n1286));
  INV_X1    g1086(.A(new_n1107), .ZN(new_n1287));
  AOI21_X1  g1087(.A(new_n1286), .B1(new_n1287), .B2(new_n1105), .ZN(new_n1288));
  INV_X1    g1088(.A(G384), .ZN(new_n1289));
  NAND2_X1  g1089(.A1(new_n1288), .A2(new_n1289), .ZN(new_n1290));
  NOR4_X1   g1090(.A1(new_n1285), .A2(new_n1290), .A3(G387), .A4(G381), .ZN(new_n1291));
  INV_X1    g1091(.A(G378), .ZN(new_n1292));
  AOI21_X1  g1092(.A(new_n1259), .B1(new_n1221), .B2(new_n1231), .ZN(new_n1293));
  NAND3_X1  g1093(.A1(new_n1291), .A2(new_n1292), .A3(new_n1293), .ZN(G407));
  INV_X1    g1094(.A(G213), .ZN(new_n1295));
  NOR2_X1   g1095(.A1(new_n1295), .A2(G343), .ZN(new_n1296));
  NAND3_X1  g1096(.A1(new_n1293), .A2(new_n1292), .A3(new_n1296), .ZN(new_n1297));
  NAND3_X1  g1097(.A1(G407), .A2(G213), .A3(new_n1297), .ZN(G409));
  OAI211_X1 g1098(.A(G390), .B(new_n983), .C1(new_n1038), .C2(new_n1013), .ZN(new_n1299));
  NAND2_X1  g1099(.A1(G387), .A2(new_n1288), .ZN(new_n1300));
  NAND2_X1  g1100(.A1(new_n1299), .A2(new_n1300), .ZN(new_n1301));
  NAND2_X1  g1101(.A1(G393), .A2(G396), .ZN(new_n1302));
  NAND2_X1  g1102(.A1(new_n1285), .A2(new_n1302), .ZN(new_n1303));
  NAND2_X1  g1103(.A1(new_n1301), .A2(new_n1303), .ZN(new_n1304));
  INV_X1    g1104(.A(KEYINPUT125), .ZN(new_n1305));
  NAND4_X1  g1105(.A1(new_n1299), .A2(new_n1300), .A3(new_n1285), .A4(new_n1302), .ZN(new_n1306));
  AND3_X1   g1106(.A1(new_n1304), .A2(new_n1305), .A3(new_n1306), .ZN(new_n1307));
  AOI21_X1  g1107(.A(new_n1305), .B1(new_n1304), .B2(new_n1306), .ZN(new_n1308));
  NOR2_X1   g1108(.A1(new_n1307), .A2(new_n1308), .ZN(new_n1309));
  INV_X1    g1109(.A(KEYINPUT60), .ZN(new_n1310));
  OAI21_X1  g1110(.A(new_n1262), .B1(new_n1187), .B2(new_n1310), .ZN(new_n1311));
  NAND3_X1  g1111(.A1(new_n1183), .A2(new_n1186), .A3(KEYINPUT60), .ZN(new_n1312));
  NAND3_X1  g1112(.A1(new_n1311), .A2(new_n679), .A3(new_n1312), .ZN(new_n1313));
  NAND3_X1  g1113(.A1(new_n1313), .A2(G384), .A3(new_n1283), .ZN(new_n1314));
  INV_X1    g1114(.A(new_n1314), .ZN(new_n1315));
  AOI21_X1  g1115(.A(G384), .B1(new_n1313), .B2(new_n1283), .ZN(new_n1316));
  NAND2_X1  g1116(.A1(new_n1296), .A2(G2897), .ZN(new_n1317));
  NOR3_X1   g1117(.A1(new_n1315), .A2(new_n1316), .A3(new_n1317), .ZN(new_n1318));
  INV_X1    g1118(.A(new_n1318), .ZN(new_n1319));
  OAI21_X1  g1119(.A(new_n1317), .B1(new_n1315), .B2(new_n1316), .ZN(new_n1320));
  NAND2_X1  g1120(.A1(new_n1319), .A2(new_n1320), .ZN(new_n1321));
  NAND4_X1  g1121(.A1(new_n1212), .A2(new_n1213), .A3(new_n1218), .A4(new_n1037), .ZN(new_n1322));
  AOI22_X1  g1122(.A1(new_n1227), .A2(new_n742), .B1(new_n1234), .B2(new_n1257), .ZN(new_n1323));
  AOI21_X1  g1123(.A(G378), .B1(new_n1322), .B2(new_n1323), .ZN(new_n1324));
  AOI21_X1  g1124(.A(new_n1324), .B1(G378), .B2(new_n1293), .ZN(new_n1325));
  OAI21_X1  g1125(.A(new_n1321), .B1(new_n1325), .B2(new_n1296), .ZN(new_n1326));
  INV_X1    g1126(.A(KEYINPUT61), .ZN(new_n1327));
  NAND3_X1  g1127(.A1(new_n1232), .A2(G378), .A3(new_n1260), .ZN(new_n1328));
  NAND2_X1  g1128(.A1(new_n1323), .A2(new_n1322), .ZN(new_n1329));
  NAND2_X1  g1129(.A1(new_n1329), .A2(new_n1292), .ZN(new_n1330));
  NAND2_X1  g1130(.A1(new_n1328), .A2(new_n1330), .ZN(new_n1331));
  INV_X1    g1131(.A(KEYINPUT62), .ZN(new_n1332));
  INV_X1    g1132(.A(new_n1296), .ZN(new_n1333));
  NOR2_X1   g1133(.A1(new_n1315), .A2(new_n1316), .ZN(new_n1334));
  NAND4_X1  g1134(.A1(new_n1331), .A2(new_n1332), .A3(new_n1333), .A4(new_n1334), .ZN(new_n1335));
  NAND3_X1  g1135(.A1(new_n1326), .A2(new_n1327), .A3(new_n1335), .ZN(new_n1336));
  XNOR2_X1  g1136(.A(KEYINPUT124), .B(KEYINPUT62), .ZN(new_n1337));
  AOI21_X1  g1137(.A(new_n1296), .B1(new_n1328), .B2(new_n1330), .ZN(new_n1338));
  AOI21_X1  g1138(.A(new_n1337), .B1(new_n1338), .B2(new_n1334), .ZN(new_n1339));
  OAI21_X1  g1139(.A(new_n1309), .B1(new_n1336), .B2(new_n1339), .ZN(new_n1340));
  INV_X1    g1140(.A(new_n1338), .ZN(new_n1341));
  NAND2_X1  g1141(.A1(new_n1321), .A2(KEYINPUT123), .ZN(new_n1342));
  INV_X1    g1142(.A(KEYINPUT123), .ZN(new_n1343));
  NAND3_X1  g1143(.A1(new_n1319), .A2(new_n1343), .A3(new_n1320), .ZN(new_n1344));
  NAND3_X1  g1144(.A1(new_n1341), .A2(new_n1342), .A3(new_n1344), .ZN(new_n1345));
  NAND2_X1  g1145(.A1(new_n1338), .A2(new_n1334), .ZN(new_n1346));
  INV_X1    g1146(.A(KEYINPUT63), .ZN(new_n1347));
  NAND2_X1  g1147(.A1(new_n1346), .A2(new_n1347), .ZN(new_n1348));
  AND3_X1   g1148(.A1(new_n1304), .A2(new_n1327), .A3(new_n1306), .ZN(new_n1349));
  NAND3_X1  g1149(.A1(new_n1338), .A2(KEYINPUT63), .A3(new_n1334), .ZN(new_n1350));
  NAND4_X1  g1150(.A1(new_n1345), .A2(new_n1348), .A3(new_n1349), .A4(new_n1350), .ZN(new_n1351));
  NAND2_X1  g1151(.A1(new_n1340), .A2(new_n1351), .ZN(G405));
  NAND2_X1  g1152(.A1(G375), .A2(new_n1292), .ZN(new_n1353));
  NAND2_X1  g1153(.A1(new_n1353), .A2(new_n1328), .ZN(new_n1354));
  NAND2_X1  g1154(.A1(new_n1334), .A2(KEYINPUT126), .ZN(new_n1355));
  OR2_X1    g1155(.A1(new_n1334), .A2(KEYINPUT126), .ZN(new_n1356));
  NAND3_X1  g1156(.A1(new_n1354), .A2(new_n1355), .A3(new_n1356), .ZN(new_n1357));
  AND2_X1   g1157(.A1(new_n1304), .A2(new_n1306), .ZN(new_n1358));
  NAND4_X1  g1158(.A1(new_n1353), .A2(KEYINPUT126), .A3(new_n1334), .A4(new_n1328), .ZN(new_n1359));
  AND3_X1   g1159(.A1(new_n1357), .A2(new_n1358), .A3(new_n1359), .ZN(new_n1360));
  AOI21_X1  g1160(.A(new_n1358), .B1(new_n1357), .B2(new_n1359), .ZN(new_n1361));
  NOR2_X1   g1161(.A1(new_n1360), .A2(new_n1361), .ZN(G402));
endmodule


