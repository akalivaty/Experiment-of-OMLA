//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 1 1 0 1 1 0 1 1 0 1 0 1 1 1 0 1 1 0 0 1 1 1 1 1 1 0 1 0 0 0 1 0 0 0 1 1 1 0 0 1 1 1 0 0 1 0 1 1 1 0 1 0 1 1 1 1 1 1 1 1 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:24:33 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n698, new_n699, new_n700, new_n701, new_n702, new_n703,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n715, new_n716, new_n718, new_n719, new_n720,
    new_n721, new_n723, new_n724, new_n725, new_n726, new_n727, new_n728,
    new_n729, new_n731, new_n732, new_n733, new_n734, new_n735, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n765, new_n766,
    new_n767, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n794, new_n795, new_n796,
    new_n797, new_n798, new_n799, new_n800, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n922, new_n923, new_n924, new_n925, new_n926, new_n927,
    new_n928, new_n929, new_n930, new_n931, new_n932, new_n933, new_n934,
    new_n936, new_n937, new_n938, new_n939, new_n940, new_n941, new_n942,
    new_n943, new_n944, new_n946, new_n947, new_n948, new_n949, new_n950,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n980,
    new_n981, new_n982, new_n983, new_n984, new_n985, new_n986, new_n987,
    new_n988, new_n989, new_n990, new_n991, new_n992, new_n993, new_n994,
    new_n995, new_n996;
  OAI21_X1  g000(.A(G210), .B1(G237), .B2(G902), .ZN(new_n187));
  INV_X1    g001(.A(G119), .ZN(new_n188));
  NAND2_X1  g002(.A1(new_n188), .A2(G116), .ZN(new_n189));
  INV_X1    g003(.A(G116), .ZN(new_n190));
  NAND2_X1  g004(.A1(new_n190), .A2(G119), .ZN(new_n191));
  NAND2_X1  g005(.A1(new_n189), .A2(new_n191), .ZN(new_n192));
  XNOR2_X1  g006(.A(KEYINPUT2), .B(G113), .ZN(new_n193));
  NOR2_X1   g007(.A1(new_n192), .A2(new_n193), .ZN(new_n194));
  NAND3_X1  g008(.A1(new_n189), .A2(new_n191), .A3(KEYINPUT5), .ZN(new_n195));
  INV_X1    g009(.A(KEYINPUT5), .ZN(new_n196));
  NAND3_X1  g010(.A1(new_n196), .A2(new_n188), .A3(G116), .ZN(new_n197));
  NAND3_X1  g011(.A1(new_n195), .A2(G113), .A3(new_n197), .ZN(new_n198));
  INV_X1    g012(.A(KEYINPUT82), .ZN(new_n199));
  AOI21_X1  g013(.A(new_n194), .B1(new_n198), .B2(new_n199), .ZN(new_n200));
  NAND4_X1  g014(.A1(new_n195), .A2(KEYINPUT82), .A3(G113), .A4(new_n197), .ZN(new_n201));
  INV_X1    g015(.A(G104), .ZN(new_n202));
  OAI21_X1  g016(.A(KEYINPUT3), .B1(new_n202), .B2(G107), .ZN(new_n203));
  INV_X1    g017(.A(KEYINPUT3), .ZN(new_n204));
  INV_X1    g018(.A(G107), .ZN(new_n205));
  NAND3_X1  g019(.A1(new_n204), .A2(new_n205), .A3(G104), .ZN(new_n206));
  INV_X1    g020(.A(G101), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n202), .A2(G107), .ZN(new_n208));
  NAND4_X1  g022(.A1(new_n203), .A2(new_n206), .A3(new_n207), .A4(new_n208), .ZN(new_n209));
  NOR2_X1   g023(.A1(new_n202), .A2(G107), .ZN(new_n210));
  NOR2_X1   g024(.A1(new_n205), .A2(G104), .ZN(new_n211));
  OAI21_X1  g025(.A(G101), .B1(new_n210), .B2(new_n211), .ZN(new_n212));
  INV_X1    g026(.A(KEYINPUT80), .ZN(new_n213));
  AND3_X1   g027(.A1(new_n209), .A2(new_n212), .A3(new_n213), .ZN(new_n214));
  AOI21_X1  g028(.A(new_n213), .B1(new_n209), .B2(new_n212), .ZN(new_n215));
  OAI211_X1 g029(.A(new_n200), .B(new_n201), .C1(new_n214), .C2(new_n215), .ZN(new_n216));
  XNOR2_X1  g030(.A(G110), .B(G122), .ZN(new_n217));
  NAND3_X1  g031(.A1(new_n203), .A2(new_n206), .A3(new_n208), .ZN(new_n218));
  INV_X1    g032(.A(KEYINPUT78), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n218), .A2(new_n219), .ZN(new_n220));
  NAND4_X1  g034(.A1(new_n203), .A2(new_n206), .A3(KEYINPUT78), .A4(new_n208), .ZN(new_n221));
  NAND3_X1  g035(.A1(new_n220), .A2(G101), .A3(new_n221), .ZN(new_n222));
  AND2_X1   g036(.A1(new_n209), .A2(KEYINPUT4), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n222), .A2(new_n223), .ZN(new_n224));
  INV_X1    g038(.A(new_n224), .ZN(new_n225));
  NOR2_X1   g039(.A1(new_n207), .A2(KEYINPUT4), .ZN(new_n226));
  NAND3_X1  g040(.A1(new_n220), .A2(new_n221), .A3(new_n226), .ZN(new_n227));
  INV_X1    g041(.A(KEYINPUT2), .ZN(new_n228));
  NOR2_X1   g042(.A1(new_n228), .A2(G113), .ZN(new_n229));
  INV_X1    g043(.A(G113), .ZN(new_n230));
  NOR2_X1   g044(.A1(new_n230), .A2(KEYINPUT2), .ZN(new_n231));
  OAI211_X1 g045(.A(new_n189), .B(new_n191), .C1(new_n229), .C2(new_n231), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n192), .A2(new_n193), .ZN(new_n233));
  AND3_X1   g047(.A1(new_n232), .A2(new_n233), .A3(KEYINPUT68), .ZN(new_n234));
  AOI21_X1  g048(.A(KEYINPUT68), .B1(new_n232), .B2(new_n233), .ZN(new_n235));
  OAI21_X1  g049(.A(new_n227), .B1(new_n234), .B2(new_n235), .ZN(new_n236));
  OAI211_X1 g050(.A(new_n216), .B(new_n217), .C1(new_n225), .C2(new_n236), .ZN(new_n237));
  INV_X1    g051(.A(KEYINPUT83), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n237), .A2(new_n238), .ZN(new_n239));
  INV_X1    g053(.A(new_n235), .ZN(new_n240));
  NAND3_X1  g054(.A1(new_n232), .A2(new_n233), .A3(KEYINPUT68), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n240), .A2(new_n241), .ZN(new_n242));
  NAND3_X1  g056(.A1(new_n242), .A2(new_n224), .A3(new_n227), .ZN(new_n243));
  NAND4_X1  g057(.A1(new_n243), .A2(KEYINPUT83), .A3(new_n216), .A4(new_n217), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n239), .A2(new_n244), .ZN(new_n245));
  INV_X1    g059(.A(KEYINPUT64), .ZN(new_n246));
  NAND3_X1  g060(.A1(new_n246), .A2(KEYINPUT0), .A3(G128), .ZN(new_n247));
  NAND2_X1  g061(.A1(KEYINPUT0), .A2(G128), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n248), .A2(KEYINPUT64), .ZN(new_n249));
  NOR2_X1   g063(.A1(KEYINPUT0), .A2(G128), .ZN(new_n250));
  OAI21_X1  g064(.A(new_n247), .B1(new_n249), .B2(new_n250), .ZN(new_n251));
  INV_X1    g065(.A(G143), .ZN(new_n252));
  OAI21_X1  g066(.A(KEYINPUT65), .B1(new_n252), .B2(G146), .ZN(new_n253));
  INV_X1    g067(.A(KEYINPUT65), .ZN(new_n254));
  INV_X1    g068(.A(G146), .ZN(new_n255));
  NAND3_X1  g069(.A1(new_n254), .A2(new_n255), .A3(G143), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n252), .A2(G146), .ZN(new_n257));
  NAND3_X1  g071(.A1(new_n253), .A2(new_n256), .A3(new_n257), .ZN(new_n258));
  XNOR2_X1  g072(.A(G143), .B(G146), .ZN(new_n259));
  INV_X1    g073(.A(new_n248), .ZN(new_n260));
  AOI22_X1  g074(.A1(new_n251), .A2(new_n258), .B1(new_n259), .B2(new_n260), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n261), .A2(G125), .ZN(new_n262));
  OAI21_X1  g076(.A(KEYINPUT1), .B1(new_n252), .B2(G146), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n263), .A2(G128), .ZN(new_n264));
  INV_X1    g078(.A(G128), .ZN(new_n265));
  NOR2_X1   g079(.A1(new_n265), .A2(KEYINPUT1), .ZN(new_n266));
  AOI22_X1  g080(.A1(new_n258), .A2(new_n264), .B1(new_n259), .B2(new_n266), .ZN(new_n267));
  OAI21_X1  g081(.A(new_n262), .B1(G125), .B2(new_n267), .ZN(new_n268));
  INV_X1    g082(.A(KEYINPUT85), .ZN(new_n269));
  INV_X1    g083(.A(G224), .ZN(new_n270));
  OAI21_X1  g084(.A(new_n269), .B1(new_n270), .B2(G953), .ZN(new_n271));
  INV_X1    g085(.A(G953), .ZN(new_n272));
  NAND3_X1  g086(.A1(new_n272), .A2(KEYINPUT85), .A3(G224), .ZN(new_n273));
  NAND3_X1  g087(.A1(new_n271), .A2(KEYINPUT7), .A3(new_n273), .ZN(new_n274));
  OR2_X1    g088(.A1(new_n268), .A2(new_n274), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n268), .A2(new_n274), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n209), .A2(new_n212), .ZN(new_n277));
  NAND3_X1  g091(.A1(new_n200), .A2(new_n277), .A3(new_n201), .ZN(new_n278));
  AOI21_X1  g092(.A(new_n277), .B1(new_n232), .B2(new_n198), .ZN(new_n279));
  XOR2_X1   g093(.A(new_n217), .B(KEYINPUT8), .Z(new_n280));
  NOR2_X1   g094(.A1(new_n279), .A2(new_n280), .ZN(new_n281));
  AOI22_X1  g095(.A1(new_n275), .A2(new_n276), .B1(new_n278), .B2(new_n281), .ZN(new_n282));
  AOI21_X1  g096(.A(G902), .B1(new_n245), .B2(new_n282), .ZN(new_n283));
  INV_X1    g097(.A(KEYINPUT86), .ZN(new_n284));
  AOI21_X1  g098(.A(new_n217), .B1(new_n243), .B2(new_n216), .ZN(new_n285));
  INV_X1    g099(.A(KEYINPUT6), .ZN(new_n286));
  NOR2_X1   g100(.A1(new_n285), .A2(new_n286), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n245), .A2(new_n287), .ZN(new_n288));
  AOI211_X1 g102(.A(KEYINPUT6), .B(new_n217), .C1(new_n243), .C2(new_n216), .ZN(new_n289));
  INV_X1    g103(.A(new_n289), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n271), .A2(new_n273), .ZN(new_n291));
  XNOR2_X1  g105(.A(new_n291), .B(KEYINPUT84), .ZN(new_n292));
  XNOR2_X1  g106(.A(new_n268), .B(new_n292), .ZN(new_n293));
  AND4_X1   g107(.A1(new_n284), .A2(new_n288), .A3(new_n290), .A4(new_n293), .ZN(new_n294));
  AOI21_X1  g108(.A(new_n289), .B1(new_n245), .B2(new_n287), .ZN(new_n295));
  AOI21_X1  g109(.A(new_n284), .B1(new_n295), .B2(new_n293), .ZN(new_n296));
  OAI211_X1 g110(.A(new_n187), .B(new_n283), .C1(new_n294), .C2(new_n296), .ZN(new_n297));
  INV_X1    g111(.A(KEYINPUT88), .ZN(new_n298));
  NAND2_X1  g112(.A1(new_n297), .A2(new_n298), .ZN(new_n299));
  OAI21_X1  g113(.A(new_n283), .B1(new_n294), .B2(new_n296), .ZN(new_n300));
  XOR2_X1   g114(.A(new_n187), .B(KEYINPUT87), .Z(new_n301));
  NAND2_X1  g115(.A1(new_n300), .A2(new_n301), .ZN(new_n302));
  NAND3_X1  g116(.A1(new_n288), .A2(new_n290), .A3(new_n293), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n303), .A2(KEYINPUT86), .ZN(new_n304));
  NAND3_X1  g118(.A1(new_n295), .A2(new_n284), .A3(new_n293), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n304), .A2(new_n305), .ZN(new_n306));
  NAND4_X1  g120(.A1(new_n306), .A2(KEYINPUT88), .A3(new_n187), .A4(new_n283), .ZN(new_n307));
  NAND3_X1  g121(.A1(new_n299), .A2(new_n302), .A3(new_n307), .ZN(new_n308));
  XOR2_X1   g122(.A(KEYINPUT89), .B(KEYINPUT20), .Z(new_n309));
  XNOR2_X1  g123(.A(G113), .B(G122), .ZN(new_n310));
  XNOR2_X1  g124(.A(new_n310), .B(new_n202), .ZN(new_n311));
  INV_X1    g125(.A(G237), .ZN(new_n312));
  NAND3_X1  g126(.A1(new_n312), .A2(new_n272), .A3(G214), .ZN(new_n313));
  XNOR2_X1  g127(.A(new_n313), .B(G143), .ZN(new_n314));
  INV_X1    g128(.A(KEYINPUT18), .ZN(new_n315));
  INV_X1    g129(.A(G131), .ZN(new_n316));
  OAI21_X1  g130(.A(new_n314), .B1(new_n315), .B2(new_n316), .ZN(new_n317));
  XNOR2_X1  g131(.A(new_n313), .B(new_n252), .ZN(new_n318));
  NAND3_X1  g132(.A1(new_n318), .A2(KEYINPUT18), .A3(G131), .ZN(new_n319));
  XNOR2_X1  g133(.A(G125), .B(G140), .ZN(new_n320));
  XNOR2_X1  g134(.A(new_n320), .B(new_n255), .ZN(new_n321));
  NAND3_X1  g135(.A1(new_n317), .A2(new_n319), .A3(new_n321), .ZN(new_n322));
  INV_X1    g136(.A(KEYINPUT75), .ZN(new_n323));
  INV_X1    g137(.A(G140), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n324), .A2(G125), .ZN(new_n325));
  INV_X1    g139(.A(G125), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n326), .A2(G140), .ZN(new_n327));
  NAND3_X1  g141(.A1(new_n325), .A2(new_n327), .A3(KEYINPUT16), .ZN(new_n328));
  OR3_X1    g142(.A1(new_n326), .A2(KEYINPUT16), .A3(G140), .ZN(new_n329));
  AOI21_X1  g143(.A(new_n323), .B1(new_n328), .B2(new_n329), .ZN(new_n330));
  NOR3_X1   g144(.A1(new_n326), .A2(KEYINPUT16), .A3(G140), .ZN(new_n331));
  NOR2_X1   g145(.A1(new_n331), .A2(KEYINPUT75), .ZN(new_n332));
  OAI21_X1  g146(.A(new_n255), .B1(new_n330), .B2(new_n332), .ZN(new_n333));
  INV_X1    g147(.A(new_n332), .ZN(new_n334));
  AOI21_X1  g148(.A(new_n331), .B1(new_n320), .B2(KEYINPUT16), .ZN(new_n335));
  OAI211_X1 g149(.A(new_n334), .B(G146), .C1(new_n335), .C2(new_n323), .ZN(new_n336));
  NAND3_X1  g150(.A1(new_n318), .A2(KEYINPUT17), .A3(G131), .ZN(new_n337));
  NAND3_X1  g151(.A1(new_n333), .A2(new_n336), .A3(new_n337), .ZN(new_n338));
  INV_X1    g152(.A(KEYINPUT91), .ZN(new_n339));
  AND2_X1   g153(.A1(new_n338), .A2(new_n339), .ZN(new_n340));
  NAND4_X1  g154(.A1(new_n333), .A2(new_n336), .A3(new_n337), .A4(KEYINPUT91), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n318), .A2(G131), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n314), .A2(new_n316), .ZN(new_n343));
  INV_X1    g157(.A(KEYINPUT17), .ZN(new_n344));
  NAND3_X1  g158(.A1(new_n342), .A2(new_n343), .A3(new_n344), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n341), .A2(new_n345), .ZN(new_n346));
  OAI211_X1 g160(.A(new_n311), .B(new_n322), .C1(new_n340), .C2(new_n346), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n342), .A2(new_n343), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n320), .A2(KEYINPUT90), .ZN(new_n349));
  XNOR2_X1  g163(.A(new_n349), .B(KEYINPUT19), .ZN(new_n350));
  OAI211_X1 g164(.A(new_n348), .B(new_n336), .C1(G146), .C2(new_n350), .ZN(new_n351));
  NAND2_X1  g165(.A1(new_n351), .A2(new_n322), .ZN(new_n352));
  INV_X1    g166(.A(new_n311), .ZN(new_n353));
  NAND2_X1  g167(.A1(new_n352), .A2(new_n353), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n347), .A2(new_n354), .ZN(new_n355));
  NOR2_X1   g169(.A1(G475), .A2(G902), .ZN(new_n356));
  AOI21_X1  g170(.A(new_n309), .B1(new_n355), .B2(new_n356), .ZN(new_n357));
  INV_X1    g171(.A(new_n356), .ZN(new_n358));
  AOI211_X1 g172(.A(KEYINPUT20), .B(new_n358), .C1(new_n347), .C2(new_n354), .ZN(new_n359));
  OAI21_X1  g173(.A(new_n322), .B1(new_n340), .B2(new_n346), .ZN(new_n360));
  NAND2_X1  g174(.A1(new_n360), .A2(new_n353), .ZN(new_n361));
  AOI21_X1  g175(.A(G902), .B1(new_n361), .B2(new_n347), .ZN(new_n362));
  INV_X1    g176(.A(G475), .ZN(new_n363));
  OAI22_X1  g177(.A1(new_n357), .A2(new_n359), .B1(new_n362), .B2(new_n363), .ZN(new_n364));
  INV_X1    g178(.A(new_n364), .ZN(new_n365));
  INV_X1    g179(.A(G134), .ZN(new_n366));
  NOR2_X1   g180(.A1(new_n265), .A2(G143), .ZN(new_n367));
  INV_X1    g181(.A(KEYINPUT13), .ZN(new_n368));
  AOI21_X1  g182(.A(new_n366), .B1(new_n367), .B2(new_n368), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n252), .A2(G128), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n265), .A2(G143), .ZN(new_n371));
  NAND3_X1  g185(.A1(new_n370), .A2(new_n371), .A3(KEYINPUT13), .ZN(new_n372));
  NAND3_X1  g186(.A1(new_n370), .A2(new_n371), .A3(new_n366), .ZN(new_n373));
  AOI22_X1  g187(.A1(new_n369), .A2(new_n372), .B1(new_n373), .B2(KEYINPUT93), .ZN(new_n374));
  OR2_X1    g188(.A1(new_n373), .A2(KEYINPUT93), .ZN(new_n375));
  OAI21_X1  g189(.A(KEYINPUT92), .B1(new_n190), .B2(G122), .ZN(new_n376));
  INV_X1    g190(.A(KEYINPUT92), .ZN(new_n377));
  INV_X1    g191(.A(G122), .ZN(new_n378));
  NAND3_X1  g192(.A1(new_n377), .A2(new_n378), .A3(G116), .ZN(new_n379));
  NAND2_X1  g193(.A1(new_n376), .A2(new_n379), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n190), .A2(G122), .ZN(new_n381));
  AND3_X1   g195(.A1(new_n380), .A2(new_n205), .A3(new_n381), .ZN(new_n382));
  AOI21_X1  g196(.A(new_n205), .B1(new_n380), .B2(new_n381), .ZN(new_n383));
  OAI211_X1 g197(.A(new_n374), .B(new_n375), .C1(new_n382), .C2(new_n383), .ZN(new_n384));
  AND2_X1   g198(.A1(new_n376), .A2(new_n379), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n381), .A2(KEYINPUT14), .ZN(new_n386));
  INV_X1    g200(.A(KEYINPUT14), .ZN(new_n387));
  NAND3_X1  g201(.A1(new_n387), .A2(new_n190), .A3(G122), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n386), .A2(new_n388), .ZN(new_n389));
  OAI21_X1  g203(.A(G107), .B1(new_n385), .B2(new_n389), .ZN(new_n390));
  NAND3_X1  g204(.A1(new_n380), .A2(new_n205), .A3(new_n381), .ZN(new_n391));
  INV_X1    g205(.A(new_n371), .ZN(new_n392));
  OAI21_X1  g206(.A(G134), .B1(new_n392), .B2(new_n367), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n393), .A2(new_n373), .ZN(new_n394));
  NAND3_X1  g208(.A1(new_n390), .A2(new_n391), .A3(new_n394), .ZN(new_n395));
  XNOR2_X1  g209(.A(KEYINPUT9), .B(G234), .ZN(new_n396));
  INV_X1    g210(.A(G217), .ZN(new_n397));
  NOR3_X1   g211(.A1(new_n396), .A2(new_n397), .A3(G953), .ZN(new_n398));
  NAND3_X1  g212(.A1(new_n384), .A2(new_n395), .A3(new_n398), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n399), .A2(KEYINPUT94), .ZN(new_n400));
  INV_X1    g214(.A(KEYINPUT94), .ZN(new_n401));
  NAND4_X1  g215(.A1(new_n384), .A2(new_n395), .A3(new_n401), .A4(new_n398), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n384), .A2(new_n395), .ZN(new_n403));
  INV_X1    g217(.A(new_n398), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n403), .A2(new_n404), .ZN(new_n405));
  NAND3_X1  g219(.A1(new_n400), .A2(new_n402), .A3(new_n405), .ZN(new_n406));
  INV_X1    g220(.A(G902), .ZN(new_n407));
  NAND2_X1  g221(.A1(new_n406), .A2(new_n407), .ZN(new_n408));
  NAND2_X1  g222(.A1(new_n408), .A2(KEYINPUT95), .ZN(new_n409));
  INV_X1    g223(.A(G478), .ZN(new_n410));
  NOR2_X1   g224(.A1(new_n410), .A2(KEYINPUT15), .ZN(new_n411));
  INV_X1    g225(.A(KEYINPUT95), .ZN(new_n412));
  NAND3_X1  g226(.A1(new_n406), .A2(new_n412), .A3(new_n407), .ZN(new_n413));
  NAND3_X1  g227(.A1(new_n409), .A2(new_n411), .A3(new_n413), .ZN(new_n414));
  OR2_X1    g228(.A1(new_n408), .A2(new_n411), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n414), .A2(new_n415), .ZN(new_n416));
  INV_X1    g230(.A(new_n416), .ZN(new_n417));
  NAND2_X1  g231(.A1(G234), .A2(G237), .ZN(new_n418));
  NAND3_X1  g232(.A1(new_n418), .A2(G952), .A3(new_n272), .ZN(new_n419));
  XNOR2_X1  g233(.A(KEYINPUT21), .B(G898), .ZN(new_n420));
  INV_X1    g234(.A(new_n420), .ZN(new_n421));
  NAND3_X1  g235(.A1(new_n418), .A2(G902), .A3(G953), .ZN(new_n422));
  OAI21_X1  g236(.A(new_n419), .B1(new_n421), .B2(new_n422), .ZN(new_n423));
  NAND4_X1  g237(.A1(new_n365), .A2(KEYINPUT96), .A3(new_n417), .A4(new_n423), .ZN(new_n424));
  INV_X1    g238(.A(KEYINPUT96), .ZN(new_n425));
  NAND3_X1  g239(.A1(new_n414), .A2(new_n415), .A3(new_n423), .ZN(new_n426));
  OAI21_X1  g240(.A(new_n425), .B1(new_n364), .B2(new_n426), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n424), .A2(new_n427), .ZN(new_n428));
  OAI21_X1  g242(.A(G214), .B1(G237), .B2(G902), .ZN(new_n429));
  INV_X1    g243(.A(G469), .ZN(new_n430));
  NAND3_X1  g244(.A1(new_n224), .A2(new_n261), .A3(new_n227), .ZN(new_n431));
  INV_X1    g245(.A(KEYINPUT10), .ZN(new_n432));
  AND2_X1   g246(.A1(new_n259), .A2(new_n266), .ZN(new_n433));
  INV_X1    g247(.A(KEYINPUT79), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n263), .A2(new_n434), .ZN(new_n435));
  OAI211_X1 g249(.A(KEYINPUT79), .B(KEYINPUT1), .C1(new_n252), .C2(G146), .ZN(new_n436));
  NAND3_X1  g250(.A1(new_n435), .A2(G128), .A3(new_n436), .ZN(new_n437));
  INV_X1    g251(.A(new_n259), .ZN(new_n438));
  AOI21_X1  g252(.A(new_n433), .B1(new_n437), .B2(new_n438), .ZN(new_n439));
  OAI21_X1  g253(.A(new_n432), .B1(new_n439), .B2(new_n277), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n258), .A2(new_n264), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n259), .A2(new_n266), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n441), .A2(new_n442), .ZN(new_n443));
  OAI211_X1 g257(.A(KEYINPUT10), .B(new_n443), .C1(new_n214), .C2(new_n215), .ZN(new_n444));
  INV_X1    g258(.A(KEYINPUT11), .ZN(new_n445));
  OAI21_X1  g259(.A(new_n445), .B1(new_n366), .B2(G137), .ZN(new_n446));
  INV_X1    g260(.A(G137), .ZN(new_n447));
  NAND3_X1  g261(.A1(new_n447), .A2(KEYINPUT11), .A3(G134), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n366), .A2(G137), .ZN(new_n449));
  NAND3_X1  g263(.A1(new_n446), .A2(new_n448), .A3(new_n449), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n450), .A2(G131), .ZN(new_n451));
  INV_X1    g265(.A(KEYINPUT81), .ZN(new_n452));
  NAND4_X1  g266(.A1(new_n446), .A2(new_n448), .A3(new_n316), .A4(new_n449), .ZN(new_n453));
  AND3_X1   g267(.A1(new_n451), .A2(new_n452), .A3(new_n453), .ZN(new_n454));
  AOI21_X1  g268(.A(new_n452), .B1(new_n451), .B2(new_n453), .ZN(new_n455));
  NOR2_X1   g269(.A1(new_n454), .A2(new_n455), .ZN(new_n456));
  NAND4_X1  g270(.A1(new_n431), .A2(new_n440), .A3(new_n444), .A4(new_n456), .ZN(new_n457));
  XNOR2_X1  g271(.A(G110), .B(G140), .ZN(new_n458));
  AND2_X1   g272(.A1(new_n272), .A2(G227), .ZN(new_n459));
  XNOR2_X1  g273(.A(new_n458), .B(new_n459), .ZN(new_n460));
  INV_X1    g274(.A(new_n460), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n267), .A2(new_n277), .ZN(new_n462));
  OAI21_X1  g276(.A(new_n462), .B1(new_n439), .B2(new_n277), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n451), .A2(new_n453), .ZN(new_n464));
  AND3_X1   g278(.A1(new_n463), .A2(KEYINPUT12), .A3(new_n464), .ZN(new_n465));
  AOI21_X1  g279(.A(KEYINPUT12), .B1(new_n463), .B2(new_n464), .ZN(new_n466));
  OAI211_X1 g280(.A(new_n457), .B(new_n461), .C1(new_n465), .C2(new_n466), .ZN(new_n467));
  INV_X1    g281(.A(new_n467), .ZN(new_n468));
  NAND3_X1  g282(.A1(new_n431), .A2(new_n440), .A3(new_n444), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n469), .A2(new_n464), .ZN(new_n470));
  AOI21_X1  g284(.A(new_n461), .B1(new_n470), .B2(new_n457), .ZN(new_n471));
  OAI211_X1 g285(.A(new_n430), .B(new_n407), .C1(new_n468), .C2(new_n471), .ZN(new_n472));
  NAND2_X1  g286(.A1(G469), .A2(G902), .ZN(new_n473));
  OAI21_X1  g287(.A(new_n457), .B1(new_n465), .B2(new_n466), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n474), .A2(new_n460), .ZN(new_n475));
  NAND3_X1  g289(.A1(new_n470), .A2(new_n457), .A3(new_n461), .ZN(new_n476));
  NAND3_X1  g290(.A1(new_n475), .A2(G469), .A3(new_n476), .ZN(new_n477));
  NAND3_X1  g291(.A1(new_n472), .A2(new_n473), .A3(new_n477), .ZN(new_n478));
  OAI21_X1  g292(.A(G221), .B1(new_n396), .B2(G902), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n478), .A2(new_n479), .ZN(new_n480));
  INV_X1    g294(.A(new_n480), .ZN(new_n481));
  NAND4_X1  g295(.A1(new_n308), .A2(new_n428), .A3(new_n429), .A4(new_n481), .ZN(new_n482));
  INV_X1    g296(.A(KEYINPUT72), .ZN(new_n483));
  INV_X1    g297(.A(KEYINPUT67), .ZN(new_n484));
  INV_X1    g298(.A(KEYINPUT66), .ZN(new_n485));
  NOR2_X1   g299(.A1(new_n366), .A2(G137), .ZN(new_n486));
  NOR2_X1   g300(.A1(new_n447), .A2(G134), .ZN(new_n487));
  OAI21_X1  g301(.A(G131), .B1(new_n486), .B2(new_n487), .ZN(new_n488));
  AOI21_X1  g302(.A(new_n485), .B1(new_n453), .B2(new_n488), .ZN(new_n489));
  NOR2_X1   g303(.A1(new_n489), .A2(new_n267), .ZN(new_n490));
  AND3_X1   g304(.A1(new_n453), .A2(new_n488), .A3(new_n485), .ZN(new_n491));
  INV_X1    g305(.A(new_n491), .ZN(new_n492));
  AOI22_X1  g306(.A1(new_n490), .A2(new_n492), .B1(new_n261), .B2(new_n464), .ZN(new_n493));
  OAI21_X1  g307(.A(new_n484), .B1(new_n493), .B2(KEYINPUT30), .ZN(new_n494));
  INV_X1    g308(.A(KEYINPUT30), .ZN(new_n495));
  NOR3_X1   g309(.A1(new_n491), .A2(new_n489), .A3(new_n267), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n464), .A2(new_n261), .ZN(new_n497));
  INV_X1    g311(.A(new_n497), .ZN(new_n498));
  OAI211_X1 g312(.A(KEYINPUT67), .B(new_n495), .C1(new_n496), .C2(new_n498), .ZN(new_n499));
  INV_X1    g313(.A(KEYINPUT69), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n497), .A2(new_n500), .ZN(new_n501));
  NAND3_X1  g315(.A1(new_n464), .A2(new_n261), .A3(KEYINPUT69), .ZN(new_n502));
  AND2_X1   g316(.A1(new_n453), .A2(new_n488), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n443), .A2(new_n503), .ZN(new_n504));
  NAND4_X1  g318(.A1(new_n501), .A2(KEYINPUT30), .A3(new_n502), .A4(new_n504), .ZN(new_n505));
  NAND4_X1  g319(.A1(new_n494), .A2(new_n499), .A3(new_n242), .A4(new_n505), .ZN(new_n506));
  NOR2_X1   g320(.A1(new_n234), .A2(new_n235), .ZN(new_n507));
  NAND4_X1  g321(.A1(new_n501), .A2(new_n507), .A3(new_n502), .A4(new_n504), .ZN(new_n508));
  NAND3_X1  g322(.A1(new_n312), .A2(new_n272), .A3(G210), .ZN(new_n509));
  XOR2_X1   g323(.A(new_n509), .B(KEYINPUT27), .Z(new_n510));
  XNOR2_X1  g324(.A(KEYINPUT26), .B(G101), .ZN(new_n511));
  XNOR2_X1  g325(.A(new_n510), .B(new_n511), .ZN(new_n512));
  INV_X1    g326(.A(KEYINPUT70), .ZN(new_n513));
  NOR2_X1   g327(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  NAND3_X1  g328(.A1(new_n506), .A2(new_n508), .A3(new_n514), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n515), .A2(KEYINPUT31), .ZN(new_n516));
  OAI21_X1  g330(.A(new_n508), .B1(new_n507), .B2(new_n493), .ZN(new_n517));
  AND2_X1   g331(.A1(new_n517), .A2(KEYINPUT28), .ZN(new_n518));
  NAND3_X1  g332(.A1(new_n507), .A2(new_n497), .A3(new_n504), .ZN(new_n519));
  INV_X1    g333(.A(KEYINPUT28), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  INV_X1    g335(.A(new_n521), .ZN(new_n522));
  OAI21_X1  g336(.A(new_n512), .B1(new_n518), .B2(new_n522), .ZN(new_n523));
  NOR3_X1   g337(.A1(new_n512), .A2(new_n513), .A3(KEYINPUT31), .ZN(new_n524));
  NAND3_X1  g338(.A1(new_n506), .A2(new_n508), .A3(new_n524), .ZN(new_n525));
  NAND3_X1  g339(.A1(new_n516), .A2(new_n523), .A3(new_n525), .ZN(new_n526));
  NOR2_X1   g340(.A1(G472), .A2(G902), .ZN(new_n527));
  INV_X1    g341(.A(new_n527), .ZN(new_n528));
  INV_X1    g342(.A(KEYINPUT32), .ZN(new_n529));
  NOR2_X1   g343(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n526), .A2(new_n530), .ZN(new_n531));
  INV_X1    g345(.A(KEYINPUT29), .ZN(new_n532));
  NAND4_X1  g346(.A1(new_n506), .A2(new_n532), .A3(new_n508), .A4(new_n512), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n533), .A2(new_n407), .ZN(new_n534));
  NAND2_X1  g348(.A1(new_n502), .A2(new_n504), .ZN(new_n535));
  AOI21_X1  g349(.A(KEYINPUT69), .B1(new_n464), .B2(new_n261), .ZN(new_n536));
  OAI21_X1  g350(.A(new_n242), .B1(new_n535), .B2(new_n536), .ZN(new_n537));
  OAI21_X1  g351(.A(new_n537), .B1(new_n508), .B2(KEYINPUT71), .ZN(new_n538));
  INV_X1    g352(.A(KEYINPUT71), .ZN(new_n539));
  NOR2_X1   g353(.A1(new_n535), .A2(new_n536), .ZN(new_n540));
  AOI21_X1  g354(.A(new_n539), .B1(new_n540), .B2(new_n507), .ZN(new_n541));
  OAI21_X1  g355(.A(KEYINPUT28), .B1(new_n538), .B2(new_n541), .ZN(new_n542));
  NAND2_X1  g356(.A1(new_n542), .A2(new_n521), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n543), .A2(KEYINPUT29), .ZN(new_n544));
  AOI21_X1  g358(.A(new_n522), .B1(new_n517), .B2(KEYINPUT28), .ZN(new_n545));
  AOI21_X1  g359(.A(new_n512), .B1(new_n545), .B2(new_n532), .ZN(new_n546));
  AOI21_X1  g360(.A(new_n534), .B1(new_n544), .B2(new_n546), .ZN(new_n547));
  INV_X1    g361(.A(G472), .ZN(new_n548));
  OAI21_X1  g362(.A(new_n531), .B1(new_n547), .B2(new_n548), .ZN(new_n549));
  AOI21_X1  g363(.A(KEYINPUT32), .B1(new_n526), .B2(new_n527), .ZN(new_n550));
  OAI21_X1  g364(.A(new_n483), .B1(new_n549), .B2(new_n550), .ZN(new_n551));
  XNOR2_X1  g365(.A(KEYINPUT22), .B(G137), .ZN(new_n552));
  NAND3_X1  g366(.A1(new_n272), .A2(G221), .A3(G234), .ZN(new_n553));
  XNOR2_X1  g367(.A(new_n552), .B(new_n553), .ZN(new_n554));
  INV_X1    g368(.A(new_n554), .ZN(new_n555));
  XNOR2_X1  g369(.A(KEYINPUT24), .B(G110), .ZN(new_n556));
  INV_X1    g370(.A(KEYINPUT73), .ZN(new_n557));
  XNOR2_X1  g371(.A(new_n556), .B(new_n557), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n188), .A2(G128), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n265), .A2(G119), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n559), .A2(new_n560), .ZN(new_n561));
  INV_X1    g375(.A(new_n561), .ZN(new_n562));
  INV_X1    g376(.A(KEYINPUT74), .ZN(new_n563));
  OAI21_X1  g377(.A(new_n563), .B1(new_n188), .B2(G128), .ZN(new_n564));
  NAND3_X1  g378(.A1(new_n564), .A2(KEYINPUT23), .A3(new_n559), .ZN(new_n565));
  OAI21_X1  g379(.A(KEYINPUT23), .B1(new_n265), .B2(G119), .ZN(new_n566));
  NAND3_X1  g380(.A1(new_n566), .A2(new_n563), .A3(new_n560), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n565), .A2(new_n567), .ZN(new_n568));
  OAI22_X1  g382(.A1(new_n558), .A2(new_n562), .B1(G110), .B2(new_n568), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n320), .A2(new_n255), .ZN(new_n570));
  AND3_X1   g384(.A1(new_n569), .A2(new_n336), .A3(new_n570), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n568), .A2(G110), .ZN(new_n572));
  XNOR2_X1  g386(.A(new_n556), .B(KEYINPUT73), .ZN(new_n573));
  OAI21_X1  g387(.A(new_n572), .B1(new_n573), .B2(new_n561), .ZN(new_n574));
  AOI21_X1  g388(.A(new_n574), .B1(new_n336), .B2(new_n333), .ZN(new_n575));
  OAI21_X1  g389(.A(new_n555), .B1(new_n571), .B2(new_n575), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n333), .A2(new_n336), .ZN(new_n577));
  OAI211_X1 g391(.A(new_n577), .B(new_n572), .C1(new_n561), .C2(new_n573), .ZN(new_n578));
  NAND3_X1  g392(.A1(new_n569), .A2(new_n336), .A3(new_n570), .ZN(new_n579));
  NAND3_X1  g393(.A1(new_n578), .A2(new_n579), .A3(new_n554), .ZN(new_n580));
  AND2_X1   g394(.A1(new_n576), .A2(new_n580), .ZN(new_n581));
  AOI21_X1  g395(.A(new_n397), .B1(G234), .B2(new_n407), .ZN(new_n582));
  NOR2_X1   g396(.A1(new_n582), .A2(G902), .ZN(new_n583));
  XNOR2_X1  g397(.A(new_n583), .B(KEYINPUT77), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n581), .A2(new_n584), .ZN(new_n585));
  INV_X1    g399(.A(new_n585), .ZN(new_n586));
  NAND3_X1  g400(.A1(new_n576), .A2(new_n407), .A3(new_n580), .ZN(new_n587));
  INV_X1    g401(.A(KEYINPUT76), .ZN(new_n588));
  AOI21_X1  g402(.A(KEYINPUT25), .B1(new_n587), .B2(new_n588), .ZN(new_n589));
  INV_X1    g403(.A(new_n582), .ZN(new_n590));
  NOR2_X1   g404(.A1(new_n589), .A2(new_n590), .ZN(new_n591));
  NAND3_X1  g405(.A1(new_n587), .A2(new_n588), .A3(KEYINPUT25), .ZN(new_n592));
  AOI21_X1  g406(.A(new_n586), .B1(new_n591), .B2(new_n592), .ZN(new_n593));
  NAND2_X1  g407(.A1(new_n526), .A2(new_n527), .ZN(new_n594));
  NAND2_X1  g408(.A1(new_n594), .A2(new_n529), .ZN(new_n595));
  NAND3_X1  g409(.A1(new_n540), .A2(new_n539), .A3(new_n507), .ZN(new_n596));
  NAND2_X1  g410(.A1(new_n508), .A2(KEYINPUT71), .ZN(new_n597));
  NAND3_X1  g411(.A1(new_n596), .A2(new_n597), .A3(new_n537), .ZN(new_n598));
  AOI21_X1  g412(.A(new_n522), .B1(new_n598), .B2(KEYINPUT28), .ZN(new_n599));
  OAI21_X1  g413(.A(new_n546), .B1(new_n599), .B2(new_n532), .ZN(new_n600));
  INV_X1    g414(.A(new_n534), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n602), .A2(G472), .ZN(new_n603));
  NAND4_X1  g417(.A1(new_n595), .A2(new_n603), .A3(KEYINPUT72), .A4(new_n531), .ZN(new_n604));
  NAND3_X1  g418(.A1(new_n551), .A2(new_n593), .A3(new_n604), .ZN(new_n605));
  NOR2_X1   g419(.A1(new_n482), .A2(new_n605), .ZN(new_n606));
  XNOR2_X1  g420(.A(new_n606), .B(new_n207), .ZN(G3));
  INV_X1    g421(.A(new_n429), .ZN(new_n608));
  AOI21_X1  g422(.A(new_n187), .B1(new_n306), .B2(new_n283), .ZN(new_n609));
  AOI21_X1  g423(.A(new_n608), .B1(new_n609), .B2(KEYINPUT97), .ZN(new_n610));
  NAND3_X1  g424(.A1(new_n409), .A2(new_n410), .A3(new_n413), .ZN(new_n611));
  NOR2_X1   g425(.A1(new_n410), .A2(G902), .ZN(new_n612));
  INV_X1    g426(.A(KEYINPUT33), .ZN(new_n613));
  NOR2_X1   g427(.A1(new_n399), .A2(KEYINPUT98), .ZN(new_n614));
  AOI21_X1  g428(.A(new_n398), .B1(new_n384), .B2(new_n395), .ZN(new_n615));
  NOR2_X1   g429(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  NAND2_X1  g430(.A1(new_n399), .A2(KEYINPUT98), .ZN(new_n617));
  AOI21_X1  g431(.A(new_n613), .B1(new_n616), .B2(new_n617), .ZN(new_n618));
  NOR2_X1   g432(.A1(new_n406), .A2(KEYINPUT33), .ZN(new_n619));
  OAI21_X1  g433(.A(new_n612), .B1(new_n618), .B2(new_n619), .ZN(new_n620));
  NAND2_X1  g434(.A1(new_n611), .A2(new_n620), .ZN(new_n621));
  NAND2_X1  g435(.A1(new_n364), .A2(new_n621), .ZN(new_n622));
  XNOR2_X1  g436(.A(new_n622), .B(KEYINPUT99), .ZN(new_n623));
  INV_X1    g437(.A(new_n187), .ZN(new_n624));
  NAND2_X1  g438(.A1(new_n300), .A2(new_n624), .ZN(new_n625));
  INV_X1    g439(.A(KEYINPUT97), .ZN(new_n626));
  NAND3_X1  g440(.A1(new_n625), .A2(new_n626), .A3(new_n297), .ZN(new_n627));
  NAND4_X1  g441(.A1(new_n610), .A2(new_n623), .A3(new_n627), .A4(new_n423), .ZN(new_n628));
  AOI21_X1  g442(.A(new_n548), .B1(new_n526), .B2(new_n407), .ZN(new_n629));
  INV_X1    g443(.A(new_n629), .ZN(new_n630));
  NAND2_X1  g444(.A1(new_n630), .A2(new_n594), .ZN(new_n631));
  NAND3_X1  g445(.A1(new_n593), .A2(new_n479), .A3(new_n478), .ZN(new_n632));
  NOR3_X1   g446(.A1(new_n628), .A2(new_n631), .A3(new_n632), .ZN(new_n633));
  XNOR2_X1  g447(.A(KEYINPUT34), .B(G104), .ZN(new_n634));
  XNOR2_X1  g448(.A(new_n633), .B(new_n634), .ZN(G6));
  INV_X1    g449(.A(new_n347), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n338), .A2(new_n339), .ZN(new_n637));
  NAND3_X1  g451(.A1(new_n637), .A2(new_n345), .A3(new_n341), .ZN(new_n638));
  AOI21_X1  g452(.A(new_n311), .B1(new_n638), .B2(new_n322), .ZN(new_n639));
  OAI21_X1  g453(.A(new_n407), .B1(new_n636), .B2(new_n639), .ZN(new_n640));
  NAND2_X1  g454(.A1(new_n640), .A2(G475), .ZN(new_n641));
  AOI21_X1  g455(.A(new_n358), .B1(new_n347), .B2(new_n354), .ZN(new_n642));
  AND2_X1   g456(.A1(new_n642), .A2(new_n309), .ZN(new_n643));
  OAI21_X1  g457(.A(new_n641), .B1(new_n643), .B2(new_n357), .ZN(new_n644));
  NOR2_X1   g458(.A1(new_n417), .A2(new_n644), .ZN(new_n645));
  NAND4_X1  g459(.A1(new_n610), .A2(new_n627), .A3(new_n423), .A4(new_n645), .ZN(new_n646));
  NOR3_X1   g460(.A1(new_n646), .A2(new_n631), .A3(new_n632), .ZN(new_n647));
  XNOR2_X1  g461(.A(KEYINPUT35), .B(G107), .ZN(new_n648));
  XNOR2_X1  g462(.A(new_n647), .B(new_n648), .ZN(G9));
  INV_X1    g463(.A(KEYINPUT100), .ZN(new_n650));
  AND3_X1   g464(.A1(new_n587), .A2(new_n588), .A3(KEYINPUT25), .ZN(new_n651));
  NOR3_X1   g465(.A1(new_n651), .A2(new_n589), .A3(new_n590), .ZN(new_n652));
  NAND2_X1  g466(.A1(new_n578), .A2(new_n579), .ZN(new_n653));
  NOR2_X1   g467(.A1(new_n555), .A2(KEYINPUT36), .ZN(new_n654));
  XNOR2_X1  g468(.A(new_n653), .B(new_n654), .ZN(new_n655));
  NAND2_X1  g469(.A1(new_n655), .A2(new_n584), .ZN(new_n656));
  INV_X1    g470(.A(new_n656), .ZN(new_n657));
  OAI21_X1  g471(.A(new_n650), .B1(new_n652), .B2(new_n657), .ZN(new_n658));
  NAND2_X1  g472(.A1(new_n587), .A2(new_n588), .ZN(new_n659));
  INV_X1    g473(.A(KEYINPUT25), .ZN(new_n660));
  NAND2_X1  g474(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  NAND3_X1  g475(.A1(new_n661), .A2(new_n582), .A3(new_n592), .ZN(new_n662));
  NAND3_X1  g476(.A1(new_n662), .A2(KEYINPUT100), .A3(new_n656), .ZN(new_n663));
  NAND3_X1  g477(.A1(new_n481), .A2(new_n658), .A3(new_n663), .ZN(new_n664));
  NOR2_X1   g478(.A1(new_n664), .A2(new_n631), .ZN(new_n665));
  NAND4_X1  g479(.A1(new_n665), .A2(new_n429), .A3(new_n308), .A4(new_n428), .ZN(new_n666));
  XOR2_X1   g480(.A(KEYINPUT37), .B(G110), .Z(new_n667));
  XNOR2_X1  g481(.A(new_n666), .B(new_n667), .ZN(G12));
  NAND2_X1  g482(.A1(new_n610), .A2(new_n627), .ZN(new_n669));
  XNOR2_X1  g483(.A(new_n419), .B(KEYINPUT101), .ZN(new_n670));
  OAI21_X1  g484(.A(new_n670), .B1(G900), .B2(new_n422), .ZN(new_n671));
  INV_X1    g485(.A(new_n671), .ZN(new_n672));
  OR2_X1    g486(.A1(new_n644), .A2(new_n672), .ZN(new_n673));
  NOR3_X1   g487(.A1(new_n669), .A2(new_n417), .A3(new_n673), .ZN(new_n674));
  NAND2_X1  g488(.A1(new_n551), .A2(new_n604), .ZN(new_n675));
  NOR2_X1   g489(.A1(new_n675), .A2(new_n664), .ZN(new_n676));
  NAND2_X1  g490(.A1(new_n674), .A2(new_n676), .ZN(new_n677));
  XNOR2_X1  g491(.A(new_n677), .B(G128), .ZN(G30));
  AND2_X1   g492(.A1(new_n506), .A2(new_n508), .ZN(new_n679));
  NOR2_X1   g493(.A1(new_n679), .A2(new_n512), .ZN(new_n680));
  INV_X1    g494(.A(new_n512), .ZN(new_n681));
  OAI21_X1  g495(.A(new_n407), .B1(new_n598), .B2(new_n681), .ZN(new_n682));
  OAI21_X1  g496(.A(G472), .B1(new_n680), .B2(new_n682), .ZN(new_n683));
  AND3_X1   g497(.A1(new_n595), .A2(new_n531), .A3(new_n683), .ZN(new_n684));
  NOR2_X1   g498(.A1(new_n652), .A2(new_n657), .ZN(new_n685));
  INV_X1    g499(.A(new_n685), .ZN(new_n686));
  NOR2_X1   g500(.A1(new_n686), .A2(new_n608), .ZN(new_n687));
  NOR2_X1   g501(.A1(new_n365), .A2(new_n417), .ZN(new_n688));
  XOR2_X1   g502(.A(new_n671), .B(KEYINPUT39), .Z(new_n689));
  NOR2_X1   g503(.A1(new_n480), .A2(new_n689), .ZN(new_n690));
  INV_X1    g504(.A(new_n690), .ZN(new_n691));
  OAI211_X1 g505(.A(new_n687), .B(new_n688), .C1(KEYINPUT40), .C2(new_n691), .ZN(new_n692));
  AOI211_X1 g506(.A(new_n684), .B(new_n692), .C1(KEYINPUT40), .C2(new_n691), .ZN(new_n693));
  XOR2_X1   g507(.A(new_n308), .B(KEYINPUT38), .Z(new_n694));
  INV_X1    g508(.A(new_n694), .ZN(new_n695));
  NAND2_X1  g509(.A1(new_n693), .A2(new_n695), .ZN(new_n696));
  XNOR2_X1  g510(.A(new_n696), .B(G143), .ZN(G45));
  NOR2_X1   g511(.A1(new_n622), .A2(new_n672), .ZN(new_n698));
  INV_X1    g512(.A(new_n698), .ZN(new_n699));
  OAI21_X1  g513(.A(KEYINPUT102), .B1(new_n669), .B2(new_n699), .ZN(new_n700));
  INV_X1    g514(.A(KEYINPUT102), .ZN(new_n701));
  NAND4_X1  g515(.A1(new_n610), .A2(new_n627), .A3(new_n701), .A4(new_n698), .ZN(new_n702));
  NAND3_X1  g516(.A1(new_n700), .A2(new_n676), .A3(new_n702), .ZN(new_n703));
  XNOR2_X1  g517(.A(new_n703), .B(G146), .ZN(G48));
  NOR2_X1   g518(.A1(new_n468), .A2(new_n471), .ZN(new_n705));
  OAI21_X1  g519(.A(G469), .B1(new_n705), .B2(G902), .ZN(new_n706));
  AND2_X1   g520(.A1(new_n706), .A2(new_n472), .ZN(new_n707));
  INV_X1    g521(.A(new_n707), .ZN(new_n708));
  INV_X1    g522(.A(new_n479), .ZN(new_n709));
  NOR2_X1   g523(.A1(new_n708), .A2(new_n709), .ZN(new_n710));
  NAND4_X1  g524(.A1(new_n551), .A2(new_n593), .A3(new_n604), .A4(new_n710), .ZN(new_n711));
  NOR2_X1   g525(.A1(new_n628), .A2(new_n711), .ZN(new_n712));
  XOR2_X1   g526(.A(KEYINPUT41), .B(G113), .Z(new_n713));
  XNOR2_X1  g527(.A(new_n712), .B(new_n713), .ZN(G15));
  NOR2_X1   g528(.A1(new_n711), .A2(new_n646), .ZN(new_n715));
  XNOR2_X1  g529(.A(KEYINPUT103), .B(G116), .ZN(new_n716));
  XNOR2_X1  g530(.A(new_n715), .B(new_n716), .ZN(G18));
  NAND2_X1  g531(.A1(new_n658), .A2(new_n663), .ZN(new_n718));
  AOI21_X1  g532(.A(new_n718), .B1(new_n427), .B2(new_n424), .ZN(new_n719));
  NAND4_X1  g533(.A1(new_n719), .A2(new_n627), .A3(new_n610), .A4(new_n710), .ZN(new_n720));
  NOR2_X1   g534(.A1(new_n720), .A2(new_n675), .ZN(new_n721));
  XNOR2_X1  g535(.A(new_n721), .B(new_n188), .ZN(G21));
  NAND4_X1  g536(.A1(new_n706), .A2(new_n423), .A3(new_n479), .A4(new_n472), .ZN(new_n723));
  AOI22_X1  g537(.A1(new_n679), .A2(new_n524), .B1(new_n515), .B2(KEYINPUT31), .ZN(new_n724));
  NAND2_X1  g538(.A1(new_n543), .A2(new_n512), .ZN(new_n725));
  AOI21_X1  g539(.A(new_n528), .B1(new_n724), .B2(new_n725), .ZN(new_n726));
  NAND2_X1  g540(.A1(new_n662), .A2(new_n585), .ZN(new_n727));
  NOR4_X1   g541(.A1(new_n629), .A2(new_n723), .A3(new_n726), .A4(new_n727), .ZN(new_n728));
  NAND4_X1  g542(.A1(new_n728), .A2(new_n627), .A3(new_n610), .A4(new_n688), .ZN(new_n729));
  XNOR2_X1  g543(.A(new_n729), .B(G122), .ZN(G24));
  INV_X1    g544(.A(new_n710), .ZN(new_n731));
  NOR2_X1   g545(.A1(new_n669), .A2(new_n731), .ZN(new_n732));
  NOR3_X1   g546(.A1(new_n685), .A2(new_n629), .A3(new_n726), .ZN(new_n733));
  AND2_X1   g547(.A1(new_n733), .A2(new_n698), .ZN(new_n734));
  NAND2_X1  g548(.A1(new_n732), .A2(new_n734), .ZN(new_n735));
  XNOR2_X1  g549(.A(new_n735), .B(G125), .ZN(G27));
  INV_X1    g550(.A(KEYINPUT106), .ZN(new_n737));
  AND2_X1   g551(.A1(new_n299), .A2(new_n307), .ZN(new_n738));
  AOI21_X1  g552(.A(new_n608), .B1(new_n300), .B2(new_n301), .ZN(new_n739));
  INV_X1    g553(.A(new_n464), .ZN(new_n740));
  AND2_X1   g554(.A1(new_n440), .A2(new_n444), .ZN(new_n741));
  AOI21_X1  g555(.A(new_n740), .B1(new_n741), .B2(new_n431), .ZN(new_n742));
  INV_X1    g556(.A(new_n457), .ZN(new_n743));
  OAI21_X1  g557(.A(new_n460), .B1(new_n742), .B2(new_n743), .ZN(new_n744));
  AOI211_X1 g558(.A(G469), .B(G902), .C1(new_n744), .C2(new_n467), .ZN(new_n745));
  NAND2_X1  g559(.A1(new_n477), .A2(new_n473), .ZN(new_n746));
  OAI21_X1  g560(.A(KEYINPUT104), .B1(new_n745), .B2(new_n746), .ZN(new_n747));
  INV_X1    g561(.A(KEYINPUT104), .ZN(new_n748));
  NAND4_X1  g562(.A1(new_n472), .A2(new_n748), .A3(new_n473), .A4(new_n477), .ZN(new_n749));
  AND3_X1   g563(.A1(new_n747), .A2(new_n479), .A3(new_n749), .ZN(new_n750));
  NAND4_X1  g564(.A1(new_n738), .A2(KEYINPUT105), .A3(new_n739), .A4(new_n750), .ZN(new_n751));
  NAND4_X1  g565(.A1(new_n750), .A2(new_n739), .A3(new_n299), .A4(new_n307), .ZN(new_n752));
  INV_X1    g566(.A(KEYINPUT105), .ZN(new_n753));
  NAND2_X1  g567(.A1(new_n752), .A2(new_n753), .ZN(new_n754));
  NAND2_X1  g568(.A1(new_n751), .A2(new_n754), .ZN(new_n755));
  INV_X1    g569(.A(KEYINPUT42), .ZN(new_n756));
  NOR3_X1   g570(.A1(new_n622), .A2(new_n756), .A3(new_n672), .ZN(new_n757));
  OAI211_X1 g571(.A(new_n757), .B(new_n593), .C1(new_n550), .C2(new_n549), .ZN(new_n758));
  INV_X1    g572(.A(new_n758), .ZN(new_n759));
  AOI21_X1  g573(.A(new_n737), .B1(new_n755), .B2(new_n759), .ZN(new_n760));
  AOI211_X1 g574(.A(KEYINPUT106), .B(new_n758), .C1(new_n751), .C2(new_n754), .ZN(new_n761));
  AOI211_X1 g575(.A(new_n699), .B(new_n605), .C1(new_n751), .C2(new_n754), .ZN(new_n762));
  OAI22_X1  g576(.A1(new_n760), .A2(new_n761), .B1(new_n762), .B2(KEYINPUT42), .ZN(new_n763));
  XNOR2_X1  g577(.A(new_n763), .B(G131), .ZN(G33));
  INV_X1    g578(.A(new_n605), .ZN(new_n765));
  NOR2_X1   g579(.A1(new_n673), .A2(new_n417), .ZN(new_n766));
  NAND3_X1  g580(.A1(new_n755), .A2(new_n765), .A3(new_n766), .ZN(new_n767));
  XNOR2_X1  g581(.A(new_n767), .B(G134), .ZN(G36));
  INV_X1    g582(.A(KEYINPUT20), .ZN(new_n769));
  NAND3_X1  g583(.A1(new_n355), .A2(new_n769), .A3(new_n356), .ZN(new_n770));
  OAI21_X1  g584(.A(new_n770), .B1(new_n309), .B2(new_n642), .ZN(new_n771));
  AND3_X1   g585(.A1(new_n621), .A2(new_n771), .A3(new_n641), .ZN(new_n772));
  XNOR2_X1  g586(.A(new_n772), .B(KEYINPUT43), .ZN(new_n773));
  NAND3_X1  g587(.A1(new_n773), .A2(new_n631), .A3(new_n686), .ZN(new_n774));
  INV_X1    g588(.A(KEYINPUT44), .ZN(new_n775));
  NAND2_X1  g589(.A1(new_n774), .A2(new_n775), .ZN(new_n776));
  XOR2_X1   g590(.A(new_n776), .B(KEYINPUT108), .Z(new_n777));
  AND2_X1   g591(.A1(new_n475), .A2(new_n476), .ZN(new_n778));
  OR2_X1    g592(.A1(new_n778), .A2(KEYINPUT45), .ZN(new_n779));
  NAND2_X1  g593(.A1(new_n778), .A2(KEYINPUT45), .ZN(new_n780));
  NAND3_X1  g594(.A1(new_n779), .A2(G469), .A3(new_n780), .ZN(new_n781));
  AND2_X1   g595(.A1(new_n781), .A2(new_n473), .ZN(new_n782));
  AND2_X1   g596(.A1(new_n782), .A2(KEYINPUT46), .ZN(new_n783));
  OAI21_X1  g597(.A(new_n472), .B1(new_n782), .B2(KEYINPUT46), .ZN(new_n784));
  OAI21_X1  g598(.A(new_n479), .B1(new_n783), .B2(new_n784), .ZN(new_n785));
  NOR2_X1   g599(.A1(new_n785), .A2(new_n689), .ZN(new_n786));
  NAND2_X1  g600(.A1(new_n738), .A2(new_n739), .ZN(new_n787));
  INV_X1    g601(.A(new_n787), .ZN(new_n788));
  OAI21_X1  g602(.A(new_n788), .B1(new_n774), .B2(new_n775), .ZN(new_n789));
  OR2_X1    g603(.A1(new_n789), .A2(KEYINPUT107), .ZN(new_n790));
  NAND2_X1  g604(.A1(new_n789), .A2(KEYINPUT107), .ZN(new_n791));
  NAND4_X1  g605(.A1(new_n777), .A2(new_n786), .A3(new_n790), .A4(new_n791), .ZN(new_n792));
  XNOR2_X1  g606(.A(new_n792), .B(G137), .ZN(G39));
  INV_X1    g607(.A(new_n675), .ZN(new_n794));
  NOR4_X1   g608(.A1(new_n794), .A2(new_n787), .A3(new_n593), .A4(new_n699), .ZN(new_n795));
  AND2_X1   g609(.A1(new_n795), .A2(KEYINPUT109), .ZN(new_n796));
  XNOR2_X1  g610(.A(new_n785), .B(KEYINPUT47), .ZN(new_n797));
  NOR2_X1   g611(.A1(new_n796), .A2(new_n797), .ZN(new_n798));
  OAI21_X1  g612(.A(new_n798), .B1(KEYINPUT109), .B2(new_n795), .ZN(new_n799));
  XNOR2_X1  g613(.A(KEYINPUT110), .B(G140), .ZN(new_n800));
  XNOR2_X1  g614(.A(new_n799), .B(new_n800), .ZN(G42));
  INV_X1    g615(.A(new_n670), .ZN(new_n802));
  NAND2_X1  g616(.A1(new_n773), .A2(new_n802), .ZN(new_n803));
  NOR4_X1   g617(.A1(new_n803), .A2(new_n727), .A3(new_n629), .A4(new_n726), .ZN(new_n804));
  NOR2_X1   g618(.A1(new_n731), .A2(new_n429), .ZN(new_n805));
  NAND3_X1  g619(.A1(new_n804), .A2(new_n694), .A3(new_n805), .ZN(new_n806));
  INV_X1    g620(.A(KEYINPUT50), .ZN(new_n807));
  XNOR2_X1  g621(.A(new_n806), .B(new_n807), .ZN(new_n808));
  NAND2_X1  g622(.A1(new_n788), .A2(new_n710), .ZN(new_n809));
  NAND2_X1  g623(.A1(new_n684), .A2(new_n593), .ZN(new_n810));
  NOR3_X1   g624(.A1(new_n809), .A2(new_n419), .A3(new_n810), .ZN(new_n811));
  NOR2_X1   g625(.A1(new_n364), .A2(new_n621), .ZN(new_n812));
  NOR2_X1   g626(.A1(new_n809), .A2(new_n803), .ZN(new_n813));
  AOI22_X1  g627(.A1(new_n811), .A2(new_n812), .B1(new_n813), .B2(new_n733), .ZN(new_n814));
  NAND2_X1  g628(.A1(new_n808), .A2(new_n814), .ZN(new_n815));
  OR2_X1    g629(.A1(new_n815), .A2(KEYINPUT116), .ZN(new_n816));
  NAND2_X1  g630(.A1(new_n815), .A2(KEYINPUT116), .ZN(new_n817));
  OAI21_X1  g631(.A(new_n797), .B1(new_n479), .B2(new_n708), .ZN(new_n818));
  NAND3_X1  g632(.A1(new_n818), .A2(new_n788), .A3(new_n804), .ZN(new_n819));
  AND2_X1   g633(.A1(new_n819), .A2(KEYINPUT51), .ZN(new_n820));
  NAND3_X1  g634(.A1(new_n816), .A2(new_n817), .A3(new_n820), .ZN(new_n821));
  INV_X1    g635(.A(KEYINPUT117), .ZN(new_n822));
  XNOR2_X1  g636(.A(new_n821), .B(new_n822), .ZN(new_n823));
  XOR2_X1   g637(.A(KEYINPUT114), .B(KEYINPUT51), .Z(new_n824));
  XNOR2_X1  g638(.A(new_n819), .B(KEYINPUT115), .ZN(new_n825));
  OAI21_X1  g639(.A(new_n824), .B1(new_n825), .B2(new_n815), .ZN(new_n826));
  NAND2_X1  g640(.A1(new_n811), .A2(new_n623), .ZN(new_n827));
  NAND2_X1  g641(.A1(new_n804), .A2(new_n732), .ZN(new_n828));
  NAND4_X1  g642(.A1(new_n827), .A2(G952), .A3(new_n272), .A4(new_n828), .ZN(new_n829));
  INV_X1    g643(.A(new_n549), .ZN(new_n830));
  AOI21_X1  g644(.A(new_n727), .B1(new_n830), .B2(new_n595), .ZN(new_n831));
  AND2_X1   g645(.A1(new_n813), .A2(new_n831), .ZN(new_n832));
  INV_X1    g646(.A(KEYINPUT118), .ZN(new_n833));
  NOR3_X1   g647(.A1(new_n832), .A2(new_n833), .A3(KEYINPUT48), .ZN(new_n834));
  XNOR2_X1  g648(.A(KEYINPUT118), .B(KEYINPUT48), .ZN(new_n835));
  AOI211_X1 g649(.A(new_n829), .B(new_n834), .C1(new_n832), .C2(new_n835), .ZN(new_n836));
  NAND3_X1  g650(.A1(new_n823), .A2(new_n826), .A3(new_n836), .ZN(new_n837));
  INV_X1    g651(.A(new_n669), .ZN(new_n838));
  NAND3_X1  g652(.A1(new_n750), .A2(new_n685), .A3(new_n671), .ZN(new_n839));
  NOR2_X1   g653(.A1(new_n839), .A2(new_n684), .ZN(new_n840));
  NAND3_X1  g654(.A1(new_n838), .A2(new_n840), .A3(new_n688), .ZN(new_n841));
  NAND4_X1  g655(.A1(new_n703), .A2(new_n677), .A3(new_n735), .A4(new_n841), .ZN(new_n842));
  NAND2_X1  g656(.A1(new_n842), .A2(KEYINPUT52), .ZN(new_n843));
  AOI22_X1  g657(.A1(new_n674), .A2(new_n676), .B1(new_n732), .B2(new_n734), .ZN(new_n844));
  INV_X1    g658(.A(KEYINPUT52), .ZN(new_n845));
  NAND4_X1  g659(.A1(new_n844), .A2(new_n845), .A3(new_n703), .A4(new_n841), .ZN(new_n846));
  NAND2_X1  g660(.A1(new_n843), .A2(new_n846), .ZN(new_n847));
  OAI21_X1  g661(.A(new_n666), .B1(new_n720), .B2(new_n675), .ZN(new_n848));
  AOI21_X1  g662(.A(new_n711), .B1(new_n628), .B2(new_n646), .ZN(new_n849));
  INV_X1    g663(.A(new_n423), .ZN(new_n850));
  INV_X1    g664(.A(KEYINPUT111), .ZN(new_n851));
  NAND4_X1  g665(.A1(new_n416), .A2(new_n771), .A3(new_n641), .A4(new_n851), .ZN(new_n852));
  AND2_X1   g666(.A1(new_n852), .A2(new_n622), .ZN(new_n853));
  OAI21_X1  g667(.A(KEYINPUT111), .B1(new_n417), .B2(new_n364), .ZN(new_n854));
  AOI21_X1  g668(.A(new_n850), .B1(new_n853), .B2(new_n854), .ZN(new_n855));
  INV_X1    g669(.A(new_n594), .ZN(new_n856));
  NOR3_X1   g670(.A1(new_n632), .A2(new_n856), .A3(new_n629), .ZN(new_n857));
  NAND4_X1  g671(.A1(new_n855), .A2(new_n429), .A3(new_n857), .A4(new_n308), .ZN(new_n858));
  NAND2_X1  g672(.A1(new_n858), .A2(new_n729), .ZN(new_n859));
  NOR4_X1   g673(.A1(new_n848), .A2(new_n849), .A3(new_n859), .A4(new_n606), .ZN(new_n860));
  NOR2_X1   g674(.A1(new_n673), .A2(new_n416), .ZN(new_n861));
  NAND3_X1  g675(.A1(new_n676), .A2(new_n788), .A3(new_n861), .ZN(new_n862));
  NAND2_X1  g676(.A1(new_n755), .A2(new_n734), .ZN(new_n863));
  AND3_X1   g677(.A1(new_n767), .A2(new_n862), .A3(new_n863), .ZN(new_n864));
  NAND3_X1  g678(.A1(new_n763), .A2(new_n860), .A3(new_n864), .ZN(new_n865));
  INV_X1    g679(.A(KEYINPUT112), .ZN(new_n866));
  NAND2_X1  g680(.A1(new_n865), .A2(new_n866), .ZN(new_n867));
  NAND4_X1  g681(.A1(new_n763), .A2(new_n860), .A3(new_n864), .A4(KEYINPUT112), .ZN(new_n868));
  AOI21_X1  g682(.A(new_n847), .B1(new_n867), .B2(new_n868), .ZN(new_n869));
  INV_X1    g683(.A(KEYINPUT53), .ZN(new_n870));
  NAND2_X1  g684(.A1(new_n867), .A2(new_n868), .ZN(new_n871));
  NAND2_X1  g685(.A1(new_n871), .A2(new_n870), .ZN(new_n872));
  AOI21_X1  g686(.A(KEYINPUT113), .B1(new_n843), .B2(new_n846), .ZN(new_n873));
  INV_X1    g687(.A(new_n873), .ZN(new_n874));
  NAND3_X1  g688(.A1(new_n843), .A2(KEYINPUT113), .A3(new_n846), .ZN(new_n875));
  NAND2_X1  g689(.A1(new_n874), .A2(new_n875), .ZN(new_n876));
  INV_X1    g690(.A(new_n876), .ZN(new_n877));
  OAI221_X1 g691(.A(KEYINPUT54), .B1(new_n869), .B2(new_n870), .C1(new_n872), .C2(new_n877), .ZN(new_n878));
  INV_X1    g692(.A(KEYINPUT54), .ZN(new_n879));
  INV_X1    g693(.A(new_n865), .ZN(new_n880));
  AND3_X1   g694(.A1(new_n843), .A2(KEYINPUT113), .A3(new_n846), .ZN(new_n881));
  OAI211_X1 g695(.A(new_n880), .B(KEYINPUT53), .C1(new_n881), .C2(new_n873), .ZN(new_n882));
  OAI211_X1 g696(.A(new_n879), .B(new_n882), .C1(new_n869), .C2(KEYINPUT53), .ZN(new_n883));
  NAND2_X1  g697(.A1(new_n878), .A2(new_n883), .ZN(new_n884));
  OAI22_X1  g698(.A1(new_n837), .A2(new_n884), .B1(G952), .B2(G953), .ZN(new_n885));
  OR2_X1    g699(.A1(new_n708), .A2(KEYINPUT49), .ZN(new_n886));
  NAND2_X1  g700(.A1(new_n708), .A2(KEYINPUT49), .ZN(new_n887));
  NOR2_X1   g701(.A1(new_n709), .A2(new_n608), .ZN(new_n888));
  NAND4_X1  g702(.A1(new_n886), .A2(new_n887), .A3(new_n772), .A4(new_n888), .ZN(new_n889));
  OR3_X1    g703(.A1(new_n695), .A2(new_n810), .A3(new_n889), .ZN(new_n890));
  NAND2_X1  g704(.A1(new_n885), .A2(new_n890), .ZN(G75));
  NOR2_X1   g705(.A1(new_n272), .A2(G952), .ZN(new_n892));
  XOR2_X1   g706(.A(new_n892), .B(KEYINPUT119), .Z(new_n893));
  INV_X1    g707(.A(new_n893), .ZN(new_n894));
  XOR2_X1   g708(.A(new_n295), .B(new_n293), .Z(new_n895));
  XNOR2_X1  g709(.A(new_n895), .B(KEYINPUT55), .ZN(new_n896));
  OAI21_X1  g710(.A(new_n882), .B1(new_n869), .B2(KEYINPUT53), .ZN(new_n897));
  NAND3_X1  g711(.A1(new_n897), .A2(G210), .A3(G902), .ZN(new_n898));
  INV_X1    g712(.A(KEYINPUT56), .ZN(new_n899));
  AOI21_X1  g713(.A(new_n896), .B1(new_n898), .B2(new_n899), .ZN(new_n900));
  NAND3_X1  g714(.A1(new_n897), .A2(G902), .A3(new_n301), .ZN(new_n901));
  AND2_X1   g715(.A1(new_n896), .A2(new_n899), .ZN(new_n902));
  AOI211_X1 g716(.A(new_n894), .B(new_n900), .C1(new_n901), .C2(new_n902), .ZN(G51));
  OR2_X1    g717(.A1(new_n869), .A2(KEYINPUT53), .ZN(new_n904));
  AOI211_X1 g718(.A(new_n407), .B(new_n781), .C1(new_n904), .C2(new_n882), .ZN(new_n905));
  NAND2_X1  g719(.A1(new_n897), .A2(KEYINPUT54), .ZN(new_n906));
  NAND2_X1  g720(.A1(new_n906), .A2(new_n883), .ZN(new_n907));
  XOR2_X1   g721(.A(new_n473), .B(KEYINPUT57), .Z(new_n908));
  AOI21_X1  g722(.A(new_n705), .B1(new_n907), .B2(new_n908), .ZN(new_n909));
  AOI21_X1  g723(.A(new_n905), .B1(new_n909), .B2(KEYINPUT120), .ZN(new_n910));
  INV_X1    g724(.A(KEYINPUT120), .ZN(new_n911));
  INV_X1    g725(.A(new_n908), .ZN(new_n912));
  AOI21_X1  g726(.A(new_n912), .B1(new_n906), .B2(new_n883), .ZN(new_n913));
  OAI21_X1  g727(.A(new_n911), .B1(new_n913), .B2(new_n705), .ZN(new_n914));
  AOI21_X1  g728(.A(new_n892), .B1(new_n910), .B2(new_n914), .ZN(G54));
  NAND4_X1  g729(.A1(new_n897), .A2(KEYINPUT58), .A3(G475), .A4(G902), .ZN(new_n916));
  INV_X1    g730(.A(new_n355), .ZN(new_n917));
  AND3_X1   g731(.A1(new_n916), .A2(KEYINPUT121), .A3(new_n917), .ZN(new_n918));
  AOI21_X1  g732(.A(KEYINPUT121), .B1(new_n916), .B2(new_n917), .ZN(new_n919));
  NOR2_X1   g733(.A1(new_n916), .A2(new_n917), .ZN(new_n920));
  NOR4_X1   g734(.A1(new_n918), .A2(new_n919), .A3(new_n920), .A4(new_n892), .ZN(G60));
  INV_X1    g735(.A(new_n618), .ZN(new_n922));
  INV_X1    g736(.A(new_n619), .ZN(new_n923));
  NAND2_X1  g737(.A1(new_n922), .A2(new_n923), .ZN(new_n924));
  NAND2_X1  g738(.A1(G478), .A2(G902), .ZN(new_n925));
  XOR2_X1   g739(.A(new_n925), .B(KEYINPUT59), .Z(new_n926));
  INV_X1    g740(.A(new_n926), .ZN(new_n927));
  NAND3_X1  g741(.A1(new_n907), .A2(new_n924), .A3(new_n927), .ZN(new_n928));
  NAND2_X1  g742(.A1(new_n928), .A2(new_n893), .ZN(new_n929));
  NAND2_X1  g743(.A1(new_n884), .A2(new_n927), .ZN(new_n930));
  INV_X1    g744(.A(KEYINPUT122), .ZN(new_n931));
  NAND4_X1  g745(.A1(new_n930), .A2(new_n931), .A3(new_n922), .A4(new_n923), .ZN(new_n932));
  AOI21_X1  g746(.A(new_n926), .B1(new_n878), .B2(new_n883), .ZN(new_n933));
  OAI21_X1  g747(.A(KEYINPUT122), .B1(new_n933), .B2(new_n924), .ZN(new_n934));
  AOI21_X1  g748(.A(new_n929), .B1(new_n932), .B2(new_n934), .ZN(G63));
  NAND2_X1  g749(.A1(G217), .A2(G902), .ZN(new_n936));
  XNOR2_X1  g750(.A(new_n936), .B(KEYINPUT60), .ZN(new_n937));
  AOI21_X1  g751(.A(new_n937), .B1(new_n904), .B2(new_n882), .ZN(new_n938));
  NAND2_X1  g752(.A1(new_n938), .A2(new_n655), .ZN(new_n939));
  OAI211_X1 g753(.A(new_n939), .B(new_n893), .C1(new_n581), .C2(new_n938), .ZN(new_n940));
  INV_X1    g754(.A(KEYINPUT61), .ZN(new_n941));
  NAND2_X1  g755(.A1(new_n940), .A2(new_n941), .ZN(new_n942));
  OR2_X1    g756(.A1(new_n938), .A2(new_n581), .ZN(new_n943));
  NAND4_X1  g757(.A1(new_n943), .A2(KEYINPUT61), .A3(new_n893), .A4(new_n939), .ZN(new_n944));
  NAND2_X1  g758(.A1(new_n942), .A2(new_n944), .ZN(G66));
  AOI21_X1  g759(.A(new_n272), .B1(new_n421), .B2(G224), .ZN(new_n946));
  INV_X1    g760(.A(new_n860), .ZN(new_n947));
  AOI21_X1  g761(.A(new_n946), .B1(new_n947), .B2(new_n272), .ZN(new_n948));
  INV_X1    g762(.A(G898), .ZN(new_n949));
  AOI21_X1  g763(.A(new_n295), .B1(new_n949), .B2(G953), .ZN(new_n950));
  XNOR2_X1  g764(.A(new_n948), .B(new_n950), .ZN(G69));
  NAND3_X1  g765(.A1(new_n494), .A2(new_n505), .A3(new_n499), .ZN(new_n952));
  XOR2_X1   g766(.A(new_n952), .B(new_n350), .Z(new_n953));
  NAND2_X1  g767(.A1(new_n853), .A2(new_n854), .ZN(new_n954));
  NAND4_X1  g768(.A1(new_n788), .A2(new_n765), .A3(new_n690), .A4(new_n954), .ZN(new_n955));
  AND3_X1   g769(.A1(new_n799), .A2(new_n792), .A3(new_n955), .ZN(new_n956));
  AND2_X1   g770(.A1(new_n844), .A2(new_n703), .ZN(new_n957));
  NAND2_X1  g771(.A1(new_n957), .A2(new_n696), .ZN(new_n958));
  OR2_X1    g772(.A1(new_n958), .A2(KEYINPUT62), .ZN(new_n959));
  NAND2_X1  g773(.A1(new_n958), .A2(KEYINPUT62), .ZN(new_n960));
  AND3_X1   g774(.A1(new_n956), .A2(new_n959), .A3(new_n960), .ZN(new_n961));
  OAI21_X1  g775(.A(new_n953), .B1(new_n961), .B2(G953), .ZN(new_n962));
  OR2_X1    g776(.A1(new_n272), .A2(G900), .ZN(new_n963));
  NAND2_X1  g777(.A1(new_n962), .A2(new_n963), .ZN(new_n964));
  NAND4_X1  g778(.A1(new_n786), .A2(new_n838), .A3(new_n688), .A4(new_n831), .ZN(new_n965));
  NAND4_X1  g779(.A1(new_n799), .A2(new_n792), .A3(new_n957), .A4(new_n965), .ZN(new_n966));
  AND2_X1   g780(.A1(new_n763), .A2(new_n767), .ZN(new_n967));
  OR2_X1    g781(.A1(new_n967), .A2(KEYINPUT123), .ZN(new_n968));
  NAND2_X1  g782(.A1(new_n967), .A2(KEYINPUT123), .ZN(new_n969));
  AOI21_X1  g783(.A(new_n966), .B1(new_n968), .B2(new_n969), .ZN(new_n970));
  NOR3_X1   g784(.A1(new_n970), .A2(G953), .A3(new_n953), .ZN(new_n971));
  AOI21_X1  g785(.A(new_n272), .B1(G227), .B2(G900), .ZN(new_n972));
  OAI22_X1  g786(.A1(new_n964), .A2(new_n971), .B1(KEYINPUT124), .B2(new_n972), .ZN(new_n973));
  NAND2_X1  g787(.A1(new_n972), .A2(KEYINPUT124), .ZN(new_n974));
  XOR2_X1   g788(.A(new_n974), .B(KEYINPUT125), .Z(new_n975));
  INV_X1    g789(.A(new_n975), .ZN(new_n976));
  NAND2_X1  g790(.A1(new_n973), .A2(new_n976), .ZN(new_n977));
  OAI221_X1 g791(.A(new_n975), .B1(KEYINPUT124), .B2(new_n972), .C1(new_n964), .C2(new_n971), .ZN(new_n978));
  NAND2_X1  g792(.A1(new_n977), .A2(new_n978), .ZN(G72));
  INV_X1    g793(.A(new_n679), .ZN(new_n980));
  NOR2_X1   g794(.A1(new_n980), .A2(new_n681), .ZN(new_n981));
  AND2_X1   g795(.A1(new_n970), .A2(new_n860), .ZN(new_n982));
  NAND2_X1  g796(.A1(G472), .A2(G902), .ZN(new_n983));
  XOR2_X1   g797(.A(new_n983), .B(KEYINPUT63), .Z(new_n984));
  INV_X1    g798(.A(new_n984), .ZN(new_n985));
  OAI21_X1  g799(.A(new_n981), .B1(new_n982), .B2(new_n985), .ZN(new_n986));
  NOR3_X1   g800(.A1(new_n981), .A2(new_n680), .A3(new_n985), .ZN(new_n987));
  XNOR2_X1  g801(.A(new_n987), .B(KEYINPUT126), .ZN(new_n988));
  OAI221_X1 g802(.A(new_n988), .B1(new_n869), .B2(new_n870), .C1(new_n872), .C2(new_n877), .ZN(new_n989));
  NAND3_X1  g803(.A1(new_n956), .A2(new_n959), .A3(new_n960), .ZN(new_n990));
  OAI21_X1  g804(.A(new_n984), .B1(new_n990), .B2(new_n947), .ZN(new_n991));
  AOI21_X1  g805(.A(new_n892), .B1(new_n991), .B2(new_n680), .ZN(new_n992));
  NAND3_X1  g806(.A1(new_n986), .A2(new_n989), .A3(new_n992), .ZN(new_n993));
  INV_X1    g807(.A(KEYINPUT127), .ZN(new_n994));
  NAND2_X1  g808(.A1(new_n993), .A2(new_n994), .ZN(new_n995));
  NAND4_X1  g809(.A1(new_n986), .A2(new_n992), .A3(KEYINPUT127), .A4(new_n989), .ZN(new_n996));
  NAND2_X1  g810(.A1(new_n995), .A2(new_n996), .ZN(G57));
endmodule


