

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n352, n353, n354, n355, n356, n357, n358, n359, n360, n361, n362,
         n363, n364, n365, n366, n367, n368, n369, n370, n371, n372, n373,
         n374, n375, n376, n377, n378, n379, n380, n381, n382, n383, n384,
         n385, n386, n387, n388, n389, n390, n391, n392, n393, n394, n395,
         n396, n397, n398, n399, n400, n401, n402, n403, n404, n405, n406,
         n407, n408, n409, n410, n411, n412, n413, n414, n415, n416, n417,
         n418, n419, n420, n421, n422, n423, n424, n425, n426, n427, n428,
         n429, n430, n431, n432, n433, n434, n435, n436, n437, n438, n439,
         n440, n441, n442, n443, n444, n445, n446, n447, n448, n449, n450,
         n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, n461,
         n462, n463, n464, n465, n466, n467, n468, n469, n470, n471, n472,
         n473, n474, n475, n476, n477, n478, n479, n480, n481, n482, n483,
         n484, n485, n486, n487, n488, n489, n490, n491, n492, n493, n494,
         n495, n496, n497, n498, n499, n500, n501, n502, n503, n504, n505,
         n506, n507, n508, n509, n510, n511, n512, n513, n514, n515, n516,
         n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527,
         n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538,
         n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549,
         n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560,
         n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571,
         n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582,
         n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593,
         n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604,
         n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615,
         n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626,
         n627, n628, n629, n630, n631, n632, n633, n634, n635, n636, n637,
         n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, n648,
         n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659,
         n660, n661, n662, n663, n664, n665, n666, n667, n668, n669, n670,
         n671, n672, n673, n674, n675, n676, n677, n678, n679, n680, n681,
         n682, n683, n684, n685, n686, n687, n688, n689, n690, n691, n692,
         n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, n703,
         n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, n714,
         n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, n725,
         n726, n727, n728, n729, n730, n731, n732, n733, n734, n735, n736,
         n737, n738, n739, n740, n741, n742, n743, n744, n745, n746, n747,
         n748, n749, n750, n751, n752, n753, n754, n755, n756, n757, n758;

  XNOR2_X1 U373 ( .A(n573), .B(n572), .ZN(n581) );
  AND2_X1 U374 ( .A1(n571), .A2(n570), .ZN(n573) );
  NOR2_X1 U375 ( .A1(n616), .A2(n449), .ZN(n419) );
  NOR2_X2 U376 ( .A1(n673), .A2(n672), .ZN(n575) );
  NOR2_X2 U377 ( .A1(n757), .A2(n758), .ZN(n422) );
  AND2_X4 U378 ( .A1(n398), .A2(n410), .ZN(n710) );
  AND2_X2 U379 ( .A1(n370), .A2(n362), .ZN(n398) );
  AND2_X2 U380 ( .A1(n600), .A2(n421), .ZN(n420) );
  OR2_X2 U381 ( .A1(n696), .A2(n642), .ZN(n447) );
  XNOR2_X2 U382 ( .A(n500), .B(n465), .ZN(n746) );
  NOR2_X2 U383 ( .A1(n533), .A2(n532), .ZN(n534) );
  XNOR2_X2 U384 ( .A(n565), .B(KEYINPUT38), .ZN(n670) );
  XNOR2_X1 U385 ( .A(n553), .B(n552), .ZN(n616) );
  NAND2_X1 U386 ( .A1(n655), .A2(n747), .ZN(n652) );
  XNOR2_X1 U387 ( .A(n636), .B(KEYINPUT45), .ZN(n655) );
  NOR2_X1 U388 ( .A1(n599), .A2(n428), .ZN(n600) );
  XNOR2_X1 U389 ( .A(n402), .B(KEYINPUT72), .ZN(n587) );
  XNOR2_X1 U390 ( .A(n544), .B(n543), .ZN(n631) );
  NOR2_X1 U391 ( .A1(n616), .A2(n593), .ZN(n569) );
  AND2_X1 U392 ( .A1(n408), .A2(n407), .ZN(n406) );
  XNOR2_X1 U393 ( .A(n484), .B(n483), .ZN(n662) );
  XNOR2_X1 U394 ( .A(n424), .B(n423), .ZN(n495) );
  XNOR2_X1 U395 ( .A(n430), .B(KEYINPUT3), .ZN(n424) );
  XNOR2_X1 U396 ( .A(KEYINPUT71), .B(KEYINPUT16), .ZN(n431) );
  XNOR2_X1 U397 ( .A(n624), .B(n623), .ZN(n677) );
  BUF_X1 U398 ( .A(n757), .Z(n352) );
  BUF_X1 U399 ( .A(n577), .Z(n353) );
  XNOR2_X1 U400 ( .A(n399), .B(G472), .ZN(n354) );
  XNOR2_X1 U401 ( .A(n395), .B(n579), .ZN(n757) );
  XNOR2_X1 U402 ( .A(n399), .B(G472), .ZN(n553) );
  NOR2_X1 U403 ( .A1(n677), .A2(n533), .ZN(n413) );
  XOR2_X2 U404 ( .A(KEYINPUT42), .B(n576), .Z(n758) );
  XNOR2_X2 U405 ( .A(n411), .B(n626), .ZN(n702) );
  XNOR2_X1 U406 ( .A(n511), .B(n510), .ZN(n647) );
  XNOR2_X1 U407 ( .A(n659), .B(KEYINPUT50), .ZN(n380) );
  NAND2_X1 U408 ( .A1(n721), .A2(n631), .ZN(n394) );
  NAND2_X1 U409 ( .A1(n383), .A2(n382), .ZN(n381) );
  XNOR2_X1 U410 ( .A(n668), .B(n384), .ZN(n383) );
  XNOR2_X1 U411 ( .A(n385), .B(KEYINPUT51), .ZN(n384) );
  XNOR2_X1 U412 ( .A(G128), .B(KEYINPUT90), .ZN(n467) );
  INV_X1 U413 ( .A(G237), .ZN(n444) );
  BUF_X1 U414 ( .A(n541), .Z(n377) );
  INV_X1 U415 ( .A(n564), .ZN(n405) );
  XNOR2_X1 U416 ( .A(KEYINPUT68), .B(KEYINPUT0), .ZN(n455) );
  XNOR2_X1 U417 ( .A(n514), .B(n513), .ZN(n563) );
  XNOR2_X1 U418 ( .A(n379), .B(n378), .ZN(n667) );
  INV_X1 U419 ( .A(KEYINPUT115), .ZN(n378) );
  NAND2_X1 U420 ( .A1(n380), .A2(n359), .ZN(n379) );
  INV_X1 U421 ( .A(KEYINPUT116), .ZN(n385) );
  NAND2_X1 U422 ( .A1(n725), .A2(n356), .ZN(n402) );
  INV_X1 U423 ( .A(n674), .ZN(n391) );
  XNOR2_X1 U424 ( .A(n394), .B(n393), .ZN(n392) );
  INV_X1 U425 ( .A(KEYINPUT97), .ZN(n393) );
  NOR2_X1 U426 ( .A1(G237), .A2(G953), .ZN(n496) );
  XNOR2_X1 U427 ( .A(n381), .B(KEYINPUT117), .ZN(n680) );
  AND2_X1 U428 ( .A1(n540), .A2(n620), .ZN(n417) );
  XNOR2_X1 U429 ( .A(KEYINPUT95), .B(KEYINPUT5), .ZN(n492) );
  XOR2_X1 U430 ( .A(G101), .B(G137), .Z(n493) );
  XOR2_X1 U431 ( .A(KEYINPUT84), .B(KEYINPUT8), .Z(n472) );
  XNOR2_X1 U432 ( .A(G113), .B(G143), .ZN(n507) );
  INV_X1 U433 ( .A(G128), .ZN(n437) );
  XNOR2_X1 U434 ( .A(G119), .B(G116), .ZN(n423) );
  XNOR2_X1 U435 ( .A(G119), .B(G110), .ZN(n466) );
  XOR2_X1 U436 ( .A(G122), .B(G107), .Z(n521) );
  XNOR2_X1 U437 ( .A(G107), .B(G104), .ZN(n433) );
  XNOR2_X1 U438 ( .A(KEYINPUT17), .B(KEYINPUT18), .ZN(n440) );
  XNOR2_X1 U439 ( .A(G146), .B(G125), .ZN(n475) );
  XNOR2_X1 U440 ( .A(n373), .B(n372), .ZN(n683) );
  INV_X1 U441 ( .A(KEYINPUT118), .ZN(n372) );
  NAND2_X1 U442 ( .A1(n374), .A2(n355), .ZN(n373) );
  NOR2_X1 U443 ( .A1(n607), .A2(n377), .ZN(n609) );
  XNOR2_X1 U444 ( .A(n561), .B(KEYINPUT75), .ZN(n577) );
  XNOR2_X1 U445 ( .A(n419), .B(KEYINPUT30), .ZN(n560) );
  NAND2_X1 U446 ( .A1(n405), .A2(n404), .ZN(n403) );
  XNOR2_X1 U447 ( .A(n647), .B(n646), .ZN(n648) );
  NAND2_X1 U448 ( .A1(n652), .A2(n641), .ZN(n410) );
  NOR2_X1 U449 ( .A1(n748), .A2(G952), .ZN(n718) );
  OR2_X1 U450 ( .A1(n683), .A2(KEYINPUT119), .ZN(n368) );
  INV_X2 U451 ( .A(G953), .ZN(n748) );
  NAND2_X1 U452 ( .A1(n597), .A2(n377), .ZN(n731) );
  NAND2_X1 U453 ( .A1(n405), .A2(n669), .ZN(n594) );
  XNOR2_X1 U454 ( .A(n426), .B(n425), .ZN(n629) );
  INV_X1 U455 ( .A(KEYINPUT105), .ZN(n425) );
  NAND2_X1 U456 ( .A1(n427), .A2(n619), .ZN(n426) );
  XNOR2_X1 U457 ( .A(n618), .B(KEYINPUT65), .ZN(n427) );
  INV_X1 U458 ( .A(G110), .ZN(n687) );
  NAND2_X1 U459 ( .A1(n501), .A2(n660), .ZN(n721) );
  OR2_X1 U460 ( .A1(n682), .A2(n677), .ZN(n355) );
  XNOR2_X1 U461 ( .A(n575), .B(n574), .ZN(n682) );
  NOR2_X1 U462 ( .A1(n674), .A2(KEYINPUT47), .ZN(n356) );
  AND2_X1 U463 ( .A1(n548), .A2(n658), .ZN(n617) );
  AND2_X1 U464 ( .A1(n747), .A2(n654), .ZN(n357) );
  NAND2_X1 U465 ( .A1(n683), .A2(KEYINPUT119), .ZN(n358) );
  NOR2_X1 U466 ( .A1(n665), .A2(n354), .ZN(n359) );
  BUF_X1 U467 ( .A(n564), .Z(n565) );
  AND2_X1 U468 ( .A1(n368), .A2(n748), .ZN(n360) );
  AND2_X1 U469 ( .A1(G952), .A2(n656), .ZN(n361) );
  OR2_X1 U470 ( .A1(n643), .A2(n642), .ZN(n362) );
  AND2_X1 U471 ( .A1(n536), .A2(n541), .ZN(n537) );
  NAND2_X1 U472 ( .A1(n601), .A2(n729), .ZN(n395) );
  AND2_X1 U473 ( .A1(n416), .A2(n622), .ZN(n415) );
  NAND2_X1 U474 ( .A1(n621), .A2(KEYINPUT106), .ZN(n414) );
  AND2_X2 U475 ( .A1(n702), .A2(n627), .ZN(n628) );
  AND2_X1 U476 ( .A1(n616), .A2(n658), .ZN(n363) );
  NAND2_X1 U477 ( .A1(n406), .A2(n403), .ZN(n580) );
  NAND2_X1 U478 ( .A1(n652), .A2(n644), .ZN(n388) );
  NAND2_X1 U479 ( .A1(n364), .A2(n360), .ZN(n685) );
  NAND2_X1 U480 ( .A1(n366), .A2(n365), .ZN(n364) );
  NAND2_X1 U481 ( .A1(n710), .A2(G475), .ZN(n397) );
  XNOR2_X1 U482 ( .A(n397), .B(n648), .ZN(n649) );
  NAND2_X1 U483 ( .A1(n369), .A2(n358), .ZN(n365) );
  NAND2_X1 U484 ( .A1(n367), .A2(KEYINPUT119), .ZN(n366) );
  INV_X1 U485 ( .A(n369), .ZN(n367) );
  XNOR2_X1 U486 ( .A(n418), .B(KEYINPUT86), .ZN(n369) );
  NAND2_X1 U487 ( .A1(n386), .A2(n370), .ZN(n418) );
  NAND2_X1 U488 ( .A1(n401), .A2(KEYINPUT2), .ZN(n370) );
  NAND2_X1 U489 ( .A1(n628), .A2(n629), .ZN(n371) );
  XNOR2_X1 U490 ( .A(n371), .B(n630), .ZN(n635) );
  NAND2_X1 U491 ( .A1(n415), .A2(n414), .ZN(n624) );
  INV_X1 U492 ( .A(n682), .ZN(n382) );
  NAND2_X1 U493 ( .A1(n375), .A2(n361), .ZN(n374) );
  XNOR2_X1 U494 ( .A(n681), .B(n376), .ZN(n375) );
  INV_X1 U495 ( .A(KEYINPUT52), .ZN(n376) );
  INV_X1 U496 ( .A(n377), .ZN(n658) );
  NAND2_X1 U497 ( .A1(n389), .A2(n387), .ZN(n386) );
  NAND2_X1 U498 ( .A1(n388), .A2(n653), .ZN(n387) );
  NAND2_X1 U499 ( .A1(n390), .A2(n357), .ZN(n389) );
  INV_X1 U500 ( .A(n734), .ZN(n390) );
  NAND2_X1 U501 ( .A1(n392), .A2(n391), .ZN(n632) );
  AND2_X2 U502 ( .A1(n615), .A2(n614), .ZN(n747) );
  XNOR2_X2 U503 ( .A(n396), .B(n578), .ZN(n601) );
  NAND2_X1 U504 ( .A1(n577), .A2(n670), .ZN(n396) );
  NAND2_X1 U505 ( .A1(n688), .A2(n527), .ZN(n399) );
  XNOR2_X1 U506 ( .A(n400), .B(n500), .ZN(n688) );
  XNOR2_X1 U507 ( .A(n499), .B(n498), .ZN(n400) );
  INV_X1 U508 ( .A(n652), .ZN(n401) );
  INV_X1 U509 ( .A(n725), .ZN(n585) );
  XNOR2_X2 U510 ( .A(n582), .B(KEYINPUT79), .ZN(n725) );
  NOR2_X1 U511 ( .A1(n449), .A2(n450), .ZN(n404) );
  NAND2_X1 U512 ( .A1(n449), .A2(n450), .ZN(n407) );
  NAND2_X1 U513 ( .A1(n564), .A2(n450), .ZN(n408) );
  XNOR2_X2 U514 ( .A(n409), .B(n455), .ZN(n533) );
  NAND2_X1 U515 ( .A1(n580), .A2(n454), .ZN(n409) );
  NAND2_X1 U516 ( .A1(n635), .A2(n634), .ZN(n636) );
  NAND2_X1 U517 ( .A1(n710), .A2(G210), .ZN(n698) );
  NAND2_X1 U518 ( .A1(n412), .A2(n625), .ZN(n411) );
  XNOR2_X1 U519 ( .A(n413), .B(KEYINPUT34), .ZN(n412) );
  NAND2_X1 U520 ( .A1(n417), .A2(n541), .ZN(n416) );
  NAND2_X1 U521 ( .A1(n541), .A2(n540), .ZN(n621) );
  XNOR2_X2 U522 ( .A(n570), .B(KEYINPUT1), .ZN(n541) );
  XNOR2_X1 U523 ( .A(n420), .B(KEYINPUT48), .ZN(n615) );
  XNOR2_X1 U524 ( .A(n422), .B(KEYINPUT46), .ZN(n421) );
  INV_X1 U525 ( .A(n629), .ZN(n686) );
  BUF_X1 U526 ( .A(n655), .Z(n734) );
  XNOR2_X2 U527 ( .A(n516), .B(KEYINPUT4), .ZN(n457) );
  XNOR2_X2 U528 ( .A(n438), .B(n437), .ZN(n516) );
  BUF_X1 U529 ( .A(n739), .Z(n740) );
  NAND2_X1 U530 ( .A1(n598), .A2(n731), .ZN(n428) );
  AND2_X1 U531 ( .A1(G214), .A2(n506), .ZN(n429) );
  INV_X1 U532 ( .A(n657), .ZN(n540) );
  XNOR2_X1 U533 ( .A(n429), .B(n509), .ZN(n510) );
  XNOR2_X1 U534 ( .A(n512), .B(G475), .ZN(n513) );
  INV_X1 U535 ( .A(KEYINPUT40), .ZN(n579) );
  XNOR2_X2 U536 ( .A(G113), .B(KEYINPUT70), .ZN(n430) );
  XNOR2_X1 U537 ( .A(n431), .B(G122), .ZN(n432) );
  XNOR2_X1 U538 ( .A(n495), .B(n432), .ZN(n436) );
  XNOR2_X1 U539 ( .A(n433), .B(n687), .ZN(n435) );
  XNOR2_X1 U540 ( .A(G101), .B(KEYINPUT73), .ZN(n434) );
  XNOR2_X1 U541 ( .A(n435), .B(n434), .ZN(n460) );
  XNOR2_X1 U542 ( .A(n436), .B(n460), .ZN(n739) );
  XNOR2_X2 U543 ( .A(G143), .B(KEYINPUT64), .ZN(n438) );
  NAND2_X1 U544 ( .A1(n748), .A2(G224), .ZN(n439) );
  XNOR2_X1 U545 ( .A(n440), .B(n439), .ZN(n441) );
  XNOR2_X1 U546 ( .A(n475), .B(n441), .ZN(n442) );
  XNOR2_X1 U547 ( .A(n457), .B(n442), .ZN(n443) );
  XNOR2_X1 U548 ( .A(n739), .B(n443), .ZN(n696) );
  XNOR2_X1 U549 ( .A(G902), .B(KEYINPUT15), .ZN(n637) );
  INV_X1 U550 ( .A(n637), .ZN(n642) );
  INV_X1 U551 ( .A(G902), .ZN(n527) );
  NAND2_X1 U552 ( .A1(n527), .A2(n444), .ZN(n448) );
  NAND2_X1 U553 ( .A1(n448), .A2(G210), .ZN(n445) );
  XNOR2_X1 U554 ( .A(n445), .B(KEYINPUT80), .ZN(n446) );
  XNOR2_X2 U555 ( .A(n447), .B(n446), .ZN(n564) );
  NAND2_X1 U556 ( .A1(n448), .A2(G214), .ZN(n669) );
  INV_X1 U557 ( .A(n669), .ZN(n449) );
  XNOR2_X1 U558 ( .A(KEYINPUT76), .B(KEYINPUT19), .ZN(n450) );
  NOR2_X1 U559 ( .A1(G898), .A2(n748), .ZN(n741) );
  NAND2_X1 U560 ( .A1(n741), .A2(G902), .ZN(n451) );
  NAND2_X1 U561 ( .A1(n748), .A2(G952), .ZN(n556) );
  NAND2_X1 U562 ( .A1(n451), .A2(n556), .ZN(n453) );
  NAND2_X1 U563 ( .A1(G237), .A2(G234), .ZN(n452) );
  XNOR2_X1 U564 ( .A(n452), .B(KEYINPUT14), .ZN(n656) );
  AND2_X1 U565 ( .A1(n453), .A2(n656), .ZN(n454) );
  XNOR2_X1 U566 ( .A(G134), .B(G131), .ZN(n456) );
  XNOR2_X2 U567 ( .A(n457), .B(n456), .ZN(n500) );
  XNOR2_X2 U568 ( .A(G140), .B(G137), .ZN(n465) );
  NAND2_X1 U569 ( .A1(n748), .A2(G227), .ZN(n458) );
  XNOR2_X1 U570 ( .A(n458), .B(G146), .ZN(n459) );
  XNOR2_X1 U571 ( .A(n460), .B(n459), .ZN(n461) );
  XNOR2_X1 U572 ( .A(n746), .B(n461), .ZN(n711) );
  OR2_X2 U573 ( .A1(n711), .A2(G902), .ZN(n464) );
  INV_X1 U574 ( .A(KEYINPUT69), .ZN(n462) );
  XNOR2_X1 U575 ( .A(n462), .B(G469), .ZN(n463) );
  XNOR2_X2 U576 ( .A(n464), .B(n463), .ZN(n570) );
  INV_X1 U577 ( .A(n570), .ZN(n488) );
  XNOR2_X1 U578 ( .A(n466), .B(n465), .ZN(n470) );
  XOR2_X1 U579 ( .A(KEYINPUT91), .B(KEYINPUT24), .Z(n468) );
  XNOR2_X1 U580 ( .A(n468), .B(n467), .ZN(n469) );
  XNOR2_X1 U581 ( .A(n470), .B(n469), .ZN(n474) );
  NAND2_X1 U582 ( .A1(G234), .A2(n748), .ZN(n471) );
  XNOR2_X1 U583 ( .A(n472), .B(n471), .ZN(n515) );
  NAND2_X1 U584 ( .A1(G221), .A2(n515), .ZN(n473) );
  XNOR2_X1 U585 ( .A(n474), .B(n473), .ZN(n478) );
  XNOR2_X1 U586 ( .A(n475), .B(KEYINPUT10), .ZN(n745) );
  XNOR2_X1 U587 ( .A(KEYINPUT83), .B(KEYINPUT23), .ZN(n476) );
  XNOR2_X1 U588 ( .A(n745), .B(n476), .ZN(n477) );
  XNOR2_X1 U589 ( .A(n478), .B(n477), .ZN(n704) );
  NAND2_X1 U590 ( .A1(n704), .A2(n527), .ZN(n484) );
  NAND2_X1 U591 ( .A1(n637), .A2(G234), .ZN(n479) );
  XNOR2_X1 U592 ( .A(n479), .B(KEYINPUT20), .ZN(n485) );
  NAND2_X1 U593 ( .A1(n485), .A2(G217), .ZN(n482) );
  XNOR2_X1 U594 ( .A(KEYINPUT92), .B(KEYINPUT25), .ZN(n480) );
  XNOR2_X1 U595 ( .A(n480), .B(KEYINPUT77), .ZN(n481) );
  XNOR2_X1 U596 ( .A(n482), .B(n481), .ZN(n483) );
  NAND2_X1 U597 ( .A1(n485), .A2(G221), .ZN(n487) );
  XNOR2_X1 U598 ( .A(KEYINPUT21), .B(KEYINPUT93), .ZN(n486) );
  XNOR2_X1 U599 ( .A(n487), .B(n486), .ZN(n661) );
  NAND2_X1 U600 ( .A1(n662), .A2(n661), .ZN(n657) );
  OR2_X1 U601 ( .A1(n488), .A2(n657), .ZN(n489) );
  OR2_X1 U602 ( .A1(n533), .A2(n489), .ZN(n491) );
  INV_X1 U603 ( .A(KEYINPUT94), .ZN(n490) );
  XNOR2_X1 U604 ( .A(n491), .B(n490), .ZN(n501) );
  XNOR2_X1 U605 ( .A(n493), .B(n492), .ZN(n494) );
  XNOR2_X1 U606 ( .A(n495), .B(n494), .ZN(n499) );
  XNOR2_X1 U607 ( .A(n496), .B(KEYINPUT74), .ZN(n506) );
  NAND2_X1 U608 ( .A1(G210), .A2(n506), .ZN(n497) );
  XNOR2_X1 U609 ( .A(n497), .B(G146), .ZN(n498) );
  INV_X1 U610 ( .A(n354), .ZN(n660) );
  XOR2_X1 U611 ( .A(KEYINPUT12), .B(KEYINPUT98), .Z(n505) );
  XNOR2_X1 U612 ( .A(G104), .B(G122), .ZN(n502) );
  XNOR2_X1 U613 ( .A(n502), .B(KEYINPUT11), .ZN(n503) );
  XNOR2_X1 U614 ( .A(n745), .B(n503), .ZN(n504) );
  XNOR2_X1 U615 ( .A(n505), .B(n504), .ZN(n511) );
  XOR2_X1 U616 ( .A(G140), .B(G131), .Z(n508) );
  XNOR2_X1 U617 ( .A(n508), .B(n507), .ZN(n509) );
  NOR2_X1 U618 ( .A1(G902), .A2(n647), .ZN(n514) );
  XNOR2_X1 U619 ( .A(KEYINPUT99), .B(KEYINPUT13), .ZN(n512) );
  NAND2_X1 U620 ( .A1(G217), .A2(n515), .ZN(n518) );
  INV_X1 U621 ( .A(n516), .ZN(n517) );
  XNOR2_X1 U622 ( .A(n518), .B(n517), .ZN(n526) );
  XOR2_X1 U623 ( .A(KEYINPUT100), .B(KEYINPUT9), .Z(n520) );
  XNOR2_X1 U624 ( .A(KEYINPUT101), .B(KEYINPUT7), .ZN(n519) );
  XNOR2_X1 U625 ( .A(n520), .B(n519), .ZN(n524) );
  XNOR2_X1 U626 ( .A(G116), .B(G134), .ZN(n522) );
  XNOR2_X1 U627 ( .A(n522), .B(n521), .ZN(n523) );
  XNOR2_X1 U628 ( .A(n524), .B(n523), .ZN(n525) );
  XNOR2_X1 U629 ( .A(n526), .B(n525), .ZN(n706) );
  NAND2_X1 U630 ( .A1(n706), .A2(n527), .ZN(n529) );
  INV_X1 U631 ( .A(G478), .ZN(n528) );
  XNOR2_X1 U632 ( .A(n529), .B(n528), .ZN(n562) );
  INV_X1 U633 ( .A(n562), .ZN(n546) );
  OR2_X1 U634 ( .A1(n563), .A2(n546), .ZN(n584) );
  NOR2_X1 U635 ( .A1(n721), .A2(n584), .ZN(n530) );
  XOR2_X1 U636 ( .A(G104), .B(n530), .Z(G6) );
  NAND2_X1 U637 ( .A1(n563), .A2(n562), .ZN(n672) );
  INV_X1 U638 ( .A(n661), .ZN(n531) );
  OR2_X1 U639 ( .A1(n672), .A2(n531), .ZN(n532) );
  XNOR2_X1 U640 ( .A(n534), .B(KEYINPUT22), .ZN(n548) );
  INV_X1 U641 ( .A(KEYINPUT6), .ZN(n535) );
  XNOR2_X1 U642 ( .A(n354), .B(n535), .ZN(n622) );
  NOR2_X1 U643 ( .A1(n622), .A2(n662), .ZN(n536) );
  XNOR2_X1 U644 ( .A(n537), .B(KEYINPUT78), .ZN(n538) );
  NAND2_X1 U645 ( .A1(n548), .A2(n538), .ZN(n539) );
  XNOR2_X1 U646 ( .A(n539), .B(KEYINPUT32), .ZN(n627) );
  XNOR2_X1 U647 ( .A(n627), .B(G119), .ZN(G21) );
  OR2_X1 U648 ( .A1(n621), .A2(n660), .ZN(n666) );
  OR2_X1 U649 ( .A1(n666), .A2(n533), .ZN(n544) );
  INV_X1 U650 ( .A(KEYINPUT96), .ZN(n542) );
  XNOR2_X1 U651 ( .A(n542), .B(KEYINPUT31), .ZN(n543) );
  NOR2_X1 U652 ( .A1(n631), .A2(n584), .ZN(n545) );
  XOR2_X1 U653 ( .A(G113), .B(n545), .Z(G15) );
  AND2_X1 U654 ( .A1(n563), .A2(n546), .ZN(n726) );
  INV_X1 U655 ( .A(n726), .ZN(n720) );
  NOR2_X1 U656 ( .A1(n631), .A2(n720), .ZN(n547) );
  XOR2_X1 U657 ( .A(G116), .B(n547), .Z(G18) );
  INV_X1 U658 ( .A(n662), .ZN(n619) );
  NOR2_X1 U659 ( .A1(n622), .A2(n619), .ZN(n549) );
  NAND2_X1 U660 ( .A1(n617), .A2(n549), .ZN(n551) );
  INV_X1 U661 ( .A(KEYINPUT103), .ZN(n550) );
  XNOR2_X1 U662 ( .A(n551), .B(n550), .ZN(n633) );
  XNOR2_X1 U663 ( .A(n633), .B(G101), .ZN(G3) );
  INV_X1 U664 ( .A(KEYINPUT104), .ZN(n552) );
  NOR2_X1 U665 ( .A1(G900), .A2(n748), .ZN(n554) );
  NAND2_X1 U666 ( .A1(G902), .A2(n554), .ZN(n555) );
  NAND2_X1 U667 ( .A1(n556), .A2(n555), .ZN(n557) );
  NAND2_X1 U668 ( .A1(n557), .A2(n656), .ZN(n567) );
  NOR2_X1 U669 ( .A1(n657), .A2(n567), .ZN(n558) );
  AND2_X1 U670 ( .A1(n570), .A2(n558), .ZN(n559) );
  NAND2_X1 U671 ( .A1(n560), .A2(n559), .ZN(n561) );
  NOR2_X1 U672 ( .A1(n563), .A2(n562), .ZN(n625) );
  AND2_X1 U673 ( .A1(n625), .A2(n405), .ZN(n566) );
  NAND2_X1 U674 ( .A1(n353), .A2(n566), .ZN(n589) );
  XNOR2_X1 U675 ( .A(n589), .B(G143), .ZN(G45) );
  NOR2_X1 U676 ( .A1(n662), .A2(n567), .ZN(n568) );
  NAND2_X1 U677 ( .A1(n568), .A2(n661), .ZN(n593) );
  XNOR2_X1 U678 ( .A(KEYINPUT28), .B(n569), .ZN(n571) );
  INV_X1 U679 ( .A(KEYINPUT109), .ZN(n572) );
  NAND2_X1 U680 ( .A1(n670), .A2(n669), .ZN(n673) );
  XNOR2_X1 U681 ( .A(KEYINPUT110), .B(KEYINPUT41), .ZN(n574) );
  NAND2_X1 U682 ( .A1(n581), .A2(n382), .ZN(n576) );
  XOR2_X1 U683 ( .A(KEYINPUT87), .B(KEYINPUT39), .Z(n578) );
  INV_X1 U684 ( .A(n584), .ZN(n729) );
  NAND2_X1 U685 ( .A1(n581), .A2(n580), .ZN(n582) );
  INV_X1 U686 ( .A(KEYINPUT102), .ZN(n583) );
  XNOR2_X1 U687 ( .A(n726), .B(n583), .ZN(n602) );
  AND2_X1 U688 ( .A1(n602), .A2(n584), .ZN(n674) );
  NAND2_X1 U689 ( .A1(n585), .A2(KEYINPUT47), .ZN(n586) );
  NAND2_X1 U690 ( .A1(n587), .A2(n586), .ZN(n599) );
  NAND2_X1 U691 ( .A1(n674), .A2(KEYINPUT47), .ZN(n588) );
  XNOR2_X1 U692 ( .A(KEYINPUT82), .B(n588), .ZN(n590) );
  NAND2_X1 U693 ( .A1(n590), .A2(n589), .ZN(n591) );
  XNOR2_X1 U694 ( .A(n591), .B(KEYINPUT81), .ZN(n598) );
  NAND2_X1 U695 ( .A1(n622), .A2(n729), .ZN(n592) );
  NOR2_X1 U696 ( .A1(n593), .A2(n592), .ZN(n605) );
  XNOR2_X1 U697 ( .A(KEYINPUT111), .B(n605), .ZN(n595) );
  NOR2_X1 U698 ( .A1(n595), .A2(n594), .ZN(n596) );
  XNOR2_X1 U699 ( .A(n596), .B(KEYINPUT36), .ZN(n597) );
  BUF_X1 U700 ( .A(n601), .Z(n604) );
  INV_X1 U701 ( .A(n602), .ZN(n603) );
  NAND2_X1 U702 ( .A1(n604), .A2(n603), .ZN(n733) );
  INV_X1 U703 ( .A(n733), .ZN(n613) );
  NAND2_X1 U704 ( .A1(n605), .A2(n669), .ZN(n606) );
  XOR2_X1 U705 ( .A(KEYINPUT107), .B(n606), .Z(n607) );
  INV_X1 U706 ( .A(KEYINPUT43), .ZN(n608) );
  XNOR2_X1 U707 ( .A(n609), .B(n608), .ZN(n610) );
  NAND2_X1 U708 ( .A1(n610), .A2(n565), .ZN(n612) );
  INV_X1 U709 ( .A(KEYINPUT108), .ZN(n611) );
  XNOR2_X1 U710 ( .A(n612), .B(n611), .ZN(n755) );
  NOR2_X1 U711 ( .A1(n613), .A2(n755), .ZN(n614) );
  NAND2_X1 U712 ( .A1(n363), .A2(n548), .ZN(n618) );
  INV_X1 U713 ( .A(KEYINPUT106), .ZN(n620) );
  INV_X1 U714 ( .A(KEYINPUT33), .ZN(n623) );
  INV_X1 U715 ( .A(KEYINPUT35), .ZN(n626) );
  INV_X1 U716 ( .A(KEYINPUT44), .ZN(n630) );
  AND2_X1 U717 ( .A1(n633), .A2(n632), .ZN(n634) );
  NAND2_X1 U718 ( .A1(KEYINPUT2), .A2(KEYINPUT66), .ZN(n640) );
  INV_X1 U719 ( .A(KEYINPUT2), .ZN(n644) );
  NOR2_X1 U720 ( .A1(n637), .A2(n644), .ZN(n638) );
  NOR2_X1 U721 ( .A1(n638), .A2(KEYINPUT66), .ZN(n643) );
  INV_X1 U722 ( .A(n643), .ZN(n639) );
  AND2_X1 U723 ( .A1(n640), .A2(n639), .ZN(n641) );
  XNOR2_X1 U724 ( .A(KEYINPUT89), .B(KEYINPUT124), .ZN(n645) );
  XNOR2_X1 U725 ( .A(n645), .B(KEYINPUT59), .ZN(n646) );
  NOR2_X2 U726 ( .A1(n649), .A2(n718), .ZN(n651) );
  XOR2_X1 U727 ( .A(KEYINPUT67), .B(KEYINPUT60), .Z(n650) );
  XNOR2_X1 U728 ( .A(n651), .B(n650), .ZN(G60) );
  INV_X1 U729 ( .A(KEYINPUT85), .ZN(n653) );
  NOR2_X1 U730 ( .A1(n653), .A2(KEYINPUT2), .ZN(n654) );
  NAND2_X1 U731 ( .A1(n658), .A2(n657), .ZN(n659) );
  OR2_X1 U732 ( .A1(n662), .A2(n661), .ZN(n663) );
  XNOR2_X1 U733 ( .A(n663), .B(KEYINPUT49), .ZN(n664) );
  XNOR2_X1 U734 ( .A(n664), .B(KEYINPUT114), .ZN(n665) );
  NAND2_X1 U735 ( .A1(n667), .A2(n666), .ZN(n668) );
  NOR2_X1 U736 ( .A1(n670), .A2(n669), .ZN(n671) );
  NOR2_X1 U737 ( .A1(n672), .A2(n671), .ZN(n676) );
  NOR2_X1 U738 ( .A1(n674), .A2(n673), .ZN(n675) );
  NOR2_X1 U739 ( .A1(n676), .A2(n675), .ZN(n678) );
  NOR2_X1 U740 ( .A1(n678), .A2(n677), .ZN(n679) );
  NOR2_X1 U741 ( .A1(n680), .A2(n679), .ZN(n681) );
  XOR2_X1 U742 ( .A(KEYINPUT120), .B(KEYINPUT53), .Z(n684) );
  XNOR2_X1 U743 ( .A(n685), .B(n684), .ZN(G75) );
  XNOR2_X1 U744 ( .A(n686), .B(n687), .ZN(G12) );
  NAND2_X1 U745 ( .A1(n710), .A2(G472), .ZN(n691) );
  XOR2_X1 U746 ( .A(KEYINPUT88), .B(KEYINPUT62), .Z(n689) );
  XNOR2_X1 U747 ( .A(n688), .B(n689), .ZN(n690) );
  XNOR2_X1 U748 ( .A(n691), .B(n690), .ZN(n692) );
  NOR2_X2 U749 ( .A1(n692), .A2(n718), .ZN(n694) );
  XOR2_X1 U750 ( .A(KEYINPUT112), .B(KEYINPUT63), .Z(n693) );
  XNOR2_X1 U751 ( .A(n694), .B(n693), .ZN(G57) );
  XOR2_X1 U752 ( .A(KEYINPUT54), .B(KEYINPUT55), .Z(n695) );
  XNOR2_X1 U753 ( .A(n696), .B(n695), .ZN(n697) );
  XNOR2_X1 U754 ( .A(n698), .B(n697), .ZN(n699) );
  NOR2_X2 U755 ( .A1(n699), .A2(n718), .ZN(n700) );
  XNOR2_X1 U756 ( .A(n700), .B(KEYINPUT56), .ZN(G51) );
  XOR2_X1 U757 ( .A(G122), .B(KEYINPUT127), .Z(n701) );
  XNOR2_X1 U758 ( .A(n702), .B(n701), .ZN(G24) );
  NAND2_X1 U759 ( .A1(n710), .A2(G217), .ZN(n703) );
  XOR2_X1 U760 ( .A(n704), .B(n703), .Z(n705) );
  NOR2_X1 U761 ( .A1(n705), .A2(n718), .ZN(G66) );
  NAND2_X1 U762 ( .A1(n710), .A2(G478), .ZN(n708) );
  XNOR2_X1 U763 ( .A(n706), .B(KEYINPUT125), .ZN(n707) );
  XNOR2_X1 U764 ( .A(n708), .B(n707), .ZN(n709) );
  NOR2_X1 U765 ( .A1(n709), .A2(n718), .ZN(G63) );
  NAND2_X1 U766 ( .A1(n710), .A2(G469), .ZN(n717) );
  XNOR2_X1 U767 ( .A(KEYINPUT122), .B(KEYINPUT123), .ZN(n712) );
  XNOR2_X1 U768 ( .A(n712), .B(KEYINPUT121), .ZN(n714) );
  XOR2_X1 U769 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n713) );
  XNOR2_X1 U770 ( .A(n714), .B(n713), .ZN(n715) );
  XNOR2_X1 U771 ( .A(n711), .B(n715), .ZN(n716) );
  XNOR2_X1 U772 ( .A(n717), .B(n716), .ZN(n719) );
  NOR2_X1 U773 ( .A1(n719), .A2(n718), .ZN(G54) );
  XOR2_X1 U774 ( .A(KEYINPUT27), .B(KEYINPUT26), .Z(n723) );
  NOR2_X1 U775 ( .A1(n721), .A2(n720), .ZN(n722) );
  XOR2_X1 U776 ( .A(n723), .B(n722), .Z(n724) );
  XNOR2_X1 U777 ( .A(G107), .B(n724), .ZN(G9) );
  XOR2_X1 U778 ( .A(G128), .B(KEYINPUT29), .Z(n728) );
  NAND2_X1 U779 ( .A1(n725), .A2(n726), .ZN(n727) );
  XNOR2_X1 U780 ( .A(n728), .B(n727), .ZN(G30) );
  NAND2_X1 U781 ( .A1(n725), .A2(n729), .ZN(n730) );
  XNOR2_X1 U782 ( .A(n730), .B(G146), .ZN(G48) );
  XOR2_X1 U783 ( .A(G125), .B(n731), .Z(n732) );
  XNOR2_X1 U784 ( .A(n732), .B(KEYINPUT37), .ZN(G27) );
  XNOR2_X1 U785 ( .A(G134), .B(n733), .ZN(G36) );
  NAND2_X1 U786 ( .A1(n734), .A2(n748), .ZN(n738) );
  NAND2_X1 U787 ( .A1(G953), .A2(G224), .ZN(n735) );
  XNOR2_X1 U788 ( .A(KEYINPUT61), .B(n735), .ZN(n736) );
  NAND2_X1 U789 ( .A1(n736), .A2(G898), .ZN(n737) );
  NAND2_X1 U790 ( .A1(n738), .A2(n737), .ZN(n744) );
  XOR2_X1 U791 ( .A(KEYINPUT126), .B(n740), .Z(n742) );
  NOR2_X1 U792 ( .A1(n742), .A2(n741), .ZN(n743) );
  XNOR2_X1 U793 ( .A(n744), .B(n743), .ZN(G69) );
  XOR2_X1 U794 ( .A(n746), .B(n745), .Z(n750) );
  XNOR2_X1 U795 ( .A(n747), .B(n750), .ZN(n749) );
  NAND2_X1 U796 ( .A1(n749), .A2(n748), .ZN(n754) );
  XOR2_X1 U797 ( .A(G227), .B(n750), .Z(n751) );
  NAND2_X1 U798 ( .A1(n751), .A2(G900), .ZN(n752) );
  NAND2_X1 U799 ( .A1(n752), .A2(G953), .ZN(n753) );
  NAND2_X1 U800 ( .A1(n754), .A2(n753), .ZN(G72) );
  XNOR2_X1 U801 ( .A(G140), .B(KEYINPUT113), .ZN(n756) );
  XNOR2_X1 U802 ( .A(n756), .B(n755), .ZN(G42) );
  XOR2_X1 U803 ( .A(n352), .B(G131), .Z(G33) );
  XOR2_X1 U804 ( .A(G137), .B(n758), .Z(G39) );
endmodule

