

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n295, n296, n297, n298, n299, n300, n301, n302, n303, n304, n305,
         n306, n307, n308, n309, n310, n311, n312, n313, n314, n315, n316,
         n317, n318, n319, n320, n321, n322, n323, n324, n325, n326, n327,
         n328, n329, n330, n331, n332, n333, n334, n335, n336, n337, n338,
         n339, n340, n341, n342, n343, n344, n345, n346, n347, n348, n349,
         n350, n351, n352, n353, n354, n355, n356, n357, n358, n359, n360,
         n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, n371,
         n372, n373, n374, n375, n376, n377, n378, n379, n380, n381, n382,
         n383, n384, n385, n386, n387, n388, n389, n390, n391, n392, n393,
         n394, n395, n396, n397, n398, n399, n400, n401, n402, n403, n404,
         n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, n415,
         n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426,
         n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437,
         n438, n439, n440, n441, n442, n443, n444, n445, n446, n447, n448,
         n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, n459,
         n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, n470,
         n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481,
         n482, n483, n484, n485, n486, n487, n488, n489, n490, n491, n492,
         n493, n494, n495, n496, n497, n498, n499, n500, n501, n502, n503,
         n504, n505, n506, n507, n508, n509, n510, n511, n512, n513, n514,
         n515, n516, n517, n518, n519, n520, n521, n522, n523, n524, n525,
         n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536,
         n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547,
         n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558,
         n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569,
         n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580,
         n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591,
         n592;

  XNOR2_X1 U327 ( .A(KEYINPUT64), .B(KEYINPUT48), .ZN(n477) );
  XNOR2_X1 U328 ( .A(n423), .B(n422), .ZN(n530) );
  XNOR2_X1 U329 ( .A(G29GAT), .B(KEYINPUT72), .ZN(n321) );
  XNOR2_X1 U330 ( .A(n322), .B(n321), .ZN(n324) );
  INV_X1 U331 ( .A(KEYINPUT37), .ZN(n421) );
  XNOR2_X1 U332 ( .A(n421), .B(KEYINPUT105), .ZN(n422) );
  XNOR2_X1 U333 ( .A(n330), .B(n329), .ZN(n331) );
  XNOR2_X1 U334 ( .A(n304), .B(n303), .ZN(n305) );
  XNOR2_X1 U335 ( .A(n332), .B(n331), .ZN(n333) );
  XNOR2_X1 U336 ( .A(n478), .B(n477), .ZN(n560) );
  XNOR2_X1 U337 ( .A(n306), .B(n305), .ZN(n310) );
  NOR2_X1 U338 ( .A1(n486), .A2(n485), .ZN(n574) );
  INV_X1 U339 ( .A(G43GAT), .ZN(n460) );
  XNOR2_X1 U340 ( .A(n491), .B(n490), .ZN(n492) );
  XNOR2_X1 U341 ( .A(n460), .B(KEYINPUT40), .ZN(n461) );
  XNOR2_X1 U342 ( .A(n493), .B(n492), .ZN(G1351GAT) );
  XNOR2_X1 U343 ( .A(n462), .B(n461), .ZN(G1330GAT) );
  XOR2_X1 U344 ( .A(G190GAT), .B(G134GAT), .Z(n296) );
  XOR2_X1 U345 ( .A(G15GAT), .B(G127GAT), .Z(n341) );
  XOR2_X1 U346 ( .A(G113GAT), .B(KEYINPUT0), .Z(n410) );
  XNOR2_X1 U347 ( .A(n341), .B(n410), .ZN(n295) );
  XNOR2_X1 U348 ( .A(n296), .B(n295), .ZN(n297) );
  XOR2_X1 U349 ( .A(G120GAT), .B(G71GAT), .Z(n453) );
  XOR2_X1 U350 ( .A(n297), .B(n453), .Z(n306) );
  XOR2_X1 U351 ( .A(G176GAT), .B(KEYINPUT20), .Z(n299) );
  NAND2_X1 U352 ( .A1(G227GAT), .A2(G233GAT), .ZN(n298) );
  XNOR2_X1 U353 ( .A(n299), .B(n298), .ZN(n300) );
  XNOR2_X1 U354 ( .A(G169GAT), .B(n300), .ZN(n304) );
  XOR2_X1 U355 ( .A(KEYINPUT90), .B(KEYINPUT91), .Z(n302) );
  XNOR2_X1 U356 ( .A(G43GAT), .B(G99GAT), .ZN(n301) );
  XNOR2_X1 U357 ( .A(n302), .B(n301), .ZN(n303) );
  XOR2_X1 U358 ( .A(KEYINPUT89), .B(KEYINPUT17), .Z(n308) );
  XNOR2_X1 U359 ( .A(KEYINPUT18), .B(G183GAT), .ZN(n307) );
  XNOR2_X1 U360 ( .A(n308), .B(n307), .ZN(n309) );
  XOR2_X1 U361 ( .A(KEYINPUT19), .B(n309), .Z(n382) );
  XOR2_X1 U362 ( .A(n310), .B(n382), .Z(n486) );
  XNOR2_X1 U363 ( .A(G50GAT), .B(KEYINPUT79), .ZN(n311) );
  XNOR2_X1 U364 ( .A(n311), .B(G162GAT), .ZN(n360) );
  XNOR2_X1 U365 ( .A(G99GAT), .B(G85GAT), .ZN(n312) );
  XNOR2_X1 U366 ( .A(n312), .B(KEYINPUT75), .ZN(n443) );
  XNOR2_X1 U367 ( .A(n360), .B(n443), .ZN(n334) );
  XOR2_X1 U368 ( .A(KEYINPUT82), .B(KEYINPUT10), .Z(n314) );
  XNOR2_X1 U369 ( .A(KEYINPUT67), .B(KEYINPUT9), .ZN(n313) );
  XNOR2_X1 U370 ( .A(n314), .B(n313), .ZN(n316) );
  INV_X1 U371 ( .A(G92GAT), .ZN(n315) );
  XNOR2_X1 U372 ( .A(n316), .B(n315), .ZN(n318) );
  NAND2_X1 U373 ( .A1(G232GAT), .A2(G233GAT), .ZN(n317) );
  XNOR2_X1 U374 ( .A(n318), .B(n317), .ZN(n320) );
  INV_X1 U375 ( .A(KEYINPUT80), .ZN(n319) );
  XNOR2_X1 U376 ( .A(n320), .B(n319), .ZN(n326) );
  XNOR2_X1 U377 ( .A(G43GAT), .B(KEYINPUT7), .ZN(n322) );
  XOR2_X1 U378 ( .A(KEYINPUT71), .B(KEYINPUT8), .Z(n323) );
  XNOR2_X1 U379 ( .A(n324), .B(n323), .ZN(n438) );
  XNOR2_X1 U380 ( .A(n438), .B(G106GAT), .ZN(n325) );
  XNOR2_X1 U381 ( .A(n326), .B(n325), .ZN(n332) );
  XOR2_X1 U382 ( .A(KEYINPUT84), .B(KEYINPUT11), .Z(n328) );
  XOR2_X1 U383 ( .A(G134GAT), .B(KEYINPUT83), .Z(n407) );
  XOR2_X1 U384 ( .A(G36GAT), .B(G190GAT), .Z(n380) );
  XNOR2_X1 U385 ( .A(n407), .B(n380), .ZN(n327) );
  XOR2_X1 U386 ( .A(n328), .B(n327), .Z(n330) );
  XNOR2_X1 U387 ( .A(G218GAT), .B(KEYINPUT81), .ZN(n329) );
  XNOR2_X1 U388 ( .A(n334), .B(n333), .ZN(n569) );
  XOR2_X1 U389 ( .A(KEYINPUT36), .B(KEYINPUT104), .Z(n335) );
  XNOR2_X1 U390 ( .A(n569), .B(n335), .ZN(n590) );
  XOR2_X1 U391 ( .A(KEYINPUT87), .B(KEYINPUT15), .Z(n337) );
  XNOR2_X1 U392 ( .A(KEYINPUT12), .B(KEYINPUT86), .ZN(n336) );
  XNOR2_X1 U393 ( .A(n337), .B(n336), .ZN(n353) );
  XOR2_X1 U394 ( .A(G22GAT), .B(G155GAT), .Z(n357) );
  XOR2_X1 U395 ( .A(n357), .B(KEYINPUT14), .Z(n339) );
  NAND2_X1 U396 ( .A1(G231GAT), .A2(G233GAT), .ZN(n338) );
  XNOR2_X1 U397 ( .A(n339), .B(n338), .ZN(n340) );
  XNOR2_X1 U398 ( .A(n341), .B(n340), .ZN(n351) );
  XOR2_X1 U399 ( .A(G78GAT), .B(G211GAT), .Z(n343) );
  XNOR2_X1 U400 ( .A(G183GAT), .B(G71GAT), .ZN(n342) );
  XNOR2_X1 U401 ( .A(n343), .B(n342), .ZN(n347) );
  XOR2_X1 U402 ( .A(KEYINPUT85), .B(KEYINPUT88), .Z(n345) );
  XNOR2_X1 U403 ( .A(G8GAT), .B(G64GAT), .ZN(n344) );
  XNOR2_X1 U404 ( .A(n345), .B(n344), .ZN(n346) );
  XOR2_X1 U405 ( .A(n347), .B(n346), .Z(n349) );
  XOR2_X1 U406 ( .A(KEYINPUT73), .B(G1GAT), .Z(n425) );
  XOR2_X1 U407 ( .A(G57GAT), .B(KEYINPUT13), .Z(n452) );
  XNOR2_X1 U408 ( .A(n425), .B(n452), .ZN(n348) );
  XNOR2_X1 U409 ( .A(n349), .B(n348), .ZN(n350) );
  XNOR2_X1 U410 ( .A(n351), .B(n350), .ZN(n352) );
  XOR2_X1 U411 ( .A(n353), .B(n352), .Z(n586) );
  INV_X1 U412 ( .A(n586), .ZN(n494) );
  XOR2_X1 U413 ( .A(KEYINPUT94), .B(KEYINPUT93), .Z(n355) );
  XNOR2_X1 U414 ( .A(KEYINPUT92), .B(KEYINPUT24), .ZN(n354) );
  XNOR2_X1 U415 ( .A(n355), .B(n354), .ZN(n371) );
  XNOR2_X1 U416 ( .A(G106GAT), .B(G78GAT), .ZN(n356) );
  XNOR2_X1 U417 ( .A(n356), .B(G148GAT), .ZN(n444) );
  XOR2_X1 U418 ( .A(n357), .B(n444), .Z(n359) );
  XNOR2_X1 U419 ( .A(KEYINPUT23), .B(G204GAT), .ZN(n358) );
  XNOR2_X1 U420 ( .A(n359), .B(n358), .ZN(n364) );
  XOR2_X1 U421 ( .A(KEYINPUT22), .B(n360), .Z(n362) );
  NAND2_X1 U422 ( .A1(G228GAT), .A2(G233GAT), .ZN(n361) );
  XNOR2_X1 U423 ( .A(n362), .B(n361), .ZN(n363) );
  XOR2_X1 U424 ( .A(n364), .B(n363), .Z(n369) );
  XNOR2_X1 U425 ( .A(G141GAT), .B(KEYINPUT3), .ZN(n365) );
  XNOR2_X1 U426 ( .A(n365), .B(KEYINPUT2), .ZN(n409) );
  XOR2_X1 U427 ( .A(G211GAT), .B(KEYINPUT21), .Z(n367) );
  XNOR2_X1 U428 ( .A(G197GAT), .B(G218GAT), .ZN(n366) );
  XNOR2_X1 U429 ( .A(n367), .B(n366), .ZN(n377) );
  XNOR2_X1 U430 ( .A(n409), .B(n377), .ZN(n368) );
  XNOR2_X1 U431 ( .A(n369), .B(n368), .ZN(n370) );
  XNOR2_X1 U432 ( .A(n371), .B(n370), .ZN(n483) );
  INV_X1 U433 ( .A(n486), .ZN(n545) );
  XOR2_X1 U434 ( .A(KEYINPUT97), .B(KEYINPUT98), .Z(n373) );
  NAND2_X1 U435 ( .A1(G226GAT), .A2(G233GAT), .ZN(n372) );
  XNOR2_X1 U436 ( .A(n373), .B(n372), .ZN(n374) );
  XOR2_X1 U437 ( .A(n374), .B(KEYINPUT85), .Z(n379) );
  XOR2_X1 U438 ( .A(G64GAT), .B(G92GAT), .Z(n376) );
  XNOR2_X1 U439 ( .A(G176GAT), .B(G204GAT), .ZN(n375) );
  XNOR2_X1 U440 ( .A(n376), .B(n375), .ZN(n450) );
  XNOR2_X1 U441 ( .A(n377), .B(n450), .ZN(n378) );
  XNOR2_X1 U442 ( .A(n379), .B(n378), .ZN(n381) );
  XOR2_X1 U443 ( .A(n381), .B(n380), .Z(n385) );
  XOR2_X1 U444 ( .A(G169GAT), .B(G8GAT), .Z(n424) );
  INV_X1 U445 ( .A(n382), .ZN(n383) );
  XOR2_X1 U446 ( .A(n424), .B(n383), .Z(n384) );
  XOR2_X1 U447 ( .A(n385), .B(n384), .Z(n511) );
  INV_X1 U448 ( .A(n511), .ZN(n536) );
  AND2_X1 U449 ( .A1(n545), .A2(n536), .ZN(n386) );
  XNOR2_X1 U450 ( .A(KEYINPUT100), .B(n386), .ZN(n387) );
  NOR2_X1 U451 ( .A1(n483), .A2(n387), .ZN(n389) );
  XOR2_X1 U452 ( .A(KEYINPUT25), .B(KEYINPUT101), .Z(n388) );
  XNOR2_X1 U453 ( .A(n389), .B(n388), .ZN(n393) );
  NAND2_X1 U454 ( .A1(n483), .A2(n486), .ZN(n390) );
  XNOR2_X1 U455 ( .A(n390), .B(KEYINPUT26), .ZN(n576) );
  XNOR2_X1 U456 ( .A(n511), .B(KEYINPUT27), .ZN(n416) );
  NOR2_X1 U457 ( .A1(n576), .A2(n416), .ZN(n391) );
  XNOR2_X1 U458 ( .A(n391), .B(KEYINPUT99), .ZN(n392) );
  NAND2_X1 U459 ( .A1(n393), .A2(n392), .ZN(n415) );
  XOR2_X1 U460 ( .A(KEYINPUT95), .B(KEYINPUT6), .Z(n395) );
  XNOR2_X1 U461 ( .A(G57GAT), .B(KEYINPUT96), .ZN(n394) );
  XNOR2_X1 U462 ( .A(n395), .B(n394), .ZN(n414) );
  XOR2_X1 U463 ( .A(G85GAT), .B(G162GAT), .Z(n397) );
  XNOR2_X1 U464 ( .A(G29GAT), .B(G120GAT), .ZN(n396) );
  XNOR2_X1 U465 ( .A(n397), .B(n396), .ZN(n401) );
  XOR2_X1 U466 ( .A(G155GAT), .B(G148GAT), .Z(n399) );
  XNOR2_X1 U467 ( .A(G1GAT), .B(G127GAT), .ZN(n398) );
  XNOR2_X1 U468 ( .A(n399), .B(n398), .ZN(n400) );
  XOR2_X1 U469 ( .A(n401), .B(n400), .Z(n406) );
  XOR2_X1 U470 ( .A(KEYINPUT4), .B(KEYINPUT1), .Z(n403) );
  NAND2_X1 U471 ( .A1(G225GAT), .A2(G233GAT), .ZN(n402) );
  XNOR2_X1 U472 ( .A(n403), .B(n402), .ZN(n404) );
  XNOR2_X1 U473 ( .A(KEYINPUT5), .B(n404), .ZN(n405) );
  XNOR2_X1 U474 ( .A(n406), .B(n405), .ZN(n408) );
  XOR2_X1 U475 ( .A(n408), .B(n407), .Z(n412) );
  XNOR2_X1 U476 ( .A(n410), .B(n409), .ZN(n411) );
  XNOR2_X1 U477 ( .A(n412), .B(n411), .ZN(n413) );
  XNOR2_X1 U478 ( .A(n414), .B(n413), .ZN(n532) );
  INV_X1 U479 ( .A(n532), .ZN(n508) );
  NAND2_X1 U480 ( .A1(n415), .A2(n508), .ZN(n419) );
  OR2_X1 U481 ( .A1(n508), .A2(n416), .ZN(n559) );
  XNOR2_X1 U482 ( .A(KEYINPUT28), .B(KEYINPUT68), .ZN(n417) );
  XOR2_X1 U483 ( .A(n417), .B(n483), .Z(n514) );
  INV_X1 U484 ( .A(n514), .ZN(n540) );
  NOR2_X1 U485 ( .A1(n559), .A2(n540), .ZN(n544) );
  NAND2_X1 U486 ( .A1(n544), .A2(n486), .ZN(n418) );
  NAND2_X1 U487 ( .A1(n419), .A2(n418), .ZN(n496) );
  NAND2_X1 U488 ( .A1(n494), .A2(n496), .ZN(n420) );
  NOR2_X1 U489 ( .A1(n590), .A2(n420), .ZN(n423) );
  XOR2_X1 U490 ( .A(G113GAT), .B(G15GAT), .Z(n427) );
  XNOR2_X1 U491 ( .A(n425), .B(n424), .ZN(n426) );
  XNOR2_X1 U492 ( .A(n427), .B(n426), .ZN(n428) );
  XOR2_X1 U493 ( .A(n428), .B(G36GAT), .Z(n433) );
  XOR2_X1 U494 ( .A(KEYINPUT70), .B(G22GAT), .Z(n430) );
  XNOR2_X1 U495 ( .A(G141GAT), .B(G197GAT), .ZN(n429) );
  XNOR2_X1 U496 ( .A(n430), .B(n429), .ZN(n431) );
  XNOR2_X1 U497 ( .A(n431), .B(G50GAT), .ZN(n432) );
  XNOR2_X1 U498 ( .A(n433), .B(n432), .ZN(n437) );
  XOR2_X1 U499 ( .A(KEYINPUT69), .B(KEYINPUT30), .Z(n435) );
  NAND2_X1 U500 ( .A1(G229GAT), .A2(G233GAT), .ZN(n434) );
  XNOR2_X1 U501 ( .A(n435), .B(n434), .ZN(n436) );
  XNOR2_X1 U502 ( .A(n437), .B(n436), .ZN(n440) );
  XOR2_X1 U503 ( .A(n438), .B(KEYINPUT29), .Z(n439) );
  XOR2_X1 U504 ( .A(n440), .B(n439), .Z(n517) );
  INV_X1 U505 ( .A(n517), .ZN(n578) );
  XOR2_X1 U506 ( .A(KEYINPUT76), .B(KEYINPUT74), .Z(n442) );
  XNOR2_X1 U507 ( .A(KEYINPUT78), .B(KEYINPUT31), .ZN(n441) );
  XNOR2_X1 U508 ( .A(n442), .B(n441), .ZN(n457) );
  XNOR2_X1 U509 ( .A(n444), .B(n443), .ZN(n449) );
  XNOR2_X1 U510 ( .A(KEYINPUT77), .B(KEYINPUT33), .ZN(n446) );
  AND2_X1 U511 ( .A1(G230GAT), .A2(G233GAT), .ZN(n445) );
  XNOR2_X1 U512 ( .A(n446), .B(n445), .ZN(n447) );
  XOR2_X1 U513 ( .A(KEYINPUT32), .B(n447), .Z(n448) );
  XNOR2_X1 U514 ( .A(n449), .B(n448), .ZN(n451) );
  XOR2_X1 U515 ( .A(n451), .B(n450), .Z(n455) );
  XNOR2_X1 U516 ( .A(n453), .B(n452), .ZN(n454) );
  XNOR2_X1 U517 ( .A(n455), .B(n454), .ZN(n456) );
  XNOR2_X1 U518 ( .A(n457), .B(n456), .ZN(n583) );
  NAND2_X1 U519 ( .A1(n578), .A2(n583), .ZN(n498) );
  NOR2_X1 U520 ( .A1(n530), .A2(n498), .ZN(n458) );
  XOR2_X1 U521 ( .A(KEYINPUT106), .B(n458), .Z(n459) );
  XNOR2_X1 U522 ( .A(KEYINPUT38), .B(n459), .ZN(n513) );
  NOR2_X1 U523 ( .A1(n486), .A2(n513), .ZN(n462) );
  XOR2_X1 U524 ( .A(KEYINPUT65), .B(KEYINPUT41), .Z(n463) );
  XNOR2_X1 U525 ( .A(n583), .B(n463), .ZN(n563) );
  XOR2_X1 U526 ( .A(n563), .B(KEYINPUT109), .Z(n548) );
  NAND2_X1 U527 ( .A1(n578), .A2(n563), .ZN(n466) );
  XOR2_X1 U528 ( .A(KEYINPUT46), .B(KEYINPUT117), .Z(n464) );
  XNOR2_X1 U529 ( .A(KEYINPUT116), .B(n464), .ZN(n465) );
  XNOR2_X1 U530 ( .A(n466), .B(n465), .ZN(n468) );
  NOR2_X1 U531 ( .A1(n569), .A2(n586), .ZN(n467) );
  AND2_X1 U532 ( .A1(n468), .A2(n467), .ZN(n470) );
  XNOR2_X1 U533 ( .A(KEYINPUT118), .B(KEYINPUT119), .ZN(n469) );
  XNOR2_X1 U534 ( .A(n470), .B(n469), .ZN(n471) );
  XNOR2_X1 U535 ( .A(n471), .B(KEYINPUT47), .ZN(n476) );
  NOR2_X1 U536 ( .A1(n590), .A2(n494), .ZN(n472) );
  XNOR2_X1 U537 ( .A(n472), .B(KEYINPUT45), .ZN(n473) );
  NAND2_X1 U538 ( .A1(n473), .A2(n583), .ZN(n474) );
  NOR2_X1 U539 ( .A1(n474), .A2(n578), .ZN(n475) );
  NOR2_X1 U540 ( .A1(n476), .A2(n475), .ZN(n478) );
  XOR2_X1 U541 ( .A(n511), .B(KEYINPUT125), .Z(n479) );
  NOR2_X1 U542 ( .A1(n560), .A2(n479), .ZN(n480) );
  XNOR2_X1 U543 ( .A(n480), .B(KEYINPUT54), .ZN(n481) );
  NAND2_X1 U544 ( .A1(n481), .A2(n508), .ZN(n482) );
  XNOR2_X1 U545 ( .A(n482), .B(KEYINPUT66), .ZN(n577) );
  NOR2_X1 U546 ( .A1(n577), .A2(n483), .ZN(n484) );
  XNOR2_X1 U547 ( .A(n484), .B(KEYINPUT55), .ZN(n485) );
  NAND2_X1 U548 ( .A1(n548), .A2(n574), .ZN(n489) );
  XOR2_X1 U549 ( .A(KEYINPUT56), .B(KEYINPUT57), .Z(n487) );
  XNOR2_X1 U550 ( .A(n487), .B(G176GAT), .ZN(n488) );
  XNOR2_X1 U551 ( .A(n489), .B(n488), .ZN(G1349GAT) );
  NAND2_X1 U552 ( .A1(n574), .A2(n569), .ZN(n493) );
  XOR2_X1 U553 ( .A(KEYINPUT58), .B(KEYINPUT126), .Z(n491) );
  INV_X1 U554 ( .A(G190GAT), .ZN(n490) );
  XOR2_X1 U555 ( .A(KEYINPUT102), .B(KEYINPUT34), .Z(n500) );
  NOR2_X1 U556 ( .A1(n569), .A2(n494), .ZN(n495) );
  XNOR2_X1 U557 ( .A(n495), .B(KEYINPUT16), .ZN(n497) );
  NAND2_X1 U558 ( .A1(n497), .A2(n496), .ZN(n519) );
  NOR2_X1 U559 ( .A1(n498), .A2(n519), .ZN(n506) );
  NAND2_X1 U560 ( .A1(n506), .A2(n532), .ZN(n499) );
  XNOR2_X1 U561 ( .A(n500), .B(n499), .ZN(n501) );
  XOR2_X1 U562 ( .A(G1GAT), .B(n501), .Z(G1324GAT) );
  XOR2_X1 U563 ( .A(G8GAT), .B(KEYINPUT103), .Z(n503) );
  NAND2_X1 U564 ( .A1(n506), .A2(n536), .ZN(n502) );
  XNOR2_X1 U565 ( .A(n503), .B(n502), .ZN(G1325GAT) );
  XOR2_X1 U566 ( .A(G15GAT), .B(KEYINPUT35), .Z(n505) );
  NAND2_X1 U567 ( .A1(n506), .A2(n545), .ZN(n504) );
  XNOR2_X1 U568 ( .A(n505), .B(n504), .ZN(G1326GAT) );
  NAND2_X1 U569 ( .A1(n540), .A2(n506), .ZN(n507) );
  XNOR2_X1 U570 ( .A(n507), .B(G22GAT), .ZN(G1327GAT) );
  NOR2_X1 U571 ( .A1(n508), .A2(n513), .ZN(n509) );
  XNOR2_X1 U572 ( .A(n509), .B(KEYINPUT39), .ZN(n510) );
  XNOR2_X1 U573 ( .A(G29GAT), .B(n510), .ZN(G1328GAT) );
  NOR2_X1 U574 ( .A1(n511), .A2(n513), .ZN(n512) );
  XOR2_X1 U575 ( .A(G36GAT), .B(n512), .Z(G1329GAT) );
  NOR2_X1 U576 ( .A1(n514), .A2(n513), .ZN(n516) );
  XNOR2_X1 U577 ( .A(G50GAT), .B(KEYINPUT107), .ZN(n515) );
  XNOR2_X1 U578 ( .A(n516), .B(n515), .ZN(G1331GAT) );
  XOR2_X1 U579 ( .A(KEYINPUT108), .B(KEYINPUT42), .Z(n521) );
  NAND2_X1 U580 ( .A1(n517), .A2(n548), .ZN(n518) );
  XNOR2_X1 U581 ( .A(n518), .B(KEYINPUT110), .ZN(n529) );
  NOR2_X1 U582 ( .A1(n529), .A2(n519), .ZN(n525) );
  NAND2_X1 U583 ( .A1(n525), .A2(n532), .ZN(n520) );
  XNOR2_X1 U584 ( .A(n521), .B(n520), .ZN(n522) );
  XOR2_X1 U585 ( .A(G57GAT), .B(n522), .Z(G1332GAT) );
  NAND2_X1 U586 ( .A1(n525), .A2(n536), .ZN(n523) );
  XNOR2_X1 U587 ( .A(n523), .B(G64GAT), .ZN(G1333GAT) );
  NAND2_X1 U588 ( .A1(n525), .A2(n545), .ZN(n524) );
  XNOR2_X1 U589 ( .A(n524), .B(G71GAT), .ZN(G1334GAT) );
  XOR2_X1 U590 ( .A(KEYINPUT111), .B(KEYINPUT43), .Z(n527) );
  NAND2_X1 U591 ( .A1(n525), .A2(n540), .ZN(n526) );
  XNOR2_X1 U592 ( .A(n527), .B(n526), .ZN(n528) );
  XOR2_X1 U593 ( .A(G78GAT), .B(n528), .Z(G1335GAT) );
  XOR2_X1 U594 ( .A(KEYINPUT113), .B(KEYINPUT114), .Z(n534) );
  NOR2_X1 U595 ( .A1(n530), .A2(n529), .ZN(n531) );
  XNOR2_X1 U596 ( .A(n531), .B(KEYINPUT112), .ZN(n541) );
  NAND2_X1 U597 ( .A1(n541), .A2(n532), .ZN(n533) );
  XNOR2_X1 U598 ( .A(n534), .B(n533), .ZN(n535) );
  XNOR2_X1 U599 ( .A(G85GAT), .B(n535), .ZN(G1336GAT) );
  NAND2_X1 U600 ( .A1(n541), .A2(n536), .ZN(n537) );
  XNOR2_X1 U601 ( .A(n537), .B(G92GAT), .ZN(G1337GAT) );
  XOR2_X1 U602 ( .A(G99GAT), .B(KEYINPUT115), .Z(n539) );
  NAND2_X1 U603 ( .A1(n545), .A2(n541), .ZN(n538) );
  XNOR2_X1 U604 ( .A(n539), .B(n538), .ZN(G1338GAT) );
  NAND2_X1 U605 ( .A1(n541), .A2(n540), .ZN(n542) );
  XNOR2_X1 U606 ( .A(n542), .B(KEYINPUT44), .ZN(n543) );
  XNOR2_X1 U607 ( .A(G106GAT), .B(n543), .ZN(G1339GAT) );
  NAND2_X1 U608 ( .A1(n545), .A2(n544), .ZN(n546) );
  NOR2_X1 U609 ( .A1(n560), .A2(n546), .ZN(n556) );
  NAND2_X1 U610 ( .A1(n556), .A2(n578), .ZN(n547) );
  XNOR2_X1 U611 ( .A(n547), .B(G113GAT), .ZN(G1340GAT) );
  XOR2_X1 U612 ( .A(KEYINPUT120), .B(KEYINPUT49), .Z(n550) );
  NAND2_X1 U613 ( .A1(n556), .A2(n548), .ZN(n549) );
  XNOR2_X1 U614 ( .A(n550), .B(n549), .ZN(n551) );
  XNOR2_X1 U615 ( .A(G120GAT), .B(n551), .ZN(G1341GAT) );
  XNOR2_X1 U616 ( .A(G127GAT), .B(KEYINPUT122), .ZN(n555) );
  XOR2_X1 U617 ( .A(KEYINPUT50), .B(KEYINPUT121), .Z(n553) );
  NAND2_X1 U618 ( .A1(n556), .A2(n586), .ZN(n552) );
  XNOR2_X1 U619 ( .A(n553), .B(n552), .ZN(n554) );
  XNOR2_X1 U620 ( .A(n555), .B(n554), .ZN(G1342GAT) );
  XOR2_X1 U621 ( .A(G134GAT), .B(KEYINPUT51), .Z(n558) );
  NAND2_X1 U622 ( .A1(n556), .A2(n569), .ZN(n557) );
  XNOR2_X1 U623 ( .A(n558), .B(n557), .ZN(G1343GAT) );
  OR2_X1 U624 ( .A1(n576), .A2(n559), .ZN(n561) );
  NOR2_X1 U625 ( .A1(n561), .A2(n560), .ZN(n570) );
  AND2_X1 U626 ( .A1(n578), .A2(n570), .ZN(n562) );
  XOR2_X1 U627 ( .A(G141GAT), .B(n562), .Z(G1344GAT) );
  XOR2_X1 U628 ( .A(G148GAT), .B(KEYINPUT123), .Z(n565) );
  NAND2_X1 U629 ( .A1(n570), .A2(n563), .ZN(n564) );
  XNOR2_X1 U630 ( .A(n565), .B(n564), .ZN(n567) );
  XOR2_X1 U631 ( .A(KEYINPUT53), .B(KEYINPUT52), .Z(n566) );
  XNOR2_X1 U632 ( .A(n567), .B(n566), .ZN(G1345GAT) );
  NAND2_X1 U633 ( .A1(n570), .A2(n586), .ZN(n568) );
  XNOR2_X1 U634 ( .A(n568), .B(G155GAT), .ZN(G1346GAT) );
  NAND2_X1 U635 ( .A1(n570), .A2(n569), .ZN(n571) );
  XNOR2_X1 U636 ( .A(n571), .B(KEYINPUT124), .ZN(n572) );
  XNOR2_X1 U637 ( .A(G162GAT), .B(n572), .ZN(G1347GAT) );
  NAND2_X1 U638 ( .A1(n574), .A2(n578), .ZN(n573) );
  XNOR2_X1 U639 ( .A(n573), .B(G169GAT), .ZN(G1348GAT) );
  NAND2_X1 U640 ( .A1(n574), .A2(n586), .ZN(n575) );
  XNOR2_X1 U641 ( .A(n575), .B(G183GAT), .ZN(G1350GAT) );
  XOR2_X1 U642 ( .A(G197GAT), .B(KEYINPUT127), .Z(n580) );
  NOR2_X1 U643 ( .A1(n577), .A2(n576), .ZN(n587) );
  NAND2_X1 U644 ( .A1(n587), .A2(n578), .ZN(n579) );
  XNOR2_X1 U645 ( .A(n580), .B(n579), .ZN(n582) );
  XOR2_X1 U646 ( .A(KEYINPUT60), .B(KEYINPUT59), .Z(n581) );
  XNOR2_X1 U647 ( .A(n582), .B(n581), .ZN(G1352GAT) );
  XOR2_X1 U648 ( .A(G204GAT), .B(KEYINPUT61), .Z(n585) );
  INV_X1 U649 ( .A(n587), .ZN(n589) );
  OR2_X1 U650 ( .A1(n589), .A2(n583), .ZN(n584) );
  XNOR2_X1 U651 ( .A(n585), .B(n584), .ZN(G1353GAT) );
  NAND2_X1 U652 ( .A1(n587), .A2(n586), .ZN(n588) );
  XNOR2_X1 U653 ( .A(n588), .B(G211GAT), .ZN(G1354GAT) );
  NOR2_X1 U654 ( .A1(n590), .A2(n589), .ZN(n591) );
  XOR2_X1 U655 ( .A(KEYINPUT62), .B(n591), .Z(n592) );
  XNOR2_X1 U656 ( .A(G218GAT), .B(n592), .ZN(G1355GAT) );
endmodule

