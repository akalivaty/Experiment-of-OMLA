//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 0 1 1 1 1 1 0 1 1 1 0 0 1 0 1 1 1 0 0 1 0 0 1 1 0 0 0 1 0 0 1 1 1 1 0 0 0 0 1 0 1 1 0 1 0 1 0 1 1 0 1 0 1 1 0 0 1 1 1 0 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:25:26 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n614, new_n615,
    new_n616, new_n617, new_n619, new_n620, new_n621, new_n622, new_n623,
    new_n624, new_n625, new_n626, new_n627, new_n628, new_n629, new_n631,
    new_n632, new_n633, new_n634, new_n635, new_n636, new_n637, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n677,
    new_n678, new_n680, new_n681, new_n682, new_n683, new_n684, new_n685,
    new_n686, new_n687, new_n689, new_n690, new_n691, new_n692, new_n693,
    new_n694, new_n695, new_n696, new_n697, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n728, new_n729, new_n730, new_n731,
    new_n732, new_n733, new_n734, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n887, new_n888, new_n890, new_n891, new_n892,
    new_n893, new_n894, new_n895, new_n896, new_n897, new_n898, new_n899,
    new_n900, new_n901, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n931, new_n932, new_n933, new_n934, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n956, new_n957, new_n958, new_n959,
    new_n960, new_n961, new_n962, new_n963, new_n964;
  INV_X1    g000(.A(G469), .ZN(new_n187));
  INV_X1    g001(.A(G902), .ZN(new_n188));
  XNOR2_X1  g002(.A(G110), .B(G140), .ZN(new_n189));
  INV_X1    g003(.A(G953), .ZN(new_n190));
  AND2_X1   g004(.A1(new_n190), .A2(G227), .ZN(new_n191));
  XOR2_X1   g005(.A(new_n189), .B(new_n191), .Z(new_n192));
  INV_X1    g006(.A(KEYINPUT10), .ZN(new_n193));
  INV_X1    g007(.A(G146), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n194), .A2(KEYINPUT64), .ZN(new_n195));
  INV_X1    g009(.A(KEYINPUT64), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n196), .A2(G146), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n195), .A2(new_n197), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n198), .A2(G143), .ZN(new_n199));
  INV_X1    g013(.A(KEYINPUT1), .ZN(new_n200));
  NOR2_X1   g014(.A1(new_n194), .A2(G143), .ZN(new_n201));
  INV_X1    g015(.A(new_n201), .ZN(new_n202));
  NAND4_X1  g016(.A1(new_n199), .A2(new_n200), .A3(G128), .A4(new_n202), .ZN(new_n203));
  INV_X1    g017(.A(G143), .ZN(new_n204));
  NOR2_X1   g018(.A1(new_n204), .A2(G146), .ZN(new_n205));
  OAI21_X1  g019(.A(G128), .B1(new_n205), .B2(new_n200), .ZN(new_n206));
  AOI21_X1  g020(.A(new_n204), .B1(new_n195), .B2(new_n197), .ZN(new_n207));
  OAI21_X1  g021(.A(new_n206), .B1(new_n207), .B2(new_n201), .ZN(new_n208));
  AND2_X1   g022(.A1(new_n203), .A2(new_n208), .ZN(new_n209));
  INV_X1    g023(.A(G101), .ZN(new_n210));
  INV_X1    g024(.A(G104), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n211), .A2(G107), .ZN(new_n212));
  INV_X1    g026(.A(G107), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n213), .A2(G104), .ZN(new_n214));
  AOI21_X1  g028(.A(new_n210), .B1(new_n212), .B2(new_n214), .ZN(new_n215));
  INV_X1    g029(.A(new_n215), .ZN(new_n216));
  OAI21_X1  g030(.A(KEYINPUT3), .B1(new_n211), .B2(G107), .ZN(new_n217));
  INV_X1    g031(.A(KEYINPUT3), .ZN(new_n218));
  NAND3_X1  g032(.A1(new_n218), .A2(new_n213), .A3(G104), .ZN(new_n219));
  NAND4_X1  g033(.A1(new_n217), .A2(new_n219), .A3(new_n210), .A4(new_n212), .ZN(new_n220));
  AND2_X1   g034(.A1(new_n220), .A2(KEYINPUT81), .ZN(new_n221));
  NOR2_X1   g035(.A1(new_n220), .A2(KEYINPUT81), .ZN(new_n222));
  OAI21_X1  g036(.A(new_n216), .B1(new_n221), .B2(new_n222), .ZN(new_n223));
  OAI21_X1  g037(.A(new_n193), .B1(new_n209), .B2(new_n223), .ZN(new_n224));
  OR2_X1    g038(.A1(new_n220), .A2(KEYINPUT81), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n220), .A2(KEYINPUT81), .ZN(new_n226));
  AOI21_X1  g040(.A(new_n215), .B1(new_n225), .B2(new_n226), .ZN(new_n227));
  OAI21_X1  g041(.A(G128), .B1(new_n207), .B2(new_n200), .ZN(new_n228));
  INV_X1    g042(.A(new_n205), .ZN(new_n229));
  OAI21_X1  g043(.A(new_n229), .B1(new_n198), .B2(G143), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n228), .A2(new_n230), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n231), .A2(new_n203), .ZN(new_n232));
  NAND3_X1  g046(.A1(new_n227), .A2(new_n232), .A3(KEYINPUT10), .ZN(new_n233));
  NAND3_X1  g047(.A1(new_n217), .A2(new_n219), .A3(new_n212), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n234), .A2(G101), .ZN(new_n235));
  INV_X1    g049(.A(new_n235), .ZN(new_n236));
  XOR2_X1   g050(.A(KEYINPUT82), .B(KEYINPUT4), .Z(new_n237));
  NAND2_X1  g051(.A1(new_n236), .A2(new_n237), .ZN(new_n238));
  INV_X1    g052(.A(KEYINPUT80), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n235), .A2(new_n239), .ZN(new_n240));
  OAI21_X1  g054(.A(new_n240), .B1(new_n221), .B2(new_n222), .ZN(new_n241));
  OAI21_X1  g055(.A(KEYINPUT4), .B1(new_n235), .B2(new_n239), .ZN(new_n242));
  OAI21_X1  g056(.A(new_n238), .B1(new_n241), .B2(new_n242), .ZN(new_n243));
  AND2_X1   g057(.A1(KEYINPUT0), .A2(G128), .ZN(new_n244));
  XNOR2_X1  g058(.A(KEYINPUT64), .B(G146), .ZN(new_n245));
  OAI211_X1 g059(.A(new_n202), .B(new_n244), .C1(new_n245), .C2(new_n204), .ZN(new_n246));
  AOI21_X1  g060(.A(new_n205), .B1(new_n245), .B2(new_n204), .ZN(new_n247));
  NOR2_X1   g061(.A1(KEYINPUT0), .A2(G128), .ZN(new_n248));
  NOR2_X1   g062(.A1(new_n244), .A2(new_n248), .ZN(new_n249));
  INV_X1    g063(.A(new_n249), .ZN(new_n250));
  OAI21_X1  g064(.A(new_n246), .B1(new_n247), .B2(new_n250), .ZN(new_n251));
  NOR2_X1   g065(.A1(new_n251), .A2(KEYINPUT66), .ZN(new_n252));
  INV_X1    g066(.A(KEYINPUT66), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n230), .A2(new_n249), .ZN(new_n254));
  AOI21_X1  g068(.A(new_n253), .B1(new_n254), .B2(new_n246), .ZN(new_n255));
  NOR2_X1   g069(.A1(new_n252), .A2(new_n255), .ZN(new_n256));
  OAI211_X1 g070(.A(new_n224), .B(new_n233), .C1(new_n243), .C2(new_n256), .ZN(new_n257));
  INV_X1    g071(.A(KEYINPUT11), .ZN(new_n258));
  INV_X1    g072(.A(G134), .ZN(new_n259));
  OAI21_X1  g073(.A(new_n258), .B1(new_n259), .B2(G137), .ZN(new_n260));
  INV_X1    g074(.A(G137), .ZN(new_n261));
  NAND3_X1  g075(.A1(new_n261), .A2(KEYINPUT11), .A3(G134), .ZN(new_n262));
  INV_X1    g076(.A(G131), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n259), .A2(G137), .ZN(new_n264));
  NAND4_X1  g078(.A1(new_n260), .A2(new_n262), .A3(new_n263), .A4(new_n264), .ZN(new_n265));
  XNOR2_X1  g079(.A(new_n265), .B(KEYINPUT65), .ZN(new_n266));
  NAND3_X1  g080(.A1(new_n260), .A2(new_n264), .A3(new_n262), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n267), .A2(G131), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n266), .A2(new_n268), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n257), .A2(new_n269), .ZN(new_n270));
  INV_X1    g084(.A(KEYINPUT83), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n270), .A2(new_n271), .ZN(new_n272));
  NAND3_X1  g086(.A1(new_n257), .A2(KEYINPUT83), .A3(new_n269), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n272), .A2(new_n273), .ZN(new_n274));
  XNOR2_X1  g088(.A(new_n220), .B(KEYINPUT81), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n236), .A2(KEYINPUT80), .ZN(new_n276));
  NAND4_X1  g090(.A1(new_n275), .A2(new_n276), .A3(KEYINPUT4), .A4(new_n240), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n251), .A2(KEYINPUT66), .ZN(new_n278));
  NAND3_X1  g092(.A1(new_n254), .A2(new_n253), .A3(new_n246), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n278), .A2(new_n279), .ZN(new_n280));
  NAND3_X1  g094(.A1(new_n277), .A2(new_n280), .A3(new_n238), .ZN(new_n281));
  AND2_X1   g095(.A1(new_n266), .A2(new_n268), .ZN(new_n282));
  NAND4_X1  g096(.A1(new_n281), .A2(new_n282), .A3(new_n224), .A4(new_n233), .ZN(new_n283));
  AOI21_X1  g097(.A(new_n192), .B1(new_n274), .B2(new_n283), .ZN(new_n284));
  INV_X1    g098(.A(KEYINPUT12), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n203), .A2(new_n208), .ZN(new_n286));
  NAND2_X1  g100(.A1(new_n227), .A2(new_n286), .ZN(new_n287));
  INV_X1    g101(.A(G128), .ZN(new_n288));
  NOR3_X1   g102(.A1(new_n207), .A2(new_n288), .A3(new_n201), .ZN(new_n289));
  AOI22_X1  g103(.A1(new_n200), .A2(new_n289), .B1(new_n228), .B2(new_n230), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n290), .A2(new_n223), .ZN(new_n291));
  AOI211_X1 g105(.A(new_n285), .B(new_n282), .C1(new_n287), .C2(new_n291), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n287), .A2(new_n291), .ZN(new_n293));
  AOI21_X1  g107(.A(KEYINPUT12), .B1(new_n293), .B2(new_n269), .ZN(new_n294));
  NOR2_X1   g108(.A1(new_n292), .A2(new_n294), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n283), .A2(new_n192), .ZN(new_n296));
  NOR2_X1   g110(.A1(new_n295), .A2(new_n296), .ZN(new_n297));
  OAI211_X1 g111(.A(new_n187), .B(new_n188), .C1(new_n284), .C2(new_n297), .ZN(new_n298));
  NAND2_X1  g112(.A1(G469), .A2(G902), .ZN(new_n299));
  OR2_X1    g113(.A1(new_n292), .A2(new_n294), .ZN(new_n300));
  AOI21_X1  g114(.A(new_n192), .B1(new_n300), .B2(new_n283), .ZN(new_n301));
  AOI21_X1  g115(.A(new_n296), .B1(new_n272), .B2(new_n273), .ZN(new_n302));
  NOR2_X1   g116(.A1(new_n301), .A2(new_n302), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n303), .A2(G469), .ZN(new_n304));
  NAND3_X1  g118(.A1(new_n298), .A2(new_n299), .A3(new_n304), .ZN(new_n305));
  XOR2_X1   g119(.A(KEYINPUT9), .B(G234), .Z(new_n306));
  XNOR2_X1  g120(.A(new_n306), .B(KEYINPUT78), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n307), .A2(new_n188), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n308), .A2(G221), .ZN(new_n309));
  XOR2_X1   g123(.A(new_n309), .B(KEYINPUT79), .Z(new_n310));
  NAND2_X1  g124(.A1(new_n305), .A2(new_n310), .ZN(new_n311));
  INV_X1    g125(.A(new_n311), .ZN(new_n312));
  INV_X1    g126(.A(KEYINPUT90), .ZN(new_n313));
  AOI21_X1  g127(.A(KEYINPUT91), .B1(new_n313), .B2(new_n204), .ZN(new_n314));
  INV_X1    g128(.A(KEYINPUT91), .ZN(new_n315));
  OAI21_X1  g129(.A(G214), .B1(new_n315), .B2(G143), .ZN(new_n316));
  OR2_X1    g130(.A1(G237), .A2(G953), .ZN(new_n317));
  OAI21_X1  g131(.A(new_n314), .B1(new_n316), .B2(new_n317), .ZN(new_n318));
  OAI21_X1  g132(.A(new_n315), .B1(KEYINPUT90), .B2(G143), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n204), .A2(KEYINPUT91), .ZN(new_n320));
  NOR2_X1   g134(.A1(G237), .A2(G953), .ZN(new_n321));
  NAND4_X1  g135(.A1(new_n319), .A2(G214), .A3(new_n320), .A4(new_n321), .ZN(new_n322));
  NAND3_X1  g136(.A1(new_n318), .A2(new_n322), .A3(G131), .ZN(new_n323));
  INV_X1    g137(.A(KEYINPUT92), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n323), .A2(new_n324), .ZN(new_n325));
  NAND4_X1  g139(.A1(new_n318), .A2(new_n322), .A3(KEYINPUT92), .A4(G131), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n325), .A2(new_n326), .ZN(new_n327));
  INV_X1    g141(.A(KEYINPUT17), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n318), .A2(new_n322), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n329), .A2(new_n263), .ZN(new_n330));
  NAND3_X1  g144(.A1(new_n327), .A2(new_n328), .A3(new_n330), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n331), .A2(KEYINPUT95), .ZN(new_n332));
  INV_X1    g146(.A(KEYINPUT16), .ZN(new_n333));
  INV_X1    g147(.A(G125), .ZN(new_n334));
  OAI21_X1  g148(.A(G140), .B1(new_n334), .B2(KEYINPUT72), .ZN(new_n335));
  INV_X1    g149(.A(KEYINPUT72), .ZN(new_n336));
  INV_X1    g150(.A(G140), .ZN(new_n337));
  NAND3_X1  g151(.A1(new_n336), .A2(new_n337), .A3(G125), .ZN(new_n338));
  AOI21_X1  g152(.A(new_n333), .B1(new_n335), .B2(new_n338), .ZN(new_n339));
  AOI21_X1  g153(.A(KEYINPUT16), .B1(new_n337), .B2(G125), .ZN(new_n340));
  OR2_X1    g154(.A1(new_n339), .A2(new_n340), .ZN(new_n341));
  XNOR2_X1  g155(.A(new_n341), .B(G146), .ZN(new_n342));
  INV_X1    g156(.A(new_n342), .ZN(new_n343));
  AOI22_X1  g157(.A1(new_n325), .A2(new_n326), .B1(new_n329), .B2(new_n263), .ZN(new_n344));
  INV_X1    g158(.A(KEYINPUT95), .ZN(new_n345));
  NAND3_X1  g159(.A1(new_n344), .A2(new_n345), .A3(new_n328), .ZN(new_n346));
  NAND3_X1  g160(.A1(new_n325), .A2(KEYINPUT17), .A3(new_n326), .ZN(new_n347));
  NAND4_X1  g161(.A1(new_n332), .A2(new_n343), .A3(new_n346), .A4(new_n347), .ZN(new_n348));
  INV_X1    g162(.A(KEYINPUT18), .ZN(new_n349));
  OAI21_X1  g163(.A(new_n329), .B1(new_n349), .B2(new_n263), .ZN(new_n350));
  XNOR2_X1  g164(.A(G125), .B(G140), .ZN(new_n351));
  NAND2_X1  g165(.A1(new_n198), .A2(new_n351), .ZN(new_n352));
  AND2_X1   g166(.A1(new_n335), .A2(new_n338), .ZN(new_n353));
  OAI21_X1  g167(.A(new_n352), .B1(new_n353), .B2(new_n194), .ZN(new_n354));
  OAI211_X1 g168(.A(new_n350), .B(new_n354), .C1(new_n349), .C2(new_n323), .ZN(new_n355));
  XNOR2_X1  g169(.A(G113), .B(G122), .ZN(new_n356));
  XNOR2_X1  g170(.A(KEYINPUT94), .B(G104), .ZN(new_n357));
  XNOR2_X1  g171(.A(new_n356), .B(new_n357), .ZN(new_n358));
  NAND3_X1  g172(.A1(new_n348), .A2(new_n355), .A3(new_n358), .ZN(new_n359));
  NAND2_X1  g173(.A1(new_n341), .A2(G146), .ZN(new_n360));
  INV_X1    g174(.A(KEYINPUT19), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n351), .A2(new_n361), .ZN(new_n362));
  OAI21_X1  g176(.A(new_n362), .B1(new_n353), .B2(new_n361), .ZN(new_n363));
  OAI21_X1  g177(.A(new_n360), .B1(new_n363), .B2(new_n245), .ZN(new_n364));
  OAI21_X1  g178(.A(new_n355), .B1(new_n364), .B2(new_n344), .ZN(new_n365));
  INV_X1    g179(.A(KEYINPUT93), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n365), .A2(new_n366), .ZN(new_n367));
  INV_X1    g181(.A(new_n358), .ZN(new_n368));
  OAI211_X1 g182(.A(KEYINPUT93), .B(new_n355), .C1(new_n364), .C2(new_n344), .ZN(new_n369));
  NAND3_X1  g183(.A1(new_n367), .A2(new_n368), .A3(new_n369), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n359), .A2(new_n370), .ZN(new_n371));
  INV_X1    g185(.A(G475), .ZN(new_n372));
  NAND3_X1  g186(.A1(new_n371), .A2(new_n372), .A3(new_n188), .ZN(new_n373));
  INV_X1    g187(.A(KEYINPUT20), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n373), .A2(new_n374), .ZN(new_n375));
  AND3_X1   g189(.A1(new_n348), .A2(new_n355), .A3(new_n358), .ZN(new_n376));
  AOI21_X1  g190(.A(new_n358), .B1(new_n348), .B2(new_n355), .ZN(new_n377));
  OAI21_X1  g191(.A(new_n188), .B1(new_n376), .B2(new_n377), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n378), .A2(G475), .ZN(new_n379));
  NAND4_X1  g193(.A1(new_n371), .A2(KEYINPUT20), .A3(new_n372), .A4(new_n188), .ZN(new_n380));
  NAND3_X1  g194(.A1(new_n375), .A2(new_n379), .A3(new_n380), .ZN(new_n381));
  INV_X1    g195(.A(new_n381), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n190), .A2(G952), .ZN(new_n383));
  AOI21_X1  g197(.A(new_n383), .B1(G234), .B2(G237), .ZN(new_n384));
  INV_X1    g198(.A(new_n384), .ZN(new_n385));
  XOR2_X1   g199(.A(KEYINPUT21), .B(G898), .Z(new_n386));
  NAND2_X1  g200(.A1(G234), .A2(G237), .ZN(new_n387));
  NAND3_X1  g201(.A1(new_n387), .A2(G902), .A3(G953), .ZN(new_n388));
  OAI21_X1  g202(.A(new_n385), .B1(new_n386), .B2(new_n388), .ZN(new_n389));
  INV_X1    g203(.A(G478), .ZN(new_n390));
  NOR2_X1   g204(.A1(new_n390), .A2(KEYINPUT15), .ZN(new_n391));
  NAND2_X1  g205(.A1(new_n288), .A2(G143), .ZN(new_n392));
  XNOR2_X1  g206(.A(new_n392), .B(KEYINPUT96), .ZN(new_n393));
  OAI21_X1  g207(.A(new_n393), .B1(new_n288), .B2(G143), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n394), .A2(new_n259), .ZN(new_n395));
  INV_X1    g209(.A(G116), .ZN(new_n396));
  NAND3_X1  g210(.A1(new_n396), .A2(KEYINPUT14), .A3(G122), .ZN(new_n397));
  XNOR2_X1  g211(.A(G116), .B(G122), .ZN(new_n398));
  INV_X1    g212(.A(new_n398), .ZN(new_n399));
  OAI211_X1 g213(.A(G107), .B(new_n397), .C1(new_n399), .C2(KEYINPUT14), .ZN(new_n400));
  OAI211_X1 g214(.A(new_n393), .B(G134), .C1(new_n288), .C2(G143), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n398), .A2(new_n213), .ZN(new_n402));
  NAND4_X1  g216(.A1(new_n395), .A2(new_n400), .A3(new_n401), .A4(new_n402), .ZN(new_n403));
  INV_X1    g217(.A(KEYINPUT13), .ZN(new_n404));
  AOI21_X1  g218(.A(new_n259), .B1(new_n393), .B2(new_n404), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n405), .A2(new_n394), .ZN(new_n406));
  XNOR2_X1  g220(.A(new_n398), .B(new_n213), .ZN(new_n407));
  OAI221_X1 g221(.A(new_n393), .B1(new_n404), .B2(new_n259), .C1(new_n288), .C2(G143), .ZN(new_n408));
  NAND3_X1  g222(.A1(new_n406), .A2(new_n407), .A3(new_n408), .ZN(new_n409));
  NAND2_X1  g223(.A1(new_n403), .A2(new_n409), .ZN(new_n410));
  NAND3_X1  g224(.A1(new_n307), .A2(G217), .A3(new_n190), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n410), .A2(new_n411), .ZN(new_n412));
  INV_X1    g226(.A(new_n411), .ZN(new_n413));
  NAND3_X1  g227(.A1(new_n403), .A2(new_n409), .A3(new_n413), .ZN(new_n414));
  NAND2_X1  g228(.A1(new_n412), .A2(new_n414), .ZN(new_n415));
  INV_X1    g229(.A(KEYINPUT97), .ZN(new_n416));
  NAND3_X1  g230(.A1(new_n415), .A2(new_n416), .A3(new_n188), .ZN(new_n417));
  INV_X1    g231(.A(new_n417), .ZN(new_n418));
  AOI21_X1  g232(.A(new_n416), .B1(new_n415), .B2(new_n188), .ZN(new_n419));
  OAI21_X1  g233(.A(new_n391), .B1(new_n418), .B2(new_n419), .ZN(new_n420));
  OR2_X1    g234(.A1(new_n419), .A2(new_n391), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n420), .A2(new_n421), .ZN(new_n422));
  INV_X1    g236(.A(new_n422), .ZN(new_n423));
  AND3_X1   g237(.A1(new_n382), .A2(new_n389), .A3(new_n423), .ZN(new_n424));
  OAI21_X1  g238(.A(G214), .B1(G237), .B2(G902), .ZN(new_n425));
  INV_X1    g239(.A(new_n425), .ZN(new_n426));
  XNOR2_X1  g240(.A(KEYINPUT2), .B(G113), .ZN(new_n427));
  INV_X1    g241(.A(new_n427), .ZN(new_n428));
  XNOR2_X1  g242(.A(G116), .B(G119), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n428), .A2(new_n429), .ZN(new_n430));
  INV_X1    g244(.A(new_n429), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n431), .A2(new_n427), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n430), .A2(new_n432), .ZN(new_n433));
  OAI211_X1 g247(.A(new_n433), .B(new_n238), .C1(new_n241), .C2(new_n242), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n434), .A2(KEYINPUT84), .ZN(new_n435));
  INV_X1    g249(.A(KEYINPUT84), .ZN(new_n436));
  NAND4_X1  g250(.A1(new_n277), .A2(new_n436), .A3(new_n433), .A4(new_n238), .ZN(new_n437));
  INV_X1    g251(.A(KEYINPUT5), .ZN(new_n438));
  NOR2_X1   g252(.A1(new_n431), .A2(new_n438), .ZN(new_n439));
  INV_X1    g253(.A(new_n439), .ZN(new_n440));
  INV_X1    g254(.A(G113), .ZN(new_n441));
  NOR2_X1   g255(.A1(new_n396), .A2(G119), .ZN(new_n442));
  AOI21_X1  g256(.A(new_n441), .B1(new_n442), .B2(new_n438), .ZN(new_n443));
  AOI22_X1  g257(.A1(new_n440), .A2(new_n443), .B1(new_n428), .B2(new_n429), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n444), .A2(new_n227), .ZN(new_n445));
  NAND3_X1  g259(.A1(new_n435), .A2(new_n437), .A3(new_n445), .ZN(new_n446));
  XOR2_X1   g260(.A(G110), .B(G122), .Z(new_n447));
  NAND2_X1  g261(.A1(new_n446), .A2(new_n447), .ZN(new_n448));
  INV_X1    g262(.A(new_n447), .ZN(new_n449));
  NAND4_X1  g263(.A1(new_n435), .A2(new_n437), .A3(new_n449), .A4(new_n445), .ZN(new_n450));
  NAND3_X1  g264(.A1(new_n448), .A2(KEYINPUT6), .A3(new_n450), .ZN(new_n451));
  INV_X1    g265(.A(KEYINPUT6), .ZN(new_n452));
  NAND3_X1  g266(.A1(new_n446), .A2(new_n452), .A3(new_n447), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n290), .A2(new_n334), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n251), .A2(G125), .ZN(new_n455));
  AND2_X1   g269(.A1(new_n455), .A2(KEYINPUT85), .ZN(new_n456));
  NOR2_X1   g270(.A1(new_n455), .A2(KEYINPUT85), .ZN(new_n457));
  OAI21_X1  g271(.A(new_n454), .B1(new_n456), .B2(new_n457), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n190), .A2(G224), .ZN(new_n459));
  XNOR2_X1  g273(.A(new_n459), .B(KEYINPUT86), .ZN(new_n460));
  XNOR2_X1  g274(.A(new_n458), .B(new_n460), .ZN(new_n461));
  NAND3_X1  g275(.A1(new_n451), .A2(new_n453), .A3(new_n461), .ZN(new_n462));
  XNOR2_X1  g276(.A(new_n443), .B(KEYINPUT87), .ZN(new_n463));
  OAI21_X1  g277(.A(new_n430), .B1(new_n463), .B2(new_n439), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n464), .A2(new_n227), .ZN(new_n465));
  XOR2_X1   g279(.A(new_n447), .B(KEYINPUT8), .Z(new_n466));
  NAND2_X1  g280(.A1(new_n444), .A2(new_n223), .ZN(new_n467));
  AND3_X1   g281(.A1(new_n465), .A2(new_n466), .A3(new_n467), .ZN(new_n468));
  OR2_X1    g282(.A1(new_n468), .A2(KEYINPUT88), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n459), .A2(KEYINPUT7), .ZN(new_n470));
  NAND2_X1  g284(.A1(new_n454), .A2(new_n455), .ZN(new_n471));
  AOI22_X1  g285(.A1(new_n468), .A2(KEYINPUT88), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  OR2_X1    g286(.A1(new_n458), .A2(new_n470), .ZN(new_n473));
  NAND4_X1  g287(.A1(new_n469), .A2(new_n472), .A3(new_n450), .A4(new_n473), .ZN(new_n474));
  NAND3_X1  g288(.A1(new_n462), .A2(new_n188), .A3(new_n474), .ZN(new_n475));
  OAI21_X1  g289(.A(G210), .B1(G237), .B2(G902), .ZN(new_n476));
  XOR2_X1   g290(.A(new_n476), .B(KEYINPUT89), .Z(new_n477));
  NAND2_X1  g291(.A1(new_n475), .A2(new_n477), .ZN(new_n478));
  INV_X1    g292(.A(new_n477), .ZN(new_n479));
  NAND4_X1  g293(.A1(new_n462), .A2(new_n188), .A3(new_n479), .A4(new_n474), .ZN(new_n480));
  AOI21_X1  g294(.A(new_n426), .B1(new_n478), .B2(new_n480), .ZN(new_n481));
  NAND3_X1  g295(.A1(new_n312), .A2(new_n424), .A3(new_n481), .ZN(new_n482));
  INV_X1    g296(.A(new_n482), .ZN(new_n483));
  INV_X1    g297(.A(KEYINPUT32), .ZN(new_n484));
  XNOR2_X1  g298(.A(KEYINPUT69), .B(KEYINPUT27), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n321), .A2(G210), .ZN(new_n486));
  XNOR2_X1  g300(.A(new_n485), .B(new_n486), .ZN(new_n487));
  XNOR2_X1  g301(.A(KEYINPUT26), .B(G101), .ZN(new_n488));
  XNOR2_X1  g302(.A(new_n487), .B(new_n488), .ZN(new_n489));
  INV_X1    g303(.A(new_n489), .ZN(new_n490));
  INV_X1    g304(.A(KEYINPUT28), .ZN(new_n491));
  INV_X1    g305(.A(new_n264), .ZN(new_n492));
  NOR2_X1   g306(.A1(new_n259), .A2(G137), .ZN(new_n493));
  OAI21_X1  g307(.A(G131), .B1(new_n492), .B2(new_n493), .ZN(new_n494));
  AND2_X1   g308(.A1(new_n265), .A2(KEYINPUT65), .ZN(new_n495));
  NOR2_X1   g309(.A1(new_n265), .A2(KEYINPUT65), .ZN(new_n496));
  OAI21_X1  g310(.A(new_n494), .B1(new_n495), .B2(new_n496), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n497), .A2(KEYINPUT67), .ZN(new_n498));
  INV_X1    g312(.A(KEYINPUT67), .ZN(new_n499));
  NAND3_X1  g313(.A1(new_n266), .A2(new_n499), .A3(new_n494), .ZN(new_n500));
  NAND3_X1  g314(.A1(new_n498), .A2(new_n232), .A3(new_n500), .ZN(new_n501));
  INV_X1    g315(.A(KEYINPUT68), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  AOI21_X1  g317(.A(new_n433), .B1(new_n280), .B2(new_n269), .ZN(new_n504));
  NAND4_X1  g318(.A1(new_n498), .A2(new_n500), .A3(KEYINPUT68), .A4(new_n232), .ZN(new_n505));
  NAND3_X1  g319(.A1(new_n503), .A2(new_n504), .A3(new_n505), .ZN(new_n506));
  OAI22_X1  g320(.A1(new_n282), .A2(new_n251), .B1(new_n290), .B2(new_n497), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n507), .A2(new_n433), .ZN(new_n508));
  AOI21_X1  g322(.A(new_n491), .B1(new_n506), .B2(new_n508), .ZN(new_n509));
  AOI21_X1  g323(.A(KEYINPUT28), .B1(new_n504), .B2(new_n501), .ZN(new_n510));
  OAI21_X1  g324(.A(new_n490), .B1(new_n509), .B2(new_n510), .ZN(new_n511));
  AND2_X1   g325(.A1(new_n506), .A2(new_n489), .ZN(new_n512));
  INV_X1    g326(.A(KEYINPUT31), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n280), .A2(new_n269), .ZN(new_n514));
  NAND4_X1  g328(.A1(new_n503), .A2(KEYINPUT30), .A3(new_n514), .A4(new_n505), .ZN(new_n515));
  INV_X1    g329(.A(KEYINPUT30), .ZN(new_n516));
  AOI22_X1  g330(.A1(new_n507), .A2(new_n516), .B1(new_n430), .B2(new_n432), .ZN(new_n517));
  NAND2_X1  g331(.A1(new_n515), .A2(new_n517), .ZN(new_n518));
  NAND3_X1  g332(.A1(new_n512), .A2(new_n513), .A3(new_n518), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n511), .A2(new_n519), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n512), .A2(new_n518), .ZN(new_n521));
  AOI21_X1  g335(.A(KEYINPUT70), .B1(new_n521), .B2(KEYINPUT31), .ZN(new_n522));
  INV_X1    g336(.A(KEYINPUT70), .ZN(new_n523));
  AOI211_X1 g337(.A(new_n523), .B(new_n513), .C1(new_n512), .C2(new_n518), .ZN(new_n524));
  NOR3_X1   g338(.A1(new_n520), .A2(new_n522), .A3(new_n524), .ZN(new_n525));
  NOR2_X1   g339(.A1(G472), .A2(G902), .ZN(new_n526));
  INV_X1    g340(.A(new_n526), .ZN(new_n527));
  OAI21_X1  g341(.A(new_n484), .B1(new_n525), .B2(new_n527), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n506), .A2(new_n489), .ZN(new_n529));
  AOI21_X1  g343(.A(new_n529), .B1(new_n515), .B2(new_n517), .ZN(new_n530));
  OAI21_X1  g344(.A(new_n523), .B1(new_n530), .B2(new_n513), .ZN(new_n531));
  NAND3_X1  g345(.A1(new_n521), .A2(KEYINPUT70), .A3(KEYINPUT31), .ZN(new_n532));
  NAND4_X1  g346(.A1(new_n531), .A2(new_n511), .A3(new_n519), .A4(new_n532), .ZN(new_n533));
  NAND3_X1  g347(.A1(new_n533), .A2(KEYINPUT32), .A3(new_n526), .ZN(new_n534));
  NAND3_X1  g348(.A1(new_n503), .A2(new_n514), .A3(new_n505), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n535), .A2(new_n433), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n536), .A2(new_n506), .ZN(new_n537));
  AOI21_X1  g351(.A(new_n510), .B1(new_n537), .B2(KEYINPUT28), .ZN(new_n538));
  NAND3_X1  g352(.A1(new_n538), .A2(KEYINPUT29), .A3(new_n489), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n539), .A2(new_n188), .ZN(new_n540));
  NOR3_X1   g354(.A1(new_n509), .A2(new_n510), .A3(new_n490), .ZN(new_n541));
  AOI21_X1  g355(.A(new_n489), .B1(new_n518), .B2(new_n506), .ZN(new_n542));
  NOR3_X1   g356(.A1(new_n541), .A2(new_n542), .A3(KEYINPUT29), .ZN(new_n543));
  OAI21_X1  g357(.A(G472), .B1(new_n540), .B2(new_n543), .ZN(new_n544));
  NAND3_X1  g358(.A1(new_n528), .A2(new_n534), .A3(new_n544), .ZN(new_n545));
  INV_X1    g359(.A(KEYINPUT77), .ZN(new_n546));
  XOR2_X1   g360(.A(KEYINPUT73), .B(KEYINPUT74), .Z(new_n547));
  NAND3_X1  g361(.A1(new_n190), .A2(G221), .A3(G234), .ZN(new_n548));
  XNOR2_X1  g362(.A(new_n547), .B(new_n548), .ZN(new_n549));
  XNOR2_X1  g363(.A(KEYINPUT22), .B(G137), .ZN(new_n550));
  XNOR2_X1  g364(.A(new_n549), .B(new_n550), .ZN(new_n551));
  INV_X1    g365(.A(KEYINPUT75), .ZN(new_n552));
  XNOR2_X1  g366(.A(new_n551), .B(new_n552), .ZN(new_n553));
  INV_X1    g367(.A(G119), .ZN(new_n554));
  NOR2_X1   g368(.A1(new_n554), .A2(G128), .ZN(new_n555));
  OR2_X1    g369(.A1(new_n555), .A2(KEYINPUT23), .ZN(new_n556));
  NOR2_X1   g370(.A1(new_n288), .A2(G119), .ZN(new_n557));
  INV_X1    g371(.A(new_n557), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n555), .A2(KEYINPUT23), .ZN(new_n559));
  NAND3_X1  g373(.A1(new_n556), .A2(new_n558), .A3(new_n559), .ZN(new_n560));
  XNOR2_X1  g374(.A(new_n560), .B(KEYINPUT71), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n561), .A2(G110), .ZN(new_n562));
  NOR2_X1   g376(.A1(new_n557), .A2(new_n555), .ZN(new_n563));
  XOR2_X1   g377(.A(KEYINPUT24), .B(G110), .Z(new_n564));
  NAND2_X1  g378(.A1(new_n563), .A2(new_n564), .ZN(new_n565));
  NAND3_X1  g379(.A1(new_n562), .A2(new_n342), .A3(new_n565), .ZN(new_n566));
  OAI22_X1  g380(.A1(new_n560), .A2(G110), .B1(new_n563), .B2(new_n564), .ZN(new_n567));
  NAND3_X1  g381(.A1(new_n567), .A2(new_n360), .A3(new_n352), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n566), .A2(new_n568), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n553), .A2(new_n569), .ZN(new_n570));
  INV_X1    g384(.A(new_n551), .ZN(new_n571));
  OAI21_X1  g385(.A(new_n570), .B1(new_n569), .B2(new_n571), .ZN(new_n572));
  NAND2_X1  g386(.A1(new_n572), .A2(new_n188), .ZN(new_n573));
  NAND2_X1  g387(.A1(new_n573), .A2(KEYINPUT25), .ZN(new_n574));
  INV_X1    g388(.A(G217), .ZN(new_n575));
  AOI21_X1  g389(.A(new_n575), .B1(G234), .B2(new_n188), .ZN(new_n576));
  INV_X1    g390(.A(KEYINPUT25), .ZN(new_n577));
  NAND3_X1  g391(.A1(new_n572), .A2(new_n577), .A3(new_n188), .ZN(new_n578));
  NAND3_X1  g392(.A1(new_n574), .A2(new_n576), .A3(new_n578), .ZN(new_n579));
  OR2_X1    g393(.A1(new_n572), .A2(KEYINPUT76), .ZN(new_n580));
  NOR2_X1   g394(.A1(new_n576), .A2(G902), .ZN(new_n581));
  NAND2_X1  g395(.A1(new_n572), .A2(KEYINPUT76), .ZN(new_n582));
  NAND3_X1  g396(.A1(new_n580), .A2(new_n581), .A3(new_n582), .ZN(new_n583));
  AND2_X1   g397(.A1(new_n579), .A2(new_n583), .ZN(new_n584));
  NAND3_X1  g398(.A1(new_n545), .A2(new_n546), .A3(new_n584), .ZN(new_n585));
  INV_X1    g399(.A(new_n585), .ZN(new_n586));
  AOI21_X1  g400(.A(new_n546), .B1(new_n545), .B2(new_n584), .ZN(new_n587));
  OAI21_X1  g401(.A(new_n483), .B1(new_n586), .B2(new_n587), .ZN(new_n588));
  XNOR2_X1  g402(.A(new_n588), .B(G101), .ZN(G3));
  NAND2_X1  g403(.A1(new_n533), .A2(new_n188), .ZN(new_n590));
  NAND2_X1  g404(.A1(KEYINPUT98), .A2(G472), .ZN(new_n591));
  XNOR2_X1  g405(.A(new_n590), .B(new_n591), .ZN(new_n592));
  NAND3_X1  g406(.A1(new_n592), .A2(new_n584), .A3(new_n312), .ZN(new_n593));
  NAND2_X1  g407(.A1(new_n411), .A2(KEYINPUT100), .ZN(new_n594));
  NAND2_X1  g408(.A1(new_n594), .A2(KEYINPUT33), .ZN(new_n595));
  INV_X1    g409(.A(new_n414), .ZN(new_n596));
  AOI21_X1  g410(.A(new_n413), .B1(new_n403), .B2(new_n409), .ZN(new_n597));
  OAI21_X1  g411(.A(new_n595), .B1(new_n596), .B2(new_n597), .ZN(new_n598));
  NAND4_X1  g412(.A1(new_n412), .A2(KEYINPUT33), .A3(new_n414), .A4(new_n594), .ZN(new_n599));
  NAND4_X1  g413(.A1(new_n598), .A2(new_n599), .A3(G478), .A4(new_n188), .ZN(new_n600));
  OR2_X1    g414(.A1(new_n600), .A2(KEYINPUT101), .ZN(new_n601));
  INV_X1    g415(.A(new_n415), .ZN(new_n602));
  OAI21_X1  g416(.A(new_n390), .B1(new_n602), .B2(G902), .ZN(new_n603));
  NAND2_X1  g417(.A1(new_n600), .A2(KEYINPUT101), .ZN(new_n604));
  NAND3_X1  g418(.A1(new_n601), .A2(new_n603), .A3(new_n604), .ZN(new_n605));
  NAND2_X1  g419(.A1(new_n381), .A2(new_n605), .ZN(new_n606));
  NAND3_X1  g420(.A1(new_n478), .A2(KEYINPUT99), .A3(new_n480), .ZN(new_n607));
  INV_X1    g421(.A(KEYINPUT99), .ZN(new_n608));
  NAND3_X1  g422(.A1(new_n475), .A2(new_n608), .A3(new_n477), .ZN(new_n609));
  NAND4_X1  g423(.A1(new_n607), .A2(new_n389), .A3(new_n425), .A4(new_n609), .ZN(new_n610));
  NOR3_X1   g424(.A1(new_n593), .A2(new_n606), .A3(new_n610), .ZN(new_n611));
  XNOR2_X1  g425(.A(KEYINPUT34), .B(G104), .ZN(new_n612));
  XNOR2_X1  g426(.A(new_n611), .B(new_n612), .ZN(G6));
  NOR2_X1   g427(.A1(new_n381), .A2(new_n423), .ZN(new_n614));
  INV_X1    g428(.A(new_n614), .ZN(new_n615));
  NOR3_X1   g429(.A1(new_n593), .A2(new_n610), .A3(new_n615), .ZN(new_n616));
  XNOR2_X1  g430(.A(KEYINPUT35), .B(G107), .ZN(new_n617));
  XNOR2_X1  g431(.A(new_n616), .B(new_n617), .ZN(G9));
  NOR2_X1   g432(.A1(new_n522), .A2(new_n524), .ZN(new_n619));
  INV_X1    g433(.A(new_n520), .ZN(new_n620));
  AOI21_X1  g434(.A(G902), .B1(new_n619), .B2(new_n620), .ZN(new_n621));
  XNOR2_X1  g435(.A(new_n621), .B(new_n591), .ZN(new_n622));
  INV_X1    g436(.A(KEYINPUT36), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n553), .A2(new_n623), .ZN(new_n624));
  XOR2_X1   g438(.A(new_n624), .B(new_n569), .Z(new_n625));
  NAND2_X1  g439(.A1(new_n625), .A2(new_n581), .ZN(new_n626));
  AND2_X1   g440(.A1(new_n579), .A2(new_n626), .ZN(new_n627));
  NOR3_X1   g441(.A1(new_n482), .A2(new_n622), .A3(new_n627), .ZN(new_n628));
  XNOR2_X1  g442(.A(KEYINPUT37), .B(G110), .ZN(new_n629));
  XNOR2_X1  g443(.A(new_n628), .B(new_n629), .ZN(G12));
  AND3_X1   g444(.A1(new_n478), .A2(KEYINPUT99), .A3(new_n480), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n609), .A2(new_n425), .ZN(new_n632));
  NOR3_X1   g446(.A1(new_n631), .A2(new_n627), .A3(new_n632), .ZN(new_n633));
  OAI21_X1  g447(.A(new_n385), .B1(new_n388), .B2(G900), .ZN(new_n634));
  AND2_X1   g448(.A1(new_n614), .A2(new_n634), .ZN(new_n635));
  NAND4_X1  g449(.A1(new_n633), .A2(new_n545), .A3(new_n312), .A4(new_n635), .ZN(new_n636));
  XOR2_X1   g450(.A(KEYINPUT102), .B(G128), .Z(new_n637));
  XNOR2_X1  g451(.A(new_n636), .B(new_n637), .ZN(G30));
  NAND2_X1  g452(.A1(new_n381), .A2(new_n422), .ZN(new_n639));
  XNOR2_X1  g453(.A(new_n634), .B(KEYINPUT39), .ZN(new_n640));
  NAND2_X1  g454(.A1(new_n312), .A2(new_n640), .ZN(new_n641));
  AOI211_X1 g455(.A(new_n426), .B(new_n639), .C1(new_n641), .C2(KEYINPUT40), .ZN(new_n642));
  NAND2_X1  g456(.A1(new_n478), .A2(new_n480), .ZN(new_n643));
  XNOR2_X1  g457(.A(KEYINPUT103), .B(KEYINPUT38), .ZN(new_n644));
  XNOR2_X1  g458(.A(new_n643), .B(new_n644), .ZN(new_n645));
  INV_X1    g459(.A(new_n645), .ZN(new_n646));
  OAI211_X1 g460(.A(new_n642), .B(new_n646), .C1(KEYINPUT40), .C2(new_n641), .ZN(new_n647));
  NAND2_X1  g461(.A1(new_n579), .A2(new_n626), .ZN(new_n648));
  OAI21_X1  g462(.A(new_n188), .B1(new_n537), .B2(new_n489), .ZN(new_n649));
  AOI21_X1  g463(.A(new_n490), .B1(new_n518), .B2(new_n506), .ZN(new_n650));
  OAI21_X1  g464(.A(G472), .B1(new_n649), .B2(new_n650), .ZN(new_n651));
  NAND3_X1  g465(.A1(new_n528), .A2(new_n534), .A3(new_n651), .ZN(new_n652));
  INV_X1    g466(.A(new_n652), .ZN(new_n653));
  NOR3_X1   g467(.A1(new_n647), .A2(new_n648), .A3(new_n653), .ZN(new_n654));
  XNOR2_X1  g468(.A(new_n654), .B(new_n204), .ZN(G45));
  NAND3_X1  g469(.A1(new_n381), .A2(new_n605), .A3(new_n634), .ZN(new_n656));
  NAND2_X1  g470(.A1(new_n656), .A2(KEYINPUT104), .ZN(new_n657));
  INV_X1    g471(.A(KEYINPUT104), .ZN(new_n658));
  NAND4_X1  g472(.A1(new_n381), .A2(new_n605), .A3(new_n658), .A4(new_n634), .ZN(new_n659));
  AND2_X1   g473(.A1(new_n657), .A2(new_n659), .ZN(new_n660));
  NAND4_X1  g474(.A1(new_n660), .A2(new_n633), .A3(new_n545), .A4(new_n312), .ZN(new_n661));
  XNOR2_X1  g475(.A(new_n661), .B(G146), .ZN(G48));
  NOR2_X1   g476(.A1(new_n610), .A2(new_n606), .ZN(new_n663));
  NOR2_X1   g477(.A1(new_n187), .A2(KEYINPUT105), .ZN(new_n664));
  AND3_X1   g478(.A1(new_n257), .A2(KEYINPUT83), .A3(new_n269), .ZN(new_n665));
  AOI21_X1  g479(.A(KEYINPUT83), .B1(new_n257), .B2(new_n269), .ZN(new_n666));
  OAI21_X1  g480(.A(new_n283), .B1(new_n665), .B2(new_n666), .ZN(new_n667));
  INV_X1    g481(.A(new_n192), .ZN(new_n668));
  AOI21_X1  g482(.A(new_n297), .B1(new_n667), .B2(new_n668), .ZN(new_n669));
  OAI21_X1  g483(.A(new_n664), .B1(new_n669), .B2(G902), .ZN(new_n670));
  INV_X1    g484(.A(new_n664), .ZN(new_n671));
  OAI211_X1 g485(.A(new_n188), .B(new_n671), .C1(new_n284), .C2(new_n297), .ZN(new_n672));
  AND3_X1   g486(.A1(new_n670), .A2(new_n672), .A3(new_n309), .ZN(new_n673));
  NAND4_X1  g487(.A1(new_n663), .A2(new_n584), .A3(new_n545), .A4(new_n673), .ZN(new_n674));
  XNOR2_X1  g488(.A(KEYINPUT41), .B(G113), .ZN(new_n675));
  XNOR2_X1  g489(.A(new_n674), .B(new_n675), .ZN(G15));
  NOR2_X1   g490(.A1(new_n610), .A2(new_n615), .ZN(new_n677));
  NAND4_X1  g491(.A1(new_n677), .A2(new_n584), .A3(new_n545), .A4(new_n673), .ZN(new_n678));
  XNOR2_X1  g492(.A(new_n678), .B(G116), .ZN(G18));
  NAND2_X1  g493(.A1(new_n545), .A2(new_n424), .ZN(new_n680));
  INV_X1    g494(.A(new_n632), .ZN(new_n681));
  NAND4_X1  g495(.A1(new_n681), .A2(new_n673), .A3(new_n607), .A4(new_n648), .ZN(new_n682));
  OAI21_X1  g496(.A(KEYINPUT106), .B1(new_n680), .B2(new_n682), .ZN(new_n683));
  INV_X1    g497(.A(new_n682), .ZN(new_n684));
  INV_X1    g498(.A(KEYINPUT106), .ZN(new_n685));
  NAND4_X1  g499(.A1(new_n684), .A2(new_n685), .A3(new_n545), .A4(new_n424), .ZN(new_n686));
  NAND2_X1  g500(.A1(new_n683), .A2(new_n686), .ZN(new_n687));
  XNOR2_X1  g501(.A(new_n687), .B(G119), .ZN(G21));
  NOR2_X1   g502(.A1(new_n538), .A2(new_n489), .ZN(new_n689));
  NAND2_X1  g503(.A1(new_n521), .A2(KEYINPUT31), .ZN(new_n690));
  NAND2_X1  g504(.A1(new_n690), .A2(new_n519), .ZN(new_n691));
  OAI21_X1  g505(.A(new_n526), .B1(new_n689), .B2(new_n691), .ZN(new_n692));
  INV_X1    g506(.A(G472), .ZN(new_n693));
  OAI211_X1 g507(.A(new_n584), .B(new_n692), .C1(new_n621), .C2(new_n693), .ZN(new_n694));
  INV_X1    g508(.A(new_n639), .ZN(new_n695));
  NAND2_X1  g509(.A1(new_n673), .A2(new_n695), .ZN(new_n696));
  NOR3_X1   g510(.A1(new_n694), .A2(new_n696), .A3(new_n610), .ZN(new_n697));
  XOR2_X1   g511(.A(new_n697), .B(G122), .Z(G24));
  NAND3_X1  g512(.A1(new_n670), .A2(new_n672), .A3(new_n309), .ZN(new_n699));
  NOR3_X1   g513(.A1(new_n631), .A2(new_n632), .A3(new_n699), .ZN(new_n700));
  INV_X1    g514(.A(new_n689), .ZN(new_n701));
  INV_X1    g515(.A(new_n691), .ZN(new_n702));
  AOI21_X1  g516(.A(new_n527), .B1(new_n701), .B2(new_n702), .ZN(new_n703));
  AOI21_X1  g517(.A(new_n703), .B1(G472), .B2(new_n590), .ZN(new_n704));
  NAND4_X1  g518(.A1(new_n660), .A2(new_n700), .A3(new_n704), .A4(new_n648), .ZN(new_n705));
  XNOR2_X1  g519(.A(KEYINPUT107), .B(G125), .ZN(new_n706));
  XNOR2_X1  g520(.A(new_n705), .B(new_n706), .ZN(G27));
  INV_X1    g521(.A(KEYINPUT42), .ZN(new_n708));
  INV_X1    g522(.A(new_n309), .ZN(new_n709));
  INV_X1    g523(.A(KEYINPUT108), .ZN(new_n710));
  NAND2_X1  g524(.A1(new_n305), .A2(new_n710), .ZN(new_n711));
  NAND4_X1  g525(.A1(new_n298), .A2(new_n304), .A3(KEYINPUT108), .A4(new_n299), .ZN(new_n712));
  AOI21_X1  g526(.A(new_n709), .B1(new_n711), .B2(new_n712), .ZN(new_n713));
  NAND3_X1  g527(.A1(new_n478), .A2(new_n425), .A3(new_n480), .ZN(new_n714));
  INV_X1    g528(.A(new_n714), .ZN(new_n715));
  NAND3_X1  g529(.A1(new_n660), .A2(new_n713), .A3(new_n715), .ZN(new_n716));
  NAND2_X1  g530(.A1(new_n545), .A2(new_n584), .ZN(new_n717));
  OAI21_X1  g531(.A(new_n708), .B1(new_n716), .B2(new_n717), .ZN(new_n718));
  INV_X1    g532(.A(new_n584), .ZN(new_n719));
  AND3_X1   g533(.A1(new_n533), .A2(KEYINPUT32), .A3(new_n526), .ZN(new_n720));
  AOI21_X1  g534(.A(KEYINPUT32), .B1(new_n533), .B2(new_n526), .ZN(new_n721));
  NOR2_X1   g535(.A1(new_n720), .A2(new_n721), .ZN(new_n722));
  AOI21_X1  g536(.A(new_n719), .B1(new_n722), .B2(new_n544), .ZN(new_n723));
  AOI211_X1 g537(.A(new_n709), .B(new_n714), .C1(new_n711), .C2(new_n712), .ZN(new_n724));
  NAND4_X1  g538(.A1(new_n723), .A2(KEYINPUT42), .A3(new_n660), .A4(new_n724), .ZN(new_n725));
  NAND2_X1  g539(.A1(new_n718), .A2(new_n725), .ZN(new_n726));
  XNOR2_X1  g540(.A(new_n726), .B(G131), .ZN(G33));
  INV_X1    g541(.A(KEYINPUT109), .ZN(new_n728));
  NAND4_X1  g542(.A1(new_n723), .A2(new_n728), .A3(new_n635), .A4(new_n724), .ZN(new_n729));
  NAND3_X1  g543(.A1(new_n545), .A2(new_n584), .A3(new_n635), .ZN(new_n730));
  NAND2_X1  g544(.A1(new_n711), .A2(new_n712), .ZN(new_n731));
  NAND3_X1  g545(.A1(new_n731), .A2(new_n309), .A3(new_n715), .ZN(new_n732));
  OAI21_X1  g546(.A(KEYINPUT109), .B1(new_n730), .B2(new_n732), .ZN(new_n733));
  NAND2_X1  g547(.A1(new_n729), .A2(new_n733), .ZN(new_n734));
  XNOR2_X1  g548(.A(new_n734), .B(G134), .ZN(G36));
  OAI211_X1 g549(.A(KEYINPUT110), .B(G469), .C1(new_n303), .C2(KEYINPUT45), .ZN(new_n736));
  INV_X1    g550(.A(KEYINPUT110), .ZN(new_n737));
  OAI211_X1 g551(.A(new_n283), .B(new_n192), .C1(new_n665), .C2(new_n666), .ZN(new_n738));
  INV_X1    g552(.A(new_n283), .ZN(new_n739));
  OAI21_X1  g553(.A(new_n668), .B1(new_n295), .B2(new_n739), .ZN(new_n740));
  AOI21_X1  g554(.A(KEYINPUT45), .B1(new_n738), .B2(new_n740), .ZN(new_n741));
  OAI21_X1  g555(.A(new_n737), .B1(new_n741), .B2(new_n187), .ZN(new_n742));
  NAND2_X1  g556(.A1(new_n303), .A2(KEYINPUT45), .ZN(new_n743));
  NAND3_X1  g557(.A1(new_n736), .A2(new_n742), .A3(new_n743), .ZN(new_n744));
  AOI21_X1  g558(.A(KEYINPUT46), .B1(new_n744), .B2(new_n299), .ZN(new_n745));
  OR2_X1    g559(.A1(new_n745), .A2(KEYINPUT111), .ZN(new_n746));
  NAND3_X1  g560(.A1(new_n744), .A2(KEYINPUT46), .A3(new_n299), .ZN(new_n747));
  NAND2_X1  g561(.A1(new_n745), .A2(KEYINPUT111), .ZN(new_n748));
  NAND4_X1  g562(.A1(new_n746), .A2(new_n747), .A3(new_n298), .A4(new_n748), .ZN(new_n749));
  INV_X1    g563(.A(new_n749), .ZN(new_n750));
  NOR2_X1   g564(.A1(new_n750), .A2(new_n709), .ZN(new_n751));
  AND2_X1   g565(.A1(new_n751), .A2(new_n640), .ZN(new_n752));
  NAND2_X1  g566(.A1(new_n382), .A2(new_n605), .ZN(new_n753));
  XOR2_X1   g567(.A(new_n753), .B(KEYINPUT43), .Z(new_n754));
  NAND3_X1  g568(.A1(new_n754), .A2(new_n622), .A3(new_n648), .ZN(new_n755));
  XNOR2_X1  g569(.A(new_n755), .B(KEYINPUT44), .ZN(new_n756));
  XOR2_X1   g570(.A(new_n714), .B(KEYINPUT112), .Z(new_n757));
  INV_X1    g571(.A(new_n757), .ZN(new_n758));
  NAND3_X1  g572(.A1(new_n752), .A2(new_n756), .A3(new_n758), .ZN(new_n759));
  XNOR2_X1  g573(.A(new_n759), .B(G137), .ZN(G39));
  AND3_X1   g574(.A1(new_n749), .A2(KEYINPUT47), .A3(new_n309), .ZN(new_n761));
  INV_X1    g575(.A(new_n761), .ZN(new_n762));
  AOI21_X1  g576(.A(KEYINPUT47), .B1(new_n749), .B2(new_n309), .ZN(new_n763));
  INV_X1    g577(.A(new_n763), .ZN(new_n764));
  AOI21_X1  g578(.A(new_n545), .B1(new_n762), .B2(new_n764), .ZN(new_n765));
  NAND4_X1  g579(.A1(new_n765), .A2(new_n719), .A3(new_n660), .A4(new_n715), .ZN(new_n766));
  XNOR2_X1  g580(.A(new_n766), .B(G140), .ZN(G42));
  AND3_X1   g581(.A1(new_n545), .A2(new_n584), .A3(new_n673), .ZN(new_n768));
  AOI21_X1  g582(.A(new_n697), .B1(new_n768), .B2(new_n663), .ZN(new_n769));
  NAND2_X1  g583(.A1(new_n615), .A2(new_n606), .ZN(new_n770));
  AND3_X1   g584(.A1(new_n770), .A2(new_n389), .A3(new_n481), .ZN(new_n771));
  NAND4_X1  g585(.A1(new_n771), .A2(new_n584), .A3(new_n312), .A4(new_n592), .ZN(new_n772));
  NAND4_X1  g586(.A1(new_n687), .A2(new_n769), .A3(new_n678), .A4(new_n772), .ZN(new_n773));
  INV_X1    g587(.A(new_n628), .ZN(new_n774));
  NAND2_X1  g588(.A1(new_n588), .A2(new_n774), .ZN(new_n775));
  NOR2_X1   g589(.A1(new_n773), .A2(new_n775), .ZN(new_n776));
  NAND2_X1  g590(.A1(new_n590), .A2(G472), .ZN(new_n777));
  NAND4_X1  g591(.A1(new_n777), .A2(new_n657), .A3(new_n659), .A4(new_n692), .ZN(new_n778));
  NOR2_X1   g592(.A1(new_n732), .A2(new_n778), .ZN(new_n779));
  AND3_X1   g593(.A1(new_n382), .A2(new_n423), .A3(new_n634), .ZN(new_n780));
  AND4_X1   g594(.A1(new_n545), .A2(new_n780), .A3(new_n312), .A4(new_n715), .ZN(new_n781));
  OAI21_X1  g595(.A(new_n648), .B1(new_n779), .B2(new_n781), .ZN(new_n782));
  AND3_X1   g596(.A1(new_n726), .A2(new_n734), .A3(new_n782), .ZN(new_n783));
  INV_X1    g597(.A(KEYINPUT52), .ZN(new_n784));
  NAND3_X1  g598(.A1(new_n661), .A2(new_n705), .A3(new_n636), .ZN(new_n785));
  NAND3_X1  g599(.A1(new_n652), .A2(new_n627), .A3(new_n634), .ZN(new_n786));
  NOR3_X1   g600(.A1(new_n631), .A2(new_n632), .A3(new_n639), .ZN(new_n787));
  NAND2_X1  g601(.A1(new_n713), .A2(new_n787), .ZN(new_n788));
  NOR2_X1   g602(.A1(new_n786), .A2(new_n788), .ZN(new_n789));
  OAI21_X1  g603(.A(new_n784), .B1(new_n785), .B2(new_n789), .ZN(new_n790));
  AOI21_X1  g604(.A(new_n311), .B1(new_n722), .B2(new_n544), .ZN(new_n791));
  OAI211_X1 g605(.A(new_n791), .B(new_n633), .C1(new_n635), .C2(new_n660), .ZN(new_n792));
  AND3_X1   g606(.A1(new_n652), .A2(new_n627), .A3(new_n634), .ZN(new_n793));
  AND2_X1   g607(.A1(new_n713), .A2(new_n787), .ZN(new_n794));
  NAND2_X1  g608(.A1(new_n793), .A2(new_n794), .ZN(new_n795));
  NAND4_X1  g609(.A1(new_n792), .A2(new_n795), .A3(KEYINPUT52), .A4(new_n705), .ZN(new_n796));
  NAND2_X1  g610(.A1(new_n790), .A2(new_n796), .ZN(new_n797));
  NAND3_X1  g611(.A1(new_n776), .A2(new_n783), .A3(new_n797), .ZN(new_n798));
  INV_X1    g612(.A(KEYINPUT53), .ZN(new_n799));
  NAND2_X1  g613(.A1(new_n798), .A2(new_n799), .ZN(new_n800));
  INV_X1    g614(.A(KEYINPUT54), .ZN(new_n801));
  NAND4_X1  g615(.A1(new_n776), .A2(new_n783), .A3(KEYINPUT53), .A4(new_n797), .ZN(new_n802));
  NAND3_X1  g616(.A1(new_n800), .A2(new_n801), .A3(new_n802), .ZN(new_n803));
  NAND3_X1  g617(.A1(new_n800), .A2(KEYINPUT114), .A3(new_n802), .ZN(new_n804));
  INV_X1    g618(.A(KEYINPUT114), .ZN(new_n805));
  NAND3_X1  g619(.A1(new_n798), .A2(new_n805), .A3(new_n799), .ZN(new_n806));
  NAND2_X1  g620(.A1(new_n804), .A2(new_n806), .ZN(new_n807));
  OAI21_X1  g621(.A(new_n803), .B1(new_n807), .B2(new_n801), .ZN(new_n808));
  NOR3_X1   g622(.A1(new_n699), .A2(new_n714), .A3(new_n385), .ZN(new_n809));
  AND2_X1   g623(.A1(new_n754), .A2(new_n809), .ZN(new_n810));
  NAND2_X1  g624(.A1(new_n810), .A2(new_n723), .ZN(new_n811));
  AND2_X1   g625(.A1(new_n811), .A2(KEYINPUT119), .ZN(new_n812));
  INV_X1    g626(.A(KEYINPUT48), .ZN(new_n813));
  NAND2_X1  g627(.A1(new_n812), .A2(new_n813), .ZN(new_n814));
  NAND2_X1  g628(.A1(new_n653), .A2(new_n584), .ZN(new_n815));
  INV_X1    g629(.A(new_n809), .ZN(new_n816));
  NOR3_X1   g630(.A1(new_n815), .A2(new_n606), .A3(new_n816), .ZN(new_n817));
  NOR2_X1   g631(.A1(new_n817), .A2(new_n383), .ZN(new_n818));
  OAI21_X1  g632(.A(KEYINPUT48), .B1(new_n811), .B2(KEYINPUT119), .ZN(new_n819));
  OAI211_X1 g633(.A(new_n814), .B(new_n818), .C1(new_n819), .C2(new_n812), .ZN(new_n820));
  INV_X1    g634(.A(KEYINPUT118), .ZN(new_n821));
  NOR2_X1   g635(.A1(new_n821), .A2(KEYINPUT50), .ZN(new_n822));
  INV_X1    g636(.A(new_n694), .ZN(new_n823));
  NAND3_X1  g637(.A1(new_n754), .A2(new_n384), .A3(new_n823), .ZN(new_n824));
  AOI21_X1  g638(.A(KEYINPUT117), .B1(new_n673), .B2(new_n426), .ZN(new_n825));
  NOR2_X1   g639(.A1(new_n824), .A2(new_n825), .ZN(new_n826));
  INV_X1    g640(.A(new_n826), .ZN(new_n827));
  INV_X1    g641(.A(KEYINPUT117), .ZN(new_n828));
  NAND2_X1  g642(.A1(new_n673), .A2(new_n426), .ZN(new_n829));
  OAI21_X1  g643(.A(new_n645), .B1(new_n828), .B2(new_n829), .ZN(new_n830));
  OAI21_X1  g644(.A(new_n822), .B1(new_n827), .B2(new_n830), .ZN(new_n831));
  OR4_X1    g645(.A1(new_n824), .A2(new_n822), .A3(new_n830), .A4(new_n825), .ZN(new_n832));
  NAND2_X1  g646(.A1(new_n831), .A2(new_n832), .ZN(new_n833));
  NOR4_X1   g647(.A1(new_n815), .A2(new_n381), .A3(new_n605), .A4(new_n816), .ZN(new_n834));
  INV_X1    g648(.A(new_n834), .ZN(new_n835));
  NAND3_X1  g649(.A1(new_n810), .A2(new_n648), .A3(new_n704), .ZN(new_n836));
  AND3_X1   g650(.A1(new_n833), .A2(new_n835), .A3(new_n836), .ZN(new_n837));
  INV_X1    g651(.A(KEYINPUT51), .ZN(new_n838));
  NAND2_X1  g652(.A1(new_n670), .A2(new_n672), .ZN(new_n839));
  NOR2_X1   g653(.A1(new_n839), .A2(new_n310), .ZN(new_n840));
  OR3_X1    g654(.A1(new_n761), .A2(new_n763), .A3(new_n840), .ZN(new_n841));
  NOR2_X1   g655(.A1(new_n824), .A2(new_n757), .ZN(new_n842));
  AOI21_X1  g656(.A(new_n838), .B1(new_n841), .B2(new_n842), .ZN(new_n843));
  AOI21_X1  g657(.A(new_n820), .B1(new_n837), .B2(new_n843), .ZN(new_n844));
  NAND4_X1  g658(.A1(new_n754), .A2(new_n384), .A3(new_n700), .A4(new_n823), .ZN(new_n845));
  NAND3_X1  g659(.A1(new_n833), .A2(new_n835), .A3(new_n836), .ZN(new_n846));
  NAND3_X1  g660(.A1(new_n762), .A2(KEYINPUT115), .A3(new_n764), .ZN(new_n847));
  OR2_X1    g661(.A1(new_n840), .A2(KEYINPUT116), .ZN(new_n848));
  INV_X1    g662(.A(KEYINPUT115), .ZN(new_n849));
  OAI21_X1  g663(.A(new_n849), .B1(new_n761), .B2(new_n763), .ZN(new_n850));
  NAND2_X1  g664(.A1(new_n840), .A2(KEYINPUT116), .ZN(new_n851));
  NAND4_X1  g665(.A1(new_n847), .A2(new_n848), .A3(new_n850), .A4(new_n851), .ZN(new_n852));
  AOI21_X1  g666(.A(new_n846), .B1(new_n852), .B2(new_n842), .ZN(new_n853));
  OAI211_X1 g667(.A(new_n844), .B(new_n845), .C1(new_n853), .C2(KEYINPUT51), .ZN(new_n854));
  OAI22_X1  g668(.A1(new_n808), .A2(new_n854), .B1(G952), .B2(G953), .ZN(new_n855));
  AND3_X1   g669(.A1(new_n584), .A2(new_n425), .A3(new_n310), .ZN(new_n856));
  INV_X1    g670(.A(new_n856), .ZN(new_n857));
  AOI21_X1  g671(.A(new_n753), .B1(new_n857), .B2(KEYINPUT113), .ZN(new_n858));
  OR2_X1    g672(.A1(new_n839), .A2(KEYINPUT49), .ZN(new_n859));
  NAND2_X1  g673(.A1(new_n858), .A2(new_n859), .ZN(new_n860));
  AOI21_X1  g674(.A(new_n860), .B1(KEYINPUT49), .B2(new_n839), .ZN(new_n861));
  OR2_X1    g675(.A1(new_n857), .A2(KEYINPUT113), .ZN(new_n862));
  NAND4_X1  g676(.A1(new_n861), .A2(new_n653), .A3(new_n645), .A4(new_n862), .ZN(new_n863));
  NAND2_X1  g677(.A1(new_n855), .A2(new_n863), .ZN(new_n864));
  INV_X1    g678(.A(KEYINPUT120), .ZN(new_n865));
  NAND2_X1  g679(.A1(new_n864), .A2(new_n865), .ZN(new_n866));
  NAND3_X1  g680(.A1(new_n855), .A2(KEYINPUT120), .A3(new_n863), .ZN(new_n867));
  NAND2_X1  g681(.A1(new_n866), .A2(new_n867), .ZN(G75));
  AOI21_X1  g682(.A(new_n188), .B1(new_n800), .B2(new_n802), .ZN(new_n869));
  AOI21_X1  g683(.A(KEYINPUT56), .B1(new_n869), .B2(new_n477), .ZN(new_n870));
  NAND2_X1  g684(.A1(new_n451), .A2(new_n453), .ZN(new_n871));
  XNOR2_X1  g685(.A(new_n871), .B(new_n461), .ZN(new_n872));
  XNOR2_X1  g686(.A(new_n872), .B(KEYINPUT121), .ZN(new_n873));
  XNOR2_X1  g687(.A(new_n873), .B(KEYINPUT55), .ZN(new_n874));
  NOR2_X1   g688(.A1(KEYINPUT122), .A2(KEYINPUT56), .ZN(new_n875));
  NOR2_X1   g689(.A1(new_n874), .A2(new_n875), .ZN(new_n876));
  XNOR2_X1  g690(.A(new_n870), .B(new_n876), .ZN(new_n877));
  NOR2_X1   g691(.A1(new_n190), .A2(G952), .ZN(new_n878));
  NOR2_X1   g692(.A1(new_n877), .A2(new_n878), .ZN(G51));
  NAND2_X1  g693(.A1(new_n800), .A2(new_n802), .ZN(new_n880));
  XNOR2_X1  g694(.A(new_n880), .B(new_n801), .ZN(new_n881));
  XNOR2_X1  g695(.A(new_n299), .B(KEYINPUT57), .ZN(new_n882));
  OAI22_X1  g696(.A1(new_n881), .A2(new_n882), .B1(new_n284), .B2(new_n297), .ZN(new_n883));
  XOR2_X1   g697(.A(new_n744), .B(KEYINPUT123), .Z(new_n884));
  NAND2_X1  g698(.A1(new_n869), .A2(new_n884), .ZN(new_n885));
  AOI21_X1  g699(.A(new_n878), .B1(new_n883), .B2(new_n885), .ZN(G54));
  NAND3_X1  g700(.A1(new_n869), .A2(KEYINPUT58), .A3(G475), .ZN(new_n887));
  XOR2_X1   g701(.A(new_n887), .B(new_n371), .Z(new_n888));
  NOR2_X1   g702(.A1(new_n888), .A2(new_n878), .ZN(G60));
  NAND2_X1  g703(.A1(new_n598), .A2(new_n599), .ZN(new_n890));
  NAND2_X1  g704(.A1(G478), .A2(G902), .ZN(new_n891));
  XOR2_X1   g705(.A(new_n891), .B(KEYINPUT59), .Z(new_n892));
  OR3_X1    g706(.A1(new_n881), .A2(new_n890), .A3(new_n892), .ZN(new_n893));
  INV_X1    g707(.A(new_n878), .ZN(new_n894));
  NAND2_X1  g708(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  INV_X1    g709(.A(new_n892), .ZN(new_n896));
  NAND2_X1  g710(.A1(new_n808), .A2(new_n896), .ZN(new_n897));
  NAND2_X1  g711(.A1(new_n897), .A2(new_n890), .ZN(new_n898));
  NAND2_X1  g712(.A1(new_n898), .A2(KEYINPUT124), .ZN(new_n899));
  INV_X1    g713(.A(KEYINPUT124), .ZN(new_n900));
  NAND3_X1  g714(.A1(new_n897), .A2(new_n900), .A3(new_n890), .ZN(new_n901));
  AOI21_X1  g715(.A(new_n895), .B1(new_n899), .B2(new_n901), .ZN(G63));
  NAND2_X1  g716(.A1(G217), .A2(G902), .ZN(new_n903));
  XNOR2_X1  g717(.A(new_n903), .B(KEYINPUT60), .ZN(new_n904));
  INV_X1    g718(.A(new_n904), .ZN(new_n905));
  AND2_X1   g719(.A1(new_n790), .A2(new_n796), .ZN(new_n906));
  NAND2_X1  g720(.A1(new_n717), .A2(KEYINPUT77), .ZN(new_n907));
  NAND2_X1  g721(.A1(new_n907), .A2(new_n585), .ZN(new_n908));
  AOI21_X1  g722(.A(new_n628), .B1(new_n908), .B2(new_n483), .ZN(new_n909));
  INV_X1    g723(.A(new_n697), .ZN(new_n910));
  AND3_X1   g724(.A1(new_n910), .A2(new_n674), .A3(new_n678), .ZN(new_n911));
  NAND4_X1  g725(.A1(new_n909), .A2(new_n687), .A3(new_n911), .A4(new_n772), .ZN(new_n912));
  NOR2_X1   g726(.A1(new_n906), .A2(new_n912), .ZN(new_n913));
  AOI21_X1  g727(.A(KEYINPUT53), .B1(new_n913), .B2(new_n783), .ZN(new_n914));
  INV_X1    g728(.A(new_n802), .ZN(new_n915));
  OAI21_X1  g729(.A(new_n905), .B1(new_n914), .B2(new_n915), .ZN(new_n916));
  INV_X1    g730(.A(KEYINPUT126), .ZN(new_n917));
  NAND2_X1  g731(.A1(new_n916), .A2(new_n917), .ZN(new_n918));
  NAND2_X1  g732(.A1(new_n580), .A2(new_n582), .ZN(new_n919));
  NAND3_X1  g733(.A1(new_n880), .A2(KEYINPUT126), .A3(new_n905), .ZN(new_n920));
  NAND3_X1  g734(.A1(new_n918), .A2(new_n919), .A3(new_n920), .ZN(new_n921));
  AOI21_X1  g735(.A(KEYINPUT126), .B1(new_n880), .B2(new_n905), .ZN(new_n922));
  AOI211_X1 g736(.A(new_n917), .B(new_n904), .C1(new_n800), .C2(new_n802), .ZN(new_n923));
  OAI21_X1  g737(.A(new_n625), .B1(new_n922), .B2(new_n923), .ZN(new_n924));
  NAND3_X1  g738(.A1(new_n921), .A2(new_n924), .A3(new_n894), .ZN(new_n925));
  INV_X1    g739(.A(KEYINPUT125), .ZN(new_n926));
  XNOR2_X1  g740(.A(KEYINPUT127), .B(KEYINPUT61), .ZN(new_n927));
  AND3_X1   g741(.A1(new_n925), .A2(new_n926), .A3(new_n927), .ZN(new_n928));
  AOI21_X1  g742(.A(new_n927), .B1(new_n925), .B2(new_n926), .ZN(new_n929));
  NOR2_X1   g743(.A1(new_n928), .A2(new_n929), .ZN(G66));
  NAND2_X1  g744(.A1(new_n386), .A2(G224), .ZN(new_n931));
  NAND2_X1  g745(.A1(new_n931), .A2(G953), .ZN(new_n932));
  OAI21_X1  g746(.A(new_n932), .B1(new_n776), .B2(G953), .ZN(new_n933));
  OAI21_X1  g747(.A(new_n871), .B1(G898), .B2(new_n190), .ZN(new_n934));
  XNOR2_X1  g748(.A(new_n933), .B(new_n934), .ZN(G69));
  NOR2_X1   g749(.A1(new_n654), .A2(new_n785), .ZN(new_n936));
  XNOR2_X1  g750(.A(new_n936), .B(KEYINPUT62), .ZN(new_n937));
  NAND3_X1  g751(.A1(new_n908), .A2(new_n715), .A3(new_n770), .ZN(new_n938));
  OR2_X1    g752(.A1(new_n938), .A2(new_n641), .ZN(new_n939));
  NAND4_X1  g753(.A1(new_n937), .A2(new_n759), .A3(new_n766), .A4(new_n939), .ZN(new_n940));
  NAND2_X1  g754(.A1(new_n940), .A2(new_n190), .ZN(new_n941));
  NAND2_X1  g755(.A1(new_n507), .A2(new_n516), .ZN(new_n942));
  NAND2_X1  g756(.A1(new_n515), .A2(new_n942), .ZN(new_n943));
  XNOR2_X1  g757(.A(new_n943), .B(new_n363), .ZN(new_n944));
  INV_X1    g758(.A(new_n944), .ZN(new_n945));
  NAND2_X1  g759(.A1(new_n941), .A2(new_n945), .ZN(new_n946));
  NAND2_X1  g760(.A1(G900), .A2(G953), .ZN(new_n947));
  NAND3_X1  g761(.A1(new_n752), .A2(new_n723), .A3(new_n787), .ZN(new_n948));
  AND3_X1   g762(.A1(new_n948), .A2(new_n726), .A3(new_n734), .ZN(new_n949));
  INV_X1    g763(.A(new_n785), .ZN(new_n950));
  NAND4_X1  g764(.A1(new_n949), .A2(new_n766), .A3(new_n759), .A4(new_n950), .ZN(new_n951));
  OAI211_X1 g765(.A(new_n944), .B(new_n947), .C1(new_n951), .C2(G953), .ZN(new_n952));
  NAND2_X1  g766(.A1(new_n946), .A2(new_n952), .ZN(new_n953));
  AOI21_X1  g767(.A(new_n190), .B1(G227), .B2(G900), .ZN(new_n954));
  XNOR2_X1  g768(.A(new_n953), .B(new_n954), .ZN(G72));
  NAND2_X1  g769(.A1(G472), .A2(G902), .ZN(new_n956));
  XOR2_X1   g770(.A(new_n956), .B(KEYINPUT63), .Z(new_n957));
  OAI21_X1  g771(.A(new_n957), .B1(new_n940), .B2(new_n912), .ZN(new_n958));
  AND2_X1   g772(.A1(new_n958), .A2(new_n650), .ZN(new_n959));
  OAI21_X1  g773(.A(new_n957), .B1(new_n951), .B2(new_n912), .ZN(new_n960));
  AND3_X1   g774(.A1(new_n518), .A2(new_n506), .A3(new_n490), .ZN(new_n961));
  AND2_X1   g775(.A1(new_n960), .A2(new_n961), .ZN(new_n962));
  INV_X1    g776(.A(new_n957), .ZN(new_n963));
  NOR4_X1   g777(.A1(new_n807), .A2(new_n650), .A3(new_n963), .A4(new_n961), .ZN(new_n964));
  NOR4_X1   g778(.A1(new_n959), .A2(new_n962), .A3(new_n878), .A4(new_n964), .ZN(G57));
endmodule


