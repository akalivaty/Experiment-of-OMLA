//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 0 0 0 1 1 1 1 0 0 0 0 1 1 1 0 1 0 0 0 0 1 1 0 0 1 0 0 1 1 1 1 0 1 0 1 0 1 1 1 1 0 0 1 1 1 0 0 1 1 1 1 1 0 0 1 1 0 0 0 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:21:09 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n711, new_n712, new_n713, new_n714,
    new_n715, new_n717, new_n718, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n743, new_n744, new_n745,
    new_n747, new_n748, new_n749, new_n750, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n786, new_n787, new_n788, new_n789, new_n790, new_n791, new_n792,
    new_n793, new_n794, new_n795, new_n796, new_n797, new_n798, new_n800,
    new_n802, new_n803, new_n804, new_n805, new_n806, new_n807, new_n808,
    new_n809, new_n810, new_n811, new_n813, new_n814, new_n815, new_n816,
    new_n818, new_n819, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n877, new_n878, new_n880, new_n881, new_n882, new_n883, new_n885,
    new_n886, new_n887, new_n888, new_n889, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n939, new_n940, new_n941, new_n942,
    new_n944, new_n945, new_n946, new_n947, new_n948, new_n949, new_n950,
    new_n951, new_n952, new_n953, new_n954, new_n955, new_n956, new_n957,
    new_n958, new_n959, new_n960, new_n961, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n972, new_n973,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n982,
    new_n983, new_n984, new_n986, new_n987, new_n988, new_n990, new_n991,
    new_n992, new_n994, new_n995, new_n996, new_n997, new_n998, new_n999,
    new_n1000, new_n1002, new_n1003, new_n1004, new_n1005, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1018, new_n1019, new_n1020;
  INV_X1    g000(.A(KEYINPUT87), .ZN(new_n202));
  XNOR2_X1  g001(.A(G78gat), .B(G106gat), .ZN(new_n203));
  XNOR2_X1  g002(.A(new_n203), .B(G22gat), .ZN(new_n204));
  INV_X1    g003(.A(new_n204), .ZN(new_n205));
  INV_X1    g004(.A(G148gat), .ZN(new_n206));
  OAI21_X1  g005(.A(KEYINPUT75), .B1(new_n206), .B2(G141gat), .ZN(new_n207));
  INV_X1    g006(.A(KEYINPUT75), .ZN(new_n208));
  INV_X1    g007(.A(G141gat), .ZN(new_n209));
  NAND3_X1  g008(.A1(new_n208), .A2(new_n209), .A3(G148gat), .ZN(new_n210));
  OAI211_X1 g009(.A(new_n207), .B(new_n210), .C1(new_n209), .C2(G148gat), .ZN(new_n211));
  NAND2_X1  g010(.A1(G155gat), .A2(G162gat), .ZN(new_n212));
  INV_X1    g011(.A(G155gat), .ZN(new_n213));
  INV_X1    g012(.A(G162gat), .ZN(new_n214));
  NAND2_X1  g013(.A1(new_n213), .A2(new_n214), .ZN(new_n215));
  OAI21_X1  g014(.A(new_n212), .B1(new_n215), .B2(KEYINPUT2), .ZN(new_n216));
  NAND2_X1  g015(.A1(new_n211), .A2(new_n216), .ZN(new_n217));
  INV_X1    g016(.A(KEYINPUT2), .ZN(new_n218));
  NOR2_X1   g017(.A1(new_n206), .A2(G141gat), .ZN(new_n219));
  NOR2_X1   g018(.A1(new_n209), .A2(G148gat), .ZN(new_n220));
  OAI21_X1  g019(.A(new_n218), .B1(new_n219), .B2(new_n220), .ZN(new_n221));
  AND2_X1   g020(.A1(new_n215), .A2(new_n212), .ZN(new_n222));
  NAND2_X1  g021(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  NAND2_X1  g022(.A1(new_n217), .A2(new_n223), .ZN(new_n224));
  INV_X1    g023(.A(new_n224), .ZN(new_n225));
  INV_X1    g024(.A(KEYINPUT3), .ZN(new_n226));
  AOI21_X1  g025(.A(KEYINPUT29), .B1(new_n225), .B2(new_n226), .ZN(new_n227));
  NAND2_X1  g026(.A1(new_n227), .A2(KEYINPUT81), .ZN(new_n228));
  INV_X1    g027(.A(KEYINPUT22), .ZN(new_n229));
  XOR2_X1   g028(.A(KEYINPUT72), .B(G211gat), .Z(new_n230));
  INV_X1    g029(.A(G218gat), .ZN(new_n231));
  OAI21_X1  g030(.A(new_n229), .B1(new_n230), .B2(new_n231), .ZN(new_n232));
  XNOR2_X1  g031(.A(G197gat), .B(G204gat), .ZN(new_n233));
  XNOR2_X1  g032(.A(G211gat), .B(G218gat), .ZN(new_n234));
  NAND3_X1  g033(.A1(new_n232), .A2(new_n233), .A3(new_n234), .ZN(new_n235));
  INV_X1    g034(.A(new_n235), .ZN(new_n236));
  AOI21_X1  g035(.A(new_n234), .B1(new_n232), .B2(new_n233), .ZN(new_n237));
  NOR2_X1   g036(.A1(new_n236), .A2(new_n237), .ZN(new_n238));
  INV_X1    g037(.A(KEYINPUT29), .ZN(new_n239));
  OAI21_X1  g038(.A(new_n239), .B1(new_n224), .B2(KEYINPUT3), .ZN(new_n240));
  INV_X1    g039(.A(KEYINPUT81), .ZN(new_n241));
  NAND2_X1  g040(.A1(new_n240), .A2(new_n241), .ZN(new_n242));
  NAND3_X1  g041(.A1(new_n228), .A2(new_n238), .A3(new_n242), .ZN(new_n243));
  INV_X1    g042(.A(G228gat), .ZN(new_n244));
  INV_X1    g043(.A(G233gat), .ZN(new_n245));
  NOR2_X1   g044(.A1(new_n244), .A2(new_n245), .ZN(new_n246));
  INV_X1    g045(.A(KEYINPUT76), .ZN(new_n247));
  AOI21_X1  g046(.A(new_n247), .B1(new_n217), .B2(new_n223), .ZN(new_n248));
  INV_X1    g047(.A(new_n248), .ZN(new_n249));
  NAND3_X1  g048(.A1(new_n217), .A2(new_n223), .A3(new_n247), .ZN(new_n250));
  NAND2_X1  g049(.A1(new_n249), .A2(new_n250), .ZN(new_n251));
  OAI21_X1  g050(.A(new_n239), .B1(new_n236), .B2(new_n237), .ZN(new_n252));
  AND2_X1   g051(.A1(new_n252), .A2(new_n226), .ZN(new_n253));
  OAI211_X1 g052(.A(new_n243), .B(new_n246), .C1(new_n251), .C2(new_n253), .ZN(new_n254));
  INV_X1    g053(.A(KEYINPUT78), .ZN(new_n255));
  XNOR2_X1  g054(.A(new_n224), .B(new_n255), .ZN(new_n256));
  AOI21_X1  g055(.A(new_n256), .B1(new_n226), .B2(new_n252), .ZN(new_n257));
  INV_X1    g056(.A(new_n238), .ZN(new_n258));
  NOR2_X1   g057(.A1(new_n258), .A2(new_n227), .ZN(new_n259));
  OAI22_X1  g058(.A1(new_n257), .A2(new_n259), .B1(new_n244), .B2(new_n245), .ZN(new_n260));
  XNOR2_X1  g059(.A(KEYINPUT31), .B(G50gat), .ZN(new_n261));
  INV_X1    g060(.A(new_n261), .ZN(new_n262));
  NAND3_X1  g061(.A1(new_n254), .A2(new_n260), .A3(new_n262), .ZN(new_n263));
  INV_X1    g062(.A(new_n263), .ZN(new_n264));
  AOI21_X1  g063(.A(new_n262), .B1(new_n254), .B2(new_n260), .ZN(new_n265));
  OAI21_X1  g064(.A(new_n205), .B1(new_n264), .B2(new_n265), .ZN(new_n266));
  NAND2_X1  g065(.A1(new_n254), .A2(new_n260), .ZN(new_n267));
  NAND2_X1  g066(.A1(new_n267), .A2(new_n261), .ZN(new_n268));
  NAND3_X1  g067(.A1(new_n268), .A2(new_n204), .A3(new_n263), .ZN(new_n269));
  AND2_X1   g068(.A1(new_n266), .A2(new_n269), .ZN(new_n270));
  XNOR2_X1  g069(.A(G1gat), .B(G29gat), .ZN(new_n271));
  XNOR2_X1  g070(.A(new_n271), .B(KEYINPUT0), .ZN(new_n272));
  XNOR2_X1  g071(.A(new_n272), .B(G57gat), .ZN(new_n273));
  INV_X1    g072(.A(G85gat), .ZN(new_n274));
  XNOR2_X1  g073(.A(new_n273), .B(new_n274), .ZN(new_n275));
  INV_X1    g074(.A(new_n275), .ZN(new_n276));
  INV_X1    g075(.A(G134gat), .ZN(new_n277));
  INV_X1    g076(.A(KEYINPUT68), .ZN(new_n278));
  INV_X1    g077(.A(G127gat), .ZN(new_n279));
  INV_X1    g078(.A(KEYINPUT1), .ZN(new_n280));
  OAI21_X1  g079(.A(new_n280), .B1(G113gat), .B2(G120gat), .ZN(new_n281));
  NAND2_X1  g080(.A1(G113gat), .A2(G120gat), .ZN(new_n282));
  INV_X1    g081(.A(new_n282), .ZN(new_n283));
  OAI211_X1 g082(.A(new_n278), .B(new_n279), .C1(new_n281), .C2(new_n283), .ZN(new_n284));
  INV_X1    g083(.A(new_n284), .ZN(new_n285));
  INV_X1    g084(.A(G113gat), .ZN(new_n286));
  INV_X1    g085(.A(G120gat), .ZN(new_n287));
  NAND2_X1  g086(.A1(new_n286), .A2(new_n287), .ZN(new_n288));
  NAND3_X1  g087(.A1(new_n288), .A2(new_n280), .A3(new_n282), .ZN(new_n289));
  AOI21_X1  g088(.A(new_n279), .B1(new_n289), .B2(new_n278), .ZN(new_n290));
  OAI21_X1  g089(.A(new_n277), .B1(new_n285), .B2(new_n290), .ZN(new_n291));
  OAI21_X1  g090(.A(new_n278), .B1(new_n281), .B2(new_n283), .ZN(new_n292));
  NAND2_X1  g091(.A1(new_n292), .A2(G127gat), .ZN(new_n293));
  NAND3_X1  g092(.A1(new_n293), .A2(G134gat), .A3(new_n284), .ZN(new_n294));
  NAND2_X1  g093(.A1(new_n291), .A2(new_n294), .ZN(new_n295));
  NAND2_X1  g094(.A1(new_n295), .A2(new_n225), .ZN(new_n296));
  OAI21_X1  g095(.A(new_n296), .B1(new_n251), .B2(new_n295), .ZN(new_n297));
  NAND2_X1  g096(.A1(G225gat), .A2(G233gat), .ZN(new_n298));
  INV_X1    g097(.A(new_n298), .ZN(new_n299));
  NAND2_X1  g098(.A1(new_n297), .A2(new_n299), .ZN(new_n300));
  NAND2_X1  g099(.A1(new_n300), .A2(KEYINPUT5), .ZN(new_n301));
  INV_X1    g100(.A(new_n250), .ZN(new_n302));
  NOR3_X1   g101(.A1(new_n302), .A2(new_n226), .A3(new_n248), .ZN(new_n303));
  OAI211_X1 g102(.A(new_n291), .B(new_n294), .C1(KEYINPUT3), .C2(new_n224), .ZN(new_n304));
  OAI21_X1  g103(.A(KEYINPUT77), .B1(new_n303), .B2(new_n304), .ZN(new_n305));
  INV_X1    g104(.A(new_n304), .ZN(new_n306));
  INV_X1    g105(.A(KEYINPUT77), .ZN(new_n307));
  NAND3_X1  g106(.A1(new_n249), .A2(KEYINPUT3), .A3(new_n250), .ZN(new_n308));
  NAND3_X1  g107(.A1(new_n306), .A2(new_n307), .A3(new_n308), .ZN(new_n309));
  AOI21_X1  g108(.A(new_n299), .B1(new_n305), .B2(new_n309), .ZN(new_n310));
  XNOR2_X1  g109(.A(new_n224), .B(KEYINPUT78), .ZN(new_n311));
  INV_X1    g110(.A(new_n295), .ZN(new_n312));
  OAI21_X1  g111(.A(KEYINPUT4), .B1(new_n311), .B2(new_n312), .ZN(new_n313));
  INV_X1    g112(.A(KEYINPUT79), .ZN(new_n314));
  OAI21_X1  g113(.A(new_n314), .B1(new_n296), .B2(KEYINPUT4), .ZN(new_n315));
  AOI21_X1  g114(.A(new_n224), .B1(new_n291), .B2(new_n294), .ZN(new_n316));
  INV_X1    g115(.A(KEYINPUT4), .ZN(new_n317));
  NAND3_X1  g116(.A1(new_n316), .A2(KEYINPUT79), .A3(new_n317), .ZN(new_n318));
  NAND3_X1  g117(.A1(new_n313), .A2(new_n315), .A3(new_n318), .ZN(new_n319));
  AOI21_X1  g118(.A(new_n301), .B1(new_n310), .B2(new_n319), .ZN(new_n320));
  NAND2_X1  g119(.A1(new_n305), .A2(new_n309), .ZN(new_n321));
  NAND3_X1  g120(.A1(new_n256), .A2(new_n317), .A3(new_n295), .ZN(new_n322));
  INV_X1    g121(.A(KEYINPUT80), .ZN(new_n323));
  NAND3_X1  g122(.A1(new_n296), .A2(new_n323), .A3(KEYINPUT4), .ZN(new_n324));
  OAI21_X1  g123(.A(KEYINPUT80), .B1(new_n316), .B2(new_n317), .ZN(new_n325));
  NAND3_X1  g124(.A1(new_n322), .A2(new_n324), .A3(new_n325), .ZN(new_n326));
  NOR2_X1   g125(.A1(new_n299), .A2(KEYINPUT5), .ZN(new_n327));
  NAND3_X1  g126(.A1(new_n321), .A2(new_n326), .A3(new_n327), .ZN(new_n328));
  INV_X1    g127(.A(new_n328), .ZN(new_n329));
  OAI21_X1  g128(.A(new_n276), .B1(new_n320), .B2(new_n329), .ZN(new_n330));
  INV_X1    g129(.A(KEYINPUT5), .ZN(new_n331));
  AOI21_X1  g130(.A(new_n331), .B1(new_n297), .B2(new_n299), .ZN(new_n332));
  NOR3_X1   g131(.A1(new_n303), .A2(KEYINPUT77), .A3(new_n304), .ZN(new_n333));
  AOI21_X1  g132(.A(new_n307), .B1(new_n306), .B2(new_n308), .ZN(new_n334));
  OAI21_X1  g133(.A(new_n298), .B1(new_n333), .B2(new_n334), .ZN(new_n335));
  AND3_X1   g134(.A1(new_n313), .A2(new_n315), .A3(new_n318), .ZN(new_n336));
  OAI21_X1  g135(.A(new_n332), .B1(new_n335), .B2(new_n336), .ZN(new_n337));
  NAND3_X1  g136(.A1(new_n337), .A2(new_n275), .A3(new_n328), .ZN(new_n338));
  INV_X1    g137(.A(KEYINPUT6), .ZN(new_n339));
  NAND3_X1  g138(.A1(new_n330), .A2(new_n338), .A3(new_n339), .ZN(new_n340));
  OAI211_X1 g139(.A(KEYINPUT6), .B(new_n276), .C1(new_n320), .C2(new_n329), .ZN(new_n341));
  AND2_X1   g140(.A1(new_n340), .A2(new_n341), .ZN(new_n342));
  XNOR2_X1  g141(.A(KEYINPUT65), .B(KEYINPUT23), .ZN(new_n343));
  INV_X1    g142(.A(G169gat), .ZN(new_n344));
  INV_X1    g143(.A(G176gat), .ZN(new_n345));
  NAND2_X1  g144(.A1(new_n344), .A2(new_n345), .ZN(new_n346));
  NAND2_X1  g145(.A1(new_n343), .A2(new_n346), .ZN(new_n347));
  NAND2_X1  g146(.A1(G169gat), .A2(G176gat), .ZN(new_n348));
  INV_X1    g147(.A(KEYINPUT66), .ZN(new_n349));
  XNOR2_X1  g148(.A(new_n348), .B(new_n349), .ZN(new_n350));
  NAND3_X1  g149(.A1(new_n344), .A2(new_n345), .A3(KEYINPUT23), .ZN(new_n351));
  NAND3_X1  g150(.A1(new_n347), .A2(new_n350), .A3(new_n351), .ZN(new_n352));
  NAND2_X1  g151(.A1(G183gat), .A2(G190gat), .ZN(new_n353));
  NOR2_X1   g152(.A1(new_n353), .A2(KEYINPUT24), .ZN(new_n354));
  INV_X1    g153(.A(new_n354), .ZN(new_n355));
  XNOR2_X1  g154(.A(G183gat), .B(G190gat), .ZN(new_n356));
  INV_X1    g155(.A(KEYINPUT24), .ZN(new_n357));
  OAI21_X1  g156(.A(new_n355), .B1(new_n356), .B2(new_n357), .ZN(new_n358));
  OAI21_X1  g157(.A(KEYINPUT25), .B1(new_n352), .B2(new_n358), .ZN(new_n359));
  XNOR2_X1  g158(.A(KEYINPUT27), .B(G183gat), .ZN(new_n360));
  INV_X1    g159(.A(G190gat), .ZN(new_n361));
  NAND2_X1  g160(.A1(new_n360), .A2(new_n361), .ZN(new_n362));
  XOR2_X1   g161(.A(KEYINPUT67), .B(KEYINPUT28), .Z(new_n363));
  NAND2_X1  g162(.A1(new_n362), .A2(new_n363), .ZN(new_n364));
  INV_X1    g163(.A(new_n348), .ZN(new_n365));
  AOI21_X1  g164(.A(new_n365), .B1(KEYINPUT26), .B2(new_n346), .ZN(new_n366));
  OR3_X1    g165(.A1(KEYINPUT26), .A2(G169gat), .A3(G176gat), .ZN(new_n367));
  NAND2_X1  g166(.A1(new_n366), .A2(new_n367), .ZN(new_n368));
  NOR2_X1   g167(.A1(KEYINPUT67), .A2(KEYINPUT28), .ZN(new_n369));
  NAND3_X1  g168(.A1(new_n360), .A2(new_n361), .A3(new_n369), .ZN(new_n370));
  NAND4_X1  g169(.A1(new_n364), .A2(new_n368), .A3(new_n353), .A4(new_n370), .ZN(new_n371));
  XOR2_X1   g170(.A(G183gat), .B(G190gat), .Z(new_n372));
  AOI21_X1  g171(.A(new_n354), .B1(new_n372), .B2(KEYINPUT24), .ZN(new_n373));
  OR2_X1    g172(.A1(KEYINPUT64), .A2(G169gat), .ZN(new_n374));
  NAND2_X1  g173(.A1(KEYINPUT64), .A2(G169gat), .ZN(new_n375));
  NAND4_X1  g174(.A1(new_n374), .A2(KEYINPUT23), .A3(new_n345), .A4(new_n375), .ZN(new_n376));
  NOR2_X1   g175(.A1(new_n365), .A2(KEYINPUT25), .ZN(new_n377));
  NAND4_X1  g176(.A1(new_n373), .A2(new_n347), .A3(new_n376), .A4(new_n377), .ZN(new_n378));
  NAND3_X1  g177(.A1(new_n359), .A2(new_n371), .A3(new_n378), .ZN(new_n379));
  INV_X1    g178(.A(G226gat), .ZN(new_n380));
  NOR2_X1   g179(.A1(new_n380), .A2(new_n245), .ZN(new_n381));
  NAND2_X1  g180(.A1(new_n379), .A2(new_n381), .ZN(new_n382));
  AND2_X1   g181(.A1(new_n370), .A2(new_n353), .ZN(new_n383));
  AOI22_X1  g182(.A1(new_n362), .A2(new_n363), .B1(new_n366), .B2(new_n367), .ZN(new_n384));
  AND3_X1   g183(.A1(new_n347), .A2(new_n376), .A3(new_n377), .ZN(new_n385));
  AOI22_X1  g184(.A1(new_n383), .A2(new_n384), .B1(new_n385), .B2(new_n373), .ZN(new_n386));
  AOI21_X1  g185(.A(KEYINPUT29), .B1(new_n386), .B2(new_n359), .ZN(new_n387));
  OAI211_X1 g186(.A(new_n258), .B(new_n382), .C1(new_n387), .C2(new_n381), .ZN(new_n388));
  AOI21_X1  g187(.A(new_n381), .B1(new_n379), .B2(new_n239), .ZN(new_n389));
  INV_X1    g188(.A(new_n381), .ZN(new_n390));
  AOI21_X1  g189(.A(new_n390), .B1(new_n386), .B2(new_n359), .ZN(new_n391));
  OAI21_X1  g190(.A(new_n238), .B1(new_n389), .B2(new_n391), .ZN(new_n392));
  INV_X1    g191(.A(KEYINPUT73), .ZN(new_n393));
  NAND3_X1  g192(.A1(new_n388), .A2(new_n392), .A3(new_n393), .ZN(new_n394));
  INV_X1    g193(.A(new_n389), .ZN(new_n395));
  NAND4_X1  g194(.A1(new_n395), .A2(KEYINPUT73), .A3(new_n258), .A4(new_n382), .ZN(new_n396));
  XNOR2_X1  g195(.A(G8gat), .B(G36gat), .ZN(new_n397));
  XNOR2_X1  g196(.A(new_n397), .B(G64gat), .ZN(new_n398));
  INV_X1    g197(.A(G92gat), .ZN(new_n399));
  XNOR2_X1  g198(.A(new_n398), .B(new_n399), .ZN(new_n400));
  INV_X1    g199(.A(new_n400), .ZN(new_n401));
  AND3_X1   g200(.A1(new_n394), .A2(new_n396), .A3(new_n401), .ZN(new_n402));
  NAND2_X1  g201(.A1(new_n394), .A2(new_n396), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n403), .A2(new_n400), .ZN(new_n404));
  INV_X1    g203(.A(KEYINPUT30), .ZN(new_n405));
  AOI21_X1  g204(.A(new_n402), .B1(new_n404), .B2(new_n405), .ZN(new_n406));
  AOI21_X1  g205(.A(new_n401), .B1(new_n394), .B2(new_n396), .ZN(new_n407));
  NAND3_X1  g206(.A1(new_n407), .A2(KEYINPUT74), .A3(KEYINPUT30), .ZN(new_n408));
  INV_X1    g207(.A(new_n408), .ZN(new_n409));
  AOI21_X1  g208(.A(KEYINPUT74), .B1(new_n407), .B2(KEYINPUT30), .ZN(new_n410));
  OAI21_X1  g209(.A(new_n406), .B1(new_n409), .B2(new_n410), .ZN(new_n411));
  OAI21_X1  g210(.A(new_n270), .B1(new_n342), .B2(new_n411), .ZN(new_n412));
  NAND3_X1  g211(.A1(new_n312), .A2(new_n359), .A3(new_n386), .ZN(new_n413));
  INV_X1    g212(.A(G227gat), .ZN(new_n414));
  NOR2_X1   g213(.A1(new_n414), .A2(new_n245), .ZN(new_n415));
  NAND2_X1  g214(.A1(new_n379), .A2(new_n295), .ZN(new_n416));
  NAND3_X1  g215(.A1(new_n413), .A2(new_n415), .A3(new_n416), .ZN(new_n417));
  INV_X1    g216(.A(KEYINPUT32), .ZN(new_n418));
  XNOR2_X1  g217(.A(G15gat), .B(G43gat), .ZN(new_n419));
  XNOR2_X1  g218(.A(G71gat), .B(G99gat), .ZN(new_n420));
  XNOR2_X1  g219(.A(new_n419), .B(new_n420), .ZN(new_n421));
  INV_X1    g220(.A(new_n421), .ZN(new_n422));
  AOI21_X1  g221(.A(new_n418), .B1(new_n422), .B2(KEYINPUT33), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n417), .A2(new_n423), .ZN(new_n424));
  INV_X1    g223(.A(KEYINPUT69), .ZN(new_n425));
  NAND2_X1  g224(.A1(new_n418), .A2(KEYINPUT33), .ZN(new_n426));
  NAND2_X1  g225(.A1(new_n417), .A2(new_n426), .ZN(new_n427));
  AOI21_X1  g226(.A(new_n425), .B1(new_n427), .B2(new_n422), .ZN(new_n428));
  AOI211_X1 g227(.A(KEYINPUT69), .B(new_n421), .C1(new_n417), .C2(new_n426), .ZN(new_n429));
  OAI21_X1  g228(.A(new_n424), .B1(new_n428), .B2(new_n429), .ZN(new_n430));
  INV_X1    g229(.A(KEYINPUT71), .ZN(new_n431));
  NAND2_X1  g230(.A1(new_n430), .A2(new_n431), .ZN(new_n432));
  OAI211_X1 g231(.A(KEYINPUT71), .B(new_n424), .C1(new_n428), .C2(new_n429), .ZN(new_n433));
  NAND2_X1  g232(.A1(new_n413), .A2(new_n416), .ZN(new_n434));
  INV_X1    g233(.A(new_n415), .ZN(new_n435));
  NAND2_X1  g234(.A1(new_n434), .A2(new_n435), .ZN(new_n436));
  XOR2_X1   g235(.A(KEYINPUT70), .B(KEYINPUT34), .Z(new_n437));
  XNOR2_X1  g236(.A(new_n436), .B(new_n437), .ZN(new_n438));
  NAND3_X1  g237(.A1(new_n432), .A2(new_n433), .A3(new_n438), .ZN(new_n439));
  OR2_X1    g238(.A1(new_n433), .A2(new_n438), .ZN(new_n440));
  NAND3_X1  g239(.A1(new_n439), .A2(KEYINPUT36), .A3(new_n440), .ZN(new_n441));
  NAND2_X1  g240(.A1(new_n439), .A2(new_n440), .ZN(new_n442));
  INV_X1    g241(.A(KEYINPUT36), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  NAND3_X1  g243(.A1(new_n412), .A2(new_n441), .A3(new_n444), .ZN(new_n445));
  INV_X1    g244(.A(KEYINPUT82), .ZN(new_n446));
  NAND2_X1  g245(.A1(new_n411), .A2(new_n446), .ZN(new_n447));
  INV_X1    g246(.A(KEYINPUT74), .ZN(new_n448));
  OAI21_X1  g247(.A(new_n448), .B1(new_n404), .B2(new_n405), .ZN(new_n449));
  NAND2_X1  g248(.A1(new_n449), .A2(new_n408), .ZN(new_n450));
  NAND3_X1  g249(.A1(new_n450), .A2(KEYINPUT82), .A3(new_n406), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n447), .A2(new_n451), .ZN(new_n452));
  AOI21_X1  g251(.A(new_n298), .B1(new_n321), .B2(new_n326), .ZN(new_n453));
  INV_X1    g252(.A(KEYINPUT39), .ZN(new_n454));
  NAND2_X1  g253(.A1(new_n453), .A2(new_n454), .ZN(new_n455));
  OAI211_X1 g254(.A(new_n296), .B(new_n298), .C1(new_n251), .C2(new_n295), .ZN(new_n456));
  NAND2_X1  g255(.A1(new_n456), .A2(KEYINPUT39), .ZN(new_n457));
  INV_X1    g256(.A(KEYINPUT83), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  NAND3_X1  g258(.A1(new_n456), .A2(KEYINPUT83), .A3(KEYINPUT39), .ZN(new_n460));
  NAND2_X1  g259(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  OAI211_X1 g260(.A(new_n455), .B(new_n275), .C1(new_n453), .C2(new_n461), .ZN(new_n462));
  INV_X1    g261(.A(KEYINPUT40), .ZN(new_n463));
  OAI21_X1  g262(.A(new_n330), .B1(new_n462), .B2(new_n463), .ZN(new_n464));
  OAI21_X1  g263(.A(new_n275), .B1(new_n461), .B2(new_n453), .ZN(new_n465));
  INV_X1    g264(.A(new_n455), .ZN(new_n466));
  OAI21_X1  g265(.A(new_n463), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  INV_X1    g266(.A(KEYINPUT84), .ZN(new_n468));
  NAND2_X1  g267(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  NAND3_X1  g268(.A1(new_n462), .A2(KEYINPUT84), .A3(new_n463), .ZN(new_n470));
  AOI21_X1  g269(.A(new_n464), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  AOI21_X1  g270(.A(new_n270), .B1(new_n452), .B2(new_n471), .ZN(new_n472));
  INV_X1    g271(.A(KEYINPUT37), .ZN(new_n473));
  NAND2_X1  g272(.A1(new_n403), .A2(new_n473), .ZN(new_n474));
  NAND2_X1  g273(.A1(new_n474), .A2(KEYINPUT85), .ZN(new_n475));
  INV_X1    g274(.A(KEYINPUT85), .ZN(new_n476));
  NAND3_X1  g275(.A1(new_n403), .A2(new_n476), .A3(new_n473), .ZN(new_n477));
  NAND3_X1  g276(.A1(new_n475), .A2(new_n477), .A3(new_n401), .ZN(new_n478));
  AOI21_X1  g277(.A(new_n473), .B1(new_n388), .B2(new_n392), .ZN(new_n479));
  OR2_X1    g278(.A1(new_n479), .A2(KEYINPUT38), .ZN(new_n480));
  OR2_X1    g279(.A1(new_n478), .A2(new_n480), .ZN(new_n481));
  NOR2_X1   g280(.A1(new_n403), .A2(new_n473), .ZN(new_n482));
  OAI21_X1  g281(.A(KEYINPUT38), .B1(new_n478), .B2(new_n482), .ZN(new_n483));
  NAND4_X1  g282(.A1(new_n481), .A2(new_n483), .A3(new_n342), .A4(new_n404), .ZN(new_n484));
  AOI21_X1  g283(.A(new_n445), .B1(new_n472), .B2(new_n484), .ZN(new_n485));
  NAND2_X1  g284(.A1(new_n340), .A2(new_n341), .ZN(new_n486));
  NAND3_X1  g285(.A1(new_n394), .A2(new_n396), .A3(new_n401), .ZN(new_n487));
  OAI21_X1  g286(.A(new_n487), .B1(new_n407), .B2(KEYINPUT30), .ZN(new_n488));
  AOI21_X1  g287(.A(new_n488), .B1(new_n449), .B2(new_n408), .ZN(new_n489));
  NAND2_X1  g288(.A1(new_n266), .A2(new_n269), .ZN(new_n490));
  NAND4_X1  g289(.A1(new_n442), .A2(new_n486), .A3(new_n489), .A4(new_n490), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n491), .A2(KEYINPUT35), .ZN(new_n492));
  AOI21_X1  g291(.A(new_n270), .B1(new_n439), .B2(new_n440), .ZN(new_n493));
  XNOR2_X1  g292(.A(KEYINPUT86), .B(KEYINPUT35), .ZN(new_n494));
  AOI21_X1  g293(.A(new_n494), .B1(new_n340), .B2(new_n341), .ZN(new_n495));
  NAND4_X1  g294(.A1(new_n493), .A2(new_n447), .A3(new_n451), .A4(new_n495), .ZN(new_n496));
  AND2_X1   g295(.A1(new_n492), .A2(new_n496), .ZN(new_n497));
  OAI21_X1  g296(.A(new_n202), .B1(new_n485), .B2(new_n497), .ZN(new_n498));
  NOR2_X1   g297(.A1(new_n411), .A2(new_n446), .ZN(new_n499));
  AOI21_X1  g298(.A(KEYINPUT82), .B1(new_n450), .B2(new_n406), .ZN(new_n500));
  OAI21_X1  g299(.A(new_n471), .B1(new_n499), .B2(new_n500), .ZN(new_n501));
  NAND3_X1  g300(.A1(new_n501), .A2(new_n484), .A3(new_n490), .ZN(new_n502));
  AND3_X1   g301(.A1(new_n412), .A2(new_n441), .A3(new_n444), .ZN(new_n503));
  NAND2_X1  g302(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  NAND2_X1  g303(.A1(new_n492), .A2(new_n496), .ZN(new_n505));
  NAND3_X1  g304(.A1(new_n504), .A2(KEYINPUT87), .A3(new_n505), .ZN(new_n506));
  XNOR2_X1  g305(.A(G113gat), .B(G141gat), .ZN(new_n507));
  XNOR2_X1  g306(.A(new_n507), .B(KEYINPUT11), .ZN(new_n508));
  NAND2_X1  g307(.A1(new_n508), .A2(G169gat), .ZN(new_n509));
  OR2_X1    g308(.A1(new_n507), .A2(KEYINPUT11), .ZN(new_n510));
  NAND2_X1  g309(.A1(new_n507), .A2(KEYINPUT11), .ZN(new_n511));
  NAND3_X1  g310(.A1(new_n510), .A2(new_n344), .A3(new_n511), .ZN(new_n512));
  AOI21_X1  g311(.A(G197gat), .B1(new_n509), .B2(new_n512), .ZN(new_n513));
  INV_X1    g312(.A(new_n513), .ZN(new_n514));
  NAND3_X1  g313(.A1(new_n509), .A2(G197gat), .A3(new_n512), .ZN(new_n515));
  AND3_X1   g314(.A1(new_n514), .A2(KEYINPUT12), .A3(new_n515), .ZN(new_n516));
  AOI21_X1  g315(.A(KEYINPUT12), .B1(new_n514), .B2(new_n515), .ZN(new_n517));
  NOR2_X1   g316(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  INV_X1    g317(.A(new_n518), .ZN(new_n519));
  INV_X1    g318(.A(KEYINPUT90), .ZN(new_n520));
  AND2_X1   g319(.A1(G43gat), .A2(G50gat), .ZN(new_n521));
  NOR2_X1   g320(.A1(G43gat), .A2(G50gat), .ZN(new_n522));
  OAI21_X1  g321(.A(KEYINPUT15), .B1(new_n521), .B2(new_n522), .ZN(new_n523));
  INV_X1    g322(.A(G43gat), .ZN(new_n524));
  INV_X1    g323(.A(G50gat), .ZN(new_n525));
  NAND2_X1  g324(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  INV_X1    g325(.A(KEYINPUT15), .ZN(new_n527));
  NAND2_X1  g326(.A1(G43gat), .A2(G50gat), .ZN(new_n528));
  NAND3_X1  g327(.A1(new_n526), .A2(new_n527), .A3(new_n528), .ZN(new_n529));
  NAND2_X1  g328(.A1(G29gat), .A2(G36gat), .ZN(new_n530));
  AND3_X1   g329(.A1(new_n523), .A2(new_n529), .A3(new_n530), .ZN(new_n531));
  OAI21_X1  g330(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n532));
  INV_X1    g331(.A(KEYINPUT88), .ZN(new_n533));
  NAND2_X1  g332(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  OAI211_X1 g333(.A(KEYINPUT88), .B(KEYINPUT14), .C1(G29gat), .C2(G36gat), .ZN(new_n535));
  NAND2_X1  g334(.A1(new_n534), .A2(new_n535), .ZN(new_n536));
  INV_X1    g335(.A(KEYINPUT14), .ZN(new_n537));
  INV_X1    g336(.A(G29gat), .ZN(new_n538));
  INV_X1    g337(.A(G36gat), .ZN(new_n539));
  NAND3_X1  g338(.A1(new_n537), .A2(new_n538), .A3(new_n539), .ZN(new_n540));
  NAND2_X1  g339(.A1(new_n536), .A2(new_n540), .ZN(new_n541));
  AOI21_X1  g340(.A(new_n520), .B1(new_n531), .B2(new_n541), .ZN(new_n542));
  NAND3_X1  g341(.A1(new_n523), .A2(new_n529), .A3(new_n530), .ZN(new_n543));
  NOR3_X1   g342(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n544));
  AOI21_X1  g343(.A(new_n544), .B1(new_n534), .B2(new_n535), .ZN(new_n545));
  NOR3_X1   g344(.A1(new_n543), .A2(new_n545), .A3(KEYINPUT90), .ZN(new_n546));
  NOR4_X1   g345(.A1(KEYINPUT89), .A2(KEYINPUT14), .A3(G29gat), .A4(G36gat), .ZN(new_n547));
  INV_X1    g346(.A(KEYINPUT89), .ZN(new_n548));
  NOR2_X1   g347(.A1(KEYINPUT14), .A2(G29gat), .ZN(new_n549));
  AOI21_X1  g348(.A(new_n548), .B1(new_n549), .B2(new_n539), .ZN(new_n550));
  NOR2_X1   g349(.A1(new_n547), .A2(new_n550), .ZN(new_n551));
  AOI22_X1  g350(.A1(new_n551), .A2(new_n536), .B1(G29gat), .B2(G36gat), .ZN(new_n552));
  OAI22_X1  g351(.A1(new_n542), .A2(new_n546), .B1(new_n523), .B2(new_n552), .ZN(new_n553));
  XNOR2_X1  g352(.A(G15gat), .B(G22gat), .ZN(new_n554));
  INV_X1    g353(.A(G1gat), .ZN(new_n555));
  NAND2_X1  g354(.A1(new_n555), .A2(KEYINPUT16), .ZN(new_n556));
  NAND2_X1  g355(.A1(new_n554), .A2(new_n556), .ZN(new_n557));
  OAI21_X1  g356(.A(new_n557), .B1(G1gat), .B2(new_n554), .ZN(new_n558));
  NAND2_X1  g357(.A1(new_n558), .A2(G8gat), .ZN(new_n559));
  INV_X1    g358(.A(G8gat), .ZN(new_n560));
  OAI211_X1 g359(.A(new_n557), .B(new_n560), .C1(G1gat), .C2(new_n554), .ZN(new_n561));
  NAND2_X1  g360(.A1(new_n559), .A2(new_n561), .ZN(new_n562));
  NAND2_X1  g361(.A1(new_n553), .A2(new_n562), .ZN(new_n563));
  NAND3_X1  g362(.A1(new_n531), .A2(new_n520), .A3(new_n541), .ZN(new_n564));
  OAI21_X1  g363(.A(KEYINPUT90), .B1(new_n543), .B2(new_n545), .ZN(new_n565));
  AND2_X1   g364(.A1(new_n534), .A2(new_n535), .ZN(new_n566));
  NAND2_X1  g365(.A1(new_n540), .A2(KEYINPUT89), .ZN(new_n567));
  NAND3_X1  g366(.A1(new_n549), .A2(new_n548), .A3(new_n539), .ZN(new_n568));
  NAND2_X1  g367(.A1(new_n567), .A2(new_n568), .ZN(new_n569));
  OAI21_X1  g368(.A(new_n530), .B1(new_n566), .B2(new_n569), .ZN(new_n570));
  INV_X1    g369(.A(new_n523), .ZN(new_n571));
  AOI22_X1  g370(.A1(new_n564), .A2(new_n565), .B1(new_n570), .B2(new_n571), .ZN(new_n572));
  INV_X1    g371(.A(new_n562), .ZN(new_n573));
  NAND2_X1  g372(.A1(new_n572), .A2(new_n573), .ZN(new_n574));
  NAND2_X1  g373(.A1(new_n563), .A2(new_n574), .ZN(new_n575));
  NAND2_X1  g374(.A1(G229gat), .A2(G233gat), .ZN(new_n576));
  XOR2_X1   g375(.A(new_n576), .B(KEYINPUT13), .Z(new_n577));
  NAND2_X1  g376(.A1(new_n575), .A2(new_n577), .ZN(new_n578));
  OAI21_X1  g377(.A(new_n573), .B1(new_n572), .B2(KEYINPUT17), .ZN(new_n579));
  NAND2_X1  g378(.A1(new_n564), .A2(new_n565), .ZN(new_n580));
  NAND2_X1  g379(.A1(new_n570), .A2(new_n571), .ZN(new_n581));
  AND3_X1   g380(.A1(new_n580), .A2(KEYINPUT17), .A3(new_n581), .ZN(new_n582));
  OAI211_X1 g381(.A(new_n576), .B(new_n563), .C1(new_n579), .C2(new_n582), .ZN(new_n583));
  INV_X1    g382(.A(KEYINPUT18), .ZN(new_n584));
  OAI21_X1  g383(.A(new_n578), .B1(new_n583), .B2(new_n584), .ZN(new_n585));
  XNOR2_X1  g384(.A(KEYINPUT91), .B(KEYINPUT18), .ZN(new_n586));
  INV_X1    g385(.A(new_n586), .ZN(new_n587));
  NOR2_X1   g386(.A1(new_n572), .A2(new_n573), .ZN(new_n588));
  INV_X1    g387(.A(KEYINPUT17), .ZN(new_n589));
  AOI21_X1  g388(.A(new_n562), .B1(new_n553), .B2(new_n589), .ZN(new_n590));
  NAND3_X1  g389(.A1(new_n580), .A2(KEYINPUT17), .A3(new_n581), .ZN(new_n591));
  AOI21_X1  g390(.A(new_n588), .B1(new_n590), .B2(new_n591), .ZN(new_n592));
  AOI21_X1  g391(.A(new_n587), .B1(new_n592), .B2(new_n576), .ZN(new_n593));
  OAI21_X1  g392(.A(new_n519), .B1(new_n585), .B2(new_n593), .ZN(new_n594));
  NAND2_X1  g393(.A1(new_n583), .A2(new_n586), .ZN(new_n595));
  NAND2_X1  g394(.A1(new_n553), .A2(new_n589), .ZN(new_n596));
  NAND3_X1  g395(.A1(new_n596), .A2(new_n573), .A3(new_n591), .ZN(new_n597));
  NAND4_X1  g396(.A1(new_n597), .A2(KEYINPUT18), .A3(new_n576), .A4(new_n563), .ZN(new_n598));
  NAND4_X1  g397(.A1(new_n595), .A2(new_n518), .A3(new_n598), .A4(new_n578), .ZN(new_n599));
  NAND2_X1  g398(.A1(new_n594), .A2(new_n599), .ZN(new_n600));
  INV_X1    g399(.A(KEYINPUT92), .ZN(new_n601));
  NAND2_X1  g400(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  NAND3_X1  g401(.A1(new_n594), .A2(KEYINPUT92), .A3(new_n599), .ZN(new_n603));
  NAND2_X1  g402(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  OR2_X1    g403(.A1(G57gat), .A2(G64gat), .ZN(new_n605));
  NAND2_X1  g404(.A1(G57gat), .A2(G64gat), .ZN(new_n606));
  AND2_X1   g405(.A1(new_n605), .A2(new_n606), .ZN(new_n607));
  NAND2_X1  g406(.A1(G71gat), .A2(G78gat), .ZN(new_n608));
  INV_X1    g407(.A(KEYINPUT9), .ZN(new_n609));
  NAND2_X1  g408(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  INV_X1    g409(.A(KEYINPUT95), .ZN(new_n611));
  NAND2_X1  g410(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  NOR2_X1   g411(.A1(G71gat), .A2(G78gat), .ZN(new_n613));
  INV_X1    g412(.A(new_n613), .ZN(new_n614));
  NAND2_X1  g413(.A1(new_n614), .A2(new_n608), .ZN(new_n615));
  NAND3_X1  g414(.A1(new_n608), .A2(KEYINPUT95), .A3(new_n609), .ZN(new_n616));
  NAND4_X1  g415(.A1(new_n607), .A2(new_n612), .A3(new_n615), .A4(new_n616), .ZN(new_n617));
  NAND3_X1  g416(.A1(new_n610), .A2(new_n605), .A3(new_n606), .ZN(new_n618));
  NAND2_X1  g417(.A1(new_n608), .A2(KEYINPUT93), .ZN(new_n619));
  INV_X1    g418(.A(KEYINPUT93), .ZN(new_n620));
  NAND3_X1  g419(.A1(new_n620), .A2(G71gat), .A3(G78gat), .ZN(new_n621));
  AOI21_X1  g420(.A(new_n613), .B1(new_n619), .B2(new_n621), .ZN(new_n622));
  INV_X1    g421(.A(KEYINPUT94), .ZN(new_n623));
  OAI21_X1  g422(.A(new_n618), .B1(new_n622), .B2(new_n623), .ZN(new_n624));
  AOI211_X1 g423(.A(KEYINPUT94), .B(new_n613), .C1(new_n619), .C2(new_n621), .ZN(new_n625));
  OAI21_X1  g424(.A(new_n617), .B1(new_n624), .B2(new_n625), .ZN(new_n626));
  NAND2_X1  g425(.A1(new_n626), .A2(KEYINPUT96), .ZN(new_n627));
  INV_X1    g426(.A(KEYINPUT96), .ZN(new_n628));
  OAI211_X1 g427(.A(new_n628), .B(new_n617), .C1(new_n624), .C2(new_n625), .ZN(new_n629));
  NAND2_X1  g428(.A1(new_n627), .A2(new_n629), .ZN(new_n630));
  INV_X1    g429(.A(KEYINPUT21), .ZN(new_n631));
  OAI21_X1  g430(.A(new_n573), .B1(new_n630), .B2(new_n631), .ZN(new_n632));
  XNOR2_X1  g431(.A(new_n632), .B(G183gat), .ZN(new_n633));
  XNOR2_X1  g432(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n634));
  NAND2_X1  g433(.A1(G231gat), .A2(G233gat), .ZN(new_n635));
  XNOR2_X1  g434(.A(new_n634), .B(new_n635), .ZN(new_n636));
  XNOR2_X1  g435(.A(new_n633), .B(new_n636), .ZN(new_n637));
  NAND2_X1  g436(.A1(new_n630), .A2(new_n631), .ZN(new_n638));
  XOR2_X1   g437(.A(G127gat), .B(G155gat), .Z(new_n639));
  XNOR2_X1  g438(.A(new_n638), .B(new_n639), .ZN(new_n640));
  XNOR2_X1  g439(.A(new_n640), .B(G211gat), .ZN(new_n641));
  OR2_X1    g440(.A1(new_n637), .A2(new_n641), .ZN(new_n642));
  NAND2_X1  g441(.A1(new_n637), .A2(new_n641), .ZN(new_n643));
  NAND2_X1  g442(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  NAND2_X1  g443(.A1(G85gat), .A2(G92gat), .ZN(new_n645));
  XNOR2_X1  g444(.A(new_n645), .B(KEYINPUT7), .ZN(new_n646));
  NAND2_X1  g445(.A1(G99gat), .A2(G106gat), .ZN(new_n647));
  AOI22_X1  g446(.A1(KEYINPUT8), .A2(new_n647), .B1(new_n274), .B2(new_n399), .ZN(new_n648));
  NAND2_X1  g447(.A1(new_n646), .A2(new_n648), .ZN(new_n649));
  XNOR2_X1  g448(.A(G99gat), .B(G106gat), .ZN(new_n650));
  XNOR2_X1  g449(.A(new_n649), .B(new_n650), .ZN(new_n651));
  INV_X1    g450(.A(new_n651), .ZN(new_n652));
  NAND3_X1  g451(.A1(new_n596), .A2(new_n591), .A3(new_n652), .ZN(new_n653));
  AND2_X1   g452(.A1(G232gat), .A2(G233gat), .ZN(new_n654));
  AOI22_X1  g453(.A1(new_n553), .A2(new_n651), .B1(KEYINPUT41), .B2(new_n654), .ZN(new_n655));
  NAND2_X1  g454(.A1(new_n653), .A2(new_n655), .ZN(new_n656));
  XOR2_X1   g455(.A(G134gat), .B(G162gat), .Z(new_n657));
  XNOR2_X1  g456(.A(new_n656), .B(new_n657), .ZN(new_n658));
  NOR2_X1   g457(.A1(new_n654), .A2(KEYINPUT41), .ZN(new_n659));
  XNOR2_X1  g458(.A(G190gat), .B(G218gat), .ZN(new_n660));
  XNOR2_X1  g459(.A(new_n659), .B(new_n660), .ZN(new_n661));
  XNOR2_X1  g460(.A(new_n658), .B(new_n661), .ZN(new_n662));
  INV_X1    g461(.A(new_n662), .ZN(new_n663));
  XNOR2_X1  g462(.A(G120gat), .B(G148gat), .ZN(new_n664));
  XNOR2_X1  g463(.A(new_n664), .B(G176gat), .ZN(new_n665));
  XOR2_X1   g464(.A(new_n665), .B(G204gat), .Z(new_n666));
  INV_X1    g465(.A(new_n666), .ZN(new_n667));
  INV_X1    g466(.A(G230gat), .ZN(new_n668));
  NOR2_X1   g467(.A1(new_n668), .A2(new_n245), .ZN(new_n669));
  AND2_X1   g468(.A1(new_n619), .A2(new_n621), .ZN(new_n670));
  OAI21_X1  g469(.A(KEYINPUT94), .B1(new_n670), .B2(new_n613), .ZN(new_n671));
  NAND2_X1  g470(.A1(new_n622), .A2(new_n623), .ZN(new_n672));
  NAND3_X1  g471(.A1(new_n671), .A2(new_n672), .A3(new_n618), .ZN(new_n673));
  AOI21_X1  g472(.A(new_n628), .B1(new_n673), .B2(new_n617), .ZN(new_n674));
  INV_X1    g473(.A(new_n629), .ZN(new_n675));
  OAI21_X1  g474(.A(new_n652), .B1(new_n674), .B2(new_n675), .ZN(new_n676));
  INV_X1    g475(.A(KEYINPUT10), .ZN(new_n677));
  NOR2_X1   g476(.A1(new_n650), .A2(KEYINPUT97), .ZN(new_n678));
  AND2_X1   g477(.A1(new_n649), .A2(new_n678), .ZN(new_n679));
  NOR2_X1   g478(.A1(new_n649), .A2(new_n678), .ZN(new_n680));
  NOR3_X1   g479(.A1(new_n626), .A2(new_n679), .A3(new_n680), .ZN(new_n681));
  INV_X1    g480(.A(new_n681), .ZN(new_n682));
  NAND3_X1  g481(.A1(new_n676), .A2(new_n677), .A3(new_n682), .ZN(new_n683));
  NAND4_X1  g482(.A1(new_n627), .A2(KEYINPUT10), .A3(new_n629), .A4(new_n651), .ZN(new_n684));
  AOI21_X1  g483(.A(new_n669), .B1(new_n683), .B2(new_n684), .ZN(new_n685));
  AOI21_X1  g484(.A(new_n651), .B1(new_n627), .B2(new_n629), .ZN(new_n686));
  OAI21_X1  g485(.A(new_n669), .B1(new_n686), .B2(new_n681), .ZN(new_n687));
  INV_X1    g486(.A(new_n687), .ZN(new_n688));
  OAI21_X1  g487(.A(new_n667), .B1(new_n685), .B2(new_n688), .ZN(new_n689));
  INV_X1    g488(.A(new_n684), .ZN(new_n690));
  AOI21_X1  g489(.A(new_n681), .B1(new_n630), .B2(new_n652), .ZN(new_n691));
  AOI21_X1  g490(.A(new_n690), .B1(new_n691), .B2(new_n677), .ZN(new_n692));
  OAI211_X1 g491(.A(new_n687), .B(new_n666), .C1(new_n692), .C2(new_n669), .ZN(new_n693));
  NAND3_X1  g492(.A1(new_n689), .A2(KEYINPUT98), .A3(new_n693), .ZN(new_n694));
  INV_X1    g493(.A(KEYINPUT98), .ZN(new_n695));
  OAI211_X1 g494(.A(new_n695), .B(new_n667), .C1(new_n685), .C2(new_n688), .ZN(new_n696));
  NAND2_X1  g495(.A1(new_n694), .A2(new_n696), .ZN(new_n697));
  NAND3_X1  g496(.A1(new_n644), .A2(new_n663), .A3(new_n697), .ZN(new_n698));
  INV_X1    g497(.A(new_n698), .ZN(new_n699));
  NAND4_X1  g498(.A1(new_n498), .A2(new_n506), .A3(new_n604), .A4(new_n699), .ZN(new_n700));
  NOR2_X1   g499(.A1(new_n700), .A2(new_n486), .ZN(new_n701));
  XNOR2_X1  g500(.A(new_n701), .B(new_n555), .ZN(G1324gat));
  INV_X1    g501(.A(new_n452), .ZN(new_n703));
  NOR2_X1   g502(.A1(new_n700), .A2(new_n703), .ZN(new_n704));
  NOR2_X1   g503(.A1(new_n704), .A2(new_n560), .ZN(new_n705));
  INV_X1    g504(.A(KEYINPUT42), .ZN(new_n706));
  XOR2_X1   g505(.A(KEYINPUT16), .B(G8gat), .Z(new_n707));
  NAND2_X1  g506(.A1(new_n704), .A2(new_n707), .ZN(new_n708));
  AOI21_X1  g507(.A(new_n705), .B1(new_n706), .B2(new_n708), .ZN(new_n709));
  OAI21_X1  g508(.A(new_n709), .B1(new_n706), .B2(new_n708), .ZN(G1325gat));
  NAND2_X1  g509(.A1(new_n444), .A2(new_n441), .ZN(new_n711));
  INV_X1    g510(.A(new_n711), .ZN(new_n712));
  OAI21_X1  g511(.A(G15gat), .B1(new_n700), .B2(new_n712), .ZN(new_n713));
  INV_X1    g512(.A(new_n442), .ZN(new_n714));
  OR2_X1    g513(.A1(new_n714), .A2(G15gat), .ZN(new_n715));
  OAI21_X1  g514(.A(new_n713), .B1(new_n700), .B2(new_n715), .ZN(G1326gat));
  NOR2_X1   g515(.A1(new_n700), .A2(new_n490), .ZN(new_n717));
  XOR2_X1   g516(.A(KEYINPUT43), .B(G22gat), .Z(new_n718));
  XNOR2_X1  g517(.A(new_n717), .B(new_n718), .ZN(G1327gat));
  INV_X1    g518(.A(new_n697), .ZN(new_n720));
  NOR2_X1   g519(.A1(new_n644), .A2(new_n720), .ZN(new_n721));
  NAND2_X1  g520(.A1(new_n721), .A2(new_n662), .ZN(new_n722));
  XNOR2_X1  g521(.A(new_n722), .B(KEYINPUT99), .ZN(new_n723));
  NAND4_X1  g522(.A1(new_n498), .A2(new_n506), .A3(new_n604), .A4(new_n723), .ZN(new_n724));
  INV_X1    g523(.A(new_n724), .ZN(new_n725));
  NAND3_X1  g524(.A1(new_n725), .A2(new_n538), .A3(new_n342), .ZN(new_n726));
  XNOR2_X1  g525(.A(new_n726), .B(KEYINPUT45), .ZN(new_n727));
  NAND3_X1  g526(.A1(new_n498), .A2(new_n506), .A3(new_n662), .ZN(new_n728));
  NAND2_X1  g527(.A1(new_n728), .A2(KEYINPUT44), .ZN(new_n729));
  INV_X1    g528(.A(KEYINPUT44), .ZN(new_n730));
  OAI211_X1 g529(.A(new_n730), .B(new_n662), .C1(new_n485), .C2(new_n497), .ZN(new_n731));
  NAND2_X1  g530(.A1(new_n731), .A2(KEYINPUT100), .ZN(new_n732));
  NAND2_X1  g531(.A1(new_n504), .A2(new_n505), .ZN(new_n733));
  INV_X1    g532(.A(KEYINPUT100), .ZN(new_n734));
  NAND4_X1  g533(.A1(new_n733), .A2(new_n734), .A3(new_n730), .A4(new_n662), .ZN(new_n735));
  NAND2_X1  g534(.A1(new_n732), .A2(new_n735), .ZN(new_n736));
  NAND2_X1  g535(.A1(new_n729), .A2(new_n736), .ZN(new_n737));
  NAND2_X1  g536(.A1(new_n721), .A2(new_n600), .ZN(new_n738));
  INV_X1    g537(.A(new_n738), .ZN(new_n739));
  NAND2_X1  g538(.A1(new_n737), .A2(new_n739), .ZN(new_n740));
  OAI21_X1  g539(.A(G29gat), .B1(new_n740), .B2(new_n486), .ZN(new_n741));
  NAND2_X1  g540(.A1(new_n727), .A2(new_n741), .ZN(G1328gat));
  OAI21_X1  g541(.A(G36gat), .B1(new_n740), .B2(new_n703), .ZN(new_n743));
  NOR3_X1   g542(.A1(new_n724), .A2(G36gat), .A3(new_n703), .ZN(new_n744));
  XNOR2_X1  g543(.A(new_n744), .B(KEYINPUT46), .ZN(new_n745));
  NAND2_X1  g544(.A1(new_n743), .A2(new_n745), .ZN(G1329gat));
  NOR3_X1   g545(.A1(new_n724), .A2(G43gat), .A3(new_n714), .ZN(new_n747));
  AOI21_X1  g546(.A(new_n738), .B1(new_n729), .B2(new_n736), .ZN(new_n748));
  NAND2_X1  g547(.A1(new_n748), .A2(new_n711), .ZN(new_n749));
  AOI21_X1  g548(.A(new_n747), .B1(new_n749), .B2(G43gat), .ZN(new_n750));
  XNOR2_X1  g549(.A(new_n750), .B(KEYINPUT47), .ZN(G1330gat));
  INV_X1    g550(.A(KEYINPUT48), .ZN(new_n752));
  OAI211_X1 g551(.A(new_n525), .B(new_n270), .C1(new_n724), .C2(KEYINPUT102), .ZN(new_n753));
  INV_X1    g552(.A(new_n753), .ZN(new_n754));
  NAND2_X1  g553(.A1(new_n724), .A2(KEYINPUT102), .ZN(new_n755));
  NAND2_X1  g554(.A1(new_n754), .A2(new_n755), .ZN(new_n756));
  AOI21_X1  g555(.A(new_n525), .B1(new_n748), .B2(new_n270), .ZN(new_n757));
  INV_X1    g556(.A(KEYINPUT101), .ZN(new_n758));
  OAI21_X1  g557(.A(new_n756), .B1(new_n757), .B2(new_n758), .ZN(new_n759));
  AOI211_X1 g558(.A(KEYINPUT101), .B(new_n525), .C1(new_n748), .C2(new_n270), .ZN(new_n760));
  OAI21_X1  g559(.A(new_n752), .B1(new_n759), .B2(new_n760), .ZN(new_n761));
  OAI21_X1  g560(.A(G50gat), .B1(new_n740), .B2(new_n490), .ZN(new_n762));
  INV_X1    g561(.A(new_n755), .ZN(new_n763));
  OAI21_X1  g562(.A(KEYINPUT48), .B1(new_n763), .B2(new_n753), .ZN(new_n764));
  INV_X1    g563(.A(new_n764), .ZN(new_n765));
  INV_X1    g564(.A(KEYINPUT103), .ZN(new_n766));
  NAND3_X1  g565(.A1(new_n762), .A2(new_n765), .A3(new_n766), .ZN(new_n767));
  OAI21_X1  g566(.A(KEYINPUT103), .B1(new_n757), .B2(new_n764), .ZN(new_n768));
  NAND2_X1  g567(.A1(new_n767), .A2(new_n768), .ZN(new_n769));
  NAND2_X1  g568(.A1(new_n761), .A2(new_n769), .ZN(G1331gat));
  INV_X1    g569(.A(new_n644), .ZN(new_n771));
  NOR2_X1   g570(.A1(new_n771), .A2(new_n662), .ZN(new_n772));
  INV_X1    g571(.A(new_n600), .ZN(new_n773));
  NAND2_X1  g572(.A1(new_n772), .A2(new_n773), .ZN(new_n774));
  NOR2_X1   g573(.A1(new_n774), .A2(new_n697), .ZN(new_n775));
  AND2_X1   g574(.A1(new_n733), .A2(new_n775), .ZN(new_n776));
  XNOR2_X1  g575(.A(new_n342), .B(KEYINPUT104), .ZN(new_n777));
  NAND2_X1  g576(.A1(new_n776), .A2(new_n777), .ZN(new_n778));
  XNOR2_X1  g577(.A(new_n778), .B(G57gat), .ZN(G1332gat));
  INV_X1    g578(.A(new_n776), .ZN(new_n780));
  NOR2_X1   g579(.A1(new_n780), .A2(new_n703), .ZN(new_n781));
  NOR2_X1   g580(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n782));
  AND2_X1   g581(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n783));
  OAI21_X1  g582(.A(new_n781), .B1(new_n782), .B2(new_n783), .ZN(new_n784));
  OAI21_X1  g583(.A(new_n784), .B1(new_n781), .B2(new_n782), .ZN(G1333gat));
  INV_X1    g584(.A(KEYINPUT50), .ZN(new_n786));
  NAND3_X1  g585(.A1(new_n776), .A2(G71gat), .A3(new_n711), .ZN(new_n787));
  XNOR2_X1  g586(.A(new_n787), .B(KEYINPUT105), .ZN(new_n788));
  INV_X1    g587(.A(KEYINPUT106), .ZN(new_n789));
  INV_X1    g588(.A(G71gat), .ZN(new_n790));
  OAI21_X1  g589(.A(new_n790), .B1(new_n780), .B2(new_n714), .ZN(new_n791));
  NAND3_X1  g590(.A1(new_n788), .A2(new_n789), .A3(new_n791), .ZN(new_n792));
  INV_X1    g591(.A(new_n792), .ZN(new_n793));
  AOI21_X1  g592(.A(new_n789), .B1(new_n788), .B2(new_n791), .ZN(new_n794));
  OAI21_X1  g593(.A(new_n786), .B1(new_n793), .B2(new_n794), .ZN(new_n795));
  NAND2_X1  g594(.A1(new_n788), .A2(new_n791), .ZN(new_n796));
  NAND2_X1  g595(.A1(new_n796), .A2(KEYINPUT106), .ZN(new_n797));
  NAND3_X1  g596(.A1(new_n797), .A2(KEYINPUT50), .A3(new_n792), .ZN(new_n798));
  NAND2_X1  g597(.A1(new_n795), .A2(new_n798), .ZN(G1334gat));
  NAND2_X1  g598(.A1(new_n776), .A2(new_n270), .ZN(new_n800));
  XNOR2_X1  g599(.A(new_n800), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g600(.A1(new_n644), .A2(new_n600), .ZN(new_n802));
  NAND3_X1  g601(.A1(new_n733), .A2(new_n662), .A3(new_n802), .ZN(new_n803));
  INV_X1    g602(.A(KEYINPUT51), .ZN(new_n804));
  NAND2_X1  g603(.A1(new_n803), .A2(new_n804), .ZN(new_n805));
  NAND4_X1  g604(.A1(new_n733), .A2(KEYINPUT51), .A3(new_n662), .A4(new_n802), .ZN(new_n806));
  AOI21_X1  g605(.A(new_n697), .B1(new_n805), .B2(new_n806), .ZN(new_n807));
  NAND3_X1  g606(.A1(new_n807), .A2(new_n274), .A3(new_n342), .ZN(new_n808));
  NAND2_X1  g607(.A1(new_n802), .A2(new_n720), .ZN(new_n809));
  AOI21_X1  g608(.A(new_n809), .B1(new_n729), .B2(new_n736), .ZN(new_n810));
  AND2_X1   g609(.A1(new_n810), .A2(new_n342), .ZN(new_n811));
  OAI21_X1  g610(.A(new_n808), .B1(new_n811), .B2(new_n274), .ZN(G1336gat));
  NAND2_X1  g611(.A1(new_n810), .A2(new_n452), .ZN(new_n813));
  NOR2_X1   g612(.A1(new_n703), .A2(G92gat), .ZN(new_n814));
  AOI22_X1  g613(.A1(new_n813), .A2(G92gat), .B1(new_n807), .B2(new_n814), .ZN(new_n815));
  INV_X1    g614(.A(KEYINPUT52), .ZN(new_n816));
  XNOR2_X1  g615(.A(new_n815), .B(new_n816), .ZN(G1337gat));
  AOI21_X1  g616(.A(G99gat), .B1(new_n807), .B2(new_n442), .ZN(new_n818));
  AND2_X1   g617(.A1(new_n711), .A2(G99gat), .ZN(new_n819));
  AOI21_X1  g618(.A(new_n818), .B1(new_n810), .B2(new_n819), .ZN(G1338gat));
  XNOR2_X1  g619(.A(KEYINPUT107), .B(G106gat), .ZN(new_n821));
  AOI21_X1  g620(.A(new_n821), .B1(new_n810), .B2(new_n270), .ZN(new_n822));
  NOR2_X1   g621(.A1(new_n490), .A2(G106gat), .ZN(new_n823));
  NAND2_X1  g622(.A1(new_n807), .A2(new_n823), .ZN(new_n824));
  NAND2_X1  g623(.A1(new_n824), .A2(KEYINPUT108), .ZN(new_n825));
  NOR2_X1   g624(.A1(new_n822), .A2(new_n825), .ZN(new_n826));
  XNOR2_X1  g625(.A(KEYINPUT109), .B(KEYINPUT53), .ZN(new_n827));
  INV_X1    g626(.A(new_n827), .ZN(new_n828));
  XNOR2_X1  g627(.A(new_n826), .B(new_n828), .ZN(G1339gat));
  NAND3_X1  g628(.A1(new_n772), .A2(new_n773), .A3(new_n697), .ZN(new_n830));
  NOR3_X1   g629(.A1(new_n686), .A2(KEYINPUT10), .A3(new_n681), .ZN(new_n831));
  OAI22_X1  g630(.A1(new_n831), .A2(new_n690), .B1(new_n668), .B2(new_n245), .ZN(new_n832));
  NAND3_X1  g631(.A1(new_n683), .A2(new_n684), .A3(new_n669), .ZN(new_n833));
  NAND3_X1  g632(.A1(new_n832), .A2(KEYINPUT54), .A3(new_n833), .ZN(new_n834));
  INV_X1    g633(.A(KEYINPUT54), .ZN(new_n835));
  AOI21_X1  g634(.A(new_n666), .B1(new_n685), .B2(new_n835), .ZN(new_n836));
  NAND3_X1  g635(.A1(new_n834), .A2(new_n836), .A3(KEYINPUT55), .ZN(new_n837));
  NAND2_X1  g636(.A1(new_n837), .A2(new_n693), .ZN(new_n838));
  AOI21_X1  g637(.A(KEYINPUT55), .B1(new_n834), .B2(new_n836), .ZN(new_n839));
  NOR2_X1   g638(.A1(new_n838), .A2(new_n839), .ZN(new_n840));
  NAND2_X1  g639(.A1(new_n514), .A2(new_n515), .ZN(new_n841));
  AOI21_X1  g640(.A(new_n576), .B1(new_n597), .B2(new_n563), .ZN(new_n842));
  NOR2_X1   g641(.A1(new_n575), .A2(new_n577), .ZN(new_n843));
  OAI21_X1  g642(.A(new_n841), .B1(new_n842), .B2(new_n843), .ZN(new_n844));
  AND2_X1   g643(.A1(new_n599), .A2(new_n844), .ZN(new_n845));
  NAND3_X1  g644(.A1(new_n840), .A2(new_n662), .A3(new_n845), .ZN(new_n846));
  INV_X1    g645(.A(new_n846), .ZN(new_n847));
  AND3_X1   g646(.A1(new_n845), .A2(new_n696), .A3(new_n694), .ZN(new_n848));
  NAND2_X1  g647(.A1(new_n848), .A2(KEYINPUT110), .ZN(new_n849));
  NAND4_X1  g648(.A1(new_n694), .A2(new_n599), .A3(new_n696), .A4(new_n844), .ZN(new_n850));
  INV_X1    g649(.A(KEYINPUT110), .ZN(new_n851));
  NAND2_X1  g650(.A1(new_n850), .A2(new_n851), .ZN(new_n852));
  NAND2_X1  g651(.A1(new_n834), .A2(new_n836), .ZN(new_n853));
  INV_X1    g652(.A(KEYINPUT55), .ZN(new_n854));
  NAND2_X1  g653(.A1(new_n853), .A2(new_n854), .ZN(new_n855));
  NAND3_X1  g654(.A1(new_n855), .A2(new_n693), .A3(new_n837), .ZN(new_n856));
  OAI211_X1 g655(.A(new_n849), .B(new_n852), .C1(new_n773), .C2(new_n856), .ZN(new_n857));
  AOI21_X1  g656(.A(new_n847), .B1(new_n857), .B2(new_n663), .ZN(new_n858));
  OAI21_X1  g657(.A(new_n830), .B1(new_n858), .B2(new_n644), .ZN(new_n859));
  NAND2_X1  g658(.A1(new_n859), .A2(KEYINPUT111), .ZN(new_n860));
  INV_X1    g659(.A(KEYINPUT111), .ZN(new_n861));
  OAI211_X1 g660(.A(new_n830), .B(new_n861), .C1(new_n858), .C2(new_n644), .ZN(new_n862));
  NAND2_X1  g661(.A1(new_n860), .A2(new_n862), .ZN(new_n863));
  NOR2_X1   g662(.A1(new_n863), .A2(new_n270), .ZN(new_n864));
  NAND4_X1  g663(.A1(new_n864), .A2(new_n342), .A3(new_n703), .A4(new_n442), .ZN(new_n865));
  AND3_X1   g664(.A1(new_n594), .A2(KEYINPUT92), .A3(new_n599), .ZN(new_n866));
  AOI21_X1  g665(.A(KEYINPUT92), .B1(new_n594), .B2(new_n599), .ZN(new_n867));
  NOR2_X1   g666(.A1(new_n866), .A2(new_n867), .ZN(new_n868));
  NOR3_X1   g667(.A1(new_n865), .A2(new_n286), .A3(new_n868), .ZN(new_n869));
  INV_X1    g668(.A(new_n863), .ZN(new_n870));
  AND2_X1   g669(.A1(new_n870), .A2(new_n777), .ZN(new_n871));
  NOR3_X1   g670(.A1(new_n452), .A2(new_n270), .A3(new_n714), .ZN(new_n872));
  NAND2_X1  g671(.A1(new_n871), .A2(new_n872), .ZN(new_n873));
  INV_X1    g672(.A(new_n873), .ZN(new_n874));
  NAND2_X1  g673(.A1(new_n874), .A2(new_n600), .ZN(new_n875));
  AOI21_X1  g674(.A(new_n869), .B1(new_n875), .B2(new_n286), .ZN(G1340gat));
  NOR3_X1   g675(.A1(new_n865), .A2(new_n287), .A3(new_n697), .ZN(new_n877));
  NAND2_X1  g676(.A1(new_n874), .A2(new_n720), .ZN(new_n878));
  AOI21_X1  g677(.A(new_n877), .B1(new_n878), .B2(new_n287), .ZN(G1341gat));
  NOR3_X1   g678(.A1(new_n865), .A2(new_n279), .A3(new_n771), .ZN(new_n880));
  NAND2_X1  g679(.A1(new_n874), .A2(new_n644), .ZN(new_n881));
  OR2_X1    g680(.A1(new_n881), .A2(KEYINPUT112), .ZN(new_n882));
  AOI21_X1  g681(.A(G127gat), .B1(new_n881), .B2(KEYINPUT112), .ZN(new_n883));
  AOI21_X1  g682(.A(new_n880), .B1(new_n882), .B2(new_n883), .ZN(G1342gat));
  OAI21_X1  g683(.A(G134gat), .B1(new_n865), .B2(new_n663), .ZN(new_n885));
  XNOR2_X1  g684(.A(new_n885), .B(KEYINPUT113), .ZN(new_n886));
  NAND2_X1  g685(.A1(new_n662), .A2(new_n277), .ZN(new_n887));
  OAI21_X1  g686(.A(KEYINPUT56), .B1(new_n873), .B2(new_n887), .ZN(new_n888));
  OR3_X1    g687(.A1(new_n873), .A2(KEYINPUT56), .A3(new_n887), .ZN(new_n889));
  NAND3_X1  g688(.A1(new_n886), .A2(new_n888), .A3(new_n889), .ZN(G1343gat));
  NOR3_X1   g689(.A1(new_n711), .A2(new_n486), .A3(new_n452), .ZN(new_n891));
  INV_X1    g690(.A(new_n891), .ZN(new_n892));
  INV_X1    g691(.A(KEYINPUT117), .ZN(new_n893));
  INV_X1    g692(.A(KEYINPUT114), .ZN(new_n894));
  NAND2_X1  g693(.A1(new_n850), .A2(new_n894), .ZN(new_n895));
  NAND4_X1  g694(.A1(new_n845), .A2(KEYINPUT114), .A3(new_n694), .A4(new_n696), .ZN(new_n896));
  OAI211_X1 g695(.A(new_n895), .B(new_n896), .C1(new_n868), .C2(new_n856), .ZN(new_n897));
  NAND2_X1  g696(.A1(new_n897), .A2(KEYINPUT115), .ZN(new_n898));
  NAND2_X1  g697(.A1(new_n604), .A2(new_n840), .ZN(new_n899));
  INV_X1    g698(.A(KEYINPUT115), .ZN(new_n900));
  NAND4_X1  g699(.A1(new_n899), .A2(new_n900), .A3(new_n895), .A4(new_n896), .ZN(new_n901));
  NAND2_X1  g700(.A1(new_n898), .A2(new_n901), .ZN(new_n902));
  INV_X1    g701(.A(KEYINPUT116), .ZN(new_n903));
  NAND3_X1  g702(.A1(new_n902), .A2(new_n903), .A3(new_n663), .ZN(new_n904));
  NAND2_X1  g703(.A1(new_n904), .A2(new_n771), .ZN(new_n905));
  AOI21_X1  g704(.A(new_n662), .B1(new_n898), .B2(new_n901), .ZN(new_n906));
  NOR3_X1   g705(.A1(new_n906), .A2(new_n903), .A3(new_n847), .ZN(new_n907));
  OAI21_X1  g706(.A(new_n893), .B1(new_n905), .B2(new_n907), .ZN(new_n908));
  AOI22_X1  g707(.A1(new_n604), .A2(new_n840), .B1(new_n848), .B2(KEYINPUT114), .ZN(new_n909));
  AOI21_X1  g708(.A(new_n900), .B1(new_n909), .B2(new_n895), .ZN(new_n910));
  NOR2_X1   g709(.A1(new_n897), .A2(KEYINPUT115), .ZN(new_n911));
  OAI21_X1  g710(.A(new_n663), .B1(new_n910), .B2(new_n911), .ZN(new_n912));
  NAND3_X1  g711(.A1(new_n912), .A2(KEYINPUT116), .A3(new_n846), .ZN(new_n913));
  AOI21_X1  g712(.A(new_n644), .B1(new_n906), .B2(new_n903), .ZN(new_n914));
  NAND3_X1  g713(.A1(new_n913), .A2(KEYINPUT117), .A3(new_n914), .ZN(new_n915));
  NAND3_X1  g714(.A1(new_n908), .A2(new_n915), .A3(new_n830), .ZN(new_n916));
  INV_X1    g715(.A(KEYINPUT57), .ZN(new_n917));
  NOR2_X1   g716(.A1(new_n490), .A2(new_n917), .ZN(new_n918));
  NAND2_X1  g717(.A1(new_n916), .A2(new_n918), .ZN(new_n919));
  NAND3_X1  g718(.A1(new_n860), .A2(new_n270), .A3(new_n862), .ZN(new_n920));
  NAND2_X1  g719(.A1(new_n920), .A2(new_n917), .ZN(new_n921));
  AOI21_X1  g720(.A(new_n892), .B1(new_n919), .B2(new_n921), .ZN(new_n922));
  AOI21_X1  g721(.A(new_n209), .B1(new_n922), .B2(new_n600), .ZN(new_n923));
  NOR2_X1   g722(.A1(new_n711), .A2(new_n490), .ZN(new_n924));
  NAND4_X1  g723(.A1(new_n870), .A2(new_n703), .A3(new_n777), .A4(new_n924), .ZN(new_n925));
  NAND2_X1  g724(.A1(new_n604), .A2(new_n209), .ZN(new_n926));
  NOR2_X1   g725(.A1(new_n925), .A2(new_n926), .ZN(new_n927));
  OAI21_X1  g726(.A(KEYINPUT58), .B1(new_n923), .B2(new_n927), .ZN(new_n928));
  INV_X1    g727(.A(new_n918), .ZN(new_n929));
  INV_X1    g728(.A(new_n830), .ZN(new_n930));
  NAND2_X1  g729(.A1(new_n913), .A2(new_n914), .ZN(new_n931));
  AOI21_X1  g730(.A(new_n930), .B1(new_n931), .B2(new_n893), .ZN(new_n932));
  AOI21_X1  g731(.A(new_n929), .B1(new_n932), .B2(new_n915), .ZN(new_n933));
  INV_X1    g732(.A(new_n921), .ZN(new_n934));
  OAI211_X1 g733(.A(new_n604), .B(new_n891), .C1(new_n933), .C2(new_n934), .ZN(new_n935));
  NAND2_X1  g734(.A1(new_n935), .A2(G141gat), .ZN(new_n936));
  INV_X1    g735(.A(KEYINPUT58), .ZN(new_n937));
  OAI21_X1  g736(.A(new_n937), .B1(new_n925), .B2(new_n926), .ZN(new_n938));
  INV_X1    g737(.A(new_n938), .ZN(new_n939));
  AOI21_X1  g738(.A(KEYINPUT118), .B1(new_n936), .B2(new_n939), .ZN(new_n940));
  INV_X1    g739(.A(KEYINPUT118), .ZN(new_n941));
  AOI211_X1 g740(.A(new_n941), .B(new_n938), .C1(new_n935), .C2(G141gat), .ZN(new_n942));
  OAI21_X1  g741(.A(new_n928), .B1(new_n940), .B2(new_n942), .ZN(G1344gat));
  NOR3_X1   g742(.A1(new_n925), .A2(G148gat), .A3(new_n697), .ZN(new_n944));
  XNOR2_X1  g743(.A(new_n944), .B(KEYINPUT119), .ZN(new_n945));
  INV_X1    g744(.A(KEYINPUT59), .ZN(new_n946));
  OR3_X1    g745(.A1(new_n698), .A2(KEYINPUT121), .A3(new_n604), .ZN(new_n947));
  OAI21_X1  g746(.A(KEYINPUT121), .B1(new_n698), .B2(new_n604), .ZN(new_n948));
  NAND2_X1  g747(.A1(new_n947), .A2(new_n948), .ZN(new_n949));
  AOI21_X1  g748(.A(new_n847), .B1(new_n902), .B2(new_n663), .ZN(new_n950));
  OAI21_X1  g749(.A(new_n949), .B1(new_n950), .B2(new_n644), .ZN(new_n951));
  AOI21_X1  g750(.A(new_n490), .B1(new_n951), .B2(KEYINPUT122), .ZN(new_n952));
  INV_X1    g751(.A(KEYINPUT122), .ZN(new_n953));
  OAI211_X1 g752(.A(new_n953), .B(new_n949), .C1(new_n950), .C2(new_n644), .ZN(new_n954));
  AOI21_X1  g753(.A(KEYINPUT57), .B1(new_n952), .B2(new_n954), .ZN(new_n955));
  NOR2_X1   g754(.A1(new_n863), .A2(new_n929), .ZN(new_n956));
  OR2_X1    g755(.A1(new_n955), .A2(new_n956), .ZN(new_n957));
  XNOR2_X1  g756(.A(new_n891), .B(KEYINPUT120), .ZN(new_n958));
  NAND3_X1  g757(.A1(new_n957), .A2(new_n720), .A3(new_n958), .ZN(new_n959));
  AOI21_X1  g758(.A(new_n946), .B1(new_n959), .B2(G148gat), .ZN(new_n960));
  AOI211_X1 g759(.A(KEYINPUT59), .B(new_n206), .C1(new_n922), .C2(new_n720), .ZN(new_n961));
  OAI21_X1  g760(.A(new_n945), .B1(new_n960), .B2(new_n961), .ZN(G1345gat));
  OAI21_X1  g761(.A(new_n891), .B1(new_n933), .B2(new_n934), .ZN(new_n963));
  OAI21_X1  g762(.A(G155gat), .B1(new_n963), .B2(new_n771), .ZN(new_n964));
  NAND2_X1  g763(.A1(new_n644), .A2(new_n213), .ZN(new_n965));
  OAI211_X1 g764(.A(new_n964), .B(KEYINPUT123), .C1(new_n925), .C2(new_n965), .ZN(new_n966));
  INV_X1    g765(.A(KEYINPUT123), .ZN(new_n967));
  AOI21_X1  g766(.A(new_n213), .B1(new_n922), .B2(new_n644), .ZN(new_n968));
  NOR2_X1   g767(.A1(new_n925), .A2(new_n965), .ZN(new_n969));
  OAI21_X1  g768(.A(new_n967), .B1(new_n968), .B2(new_n969), .ZN(new_n970));
  NAND2_X1  g769(.A1(new_n966), .A2(new_n970), .ZN(G1346gat));
  OAI21_X1  g770(.A(G162gat), .B1(new_n963), .B2(new_n663), .ZN(new_n972));
  NAND2_X1  g771(.A1(new_n662), .A2(new_n214), .ZN(new_n973));
  OAI21_X1  g772(.A(new_n972), .B1(new_n925), .B2(new_n973), .ZN(G1347gat));
  NOR2_X1   g773(.A1(new_n777), .A2(new_n703), .ZN(new_n975));
  NAND3_X1  g774(.A1(new_n864), .A2(new_n442), .A3(new_n975), .ZN(new_n976));
  OAI21_X1  g775(.A(G169gat), .B1(new_n976), .B2(new_n868), .ZN(new_n977));
  INV_X1    g776(.A(new_n493), .ZN(new_n978));
  NOR4_X1   g777(.A1(new_n863), .A2(new_n342), .A3(new_n703), .A4(new_n978), .ZN(new_n979));
  NAND4_X1  g778(.A1(new_n979), .A2(new_n374), .A3(new_n375), .A4(new_n600), .ZN(new_n980));
  NAND2_X1  g779(.A1(new_n977), .A2(new_n980), .ZN(G1348gat));
  OAI21_X1  g780(.A(G176gat), .B1(new_n976), .B2(new_n697), .ZN(new_n982));
  NAND3_X1  g781(.A1(new_n979), .A2(new_n345), .A3(new_n720), .ZN(new_n983));
  NAND2_X1  g782(.A1(new_n982), .A2(new_n983), .ZN(new_n984));
  XOR2_X1   g783(.A(new_n984), .B(KEYINPUT124), .Z(G1349gat));
  OAI21_X1  g784(.A(G183gat), .B1(new_n976), .B2(new_n771), .ZN(new_n986));
  NAND3_X1  g785(.A1(new_n979), .A2(new_n360), .A3(new_n644), .ZN(new_n987));
  NAND2_X1  g786(.A1(new_n986), .A2(new_n987), .ZN(new_n988));
  XNOR2_X1  g787(.A(new_n988), .B(KEYINPUT60), .ZN(G1350gat));
  OAI21_X1  g788(.A(G190gat), .B1(new_n976), .B2(new_n663), .ZN(new_n990));
  XNOR2_X1  g789(.A(new_n990), .B(KEYINPUT61), .ZN(new_n991));
  NAND3_X1  g790(.A1(new_n979), .A2(new_n361), .A3(new_n662), .ZN(new_n992));
  NAND2_X1  g791(.A1(new_n991), .A2(new_n992), .ZN(G1351gat));
  NAND4_X1  g792(.A1(new_n870), .A2(new_n486), .A3(new_n452), .A4(new_n924), .ZN(new_n994));
  INV_X1    g793(.A(new_n994), .ZN(new_n995));
  AOI21_X1  g794(.A(G197gat), .B1(new_n995), .B2(new_n600), .ZN(new_n996));
  NOR3_X1   g795(.A1(new_n777), .A2(new_n703), .A3(new_n711), .ZN(new_n997));
  NAND2_X1  g796(.A1(new_n957), .A2(new_n997), .ZN(new_n998));
  INV_X1    g797(.A(new_n998), .ZN(new_n999));
  AND2_X1   g798(.A1(new_n604), .A2(G197gat), .ZN(new_n1000));
  AOI21_X1  g799(.A(new_n996), .B1(new_n999), .B2(new_n1000), .ZN(G1352gat));
  XNOR2_X1  g800(.A(KEYINPUT125), .B(G204gat), .ZN(new_n1002));
  OAI21_X1  g801(.A(new_n1002), .B1(new_n998), .B2(new_n697), .ZN(new_n1003));
  NOR3_X1   g802(.A1(new_n994), .A2(new_n697), .A3(new_n1002), .ZN(new_n1004));
  XNOR2_X1  g803(.A(new_n1004), .B(KEYINPUT62), .ZN(new_n1005));
  NAND2_X1  g804(.A1(new_n1003), .A2(new_n1005), .ZN(G1353gat));
  OAI211_X1 g805(.A(new_n644), .B(new_n997), .C1(new_n955), .C2(new_n956), .ZN(new_n1007));
  NAND2_X1  g806(.A1(new_n1007), .A2(G211gat), .ZN(new_n1008));
  INV_X1    g807(.A(KEYINPUT63), .ZN(new_n1009));
  NAND2_X1  g808(.A1(new_n1008), .A2(new_n1009), .ZN(new_n1010));
  NAND3_X1  g809(.A1(new_n1007), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n1011));
  NAND3_X1  g810(.A1(new_n1010), .A2(KEYINPUT126), .A3(new_n1011), .ZN(new_n1012));
  AND3_X1   g811(.A1(new_n995), .A2(new_n230), .A3(new_n644), .ZN(new_n1013));
  AOI21_X1  g812(.A(KEYINPUT63), .B1(new_n1007), .B2(G211gat), .ZN(new_n1014));
  INV_X1    g813(.A(KEYINPUT126), .ZN(new_n1015));
  AOI21_X1  g814(.A(new_n1013), .B1(new_n1014), .B2(new_n1015), .ZN(new_n1016));
  NAND2_X1  g815(.A1(new_n1012), .A2(new_n1016), .ZN(G1354gat));
  NOR3_X1   g816(.A1(new_n998), .A2(new_n231), .A3(new_n663), .ZN(new_n1018));
  OAI21_X1  g817(.A(new_n231), .B1(new_n994), .B2(new_n663), .ZN(new_n1019));
  XNOR2_X1  g818(.A(new_n1019), .B(KEYINPUT127), .ZN(new_n1020));
  NOR2_X1   g819(.A1(new_n1018), .A2(new_n1020), .ZN(G1355gat));
endmodule


