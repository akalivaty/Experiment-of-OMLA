//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 0 1 1 0 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 1 1 0 0 0 0 0 1 1 0 1 0 0 0 0 0 0 1 1 0 1 1 1 0 0 0 1 0 1 1 1 1 1 1 1 1 1 1 1 1 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:30:03 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n443, new_n447, new_n448, new_n450, new_n453, new_n454, new_n455,
    new_n456, new_n457, new_n460, new_n461, new_n462, new_n463, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n531, new_n532, new_n533,
    new_n534, new_n535, new_n536, new_n537, new_n540, new_n541, new_n542,
    new_n543, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n554, new_n555, new_n557, new_n558, new_n559, new_n560, new_n561,
    new_n562, new_n564, new_n565, new_n566, new_n568, new_n569, new_n570,
    new_n571, new_n572, new_n573, new_n574, new_n575, new_n576, new_n577,
    new_n578, new_n580, new_n581, new_n582, new_n583, new_n584, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n601, new_n602,
    new_n603, new_n606, new_n608, new_n609, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n822, new_n823, new_n824,
    new_n825, new_n826, new_n827, new_n828, new_n829, new_n830, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n899, new_n900, new_n901, new_n902, new_n903, new_n904, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1138, new_n1139;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  XOR2_X1   g011(.A(KEYINPUT64), .B(G96), .Z(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(new_n443));
  XOR2_X1   g018(.A(new_n443), .B(KEYINPUT65), .Z(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  XNOR2_X1  g021(.A(KEYINPUT66), .B(KEYINPUT1), .ZN(new_n447));
  NAND2_X1  g022(.A1(G7), .A2(G661), .ZN(new_n448));
  XNOR2_X1  g023(.A(new_n447), .B(new_n448), .ZN(G223));
  INV_X1    g024(.A(new_n448), .ZN(new_n450));
  NAND2_X1  g025(.A1(new_n450), .A2(G567), .ZN(G234));
  NAND2_X1  g026(.A1(new_n450), .A2(G2106), .ZN(G217));
  NOR4_X1   g027(.A1(G221), .A2(G220), .A3(G218), .A4(G219), .ZN(new_n453));
  XNOR2_X1  g028(.A(new_n453), .B(KEYINPUT2), .ZN(new_n454));
  NAND4_X1  g029(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n455));
  XOR2_X1   g030(.A(new_n455), .B(KEYINPUT67), .Z(new_n456));
  NAND2_X1  g031(.A1(new_n454), .A2(new_n456), .ZN(new_n457));
  INV_X1    g032(.A(new_n457), .ZN(G325));
  XNOR2_X1  g033(.A(new_n457), .B(KEYINPUT68), .ZN(G261));
  INV_X1    g034(.A(G2106), .ZN(new_n460));
  INV_X1    g035(.A(G567), .ZN(new_n461));
  OAI22_X1  g036(.A1(new_n454), .A2(new_n460), .B1(new_n461), .B2(new_n456), .ZN(new_n462));
  XNOR2_X1  g037(.A(new_n462), .B(KEYINPUT69), .ZN(new_n463));
  XOR2_X1   g038(.A(new_n463), .B(KEYINPUT70), .Z(G319));
  AND2_X1   g039(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n465));
  NOR2_X1   g040(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n466));
  NOR2_X1   g041(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  NOR2_X1   g042(.A1(new_n467), .A2(G2105), .ZN(new_n468));
  INV_X1    g043(.A(G2104), .ZN(new_n469));
  NOR2_X1   g044(.A1(new_n469), .A2(G2105), .ZN(new_n470));
  AOI22_X1  g045(.A1(new_n468), .A2(G137), .B1(G101), .B2(new_n470), .ZN(new_n471));
  INV_X1    g046(.A(G113), .ZN(new_n472));
  OAI21_X1  g047(.A(KEYINPUT71), .B1(new_n472), .B2(new_n469), .ZN(new_n473));
  INV_X1    g048(.A(KEYINPUT71), .ZN(new_n474));
  NAND3_X1  g049(.A1(new_n474), .A2(G113), .A3(G2104), .ZN(new_n475));
  INV_X1    g050(.A(G125), .ZN(new_n476));
  OAI211_X1 g051(.A(new_n473), .B(new_n475), .C1(new_n467), .C2(new_n476), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n477), .A2(G2105), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n471), .A2(new_n478), .ZN(new_n479));
  INV_X1    g054(.A(new_n479), .ZN(G160));
  NAND2_X1  g055(.A1(new_n468), .A2(G136), .ZN(new_n481));
  INV_X1    g056(.A(G2105), .ZN(new_n482));
  INV_X1    g057(.A(KEYINPUT3), .ZN(new_n483));
  NAND2_X1  g058(.A1(new_n483), .A2(new_n469), .ZN(new_n484));
  NAND2_X1  g059(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n485));
  AOI21_X1  g060(.A(new_n482), .B1(new_n484), .B2(new_n485), .ZN(new_n486));
  NAND2_X1  g061(.A1(new_n486), .A2(G124), .ZN(new_n487));
  OR2_X1    g062(.A1(G100), .A2(G2105), .ZN(new_n488));
  OAI211_X1 g063(.A(new_n488), .B(G2104), .C1(G112), .C2(new_n482), .ZN(new_n489));
  NAND3_X1  g064(.A1(new_n481), .A2(new_n487), .A3(new_n489), .ZN(new_n490));
  INV_X1    g065(.A(new_n490), .ZN(G162));
  INV_X1    g066(.A(G138), .ZN(new_n492));
  NOR2_X1   g067(.A1(new_n492), .A2(G2105), .ZN(new_n493));
  OAI21_X1  g068(.A(new_n493), .B1(new_n465), .B2(new_n466), .ZN(new_n494));
  INV_X1    g069(.A(KEYINPUT72), .ZN(new_n495));
  NAND2_X1  g070(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  XNOR2_X1  g071(.A(KEYINPUT3), .B(G2104), .ZN(new_n497));
  NAND3_X1  g072(.A1(new_n497), .A2(KEYINPUT72), .A3(new_n493), .ZN(new_n498));
  NAND3_X1  g073(.A1(new_n496), .A2(KEYINPUT4), .A3(new_n498), .ZN(new_n499));
  INV_X1    g074(.A(KEYINPUT4), .ZN(new_n500));
  NAND3_X1  g075(.A1(new_n494), .A2(new_n495), .A3(new_n500), .ZN(new_n501));
  INV_X1    g076(.A(G114), .ZN(new_n502));
  NAND2_X1  g077(.A1(new_n502), .A2(G2105), .ZN(new_n503));
  OAI21_X1  g078(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n504));
  INV_X1    g079(.A(new_n504), .ZN(new_n505));
  AOI22_X1  g080(.A1(new_n486), .A2(G126), .B1(new_n503), .B2(new_n505), .ZN(new_n506));
  NAND3_X1  g081(.A1(new_n499), .A2(new_n501), .A3(new_n506), .ZN(new_n507));
  INV_X1    g082(.A(new_n507), .ZN(G164));
  INV_X1    g083(.A(KEYINPUT73), .ZN(new_n509));
  INV_X1    g084(.A(KEYINPUT6), .ZN(new_n510));
  OAI21_X1  g085(.A(new_n509), .B1(new_n510), .B2(G651), .ZN(new_n511));
  INV_X1    g086(.A(G651), .ZN(new_n512));
  NAND3_X1  g087(.A1(new_n512), .A2(KEYINPUT73), .A3(KEYINPUT6), .ZN(new_n513));
  NAND2_X1  g088(.A1(new_n511), .A2(new_n513), .ZN(new_n514));
  NAND2_X1  g089(.A1(new_n510), .A2(G651), .ZN(new_n515));
  NAND2_X1  g090(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  INV_X1    g091(.A(G543), .ZN(new_n517));
  NOR2_X1   g092(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  NAND2_X1  g093(.A1(new_n518), .A2(G50), .ZN(new_n519));
  INV_X1    g094(.A(KEYINPUT5), .ZN(new_n520));
  NAND2_X1  g095(.A1(new_n520), .A2(new_n517), .ZN(new_n521));
  NAND2_X1  g096(.A1(KEYINPUT5), .A2(G543), .ZN(new_n522));
  NAND2_X1  g097(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  INV_X1    g098(.A(new_n523), .ZN(new_n524));
  NOR2_X1   g099(.A1(new_n516), .A2(new_n524), .ZN(new_n525));
  NAND2_X1  g100(.A1(new_n525), .A2(G88), .ZN(new_n526));
  AOI22_X1  g101(.A1(new_n523), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n527));
  OR2_X1    g102(.A1(new_n527), .A2(new_n512), .ZN(new_n528));
  NAND3_X1  g103(.A1(new_n519), .A2(new_n526), .A3(new_n528), .ZN(G303));
  INV_X1    g104(.A(G303), .ZN(G166));
  NAND2_X1  g105(.A1(new_n525), .A2(G89), .ZN(new_n531));
  NAND2_X1  g106(.A1(new_n518), .A2(G51), .ZN(new_n532));
  NAND3_X1  g107(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n533));
  OR2_X1    g108(.A1(new_n533), .A2(KEYINPUT7), .ZN(new_n534));
  NAND2_X1  g109(.A1(new_n533), .A2(KEYINPUT7), .ZN(new_n535));
  AND2_X1   g110(.A1(G63), .A2(G651), .ZN(new_n536));
  AOI22_X1  g111(.A1(new_n534), .A2(new_n535), .B1(new_n523), .B2(new_n536), .ZN(new_n537));
  NAND3_X1  g112(.A1(new_n531), .A2(new_n532), .A3(new_n537), .ZN(G286));
  INV_X1    g113(.A(G286), .ZN(G168));
  NAND2_X1  g114(.A1(new_n525), .A2(G90), .ZN(new_n540));
  NAND2_X1  g115(.A1(new_n518), .A2(G52), .ZN(new_n541));
  AOI22_X1  g116(.A1(new_n523), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n542));
  OR2_X1    g117(.A1(new_n542), .A2(new_n512), .ZN(new_n543));
  NAND3_X1  g118(.A1(new_n540), .A2(new_n541), .A3(new_n543), .ZN(G301));
  INV_X1    g119(.A(G301), .ZN(G171));
  NAND2_X1  g120(.A1(new_n525), .A2(G81), .ZN(new_n546));
  NAND2_X1  g121(.A1(new_n518), .A2(G43), .ZN(new_n547));
  AOI22_X1  g122(.A1(new_n523), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n548));
  OR2_X1    g123(.A1(new_n548), .A2(new_n512), .ZN(new_n549));
  NAND3_X1  g124(.A1(new_n546), .A2(new_n547), .A3(new_n549), .ZN(new_n550));
  INV_X1    g125(.A(new_n550), .ZN(new_n551));
  NAND2_X1  g126(.A1(new_n551), .A2(G860), .ZN(G153));
  NAND4_X1  g127(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g128(.A1(G1), .A2(G3), .ZN(new_n554));
  XNOR2_X1  g129(.A(new_n554), .B(KEYINPUT8), .ZN(new_n555));
  NAND4_X1  g130(.A1(G319), .A2(G483), .A3(G661), .A4(new_n555), .ZN(G188));
  NAND4_X1  g131(.A1(new_n514), .A2(G53), .A3(G543), .A4(new_n515), .ZN(new_n557));
  XNOR2_X1  g132(.A(new_n557), .B(KEYINPUT9), .ZN(new_n558));
  NAND2_X1  g133(.A1(G78), .A2(G543), .ZN(new_n559));
  INV_X1    g134(.A(G65), .ZN(new_n560));
  OAI21_X1  g135(.A(new_n559), .B1(new_n524), .B2(new_n560), .ZN(new_n561));
  AOI22_X1  g136(.A1(new_n525), .A2(G91), .B1(new_n561), .B2(G651), .ZN(new_n562));
  NAND2_X1  g137(.A1(new_n558), .A2(new_n562), .ZN(G299));
  NAND2_X1  g138(.A1(new_n518), .A2(G49), .ZN(new_n564));
  NAND2_X1  g139(.A1(new_n525), .A2(G87), .ZN(new_n565));
  OAI21_X1  g140(.A(G651), .B1(new_n523), .B2(G74), .ZN(new_n566));
  NAND3_X1  g141(.A1(new_n564), .A2(new_n565), .A3(new_n566), .ZN(G288));
  INV_X1    g142(.A(G61), .ZN(new_n568));
  AOI21_X1  g143(.A(new_n568), .B1(new_n521), .B2(new_n522), .ZN(new_n569));
  INV_X1    g144(.A(KEYINPUT74), .ZN(new_n570));
  NAND2_X1  g145(.A1(new_n569), .A2(new_n570), .ZN(new_n571));
  INV_X1    g146(.A(new_n571), .ZN(new_n572));
  NAND2_X1  g147(.A1(G73), .A2(G543), .ZN(new_n573));
  OAI21_X1  g148(.A(new_n573), .B1(new_n569), .B2(new_n570), .ZN(new_n574));
  OAI21_X1  g149(.A(G651), .B1(new_n572), .B2(new_n574), .ZN(new_n575));
  NAND4_X1  g150(.A1(new_n514), .A2(G86), .A3(new_n515), .A4(new_n523), .ZN(new_n576));
  NAND4_X1  g151(.A1(new_n514), .A2(G48), .A3(G543), .A4(new_n515), .ZN(new_n577));
  AND2_X1   g152(.A1(new_n576), .A2(new_n577), .ZN(new_n578));
  NAND2_X1  g153(.A1(new_n575), .A2(new_n578), .ZN(G305));
  AOI22_X1  g154(.A1(new_n523), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n580));
  NOR2_X1   g155(.A1(new_n580), .A2(new_n512), .ZN(new_n581));
  INV_X1    g156(.A(KEYINPUT75), .ZN(new_n582));
  XNOR2_X1  g157(.A(new_n581), .B(new_n582), .ZN(new_n583));
  AOI22_X1  g158(.A1(G47), .A2(new_n518), .B1(new_n525), .B2(G85), .ZN(new_n584));
  NAND2_X1  g159(.A1(new_n583), .A2(new_n584), .ZN(G290));
  NAND2_X1  g160(.A1(G301), .A2(G868), .ZN(new_n586));
  NAND2_X1  g161(.A1(new_n525), .A2(G92), .ZN(new_n587));
  XNOR2_X1  g162(.A(new_n587), .B(KEYINPUT10), .ZN(new_n588));
  NAND2_X1  g163(.A1(new_n518), .A2(G54), .ZN(new_n589));
  XNOR2_X1  g164(.A(KEYINPUT77), .B(G66), .ZN(new_n590));
  NAND2_X1  g165(.A1(new_n523), .A2(new_n590), .ZN(new_n591));
  NAND2_X1  g166(.A1(G79), .A2(G543), .ZN(new_n592));
  XNOR2_X1  g167(.A(new_n592), .B(KEYINPUT76), .ZN(new_n593));
  AOI21_X1  g168(.A(KEYINPUT78), .B1(new_n591), .B2(new_n593), .ZN(new_n594));
  NAND3_X1  g169(.A1(new_n591), .A2(new_n593), .A3(KEYINPUT78), .ZN(new_n595));
  NAND2_X1  g170(.A1(new_n595), .A2(G651), .ZN(new_n596));
  OAI21_X1  g171(.A(new_n589), .B1(new_n594), .B2(new_n596), .ZN(new_n597));
  NOR2_X1   g172(.A1(new_n588), .A2(new_n597), .ZN(new_n598));
  OAI21_X1  g173(.A(new_n586), .B1(new_n598), .B2(G868), .ZN(G284));
  XNOR2_X1  g174(.A(G284), .B(KEYINPUT79), .ZN(G321));
  INV_X1    g175(.A(G868), .ZN(new_n601));
  NOR2_X1   g176(.A1(G286), .A2(new_n601), .ZN(new_n602));
  XNOR2_X1  g177(.A(G299), .B(KEYINPUT80), .ZN(new_n603));
  AOI21_X1  g178(.A(new_n602), .B1(new_n603), .B2(new_n601), .ZN(G297));
  AOI21_X1  g179(.A(new_n602), .B1(new_n603), .B2(new_n601), .ZN(G280));
  INV_X1    g180(.A(G559), .ZN(new_n606));
  OAI21_X1  g181(.A(new_n598), .B1(new_n606), .B2(G860), .ZN(G148));
  NAND2_X1  g182(.A1(new_n598), .A2(new_n606), .ZN(new_n608));
  NAND2_X1  g183(.A1(new_n608), .A2(G868), .ZN(new_n609));
  OAI21_X1  g184(.A(new_n609), .B1(G868), .B2(new_n551), .ZN(G323));
  XNOR2_X1  g185(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g186(.A1(new_n468), .A2(G135), .ZN(new_n612));
  XNOR2_X1  g187(.A(new_n612), .B(KEYINPUT82), .ZN(new_n613));
  NAND2_X1  g188(.A1(new_n486), .A2(G123), .ZN(new_n614));
  NOR2_X1   g189(.A1(new_n482), .A2(G111), .ZN(new_n615));
  OAI21_X1  g190(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n616));
  OAI211_X1 g191(.A(new_n613), .B(new_n614), .C1(new_n615), .C2(new_n616), .ZN(new_n617));
  OR2_X1    g192(.A1(new_n617), .A2(G2096), .ZN(new_n618));
  NAND2_X1  g193(.A1(new_n497), .A2(new_n470), .ZN(new_n619));
  XOR2_X1   g194(.A(KEYINPUT81), .B(KEYINPUT12), .Z(new_n620));
  XNOR2_X1  g195(.A(new_n619), .B(new_n620), .ZN(new_n621));
  XNOR2_X1  g196(.A(new_n621), .B(KEYINPUT13), .ZN(new_n622));
  OR2_X1    g197(.A1(new_n622), .A2(G2100), .ZN(new_n623));
  NAND2_X1  g198(.A1(new_n622), .A2(G2100), .ZN(new_n624));
  NAND2_X1  g199(.A1(new_n617), .A2(G2096), .ZN(new_n625));
  NAND4_X1  g200(.A1(new_n618), .A2(new_n623), .A3(new_n624), .A4(new_n625), .ZN(G156));
  XNOR2_X1  g201(.A(KEYINPUT15), .B(G2435), .ZN(new_n627));
  XNOR2_X1  g202(.A(new_n627), .B(G2438), .ZN(new_n628));
  XNOR2_X1  g203(.A(G2427), .B(G2430), .ZN(new_n629));
  NAND2_X1  g204(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  AND3_X1   g205(.A1(new_n630), .A2(KEYINPUT83), .A3(KEYINPUT14), .ZN(new_n631));
  AOI21_X1  g206(.A(KEYINPUT83), .B1(new_n630), .B2(KEYINPUT14), .ZN(new_n632));
  OAI22_X1  g207(.A1(new_n631), .A2(new_n632), .B1(new_n628), .B2(new_n629), .ZN(new_n633));
  XOR2_X1   g208(.A(G2451), .B(G2454), .Z(new_n634));
  XNOR2_X1  g209(.A(new_n634), .B(KEYINPUT16), .ZN(new_n635));
  XNOR2_X1  g210(.A(new_n635), .B(KEYINPUT84), .ZN(new_n636));
  XNOR2_X1  g211(.A(new_n633), .B(new_n636), .ZN(new_n637));
  XNOR2_X1  g212(.A(G2443), .B(G2446), .ZN(new_n638));
  XNOR2_X1  g213(.A(new_n638), .B(KEYINPUT85), .ZN(new_n639));
  XNOR2_X1  g214(.A(new_n637), .B(new_n639), .ZN(new_n640));
  XNOR2_X1  g215(.A(G1341), .B(G1348), .ZN(new_n641));
  INV_X1    g216(.A(new_n641), .ZN(new_n642));
  OAI21_X1  g217(.A(G14), .B1(new_n640), .B2(new_n642), .ZN(new_n643));
  AOI21_X1  g218(.A(new_n643), .B1(new_n642), .B2(new_n640), .ZN(G401));
  XNOR2_X1  g219(.A(G2084), .B(G2090), .ZN(new_n645));
  XNOR2_X1  g220(.A(new_n645), .B(KEYINPUT86), .ZN(new_n646));
  INV_X1    g221(.A(new_n646), .ZN(new_n647));
  XNOR2_X1  g222(.A(G2067), .B(G2678), .ZN(new_n648));
  XNOR2_X1  g223(.A(G2072), .B(G2078), .ZN(new_n649));
  NAND3_X1  g224(.A1(new_n647), .A2(new_n648), .A3(new_n649), .ZN(new_n650));
  XOR2_X1   g225(.A(new_n650), .B(KEYINPUT18), .Z(new_n651));
  OAI21_X1  g226(.A(new_n646), .B1(new_n648), .B2(new_n649), .ZN(new_n652));
  OR2_X1    g227(.A1(new_n652), .A2(KEYINPUT87), .ZN(new_n653));
  NAND2_X1  g228(.A1(new_n652), .A2(KEYINPUT87), .ZN(new_n654));
  INV_X1    g229(.A(new_n648), .ZN(new_n655));
  XOR2_X1   g230(.A(new_n649), .B(KEYINPUT17), .Z(new_n656));
  OAI211_X1 g231(.A(new_n653), .B(new_n654), .C1(new_n655), .C2(new_n656), .ZN(new_n657));
  NAND3_X1  g232(.A1(new_n647), .A2(new_n656), .A3(new_n655), .ZN(new_n658));
  NAND3_X1  g233(.A1(new_n651), .A2(new_n657), .A3(new_n658), .ZN(new_n659));
  XOR2_X1   g234(.A(G2096), .B(G2100), .Z(new_n660));
  XNOR2_X1  g235(.A(new_n659), .B(new_n660), .ZN(G227));
  XOR2_X1   g236(.A(G1971), .B(G1976), .Z(new_n662));
  XNOR2_X1  g237(.A(KEYINPUT88), .B(KEYINPUT19), .ZN(new_n663));
  XNOR2_X1  g238(.A(new_n662), .B(new_n663), .ZN(new_n664));
  XNOR2_X1  g239(.A(G1956), .B(G2474), .ZN(new_n665));
  XNOR2_X1  g240(.A(G1961), .B(G1966), .ZN(new_n666));
  NOR2_X1   g241(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  INV_X1    g242(.A(new_n667), .ZN(new_n668));
  NOR2_X1   g243(.A1(new_n664), .A2(new_n668), .ZN(new_n669));
  XOR2_X1   g244(.A(new_n669), .B(KEYINPUT20), .Z(new_n670));
  NAND2_X1  g245(.A1(new_n665), .A2(new_n666), .ZN(new_n671));
  NAND3_X1  g246(.A1(new_n664), .A2(new_n668), .A3(new_n671), .ZN(new_n672));
  OAI211_X1 g247(.A(new_n670), .B(new_n672), .C1(new_n664), .C2(new_n671), .ZN(new_n673));
  XNOR2_X1  g248(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n674));
  XNOR2_X1  g249(.A(new_n673), .B(new_n674), .ZN(new_n675));
  XNOR2_X1  g250(.A(G1991), .B(G1996), .ZN(new_n676));
  XNOR2_X1  g251(.A(new_n675), .B(new_n676), .ZN(new_n677));
  XNOR2_X1  g252(.A(G1981), .B(G1986), .ZN(new_n678));
  XNOR2_X1  g253(.A(new_n677), .B(new_n678), .ZN(G229));
  XOR2_X1   g254(.A(KEYINPUT31), .B(G11), .Z(new_n680));
  XNOR2_X1  g255(.A(new_n680), .B(KEYINPUT100), .ZN(new_n681));
  INV_X1    g256(.A(KEYINPUT30), .ZN(new_n682));
  AND2_X1   g257(.A1(new_n682), .A2(G28), .ZN(new_n683));
  INV_X1    g258(.A(G29), .ZN(new_n684));
  OAI21_X1  g259(.A(new_n684), .B1(new_n682), .B2(G28), .ZN(new_n685));
  OAI221_X1 g260(.A(new_n681), .B1(new_n683), .B2(new_n685), .C1(new_n617), .C2(new_n684), .ZN(new_n686));
  XNOR2_X1  g261(.A(new_n686), .B(KEYINPUT101), .ZN(new_n687));
  INV_X1    g262(.A(G16), .ZN(new_n688));
  NOR2_X1   g263(.A1(G171), .A2(new_n688), .ZN(new_n689));
  AOI21_X1  g264(.A(new_n689), .B1(G5), .B2(new_n688), .ZN(new_n690));
  INV_X1    g265(.A(new_n690), .ZN(new_n691));
  OAI21_X1  g266(.A(new_n687), .B1(G1961), .B2(new_n691), .ZN(new_n692));
  NAND2_X1  g267(.A1(new_n684), .A2(G32), .ZN(new_n693));
  NAND2_X1  g268(.A1(new_n470), .A2(G105), .ZN(new_n694));
  XOR2_X1   g269(.A(new_n694), .B(KEYINPUT95), .Z(new_n695));
  NAND2_X1  g270(.A1(new_n468), .A2(G141), .ZN(new_n696));
  NAND2_X1  g271(.A1(new_n695), .A2(new_n696), .ZN(new_n697));
  XOR2_X1   g272(.A(KEYINPUT96), .B(KEYINPUT26), .Z(new_n698));
  NAND3_X1  g273(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n699));
  XNOR2_X1  g274(.A(new_n698), .B(new_n699), .ZN(new_n700));
  NAND2_X1  g275(.A1(new_n486), .A2(G129), .ZN(new_n701));
  NAND2_X1  g276(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  NOR2_X1   g277(.A1(new_n697), .A2(new_n702), .ZN(new_n703));
  OAI21_X1  g278(.A(new_n693), .B1(new_n703), .B2(new_n684), .ZN(new_n704));
  XOR2_X1   g279(.A(KEYINPUT27), .B(G1996), .Z(new_n705));
  XNOR2_X1  g280(.A(new_n705), .B(KEYINPUT97), .ZN(new_n706));
  XNOR2_X1  g281(.A(new_n704), .B(new_n706), .ZN(new_n707));
  NOR2_X1   g282(.A1(G27), .A2(G29), .ZN(new_n708));
  AOI21_X1  g283(.A(new_n708), .B1(G164), .B2(G29), .ZN(new_n709));
  XOR2_X1   g284(.A(new_n709), .B(G2078), .Z(new_n710));
  XNOR2_X1  g285(.A(KEYINPUT94), .B(KEYINPUT24), .ZN(new_n711));
  XNOR2_X1  g286(.A(new_n711), .B(G34), .ZN(new_n712));
  NAND2_X1  g287(.A1(new_n712), .A2(new_n684), .ZN(new_n713));
  OAI21_X1  g288(.A(new_n713), .B1(new_n479), .B2(new_n684), .ZN(new_n714));
  XNOR2_X1  g289(.A(new_n714), .B(G2084), .ZN(new_n715));
  NAND3_X1  g290(.A1(new_n707), .A2(new_n710), .A3(new_n715), .ZN(new_n716));
  AND2_X1   g291(.A1(new_n497), .A2(G127), .ZN(new_n717));
  AND2_X1   g292(.A1(G115), .A2(G2104), .ZN(new_n718));
  OAI21_X1  g293(.A(G2105), .B1(new_n717), .B2(new_n718), .ZN(new_n719));
  INV_X1    g294(.A(KEYINPUT93), .ZN(new_n720));
  OR2_X1    g295(.A1(new_n719), .A2(new_n720), .ZN(new_n721));
  NAND2_X1  g296(.A1(new_n719), .A2(new_n720), .ZN(new_n722));
  INV_X1    g297(.A(KEYINPUT25), .ZN(new_n723));
  NAND2_X1  g298(.A1(G103), .A2(G2104), .ZN(new_n724));
  OAI21_X1  g299(.A(new_n723), .B1(new_n724), .B2(G2105), .ZN(new_n725));
  NAND4_X1  g300(.A1(new_n482), .A2(KEYINPUT25), .A3(G103), .A4(G2104), .ZN(new_n726));
  AOI22_X1  g301(.A1(new_n468), .A2(G139), .B1(new_n725), .B2(new_n726), .ZN(new_n727));
  NAND3_X1  g302(.A1(new_n721), .A2(new_n722), .A3(new_n727), .ZN(new_n728));
  MUX2_X1   g303(.A(G33), .B(new_n728), .S(G29), .Z(new_n729));
  XNOR2_X1  g304(.A(new_n729), .B(G2072), .ZN(new_n730));
  NOR3_X1   g305(.A1(new_n692), .A2(new_n716), .A3(new_n730), .ZN(new_n731));
  NAND2_X1  g306(.A1(G168), .A2(G16), .ZN(new_n732));
  NOR2_X1   g307(.A1(G16), .A2(G21), .ZN(new_n733));
  OAI21_X1  g308(.A(new_n732), .B1(KEYINPUT98), .B2(new_n733), .ZN(new_n734));
  OAI21_X1  g309(.A(new_n734), .B1(KEYINPUT98), .B2(new_n732), .ZN(new_n735));
  XNOR2_X1  g310(.A(KEYINPUT99), .B(G1966), .ZN(new_n736));
  XOR2_X1   g311(.A(new_n735), .B(new_n736), .Z(new_n737));
  AOI21_X1  g312(.A(KEYINPUT102), .B1(new_n691), .B2(G1961), .ZN(new_n738));
  AND3_X1   g313(.A1(new_n691), .A2(KEYINPUT102), .A3(G1961), .ZN(new_n739));
  OAI211_X1 g314(.A(new_n731), .B(new_n737), .C1(new_n738), .C2(new_n739), .ZN(new_n740));
  OR2_X1    g315(.A1(new_n740), .A2(KEYINPUT103), .ZN(new_n741));
  NAND2_X1  g316(.A1(new_n688), .A2(G22), .ZN(new_n742));
  OAI21_X1  g317(.A(new_n742), .B1(G166), .B2(new_n688), .ZN(new_n743));
  INV_X1    g318(.A(G1971), .ZN(new_n744));
  XNOR2_X1  g319(.A(new_n743), .B(new_n744), .ZN(new_n745));
  NAND2_X1  g320(.A1(new_n688), .A2(G23), .ZN(new_n746));
  INV_X1    g321(.A(G288), .ZN(new_n747));
  OAI21_X1  g322(.A(new_n746), .B1(new_n747), .B2(new_n688), .ZN(new_n748));
  XOR2_X1   g323(.A(KEYINPUT33), .B(G1976), .Z(new_n749));
  XNOR2_X1  g324(.A(new_n749), .B(KEYINPUT91), .ZN(new_n750));
  XNOR2_X1  g325(.A(new_n748), .B(new_n750), .ZN(new_n751));
  MUX2_X1   g326(.A(G6), .B(G305), .S(G16), .Z(new_n752));
  XOR2_X1   g327(.A(KEYINPUT32), .B(G1981), .Z(new_n753));
  XNOR2_X1  g328(.A(new_n752), .B(new_n753), .ZN(new_n754));
  NAND3_X1  g329(.A1(new_n745), .A2(new_n751), .A3(new_n754), .ZN(new_n755));
  OR2_X1    g330(.A1(new_n755), .A2(KEYINPUT34), .ZN(new_n756));
  NAND2_X1  g331(.A1(new_n755), .A2(KEYINPUT34), .ZN(new_n757));
  MUX2_X1   g332(.A(G24), .B(G290), .S(G16), .Z(new_n758));
  NAND2_X1  g333(.A1(new_n758), .A2(G1986), .ZN(new_n759));
  NOR2_X1   g334(.A1(new_n758), .A2(G1986), .ZN(new_n760));
  NAND2_X1  g335(.A1(new_n684), .A2(G25), .ZN(new_n761));
  XNOR2_X1  g336(.A(new_n761), .B(KEYINPUT89), .ZN(new_n762));
  NAND2_X1  g337(.A1(new_n468), .A2(G131), .ZN(new_n763));
  NAND2_X1  g338(.A1(new_n486), .A2(G119), .ZN(new_n764));
  NOR2_X1   g339(.A1(new_n482), .A2(G107), .ZN(new_n765));
  OAI21_X1  g340(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n766));
  OAI211_X1 g341(.A(new_n763), .B(new_n764), .C1(new_n765), .C2(new_n766), .ZN(new_n767));
  AOI21_X1  g342(.A(new_n762), .B1(new_n767), .B2(G29), .ZN(new_n768));
  XOR2_X1   g343(.A(KEYINPUT35), .B(G1991), .Z(new_n769));
  XOR2_X1   g344(.A(new_n769), .B(KEYINPUT90), .Z(new_n770));
  XNOR2_X1  g345(.A(new_n768), .B(new_n770), .ZN(new_n771));
  NOR2_X1   g346(.A1(new_n760), .A2(new_n771), .ZN(new_n772));
  NAND4_X1  g347(.A1(new_n756), .A2(new_n757), .A3(new_n759), .A4(new_n772), .ZN(new_n773));
  XNOR2_X1  g348(.A(new_n773), .B(KEYINPUT36), .ZN(new_n774));
  NAND2_X1  g349(.A1(new_n740), .A2(KEYINPUT103), .ZN(new_n775));
  NAND2_X1  g350(.A1(new_n688), .A2(G19), .ZN(new_n776));
  OAI21_X1  g351(.A(new_n776), .B1(new_n551), .B2(new_n688), .ZN(new_n777));
  XOR2_X1   g352(.A(new_n777), .B(G1341), .Z(new_n778));
  NOR2_X1   g353(.A1(new_n598), .A2(new_n688), .ZN(new_n779));
  AOI21_X1  g354(.A(new_n779), .B1(G4), .B2(new_n688), .ZN(new_n780));
  INV_X1    g355(.A(G1348), .ZN(new_n781));
  OAI21_X1  g356(.A(new_n778), .B1(new_n780), .B2(new_n781), .ZN(new_n782));
  NAND2_X1  g357(.A1(new_n684), .A2(G26), .ZN(new_n783));
  XOR2_X1   g358(.A(new_n783), .B(KEYINPUT28), .Z(new_n784));
  NAND2_X1  g359(.A1(new_n468), .A2(G140), .ZN(new_n785));
  INV_X1    g360(.A(KEYINPUT92), .ZN(new_n786));
  XNOR2_X1  g361(.A(new_n785), .B(new_n786), .ZN(new_n787));
  OAI21_X1  g362(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n788));
  INV_X1    g363(.A(G116), .ZN(new_n789));
  AOI21_X1  g364(.A(new_n788), .B1(new_n789), .B2(G2105), .ZN(new_n790));
  AOI21_X1  g365(.A(new_n790), .B1(G128), .B2(new_n486), .ZN(new_n791));
  NAND2_X1  g366(.A1(new_n787), .A2(new_n791), .ZN(new_n792));
  AOI21_X1  g367(.A(new_n784), .B1(new_n792), .B2(G29), .ZN(new_n793));
  INV_X1    g368(.A(G2067), .ZN(new_n794));
  XNOR2_X1  g369(.A(new_n793), .B(new_n794), .ZN(new_n795));
  NOR2_X1   g370(.A1(G29), .A2(G35), .ZN(new_n796));
  AOI21_X1  g371(.A(new_n796), .B1(G162), .B2(G29), .ZN(new_n797));
  XNOR2_X1  g372(.A(new_n797), .B(KEYINPUT29), .ZN(new_n798));
  AOI21_X1  g373(.A(new_n795), .B1(G2090), .B2(new_n798), .ZN(new_n799));
  NAND2_X1  g374(.A1(new_n688), .A2(G20), .ZN(new_n800));
  XOR2_X1   g375(.A(new_n800), .B(KEYINPUT23), .Z(new_n801));
  AOI21_X1  g376(.A(new_n801), .B1(G299), .B2(G16), .ZN(new_n802));
  XNOR2_X1  g377(.A(new_n802), .B(G1956), .ZN(new_n803));
  OAI211_X1 g378(.A(new_n799), .B(new_n803), .C1(G2090), .C2(new_n798), .ZN(new_n804));
  AOI211_X1 g379(.A(new_n782), .B(new_n804), .C1(new_n781), .C2(new_n780), .ZN(new_n805));
  NAND4_X1  g380(.A1(new_n741), .A2(new_n774), .A3(new_n775), .A4(new_n805), .ZN(G150));
  INV_X1    g381(.A(G150), .ZN(G311));
  NAND2_X1  g382(.A1(new_n598), .A2(G559), .ZN(new_n808));
  XNOR2_X1  g383(.A(new_n808), .B(KEYINPUT38), .ZN(new_n809));
  NAND2_X1  g384(.A1(new_n525), .A2(G93), .ZN(new_n810));
  NAND2_X1  g385(.A1(new_n518), .A2(G55), .ZN(new_n811));
  AOI22_X1  g386(.A1(new_n523), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n812));
  OAI211_X1 g387(.A(new_n810), .B(new_n811), .C1(new_n512), .C2(new_n812), .ZN(new_n813));
  XNOR2_X1  g388(.A(new_n551), .B(new_n813), .ZN(new_n814));
  XNOR2_X1  g389(.A(new_n809), .B(new_n814), .ZN(new_n815));
  AND2_X1   g390(.A1(new_n815), .A2(KEYINPUT39), .ZN(new_n816));
  NOR2_X1   g391(.A1(new_n815), .A2(KEYINPUT39), .ZN(new_n817));
  NOR3_X1   g392(.A1(new_n816), .A2(new_n817), .A3(G860), .ZN(new_n818));
  NAND2_X1  g393(.A1(new_n813), .A2(G860), .ZN(new_n819));
  XNOR2_X1  g394(.A(new_n819), .B(KEYINPUT37), .ZN(new_n820));
  OR2_X1    g395(.A1(new_n818), .A2(new_n820), .ZN(G145));
  NOR2_X1   g396(.A1(new_n728), .A2(KEYINPUT104), .ZN(new_n822));
  XNOR2_X1  g397(.A(new_n792), .B(G164), .ZN(new_n823));
  INV_X1    g398(.A(new_n703), .ZN(new_n824));
  AOI21_X1  g399(.A(new_n822), .B1(new_n823), .B2(new_n824), .ZN(new_n825));
  OAI21_X1  g400(.A(new_n825), .B1(new_n824), .B2(new_n823), .ZN(new_n826));
  NAND2_X1  g401(.A1(new_n728), .A2(KEYINPUT104), .ZN(new_n827));
  XNOR2_X1  g402(.A(new_n826), .B(new_n827), .ZN(new_n828));
  NAND2_X1  g403(.A1(new_n486), .A2(G130), .ZN(new_n829));
  NOR2_X1   g404(.A1(new_n482), .A2(G118), .ZN(new_n830));
  OAI21_X1  g405(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n831));
  OAI21_X1  g406(.A(new_n829), .B1(new_n830), .B2(new_n831), .ZN(new_n832));
  AOI21_X1  g407(.A(new_n832), .B1(G142), .B2(new_n468), .ZN(new_n833));
  XOR2_X1   g408(.A(new_n833), .B(new_n767), .Z(new_n834));
  XOR2_X1   g409(.A(new_n834), .B(new_n621), .Z(new_n835));
  XNOR2_X1  g410(.A(new_n828), .B(new_n835), .ZN(new_n836));
  XNOR2_X1  g411(.A(new_n479), .B(new_n490), .ZN(new_n837));
  XNOR2_X1  g412(.A(new_n617), .B(new_n837), .ZN(new_n838));
  AOI21_X1  g413(.A(G37), .B1(new_n836), .B2(new_n838), .ZN(new_n839));
  OAI21_X1  g414(.A(new_n839), .B1(new_n838), .B2(new_n836), .ZN(new_n840));
  XNOR2_X1  g415(.A(new_n840), .B(KEYINPUT40), .ZN(G395));
  NAND2_X1  g416(.A1(new_n813), .A2(new_n601), .ZN(new_n842));
  XNOR2_X1  g417(.A(G290), .B(G305), .ZN(new_n843));
  XOR2_X1   g418(.A(G303), .B(G288), .Z(new_n844));
  XOR2_X1   g419(.A(new_n843), .B(new_n844), .Z(new_n845));
  NAND2_X1  g420(.A1(new_n845), .A2(KEYINPUT42), .ZN(new_n846));
  XNOR2_X1  g421(.A(new_n846), .B(KEYINPUT106), .ZN(new_n847));
  XNOR2_X1  g422(.A(new_n843), .B(new_n844), .ZN(new_n848));
  INV_X1    g423(.A(KEYINPUT42), .ZN(new_n849));
  NAND2_X1  g424(.A1(new_n848), .A2(new_n849), .ZN(new_n850));
  XNOR2_X1  g425(.A(new_n850), .B(KEYINPUT107), .ZN(new_n851));
  NAND2_X1  g426(.A1(new_n847), .A2(new_n851), .ZN(new_n852));
  OR3_X1    g427(.A1(new_n598), .A2(KEYINPUT105), .A3(G299), .ZN(new_n853));
  OAI21_X1  g428(.A(KEYINPUT105), .B1(new_n598), .B2(G299), .ZN(new_n854));
  NAND2_X1  g429(.A1(new_n598), .A2(G299), .ZN(new_n855));
  NAND3_X1  g430(.A1(new_n853), .A2(new_n854), .A3(new_n855), .ZN(new_n856));
  INV_X1    g431(.A(new_n856), .ZN(new_n857));
  XNOR2_X1  g432(.A(new_n608), .B(new_n814), .ZN(new_n858));
  NOR2_X1   g433(.A1(new_n857), .A2(new_n858), .ZN(new_n859));
  INV_X1    g434(.A(KEYINPUT41), .ZN(new_n860));
  XNOR2_X1  g435(.A(new_n856), .B(new_n860), .ZN(new_n861));
  AOI21_X1  g436(.A(new_n859), .B1(new_n861), .B2(new_n858), .ZN(new_n862));
  NAND2_X1  g437(.A1(new_n852), .A2(new_n862), .ZN(new_n863));
  INV_X1    g438(.A(new_n862), .ZN(new_n864));
  NAND3_X1  g439(.A1(new_n847), .A2(new_n864), .A3(new_n851), .ZN(new_n865));
  AND2_X1   g440(.A1(new_n863), .A2(new_n865), .ZN(new_n866));
  OAI21_X1  g441(.A(new_n842), .B1(new_n866), .B2(new_n601), .ZN(G295));
  INV_X1    g442(.A(KEYINPUT108), .ZN(new_n868));
  OAI211_X1 g443(.A(new_n868), .B(new_n842), .C1(new_n866), .C2(new_n601), .ZN(new_n869));
  AOI21_X1  g444(.A(new_n601), .B1(new_n863), .B2(new_n865), .ZN(new_n870));
  INV_X1    g445(.A(new_n842), .ZN(new_n871));
  OAI21_X1  g446(.A(KEYINPUT108), .B1(new_n870), .B2(new_n871), .ZN(new_n872));
  NAND2_X1  g447(.A1(new_n869), .A2(new_n872), .ZN(G331));
  OR2_X1    g448(.A1(new_n814), .A2(G301), .ZN(new_n874));
  NAND2_X1  g449(.A1(new_n814), .A2(G301), .ZN(new_n875));
  NAND2_X1  g450(.A1(new_n874), .A2(new_n875), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n876), .A2(G286), .ZN(new_n877));
  NAND3_X1  g452(.A1(new_n874), .A2(G168), .A3(new_n875), .ZN(new_n878));
  AOI21_X1  g453(.A(new_n857), .B1(new_n877), .B2(new_n878), .ZN(new_n879));
  AND2_X1   g454(.A1(new_n877), .A2(new_n878), .ZN(new_n880));
  AOI21_X1  g455(.A(new_n879), .B1(new_n861), .B2(new_n880), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n881), .A2(new_n845), .ZN(new_n882));
  INV_X1    g457(.A(G37), .ZN(new_n883));
  NAND2_X1  g458(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  NAND3_X1  g459(.A1(new_n857), .A2(KEYINPUT109), .A3(KEYINPUT41), .ZN(new_n885));
  OAI211_X1 g460(.A(new_n880), .B(new_n885), .C1(new_n861), .C2(KEYINPUT109), .ZN(new_n886));
  INV_X1    g461(.A(new_n879), .ZN(new_n887));
  AOI21_X1  g462(.A(new_n845), .B1(new_n886), .B2(new_n887), .ZN(new_n888));
  INV_X1    g463(.A(KEYINPUT43), .ZN(new_n889));
  NOR3_X1   g464(.A1(new_n884), .A2(new_n888), .A3(new_n889), .ZN(new_n890));
  OR2_X1    g465(.A1(new_n881), .A2(new_n845), .ZN(new_n891));
  AOI21_X1  g466(.A(G37), .B1(new_n881), .B2(new_n845), .ZN(new_n892));
  AOI21_X1  g467(.A(KEYINPUT43), .B1(new_n891), .B2(new_n892), .ZN(new_n893));
  OAI21_X1  g468(.A(KEYINPUT44), .B1(new_n890), .B2(new_n893), .ZN(new_n894));
  NOR3_X1   g469(.A1(new_n884), .A2(new_n888), .A3(KEYINPUT43), .ZN(new_n895));
  AOI21_X1  g470(.A(new_n889), .B1(new_n891), .B2(new_n892), .ZN(new_n896));
  NOR2_X1   g471(.A1(new_n895), .A2(new_n896), .ZN(new_n897));
  OAI21_X1  g472(.A(new_n894), .B1(new_n897), .B2(KEYINPUT44), .ZN(G397));
  INV_X1    g473(.A(G1384), .ZN(new_n899));
  AOI21_X1  g474(.A(KEYINPUT45), .B1(new_n507), .B2(new_n899), .ZN(new_n900));
  INV_X1    g475(.A(new_n900), .ZN(new_n901));
  XNOR2_X1  g476(.A(KEYINPUT110), .B(G40), .ZN(new_n902));
  INV_X1    g477(.A(new_n902), .ZN(new_n903));
  NAND3_X1  g478(.A1(new_n471), .A2(new_n478), .A3(new_n903), .ZN(new_n904));
  NOR2_X1   g479(.A1(new_n901), .A2(new_n904), .ZN(new_n905));
  XNOR2_X1  g480(.A(new_n792), .B(G2067), .ZN(new_n906));
  OAI21_X1  g481(.A(new_n905), .B1(new_n906), .B2(new_n824), .ZN(new_n907));
  INV_X1    g482(.A(G1996), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n905), .A2(new_n908), .ZN(new_n909));
  XNOR2_X1  g484(.A(new_n909), .B(KEYINPUT111), .ZN(new_n910));
  AND3_X1   g485(.A1(new_n910), .A2(KEYINPUT127), .A3(KEYINPUT46), .ZN(new_n911));
  AOI21_X1  g486(.A(KEYINPUT127), .B1(new_n910), .B2(KEYINPUT46), .ZN(new_n912));
  OAI221_X1 g487(.A(new_n907), .B1(KEYINPUT46), .B2(new_n910), .C1(new_n911), .C2(new_n912), .ZN(new_n913));
  XOR2_X1   g488(.A(new_n913), .B(KEYINPUT47), .Z(new_n914));
  INV_X1    g489(.A(new_n906), .ZN(new_n915));
  OAI21_X1  g490(.A(new_n915), .B1(new_n908), .B2(new_n703), .ZN(new_n916));
  AOI22_X1  g491(.A1(new_n910), .A2(new_n703), .B1(new_n916), .B2(new_n905), .ZN(new_n917));
  INV_X1    g492(.A(new_n769), .ZN(new_n918));
  AND2_X1   g493(.A1(new_n767), .A2(new_n918), .ZN(new_n919));
  NOR2_X1   g494(.A1(new_n767), .A2(new_n918), .ZN(new_n920));
  OAI21_X1  g495(.A(new_n905), .B1(new_n919), .B2(new_n920), .ZN(new_n921));
  AND2_X1   g496(.A1(new_n917), .A2(new_n921), .ZN(new_n922));
  NOR2_X1   g497(.A1(G290), .A2(G1986), .ZN(new_n923));
  NAND2_X1  g498(.A1(new_n923), .A2(new_n905), .ZN(new_n924));
  XNOR2_X1  g499(.A(new_n924), .B(KEYINPUT48), .ZN(new_n925));
  NAND2_X1  g500(.A1(new_n922), .A2(new_n925), .ZN(new_n926));
  INV_X1    g501(.A(new_n905), .ZN(new_n927));
  NOR2_X1   g502(.A1(new_n792), .A2(G2067), .ZN(new_n928));
  AOI21_X1  g503(.A(new_n928), .B1(new_n917), .B2(new_n920), .ZN(new_n929));
  OAI21_X1  g504(.A(new_n926), .B1(new_n927), .B2(new_n929), .ZN(new_n930));
  NOR2_X1   g505(.A1(new_n914), .A2(new_n930), .ZN(new_n931));
  INV_X1    g506(.A(G1956), .ZN(new_n932));
  INV_X1    g507(.A(KEYINPUT50), .ZN(new_n933));
  AND3_X1   g508(.A1(new_n496), .A2(KEYINPUT4), .A3(new_n498), .ZN(new_n934));
  NAND2_X1  g509(.A1(new_n506), .A2(new_n501), .ZN(new_n935));
  OAI21_X1  g510(.A(new_n899), .B1(new_n934), .B2(new_n935), .ZN(new_n936));
  INV_X1    g511(.A(KEYINPUT113), .ZN(new_n937));
  NAND2_X1  g512(.A1(new_n936), .A2(new_n937), .ZN(new_n938));
  NAND3_X1  g513(.A1(new_n507), .A2(KEYINPUT113), .A3(new_n899), .ZN(new_n939));
  AOI21_X1  g514(.A(new_n933), .B1(new_n938), .B2(new_n939), .ZN(new_n940));
  OAI211_X1 g515(.A(G126), .B(G2105), .C1(new_n465), .C2(new_n466), .ZN(new_n941));
  OR2_X1    g516(.A1(G102), .A2(G2105), .ZN(new_n942));
  NAND3_X1  g517(.A1(new_n942), .A2(new_n503), .A3(G2104), .ZN(new_n943));
  NAND2_X1  g518(.A1(new_n941), .A2(new_n943), .ZN(new_n944));
  AOI21_X1  g519(.A(KEYINPUT72), .B1(new_n497), .B2(new_n493), .ZN(new_n945));
  AOI21_X1  g520(.A(new_n944), .B1(new_n500), .B2(new_n945), .ZN(new_n946));
  AOI21_X1  g521(.A(G1384), .B1(new_n946), .B2(new_n499), .ZN(new_n947));
  AOI21_X1  g522(.A(new_n904), .B1(new_n947), .B2(new_n933), .ZN(new_n948));
  INV_X1    g523(.A(new_n948), .ZN(new_n949));
  OAI21_X1  g524(.A(new_n932), .B1(new_n940), .B2(new_n949), .ZN(new_n950));
  NAND3_X1  g525(.A1(new_n507), .A2(KEYINPUT45), .A3(new_n899), .ZN(new_n951));
  INV_X1    g526(.A(new_n904), .ZN(new_n952));
  NAND2_X1  g527(.A1(new_n951), .A2(new_n952), .ZN(new_n953));
  XNOR2_X1  g528(.A(KEYINPUT56), .B(G2072), .ZN(new_n954));
  INV_X1    g529(.A(new_n954), .ZN(new_n955));
  NOR3_X1   g530(.A1(new_n953), .A2(new_n900), .A3(new_n955), .ZN(new_n956));
  INV_X1    g531(.A(new_n956), .ZN(new_n957));
  NAND2_X1  g532(.A1(G299), .A2(KEYINPUT57), .ZN(new_n958));
  INV_X1    g533(.A(KEYINPUT57), .ZN(new_n959));
  NAND3_X1  g534(.A1(new_n558), .A2(new_n562), .A3(new_n959), .ZN(new_n960));
  NAND2_X1  g535(.A1(new_n958), .A2(new_n960), .ZN(new_n961));
  INV_X1    g536(.A(new_n961), .ZN(new_n962));
  NAND4_X1  g537(.A1(new_n950), .A2(new_n957), .A3(KEYINPUT124), .A4(new_n962), .ZN(new_n963));
  AOI211_X1 g538(.A(new_n937), .B(G1384), .C1(new_n946), .C2(new_n499), .ZN(new_n964));
  AOI21_X1  g539(.A(KEYINPUT113), .B1(new_n507), .B2(new_n899), .ZN(new_n965));
  OAI21_X1  g540(.A(KEYINPUT50), .B1(new_n964), .B2(new_n965), .ZN(new_n966));
  AOI21_X1  g541(.A(G1956), .B1(new_n966), .B2(new_n948), .ZN(new_n967));
  OAI21_X1  g542(.A(new_n961), .B1(new_n967), .B2(new_n956), .ZN(new_n968));
  AND3_X1   g543(.A1(new_n963), .A2(new_n968), .A3(KEYINPUT61), .ZN(new_n969));
  NOR3_X1   g544(.A1(new_n967), .A2(new_n961), .A3(new_n956), .ZN(new_n970));
  OR2_X1    g545(.A1(new_n970), .A2(KEYINPUT124), .ZN(new_n971));
  NAND3_X1  g546(.A1(new_n938), .A2(new_n952), .A3(new_n939), .ZN(new_n972));
  XOR2_X1   g547(.A(KEYINPUT58), .B(G1341), .Z(new_n973));
  NAND3_X1  g548(.A1(new_n972), .A2(KEYINPUT123), .A3(new_n973), .ZN(new_n974));
  INV_X1    g549(.A(new_n953), .ZN(new_n975));
  NAND3_X1  g550(.A1(new_n975), .A2(new_n908), .A3(new_n901), .ZN(new_n976));
  NAND2_X1  g551(.A1(new_n974), .A2(new_n976), .ZN(new_n977));
  AOI21_X1  g552(.A(KEYINPUT123), .B1(new_n972), .B2(new_n973), .ZN(new_n978));
  OAI21_X1  g553(.A(new_n551), .B1(new_n977), .B2(new_n978), .ZN(new_n979));
  NAND2_X1  g554(.A1(new_n979), .A2(KEYINPUT59), .ZN(new_n980));
  INV_X1    g555(.A(KEYINPUT59), .ZN(new_n981));
  OAI211_X1 g556(.A(new_n981), .B(new_n551), .C1(new_n977), .C2(new_n978), .ZN(new_n982));
  AOI22_X1  g557(.A1(new_n969), .A2(new_n971), .B1(new_n980), .B2(new_n982), .ZN(new_n983));
  INV_X1    g558(.A(KEYINPUT60), .ZN(new_n984));
  INV_X1    g559(.A(KEYINPUT115), .ZN(new_n985));
  AOI21_X1  g560(.A(new_n985), .B1(new_n936), .B2(KEYINPUT50), .ZN(new_n986));
  AOI211_X1 g561(.A(KEYINPUT115), .B(new_n933), .C1(new_n507), .C2(new_n899), .ZN(new_n987));
  NOR2_X1   g562(.A1(new_n986), .A2(new_n987), .ZN(new_n988));
  NAND3_X1  g563(.A1(new_n938), .A2(new_n933), .A3(new_n939), .ZN(new_n989));
  NAND2_X1  g564(.A1(new_n989), .A2(KEYINPUT114), .ZN(new_n990));
  INV_X1    g565(.A(KEYINPUT114), .ZN(new_n991));
  NAND4_X1  g566(.A1(new_n938), .A2(new_n991), .A3(new_n933), .A4(new_n939), .ZN(new_n992));
  AOI21_X1  g567(.A(new_n988), .B1(new_n990), .B2(new_n992), .ZN(new_n993));
  AOI21_X1  g568(.A(G1348), .B1(new_n993), .B2(new_n952), .ZN(new_n994));
  NOR2_X1   g569(.A1(new_n972), .A2(G2067), .ZN(new_n995));
  OAI21_X1  g570(.A(new_n984), .B1(new_n994), .B2(new_n995), .ZN(new_n996));
  INV_X1    g571(.A(new_n995), .ZN(new_n997));
  INV_X1    g572(.A(new_n986), .ZN(new_n998));
  INV_X1    g573(.A(new_n987), .ZN(new_n999));
  AOI221_X4 g574(.A(new_n904), .B1(new_n998), .B2(new_n999), .C1(new_n990), .C2(new_n992), .ZN(new_n1000));
  OAI211_X1 g575(.A(KEYINPUT60), .B(new_n997), .C1(new_n1000), .C2(G1348), .ZN(new_n1001));
  NAND3_X1  g576(.A1(new_n996), .A2(new_n1001), .A3(new_n598), .ZN(new_n1002));
  NOR2_X1   g577(.A1(new_n994), .A2(new_n995), .ZN(new_n1003));
  INV_X1    g578(.A(new_n598), .ZN(new_n1004));
  NAND3_X1  g579(.A1(new_n1003), .A2(KEYINPUT60), .A3(new_n1004), .ZN(new_n1005));
  INV_X1    g580(.A(KEYINPUT122), .ZN(new_n1006));
  NAND2_X1  g581(.A1(new_n966), .A2(new_n948), .ZN(new_n1007));
  AOI21_X1  g582(.A(new_n956), .B1(new_n1007), .B2(new_n932), .ZN(new_n1008));
  AOI21_X1  g583(.A(new_n1006), .B1(new_n1008), .B2(new_n962), .ZN(new_n1009));
  NOR4_X1   g584(.A1(new_n967), .A2(new_n956), .A3(KEYINPUT122), .A4(new_n961), .ZN(new_n1010));
  OAI21_X1  g585(.A(new_n968), .B1(new_n1009), .B2(new_n1010), .ZN(new_n1011));
  INV_X1    g586(.A(KEYINPUT61), .ZN(new_n1012));
  NAND2_X1  g587(.A1(new_n1011), .A2(new_n1012), .ZN(new_n1013));
  NAND4_X1  g588(.A1(new_n983), .A2(new_n1002), .A3(new_n1005), .A4(new_n1013), .ZN(new_n1014));
  OAI21_X1  g589(.A(new_n968), .B1(new_n1003), .B2(new_n1004), .ZN(new_n1015));
  OAI21_X1  g590(.A(new_n1015), .B1(new_n1009), .B2(new_n1010), .ZN(new_n1016));
  NAND2_X1  g591(.A1(new_n1014), .A2(new_n1016), .ZN(new_n1017));
  INV_X1    g592(.A(KEYINPUT49), .ZN(new_n1018));
  INV_X1    g593(.A(G1981), .ZN(new_n1019));
  NAND3_X1  g594(.A1(new_n575), .A2(new_n1019), .A3(new_n578), .ZN(new_n1020));
  INV_X1    g595(.A(new_n1020), .ZN(new_n1021));
  AOI21_X1  g596(.A(new_n1019), .B1(new_n575), .B2(new_n578), .ZN(new_n1022));
  OAI21_X1  g597(.A(new_n1018), .B1(new_n1021), .B2(new_n1022), .ZN(new_n1023));
  NAND2_X1  g598(.A1(G305), .A2(G1981), .ZN(new_n1024));
  NAND3_X1  g599(.A1(new_n1024), .A2(KEYINPUT49), .A3(new_n1020), .ZN(new_n1025));
  NAND4_X1  g600(.A1(new_n1023), .A2(new_n972), .A3(new_n1025), .A4(G8), .ZN(new_n1026));
  NAND2_X1  g601(.A1(new_n747), .A2(G1976), .ZN(new_n1027));
  XOR2_X1   g602(.A(KEYINPUT119), .B(G1976), .Z(new_n1028));
  AOI21_X1  g603(.A(KEYINPUT52), .B1(G288), .B2(new_n1028), .ZN(new_n1029));
  NAND4_X1  g604(.A1(new_n972), .A2(G8), .A3(new_n1027), .A4(new_n1029), .ZN(new_n1030));
  NAND2_X1  g605(.A1(new_n1026), .A2(new_n1030), .ZN(new_n1031));
  INV_X1    g606(.A(new_n1031), .ZN(new_n1032));
  NAND3_X1  g607(.A1(new_n972), .A2(G8), .A3(new_n1027), .ZN(new_n1033));
  INV_X1    g608(.A(KEYINPUT118), .ZN(new_n1034));
  AND3_X1   g609(.A1(new_n1033), .A2(new_n1034), .A3(KEYINPUT52), .ZN(new_n1035));
  AOI21_X1  g610(.A(new_n1034), .B1(new_n1033), .B2(KEYINPUT52), .ZN(new_n1036));
  OAI21_X1  g611(.A(new_n1032), .B1(new_n1035), .B2(new_n1036), .ZN(new_n1037));
  NAND2_X1  g612(.A1(G303), .A2(G8), .ZN(new_n1038));
  INV_X1    g613(.A(KEYINPUT116), .ZN(new_n1039));
  OAI21_X1  g614(.A(KEYINPUT117), .B1(new_n1038), .B2(new_n1039), .ZN(new_n1040));
  INV_X1    g615(.A(KEYINPUT117), .ZN(new_n1041));
  NAND4_X1  g616(.A1(G303), .A2(KEYINPUT116), .A3(new_n1041), .A4(G8), .ZN(new_n1042));
  NAND2_X1  g617(.A1(new_n1040), .A2(new_n1042), .ZN(new_n1043));
  NAND2_X1  g618(.A1(new_n1038), .A2(new_n1039), .ZN(new_n1044));
  NAND2_X1  g619(.A1(new_n1044), .A2(KEYINPUT55), .ZN(new_n1045));
  XNOR2_X1  g620(.A(new_n1043), .B(new_n1045), .ZN(new_n1046));
  INV_X1    g621(.A(G8), .ZN(new_n1047));
  NAND2_X1  g622(.A1(new_n998), .A2(new_n999), .ZN(new_n1048));
  NOR2_X1   g623(.A1(new_n904), .A2(G2090), .ZN(new_n1049));
  NOR2_X1   g624(.A1(new_n964), .A2(new_n965), .ZN(new_n1050));
  AOI21_X1  g625(.A(new_n991), .B1(new_n1050), .B2(new_n933), .ZN(new_n1051));
  INV_X1    g626(.A(new_n992), .ZN(new_n1052));
  OAI211_X1 g627(.A(new_n1048), .B(new_n1049), .C1(new_n1051), .C2(new_n1052), .ZN(new_n1053));
  NOR2_X1   g628(.A1(new_n953), .A2(new_n900), .ZN(new_n1054));
  NOR2_X1   g629(.A1(new_n1054), .A2(G1971), .ZN(new_n1055));
  INV_X1    g630(.A(new_n1055), .ZN(new_n1056));
  AOI21_X1  g631(.A(new_n1047), .B1(new_n1053), .B2(new_n1056), .ZN(new_n1057));
  AOI21_X1  g632(.A(new_n1037), .B1(new_n1046), .B2(new_n1057), .ZN(new_n1058));
  INV_X1    g633(.A(KEYINPUT125), .ZN(new_n1059));
  OAI21_X1  g634(.A(new_n1059), .B1(new_n1000), .B2(G1961), .ZN(new_n1060));
  NAND2_X1  g635(.A1(new_n993), .A2(new_n952), .ZN(new_n1061));
  INV_X1    g636(.A(G1961), .ZN(new_n1062));
  NAND3_X1  g637(.A1(new_n1061), .A2(KEYINPUT125), .A3(new_n1062), .ZN(new_n1063));
  INV_X1    g638(.A(KEYINPUT53), .ZN(new_n1064));
  INV_X1    g639(.A(new_n1054), .ZN(new_n1065));
  OAI21_X1  g640(.A(new_n1064), .B1(new_n1065), .B2(G2078), .ZN(new_n1066));
  XOR2_X1   g641(.A(G301), .B(KEYINPUT54), .Z(new_n1067));
  NOR2_X1   g642(.A1(new_n1064), .A2(G2078), .ZN(new_n1068));
  AND3_X1   g643(.A1(G160), .A2(G40), .A3(new_n1068), .ZN(new_n1069));
  NAND3_X1  g644(.A1(new_n1069), .A2(new_n901), .A3(new_n951), .ZN(new_n1070));
  AND3_X1   g645(.A1(new_n1066), .A2(new_n1067), .A3(new_n1070), .ZN(new_n1071));
  NAND3_X1  g646(.A1(new_n1060), .A2(new_n1063), .A3(new_n1071), .ZN(new_n1072));
  XOR2_X1   g647(.A(new_n1043), .B(new_n1045), .Z(new_n1073));
  AOI21_X1  g648(.A(G2090), .B1(new_n1007), .B2(KEYINPUT120), .ZN(new_n1074));
  OR3_X1    g649(.A1(new_n940), .A2(new_n949), .A3(KEYINPUT120), .ZN(new_n1075));
  AOI21_X1  g650(.A(new_n1055), .B1(new_n1074), .B2(new_n1075), .ZN(new_n1076));
  OAI21_X1  g651(.A(new_n1073), .B1(new_n1076), .B2(new_n1047), .ZN(new_n1077));
  INV_X1    g652(.A(new_n1067), .ZN(new_n1078));
  AOI21_X1  g653(.A(G1961), .B1(new_n993), .B2(new_n952), .ZN(new_n1079));
  OAI21_X1  g654(.A(new_n975), .B1(new_n1050), .B2(KEYINPUT45), .ZN(new_n1080));
  OR2_X1    g655(.A1(new_n1064), .A2(G2078), .ZN(new_n1081));
  OAI21_X1  g656(.A(new_n1066), .B1(new_n1080), .B2(new_n1081), .ZN(new_n1082));
  OAI21_X1  g657(.A(new_n1078), .B1(new_n1079), .B2(new_n1082), .ZN(new_n1083));
  NAND4_X1  g658(.A1(new_n1058), .A2(new_n1072), .A3(new_n1077), .A4(new_n1083), .ZN(new_n1084));
  NOR2_X1   g659(.A1(new_n904), .A2(G2084), .ZN(new_n1085));
  OAI211_X1 g660(.A(new_n1048), .B(new_n1085), .C1(new_n1051), .C2(new_n1052), .ZN(new_n1086));
  NAND2_X1  g661(.A1(new_n1080), .A2(new_n736), .ZN(new_n1087));
  NAND3_X1  g662(.A1(new_n1086), .A2(G168), .A3(new_n1087), .ZN(new_n1088));
  INV_X1    g663(.A(KEYINPUT51), .ZN(new_n1089));
  AND3_X1   g664(.A1(new_n1088), .A2(new_n1089), .A3(G8), .ZN(new_n1090));
  NAND2_X1  g665(.A1(new_n1086), .A2(new_n1087), .ZN(new_n1091));
  NAND2_X1  g666(.A1(new_n1091), .A2(G286), .ZN(new_n1092));
  NAND3_X1  g667(.A1(new_n1092), .A2(G8), .A3(new_n1088), .ZN(new_n1093));
  AOI21_X1  g668(.A(new_n1090), .B1(new_n1093), .B2(KEYINPUT51), .ZN(new_n1094));
  NOR2_X1   g669(.A1(new_n1084), .A2(new_n1094), .ZN(new_n1095));
  NAND2_X1  g670(.A1(new_n1017), .A2(new_n1095), .ZN(new_n1096));
  AOI22_X1  g671(.A1(new_n993), .A2(new_n1085), .B1(new_n736), .B2(new_n1080), .ZN(new_n1097));
  AOI21_X1  g672(.A(new_n1047), .B1(new_n1097), .B2(G168), .ZN(new_n1098));
  AOI21_X1  g673(.A(new_n1089), .B1(new_n1098), .B2(new_n1092), .ZN(new_n1099));
  OAI21_X1  g674(.A(KEYINPUT62), .B1(new_n1099), .B2(new_n1090), .ZN(new_n1100));
  NAND2_X1  g675(.A1(new_n1093), .A2(KEYINPUT51), .ZN(new_n1101));
  INV_X1    g676(.A(KEYINPUT62), .ZN(new_n1102));
  INV_X1    g677(.A(new_n1090), .ZN(new_n1103));
  NAND3_X1  g678(.A1(new_n1101), .A2(new_n1102), .A3(new_n1103), .ZN(new_n1104));
  NAND2_X1  g679(.A1(new_n1057), .A2(new_n1046), .ZN(new_n1105));
  INV_X1    g680(.A(new_n1037), .ZN(new_n1106));
  NAND3_X1  g681(.A1(new_n1077), .A2(new_n1105), .A3(new_n1106), .ZN(new_n1107));
  OAI21_X1  g682(.A(G171), .B1(new_n1079), .B2(new_n1082), .ZN(new_n1108));
  NOR2_X1   g683(.A1(new_n1107), .A2(new_n1108), .ZN(new_n1109));
  NAND3_X1  g684(.A1(new_n1100), .A2(new_n1104), .A3(new_n1109), .ZN(new_n1110));
  NOR2_X1   g685(.A1(G288), .A2(G1976), .ZN(new_n1111));
  AND2_X1   g686(.A1(new_n1026), .A2(new_n1111), .ZN(new_n1112));
  OAI211_X1 g687(.A(G8), .B(new_n972), .C1(new_n1112), .C2(new_n1021), .ZN(new_n1113));
  OAI21_X1  g688(.A(new_n1113), .B1(new_n1105), .B2(new_n1037), .ZN(new_n1114));
  INV_X1    g689(.A(KEYINPUT63), .ZN(new_n1115));
  NOR2_X1   g690(.A1(G286), .A2(new_n1047), .ZN(new_n1116));
  AOI21_X1  g691(.A(KEYINPUT121), .B1(new_n1091), .B2(new_n1116), .ZN(new_n1117));
  INV_X1    g692(.A(KEYINPUT121), .ZN(new_n1118));
  INV_X1    g693(.A(new_n1116), .ZN(new_n1119));
  AOI211_X1 g694(.A(new_n1118), .B(new_n1119), .C1(new_n1086), .C2(new_n1087), .ZN(new_n1120));
  NOR2_X1   g695(.A1(new_n1117), .A2(new_n1120), .ZN(new_n1121));
  OAI21_X1  g696(.A(new_n1115), .B1(new_n1107), .B2(new_n1121), .ZN(new_n1122));
  OAI21_X1  g697(.A(new_n1118), .B1(new_n1097), .B2(new_n1119), .ZN(new_n1123));
  NAND3_X1  g698(.A1(new_n1091), .A2(KEYINPUT121), .A3(new_n1116), .ZN(new_n1124));
  NAND2_X1  g699(.A1(new_n1123), .A2(new_n1124), .ZN(new_n1125));
  OR2_X1    g700(.A1(new_n1057), .A2(new_n1046), .ZN(new_n1126));
  NAND4_X1  g701(.A1(new_n1125), .A2(new_n1058), .A3(KEYINPUT63), .A4(new_n1126), .ZN(new_n1127));
  AOI21_X1  g702(.A(new_n1114), .B1(new_n1122), .B2(new_n1127), .ZN(new_n1128));
  NAND3_X1  g703(.A1(new_n1096), .A2(new_n1110), .A3(new_n1128), .ZN(new_n1129));
  AND2_X1   g704(.A1(G290), .A2(G1986), .ZN(new_n1130));
  OAI21_X1  g705(.A(new_n905), .B1(new_n1130), .B2(new_n923), .ZN(new_n1131));
  NAND2_X1  g706(.A1(new_n922), .A2(new_n1131), .ZN(new_n1132));
  XOR2_X1   g707(.A(new_n1132), .B(KEYINPUT112), .Z(new_n1133));
  AND3_X1   g708(.A1(new_n1129), .A2(KEYINPUT126), .A3(new_n1133), .ZN(new_n1134));
  AOI21_X1  g709(.A(KEYINPUT126), .B1(new_n1129), .B2(new_n1133), .ZN(new_n1135));
  OAI21_X1  g710(.A(new_n931), .B1(new_n1134), .B2(new_n1135), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g711(.A(new_n463), .ZN(new_n1138));
  NOR4_X1   g712(.A1(G229), .A2(G401), .A3(new_n1138), .A4(G227), .ZN(new_n1139));
  OAI211_X1 g713(.A(new_n840), .B(new_n1139), .C1(new_n895), .C2(new_n896), .ZN(G225));
  INV_X1    g714(.A(G225), .ZN(G308));
endmodule


