//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 0 1 1 1 1 1 1 0 0 0 1 0 1 1 0 1 0 1 0 1 1 0 1 0 0 0 0 0 1 0 0 1 0 0 1 1 0 0 1 1 0 0 1 0 0 1 1 0 1 0 0 0 0 0 1 1 0 0 1 0 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:33:44 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n447, new_n449, new_n452, new_n453, new_n454, new_n457,
    new_n458, new_n459, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n483, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n521, new_n522, new_n523, new_n524, new_n525,
    new_n526, new_n527, new_n529, new_n530, new_n531, new_n532, new_n533,
    new_n534, new_n537, new_n538, new_n539, new_n540, new_n541, new_n542,
    new_n543, new_n544, new_n545, new_n546, new_n547, new_n548, new_n549,
    new_n550, new_n553, new_n554, new_n556, new_n557, new_n558, new_n559,
    new_n560, new_n561, new_n562, new_n563, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n574, new_n575, new_n576, new_n577,
    new_n578, new_n579, new_n580, new_n582, new_n583, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n596, new_n599, new_n600, new_n602, new_n603, new_n604, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n621, new_n622,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n809, new_n810, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1159, new_n1160;
  XNOR2_X1  g000(.A(KEYINPUT64), .B(G452), .ZN(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  XOR2_X1   g003(.A(KEYINPUT65), .B(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  XNOR2_X1  g020(.A(KEYINPUT66), .B(KEYINPUT1), .ZN(new_n446));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XNOR2_X1  g022(.A(new_n446), .B(new_n447), .ZN(G223));
  INV_X1    g023(.A(new_n447), .ZN(new_n449));
  NAND2_X1  g024(.A1(new_n449), .A2(G567), .ZN(G234));
  NAND2_X1  g025(.A1(new_n449), .A2(G2106), .ZN(G217));
  NOR4_X1   g026(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n452));
  XNOR2_X1  g027(.A(new_n452), .B(KEYINPUT2), .ZN(new_n453));
  NOR4_X1   g028(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n454));
  NAND2_X1  g029(.A1(new_n453), .A2(new_n454), .ZN(G261));
  INV_X1    g030(.A(G261), .ZN(G325));
  INV_X1    g031(.A(G2106), .ZN(new_n457));
  INV_X1    g032(.A(G567), .ZN(new_n458));
  OAI22_X1  g033(.A1(new_n453), .A2(new_n457), .B1(new_n458), .B2(new_n454), .ZN(new_n459));
  XOR2_X1   g034(.A(new_n459), .B(KEYINPUT67), .Z(G319));
  INV_X1    g035(.A(G2105), .ZN(new_n461));
  NAND2_X1  g036(.A1(new_n461), .A2(G2104), .ZN(new_n462));
  INV_X1    g037(.A(new_n462), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n463), .A2(G101), .ZN(new_n464));
  INV_X1    g039(.A(KEYINPUT3), .ZN(new_n465));
  INV_X1    g040(.A(G2104), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  NAND2_X1  g042(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n469), .A2(new_n461), .ZN(new_n470));
  INV_X1    g045(.A(G137), .ZN(new_n471));
  OAI21_X1  g046(.A(new_n464), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  INV_X1    g047(.A(KEYINPUT68), .ZN(new_n473));
  AND2_X1   g048(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n474));
  NOR2_X1   g049(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n475));
  OAI21_X1  g050(.A(new_n473), .B1(new_n474), .B2(new_n475), .ZN(new_n476));
  NAND3_X1  g051(.A1(new_n467), .A2(KEYINPUT68), .A3(new_n468), .ZN(new_n477));
  NAND3_X1  g052(.A1(new_n476), .A2(new_n477), .A3(G125), .ZN(new_n478));
  INV_X1    g053(.A(KEYINPUT69), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n478), .A2(new_n479), .ZN(new_n480));
  NAND4_X1  g055(.A1(new_n476), .A2(new_n477), .A3(KEYINPUT69), .A4(G125), .ZN(new_n481));
  NAND2_X1  g056(.A1(G113), .A2(G2104), .ZN(new_n482));
  NAND3_X1  g057(.A1(new_n480), .A2(new_n481), .A3(new_n482), .ZN(new_n483));
  AOI21_X1  g058(.A(new_n472), .B1(new_n483), .B2(G2105), .ZN(G160));
  NOR2_X1   g059(.A1(new_n474), .A2(new_n475), .ZN(new_n485));
  NOR2_X1   g060(.A1(new_n485), .A2(G2105), .ZN(new_n486));
  NAND2_X1  g061(.A1(new_n486), .A2(G136), .ZN(new_n487));
  NOR2_X1   g062(.A1(new_n485), .A2(new_n461), .ZN(new_n488));
  NAND2_X1  g063(.A1(new_n488), .A2(G124), .ZN(new_n489));
  NOR2_X1   g064(.A1(new_n461), .A2(G112), .ZN(new_n490));
  OAI21_X1  g065(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n491));
  OAI211_X1 g066(.A(new_n487), .B(new_n489), .C1(new_n490), .C2(new_n491), .ZN(new_n492));
  XOR2_X1   g067(.A(new_n492), .B(KEYINPUT70), .Z(G162));
  NAND2_X1  g068(.A1(new_n469), .A2(G2105), .ZN(new_n494));
  INV_X1    g069(.A(G126), .ZN(new_n495));
  NOR2_X1   g070(.A1(new_n461), .A2(G114), .ZN(new_n496));
  OAI21_X1  g071(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n497));
  OAI22_X1  g072(.A1(new_n494), .A2(new_n495), .B1(new_n496), .B2(new_n497), .ZN(new_n498));
  INV_X1    g073(.A(G138), .ZN(new_n499));
  NOR3_X1   g074(.A1(new_n499), .A2(KEYINPUT4), .A3(G2105), .ZN(new_n500));
  NAND3_X1  g075(.A1(new_n476), .A2(new_n477), .A3(new_n500), .ZN(new_n501));
  INV_X1    g076(.A(KEYINPUT71), .ZN(new_n502));
  OAI211_X1 g077(.A(G138), .B(new_n461), .C1(new_n474), .C2(new_n475), .ZN(new_n503));
  AOI22_X1  g078(.A1(new_n501), .A2(new_n502), .B1(KEYINPUT4), .B2(new_n503), .ZN(new_n504));
  NAND4_X1  g079(.A1(new_n476), .A2(new_n477), .A3(KEYINPUT71), .A4(new_n500), .ZN(new_n505));
  AOI21_X1  g080(.A(new_n498), .B1(new_n504), .B2(new_n505), .ZN(G164));
  INV_X1    g081(.A(G543), .ZN(new_n507));
  OR2_X1    g082(.A1(KEYINPUT6), .A2(G651), .ZN(new_n508));
  NAND2_X1  g083(.A1(KEYINPUT6), .A2(G651), .ZN(new_n509));
  AOI21_X1  g084(.A(new_n507), .B1(new_n508), .B2(new_n509), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n510), .A2(G50), .ZN(new_n511));
  INV_X1    g086(.A(G88), .ZN(new_n512));
  NAND2_X1  g087(.A1(new_n508), .A2(new_n509), .ZN(new_n513));
  XNOR2_X1  g088(.A(KEYINPUT5), .B(G543), .ZN(new_n514));
  NAND2_X1  g089(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  OAI21_X1  g090(.A(new_n511), .B1(new_n512), .B2(new_n515), .ZN(new_n516));
  AOI22_X1  g091(.A1(new_n514), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n517));
  INV_X1    g092(.A(G651), .ZN(new_n518));
  NOR2_X1   g093(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  NOR2_X1   g094(.A1(new_n516), .A2(new_n519), .ZN(G166));
  NAND3_X1  g095(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n521));
  XNOR2_X1  g096(.A(new_n521), .B(KEYINPUT72), .ZN(new_n522));
  XOR2_X1   g097(.A(new_n522), .B(KEYINPUT7), .Z(new_n523));
  NAND2_X1  g098(.A1(new_n510), .A2(G51), .ZN(new_n524));
  NAND3_X1  g099(.A1(new_n514), .A2(G63), .A3(G651), .ZN(new_n525));
  XNOR2_X1  g100(.A(KEYINPUT73), .B(G89), .ZN(new_n526));
  OAI211_X1 g101(.A(new_n524), .B(new_n525), .C1(new_n515), .C2(new_n526), .ZN(new_n527));
  NOR2_X1   g102(.A1(new_n523), .A2(new_n527), .ZN(G168));
  AND2_X1   g103(.A1(new_n513), .A2(new_n514), .ZN(new_n529));
  AOI22_X1  g104(.A1(new_n529), .A2(G90), .B1(G52), .B2(new_n510), .ZN(new_n530));
  INV_X1    g105(.A(KEYINPUT74), .ZN(new_n531));
  XNOR2_X1  g106(.A(new_n530), .B(new_n531), .ZN(new_n532));
  AOI22_X1  g107(.A1(new_n514), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n533));
  OR2_X1    g108(.A1(new_n533), .A2(new_n518), .ZN(new_n534));
  NAND2_X1  g109(.A1(new_n532), .A2(new_n534), .ZN(G301));
  INV_X1    g110(.A(G301), .ZN(G171));
  AND2_X1   g111(.A1(KEYINPUT5), .A2(G543), .ZN(new_n537));
  NOR2_X1   g112(.A1(KEYINPUT5), .A2(G543), .ZN(new_n538));
  NOR2_X1   g113(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  INV_X1    g114(.A(G56), .ZN(new_n540));
  NOR2_X1   g115(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  AND2_X1   g116(.A1(G68), .A2(G543), .ZN(new_n542));
  OAI21_X1  g117(.A(G651), .B1(new_n541), .B2(new_n542), .ZN(new_n543));
  NAND2_X1  g118(.A1(new_n543), .A2(KEYINPUT75), .ZN(new_n544));
  INV_X1    g119(.A(KEYINPUT75), .ZN(new_n545));
  OAI211_X1 g120(.A(new_n545), .B(G651), .C1(new_n541), .C2(new_n542), .ZN(new_n546));
  AOI22_X1  g121(.A1(new_n529), .A2(G81), .B1(G43), .B2(new_n510), .ZN(new_n547));
  NAND3_X1  g122(.A1(new_n544), .A2(new_n546), .A3(new_n547), .ZN(new_n548));
  XNOR2_X1  g123(.A(new_n548), .B(KEYINPUT76), .ZN(new_n549));
  INV_X1    g124(.A(new_n549), .ZN(new_n550));
  NAND2_X1  g125(.A1(new_n550), .A2(G860), .ZN(G153));
  NAND4_X1  g126(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g127(.A1(G1), .A2(G3), .ZN(new_n553));
  XNOR2_X1  g128(.A(new_n553), .B(KEYINPUT8), .ZN(new_n554));
  NAND4_X1  g129(.A1(G319), .A2(G483), .A3(G661), .A4(new_n554), .ZN(G188));
  NAND2_X1  g130(.A1(new_n510), .A2(G53), .ZN(new_n556));
  INV_X1    g131(.A(KEYINPUT9), .ZN(new_n557));
  NOR2_X1   g132(.A1(new_n557), .A2(KEYINPUT77), .ZN(new_n558));
  XNOR2_X1  g133(.A(new_n556), .B(new_n558), .ZN(new_n559));
  NAND2_X1  g134(.A1(G78), .A2(G543), .ZN(new_n560));
  INV_X1    g135(.A(G65), .ZN(new_n561));
  OAI21_X1  g136(.A(new_n560), .B1(new_n539), .B2(new_n561), .ZN(new_n562));
  AOI22_X1  g137(.A1(G91), .A2(new_n529), .B1(new_n562), .B2(G651), .ZN(new_n563));
  NAND2_X1  g138(.A1(new_n559), .A2(new_n563), .ZN(G299));
  INV_X1    g139(.A(G168), .ZN(G286));
  INV_X1    g140(.A(G166), .ZN(G303));
  NAND2_X1  g141(.A1(new_n529), .A2(G87), .ZN(new_n567));
  OAI21_X1  g142(.A(G651), .B1(new_n514), .B2(G74), .ZN(new_n568));
  NAND2_X1  g143(.A1(new_n510), .A2(G49), .ZN(new_n569));
  NAND3_X1  g144(.A1(new_n567), .A2(new_n568), .A3(new_n569), .ZN(new_n570));
  INV_X1    g145(.A(KEYINPUT78), .ZN(new_n571));
  XNOR2_X1  g146(.A(new_n570), .B(new_n571), .ZN(new_n572));
  INV_X1    g147(.A(new_n572), .ZN(G288));
  AOI22_X1  g148(.A1(new_n529), .A2(G86), .B1(G48), .B2(new_n510), .ZN(new_n574));
  OAI21_X1  g149(.A(G61), .B1(new_n537), .B2(new_n538), .ZN(new_n575));
  NAND2_X1  g150(.A1(G73), .A2(G543), .ZN(new_n576));
  AOI21_X1  g151(.A(new_n518), .B1(new_n575), .B2(new_n576), .ZN(new_n577));
  INV_X1    g152(.A(KEYINPUT79), .ZN(new_n578));
  NOR2_X1   g153(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  AOI211_X1 g154(.A(KEYINPUT79), .B(new_n518), .C1(new_n575), .C2(new_n576), .ZN(new_n580));
  OAI21_X1  g155(.A(new_n574), .B1(new_n579), .B2(new_n580), .ZN(G305));
  AOI22_X1  g156(.A1(new_n529), .A2(G85), .B1(G47), .B2(new_n510), .ZN(new_n582));
  AOI22_X1  g157(.A1(new_n514), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n583));
  OAI21_X1  g158(.A(new_n582), .B1(new_n518), .B2(new_n583), .ZN(G290));
  AND3_X1   g159(.A1(new_n513), .A2(new_n514), .A3(G92), .ZN(new_n585));
  XNOR2_X1  g160(.A(new_n585), .B(KEYINPUT10), .ZN(new_n586));
  NAND2_X1  g161(.A1(G79), .A2(G543), .ZN(new_n587));
  INV_X1    g162(.A(G66), .ZN(new_n588));
  OAI21_X1  g163(.A(new_n587), .B1(new_n539), .B2(new_n588), .ZN(new_n589));
  AOI22_X1  g164(.A1(new_n589), .A2(G651), .B1(G54), .B2(new_n510), .ZN(new_n590));
  NAND2_X1  g165(.A1(new_n586), .A2(new_n590), .ZN(new_n591));
  INV_X1    g166(.A(G868), .ZN(new_n592));
  NAND2_X1  g167(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  OAI21_X1  g168(.A(new_n593), .B1(G171), .B2(new_n592), .ZN(G284));
  OAI21_X1  g169(.A(new_n593), .B1(G171), .B2(new_n592), .ZN(G321));
  NAND2_X1  g170(.A1(G299), .A2(new_n592), .ZN(new_n596));
  OAI21_X1  g171(.A(new_n596), .B1(new_n592), .B2(G168), .ZN(G297));
  OAI21_X1  g172(.A(new_n596), .B1(new_n592), .B2(G168), .ZN(G280));
  INV_X1    g173(.A(new_n591), .ZN(new_n599));
  INV_X1    g174(.A(G559), .ZN(new_n600));
  OAI21_X1  g175(.A(new_n599), .B1(new_n600), .B2(G860), .ZN(G148));
  NAND2_X1  g176(.A1(new_n599), .A2(new_n600), .ZN(new_n602));
  NAND2_X1  g177(.A1(new_n602), .A2(G868), .ZN(new_n603));
  OAI21_X1  g178(.A(new_n603), .B1(new_n550), .B2(G868), .ZN(new_n604));
  XOR2_X1   g179(.A(new_n604), .B(KEYINPUT80), .Z(G323));
  XNOR2_X1  g180(.A(G323), .B(KEYINPUT11), .ZN(G282));
  AND2_X1   g181(.A1(new_n476), .A2(new_n477), .ZN(new_n607));
  NAND2_X1  g182(.A1(new_n607), .A2(new_n463), .ZN(new_n608));
  XOR2_X1   g183(.A(KEYINPUT81), .B(KEYINPUT12), .Z(new_n609));
  XNOR2_X1  g184(.A(new_n608), .B(new_n609), .ZN(new_n610));
  XNOR2_X1  g185(.A(new_n610), .B(KEYINPUT13), .ZN(new_n611));
  OR2_X1    g186(.A1(new_n611), .A2(G2100), .ZN(new_n612));
  NAND2_X1  g187(.A1(new_n611), .A2(G2100), .ZN(new_n613));
  NAND2_X1  g188(.A1(new_n486), .A2(G135), .ZN(new_n614));
  NAND2_X1  g189(.A1(new_n488), .A2(G123), .ZN(new_n615));
  NOR2_X1   g190(.A1(new_n461), .A2(G111), .ZN(new_n616));
  OAI21_X1  g191(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n617));
  OAI211_X1 g192(.A(new_n614), .B(new_n615), .C1(new_n616), .C2(new_n617), .ZN(new_n618));
  XOR2_X1   g193(.A(new_n618), .B(G2096), .Z(new_n619));
  NAND3_X1  g194(.A1(new_n612), .A2(new_n613), .A3(new_n619), .ZN(G156));
  XOR2_X1   g195(.A(KEYINPUT15), .B(G2435), .Z(new_n621));
  XNOR2_X1  g196(.A(new_n621), .B(G2438), .ZN(new_n622));
  XOR2_X1   g197(.A(G2427), .B(G2430), .Z(new_n623));
  XNOR2_X1  g198(.A(new_n623), .B(KEYINPUT83), .ZN(new_n624));
  OR2_X1    g199(.A1(new_n622), .A2(new_n624), .ZN(new_n625));
  NAND2_X1  g200(.A1(new_n622), .A2(new_n624), .ZN(new_n626));
  NAND3_X1  g201(.A1(new_n625), .A2(KEYINPUT14), .A3(new_n626), .ZN(new_n627));
  XOR2_X1   g202(.A(KEYINPUT82), .B(KEYINPUT16), .Z(new_n628));
  XNOR2_X1  g203(.A(new_n627), .B(new_n628), .ZN(new_n629));
  XOR2_X1   g204(.A(G2451), .B(G2454), .Z(new_n630));
  XNOR2_X1  g205(.A(G2443), .B(G2446), .ZN(new_n631));
  XNOR2_X1  g206(.A(new_n630), .B(new_n631), .ZN(new_n632));
  XNOR2_X1  g207(.A(new_n629), .B(new_n632), .ZN(new_n633));
  XOR2_X1   g208(.A(G1341), .B(G1348), .Z(new_n634));
  NOR2_X1   g209(.A1(new_n633), .A2(new_n634), .ZN(new_n635));
  XNOR2_X1  g210(.A(new_n635), .B(KEYINPUT85), .ZN(new_n636));
  NAND2_X1  g211(.A1(new_n633), .A2(new_n634), .ZN(new_n637));
  XNOR2_X1  g212(.A(new_n637), .B(KEYINPUT84), .ZN(new_n638));
  INV_X1    g213(.A(G14), .ZN(new_n639));
  NOR3_X1   g214(.A1(new_n636), .A2(new_n638), .A3(new_n639), .ZN(G401));
  XOR2_X1   g215(.A(G2072), .B(G2078), .Z(new_n641));
  INV_X1    g216(.A(new_n641), .ZN(new_n642));
  XOR2_X1   g217(.A(G2084), .B(G2090), .Z(new_n643));
  XNOR2_X1  g218(.A(G2067), .B(G2678), .ZN(new_n644));
  NAND3_X1  g219(.A1(new_n642), .A2(new_n643), .A3(new_n644), .ZN(new_n645));
  XNOR2_X1  g220(.A(new_n645), .B(KEYINPUT18), .ZN(new_n646));
  XNOR2_X1  g221(.A(new_n641), .B(KEYINPUT17), .ZN(new_n647));
  XOR2_X1   g222(.A(new_n644), .B(KEYINPUT86), .Z(new_n648));
  AND2_X1   g223(.A1(new_n648), .A2(new_n643), .ZN(new_n649));
  AOI21_X1  g224(.A(new_n646), .B1(new_n647), .B2(new_n649), .ZN(new_n650));
  AOI21_X1  g225(.A(new_n643), .B1(new_n648), .B2(new_n641), .ZN(new_n651));
  NAND2_X1  g226(.A1(new_n651), .A2(KEYINPUT87), .ZN(new_n652));
  OAI21_X1  g227(.A(new_n652), .B1(new_n648), .B2(new_n647), .ZN(new_n653));
  NOR2_X1   g228(.A1(new_n651), .A2(KEYINPUT87), .ZN(new_n654));
  OAI21_X1  g229(.A(new_n650), .B1(new_n653), .B2(new_n654), .ZN(new_n655));
  XOR2_X1   g230(.A(G2096), .B(G2100), .Z(new_n656));
  XNOR2_X1  g231(.A(new_n655), .B(new_n656), .ZN(G227));
  XOR2_X1   g232(.A(G1971), .B(G1976), .Z(new_n658));
  XNOR2_X1  g233(.A(new_n658), .B(KEYINPUT19), .ZN(new_n659));
  XNOR2_X1  g234(.A(G1956), .B(G2474), .ZN(new_n660));
  XNOR2_X1  g235(.A(G1961), .B(G1966), .ZN(new_n661));
  NOR2_X1   g236(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  NAND2_X1  g237(.A1(new_n659), .A2(new_n662), .ZN(new_n663));
  XNOR2_X1  g238(.A(new_n663), .B(KEYINPUT20), .ZN(new_n664));
  AND2_X1   g239(.A1(new_n660), .A2(new_n661), .ZN(new_n665));
  NOR3_X1   g240(.A1(new_n659), .A2(new_n662), .A3(new_n665), .ZN(new_n666));
  AOI21_X1  g241(.A(new_n666), .B1(new_n659), .B2(new_n665), .ZN(new_n667));
  NAND2_X1  g242(.A1(new_n664), .A2(new_n667), .ZN(new_n668));
  XNOR2_X1  g243(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n669));
  XNOR2_X1  g244(.A(new_n668), .B(new_n669), .ZN(new_n670));
  XNOR2_X1  g245(.A(G1991), .B(G1996), .ZN(new_n671));
  XNOR2_X1  g246(.A(new_n670), .B(new_n671), .ZN(new_n672));
  XNOR2_X1  g247(.A(G1981), .B(G1986), .ZN(new_n673));
  XNOR2_X1  g248(.A(new_n672), .B(new_n673), .ZN(G229));
  INV_X1    g249(.A(G16), .ZN(new_n675));
  NAND2_X1  g250(.A1(new_n675), .A2(G20), .ZN(new_n676));
  XOR2_X1   g251(.A(new_n676), .B(KEYINPUT23), .Z(new_n677));
  AOI21_X1  g252(.A(new_n677), .B1(G299), .B2(G16), .ZN(new_n678));
  XNOR2_X1  g253(.A(new_n678), .B(KEYINPUT99), .ZN(new_n679));
  XOR2_X1   g254(.A(new_n679), .B(G1956), .Z(new_n680));
  NOR2_X1   g255(.A1(G29), .A2(G35), .ZN(new_n681));
  AOI21_X1  g256(.A(new_n681), .B1(G162), .B2(G29), .ZN(new_n682));
  XNOR2_X1  g257(.A(new_n682), .B(KEYINPUT29), .ZN(new_n683));
  OAI21_X1  g258(.A(new_n680), .B1(new_n683), .B2(G2090), .ZN(new_n684));
  NAND2_X1  g259(.A1(new_n683), .A2(G2090), .ZN(new_n685));
  NOR2_X1   g260(.A1(G29), .A2(G33), .ZN(new_n686));
  XOR2_X1   g261(.A(new_n686), .B(KEYINPUT96), .Z(new_n687));
  NAND3_X1  g262(.A1(new_n461), .A2(G103), .A3(G2104), .ZN(new_n688));
  XNOR2_X1  g263(.A(new_n688), .B(KEYINPUT25), .ZN(new_n689));
  NAND2_X1  g264(.A1(new_n607), .A2(G127), .ZN(new_n690));
  NAND2_X1  g265(.A1(G115), .A2(G2104), .ZN(new_n691));
  AOI21_X1  g266(.A(new_n461), .B1(new_n690), .B2(new_n691), .ZN(new_n692));
  INV_X1    g267(.A(G139), .ZN(new_n693));
  OAI21_X1  g268(.A(KEYINPUT97), .B1(new_n470), .B2(new_n693), .ZN(new_n694));
  OR3_X1    g269(.A1(new_n470), .A2(KEYINPUT97), .A3(new_n693), .ZN(new_n695));
  AOI211_X1 g270(.A(new_n689), .B(new_n692), .C1(new_n694), .C2(new_n695), .ZN(new_n696));
  AOI21_X1  g271(.A(new_n687), .B1(new_n696), .B2(G29), .ZN(new_n697));
  XNOR2_X1  g272(.A(new_n697), .B(KEYINPUT98), .ZN(new_n698));
  INV_X1    g273(.A(new_n698), .ZN(new_n699));
  OAI21_X1  g274(.A(new_n685), .B1(new_n699), .B2(G2072), .ZN(new_n700));
  NAND2_X1  g275(.A1(new_n675), .A2(G5), .ZN(new_n701));
  OAI21_X1  g276(.A(new_n701), .B1(G171), .B2(new_n675), .ZN(new_n702));
  INV_X1    g277(.A(G1961), .ZN(new_n703));
  XNOR2_X1  g278(.A(new_n702), .B(new_n703), .ZN(new_n704));
  NAND2_X1  g279(.A1(new_n463), .A2(G105), .ZN(new_n705));
  NAND2_X1  g280(.A1(new_n486), .A2(G141), .ZN(new_n706));
  NAND2_X1  g281(.A1(new_n488), .A2(G129), .ZN(new_n707));
  NAND3_X1  g282(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n708));
  XOR2_X1   g283(.A(new_n708), .B(KEYINPUT26), .Z(new_n709));
  AND4_X1   g284(.A1(new_n705), .A2(new_n706), .A3(new_n707), .A4(new_n709), .ZN(new_n710));
  INV_X1    g285(.A(G29), .ZN(new_n711));
  NOR2_X1   g286(.A1(new_n710), .A2(new_n711), .ZN(new_n712));
  AOI21_X1  g287(.A(new_n712), .B1(new_n711), .B2(G32), .ZN(new_n713));
  XNOR2_X1  g288(.A(KEYINPUT27), .B(G1996), .ZN(new_n714));
  OR2_X1    g289(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  XNOR2_X1  g290(.A(KEYINPUT30), .B(G28), .ZN(new_n716));
  OR2_X1    g291(.A1(KEYINPUT31), .A2(G11), .ZN(new_n717));
  NAND2_X1  g292(.A1(KEYINPUT31), .A2(G11), .ZN(new_n718));
  AOI22_X1  g293(.A1(new_n716), .A2(new_n711), .B1(new_n717), .B2(new_n718), .ZN(new_n719));
  OAI21_X1  g294(.A(new_n719), .B1(new_n618), .B2(new_n711), .ZN(new_n720));
  AOI21_X1  g295(.A(new_n720), .B1(new_n713), .B2(new_n714), .ZN(new_n721));
  NAND2_X1  g296(.A1(new_n675), .A2(G21), .ZN(new_n722));
  OAI21_X1  g297(.A(new_n722), .B1(G168), .B2(new_n675), .ZN(new_n723));
  INV_X1    g298(.A(G1966), .ZN(new_n724));
  XNOR2_X1  g299(.A(new_n723), .B(new_n724), .ZN(new_n725));
  NAND4_X1  g300(.A1(new_n704), .A2(new_n715), .A3(new_n721), .A4(new_n725), .ZN(new_n726));
  NOR2_X1   g301(.A1(G27), .A2(G29), .ZN(new_n727));
  AOI21_X1  g302(.A(new_n727), .B1(G164), .B2(G29), .ZN(new_n728));
  XNOR2_X1  g303(.A(new_n728), .B(G2078), .ZN(new_n729));
  NOR4_X1   g304(.A1(new_n684), .A2(new_n700), .A3(new_n726), .A4(new_n729), .ZN(new_n730));
  INV_X1    g305(.A(G160), .ZN(new_n731));
  INV_X1    g306(.A(KEYINPUT24), .ZN(new_n732));
  AND2_X1   g307(.A1(new_n732), .A2(G34), .ZN(new_n733));
  OAI21_X1  g308(.A(new_n711), .B1(new_n732), .B2(G34), .ZN(new_n734));
  OAI22_X1  g309(.A1(new_n731), .A2(new_n711), .B1(new_n733), .B2(new_n734), .ZN(new_n735));
  INV_X1    g310(.A(G2084), .ZN(new_n736));
  OR2_X1    g311(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  NAND2_X1  g312(.A1(new_n735), .A2(new_n736), .ZN(new_n738));
  NAND2_X1  g313(.A1(new_n699), .A2(G2072), .ZN(new_n739));
  NAND4_X1  g314(.A1(new_n730), .A2(new_n737), .A3(new_n738), .A4(new_n739), .ZN(new_n740));
  NAND2_X1  g315(.A1(new_n675), .A2(G19), .ZN(new_n741));
  OAI21_X1  g316(.A(new_n741), .B1(new_n550), .B2(new_n675), .ZN(new_n742));
  OR2_X1    g317(.A1(new_n742), .A2(G1341), .ZN(new_n743));
  NAND2_X1  g318(.A1(new_n742), .A2(G1341), .ZN(new_n744));
  NAND2_X1  g319(.A1(new_n675), .A2(G4), .ZN(new_n745));
  OAI21_X1  g320(.A(new_n745), .B1(new_n599), .B2(new_n675), .ZN(new_n746));
  INV_X1    g321(.A(G1348), .ZN(new_n747));
  XNOR2_X1  g322(.A(new_n746), .B(new_n747), .ZN(new_n748));
  NAND2_X1  g323(.A1(new_n711), .A2(G26), .ZN(new_n749));
  XOR2_X1   g324(.A(new_n749), .B(KEYINPUT28), .Z(new_n750));
  NAND2_X1  g325(.A1(new_n486), .A2(G140), .ZN(new_n751));
  NAND2_X1  g326(.A1(new_n488), .A2(G128), .ZN(new_n752));
  NOR2_X1   g327(.A1(new_n461), .A2(G116), .ZN(new_n753));
  OAI21_X1  g328(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n754));
  OAI211_X1 g329(.A(new_n751), .B(new_n752), .C1(new_n753), .C2(new_n754), .ZN(new_n755));
  AOI21_X1  g330(.A(new_n750), .B1(new_n755), .B2(G29), .ZN(new_n756));
  XNOR2_X1  g331(.A(new_n756), .B(G2067), .ZN(new_n757));
  NAND4_X1  g332(.A1(new_n743), .A2(new_n744), .A3(new_n748), .A4(new_n757), .ZN(new_n758));
  XOR2_X1   g333(.A(new_n758), .B(KEYINPUT95), .Z(new_n759));
  OR2_X1    g334(.A1(new_n740), .A2(new_n759), .ZN(new_n760));
  MUX2_X1   g335(.A(G6), .B(G305), .S(G16), .Z(new_n761));
  XOR2_X1   g336(.A(new_n761), .B(KEYINPUT89), .Z(new_n762));
  XNOR2_X1  g337(.A(KEYINPUT32), .B(G1981), .ZN(new_n763));
  OR2_X1    g338(.A1(new_n762), .A2(new_n763), .ZN(new_n764));
  NAND2_X1  g339(.A1(new_n762), .A2(new_n763), .ZN(new_n765));
  NOR2_X1   g340(.A1(G16), .A2(G22), .ZN(new_n766));
  AOI21_X1  g341(.A(new_n766), .B1(G166), .B2(G16), .ZN(new_n767));
  XNOR2_X1  g342(.A(KEYINPUT91), .B(G1971), .ZN(new_n768));
  XNOR2_X1  g343(.A(new_n767), .B(new_n768), .ZN(new_n769));
  INV_X1    g344(.A(KEYINPUT90), .ZN(new_n770));
  NAND2_X1  g345(.A1(new_n570), .A2(new_n770), .ZN(new_n771));
  NAND4_X1  g346(.A1(new_n567), .A2(KEYINPUT90), .A3(new_n568), .A4(new_n569), .ZN(new_n772));
  NAND2_X1  g347(.A1(new_n771), .A2(new_n772), .ZN(new_n773));
  MUX2_X1   g348(.A(G23), .B(new_n773), .S(G16), .Z(new_n774));
  XNOR2_X1  g349(.A(KEYINPUT33), .B(G1976), .ZN(new_n775));
  XNOR2_X1  g350(.A(new_n774), .B(new_n775), .ZN(new_n776));
  NAND4_X1  g351(.A1(new_n764), .A2(new_n765), .A3(new_n769), .A4(new_n776), .ZN(new_n777));
  NAND2_X1  g352(.A1(new_n777), .A2(KEYINPUT34), .ZN(new_n778));
  INV_X1    g353(.A(KEYINPUT93), .ZN(new_n779));
  XNOR2_X1  g354(.A(new_n778), .B(new_n779), .ZN(new_n780));
  NAND2_X1  g355(.A1(new_n486), .A2(G131), .ZN(new_n781));
  XNOR2_X1  g356(.A(new_n781), .B(KEYINPUT88), .ZN(new_n782));
  OAI21_X1  g357(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n783));
  INV_X1    g358(.A(G107), .ZN(new_n784));
  AOI21_X1  g359(.A(new_n783), .B1(new_n784), .B2(G2105), .ZN(new_n785));
  AOI21_X1  g360(.A(new_n785), .B1(new_n488), .B2(G119), .ZN(new_n786));
  NAND2_X1  g361(.A1(new_n782), .A2(new_n786), .ZN(new_n787));
  INV_X1    g362(.A(new_n787), .ZN(new_n788));
  NAND2_X1  g363(.A1(new_n788), .A2(G29), .ZN(new_n789));
  OAI21_X1  g364(.A(new_n789), .B1(G25), .B2(G29), .ZN(new_n790));
  XOR2_X1   g365(.A(KEYINPUT35), .B(G1991), .Z(new_n791));
  AND2_X1   g366(.A1(new_n790), .A2(new_n791), .ZN(new_n792));
  NOR2_X1   g367(.A1(new_n790), .A2(new_n791), .ZN(new_n793));
  MUX2_X1   g368(.A(G24), .B(G290), .S(G16), .Z(new_n794));
  XNOR2_X1  g369(.A(new_n794), .B(G1986), .ZN(new_n795));
  NOR3_X1   g370(.A1(new_n792), .A2(new_n793), .A3(new_n795), .ZN(new_n796));
  OAI21_X1  g371(.A(new_n796), .B1(new_n777), .B2(KEYINPUT34), .ZN(new_n797));
  NOR2_X1   g372(.A1(new_n797), .A2(KEYINPUT92), .ZN(new_n798));
  AND2_X1   g373(.A1(new_n797), .A2(KEYINPUT92), .ZN(new_n799));
  OAI21_X1  g374(.A(new_n780), .B1(new_n798), .B2(new_n799), .ZN(new_n800));
  INV_X1    g375(.A(KEYINPUT94), .ZN(new_n801));
  INV_X1    g376(.A(KEYINPUT36), .ZN(new_n802));
  NOR2_X1   g377(.A1(new_n801), .A2(new_n802), .ZN(new_n803));
  NAND2_X1  g378(.A1(new_n800), .A2(new_n803), .ZN(new_n804));
  OR2_X1    g379(.A1(new_n799), .A2(new_n798), .ZN(new_n805));
  INV_X1    g380(.A(new_n803), .ZN(new_n806));
  NAND3_X1  g381(.A1(new_n805), .A2(new_n806), .A3(new_n780), .ZN(new_n807));
  AOI21_X1  g382(.A(new_n760), .B1(new_n804), .B2(new_n807), .ZN(G311));
  NAND2_X1  g383(.A1(new_n807), .A2(new_n804), .ZN(new_n809));
  NOR2_X1   g384(.A1(new_n740), .A2(new_n759), .ZN(new_n810));
  NAND2_X1  g385(.A1(new_n809), .A2(new_n810), .ZN(G150));
  XNOR2_X1  g386(.A(KEYINPUT102), .B(G860), .ZN(new_n812));
  INV_X1    g387(.A(new_n812), .ZN(new_n813));
  AOI22_X1  g388(.A1(new_n514), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n814));
  NOR2_X1   g389(.A1(new_n814), .A2(new_n518), .ZN(new_n815));
  XOR2_X1   g390(.A(new_n815), .B(KEYINPUT100), .Z(new_n816));
  AOI22_X1  g391(.A1(new_n529), .A2(G93), .B1(G55), .B2(new_n510), .ZN(new_n817));
  XNOR2_X1  g392(.A(new_n817), .B(KEYINPUT101), .ZN(new_n818));
  NAND2_X1  g393(.A1(new_n816), .A2(new_n818), .ZN(new_n819));
  NAND2_X1  g394(.A1(new_n549), .A2(new_n819), .ZN(new_n820));
  OAI21_X1  g395(.A(new_n820), .B1(new_n548), .B2(new_n819), .ZN(new_n821));
  XOR2_X1   g396(.A(new_n821), .B(KEYINPUT38), .Z(new_n822));
  NOR2_X1   g397(.A1(new_n591), .A2(new_n600), .ZN(new_n823));
  XNOR2_X1  g398(.A(new_n822), .B(new_n823), .ZN(new_n824));
  INV_X1    g399(.A(KEYINPUT39), .ZN(new_n825));
  AOI21_X1  g400(.A(new_n813), .B1(new_n824), .B2(new_n825), .ZN(new_n826));
  OAI21_X1  g401(.A(new_n826), .B1(new_n825), .B2(new_n824), .ZN(new_n827));
  NAND2_X1  g402(.A1(new_n819), .A2(new_n813), .ZN(new_n828));
  XOR2_X1   g403(.A(new_n828), .B(KEYINPUT37), .Z(new_n829));
  NAND2_X1  g404(.A1(new_n827), .A2(new_n829), .ZN(G145));
  XOR2_X1   g405(.A(new_n710), .B(new_n755), .Z(new_n831));
  NAND2_X1  g406(.A1(new_n501), .A2(new_n502), .ZN(new_n832));
  NAND2_X1  g407(.A1(new_n503), .A2(KEYINPUT4), .ZN(new_n833));
  NAND3_X1  g408(.A1(new_n832), .A2(new_n505), .A3(new_n833), .ZN(new_n834));
  INV_X1    g409(.A(new_n498), .ZN(new_n835));
  NAND2_X1  g410(.A1(new_n834), .A2(new_n835), .ZN(new_n836));
  OR2_X1    g411(.A1(new_n831), .A2(new_n836), .ZN(new_n837));
  NAND2_X1  g412(.A1(new_n831), .A2(new_n836), .ZN(new_n838));
  OAI211_X1 g413(.A(new_n837), .B(new_n838), .C1(KEYINPUT104), .C2(new_n696), .ZN(new_n839));
  NAND2_X1  g414(.A1(new_n696), .A2(KEYINPUT104), .ZN(new_n840));
  XNOR2_X1  g415(.A(new_n839), .B(new_n840), .ZN(new_n841));
  NAND2_X1  g416(.A1(new_n488), .A2(G130), .ZN(new_n842));
  NOR2_X1   g417(.A1(new_n461), .A2(G118), .ZN(new_n843));
  OAI21_X1  g418(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n844));
  OAI21_X1  g419(.A(new_n842), .B1(new_n843), .B2(new_n844), .ZN(new_n845));
  AOI21_X1  g420(.A(new_n845), .B1(G142), .B2(new_n486), .ZN(new_n846));
  XOR2_X1   g421(.A(new_n846), .B(KEYINPUT105), .Z(new_n847));
  XNOR2_X1  g422(.A(new_n787), .B(new_n610), .ZN(new_n848));
  XOR2_X1   g423(.A(new_n847), .B(new_n848), .Z(new_n849));
  OR2_X1    g424(.A1(new_n841), .A2(new_n849), .ZN(new_n850));
  NAND2_X1  g425(.A1(new_n841), .A2(new_n849), .ZN(new_n851));
  NAND2_X1  g426(.A1(new_n850), .A2(new_n851), .ZN(new_n852));
  XNOR2_X1  g427(.A(G160), .B(KEYINPUT103), .ZN(new_n853));
  XNOR2_X1  g428(.A(new_n853), .B(G162), .ZN(new_n854));
  XNOR2_X1  g429(.A(new_n854), .B(new_n618), .ZN(new_n855));
  INV_X1    g430(.A(new_n855), .ZN(new_n856));
  NAND2_X1  g431(.A1(new_n852), .A2(new_n856), .ZN(new_n857));
  INV_X1    g432(.A(G37), .ZN(new_n858));
  NAND3_X1  g433(.A1(new_n850), .A2(new_n855), .A3(new_n851), .ZN(new_n859));
  NAND3_X1  g434(.A1(new_n857), .A2(new_n858), .A3(new_n859), .ZN(new_n860));
  XNOR2_X1  g435(.A(new_n860), .B(KEYINPUT40), .ZN(G395));
  NAND2_X1  g436(.A1(new_n819), .A2(new_n592), .ZN(new_n862));
  XNOR2_X1  g437(.A(new_n821), .B(new_n602), .ZN(new_n863));
  XNOR2_X1  g438(.A(new_n591), .B(G299), .ZN(new_n864));
  INV_X1    g439(.A(new_n864), .ZN(new_n865));
  NAND2_X1  g440(.A1(new_n863), .A2(new_n865), .ZN(new_n866));
  OR2_X1    g441(.A1(new_n866), .A2(KEYINPUT106), .ZN(new_n867));
  NAND2_X1  g442(.A1(new_n866), .A2(KEYINPUT106), .ZN(new_n868));
  INV_X1    g443(.A(KEYINPUT41), .ZN(new_n869));
  NAND2_X1  g444(.A1(new_n865), .A2(new_n869), .ZN(new_n870));
  INV_X1    g445(.A(KEYINPUT107), .ZN(new_n871));
  NAND2_X1  g446(.A1(new_n864), .A2(KEYINPUT41), .ZN(new_n872));
  NAND3_X1  g447(.A1(new_n870), .A2(new_n871), .A3(new_n872), .ZN(new_n873));
  NAND3_X1  g448(.A1(new_n865), .A2(KEYINPUT107), .A3(new_n869), .ZN(new_n874));
  NAND2_X1  g449(.A1(new_n873), .A2(new_n874), .ZN(new_n875));
  OR2_X1    g450(.A1(new_n863), .A2(new_n875), .ZN(new_n876));
  NAND3_X1  g451(.A1(new_n867), .A2(new_n868), .A3(new_n876), .ZN(new_n877));
  XNOR2_X1  g452(.A(new_n773), .B(G305), .ZN(new_n878));
  XNOR2_X1  g453(.A(G303), .B(G290), .ZN(new_n879));
  XNOR2_X1  g454(.A(new_n878), .B(new_n879), .ZN(new_n880));
  XNOR2_X1  g455(.A(new_n880), .B(KEYINPUT42), .ZN(new_n881));
  XNOR2_X1  g456(.A(new_n877), .B(new_n881), .ZN(new_n882));
  OAI21_X1  g457(.A(new_n862), .B1(new_n882), .B2(new_n592), .ZN(G295));
  OAI21_X1  g458(.A(new_n862), .B1(new_n882), .B2(new_n592), .ZN(G331));
  XNOR2_X1  g459(.A(G301), .B(G168), .ZN(new_n885));
  XNOR2_X1  g460(.A(new_n821), .B(new_n885), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n886), .A2(new_n865), .ZN(new_n887));
  OR2_X1    g462(.A1(new_n821), .A2(new_n885), .ZN(new_n888));
  NAND2_X1  g463(.A1(new_n821), .A2(new_n885), .ZN(new_n889));
  NAND4_X1  g464(.A1(new_n888), .A2(new_n874), .A3(new_n873), .A4(new_n889), .ZN(new_n890));
  NAND3_X1  g465(.A1(new_n887), .A2(new_n880), .A3(new_n890), .ZN(new_n891));
  INV_X1    g466(.A(KEYINPUT108), .ZN(new_n892));
  NAND2_X1  g467(.A1(new_n891), .A2(new_n892), .ZN(new_n893));
  NAND2_X1  g468(.A1(new_n887), .A2(new_n890), .ZN(new_n894));
  INV_X1    g469(.A(new_n880), .ZN(new_n895));
  NAND2_X1  g470(.A1(new_n894), .A2(new_n895), .ZN(new_n896));
  NAND4_X1  g471(.A1(new_n887), .A2(new_n890), .A3(KEYINPUT108), .A4(new_n880), .ZN(new_n897));
  NAND4_X1  g472(.A1(new_n893), .A2(new_n896), .A3(new_n858), .A4(new_n897), .ZN(new_n898));
  INV_X1    g473(.A(KEYINPUT43), .ZN(new_n899));
  AND2_X1   g474(.A1(new_n898), .A2(new_n899), .ZN(new_n900));
  AOI21_X1  g475(.A(G37), .B1(new_n891), .B2(new_n892), .ZN(new_n901));
  AOI21_X1  g476(.A(new_n886), .B1(new_n870), .B2(new_n872), .ZN(new_n902));
  INV_X1    g477(.A(new_n887), .ZN(new_n903));
  OAI21_X1  g478(.A(new_n895), .B1(new_n902), .B2(new_n903), .ZN(new_n904));
  AND4_X1   g479(.A1(KEYINPUT43), .A2(new_n901), .A3(new_n897), .A4(new_n904), .ZN(new_n905));
  OAI21_X1  g480(.A(KEYINPUT44), .B1(new_n900), .B2(new_n905), .ZN(new_n906));
  NAND2_X1  g481(.A1(new_n898), .A2(KEYINPUT43), .ZN(new_n907));
  NAND4_X1  g482(.A1(new_n901), .A2(new_n904), .A3(new_n899), .A4(new_n897), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n907), .A2(new_n908), .ZN(new_n909));
  INV_X1    g484(.A(KEYINPUT44), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n909), .A2(new_n910), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n906), .A2(new_n911), .ZN(G397));
  NOR2_X1   g487(.A1(KEYINPUT50), .A2(G1384), .ZN(new_n913));
  AOI21_X1  g488(.A(KEYINPUT112), .B1(new_n836), .B2(new_n913), .ZN(new_n914));
  INV_X1    g489(.A(KEYINPUT112), .ZN(new_n915));
  INV_X1    g490(.A(new_n913), .ZN(new_n916));
  AOI211_X1 g491(.A(new_n915), .B(new_n916), .C1(new_n834), .C2(new_n835), .ZN(new_n917));
  NOR2_X1   g492(.A1(new_n914), .A2(new_n917), .ZN(new_n918));
  INV_X1    g493(.A(KEYINPUT50), .ZN(new_n919));
  INV_X1    g494(.A(G1384), .ZN(new_n920));
  AOI21_X1  g495(.A(new_n919), .B1(new_n836), .B2(new_n920), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n483), .A2(G2105), .ZN(new_n922));
  INV_X1    g497(.A(new_n472), .ZN(new_n923));
  XNOR2_X1  g498(.A(KEYINPUT110), .B(G40), .ZN(new_n924));
  INV_X1    g499(.A(new_n924), .ZN(new_n925));
  NAND3_X1  g500(.A1(new_n922), .A2(new_n923), .A3(new_n925), .ZN(new_n926));
  NOR2_X1   g501(.A1(new_n921), .A2(new_n926), .ZN(new_n927));
  NAND3_X1  g502(.A1(new_n918), .A2(new_n927), .A3(new_n736), .ZN(new_n928));
  AOI21_X1  g503(.A(G1384), .B1(new_n834), .B2(new_n835), .ZN(new_n929));
  OAI211_X1 g504(.A(G160), .B(new_n925), .C1(new_n929), .C2(KEYINPUT45), .ZN(new_n930));
  XNOR2_X1  g505(.A(KEYINPUT109), .B(KEYINPUT45), .ZN(new_n931));
  NOR3_X1   g506(.A1(G164), .A2(G1384), .A3(new_n931), .ZN(new_n932));
  OAI21_X1  g507(.A(new_n724), .B1(new_n930), .B2(new_n932), .ZN(new_n933));
  NAND3_X1  g508(.A1(new_n928), .A2(G168), .A3(new_n933), .ZN(new_n934));
  NAND2_X1  g509(.A1(new_n934), .A2(G8), .ZN(new_n935));
  AOI21_X1  g510(.A(G168), .B1(new_n928), .B2(new_n933), .ZN(new_n936));
  OAI21_X1  g511(.A(KEYINPUT51), .B1(new_n935), .B2(new_n936), .ZN(new_n937));
  INV_X1    g512(.A(KEYINPUT51), .ZN(new_n938));
  NAND3_X1  g513(.A1(new_n934), .A2(new_n938), .A3(G8), .ZN(new_n939));
  NAND2_X1  g514(.A1(new_n937), .A2(new_n939), .ZN(new_n940));
  XOR2_X1   g515(.A(KEYINPUT121), .B(KEYINPUT54), .Z(new_n941));
  AOI21_X1  g516(.A(KEYINPUT45), .B1(new_n836), .B2(new_n920), .ZN(new_n942));
  NOR2_X1   g517(.A1(new_n942), .A2(new_n926), .ZN(new_n943));
  INV_X1    g518(.A(G2078), .ZN(new_n944));
  INV_X1    g519(.A(new_n931), .ZN(new_n945));
  NAND2_X1  g520(.A1(new_n929), .A2(new_n945), .ZN(new_n946));
  NAND4_X1  g521(.A1(new_n943), .A2(KEYINPUT122), .A3(new_n944), .A4(new_n946), .ZN(new_n947));
  INV_X1    g522(.A(KEYINPUT45), .ZN(new_n948));
  OAI21_X1  g523(.A(new_n948), .B1(G164), .B2(G1384), .ZN(new_n949));
  AOI211_X1 g524(.A(new_n472), .B(new_n924), .C1(new_n483), .C2(G2105), .ZN(new_n950));
  NAND4_X1  g525(.A1(new_n946), .A2(new_n949), .A3(new_n950), .A4(new_n944), .ZN(new_n951));
  INV_X1    g526(.A(KEYINPUT122), .ZN(new_n952));
  NAND2_X1  g527(.A1(new_n951), .A2(new_n952), .ZN(new_n953));
  NAND3_X1  g528(.A1(new_n947), .A2(new_n953), .A3(KEYINPUT53), .ZN(new_n954));
  NAND2_X1  g529(.A1(new_n836), .A2(new_n920), .ZN(new_n955));
  NAND2_X1  g530(.A1(new_n955), .A2(new_n931), .ZN(new_n956));
  NAND2_X1  g531(.A1(new_n929), .A2(KEYINPUT45), .ZN(new_n957));
  NAND4_X1  g532(.A1(new_n956), .A2(new_n944), .A3(new_n950), .A4(new_n957), .ZN(new_n958));
  INV_X1    g533(.A(KEYINPUT53), .ZN(new_n959));
  OAI21_X1  g534(.A(KEYINPUT50), .B1(G164), .B2(G1384), .ZN(new_n960));
  OAI21_X1  g535(.A(new_n915), .B1(G164), .B2(new_n916), .ZN(new_n961));
  NAND3_X1  g536(.A1(new_n836), .A2(KEYINPUT112), .A3(new_n913), .ZN(new_n962));
  NAND4_X1  g537(.A1(new_n960), .A2(new_n961), .A3(new_n950), .A4(new_n962), .ZN(new_n963));
  AOI22_X1  g538(.A1(new_n958), .A2(new_n959), .B1(new_n963), .B2(new_n703), .ZN(new_n964));
  AOI21_X1  g539(.A(G301), .B1(new_n954), .B2(new_n964), .ZN(new_n965));
  NAND2_X1  g540(.A1(new_n958), .A2(new_n959), .ZN(new_n966));
  NAND2_X1  g541(.A1(new_n963), .A2(new_n703), .ZN(new_n967));
  NOR2_X1   g542(.A1(new_n929), .A2(new_n945), .ZN(new_n968));
  NOR3_X1   g543(.A1(G164), .A2(new_n948), .A3(G1384), .ZN(new_n969));
  NOR2_X1   g544(.A1(new_n968), .A2(new_n969), .ZN(new_n970));
  AND3_X1   g545(.A1(new_n944), .A2(KEYINPUT53), .A3(G40), .ZN(new_n971));
  NAND3_X1  g546(.A1(new_n970), .A2(G160), .A3(new_n971), .ZN(new_n972));
  NAND3_X1  g547(.A1(new_n966), .A2(new_n967), .A3(new_n972), .ZN(new_n973));
  NOR2_X1   g548(.A1(new_n973), .A2(G171), .ZN(new_n974));
  OAI21_X1  g549(.A(new_n941), .B1(new_n965), .B2(new_n974), .ZN(new_n975));
  NAND3_X1  g550(.A1(new_n954), .A2(G301), .A3(new_n964), .ZN(new_n976));
  NAND2_X1  g551(.A1(new_n973), .A2(G171), .ZN(new_n977));
  NAND3_X1  g552(.A1(new_n976), .A2(new_n977), .A3(KEYINPUT54), .ZN(new_n978));
  AND3_X1   g553(.A1(new_n940), .A2(new_n975), .A3(new_n978), .ZN(new_n979));
  INV_X1    g554(.A(KEYINPUT123), .ZN(new_n980));
  NAND2_X1  g555(.A1(G303), .A2(G8), .ZN(new_n981));
  XNOR2_X1  g556(.A(new_n981), .B(KEYINPUT55), .ZN(new_n982));
  INV_X1    g557(.A(new_n982), .ZN(new_n983));
  AOI21_X1  g558(.A(G1971), .B1(new_n970), .B2(new_n950), .ZN(new_n984));
  NAND2_X1  g559(.A1(new_n961), .A2(new_n962), .ZN(new_n985));
  OAI211_X1 g560(.A(G160), .B(new_n925), .C1(new_n929), .C2(new_n919), .ZN(new_n986));
  NOR3_X1   g561(.A1(new_n985), .A2(new_n986), .A3(G2090), .ZN(new_n987));
  OAI211_X1 g562(.A(G8), .B(new_n983), .C1(new_n984), .C2(new_n987), .ZN(new_n988));
  NOR2_X1   g563(.A1(new_n926), .A2(new_n955), .ZN(new_n989));
  INV_X1    g564(.A(G8), .ZN(new_n990));
  NOR2_X1   g565(.A1(new_n989), .A2(new_n990), .ZN(new_n991));
  INV_X1    g566(.A(G1981), .ZN(new_n992));
  OAI211_X1 g567(.A(new_n574), .B(new_n992), .C1(new_n579), .C2(new_n580), .ZN(new_n993));
  NAND2_X1  g568(.A1(new_n510), .A2(G48), .ZN(new_n994));
  INV_X1    g569(.A(G86), .ZN(new_n995));
  OAI21_X1  g570(.A(new_n994), .B1(new_n995), .B2(new_n515), .ZN(new_n996));
  OAI21_X1  g571(.A(G1981), .B1(new_n996), .B2(new_n577), .ZN(new_n997));
  NAND3_X1  g572(.A1(new_n993), .A2(KEYINPUT49), .A3(new_n997), .ZN(new_n998));
  INV_X1    g573(.A(KEYINPUT115), .ZN(new_n999));
  XNOR2_X1  g574(.A(new_n998), .B(new_n999), .ZN(new_n1000));
  NAND2_X1  g575(.A1(new_n993), .A2(new_n997), .ZN(new_n1001));
  AOI21_X1  g576(.A(KEYINPUT49), .B1(new_n1001), .B2(KEYINPUT113), .ZN(new_n1002));
  INV_X1    g577(.A(KEYINPUT114), .ZN(new_n1003));
  INV_X1    g578(.A(KEYINPUT113), .ZN(new_n1004));
  NAND3_X1  g579(.A1(new_n993), .A2(new_n1004), .A3(new_n997), .ZN(new_n1005));
  AND3_X1   g580(.A1(new_n1002), .A2(new_n1003), .A3(new_n1005), .ZN(new_n1006));
  AOI21_X1  g581(.A(new_n1003), .B1(new_n1002), .B2(new_n1005), .ZN(new_n1007));
  OAI211_X1 g582(.A(new_n991), .B(new_n1000), .C1(new_n1006), .C2(new_n1007), .ZN(new_n1008));
  NAND3_X1  g583(.A1(new_n771), .A2(G1976), .A3(new_n772), .ZN(new_n1009));
  OAI211_X1 g584(.A(G8), .B(new_n1009), .C1(new_n926), .C2(new_n955), .ZN(new_n1010));
  NAND2_X1  g585(.A1(new_n1010), .A2(KEYINPUT52), .ZN(new_n1011));
  INV_X1    g586(.A(new_n1011), .ZN(new_n1012));
  INV_X1    g587(.A(KEYINPUT52), .ZN(new_n1013));
  OAI21_X1  g588(.A(new_n1013), .B1(new_n572), .B2(G1976), .ZN(new_n1014));
  NOR2_X1   g589(.A1(new_n1014), .A2(new_n1010), .ZN(new_n1015));
  NOR2_X1   g590(.A1(new_n1012), .A2(new_n1015), .ZN(new_n1016));
  NAND3_X1  g591(.A1(new_n988), .A2(new_n1008), .A3(new_n1016), .ZN(new_n1017));
  INV_X1    g592(.A(KEYINPUT116), .ZN(new_n1018));
  OAI21_X1  g593(.A(new_n1018), .B1(new_n921), .B2(new_n926), .ZN(new_n1019));
  NAND3_X1  g594(.A1(new_n960), .A2(new_n950), .A3(KEYINPUT116), .ZN(new_n1020));
  INV_X1    g595(.A(G2090), .ZN(new_n1021));
  NOR2_X1   g596(.A1(G164), .A2(new_n916), .ZN(new_n1022));
  INV_X1    g597(.A(new_n1022), .ZN(new_n1023));
  NAND4_X1  g598(.A1(new_n1019), .A2(new_n1020), .A3(new_n1021), .A4(new_n1023), .ZN(new_n1024));
  NAND3_X1  g599(.A1(new_n956), .A2(new_n950), .A3(new_n957), .ZN(new_n1025));
  INV_X1    g600(.A(G1971), .ZN(new_n1026));
  NAND2_X1  g601(.A1(new_n1025), .A2(new_n1026), .ZN(new_n1027));
  NAND2_X1  g602(.A1(new_n1024), .A2(new_n1027), .ZN(new_n1028));
  AOI21_X1  g603(.A(new_n983), .B1(new_n1028), .B2(G8), .ZN(new_n1029));
  OAI21_X1  g604(.A(new_n980), .B1(new_n1017), .B2(new_n1029), .ZN(new_n1030));
  NAND2_X1  g605(.A1(new_n1028), .A2(G8), .ZN(new_n1031));
  NAND2_X1  g606(.A1(new_n1031), .A2(new_n982), .ZN(new_n1032));
  OAI21_X1  g607(.A(new_n1011), .B1(new_n1010), .B2(new_n1014), .ZN(new_n1033));
  NAND2_X1  g608(.A1(new_n1002), .A2(new_n1005), .ZN(new_n1034));
  NAND2_X1  g609(.A1(new_n1034), .A2(KEYINPUT114), .ZN(new_n1035));
  NAND3_X1  g610(.A1(new_n1002), .A2(new_n1003), .A3(new_n1005), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n1035), .A2(new_n1036), .ZN(new_n1037));
  AND2_X1   g612(.A1(new_n1000), .A2(new_n991), .ZN(new_n1038));
  AOI21_X1  g613(.A(new_n1033), .B1(new_n1037), .B2(new_n1038), .ZN(new_n1039));
  NAND4_X1  g614(.A1(new_n1032), .A2(KEYINPUT123), .A3(new_n988), .A4(new_n1039), .ZN(new_n1040));
  AND2_X1   g615(.A1(new_n1030), .A2(new_n1040), .ZN(new_n1041));
  INV_X1    g616(.A(KEYINPUT124), .ZN(new_n1042));
  NAND3_X1  g617(.A1(new_n979), .A2(new_n1041), .A3(new_n1042), .ZN(new_n1043));
  NAND3_X1  g618(.A1(new_n940), .A2(new_n975), .A3(new_n978), .ZN(new_n1044));
  NAND2_X1  g619(.A1(new_n1030), .A2(new_n1040), .ZN(new_n1045));
  OAI21_X1  g620(.A(KEYINPUT124), .B1(new_n1044), .B2(new_n1045), .ZN(new_n1046));
  OR2_X1    g621(.A1(new_n559), .A2(KEYINPUT118), .ZN(new_n1047));
  NAND2_X1  g622(.A1(new_n559), .A2(KEYINPUT118), .ZN(new_n1048));
  NAND3_X1  g623(.A1(new_n1047), .A2(new_n1048), .A3(new_n563), .ZN(new_n1049));
  INV_X1    g624(.A(KEYINPUT57), .ZN(new_n1050));
  NAND2_X1  g625(.A1(new_n1049), .A2(new_n1050), .ZN(new_n1051));
  INV_X1    g626(.A(KEYINPUT119), .ZN(new_n1052));
  OAI21_X1  g627(.A(new_n1052), .B1(G299), .B2(new_n1050), .ZN(new_n1053));
  NAND4_X1  g628(.A1(new_n559), .A2(KEYINPUT119), .A3(KEYINPUT57), .A4(new_n563), .ZN(new_n1054));
  NAND2_X1  g629(.A1(new_n1053), .A2(new_n1054), .ZN(new_n1055));
  AND2_X1   g630(.A1(new_n1051), .A2(new_n1055), .ZN(new_n1056));
  XNOR2_X1  g631(.A(KEYINPUT117), .B(G1956), .ZN(new_n1057));
  INV_X1    g632(.A(new_n1057), .ZN(new_n1058));
  AOI21_X1  g633(.A(new_n1022), .B1(new_n986), .B2(new_n1018), .ZN(new_n1059));
  AOI21_X1  g634(.A(new_n1058), .B1(new_n1059), .B2(new_n1020), .ZN(new_n1060));
  XOR2_X1   g635(.A(KEYINPUT56), .B(G2072), .Z(new_n1061));
  NOR2_X1   g636(.A1(new_n1025), .A2(new_n1061), .ZN(new_n1062));
  OAI21_X1  g637(.A(new_n1056), .B1(new_n1060), .B2(new_n1062), .ZN(new_n1063));
  INV_X1    g638(.A(new_n1063), .ZN(new_n1064));
  NAND2_X1  g639(.A1(new_n963), .A2(new_n747), .ZN(new_n1065));
  INV_X1    g640(.A(G2067), .ZN(new_n1066));
  NAND2_X1  g641(.A1(new_n989), .A2(new_n1066), .ZN(new_n1067));
  NAND3_X1  g642(.A1(new_n1065), .A2(KEYINPUT120), .A3(new_n1067), .ZN(new_n1068));
  INV_X1    g643(.A(new_n1068), .ZN(new_n1069));
  AOI21_X1  g644(.A(KEYINPUT120), .B1(new_n1065), .B2(new_n1067), .ZN(new_n1070));
  NOR3_X1   g645(.A1(new_n1069), .A2(new_n591), .A3(new_n1070), .ZN(new_n1071));
  NAND2_X1  g646(.A1(new_n1059), .A2(new_n1020), .ZN(new_n1072));
  NAND2_X1  g647(.A1(new_n1072), .A2(new_n1057), .ZN(new_n1073));
  INV_X1    g648(.A(new_n1056), .ZN(new_n1074));
  INV_X1    g649(.A(new_n1062), .ZN(new_n1075));
  NAND3_X1  g650(.A1(new_n1073), .A2(new_n1074), .A3(new_n1075), .ZN(new_n1076));
  AOI21_X1  g651(.A(new_n1064), .B1(new_n1071), .B2(new_n1076), .ZN(new_n1077));
  OAI21_X1  g652(.A(KEYINPUT60), .B1(new_n1069), .B2(new_n1070), .ZN(new_n1078));
  INV_X1    g653(.A(new_n1070), .ZN(new_n1079));
  INV_X1    g654(.A(KEYINPUT60), .ZN(new_n1080));
  NAND3_X1  g655(.A1(new_n1079), .A2(new_n1080), .A3(new_n1068), .ZN(new_n1081));
  NAND3_X1  g656(.A1(new_n1078), .A2(new_n1081), .A3(new_n599), .ZN(new_n1082));
  NAND2_X1  g657(.A1(new_n1076), .A2(new_n1063), .ZN(new_n1083));
  INV_X1    g658(.A(KEYINPUT61), .ZN(new_n1084));
  NAND2_X1  g659(.A1(new_n1083), .A2(new_n1084), .ZN(new_n1085));
  NAND2_X1  g660(.A1(new_n1082), .A2(new_n1085), .ZN(new_n1086));
  XNOR2_X1  g661(.A(KEYINPUT58), .B(G1341), .ZN(new_n1087));
  OAI22_X1  g662(.A1(new_n1025), .A2(G1996), .B1(new_n989), .B2(new_n1087), .ZN(new_n1088));
  NAND2_X1  g663(.A1(new_n1088), .A2(new_n550), .ZN(new_n1089));
  XNOR2_X1  g664(.A(new_n1089), .B(KEYINPUT59), .ZN(new_n1090));
  NAND3_X1  g665(.A1(new_n1076), .A2(KEYINPUT61), .A3(new_n1063), .ZN(new_n1091));
  OAI211_X1 g666(.A(KEYINPUT60), .B(new_n591), .C1(new_n1069), .C2(new_n1070), .ZN(new_n1092));
  NAND3_X1  g667(.A1(new_n1090), .A2(new_n1091), .A3(new_n1092), .ZN(new_n1093));
  OAI21_X1  g668(.A(new_n1077), .B1(new_n1086), .B2(new_n1093), .ZN(new_n1094));
  NAND3_X1  g669(.A1(new_n1043), .A2(new_n1046), .A3(new_n1094), .ZN(new_n1095));
  INV_X1    g670(.A(new_n965), .ZN(new_n1096));
  AND3_X1   g671(.A1(new_n934), .A2(new_n938), .A3(G8), .ZN(new_n1097));
  NOR2_X1   g672(.A1(new_n963), .A2(G2084), .ZN(new_n1098));
  AOI21_X1  g673(.A(G1966), .B1(new_n943), .B2(new_n946), .ZN(new_n1099));
  OAI21_X1  g674(.A(G286), .B1(new_n1098), .B2(new_n1099), .ZN(new_n1100));
  NAND3_X1  g675(.A1(new_n1100), .A2(G8), .A3(new_n934), .ZN(new_n1101));
  AOI21_X1  g676(.A(new_n1097), .B1(KEYINPUT51), .B2(new_n1101), .ZN(new_n1102));
  INV_X1    g677(.A(KEYINPUT62), .ZN(new_n1103));
  AOI21_X1  g678(.A(new_n1096), .B1(new_n1102), .B2(new_n1103), .ZN(new_n1104));
  NAND3_X1  g679(.A1(new_n1041), .A2(new_n1104), .A3(KEYINPUT125), .ZN(new_n1105));
  NAND3_X1  g680(.A1(new_n937), .A2(new_n1103), .A3(new_n939), .ZN(new_n1106));
  NAND4_X1  g681(.A1(new_n1106), .A2(new_n1030), .A3(new_n1040), .A4(new_n965), .ZN(new_n1107));
  INV_X1    g682(.A(KEYINPUT125), .ZN(new_n1108));
  NAND2_X1  g683(.A1(new_n1107), .A2(new_n1108), .ZN(new_n1109));
  NAND2_X1  g684(.A1(new_n940), .A2(KEYINPUT62), .ZN(new_n1110));
  NAND3_X1  g685(.A1(new_n1105), .A2(new_n1109), .A3(new_n1110), .ZN(new_n1111));
  INV_X1    g686(.A(new_n1008), .ZN(new_n1112));
  NOR3_X1   g687(.A1(new_n1112), .A2(new_n988), .A3(new_n1033), .ZN(new_n1113));
  OR2_X1    g688(.A1(G288), .A2(G1976), .ZN(new_n1114));
  OAI21_X1  g689(.A(new_n993), .B1(new_n1112), .B2(new_n1114), .ZN(new_n1115));
  AOI21_X1  g690(.A(new_n1113), .B1(new_n991), .B2(new_n1115), .ZN(new_n1116));
  NOR2_X1   g691(.A1(new_n1017), .A2(new_n1029), .ZN(new_n1117));
  INV_X1    g692(.A(KEYINPUT63), .ZN(new_n1118));
  AOI211_X1 g693(.A(new_n990), .B(G286), .C1(new_n928), .C2(new_n933), .ZN(new_n1119));
  NAND3_X1  g694(.A1(new_n1117), .A2(new_n1118), .A3(new_n1119), .ZN(new_n1120));
  NAND2_X1  g695(.A1(new_n1039), .A2(new_n1119), .ZN(new_n1121));
  OAI21_X1  g696(.A(new_n1027), .B1(G2090), .B2(new_n963), .ZN(new_n1122));
  AOI21_X1  g697(.A(new_n983), .B1(new_n1122), .B2(G8), .ZN(new_n1123));
  OAI21_X1  g698(.A(KEYINPUT63), .B1(new_n1121), .B2(new_n1123), .ZN(new_n1124));
  AND3_X1   g699(.A1(new_n1116), .A2(new_n1120), .A3(new_n1124), .ZN(new_n1125));
  NAND3_X1  g700(.A1(new_n1095), .A2(new_n1111), .A3(new_n1125), .ZN(new_n1126));
  NOR2_X1   g701(.A1(new_n956), .A2(new_n926), .ZN(new_n1127));
  XNOR2_X1  g702(.A(new_n1127), .B(KEYINPUT111), .ZN(new_n1128));
  OR2_X1    g703(.A1(new_n788), .A2(new_n791), .ZN(new_n1129));
  XNOR2_X1  g704(.A(new_n755), .B(new_n1066), .ZN(new_n1130));
  XNOR2_X1  g705(.A(new_n710), .B(G1996), .ZN(new_n1131));
  NAND2_X1  g706(.A1(new_n788), .A2(new_n791), .ZN(new_n1132));
  NAND4_X1  g707(.A1(new_n1129), .A2(new_n1130), .A3(new_n1131), .A4(new_n1132), .ZN(new_n1133));
  XNOR2_X1  g708(.A(G290), .B(G1986), .ZN(new_n1134));
  OAI21_X1  g709(.A(new_n1128), .B1(new_n1133), .B2(new_n1134), .ZN(new_n1135));
  NAND2_X1  g710(.A1(new_n1126), .A2(new_n1135), .ZN(new_n1136));
  NAND2_X1  g711(.A1(new_n1131), .A2(new_n1130), .ZN(new_n1137));
  OAI22_X1  g712(.A1(new_n1137), .A2(new_n1132), .B1(G2067), .B2(new_n755), .ZN(new_n1138));
  NAND2_X1  g713(.A1(new_n1128), .A2(new_n1138), .ZN(new_n1139));
  NOR2_X1   g714(.A1(G290), .A2(G1986), .ZN(new_n1140));
  NAND3_X1  g715(.A1(new_n1128), .A2(KEYINPUT48), .A3(new_n1140), .ZN(new_n1141));
  NAND2_X1  g716(.A1(new_n1128), .A2(new_n1133), .ZN(new_n1142));
  NAND2_X1  g717(.A1(new_n1141), .A2(new_n1142), .ZN(new_n1143));
  AOI21_X1  g718(.A(KEYINPUT48), .B1(new_n1128), .B2(new_n1140), .ZN(new_n1144));
  OAI21_X1  g719(.A(new_n1139), .B1(new_n1143), .B2(new_n1144), .ZN(new_n1145));
  INV_X1    g720(.A(G1996), .ZN(new_n1146));
  NAND3_X1  g721(.A1(new_n1128), .A2(KEYINPUT46), .A3(new_n1146), .ZN(new_n1147));
  XOR2_X1   g722(.A(new_n1147), .B(KEYINPUT126), .Z(new_n1148));
  NAND2_X1  g723(.A1(new_n1130), .A2(new_n710), .ZN(new_n1149));
  NAND2_X1  g724(.A1(new_n1128), .A2(new_n1149), .ZN(new_n1150));
  XNOR2_X1  g725(.A(new_n1150), .B(KEYINPUT127), .ZN(new_n1151));
  AND2_X1   g726(.A1(new_n1128), .A2(new_n1146), .ZN(new_n1152));
  OAI211_X1 g727(.A(new_n1148), .B(new_n1151), .C1(KEYINPUT46), .C2(new_n1152), .ZN(new_n1153));
  OR2_X1    g728(.A1(new_n1153), .A2(KEYINPUT47), .ZN(new_n1154));
  NAND2_X1  g729(.A1(new_n1153), .A2(KEYINPUT47), .ZN(new_n1155));
  AOI21_X1  g730(.A(new_n1145), .B1(new_n1154), .B2(new_n1155), .ZN(new_n1156));
  NAND2_X1  g731(.A1(new_n1136), .A2(new_n1156), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g732(.A(G319), .ZN(new_n1159));
  NOR4_X1   g733(.A1(G401), .A2(new_n1159), .A3(G227), .A4(G229), .ZN(new_n1160));
  NAND3_X1  g734(.A1(new_n909), .A2(new_n1160), .A3(new_n860), .ZN(G225));
  INV_X1    g735(.A(G225), .ZN(G308));
endmodule


