//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 1 1 0 1 1 0 0 0 0 1 0 1 0 0 1 0 1 1 1 0 1 0 1 1 0 0 0 0 0 0 1 1 0 0 0 0 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 0 0 0 1 0 1 0 1 0 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:32:25 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n454, new_n458,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n497, new_n498, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n513, new_n514, new_n515, new_n516, new_n517, new_n518,
    new_n519, new_n520, new_n521, new_n522, new_n523, new_n524, new_n525,
    new_n526, new_n527, new_n528, new_n531, new_n532, new_n533, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n548, new_n549, new_n551, new_n552,
    new_n554, new_n555, new_n556, new_n557, new_n558, new_n559, new_n560,
    new_n561, new_n562, new_n563, new_n564, new_n567, new_n568, new_n570,
    new_n571, new_n572, new_n573, new_n574, new_n575, new_n576, new_n577,
    new_n578, new_n579, new_n580, new_n581, new_n582, new_n583, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n603, new_n606, new_n607, new_n609, new_n610, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n828, new_n829,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1215, new_n1216, new_n1217, new_n1218, new_n1219, new_n1220,
    new_n1221, new_n1223, new_n1224, new_n1225;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  XNOR2_X1  g005(.A(KEYINPUT64), .B(G2066), .ZN(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  XOR2_X1   g008(.A(KEYINPUT65), .B(G44), .Z(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  XOR2_X1   g011(.A(KEYINPUT66), .B(G96), .Z(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G218), .A2(G221), .A3(G219), .A4(G220), .ZN(new_n450));
  XOR2_X1   g025(.A(new_n450), .B(KEYINPUT2), .Z(new_n451));
  NAND4_X1  g026(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n452));
  XNOR2_X1  g027(.A(new_n452), .B(KEYINPUT67), .ZN(new_n453));
  OR2_X1    g028(.A1(new_n451), .A2(new_n453), .ZN(new_n454));
  XOR2_X1   g029(.A(new_n454), .B(KEYINPUT68), .Z(G261));
  INV_X1    g030(.A(G261), .ZN(G325));
  AOI22_X1  g031(.A1(new_n451), .A2(G2106), .B1(G567), .B2(new_n453), .ZN(G319));
  NAND2_X1  g032(.A1(G113), .A2(G2104), .ZN(new_n458));
  AND2_X1   g033(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n459));
  NOR2_X1   g034(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n460));
  NOR2_X1   g035(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  INV_X1    g036(.A(G125), .ZN(new_n462));
  OAI21_X1  g037(.A(new_n458), .B1(new_n461), .B2(new_n462), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n463), .A2(G2105), .ZN(new_n464));
  OR2_X1    g039(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n465));
  NAND2_X1  g040(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n466));
  AOI21_X1  g041(.A(G2105), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  INV_X1    g042(.A(G2104), .ZN(new_n468));
  NOR2_X1   g043(.A1(new_n468), .A2(G2105), .ZN(new_n469));
  AOI22_X1  g044(.A1(new_n467), .A2(G137), .B1(G101), .B2(new_n469), .ZN(new_n470));
  AND2_X1   g045(.A1(new_n464), .A2(new_n470), .ZN(G160));
  OR2_X1    g046(.A1(G100), .A2(G2105), .ZN(new_n472));
  INV_X1    g047(.A(KEYINPUT69), .ZN(new_n473));
  AOI21_X1  g048(.A(new_n468), .B1(new_n472), .B2(new_n473), .ZN(new_n474));
  INV_X1    g049(.A(G2105), .ZN(new_n475));
  OAI221_X1 g050(.A(new_n474), .B1(new_n473), .B2(new_n472), .C1(G112), .C2(new_n475), .ZN(new_n476));
  NOR2_X1   g051(.A1(new_n461), .A2(new_n475), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n477), .A2(G124), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n467), .A2(G136), .ZN(new_n479));
  NAND3_X1  g054(.A1(new_n476), .A2(new_n478), .A3(new_n479), .ZN(new_n480));
  INV_X1    g055(.A(new_n480), .ZN(G162));
  INV_X1    g056(.A(KEYINPUT70), .ZN(new_n482));
  OAI21_X1  g057(.A(new_n482), .B1(new_n475), .B2(G114), .ZN(new_n483));
  INV_X1    g058(.A(G114), .ZN(new_n484));
  NAND3_X1  g059(.A1(new_n484), .A2(KEYINPUT70), .A3(G2105), .ZN(new_n485));
  INV_X1    g060(.A(G102), .ZN(new_n486));
  NAND2_X1  g061(.A1(new_n486), .A2(new_n475), .ZN(new_n487));
  NAND4_X1  g062(.A1(new_n483), .A2(new_n485), .A3(G2104), .A4(new_n487), .ZN(new_n488));
  OAI211_X1 g063(.A(G126), .B(G2105), .C1(new_n459), .C2(new_n460), .ZN(new_n489));
  NAND2_X1  g064(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  OAI211_X1 g065(.A(G138), .B(new_n475), .C1(new_n459), .C2(new_n460), .ZN(new_n491));
  NAND2_X1  g066(.A1(new_n491), .A2(KEYINPUT4), .ZN(new_n492));
  XNOR2_X1  g067(.A(KEYINPUT3), .B(G2104), .ZN(new_n493));
  INV_X1    g068(.A(KEYINPUT4), .ZN(new_n494));
  NAND4_X1  g069(.A1(new_n493), .A2(new_n494), .A3(G138), .A4(new_n475), .ZN(new_n495));
  AOI21_X1  g070(.A(new_n490), .B1(new_n492), .B2(new_n495), .ZN(G164));
  INV_X1    g071(.A(KEYINPUT5), .ZN(new_n497));
  INV_X1    g072(.A(G543), .ZN(new_n498));
  OAI21_X1  g073(.A(new_n497), .B1(new_n498), .B2(KEYINPUT71), .ZN(new_n499));
  INV_X1    g074(.A(KEYINPUT71), .ZN(new_n500));
  NAND3_X1  g075(.A1(new_n500), .A2(KEYINPUT5), .A3(G543), .ZN(new_n501));
  NAND2_X1  g076(.A1(new_n499), .A2(new_n501), .ZN(new_n502));
  AOI22_X1  g077(.A1(new_n502), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n503));
  INV_X1    g078(.A(G651), .ZN(new_n504));
  NOR2_X1   g079(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  XNOR2_X1  g080(.A(KEYINPUT6), .B(G651), .ZN(new_n506));
  NAND2_X1  g081(.A1(new_n502), .A2(new_n506), .ZN(new_n507));
  INV_X1    g082(.A(G88), .ZN(new_n508));
  NAND2_X1  g083(.A1(new_n506), .A2(G543), .ZN(new_n509));
  INV_X1    g084(.A(G50), .ZN(new_n510));
  OAI22_X1  g085(.A1(new_n507), .A2(new_n508), .B1(new_n509), .B2(new_n510), .ZN(new_n511));
  NOR2_X1   g086(.A1(new_n505), .A2(new_n511), .ZN(G166));
  INV_X1    g087(.A(KEYINPUT72), .ZN(new_n513));
  NAND2_X1  g088(.A1(new_n502), .A2(new_n513), .ZN(new_n514));
  NAND3_X1  g089(.A1(new_n499), .A2(KEYINPUT72), .A3(new_n501), .ZN(new_n515));
  NAND2_X1  g090(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  NAND3_X1  g091(.A1(new_n516), .A2(G63), .A3(G651), .ZN(new_n517));
  INV_X1    g092(.A(new_n509), .ZN(new_n518));
  NAND2_X1  g093(.A1(new_n518), .A2(G51), .ZN(new_n519));
  OR2_X1    g094(.A1(KEYINPUT73), .A2(G89), .ZN(new_n520));
  NAND2_X1  g095(.A1(KEYINPUT73), .A2(G89), .ZN(new_n521));
  NAND4_X1  g096(.A1(new_n502), .A2(new_n506), .A3(new_n520), .A4(new_n521), .ZN(new_n522));
  INV_X1    g097(.A(KEYINPUT74), .ZN(new_n523));
  NAND3_X1  g098(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n524));
  XNOR2_X1  g099(.A(new_n524), .B(KEYINPUT7), .ZN(new_n525));
  NAND3_X1  g100(.A1(new_n522), .A2(new_n523), .A3(new_n525), .ZN(new_n526));
  INV_X1    g101(.A(new_n526), .ZN(new_n527));
  AOI21_X1  g102(.A(new_n523), .B1(new_n522), .B2(new_n525), .ZN(new_n528));
  OAI211_X1 g103(.A(new_n517), .B(new_n519), .C1(new_n527), .C2(new_n528), .ZN(G286));
  INV_X1    g104(.A(G286), .ZN(G168));
  INV_X1    g105(.A(new_n507), .ZN(new_n531));
  AOI22_X1  g106(.A1(new_n531), .A2(G90), .B1(new_n518), .B2(G52), .ZN(new_n532));
  AOI22_X1  g107(.A1(new_n516), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n533));
  OAI21_X1  g108(.A(new_n532), .B1(new_n533), .B2(new_n504), .ZN(G301));
  INV_X1    g109(.A(G301), .ZN(G171));
  INV_X1    g110(.A(G56), .ZN(new_n536));
  AOI21_X1  g111(.A(new_n536), .B1(new_n514), .B2(new_n515), .ZN(new_n537));
  AND2_X1   g112(.A1(G68), .A2(G543), .ZN(new_n538));
  OAI21_X1  g113(.A(G651), .B1(new_n537), .B2(new_n538), .ZN(new_n539));
  NAND2_X1  g114(.A1(new_n539), .A2(KEYINPUT75), .ZN(new_n540));
  INV_X1    g115(.A(KEYINPUT75), .ZN(new_n541));
  OAI211_X1 g116(.A(new_n541), .B(G651), .C1(new_n537), .C2(new_n538), .ZN(new_n542));
  NAND2_X1  g117(.A1(new_n540), .A2(new_n542), .ZN(new_n543));
  NAND2_X1  g118(.A1(new_n531), .A2(G81), .ZN(new_n544));
  NAND2_X1  g119(.A1(new_n518), .A2(G43), .ZN(new_n545));
  AND3_X1   g120(.A1(new_n543), .A2(new_n544), .A3(new_n545), .ZN(new_n546));
  NAND2_X1  g121(.A1(new_n546), .A2(G860), .ZN(G153));
  AND3_X1   g122(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n548));
  NAND2_X1  g123(.A1(new_n548), .A2(G36), .ZN(new_n549));
  XOR2_X1   g124(.A(new_n549), .B(KEYINPUT76), .Z(G176));
  NAND2_X1  g125(.A1(G1), .A2(G3), .ZN(new_n551));
  XNOR2_X1  g126(.A(new_n551), .B(KEYINPUT8), .ZN(new_n552));
  NAND2_X1  g127(.A1(new_n548), .A2(new_n552), .ZN(G188));
  INV_X1    g128(.A(G65), .ZN(new_n554));
  AOI21_X1  g129(.A(new_n554), .B1(new_n499), .B2(new_n501), .ZN(new_n555));
  AND2_X1   g130(.A1(G78), .A2(G543), .ZN(new_n556));
  OAI21_X1  g131(.A(G651), .B1(new_n555), .B2(new_n556), .ZN(new_n557));
  NAND2_X1  g132(.A1(new_n557), .A2(KEYINPUT77), .ZN(new_n558));
  INV_X1    g133(.A(KEYINPUT77), .ZN(new_n559));
  OAI211_X1 g134(.A(new_n559), .B(G651), .C1(new_n555), .C2(new_n556), .ZN(new_n560));
  NAND2_X1  g135(.A1(new_n558), .A2(new_n560), .ZN(new_n561));
  NAND2_X1  g136(.A1(new_n531), .A2(G91), .ZN(new_n562));
  NAND3_X1  g137(.A1(new_n506), .A2(G53), .A3(G543), .ZN(new_n563));
  XNOR2_X1  g138(.A(new_n563), .B(KEYINPUT9), .ZN(new_n564));
  NAND3_X1  g139(.A1(new_n561), .A2(new_n562), .A3(new_n564), .ZN(G299));
  INV_X1    g140(.A(G166), .ZN(G303));
  OAI21_X1  g141(.A(G651), .B1(new_n516), .B2(G74), .ZN(new_n567));
  AOI22_X1  g142(.A1(new_n531), .A2(G87), .B1(new_n518), .B2(G49), .ZN(new_n568));
  NAND2_X1  g143(.A1(new_n567), .A2(new_n568), .ZN(G288));
  NAND2_X1  g144(.A1(new_n518), .A2(G48), .ZN(new_n570));
  AND3_X1   g145(.A1(new_n502), .A2(G86), .A3(new_n506), .ZN(new_n571));
  INV_X1    g146(.A(new_n571), .ZN(new_n572));
  AND3_X1   g147(.A1(new_n500), .A2(KEYINPUT5), .A3(G543), .ZN(new_n573));
  AOI21_X1  g148(.A(KEYINPUT5), .B1(new_n500), .B2(G543), .ZN(new_n574));
  OAI21_X1  g149(.A(G61), .B1(new_n573), .B2(new_n574), .ZN(new_n575));
  NAND2_X1  g150(.A1(G73), .A2(G543), .ZN(new_n576));
  NAND2_X1  g151(.A1(new_n575), .A2(new_n576), .ZN(new_n577));
  AOI21_X1  g152(.A(KEYINPUT78), .B1(new_n577), .B2(G651), .ZN(new_n578));
  INV_X1    g153(.A(G61), .ZN(new_n579));
  AOI21_X1  g154(.A(new_n579), .B1(new_n499), .B2(new_n501), .ZN(new_n580));
  INV_X1    g155(.A(new_n576), .ZN(new_n581));
  OAI211_X1 g156(.A(KEYINPUT78), .B(G651), .C1(new_n580), .C2(new_n581), .ZN(new_n582));
  INV_X1    g157(.A(new_n582), .ZN(new_n583));
  OAI211_X1 g158(.A(new_n570), .B(new_n572), .C1(new_n578), .C2(new_n583), .ZN(G305));
  AOI22_X1  g159(.A1(new_n516), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n585));
  NOR2_X1   g160(.A1(new_n585), .A2(new_n504), .ZN(new_n586));
  INV_X1    g161(.A(G85), .ZN(new_n587));
  INV_X1    g162(.A(G47), .ZN(new_n588));
  OAI22_X1  g163(.A1(new_n507), .A2(new_n587), .B1(new_n509), .B2(new_n588), .ZN(new_n589));
  NOR2_X1   g164(.A1(new_n586), .A2(new_n589), .ZN(new_n590));
  INV_X1    g165(.A(new_n590), .ZN(G290));
  NAND3_X1  g166(.A1(new_n502), .A2(G92), .A3(new_n506), .ZN(new_n592));
  INV_X1    g167(.A(KEYINPUT10), .ZN(new_n593));
  XNOR2_X1  g168(.A(new_n592), .B(new_n593), .ZN(new_n594));
  NAND2_X1  g169(.A1(new_n518), .A2(G54), .ZN(new_n595));
  AOI22_X1  g170(.A1(new_n502), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n596));
  OR2_X1    g171(.A1(new_n596), .A2(new_n504), .ZN(new_n597));
  NAND3_X1  g172(.A1(new_n594), .A2(new_n595), .A3(new_n597), .ZN(new_n598));
  INV_X1    g173(.A(G868), .ZN(new_n599));
  NAND2_X1  g174(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  OAI21_X1  g175(.A(new_n600), .B1(G171), .B2(new_n599), .ZN(G284));
  OAI21_X1  g176(.A(new_n600), .B1(G171), .B2(new_n599), .ZN(G321));
  NAND2_X1  g177(.A1(G299), .A2(new_n599), .ZN(new_n603));
  OAI21_X1  g178(.A(new_n603), .B1(G168), .B2(new_n599), .ZN(G297));
  XOR2_X1   g179(.A(G297), .B(KEYINPUT79), .Z(G280));
  INV_X1    g180(.A(new_n598), .ZN(new_n606));
  INV_X1    g181(.A(G559), .ZN(new_n607));
  OAI21_X1  g182(.A(new_n606), .B1(new_n607), .B2(G860), .ZN(G148));
  NAND2_X1  g183(.A1(new_n606), .A2(new_n607), .ZN(new_n609));
  NAND2_X1  g184(.A1(new_n609), .A2(G868), .ZN(new_n610));
  OAI21_X1  g185(.A(new_n610), .B1(new_n546), .B2(G868), .ZN(G323));
  XNOR2_X1  g186(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g187(.A1(new_n493), .A2(new_n469), .ZN(new_n613));
  XNOR2_X1  g188(.A(new_n613), .B(KEYINPUT12), .ZN(new_n614));
  XNOR2_X1  g189(.A(new_n614), .B(KEYINPUT13), .ZN(new_n615));
  XNOR2_X1  g190(.A(new_n615), .B(G2100), .ZN(new_n616));
  NAND2_X1  g191(.A1(new_n477), .A2(G123), .ZN(new_n617));
  NAND2_X1  g192(.A1(new_n467), .A2(G135), .ZN(new_n618));
  NOR2_X1   g193(.A1(G99), .A2(G2105), .ZN(new_n619));
  OAI21_X1  g194(.A(G2104), .B1(new_n475), .B2(G111), .ZN(new_n620));
  OAI211_X1 g195(.A(new_n617), .B(new_n618), .C1(new_n619), .C2(new_n620), .ZN(new_n621));
  INV_X1    g196(.A(G2096), .ZN(new_n622));
  XNOR2_X1  g197(.A(new_n621), .B(new_n622), .ZN(new_n623));
  NAND2_X1  g198(.A1(new_n616), .A2(new_n623), .ZN(G156));
  XNOR2_X1  g199(.A(G2451), .B(G2454), .ZN(new_n625));
  XNOR2_X1  g200(.A(new_n625), .B(KEYINPUT16), .ZN(new_n626));
  XNOR2_X1  g201(.A(G2443), .B(G2446), .ZN(new_n627));
  XNOR2_X1  g202(.A(new_n626), .B(new_n627), .ZN(new_n628));
  XNOR2_X1  g203(.A(G1341), .B(G1348), .ZN(new_n629));
  INV_X1    g204(.A(new_n629), .ZN(new_n630));
  XNOR2_X1  g205(.A(new_n628), .B(new_n630), .ZN(new_n631));
  XNOR2_X1  g206(.A(KEYINPUT15), .B(G2430), .ZN(new_n632));
  XNOR2_X1  g207(.A(new_n632), .B(G2435), .ZN(new_n633));
  XOR2_X1   g208(.A(G2427), .B(G2438), .Z(new_n634));
  XNOR2_X1  g209(.A(new_n633), .B(new_n634), .ZN(new_n635));
  NAND2_X1  g210(.A1(new_n635), .A2(KEYINPUT14), .ZN(new_n636));
  XNOR2_X1  g211(.A(new_n631), .B(new_n636), .ZN(new_n637));
  NAND2_X1  g212(.A1(new_n637), .A2(G14), .ZN(new_n638));
  INV_X1    g213(.A(new_n638), .ZN(G401));
  XOR2_X1   g214(.A(G2084), .B(G2090), .Z(new_n640));
  XNOR2_X1  g215(.A(G2072), .B(G2078), .ZN(new_n641));
  XNOR2_X1  g216(.A(new_n641), .B(KEYINPUT17), .ZN(new_n642));
  XNOR2_X1  g217(.A(G2067), .B(G2678), .ZN(new_n643));
  AOI21_X1  g218(.A(new_n640), .B1(new_n642), .B2(new_n643), .ZN(new_n644));
  OAI21_X1  g219(.A(new_n644), .B1(new_n643), .B2(new_n641), .ZN(new_n645));
  XNOR2_X1  g220(.A(new_n645), .B(KEYINPUT80), .ZN(new_n646));
  NAND3_X1  g221(.A1(new_n640), .A2(new_n643), .A3(new_n641), .ZN(new_n647));
  XOR2_X1   g222(.A(new_n647), .B(KEYINPUT18), .Z(new_n648));
  INV_X1    g223(.A(new_n640), .ZN(new_n649));
  OR3_X1    g224(.A1(new_n642), .A2(new_n649), .A3(new_n643), .ZN(new_n650));
  NAND3_X1  g225(.A1(new_n646), .A2(new_n648), .A3(new_n650), .ZN(new_n651));
  XNOR2_X1  g226(.A(new_n651), .B(new_n622), .ZN(new_n652));
  NAND2_X1  g227(.A1(new_n652), .A2(G2100), .ZN(new_n653));
  XNOR2_X1  g228(.A(new_n651), .B(G2096), .ZN(new_n654));
  INV_X1    g229(.A(G2100), .ZN(new_n655));
  NAND2_X1  g230(.A1(new_n654), .A2(new_n655), .ZN(new_n656));
  NAND2_X1  g231(.A1(new_n653), .A2(new_n656), .ZN(G227));
  XNOR2_X1  g232(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n658));
  INV_X1    g233(.A(new_n658), .ZN(new_n659));
  XNOR2_X1  g234(.A(G1971), .B(G1976), .ZN(new_n660));
  XNOR2_X1  g235(.A(new_n660), .B(KEYINPUT81), .ZN(new_n661));
  XNOR2_X1  g236(.A(new_n661), .B(KEYINPUT19), .ZN(new_n662));
  XOR2_X1   g237(.A(G1956), .B(G2474), .Z(new_n663));
  XOR2_X1   g238(.A(G1961), .B(G1966), .Z(new_n664));
  AND2_X1   g239(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  NAND2_X1  g240(.A1(new_n662), .A2(new_n665), .ZN(new_n666));
  NAND2_X1  g241(.A1(new_n666), .A2(KEYINPUT82), .ZN(new_n667));
  INV_X1    g242(.A(KEYINPUT82), .ZN(new_n668));
  NAND3_X1  g243(.A1(new_n662), .A2(new_n668), .A3(new_n665), .ZN(new_n669));
  NAND2_X1  g244(.A1(new_n667), .A2(new_n669), .ZN(new_n670));
  INV_X1    g245(.A(KEYINPUT20), .ZN(new_n671));
  NAND2_X1  g246(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  NAND3_X1  g247(.A1(new_n667), .A2(KEYINPUT20), .A3(new_n669), .ZN(new_n673));
  NOR2_X1   g248(.A1(new_n663), .A2(new_n664), .ZN(new_n674));
  OR3_X1    g249(.A1(new_n662), .A2(new_n665), .A3(new_n674), .ZN(new_n675));
  NAND2_X1  g250(.A1(new_n662), .A2(new_n674), .ZN(new_n676));
  NAND4_X1  g251(.A1(new_n672), .A2(new_n673), .A3(new_n675), .A4(new_n676), .ZN(new_n677));
  XNOR2_X1  g252(.A(G1991), .B(G1996), .ZN(new_n678));
  INV_X1    g253(.A(new_n678), .ZN(new_n679));
  NAND2_X1  g254(.A1(new_n677), .A2(new_n679), .ZN(new_n680));
  AND2_X1   g255(.A1(new_n673), .A2(new_n676), .ZN(new_n681));
  NAND4_X1  g256(.A1(new_n681), .A2(new_n678), .A3(new_n675), .A4(new_n672), .ZN(new_n682));
  XOR2_X1   g257(.A(G1981), .B(G1986), .Z(new_n683));
  INV_X1    g258(.A(new_n683), .ZN(new_n684));
  NAND3_X1  g259(.A1(new_n680), .A2(new_n682), .A3(new_n684), .ZN(new_n685));
  INV_X1    g260(.A(new_n685), .ZN(new_n686));
  AOI21_X1  g261(.A(new_n684), .B1(new_n680), .B2(new_n682), .ZN(new_n687));
  OAI21_X1  g262(.A(new_n659), .B1(new_n686), .B2(new_n687), .ZN(new_n688));
  INV_X1    g263(.A(new_n687), .ZN(new_n689));
  NAND3_X1  g264(.A1(new_n689), .A2(new_n658), .A3(new_n685), .ZN(new_n690));
  NAND2_X1  g265(.A1(new_n688), .A2(new_n690), .ZN(new_n691));
  INV_X1    g266(.A(new_n691), .ZN(G229));
  XOR2_X1   g267(.A(KEYINPUT86), .B(KEYINPUT25), .Z(new_n693));
  NAND2_X1  g268(.A1(new_n469), .A2(G103), .ZN(new_n694));
  XNOR2_X1  g269(.A(new_n693), .B(new_n694), .ZN(new_n695));
  NAND2_X1  g270(.A1(new_n467), .A2(G139), .ZN(new_n696));
  AOI22_X1  g271(.A1(new_n493), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n697));
  OAI211_X1 g272(.A(new_n695), .B(new_n696), .C1(new_n475), .C2(new_n697), .ZN(new_n698));
  XOR2_X1   g273(.A(new_n698), .B(KEYINPUT87), .Z(new_n699));
  INV_X1    g274(.A(new_n699), .ZN(new_n700));
  NAND2_X1  g275(.A1(new_n700), .A2(G29), .ZN(new_n701));
  OAI21_X1  g276(.A(new_n701), .B1(G29), .B2(G33), .ZN(new_n702));
  XOR2_X1   g277(.A(new_n702), .B(G2072), .Z(new_n703));
  NAND3_X1  g278(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n704));
  XNOR2_X1  g279(.A(new_n704), .B(KEYINPUT90), .ZN(new_n705));
  XOR2_X1   g280(.A(new_n705), .B(KEYINPUT26), .Z(new_n706));
  AOI22_X1  g281(.A1(new_n477), .A2(G129), .B1(G141), .B2(new_n467), .ZN(new_n707));
  NAND2_X1  g282(.A1(new_n469), .A2(G105), .ZN(new_n708));
  XNOR2_X1  g283(.A(new_n708), .B(KEYINPUT89), .ZN(new_n709));
  NAND2_X1  g284(.A1(new_n707), .A2(new_n709), .ZN(new_n710));
  NOR2_X1   g285(.A1(new_n706), .A2(new_n710), .ZN(new_n711));
  NAND2_X1  g286(.A1(new_n711), .A2(G29), .ZN(new_n712));
  OAI21_X1  g287(.A(new_n712), .B1(G29), .B2(G32), .ZN(new_n713));
  INV_X1    g288(.A(new_n713), .ZN(new_n714));
  XNOR2_X1  g289(.A(KEYINPUT27), .B(G1996), .ZN(new_n715));
  XNOR2_X1  g290(.A(new_n715), .B(KEYINPUT91), .ZN(new_n716));
  NOR2_X1   g291(.A1(new_n714), .A2(new_n716), .ZN(new_n717));
  XOR2_X1   g292(.A(new_n717), .B(KEYINPUT92), .Z(new_n718));
  INV_X1    g293(.A(G16), .ZN(new_n719));
  NOR2_X1   g294(.A1(G286), .A2(new_n719), .ZN(new_n720));
  NOR2_X1   g295(.A1(G16), .A2(G21), .ZN(new_n721));
  NOR3_X1   g296(.A1(new_n720), .A2(KEYINPUT93), .A3(new_n721), .ZN(new_n722));
  AOI21_X1  g297(.A(new_n722), .B1(KEYINPUT93), .B2(new_n720), .ZN(new_n723));
  INV_X1    g298(.A(G1966), .ZN(new_n724));
  NOR2_X1   g299(.A1(new_n723), .A2(new_n724), .ZN(new_n725));
  INV_X1    g300(.A(G26), .ZN(new_n726));
  OR3_X1    g301(.A1(new_n726), .A2(KEYINPUT28), .A3(G29), .ZN(new_n727));
  NAND2_X1  g302(.A1(new_n477), .A2(G128), .ZN(new_n728));
  NAND2_X1  g303(.A1(new_n467), .A2(G140), .ZN(new_n729));
  OR2_X1    g304(.A1(G104), .A2(G2105), .ZN(new_n730));
  OAI211_X1 g305(.A(new_n730), .B(G2104), .C1(G116), .C2(new_n475), .ZN(new_n731));
  NAND3_X1  g306(.A1(new_n728), .A2(new_n729), .A3(new_n731), .ZN(new_n732));
  INV_X1    g307(.A(KEYINPUT85), .ZN(new_n733));
  OR2_X1    g308(.A1(new_n732), .A2(new_n733), .ZN(new_n734));
  NAND2_X1  g309(.A1(new_n732), .A2(new_n733), .ZN(new_n735));
  NAND2_X1  g310(.A1(new_n734), .A2(new_n735), .ZN(new_n736));
  INV_X1    g311(.A(new_n736), .ZN(new_n737));
  INV_X1    g312(.A(G29), .ZN(new_n738));
  NOR2_X1   g313(.A1(new_n737), .A2(new_n738), .ZN(new_n739));
  OAI21_X1  g314(.A(KEYINPUT28), .B1(new_n726), .B2(G29), .ZN(new_n740));
  OAI21_X1  g315(.A(new_n727), .B1(new_n739), .B2(new_n740), .ZN(new_n741));
  INV_X1    g316(.A(G2067), .ZN(new_n742));
  XNOR2_X1  g317(.A(new_n741), .B(new_n742), .ZN(new_n743));
  NOR3_X1   g318(.A1(new_n718), .A2(new_n725), .A3(new_n743), .ZN(new_n744));
  NAND2_X1  g319(.A1(new_n719), .A2(G20), .ZN(new_n745));
  INV_X1    g320(.A(G299), .ZN(new_n746));
  OAI211_X1 g321(.A(KEYINPUT23), .B(new_n745), .C1(new_n746), .C2(new_n719), .ZN(new_n747));
  OAI21_X1  g322(.A(new_n747), .B1(KEYINPUT23), .B2(new_n745), .ZN(new_n748));
  INV_X1    g323(.A(G1956), .ZN(new_n749));
  XNOR2_X1  g324(.A(new_n748), .B(new_n749), .ZN(new_n750));
  AOI21_X1  g325(.A(new_n750), .B1(new_n724), .B2(new_n723), .ZN(new_n751));
  NAND2_X1  g326(.A1(new_n719), .A2(G19), .ZN(new_n752));
  OAI21_X1  g327(.A(new_n752), .B1(new_n546), .B2(new_n719), .ZN(new_n753));
  XOR2_X1   g328(.A(new_n753), .B(G1341), .Z(new_n754));
  OR2_X1    g329(.A1(KEYINPUT24), .A2(G34), .ZN(new_n755));
  NAND2_X1  g330(.A1(KEYINPUT24), .A2(G34), .ZN(new_n756));
  NAND3_X1  g331(.A1(new_n755), .A2(new_n738), .A3(new_n756), .ZN(new_n757));
  OAI21_X1  g332(.A(new_n757), .B1(G160), .B2(new_n738), .ZN(new_n758));
  XNOR2_X1  g333(.A(new_n758), .B(KEYINPUT88), .ZN(new_n759));
  INV_X1    g334(.A(G2084), .ZN(new_n760));
  XNOR2_X1  g335(.A(new_n759), .B(new_n760), .ZN(new_n761));
  INV_X1    g336(.A(G1348), .ZN(new_n762));
  NOR2_X1   g337(.A1(new_n606), .A2(new_n719), .ZN(new_n763));
  AOI21_X1  g338(.A(new_n763), .B1(G4), .B2(new_n719), .ZN(new_n764));
  OAI21_X1  g339(.A(new_n761), .B1(new_n762), .B2(new_n764), .ZN(new_n765));
  INV_X1    g340(.A(G35), .ZN(new_n766));
  OAI21_X1  g341(.A(KEYINPUT95), .B1(new_n766), .B2(G29), .ZN(new_n767));
  OR3_X1    g342(.A1(new_n766), .A2(KEYINPUT95), .A3(G29), .ZN(new_n768));
  OAI211_X1 g343(.A(new_n767), .B(new_n768), .C1(G162), .C2(new_n738), .ZN(new_n769));
  XNOR2_X1  g344(.A(KEYINPUT96), .B(KEYINPUT29), .ZN(new_n770));
  XNOR2_X1  g345(.A(new_n770), .B(G2090), .ZN(new_n771));
  XNOR2_X1  g346(.A(new_n769), .B(new_n771), .ZN(new_n772));
  AND2_X1   g347(.A1(KEYINPUT30), .A2(G28), .ZN(new_n773));
  NOR2_X1   g348(.A1(KEYINPUT30), .A2(G28), .ZN(new_n774));
  OAI21_X1  g349(.A(new_n738), .B1(new_n773), .B2(new_n774), .ZN(new_n775));
  OAI21_X1  g350(.A(new_n775), .B1(new_n621), .B2(new_n738), .ZN(new_n776));
  NOR2_X1   g351(.A1(new_n772), .A2(new_n776), .ZN(new_n777));
  NAND2_X1  g352(.A1(new_n764), .A2(new_n762), .ZN(new_n778));
  NOR2_X1   g353(.A1(G27), .A2(G29), .ZN(new_n779));
  AOI21_X1  g354(.A(new_n779), .B1(G164), .B2(G29), .ZN(new_n780));
  XNOR2_X1  g355(.A(new_n780), .B(G2078), .ZN(new_n781));
  AOI21_X1  g356(.A(new_n781), .B1(new_n714), .B2(new_n716), .ZN(new_n782));
  XNOR2_X1  g357(.A(KEYINPUT31), .B(G11), .ZN(new_n783));
  NAND4_X1  g358(.A1(new_n777), .A2(new_n778), .A3(new_n782), .A4(new_n783), .ZN(new_n784));
  NAND2_X1  g359(.A1(new_n719), .A2(G5), .ZN(new_n785));
  OAI21_X1  g360(.A(new_n785), .B1(G171), .B2(new_n719), .ZN(new_n786));
  XOR2_X1   g361(.A(KEYINPUT94), .B(G1961), .Z(new_n787));
  XNOR2_X1  g362(.A(new_n786), .B(new_n787), .ZN(new_n788));
  NOR3_X1   g363(.A1(new_n765), .A2(new_n784), .A3(new_n788), .ZN(new_n789));
  NAND4_X1  g364(.A1(new_n744), .A2(new_n751), .A3(new_n754), .A4(new_n789), .ZN(new_n790));
  NAND2_X1  g365(.A1(new_n477), .A2(G119), .ZN(new_n791));
  NAND2_X1  g366(.A1(new_n467), .A2(G131), .ZN(new_n792));
  NOR2_X1   g367(.A1(G95), .A2(G2105), .ZN(new_n793));
  OAI21_X1  g368(.A(G2104), .B1(new_n475), .B2(G107), .ZN(new_n794));
  OAI211_X1 g369(.A(new_n791), .B(new_n792), .C1(new_n793), .C2(new_n794), .ZN(new_n795));
  MUX2_X1   g370(.A(G25), .B(new_n795), .S(G29), .Z(new_n796));
  XNOR2_X1  g371(.A(KEYINPUT35), .B(G1991), .ZN(new_n797));
  INV_X1    g372(.A(new_n797), .ZN(new_n798));
  XNOR2_X1  g373(.A(new_n796), .B(new_n798), .ZN(new_n799));
  NAND2_X1  g374(.A1(new_n719), .A2(G24), .ZN(new_n800));
  OAI21_X1  g375(.A(new_n800), .B1(new_n590), .B2(new_n719), .ZN(new_n801));
  INV_X1    g376(.A(new_n801), .ZN(new_n802));
  INV_X1    g377(.A(G1986), .ZN(new_n803));
  OAI21_X1  g378(.A(new_n799), .B1(new_n802), .B2(new_n803), .ZN(new_n804));
  NAND2_X1  g379(.A1(new_n719), .A2(G6), .ZN(new_n805));
  INV_X1    g380(.A(G305), .ZN(new_n806));
  OAI21_X1  g381(.A(new_n805), .B1(new_n806), .B2(new_n719), .ZN(new_n807));
  XNOR2_X1  g382(.A(new_n807), .B(KEYINPUT32), .ZN(new_n808));
  INV_X1    g383(.A(G1981), .ZN(new_n809));
  XNOR2_X1  g384(.A(new_n808), .B(new_n809), .ZN(new_n810));
  NAND2_X1  g385(.A1(new_n719), .A2(G22), .ZN(new_n811));
  OAI21_X1  g386(.A(new_n811), .B1(G166), .B2(new_n719), .ZN(new_n812));
  XNOR2_X1  g387(.A(new_n812), .B(KEYINPUT84), .ZN(new_n813));
  XOR2_X1   g388(.A(KEYINPUT83), .B(G1971), .Z(new_n814));
  XNOR2_X1  g389(.A(new_n813), .B(new_n814), .ZN(new_n815));
  NAND2_X1  g390(.A1(new_n719), .A2(G23), .ZN(new_n816));
  INV_X1    g391(.A(G288), .ZN(new_n817));
  OAI21_X1  g392(.A(new_n816), .B1(new_n817), .B2(new_n719), .ZN(new_n818));
  XNOR2_X1  g393(.A(new_n818), .B(KEYINPUT33), .ZN(new_n819));
  XNOR2_X1  g394(.A(new_n819), .B(G1976), .ZN(new_n820));
  NAND3_X1  g395(.A1(new_n810), .A2(new_n815), .A3(new_n820), .ZN(new_n821));
  AOI21_X1  g396(.A(new_n804), .B1(new_n821), .B2(KEYINPUT34), .ZN(new_n822));
  NAND2_X1  g397(.A1(new_n802), .A2(new_n803), .ZN(new_n823));
  OAI211_X1 g398(.A(new_n822), .B(new_n823), .C1(KEYINPUT34), .C2(new_n821), .ZN(new_n824));
  OR2_X1    g399(.A1(new_n824), .A2(KEYINPUT36), .ZN(new_n825));
  NAND2_X1  g400(.A1(new_n824), .A2(KEYINPUT36), .ZN(new_n826));
  AOI211_X1 g401(.A(new_n703), .B(new_n790), .C1(new_n825), .C2(new_n826), .ZN(G311));
  AOI21_X1  g402(.A(new_n790), .B1(new_n825), .B2(new_n826), .ZN(new_n828));
  INV_X1    g403(.A(new_n703), .ZN(new_n829));
  NAND2_X1  g404(.A1(new_n828), .A2(new_n829), .ZN(G150));
  AOI22_X1  g405(.A1(new_n516), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n831));
  NOR2_X1   g406(.A1(new_n831), .A2(new_n504), .ZN(new_n832));
  INV_X1    g407(.A(G93), .ZN(new_n833));
  INV_X1    g408(.A(G55), .ZN(new_n834));
  OAI22_X1  g409(.A1(new_n507), .A2(new_n833), .B1(new_n509), .B2(new_n834), .ZN(new_n835));
  OR2_X1    g410(.A1(new_n832), .A2(new_n835), .ZN(new_n836));
  NAND2_X1  g411(.A1(new_n836), .A2(G860), .ZN(new_n837));
  XOR2_X1   g412(.A(new_n837), .B(KEYINPUT37), .Z(new_n838));
  NAND3_X1  g413(.A1(new_n543), .A2(new_n544), .A3(new_n545), .ZN(new_n839));
  NOR2_X1   g414(.A1(new_n832), .A2(new_n835), .ZN(new_n840));
  NAND2_X1  g415(.A1(new_n839), .A2(new_n840), .ZN(new_n841));
  AOI22_X1  g416(.A1(new_n540), .A2(new_n542), .B1(G43), .B2(new_n518), .ZN(new_n842));
  NAND3_X1  g417(.A1(new_n842), .A2(new_n836), .A3(new_n544), .ZN(new_n843));
  NAND2_X1  g418(.A1(new_n841), .A2(new_n843), .ZN(new_n844));
  XNOR2_X1  g419(.A(new_n844), .B(KEYINPUT39), .ZN(new_n845));
  NAND2_X1  g420(.A1(new_n606), .A2(G559), .ZN(new_n846));
  XNOR2_X1  g421(.A(new_n846), .B(KEYINPUT38), .ZN(new_n847));
  XNOR2_X1  g422(.A(new_n845), .B(new_n847), .ZN(new_n848));
  OAI21_X1  g423(.A(new_n838), .B1(new_n848), .B2(G860), .ZN(G145));
  XNOR2_X1  g424(.A(KEYINPUT97), .B(G37), .ZN(new_n850));
  NAND2_X1  g425(.A1(new_n477), .A2(G130), .ZN(new_n851));
  NOR2_X1   g426(.A1(G106), .A2(G2105), .ZN(new_n852));
  OAI21_X1  g427(.A(G2104), .B1(new_n475), .B2(G118), .ZN(new_n853));
  OAI21_X1  g428(.A(new_n851), .B1(new_n852), .B2(new_n853), .ZN(new_n854));
  AOI21_X1  g429(.A(new_n854), .B1(G142), .B2(new_n467), .ZN(new_n855));
  XNOR2_X1  g430(.A(new_n855), .B(new_n614), .ZN(new_n856));
  XNOR2_X1  g431(.A(new_n856), .B(new_n795), .ZN(new_n857));
  INV_X1    g432(.A(new_n857), .ZN(new_n858));
  NAND2_X1  g433(.A1(new_n736), .A2(new_n711), .ZN(new_n859));
  OAI211_X1 g434(.A(new_n734), .B(new_n735), .C1(new_n710), .C2(new_n706), .ZN(new_n860));
  NAND2_X1  g435(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  NAND2_X1  g436(.A1(new_n492), .A2(new_n495), .ZN(new_n862));
  AND2_X1   g437(.A1(new_n488), .A2(new_n489), .ZN(new_n863));
  NAND2_X1  g438(.A1(new_n862), .A2(new_n863), .ZN(new_n864));
  NAND2_X1  g439(.A1(new_n861), .A2(new_n864), .ZN(new_n865));
  NAND3_X1  g440(.A1(new_n859), .A2(G164), .A3(new_n860), .ZN(new_n866));
  AND3_X1   g441(.A1(new_n865), .A2(new_n698), .A3(new_n866), .ZN(new_n867));
  AOI21_X1  g442(.A(new_n699), .B1(new_n865), .B2(new_n866), .ZN(new_n868));
  OAI21_X1  g443(.A(new_n858), .B1(new_n867), .B2(new_n868), .ZN(new_n869));
  NAND2_X1  g444(.A1(new_n865), .A2(new_n866), .ZN(new_n870));
  NAND2_X1  g445(.A1(new_n870), .A2(new_n700), .ZN(new_n871));
  NAND3_X1  g446(.A1(new_n865), .A2(new_n698), .A3(new_n866), .ZN(new_n872));
  NAND3_X1  g447(.A1(new_n871), .A2(new_n857), .A3(new_n872), .ZN(new_n873));
  NAND2_X1  g448(.A1(new_n869), .A2(new_n873), .ZN(new_n874));
  XOR2_X1   g449(.A(G160), .B(new_n480), .Z(new_n875));
  XNOR2_X1  g450(.A(new_n875), .B(new_n621), .ZN(new_n876));
  AOI21_X1  g451(.A(new_n850), .B1(new_n874), .B2(new_n876), .ZN(new_n877));
  NAND2_X1  g452(.A1(new_n869), .A2(KEYINPUT98), .ZN(new_n878));
  INV_X1    g453(.A(KEYINPUT98), .ZN(new_n879));
  OAI211_X1 g454(.A(new_n858), .B(new_n879), .C1(new_n867), .C2(new_n868), .ZN(new_n880));
  NAND3_X1  g455(.A1(new_n878), .A2(new_n873), .A3(new_n880), .ZN(new_n881));
  XOR2_X1   g456(.A(new_n876), .B(KEYINPUT99), .Z(new_n882));
  OAI21_X1  g457(.A(new_n877), .B1(new_n881), .B2(new_n882), .ZN(new_n883));
  XNOR2_X1  g458(.A(new_n883), .B(KEYINPUT40), .ZN(G395));
  XNOR2_X1  g459(.A(new_n844), .B(new_n609), .ZN(new_n885));
  XNOR2_X1  g460(.A(G299), .B(new_n598), .ZN(new_n886));
  NOR2_X1   g461(.A1(new_n885), .A2(new_n886), .ZN(new_n887));
  INV_X1    g462(.A(KEYINPUT41), .ZN(new_n888));
  NAND2_X1  g463(.A1(new_n606), .A2(G299), .ZN(new_n889));
  AOI22_X1  g464(.A1(new_n558), .A2(new_n560), .B1(G91), .B2(new_n531), .ZN(new_n890));
  NAND3_X1  g465(.A1(new_n598), .A2(new_n890), .A3(new_n564), .ZN(new_n891));
  AOI21_X1  g466(.A(KEYINPUT100), .B1(new_n889), .B2(new_n891), .ZN(new_n892));
  OAI21_X1  g467(.A(KEYINPUT100), .B1(new_n606), .B2(G299), .ZN(new_n893));
  INV_X1    g468(.A(new_n893), .ZN(new_n894));
  OAI21_X1  g469(.A(new_n888), .B1(new_n892), .B2(new_n894), .ZN(new_n895));
  INV_X1    g470(.A(new_n886), .ZN(new_n896));
  OAI21_X1  g471(.A(new_n895), .B1(new_n888), .B2(new_n896), .ZN(new_n897));
  AOI21_X1  g472(.A(new_n887), .B1(new_n885), .B2(new_n897), .ZN(new_n898));
  INV_X1    g473(.A(KEYINPUT42), .ZN(new_n899));
  NOR2_X1   g474(.A1(new_n817), .A2(G303), .ZN(new_n900));
  NOR2_X1   g475(.A1(G288), .A2(G166), .ZN(new_n901));
  OAI21_X1  g476(.A(new_n590), .B1(new_n900), .B2(new_n901), .ZN(new_n902));
  INV_X1    g477(.A(new_n902), .ZN(new_n903));
  NOR3_X1   g478(.A1(new_n900), .A2(new_n590), .A3(new_n901), .ZN(new_n904));
  NOR3_X1   g479(.A1(new_n903), .A2(G305), .A3(new_n904), .ZN(new_n905));
  OR3_X1    g480(.A1(new_n900), .A2(new_n590), .A3(new_n901), .ZN(new_n906));
  AOI21_X1  g481(.A(new_n806), .B1(new_n906), .B2(new_n902), .ZN(new_n907));
  OAI21_X1  g482(.A(new_n899), .B1(new_n905), .B2(new_n907), .ZN(new_n908));
  INV_X1    g483(.A(KEYINPUT101), .ZN(new_n909));
  OAI21_X1  g484(.A(new_n909), .B1(new_n905), .B2(new_n907), .ZN(new_n910));
  OAI21_X1  g485(.A(G305), .B1(new_n903), .B2(new_n904), .ZN(new_n911));
  NAND3_X1  g486(.A1(new_n906), .A2(new_n806), .A3(new_n902), .ZN(new_n912));
  NAND3_X1  g487(.A1(new_n911), .A2(KEYINPUT101), .A3(new_n912), .ZN(new_n913));
  NAND2_X1  g488(.A1(new_n910), .A2(new_n913), .ZN(new_n914));
  OAI21_X1  g489(.A(new_n908), .B1(new_n914), .B2(new_n899), .ZN(new_n915));
  OR2_X1    g490(.A1(new_n898), .A2(new_n915), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n898), .A2(new_n915), .ZN(new_n917));
  NAND3_X1  g492(.A1(new_n916), .A2(G868), .A3(new_n917), .ZN(new_n918));
  NOR2_X1   g493(.A1(new_n840), .A2(G868), .ZN(new_n919));
  OAI21_X1  g494(.A(new_n918), .B1(KEYINPUT102), .B2(new_n919), .ZN(new_n920));
  OAI21_X1  g495(.A(new_n920), .B1(KEYINPUT102), .B2(new_n918), .ZN(G295));
  OAI21_X1  g496(.A(new_n920), .B1(KEYINPUT102), .B2(new_n918), .ZN(G331));
  XNOR2_X1  g497(.A(G286), .B(G301), .ZN(new_n923));
  INV_X1    g498(.A(new_n923), .ZN(new_n924));
  NOR2_X1   g499(.A1(new_n839), .A2(new_n840), .ZN(new_n925));
  AOI21_X1  g500(.A(new_n836), .B1(new_n842), .B2(new_n544), .ZN(new_n926));
  OAI21_X1  g501(.A(new_n924), .B1(new_n925), .B2(new_n926), .ZN(new_n927));
  NAND3_X1  g502(.A1(new_n841), .A2(new_n923), .A3(new_n843), .ZN(new_n928));
  NAND3_X1  g503(.A1(new_n927), .A2(KEYINPUT103), .A3(new_n928), .ZN(new_n929));
  INV_X1    g504(.A(KEYINPUT103), .ZN(new_n930));
  NAND4_X1  g505(.A1(new_n841), .A2(new_n843), .A3(new_n923), .A4(new_n930), .ZN(new_n931));
  NAND3_X1  g506(.A1(new_n929), .A2(new_n897), .A3(new_n931), .ZN(new_n932));
  NAND3_X1  g507(.A1(new_n927), .A2(new_n896), .A3(new_n928), .ZN(new_n933));
  INV_X1    g508(.A(KEYINPUT104), .ZN(new_n934));
  NAND2_X1  g509(.A1(new_n933), .A2(new_n934), .ZN(new_n935));
  NAND4_X1  g510(.A1(new_n927), .A2(KEYINPUT104), .A3(new_n896), .A4(new_n928), .ZN(new_n936));
  NAND3_X1  g511(.A1(new_n932), .A2(new_n935), .A3(new_n936), .ZN(new_n937));
  INV_X1    g512(.A(new_n914), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n937), .A2(new_n938), .ZN(new_n939));
  INV_X1    g514(.A(G37), .ZN(new_n940));
  NAND4_X1  g515(.A1(new_n914), .A2(new_n932), .A3(new_n935), .A4(new_n936), .ZN(new_n941));
  NAND3_X1  g516(.A1(new_n939), .A2(new_n940), .A3(new_n941), .ZN(new_n942));
  INV_X1    g517(.A(KEYINPUT43), .ZN(new_n943));
  AND2_X1   g518(.A1(new_n942), .A2(new_n943), .ZN(new_n944));
  INV_X1    g519(.A(new_n850), .ZN(new_n945));
  OAI21_X1  g520(.A(new_n893), .B1(new_n886), .B2(KEYINPUT100), .ZN(new_n946));
  AOI211_X1 g521(.A(new_n888), .B(new_n946), .C1(new_n927), .C2(new_n928), .ZN(new_n947));
  NAND2_X1  g522(.A1(new_n946), .A2(KEYINPUT41), .ZN(new_n948));
  INV_X1    g523(.A(new_n928), .ZN(new_n949));
  AOI21_X1  g524(.A(new_n923), .B1(new_n841), .B2(new_n843), .ZN(new_n950));
  OAI21_X1  g525(.A(new_n948), .B1(new_n949), .B2(new_n950), .ZN(new_n951));
  NAND3_X1  g526(.A1(new_n951), .A2(new_n931), .A3(new_n929), .ZN(new_n952));
  AOI21_X1  g527(.A(new_n947), .B1(new_n952), .B2(new_n896), .ZN(new_n953));
  OAI211_X1 g528(.A(new_n945), .B(new_n941), .C1(new_n953), .C2(new_n914), .ZN(new_n954));
  NOR2_X1   g529(.A1(new_n954), .A2(new_n943), .ZN(new_n955));
  OAI21_X1  g530(.A(KEYINPUT44), .B1(new_n944), .B2(new_n955), .ZN(new_n956));
  AND2_X1   g531(.A1(new_n942), .A2(KEYINPUT43), .ZN(new_n957));
  NOR2_X1   g532(.A1(new_n954), .A2(KEYINPUT43), .ZN(new_n958));
  NOR2_X1   g533(.A1(new_n957), .A2(new_n958), .ZN(new_n959));
  OAI21_X1  g534(.A(new_n956), .B1(new_n959), .B2(KEYINPUT44), .ZN(G397));
  NAND2_X1  g535(.A1(G305), .A2(G1981), .ZN(new_n961));
  OAI21_X1  g536(.A(G651), .B1(new_n580), .B2(new_n581), .ZN(new_n962));
  INV_X1    g537(.A(KEYINPUT78), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n962), .A2(new_n963), .ZN(new_n964));
  AOI21_X1  g539(.A(new_n571), .B1(new_n964), .B2(new_n582), .ZN(new_n965));
  NAND3_X1  g540(.A1(new_n965), .A2(new_n809), .A3(new_n570), .ZN(new_n966));
  NAND3_X1  g541(.A1(new_n961), .A2(KEYINPUT49), .A3(new_n966), .ZN(new_n967));
  INV_X1    g542(.A(G8), .ZN(new_n968));
  NAND3_X1  g543(.A1(new_n464), .A2(G40), .A3(new_n470), .ZN(new_n969));
  INV_X1    g544(.A(new_n969), .ZN(new_n970));
  AOI21_X1  g545(.A(G1384), .B1(new_n862), .B2(new_n863), .ZN(new_n971));
  AOI21_X1  g546(.A(new_n968), .B1(new_n970), .B2(new_n971), .ZN(new_n972));
  AND2_X1   g547(.A1(new_n967), .A2(new_n972), .ZN(new_n973));
  INV_X1    g548(.A(KEYINPUT49), .ZN(new_n974));
  NOR2_X1   g549(.A1(G305), .A2(G1981), .ZN(new_n975));
  AOI21_X1  g550(.A(new_n809), .B1(new_n965), .B2(new_n570), .ZN(new_n976));
  OAI21_X1  g551(.A(new_n974), .B1(new_n975), .B2(new_n976), .ZN(new_n977));
  NAND2_X1  g552(.A1(new_n977), .A2(KEYINPUT110), .ZN(new_n978));
  NAND2_X1  g553(.A1(new_n961), .A2(new_n966), .ZN(new_n979));
  INV_X1    g554(.A(KEYINPUT110), .ZN(new_n980));
  NAND3_X1  g555(.A1(new_n979), .A2(new_n980), .A3(new_n974), .ZN(new_n981));
  NAND3_X1  g556(.A1(new_n973), .A2(new_n978), .A3(new_n981), .ZN(new_n982));
  NAND3_X1  g557(.A1(G303), .A2(KEYINPUT55), .A3(G8), .ZN(new_n983));
  INV_X1    g558(.A(KEYINPUT55), .ZN(new_n984));
  OAI21_X1  g559(.A(new_n984), .B1(G166), .B2(new_n968), .ZN(new_n985));
  NAND2_X1  g560(.A1(new_n983), .A2(new_n985), .ZN(new_n986));
  XNOR2_X1  g561(.A(KEYINPUT108), .B(KEYINPUT50), .ZN(new_n987));
  INV_X1    g562(.A(new_n987), .ZN(new_n988));
  AOI21_X1  g563(.A(new_n969), .B1(new_n971), .B2(new_n988), .ZN(new_n989));
  INV_X1    g564(.A(G2090), .ZN(new_n990));
  OAI21_X1  g565(.A(KEYINPUT50), .B1(G164), .B2(G1384), .ZN(new_n991));
  AND3_X1   g566(.A1(new_n989), .A2(new_n990), .A3(new_n991), .ZN(new_n992));
  AOI21_X1  g567(.A(new_n969), .B1(new_n971), .B2(KEYINPUT45), .ZN(new_n993));
  XOR2_X1   g568(.A(KEYINPUT106), .B(KEYINPUT45), .Z(new_n994));
  INV_X1    g569(.A(new_n994), .ZN(new_n995));
  OAI21_X1  g570(.A(new_n995), .B1(G164), .B2(G1384), .ZN(new_n996));
  AOI21_X1  g571(.A(G1971), .B1(new_n993), .B2(new_n996), .ZN(new_n997));
  OAI211_X1 g572(.A(new_n986), .B(G8), .C1(new_n992), .C2(new_n997), .ZN(new_n998));
  INV_X1    g573(.A(KEYINPUT50), .ZN(new_n999));
  INV_X1    g574(.A(G1384), .ZN(new_n1000));
  NAND3_X1  g575(.A1(new_n864), .A2(new_n999), .A3(new_n1000), .ZN(new_n1001));
  NAND2_X1  g576(.A1(new_n1001), .A2(new_n970), .ZN(new_n1002));
  NOR2_X1   g577(.A1(new_n971), .A2(new_n988), .ZN(new_n1003));
  NOR3_X1   g578(.A1(new_n1002), .A2(G2090), .A3(new_n1003), .ZN(new_n1004));
  OAI21_X1  g579(.A(G8), .B1(new_n1004), .B2(new_n997), .ZN(new_n1005));
  NAND3_X1  g580(.A1(new_n1005), .A2(new_n985), .A3(new_n983), .ZN(new_n1006));
  INV_X1    g581(.A(G1976), .ZN(new_n1007));
  OAI21_X1  g582(.A(new_n972), .B1(new_n1007), .B2(G288), .ZN(new_n1008));
  INV_X1    g583(.A(KEYINPUT109), .ZN(new_n1009));
  INV_X1    g584(.A(KEYINPUT52), .ZN(new_n1010));
  OAI21_X1  g585(.A(new_n1008), .B1(new_n1009), .B2(new_n1010), .ZN(new_n1011));
  NOR2_X1   g586(.A1(new_n1009), .A2(new_n1010), .ZN(new_n1012));
  OAI211_X1 g587(.A(new_n972), .B(new_n1012), .C1(new_n1007), .C2(G288), .ZN(new_n1013));
  NAND3_X1  g588(.A1(G288), .A2(new_n1010), .A3(new_n1007), .ZN(new_n1014));
  NAND3_X1  g589(.A1(new_n1011), .A2(new_n1013), .A3(new_n1014), .ZN(new_n1015));
  NAND4_X1  g590(.A1(new_n982), .A2(new_n998), .A3(new_n1006), .A4(new_n1015), .ZN(new_n1016));
  AND3_X1   g591(.A1(new_n989), .A2(new_n760), .A3(new_n991), .ZN(new_n1017));
  AOI21_X1  g592(.A(new_n969), .B1(new_n971), .B2(new_n994), .ZN(new_n1018));
  INV_X1    g593(.A(KEYINPUT45), .ZN(new_n1019));
  OAI21_X1  g594(.A(new_n1019), .B1(G164), .B2(G1384), .ZN(new_n1020));
  AOI21_X1  g595(.A(G1966), .B1(new_n1018), .B2(new_n1020), .ZN(new_n1021));
  OAI21_X1  g596(.A(G8), .B1(new_n1017), .B2(new_n1021), .ZN(new_n1022));
  NAND2_X1  g597(.A1(G286), .A2(G8), .ZN(new_n1023));
  INV_X1    g598(.A(KEYINPUT51), .ZN(new_n1024));
  INV_X1    g599(.A(KEYINPUT120), .ZN(new_n1025));
  AOI21_X1  g600(.A(new_n1024), .B1(new_n1023), .B2(new_n1025), .ZN(new_n1026));
  NAND3_X1  g601(.A1(new_n1022), .A2(new_n1023), .A3(new_n1026), .ZN(new_n1027));
  INV_X1    g602(.A(new_n519), .ZN(new_n1028));
  NAND2_X1  g603(.A1(new_n522), .A2(new_n525), .ZN(new_n1029));
  NAND2_X1  g604(.A1(new_n1029), .A2(KEYINPUT74), .ZN(new_n1030));
  AOI21_X1  g605(.A(new_n1028), .B1(new_n1030), .B2(new_n526), .ZN(new_n1031));
  AOI21_X1  g606(.A(new_n968), .B1(new_n1031), .B2(new_n517), .ZN(new_n1032));
  OAI21_X1  g607(.A(KEYINPUT51), .B1(new_n1032), .B2(KEYINPUT120), .ZN(new_n1033));
  NAND3_X1  g608(.A1(new_n864), .A2(new_n1000), .A3(new_n994), .ZN(new_n1034));
  NAND2_X1  g609(.A1(new_n1034), .A2(new_n970), .ZN(new_n1035));
  NOR2_X1   g610(.A1(new_n971), .A2(KEYINPUT45), .ZN(new_n1036));
  OAI21_X1  g611(.A(new_n724), .B1(new_n1035), .B2(new_n1036), .ZN(new_n1037));
  NAND3_X1  g612(.A1(new_n989), .A2(new_n760), .A3(new_n991), .ZN(new_n1038));
  NAND2_X1  g613(.A1(new_n1037), .A2(new_n1038), .ZN(new_n1039));
  OAI211_X1 g614(.A(G8), .B(new_n1033), .C1(new_n1039), .C2(G286), .ZN(new_n1040));
  AOI21_X1  g615(.A(new_n968), .B1(new_n1037), .B2(new_n1038), .ZN(new_n1041));
  NAND2_X1  g616(.A1(new_n1041), .A2(G286), .ZN(new_n1042));
  AND3_X1   g617(.A1(new_n1027), .A2(new_n1040), .A3(new_n1042), .ZN(new_n1043));
  NOR2_X1   g618(.A1(new_n1016), .A2(new_n1043), .ZN(new_n1044));
  INV_X1    g619(.A(KEYINPUT53), .ZN(new_n1045));
  NAND2_X1  g620(.A1(new_n993), .A2(new_n996), .ZN(new_n1046));
  OAI21_X1  g621(.A(new_n1045), .B1(new_n1046), .B2(G2078), .ZN(new_n1047));
  NOR2_X1   g622(.A1(new_n1045), .A2(G2078), .ZN(new_n1048));
  NAND3_X1  g623(.A1(new_n1018), .A2(new_n1048), .A3(new_n1020), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n989), .A2(new_n991), .ZN(new_n1050));
  XNOR2_X1  g625(.A(KEYINPUT121), .B(G1961), .ZN(new_n1051));
  NAND2_X1  g626(.A1(new_n1050), .A2(new_n1051), .ZN(new_n1052));
  NAND3_X1  g627(.A1(new_n1047), .A2(new_n1049), .A3(new_n1052), .ZN(new_n1053));
  NAND2_X1  g628(.A1(new_n1053), .A2(G171), .ZN(new_n1054));
  INV_X1    g629(.A(KEYINPUT105), .ZN(new_n1055));
  OAI21_X1  g630(.A(new_n1055), .B1(G164), .B2(G1384), .ZN(new_n1056));
  NAND3_X1  g631(.A1(new_n864), .A2(KEYINPUT105), .A3(new_n1000), .ZN(new_n1057));
  NAND3_X1  g632(.A1(new_n1056), .A2(new_n995), .A3(new_n1057), .ZN(new_n1058));
  NAND2_X1  g633(.A1(new_n1058), .A2(new_n970), .ZN(new_n1059));
  NAND2_X1  g634(.A1(new_n1059), .A2(KEYINPUT122), .ZN(new_n1060));
  INV_X1    g635(.A(new_n971), .ZN(new_n1061));
  NOR2_X1   g636(.A1(new_n1061), .A2(new_n1019), .ZN(new_n1062));
  INV_X1    g637(.A(new_n1062), .ZN(new_n1063));
  INV_X1    g638(.A(KEYINPUT122), .ZN(new_n1064));
  NAND3_X1  g639(.A1(new_n1058), .A2(new_n1064), .A3(new_n970), .ZN(new_n1065));
  NAND4_X1  g640(.A1(new_n1060), .A2(new_n1048), .A3(new_n1063), .A4(new_n1065), .ZN(new_n1066));
  AND2_X1   g641(.A1(new_n1047), .A2(new_n1052), .ZN(new_n1067));
  NAND2_X1  g642(.A1(new_n1066), .A2(new_n1067), .ZN(new_n1068));
  OAI21_X1  g643(.A(new_n1054), .B1(new_n1068), .B2(G171), .ZN(new_n1069));
  INV_X1    g644(.A(KEYINPUT54), .ZN(new_n1070));
  NAND2_X1  g645(.A1(new_n1069), .A2(new_n1070), .ZN(new_n1071));
  NAND2_X1  g646(.A1(new_n1068), .A2(G171), .ZN(new_n1072));
  NAND4_X1  g647(.A1(new_n1047), .A2(new_n1052), .A3(G301), .A4(new_n1049), .ZN(new_n1073));
  AND2_X1   g648(.A1(new_n1073), .A2(KEYINPUT54), .ZN(new_n1074));
  AOI21_X1  g649(.A(KEYINPUT123), .B1(new_n1072), .B2(new_n1074), .ZN(new_n1075));
  AOI21_X1  g650(.A(G301), .B1(new_n1066), .B2(new_n1067), .ZN(new_n1076));
  INV_X1    g651(.A(KEYINPUT123), .ZN(new_n1077));
  NAND2_X1  g652(.A1(new_n1073), .A2(KEYINPUT54), .ZN(new_n1078));
  NOR3_X1   g653(.A1(new_n1076), .A2(new_n1077), .A3(new_n1078), .ZN(new_n1079));
  OAI211_X1 g654(.A(new_n1044), .B(new_n1071), .C1(new_n1075), .C2(new_n1079), .ZN(new_n1080));
  OAI21_X1  g655(.A(new_n749), .B1(new_n1002), .B2(new_n1003), .ZN(new_n1081));
  XNOR2_X1  g656(.A(KEYINPUT56), .B(G2072), .ZN(new_n1082));
  NAND3_X1  g657(.A1(new_n993), .A2(new_n996), .A3(new_n1082), .ZN(new_n1083));
  NAND2_X1  g658(.A1(new_n1081), .A2(new_n1083), .ZN(new_n1084));
  INV_X1    g659(.A(KEYINPUT57), .ZN(new_n1085));
  NAND2_X1  g660(.A1(G299), .A2(new_n1085), .ZN(new_n1086));
  NAND3_X1  g661(.A1(new_n890), .A2(KEYINPUT57), .A3(new_n564), .ZN(new_n1087));
  AND2_X1   g662(.A1(new_n1086), .A2(new_n1087), .ZN(new_n1088));
  NAND2_X1  g663(.A1(new_n1084), .A2(new_n1088), .ZN(new_n1089));
  INV_X1    g664(.A(KEYINPUT114), .ZN(new_n1090));
  NAND2_X1  g665(.A1(new_n1089), .A2(new_n1090), .ZN(new_n1091));
  NAND3_X1  g666(.A1(new_n1084), .A2(new_n1088), .A3(KEYINPUT114), .ZN(new_n1092));
  NAND2_X1  g667(.A1(new_n1091), .A2(new_n1092), .ZN(new_n1093));
  AOI21_X1  g668(.A(G1348), .B1(new_n989), .B2(new_n991), .ZN(new_n1094));
  NAND2_X1  g669(.A1(new_n970), .A2(new_n971), .ZN(new_n1095));
  NOR2_X1   g670(.A1(new_n1095), .A2(G2067), .ZN(new_n1096));
  NOR2_X1   g671(.A1(new_n1094), .A2(new_n1096), .ZN(new_n1097));
  OAI21_X1  g672(.A(new_n1093), .B1(new_n598), .B2(new_n1097), .ZN(new_n1098));
  NAND2_X1  g673(.A1(new_n1086), .A2(new_n1087), .ZN(new_n1099));
  NAND3_X1  g674(.A1(new_n1099), .A2(new_n1081), .A3(new_n1083), .ZN(new_n1100));
  NAND2_X1  g675(.A1(new_n1098), .A2(new_n1100), .ZN(new_n1101));
  NAND2_X1  g676(.A1(new_n1100), .A2(KEYINPUT118), .ZN(new_n1102));
  AND3_X1   g677(.A1(new_n1084), .A2(new_n1088), .A3(KEYINPUT114), .ZN(new_n1103));
  AOI21_X1  g678(.A(KEYINPUT114), .B1(new_n1084), .B2(new_n1088), .ZN(new_n1104));
  OAI21_X1  g679(.A(new_n1102), .B1(new_n1103), .B2(new_n1104), .ZN(new_n1105));
  INV_X1    g680(.A(KEYINPUT118), .ZN(new_n1106));
  NAND4_X1  g681(.A1(new_n1099), .A2(new_n1106), .A3(new_n1081), .A4(new_n1083), .ZN(new_n1107));
  NAND2_X1  g682(.A1(new_n1107), .A2(KEYINPUT61), .ZN(new_n1108));
  OAI21_X1  g683(.A(KEYINPUT119), .B1(new_n1105), .B2(new_n1108), .ZN(new_n1109));
  NAND2_X1  g684(.A1(new_n1097), .A2(KEYINPUT60), .ZN(new_n1110));
  INV_X1    g685(.A(KEYINPUT60), .ZN(new_n1111));
  OAI21_X1  g686(.A(new_n1111), .B1(new_n1094), .B2(new_n1096), .ZN(new_n1112));
  AND3_X1   g687(.A1(new_n1110), .A2(new_n606), .A3(new_n1112), .ZN(new_n1113));
  XOR2_X1   g688(.A(KEYINPUT117), .B(KEYINPUT61), .Z(new_n1114));
  AOI21_X1  g689(.A(new_n1114), .B1(new_n1089), .B2(new_n1100), .ZN(new_n1115));
  NOR2_X1   g690(.A1(new_n1110), .A2(new_n606), .ZN(new_n1116));
  NOR3_X1   g691(.A1(new_n1113), .A2(new_n1115), .A3(new_n1116), .ZN(new_n1117));
  INV_X1    g692(.A(KEYINPUT119), .ZN(new_n1118));
  INV_X1    g693(.A(new_n1108), .ZN(new_n1119));
  NAND4_X1  g694(.A1(new_n1093), .A2(new_n1118), .A3(new_n1119), .A4(new_n1102), .ZN(new_n1120));
  XOR2_X1   g695(.A(KEYINPUT115), .B(G1341), .Z(new_n1121));
  XNOR2_X1  g696(.A(new_n1121), .B(KEYINPUT58), .ZN(new_n1122));
  NAND2_X1  g697(.A1(new_n1095), .A2(new_n1122), .ZN(new_n1123));
  OAI21_X1  g698(.A(new_n1123), .B1(new_n1046), .B2(G1996), .ZN(new_n1124));
  NAND2_X1  g699(.A1(new_n546), .A2(new_n1124), .ZN(new_n1125));
  INV_X1    g700(.A(KEYINPUT116), .ZN(new_n1126));
  OAI21_X1  g701(.A(KEYINPUT59), .B1(new_n1125), .B2(new_n1126), .ZN(new_n1127));
  NAND2_X1  g702(.A1(new_n1125), .A2(new_n1126), .ZN(new_n1128));
  NAND2_X1  g703(.A1(new_n1127), .A2(new_n1128), .ZN(new_n1129));
  NAND3_X1  g704(.A1(new_n1125), .A2(new_n1126), .A3(KEYINPUT59), .ZN(new_n1130));
  NAND2_X1  g705(.A1(new_n1129), .A2(new_n1130), .ZN(new_n1131));
  NAND4_X1  g706(.A1(new_n1109), .A2(new_n1117), .A3(new_n1120), .A4(new_n1131), .ZN(new_n1132));
  AOI21_X1  g707(.A(new_n1080), .B1(new_n1101), .B2(new_n1132), .ZN(new_n1133));
  NAND3_X1  g708(.A1(new_n982), .A2(new_n1007), .A3(new_n817), .ZN(new_n1134));
  NAND2_X1  g709(.A1(new_n1134), .A2(new_n966), .ZN(new_n1135));
  INV_X1    g710(.A(KEYINPUT112), .ZN(new_n1136));
  NAND2_X1  g711(.A1(new_n1135), .A2(new_n1136), .ZN(new_n1137));
  NAND3_X1  g712(.A1(new_n1134), .A2(KEYINPUT112), .A3(new_n966), .ZN(new_n1138));
  NAND3_X1  g713(.A1(new_n1137), .A2(new_n972), .A3(new_n1138), .ZN(new_n1139));
  NAND3_X1  g714(.A1(new_n983), .A2(KEYINPUT113), .A3(new_n985), .ZN(new_n1140));
  OAI211_X1 g715(.A(new_n1140), .B(G8), .C1(new_n992), .C2(new_n997), .ZN(new_n1141));
  NAND4_X1  g716(.A1(new_n1141), .A2(KEYINPUT63), .A3(new_n1041), .A4(G168), .ZN(new_n1142));
  OAI21_X1  g717(.A(G8), .B1(new_n992), .B2(new_n997), .ZN(new_n1143));
  INV_X1    g718(.A(new_n1140), .ZN(new_n1144));
  AOI21_X1  g719(.A(new_n1142), .B1(new_n1143), .B2(new_n1144), .ZN(new_n1145));
  INV_X1    g720(.A(KEYINPUT111), .ZN(new_n1146));
  AOI21_X1  g721(.A(new_n980), .B1(new_n979), .B2(new_n974), .ZN(new_n1147));
  AOI211_X1 g722(.A(KEYINPUT110), .B(KEYINPUT49), .C1(new_n961), .C2(new_n966), .ZN(new_n1148));
  NAND2_X1  g723(.A1(new_n967), .A2(new_n972), .ZN(new_n1149));
  NOR3_X1   g724(.A1(new_n1147), .A2(new_n1148), .A3(new_n1149), .ZN(new_n1150));
  INV_X1    g725(.A(new_n1015), .ZN(new_n1151));
  OAI21_X1  g726(.A(new_n1146), .B1(new_n1150), .B2(new_n1151), .ZN(new_n1152));
  NAND3_X1  g727(.A1(new_n982), .A2(KEYINPUT111), .A3(new_n1015), .ZN(new_n1153));
  NAND3_X1  g728(.A1(new_n1145), .A2(new_n1152), .A3(new_n1153), .ZN(new_n1154));
  INV_X1    g729(.A(KEYINPUT63), .ZN(new_n1155));
  NAND2_X1  g730(.A1(new_n1041), .A2(G168), .ZN(new_n1156));
  OAI21_X1  g731(.A(new_n1155), .B1(new_n1016), .B2(new_n1156), .ZN(new_n1157));
  NAND2_X1  g732(.A1(new_n1154), .A2(new_n1157), .ZN(new_n1158));
  INV_X1    g733(.A(new_n998), .ZN(new_n1159));
  NAND3_X1  g734(.A1(new_n1152), .A2(new_n1159), .A3(new_n1153), .ZN(new_n1160));
  NAND3_X1  g735(.A1(new_n1139), .A2(new_n1158), .A3(new_n1160), .ZN(new_n1161));
  OAI21_X1  g736(.A(KEYINPUT124), .B1(new_n1133), .B2(new_n1161), .ZN(new_n1162));
  AND3_X1   g737(.A1(new_n1139), .A2(new_n1160), .A3(new_n1158), .ZN(new_n1163));
  OAI21_X1  g738(.A(new_n1077), .B1(new_n1076), .B2(new_n1078), .ZN(new_n1164));
  NAND2_X1  g739(.A1(new_n1047), .A2(new_n1052), .ZN(new_n1165));
  AOI21_X1  g740(.A(new_n1064), .B1(new_n1058), .B2(new_n970), .ZN(new_n1166));
  INV_X1    g741(.A(new_n1048), .ZN(new_n1167));
  NOR3_X1   g742(.A1(new_n1166), .A2(new_n1167), .A3(new_n1062), .ZN(new_n1168));
  AOI21_X1  g743(.A(new_n1165), .B1(new_n1168), .B2(new_n1065), .ZN(new_n1169));
  OAI211_X1 g744(.A(new_n1074), .B(KEYINPUT123), .C1(new_n1169), .C2(G301), .ZN(new_n1170));
  NAND2_X1  g745(.A1(new_n1164), .A2(new_n1170), .ZN(new_n1171));
  AND3_X1   g746(.A1(new_n1171), .A2(new_n1071), .A3(new_n1044), .ZN(new_n1172));
  NAND2_X1  g747(.A1(new_n1132), .A2(new_n1101), .ZN(new_n1173));
  NAND2_X1  g748(.A1(new_n1172), .A2(new_n1173), .ZN(new_n1174));
  INV_X1    g749(.A(KEYINPUT124), .ZN(new_n1175));
  NAND3_X1  g750(.A1(new_n1163), .A2(new_n1174), .A3(new_n1175), .ZN(new_n1176));
  INV_X1    g751(.A(new_n1043), .ZN(new_n1177));
  AOI21_X1  g752(.A(new_n1054), .B1(new_n1177), .B2(KEYINPUT62), .ZN(new_n1178));
  INV_X1    g753(.A(new_n1016), .ZN(new_n1179));
  OAI211_X1 g754(.A(new_n1178), .B(new_n1179), .C1(KEYINPUT62), .C2(new_n1177), .ZN(new_n1180));
  NAND3_X1  g755(.A1(new_n1162), .A2(new_n1176), .A3(new_n1180), .ZN(new_n1181));
  NOR2_X1   g756(.A1(new_n1058), .A2(new_n969), .ZN(new_n1182));
  XNOR2_X1  g757(.A(new_n736), .B(new_n742), .ZN(new_n1183));
  INV_X1    g758(.A(new_n1183), .ZN(new_n1184));
  XOR2_X1   g759(.A(new_n711), .B(G1996), .Z(new_n1185));
  NOR2_X1   g760(.A1(new_n1184), .A2(new_n1185), .ZN(new_n1186));
  XNOR2_X1  g761(.A(new_n795), .B(new_n798), .ZN(new_n1187));
  NAND2_X1  g762(.A1(new_n1186), .A2(new_n1187), .ZN(new_n1188));
  NAND2_X1  g763(.A1(new_n590), .A2(new_n803), .ZN(new_n1189));
  INV_X1    g764(.A(KEYINPUT107), .ZN(new_n1190));
  NAND2_X1  g765(.A1(new_n1189), .A2(new_n1190), .ZN(new_n1191));
  NOR2_X1   g766(.A1(new_n590), .A2(new_n803), .ZN(new_n1192));
  MUX2_X1   g767(.A(new_n1191), .B(new_n1190), .S(new_n1192), .Z(new_n1193));
  OAI21_X1  g768(.A(new_n1182), .B1(new_n1188), .B2(new_n1193), .ZN(new_n1194));
  NAND2_X1  g769(.A1(new_n1181), .A2(new_n1194), .ZN(new_n1195));
  INV_X1    g770(.A(new_n1182), .ZN(new_n1196));
  NOR2_X1   g771(.A1(new_n1196), .A2(G1996), .ZN(new_n1197));
  INV_X1    g772(.A(KEYINPUT125), .ZN(new_n1198));
  NAND2_X1  g773(.A1(new_n1198), .A2(KEYINPUT46), .ZN(new_n1199));
  XNOR2_X1  g774(.A(new_n1197), .B(new_n1199), .ZN(new_n1200));
  INV_X1    g775(.A(new_n711), .ZN(new_n1201));
  OAI21_X1  g776(.A(new_n1182), .B1(new_n1184), .B2(new_n1201), .ZN(new_n1202));
  OAI211_X1 g777(.A(new_n1200), .B(new_n1202), .C1(new_n1198), .C2(KEYINPUT46), .ZN(new_n1203));
  XOR2_X1   g778(.A(new_n1203), .B(KEYINPUT47), .Z(new_n1204));
  NOR2_X1   g779(.A1(new_n1196), .A2(new_n1189), .ZN(new_n1205));
  XNOR2_X1  g780(.A(new_n1205), .B(KEYINPUT48), .ZN(new_n1206));
  AOI21_X1  g781(.A(new_n1206), .B1(new_n1188), .B2(new_n1182), .ZN(new_n1207));
  NOR2_X1   g782(.A1(new_n795), .A2(new_n797), .ZN(new_n1208));
  NAND2_X1  g783(.A1(new_n1186), .A2(new_n1208), .ZN(new_n1209));
  NAND2_X1  g784(.A1(new_n737), .A2(new_n742), .ZN(new_n1210));
  AOI21_X1  g785(.A(new_n1196), .B1(new_n1209), .B2(new_n1210), .ZN(new_n1211));
  NOR3_X1   g786(.A1(new_n1204), .A2(new_n1207), .A3(new_n1211), .ZN(new_n1212));
  NAND2_X1  g787(.A1(new_n1195), .A2(new_n1212), .ZN(G329));
  assign    G231 = 1'b0;
  AND2_X1   g788(.A1(new_n638), .A2(G319), .ZN(new_n1215));
  NAND3_X1  g789(.A1(new_n1215), .A2(new_n653), .A3(new_n656), .ZN(new_n1216));
  NAND2_X1  g790(.A1(new_n1216), .A2(KEYINPUT126), .ZN(new_n1217));
  INV_X1    g791(.A(KEYINPUT126), .ZN(new_n1218));
  NAND4_X1  g792(.A1(new_n1215), .A2(new_n653), .A3(new_n656), .A4(new_n1218), .ZN(new_n1219));
  NAND2_X1  g793(.A1(new_n1217), .A2(new_n1219), .ZN(new_n1220));
  AND3_X1   g794(.A1(new_n883), .A2(new_n691), .A3(new_n1220), .ZN(new_n1221));
  OAI21_X1  g795(.A(new_n1221), .B1(new_n957), .B2(new_n958), .ZN(G225));
  NAND2_X1  g796(.A1(G225), .A2(KEYINPUT127), .ZN(new_n1223));
  INV_X1    g797(.A(KEYINPUT127), .ZN(new_n1224));
  OAI211_X1 g798(.A(new_n1221), .B(new_n1224), .C1(new_n957), .C2(new_n958), .ZN(new_n1225));
  NAND2_X1  g799(.A1(new_n1223), .A2(new_n1225), .ZN(G308));
endmodule


