//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 1 0 0 1 1 1 1 1 0 1 1 0 0 0 1 0 1 1 0 1 0 1 0 1 0 1 0 0 1 0 1 0 0 1 1 0 1 1 0 0 1 1 1 1 0 1 0 1 0 0 1 0 1 0 1 1 0 1 0 0 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:23:41 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n634, new_n635, new_n636, new_n637,
    new_n638, new_n639, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n646, new_n647, new_n648, new_n649, new_n650, new_n651, new_n652,
    new_n653, new_n654, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n695, new_n696,
    new_n697, new_n698, new_n699, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n712,
    new_n713, new_n714, new_n716, new_n717, new_n719, new_n720, new_n721,
    new_n722, new_n723, new_n724, new_n725, new_n726, new_n727, new_n728,
    new_n729, new_n730, new_n731, new_n732, new_n734, new_n735, new_n736,
    new_n737, new_n738, new_n739, new_n740, new_n741, new_n742, new_n743,
    new_n744, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n758, new_n759,
    new_n760, new_n761, new_n762, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n784, new_n785, new_n786, new_n787, new_n788, new_n789,
    new_n790, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n906, new_n907, new_n908, new_n909, new_n910,
    new_n911, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n926, new_n927,
    new_n928, new_n929, new_n930, new_n931, new_n932, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n939, new_n940, new_n941, new_n942,
    new_n943, new_n944, new_n945, new_n947, new_n948, new_n949, new_n950,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n985, new_n986, new_n987,
    new_n988, new_n989, new_n990, new_n991, new_n992, new_n993, new_n994,
    new_n995, new_n996, new_n997;
  XOR2_X1   g000(.A(G119), .B(G128), .Z(new_n187));
  XNOR2_X1  g001(.A(KEYINPUT24), .B(G110), .ZN(new_n188));
  NAND2_X1  g002(.A1(new_n187), .A2(new_n188), .ZN(new_n189));
  INV_X1    g003(.A(KEYINPUT23), .ZN(new_n190));
  INV_X1    g004(.A(G119), .ZN(new_n191));
  OAI21_X1  g005(.A(new_n190), .B1(new_n191), .B2(G128), .ZN(new_n192));
  INV_X1    g006(.A(G128), .ZN(new_n193));
  NAND3_X1  g007(.A1(new_n193), .A2(KEYINPUT23), .A3(G119), .ZN(new_n194));
  OAI211_X1 g008(.A(new_n192), .B(new_n194), .C1(G119), .C2(new_n193), .ZN(new_n195));
  OAI21_X1  g009(.A(new_n189), .B1(new_n195), .B2(G110), .ZN(new_n196));
  INV_X1    g010(.A(KEYINPUT77), .ZN(new_n197));
  XNOR2_X1  g011(.A(new_n196), .B(new_n197), .ZN(new_n198));
  INV_X1    g012(.A(G140), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n199), .A2(G125), .ZN(new_n200));
  OR2_X1    g014(.A1(new_n200), .A2(KEYINPUT75), .ZN(new_n201));
  INV_X1    g015(.A(G125), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n202), .A2(G140), .ZN(new_n203));
  NAND3_X1  g017(.A1(new_n200), .A2(new_n203), .A3(KEYINPUT75), .ZN(new_n204));
  NAND3_X1  g018(.A1(new_n201), .A2(KEYINPUT16), .A3(new_n204), .ZN(new_n205));
  INV_X1    g019(.A(KEYINPUT16), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n200), .A2(new_n206), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n205), .A2(new_n207), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n208), .A2(G146), .ZN(new_n209));
  AND2_X1   g023(.A1(new_n200), .A2(new_n203), .ZN(new_n210));
  INV_X1    g024(.A(G146), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  NAND3_X1  g026(.A1(new_n198), .A2(new_n209), .A3(new_n212), .ZN(new_n213));
  INV_X1    g027(.A(KEYINPUT76), .ZN(new_n214));
  NAND3_X1  g028(.A1(new_n205), .A2(new_n211), .A3(new_n207), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n209), .A2(new_n215), .ZN(new_n216));
  NOR2_X1   g030(.A1(new_n187), .A2(new_n188), .ZN(new_n217));
  AOI21_X1  g031(.A(new_n217), .B1(G110), .B2(new_n195), .ZN(new_n218));
  AOI21_X1  g032(.A(new_n214), .B1(new_n216), .B2(new_n218), .ZN(new_n219));
  AND3_X1   g033(.A1(new_n205), .A2(new_n211), .A3(new_n207), .ZN(new_n220));
  AOI21_X1  g034(.A(new_n211), .B1(new_n205), .B2(new_n207), .ZN(new_n221));
  OAI211_X1 g035(.A(new_n214), .B(new_n218), .C1(new_n220), .C2(new_n221), .ZN(new_n222));
  INV_X1    g036(.A(new_n222), .ZN(new_n223));
  OAI21_X1  g037(.A(new_n213), .B1(new_n219), .B2(new_n223), .ZN(new_n224));
  XNOR2_X1  g038(.A(KEYINPUT22), .B(G137), .ZN(new_n225));
  INV_X1    g039(.A(G953), .ZN(new_n226));
  AND3_X1   g040(.A1(new_n226), .A2(G221), .A3(G234), .ZN(new_n227));
  XOR2_X1   g041(.A(new_n225), .B(new_n227), .Z(new_n228));
  INV_X1    g042(.A(new_n228), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n224), .A2(new_n229), .ZN(new_n230));
  OAI211_X1 g044(.A(new_n213), .B(new_n228), .C1(new_n219), .C2(new_n223), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n230), .A2(new_n231), .ZN(new_n232));
  INV_X1    g046(.A(G217), .ZN(new_n233));
  INV_X1    g047(.A(G902), .ZN(new_n234));
  AOI21_X1  g048(.A(new_n233), .B1(G234), .B2(new_n234), .ZN(new_n235));
  NOR3_X1   g049(.A1(new_n232), .A2(G902), .A3(new_n235), .ZN(new_n236));
  INV_X1    g050(.A(new_n236), .ZN(new_n237));
  NAND3_X1  g051(.A1(new_n230), .A2(new_n234), .A3(new_n231), .ZN(new_n238));
  INV_X1    g052(.A(KEYINPUT79), .ZN(new_n239));
  XNOR2_X1  g053(.A(KEYINPUT78), .B(KEYINPUT25), .ZN(new_n240));
  AND3_X1   g054(.A1(new_n238), .A2(new_n239), .A3(new_n240), .ZN(new_n241));
  AOI21_X1  g055(.A(new_n239), .B1(new_n238), .B2(new_n240), .ZN(new_n242));
  INV_X1    g056(.A(KEYINPUT25), .ZN(new_n243));
  NOR2_X1   g057(.A1(new_n238), .A2(new_n243), .ZN(new_n244));
  NOR3_X1   g058(.A1(new_n241), .A2(new_n242), .A3(new_n244), .ZN(new_n245));
  INV_X1    g059(.A(new_n235), .ZN(new_n246));
  OAI21_X1  g060(.A(new_n237), .B1(new_n245), .B2(new_n246), .ZN(new_n247));
  INV_X1    g061(.A(G137), .ZN(new_n248));
  AND3_X1   g062(.A1(new_n248), .A2(KEYINPUT11), .A3(G134), .ZN(new_n249));
  AND2_X1   g063(.A1(KEYINPUT65), .A2(G134), .ZN(new_n250));
  NOR2_X1   g064(.A1(KEYINPUT65), .A2(G134), .ZN(new_n251));
  OAI21_X1  g065(.A(new_n248), .B1(new_n250), .B2(new_n251), .ZN(new_n252));
  XNOR2_X1  g066(.A(KEYINPUT64), .B(KEYINPUT11), .ZN(new_n253));
  AOI21_X1  g067(.A(new_n249), .B1(new_n252), .B2(new_n253), .ZN(new_n254));
  INV_X1    g068(.A(KEYINPUT66), .ZN(new_n255));
  NOR2_X1   g069(.A1(new_n250), .A2(new_n251), .ZN(new_n256));
  AOI21_X1  g070(.A(new_n255), .B1(new_n256), .B2(G137), .ZN(new_n257));
  NOR4_X1   g071(.A1(new_n250), .A2(new_n251), .A3(KEYINPUT66), .A4(new_n248), .ZN(new_n258));
  OAI21_X1  g072(.A(new_n254), .B1(new_n257), .B2(new_n258), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n259), .A2(G131), .ZN(new_n260));
  INV_X1    g074(.A(KEYINPUT67), .ZN(new_n261));
  INV_X1    g075(.A(G131), .ZN(new_n262));
  OAI211_X1 g076(.A(new_n254), .B(new_n262), .C1(new_n257), .C2(new_n258), .ZN(new_n263));
  NAND3_X1  g077(.A1(new_n260), .A2(new_n261), .A3(new_n263), .ZN(new_n264));
  NOR2_X1   g078(.A1(KEYINPUT0), .A2(G128), .ZN(new_n265));
  INV_X1    g079(.A(new_n265), .ZN(new_n266));
  NAND2_X1  g080(.A1(new_n211), .A2(G143), .ZN(new_n267));
  INV_X1    g081(.A(G143), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n268), .A2(G146), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n267), .A2(new_n269), .ZN(new_n270));
  INV_X1    g084(.A(KEYINPUT0), .ZN(new_n271));
  NOR2_X1   g085(.A1(new_n271), .A2(new_n193), .ZN(new_n272));
  OAI21_X1  g086(.A(new_n266), .B1(new_n270), .B2(new_n272), .ZN(new_n273));
  INV_X1    g087(.A(new_n273), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n270), .A2(new_n272), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n274), .A2(new_n275), .ZN(new_n276));
  NAND3_X1  g090(.A1(new_n259), .A2(KEYINPUT67), .A3(G131), .ZN(new_n277));
  NAND3_X1  g091(.A1(new_n264), .A2(new_n276), .A3(new_n277), .ZN(new_n278));
  OAI22_X1  g092(.A1(new_n252), .A2(KEYINPUT68), .B1(G134), .B2(new_n248), .ZN(new_n279));
  INV_X1    g093(.A(KEYINPUT68), .ZN(new_n280));
  XNOR2_X1  g094(.A(KEYINPUT65), .B(G134), .ZN(new_n281));
  AOI21_X1  g095(.A(new_n280), .B1(new_n281), .B2(new_n248), .ZN(new_n282));
  OAI21_X1  g096(.A(G131), .B1(new_n279), .B2(new_n282), .ZN(new_n283));
  AND2_X1   g097(.A1(new_n267), .A2(new_n269), .ZN(new_n284));
  AOI21_X1  g098(.A(new_n193), .B1(new_n267), .B2(KEYINPUT1), .ZN(new_n285));
  XNOR2_X1  g099(.A(new_n284), .B(new_n285), .ZN(new_n286));
  NAND3_X1  g100(.A1(new_n263), .A2(new_n283), .A3(new_n286), .ZN(new_n287));
  AND2_X1   g101(.A1(new_n287), .A2(KEYINPUT30), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n278), .A2(new_n288), .ZN(new_n289));
  NOR2_X1   g103(.A1(KEYINPUT2), .A2(G113), .ZN(new_n290));
  NAND2_X1  g104(.A1(KEYINPUT2), .A2(G113), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n291), .A2(KEYINPUT69), .ZN(new_n292));
  INV_X1    g106(.A(KEYINPUT69), .ZN(new_n293));
  NAND3_X1  g107(.A1(new_n293), .A2(KEYINPUT2), .A3(G113), .ZN(new_n294));
  AOI21_X1  g108(.A(new_n290), .B1(new_n292), .B2(new_n294), .ZN(new_n295));
  XNOR2_X1  g109(.A(G116), .B(G119), .ZN(new_n296));
  NAND2_X1  g110(.A1(new_n295), .A2(new_n296), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n191), .A2(G116), .ZN(new_n298));
  INV_X1    g112(.A(G116), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n299), .A2(G119), .ZN(new_n300));
  NAND2_X1  g114(.A1(new_n298), .A2(new_n300), .ZN(new_n301));
  INV_X1    g115(.A(KEYINPUT70), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n301), .A2(new_n302), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n296), .A2(KEYINPUT70), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n303), .A2(new_n304), .ZN(new_n305));
  OAI21_X1  g119(.A(new_n297), .B1(new_n305), .B2(new_n295), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n289), .A2(new_n306), .ZN(new_n307));
  AOI21_X1  g121(.A(KEYINPUT30), .B1(new_n278), .B2(new_n287), .ZN(new_n308));
  NOR2_X1   g122(.A1(new_n307), .A2(new_n308), .ZN(new_n309));
  INV_X1    g123(.A(new_n306), .ZN(new_n310));
  NAND3_X1  g124(.A1(new_n278), .A2(new_n310), .A3(new_n287), .ZN(new_n311));
  INV_X1    g125(.A(G210), .ZN(new_n312));
  NOR3_X1   g126(.A1(new_n312), .A2(G237), .A3(G953), .ZN(new_n313));
  XNOR2_X1  g127(.A(new_n313), .B(KEYINPUT27), .ZN(new_n314));
  XNOR2_X1  g128(.A(KEYINPUT26), .B(G101), .ZN(new_n315));
  XOR2_X1   g129(.A(new_n314), .B(new_n315), .Z(new_n316));
  NAND2_X1  g130(.A1(new_n311), .A2(new_n316), .ZN(new_n317));
  OAI21_X1  g131(.A(KEYINPUT31), .B1(new_n309), .B2(new_n317), .ZN(new_n318));
  INV_X1    g132(.A(KEYINPUT28), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n311), .A2(new_n319), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n278), .A2(new_n287), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n321), .A2(new_n306), .ZN(new_n322));
  NAND4_X1  g136(.A1(new_n278), .A2(KEYINPUT28), .A3(new_n310), .A4(new_n287), .ZN(new_n323));
  NAND3_X1  g137(.A1(new_n320), .A2(new_n322), .A3(new_n323), .ZN(new_n324));
  INV_X1    g138(.A(new_n316), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n324), .A2(new_n325), .ZN(new_n326));
  INV_X1    g140(.A(KEYINPUT30), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n321), .A2(new_n327), .ZN(new_n328));
  AOI21_X1  g142(.A(new_n310), .B1(new_n278), .B2(new_n288), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n328), .A2(new_n329), .ZN(new_n330));
  XOR2_X1   g144(.A(KEYINPUT71), .B(KEYINPUT31), .Z(new_n331));
  NAND4_X1  g145(.A1(new_n330), .A2(new_n311), .A3(new_n316), .A4(new_n331), .ZN(new_n332));
  NAND3_X1  g146(.A1(new_n318), .A2(new_n326), .A3(new_n332), .ZN(new_n333));
  NOR2_X1   g147(.A1(G472), .A2(G902), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n333), .A2(new_n334), .ZN(new_n335));
  XNOR2_X1  g149(.A(KEYINPUT72), .B(KEYINPUT32), .ZN(new_n336));
  INV_X1    g150(.A(new_n336), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n335), .A2(new_n337), .ZN(new_n338));
  AOI21_X1  g152(.A(new_n310), .B1(new_n278), .B2(new_n287), .ZN(new_n339));
  AND3_X1   g153(.A1(new_n278), .A2(new_n310), .A3(new_n287), .ZN(new_n340));
  AOI21_X1  g154(.A(new_n339), .B1(new_n340), .B2(KEYINPUT73), .ZN(new_n341));
  INV_X1    g155(.A(KEYINPUT73), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n311), .A2(new_n342), .ZN(new_n343));
  AOI21_X1  g157(.A(new_n319), .B1(new_n341), .B2(new_n343), .ZN(new_n344));
  NAND3_X1  g158(.A1(new_n320), .A2(KEYINPUT29), .A3(new_n316), .ZN(new_n345));
  OAI21_X1  g159(.A(new_n234), .B1(new_n344), .B2(new_n345), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n324), .A2(new_n316), .ZN(new_n347));
  NAND3_X1  g161(.A1(new_n330), .A2(new_n311), .A3(new_n325), .ZN(new_n348));
  AOI21_X1  g162(.A(KEYINPUT29), .B1(new_n347), .B2(new_n348), .ZN(new_n349));
  OAI21_X1  g163(.A(G472), .B1(new_n346), .B2(new_n349), .ZN(new_n350));
  NAND3_X1  g164(.A1(new_n333), .A2(KEYINPUT32), .A3(new_n334), .ZN(new_n351));
  NAND3_X1  g165(.A1(new_n338), .A2(new_n350), .A3(new_n351), .ZN(new_n352));
  INV_X1    g166(.A(KEYINPUT74), .ZN(new_n353));
  NAND2_X1  g167(.A1(new_n352), .A2(new_n353), .ZN(new_n354));
  NAND4_X1  g168(.A1(new_n338), .A2(new_n350), .A3(KEYINPUT74), .A4(new_n351), .ZN(new_n355));
  AOI21_X1  g169(.A(new_n247), .B1(new_n354), .B2(new_n355), .ZN(new_n356));
  INV_X1    g170(.A(G221), .ZN(new_n357));
  XNOR2_X1  g171(.A(KEYINPUT9), .B(G234), .ZN(new_n358));
  INV_X1    g172(.A(new_n358), .ZN(new_n359));
  AOI21_X1  g173(.A(new_n357), .B1(new_n359), .B2(new_n234), .ZN(new_n360));
  OR2_X1    g174(.A1(KEYINPUT80), .A2(G107), .ZN(new_n361));
  NAND2_X1  g175(.A1(KEYINPUT80), .A2(G107), .ZN(new_n362));
  AOI21_X1  g176(.A(G104), .B1(new_n361), .B2(new_n362), .ZN(new_n363));
  INV_X1    g177(.A(G104), .ZN(new_n364));
  NOR2_X1   g178(.A1(new_n364), .A2(G107), .ZN(new_n365));
  OAI21_X1  g179(.A(G101), .B1(new_n363), .B2(new_n365), .ZN(new_n366));
  INV_X1    g180(.A(KEYINPUT3), .ZN(new_n367));
  INV_X1    g181(.A(G107), .ZN(new_n368));
  OAI21_X1  g182(.A(new_n367), .B1(new_n368), .B2(G104), .ZN(new_n369));
  OAI21_X1  g183(.A(new_n369), .B1(new_n364), .B2(G107), .ZN(new_n370));
  NAND4_X1  g184(.A1(new_n361), .A2(new_n367), .A3(G104), .A4(new_n362), .ZN(new_n371));
  INV_X1    g185(.A(G101), .ZN(new_n372));
  NAND3_X1  g186(.A1(new_n370), .A2(new_n371), .A3(new_n372), .ZN(new_n373));
  AND2_X1   g187(.A1(new_n366), .A2(new_n373), .ZN(new_n374));
  INV_X1    g188(.A(KEYINPUT10), .ZN(new_n375));
  NAND3_X1  g189(.A1(new_n374), .A2(new_n375), .A3(new_n286), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n366), .A2(new_n373), .ZN(new_n377));
  NOR2_X1   g191(.A1(new_n284), .A2(new_n285), .ZN(new_n378));
  INV_X1    g192(.A(KEYINPUT1), .ZN(new_n379));
  AND4_X1   g193(.A1(new_n379), .A2(new_n267), .A3(new_n269), .A4(G128), .ZN(new_n380));
  NOR2_X1   g194(.A1(new_n378), .A2(new_n380), .ZN(new_n381));
  OAI21_X1  g195(.A(KEYINPUT10), .B1(new_n377), .B2(new_n381), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n376), .A2(new_n382), .ZN(new_n383));
  AOI21_X1  g197(.A(new_n372), .B1(new_n370), .B2(new_n371), .ZN(new_n384));
  INV_X1    g198(.A(KEYINPUT4), .ZN(new_n385));
  AOI22_X1  g199(.A1(new_n275), .A2(new_n274), .B1(new_n384), .B2(new_n385), .ZN(new_n386));
  NAND2_X1  g200(.A1(new_n370), .A2(new_n371), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n387), .A2(G101), .ZN(new_n388));
  NAND3_X1  g202(.A1(new_n388), .A2(KEYINPUT4), .A3(new_n373), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n386), .A2(new_n389), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n383), .A2(new_n390), .ZN(new_n391));
  INV_X1    g205(.A(KEYINPUT83), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n391), .A2(new_n392), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n264), .A2(new_n277), .ZN(new_n394));
  INV_X1    g208(.A(new_n394), .ZN(new_n395));
  AOI22_X1  g209(.A1(new_n376), .A2(new_n382), .B1(new_n389), .B2(new_n386), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n396), .A2(KEYINPUT83), .ZN(new_n397));
  NAND3_X1  g211(.A1(new_n393), .A2(new_n395), .A3(new_n397), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n394), .A2(KEYINPUT81), .ZN(new_n399));
  INV_X1    g213(.A(KEYINPUT81), .ZN(new_n400));
  NAND3_X1  g214(.A1(new_n264), .A2(new_n400), .A3(new_n277), .ZN(new_n401));
  NAND3_X1  g215(.A1(new_n399), .A2(new_n401), .A3(new_n396), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n398), .A2(new_n402), .ZN(new_n403));
  XNOR2_X1  g217(.A(G110), .B(G140), .ZN(new_n404));
  AND2_X1   g218(.A1(new_n226), .A2(G227), .ZN(new_n405));
  XNOR2_X1  g219(.A(new_n404), .B(new_n405), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n403), .A2(new_n406), .ZN(new_n407));
  INV_X1    g221(.A(new_n406), .ZN(new_n408));
  NAND3_X1  g222(.A1(new_n402), .A2(KEYINPUT84), .A3(new_n408), .ZN(new_n409));
  NAND2_X1  g223(.A1(new_n374), .A2(new_n286), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n377), .A2(new_n381), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n410), .A2(new_n411), .ZN(new_n412));
  INV_X1    g226(.A(KEYINPUT82), .ZN(new_n413));
  OAI211_X1 g227(.A(new_n395), .B(new_n412), .C1(new_n413), .C2(KEYINPUT12), .ZN(new_n414));
  NAND3_X1  g228(.A1(new_n412), .A2(new_n264), .A3(new_n277), .ZN(new_n415));
  NAND3_X1  g229(.A1(new_n264), .A2(new_n413), .A3(new_n277), .ZN(new_n416));
  INV_X1    g230(.A(KEYINPUT12), .ZN(new_n417));
  NAND3_X1  g231(.A1(new_n415), .A2(new_n416), .A3(new_n417), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n414), .A2(new_n418), .ZN(new_n419));
  NAND2_X1  g233(.A1(new_n409), .A2(new_n419), .ZN(new_n420));
  AOI21_X1  g234(.A(KEYINPUT84), .B1(new_n402), .B2(new_n408), .ZN(new_n421));
  OAI21_X1  g235(.A(new_n407), .B1(new_n420), .B2(new_n421), .ZN(new_n422));
  INV_X1    g236(.A(G469), .ZN(new_n423));
  NAND3_X1  g237(.A1(new_n422), .A2(new_n423), .A3(new_n234), .ZN(new_n424));
  NOR2_X1   g238(.A1(new_n423), .A2(new_n234), .ZN(new_n425));
  INV_X1    g239(.A(new_n418), .ZN(new_n426));
  AOI21_X1  g240(.A(new_n415), .B1(new_n417), .B2(new_n416), .ZN(new_n427));
  OAI21_X1  g241(.A(new_n402), .B1(new_n426), .B2(new_n427), .ZN(new_n428));
  AOI21_X1  g242(.A(new_n400), .B1(new_n264), .B2(new_n277), .ZN(new_n429));
  NOR2_X1   g243(.A1(new_n391), .A2(new_n429), .ZN(new_n430));
  AOI21_X1  g244(.A(new_n406), .B1(new_n430), .B2(new_n401), .ZN(new_n431));
  AOI22_X1  g245(.A1(new_n428), .A2(new_n406), .B1(new_n431), .B2(new_n398), .ZN(new_n432));
  AOI21_X1  g246(.A(new_n425), .B1(new_n432), .B2(G469), .ZN(new_n433));
  AOI21_X1  g247(.A(new_n360), .B1(new_n424), .B2(new_n433), .ZN(new_n434));
  INV_X1    g248(.A(KEYINPUT85), .ZN(new_n435));
  NOR2_X1   g249(.A1(new_n434), .A2(new_n435), .ZN(new_n436));
  AOI211_X1 g250(.A(KEYINPUT85), .B(new_n360), .C1(new_n424), .C2(new_n433), .ZN(new_n437));
  NAND2_X1  g251(.A1(new_n384), .A2(new_n385), .ZN(new_n438));
  NAND3_X1  g252(.A1(new_n389), .A2(new_n306), .A3(new_n438), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n439), .A2(KEYINPUT86), .ZN(new_n440));
  INV_X1    g254(.A(KEYINPUT86), .ZN(new_n441));
  NAND4_X1  g255(.A1(new_n389), .A2(new_n306), .A3(new_n441), .A4(new_n438), .ZN(new_n442));
  INV_X1    g256(.A(KEYINPUT5), .ZN(new_n443));
  AOI21_X1  g257(.A(new_n443), .B1(new_n303), .B2(new_n304), .ZN(new_n444));
  NAND3_X1  g258(.A1(new_n443), .A2(new_n191), .A3(G116), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n445), .A2(G113), .ZN(new_n446));
  OAI21_X1  g260(.A(new_n297), .B1(new_n444), .B2(new_n446), .ZN(new_n447));
  OR2_X1    g261(.A1(new_n447), .A2(new_n377), .ZN(new_n448));
  NAND3_X1  g262(.A1(new_n440), .A2(new_n442), .A3(new_n448), .ZN(new_n449));
  XNOR2_X1  g263(.A(G110), .B(G122), .ZN(new_n450));
  INV_X1    g264(.A(new_n450), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n449), .A2(new_n451), .ZN(new_n452));
  NAND4_X1  g266(.A1(new_n440), .A2(new_n450), .A3(new_n448), .A4(new_n442), .ZN(new_n453));
  NAND3_X1  g267(.A1(new_n452), .A2(KEYINPUT6), .A3(new_n453), .ZN(new_n454));
  INV_X1    g268(.A(KEYINPUT6), .ZN(new_n455));
  NAND3_X1  g269(.A1(new_n449), .A2(new_n455), .A3(new_n451), .ZN(new_n456));
  OAI21_X1  g270(.A(new_n202), .B1(new_n378), .B2(new_n380), .ZN(new_n457));
  INV_X1    g271(.A(new_n275), .ZN(new_n458));
  OAI21_X1  g272(.A(G125), .B1(new_n458), .B2(new_n273), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n457), .A2(new_n459), .ZN(new_n460));
  NAND2_X1  g274(.A1(new_n226), .A2(G224), .ZN(new_n461));
  XNOR2_X1  g275(.A(new_n460), .B(new_n461), .ZN(new_n462));
  NAND3_X1  g276(.A1(new_n454), .A2(new_n456), .A3(new_n462), .ZN(new_n463));
  XNOR2_X1  g277(.A(new_n450), .B(KEYINPUT8), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n447), .A2(new_n377), .ZN(new_n465));
  INV_X1    g279(.A(KEYINPUT87), .ZN(new_n466));
  OAI211_X1 g280(.A(G113), .B(new_n445), .C1(new_n301), .C2(new_n443), .ZN(new_n467));
  NAND2_X1  g281(.A1(new_n297), .A2(new_n467), .ZN(new_n468));
  OAI21_X1  g282(.A(new_n466), .B1(new_n377), .B2(new_n468), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n465), .A2(new_n469), .ZN(new_n470));
  NOR3_X1   g284(.A1(new_n377), .A2(new_n468), .A3(new_n466), .ZN(new_n471));
  OAI21_X1  g285(.A(new_n464), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  NAND3_X1  g286(.A1(new_n461), .A2(KEYINPUT88), .A3(KEYINPUT7), .ZN(new_n473));
  NAND3_X1  g287(.A1(new_n457), .A2(new_n459), .A3(new_n473), .ZN(new_n474));
  AOI21_X1  g288(.A(KEYINPUT88), .B1(new_n461), .B2(KEYINPUT7), .ZN(new_n475));
  XNOR2_X1  g289(.A(new_n474), .B(new_n475), .ZN(new_n476));
  NAND3_X1  g290(.A1(new_n453), .A2(new_n472), .A3(new_n476), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n477), .A2(new_n234), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n478), .A2(KEYINPUT89), .ZN(new_n479));
  INV_X1    g293(.A(KEYINPUT89), .ZN(new_n480));
  NAND3_X1  g294(.A1(new_n477), .A2(new_n480), .A3(new_n234), .ZN(new_n481));
  NAND3_X1  g295(.A1(new_n463), .A2(new_n479), .A3(new_n481), .ZN(new_n482));
  OAI21_X1  g296(.A(G210), .B1(G237), .B2(G902), .ZN(new_n483));
  INV_X1    g297(.A(new_n483), .ZN(new_n484));
  NAND2_X1  g298(.A1(new_n482), .A2(new_n484), .ZN(new_n485));
  NAND4_X1  g299(.A1(new_n463), .A2(new_n479), .A3(new_n483), .A4(new_n481), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n485), .A2(new_n486), .ZN(new_n487));
  OAI21_X1  g301(.A(G214), .B1(G237), .B2(G902), .ZN(new_n488));
  NAND2_X1  g302(.A1(new_n487), .A2(new_n488), .ZN(new_n489));
  NOR3_X1   g303(.A1(new_n436), .A2(new_n437), .A3(new_n489), .ZN(new_n490));
  XNOR2_X1  g304(.A(G113), .B(G122), .ZN(new_n491));
  XNOR2_X1  g305(.A(KEYINPUT94), .B(G104), .ZN(new_n492));
  XOR2_X1   g306(.A(new_n491), .B(new_n492), .Z(new_n493));
  INV_X1    g307(.A(G237), .ZN(new_n494));
  NAND4_X1  g308(.A1(new_n494), .A2(new_n226), .A3(G143), .A4(G214), .ZN(new_n495));
  XNOR2_X1  g309(.A(new_n495), .B(KEYINPUT91), .ZN(new_n496));
  INV_X1    g310(.A(KEYINPUT90), .ZN(new_n497));
  INV_X1    g311(.A(G214), .ZN(new_n498));
  NOR3_X1   g312(.A1(new_n498), .A2(G237), .A3(G953), .ZN(new_n499));
  OAI21_X1  g313(.A(new_n497), .B1(new_n499), .B2(G143), .ZN(new_n500));
  NAND3_X1  g314(.A1(new_n494), .A2(new_n226), .A3(G214), .ZN(new_n501));
  NAND3_X1  g315(.A1(new_n501), .A2(KEYINPUT90), .A3(new_n268), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n500), .A2(new_n502), .ZN(new_n503));
  AOI21_X1  g317(.A(new_n262), .B1(new_n496), .B2(new_n503), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n504), .A2(KEYINPUT17), .ZN(new_n505));
  NAND3_X1  g319(.A1(new_n505), .A2(new_n215), .A3(new_n209), .ZN(new_n506));
  INV_X1    g320(.A(new_n502), .ZN(new_n507));
  AOI21_X1  g321(.A(KEYINPUT90), .B1(new_n501), .B2(new_n268), .ZN(new_n508));
  NOR2_X1   g322(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  INV_X1    g323(.A(KEYINPUT91), .ZN(new_n510));
  XNOR2_X1  g324(.A(new_n495), .B(new_n510), .ZN(new_n511));
  NOR3_X1   g325(.A1(new_n509), .A2(new_n511), .A3(G131), .ZN(new_n512));
  NOR3_X1   g326(.A1(new_n512), .A2(new_n504), .A3(KEYINPUT17), .ZN(new_n513));
  OR2_X1    g327(.A1(new_n506), .A2(new_n513), .ZN(new_n514));
  NOR2_X1   g328(.A1(new_n509), .A2(new_n511), .ZN(new_n515));
  NAND2_X1  g329(.A1(KEYINPUT18), .A2(G131), .ZN(new_n516));
  AND2_X1   g330(.A1(new_n201), .A2(new_n204), .ZN(new_n517));
  NAND2_X1  g331(.A1(new_n517), .A2(G146), .ZN(new_n518));
  AOI22_X1  g332(.A1(new_n515), .A2(new_n516), .B1(new_n518), .B2(new_n212), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n504), .A2(KEYINPUT18), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  AOI21_X1  g335(.A(new_n493), .B1(new_n514), .B2(new_n521), .ZN(new_n522));
  OAI211_X1 g336(.A(new_n521), .B(new_n493), .C1(new_n513), .C2(new_n506), .ZN(new_n523));
  INV_X1    g337(.A(new_n523), .ZN(new_n524));
  OAI21_X1  g338(.A(new_n234), .B1(new_n522), .B2(new_n524), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n525), .A2(G475), .ZN(new_n526));
  INV_X1    g340(.A(KEYINPUT20), .ZN(new_n527));
  INV_X1    g341(.A(KEYINPUT93), .ZN(new_n528));
  OR2_X1    g342(.A1(new_n528), .A2(KEYINPUT19), .ZN(new_n529));
  NAND2_X1  g343(.A1(new_n528), .A2(KEYINPUT19), .ZN(new_n530));
  NAND3_X1  g344(.A1(new_n210), .A2(new_n529), .A3(new_n530), .ZN(new_n531));
  AOI21_X1  g345(.A(KEYINPUT92), .B1(new_n517), .B2(KEYINPUT19), .ZN(new_n532));
  AND4_X1   g346(.A1(KEYINPUT92), .A2(new_n201), .A3(KEYINPUT19), .A4(new_n204), .ZN(new_n533));
  OAI211_X1 g347(.A(new_n211), .B(new_n531), .C1(new_n532), .C2(new_n533), .ZN(new_n534));
  OAI211_X1 g348(.A(new_n534), .B(new_n209), .C1(new_n504), .C2(new_n512), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n535), .A2(new_n521), .ZN(new_n536));
  INV_X1    g350(.A(new_n493), .ZN(new_n537));
  NAND2_X1  g351(.A1(new_n536), .A2(new_n537), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n538), .A2(new_n523), .ZN(new_n539));
  NOR2_X1   g353(.A1(G475), .A2(G902), .ZN(new_n540));
  AOI21_X1  g354(.A(new_n527), .B1(new_n539), .B2(new_n540), .ZN(new_n541));
  INV_X1    g355(.A(new_n540), .ZN(new_n542));
  AOI211_X1 g356(.A(KEYINPUT20), .B(new_n542), .C1(new_n538), .C2(new_n523), .ZN(new_n543));
  OAI21_X1  g357(.A(new_n526), .B1(new_n541), .B2(new_n543), .ZN(new_n544));
  INV_X1    g358(.A(KEYINPUT96), .ZN(new_n545));
  INV_X1    g359(.A(KEYINPUT95), .ZN(new_n546));
  INV_X1    g360(.A(G122), .ZN(new_n547));
  OAI21_X1  g361(.A(new_n546), .B1(new_n547), .B2(G116), .ZN(new_n548));
  NAND3_X1  g362(.A1(new_n299), .A2(KEYINPUT95), .A3(G122), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n548), .A2(new_n549), .ZN(new_n550));
  OAI21_X1  g364(.A(new_n545), .B1(new_n550), .B2(KEYINPUT14), .ZN(new_n551));
  INV_X1    g365(.A(KEYINPUT14), .ZN(new_n552));
  NAND4_X1  g366(.A1(new_n548), .A2(new_n549), .A3(KEYINPUT96), .A4(new_n552), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n550), .A2(KEYINPUT14), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n547), .A2(G116), .ZN(new_n555));
  NAND4_X1  g369(.A1(new_n551), .A2(new_n553), .A3(new_n554), .A4(new_n555), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n556), .A2(G107), .ZN(new_n557));
  XOR2_X1   g371(.A(G128), .B(G143), .Z(new_n558));
  XNOR2_X1  g372(.A(new_n558), .B(new_n281), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n550), .A2(new_n555), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n361), .A2(new_n362), .ZN(new_n561));
  OR2_X1    g375(.A1(new_n560), .A2(new_n561), .ZN(new_n562));
  NAND3_X1  g376(.A1(new_n557), .A2(new_n559), .A3(new_n562), .ZN(new_n563));
  NAND3_X1  g377(.A1(new_n268), .A2(KEYINPUT13), .A3(G128), .ZN(new_n564));
  OAI21_X1  g378(.A(new_n564), .B1(G128), .B2(new_n268), .ZN(new_n565));
  AOI21_X1  g379(.A(KEYINPUT13), .B1(new_n268), .B2(G128), .ZN(new_n566));
  OAI21_X1  g380(.A(G134), .B1(new_n565), .B2(new_n566), .ZN(new_n567));
  AND2_X1   g381(.A1(new_n560), .A2(new_n561), .ZN(new_n568));
  NOR2_X1   g382(.A1(new_n560), .A2(new_n561), .ZN(new_n569));
  OAI221_X1 g383(.A(new_n567), .B1(new_n281), .B2(new_n558), .C1(new_n568), .C2(new_n569), .ZN(new_n570));
  NOR3_X1   g384(.A1(new_n358), .A2(new_n233), .A3(G953), .ZN(new_n571));
  AND3_X1   g385(.A1(new_n563), .A2(new_n570), .A3(new_n571), .ZN(new_n572));
  AOI21_X1  g386(.A(new_n571), .B1(new_n563), .B2(new_n570), .ZN(new_n573));
  OAI21_X1  g387(.A(new_n234), .B1(new_n572), .B2(new_n573), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n574), .A2(KEYINPUT97), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n563), .A2(new_n570), .ZN(new_n576));
  INV_X1    g390(.A(new_n571), .ZN(new_n577));
  NAND2_X1  g391(.A1(new_n576), .A2(new_n577), .ZN(new_n578));
  NAND3_X1  g392(.A1(new_n563), .A2(new_n570), .A3(new_n571), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  INV_X1    g394(.A(KEYINPUT97), .ZN(new_n581));
  NAND3_X1  g395(.A1(new_n580), .A2(new_n581), .A3(new_n234), .ZN(new_n582));
  INV_X1    g396(.A(G478), .ZN(new_n583));
  NOR2_X1   g397(.A1(new_n583), .A2(KEYINPUT15), .ZN(new_n584));
  NAND3_X1  g398(.A1(new_n575), .A2(new_n582), .A3(new_n584), .ZN(new_n585));
  OR3_X1    g399(.A1(new_n574), .A2(KEYINPUT98), .A3(new_n584), .ZN(new_n586));
  OAI21_X1  g400(.A(KEYINPUT98), .B1(new_n574), .B2(new_n584), .ZN(new_n587));
  NAND3_X1  g401(.A1(new_n585), .A2(new_n586), .A3(new_n587), .ZN(new_n588));
  NOR2_X1   g402(.A1(new_n544), .A2(new_n588), .ZN(new_n589));
  INV_X1    g403(.A(G952), .ZN(new_n590));
  NOR2_X1   g404(.A1(new_n590), .A2(G953), .ZN(new_n591));
  NAND2_X1  g405(.A1(G234), .A2(G237), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  XOR2_X1   g407(.A(KEYINPUT21), .B(G898), .Z(new_n594));
  NAND3_X1  g408(.A1(new_n592), .A2(G902), .A3(G953), .ZN(new_n595));
  OAI21_X1  g409(.A(new_n593), .B1(new_n594), .B2(new_n595), .ZN(new_n596));
  XNOR2_X1  g410(.A(new_n596), .B(KEYINPUT99), .ZN(new_n597));
  AND2_X1   g411(.A1(new_n589), .A2(new_n597), .ZN(new_n598));
  NAND3_X1  g412(.A1(new_n356), .A2(new_n490), .A3(new_n598), .ZN(new_n599));
  XNOR2_X1  g413(.A(new_n599), .B(G101), .ZN(G3));
  NAND2_X1  g414(.A1(new_n333), .A2(new_n234), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n601), .A2(G472), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n602), .A2(new_n335), .ZN(new_n603));
  NOR4_X1   g417(.A1(new_n436), .A2(new_n437), .A3(new_n603), .A4(new_n247), .ZN(new_n604));
  INV_X1    g418(.A(new_n488), .ZN(new_n605));
  INV_X1    g419(.A(new_n486), .ZN(new_n606));
  INV_X1    g420(.A(KEYINPUT100), .ZN(new_n607));
  AOI21_X1  g421(.A(new_n605), .B1(new_n606), .B2(new_n607), .ZN(new_n608));
  NAND3_X1  g422(.A1(new_n485), .A2(new_n486), .A3(KEYINPUT100), .ZN(new_n609));
  NAND2_X1  g423(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  INV_X1    g424(.A(new_n610), .ZN(new_n611));
  AND2_X1   g425(.A1(new_n575), .A2(new_n582), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n612), .A2(new_n583), .ZN(new_n613));
  XNOR2_X1  g427(.A(new_n580), .B(KEYINPUT33), .ZN(new_n614));
  NOR2_X1   g428(.A1(new_n583), .A2(G902), .ZN(new_n615));
  NAND2_X1  g429(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  NAND2_X1  g430(.A1(new_n613), .A2(new_n616), .ZN(new_n617));
  AND3_X1   g431(.A1(new_n617), .A2(new_n597), .A3(new_n544), .ZN(new_n618));
  AND2_X1   g432(.A1(new_n611), .A2(new_n618), .ZN(new_n619));
  NAND2_X1  g433(.A1(new_n604), .A2(new_n619), .ZN(new_n620));
  XNOR2_X1  g434(.A(new_n620), .B(KEYINPUT101), .ZN(new_n621));
  XNOR2_X1  g435(.A(KEYINPUT34), .B(G104), .ZN(new_n622));
  XNOR2_X1  g436(.A(new_n621), .B(new_n622), .ZN(G6));
  NAND3_X1  g437(.A1(new_n539), .A2(new_n527), .A3(new_n540), .ZN(new_n624));
  AOI21_X1  g438(.A(new_n493), .B1(new_n535), .B2(new_n521), .ZN(new_n625));
  OAI21_X1  g439(.A(new_n540), .B1(new_n524), .B2(new_n625), .ZN(new_n626));
  NAND2_X1  g440(.A1(new_n626), .A2(KEYINPUT20), .ZN(new_n627));
  NAND2_X1  g441(.A1(new_n624), .A2(new_n627), .ZN(new_n628));
  NAND4_X1  g442(.A1(new_n588), .A2(new_n628), .A3(new_n597), .A4(new_n526), .ZN(new_n629));
  NOR2_X1   g443(.A1(new_n610), .A2(new_n629), .ZN(new_n630));
  NAND2_X1  g444(.A1(new_n604), .A2(new_n630), .ZN(new_n631));
  XOR2_X1   g445(.A(KEYINPUT35), .B(G107), .Z(new_n632));
  XNOR2_X1  g446(.A(new_n631), .B(new_n632), .ZN(G9));
  NOR2_X1   g447(.A1(new_n229), .A2(KEYINPUT36), .ZN(new_n634));
  XNOR2_X1  g448(.A(new_n224), .B(new_n634), .ZN(new_n635));
  NOR2_X1   g449(.A1(new_n235), .A2(G902), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n635), .A2(new_n636), .ZN(new_n637));
  OAI21_X1  g451(.A(new_n637), .B1(new_n245), .B2(new_n246), .ZN(new_n638));
  NAND2_X1  g452(.A1(new_n598), .A2(new_n638), .ZN(new_n639));
  NOR2_X1   g453(.A1(new_n639), .A2(new_n603), .ZN(new_n640));
  NAND2_X1  g454(.A1(new_n640), .A2(new_n490), .ZN(new_n641));
  XOR2_X1   g455(.A(KEYINPUT37), .B(G110), .Z(new_n642));
  XNOR2_X1  g456(.A(new_n641), .B(new_n642), .ZN(new_n643));
  XNOR2_X1  g457(.A(KEYINPUT102), .B(KEYINPUT103), .ZN(new_n644));
  XNOR2_X1  g458(.A(new_n643), .B(new_n644), .ZN(G12));
  INV_X1    g459(.A(KEYINPUT104), .ZN(new_n646));
  AND3_X1   g460(.A1(new_n333), .A2(KEYINPUT32), .A3(new_n334), .ZN(new_n647));
  AOI21_X1  g461(.A(new_n336), .B1(new_n333), .B2(new_n334), .ZN(new_n648));
  NOR2_X1   g462(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  AOI21_X1  g463(.A(KEYINPUT74), .B1(new_n649), .B2(new_n350), .ZN(new_n650));
  INV_X1    g464(.A(new_n355), .ZN(new_n651));
  OAI21_X1  g465(.A(new_n611), .B1(new_n650), .B2(new_n651), .ZN(new_n652));
  INV_X1    g466(.A(new_n437), .ZN(new_n653));
  OAI21_X1  g467(.A(new_n593), .B1(G900), .B2(new_n595), .ZN(new_n654));
  AND4_X1   g468(.A1(new_n588), .A2(new_n628), .A3(new_n526), .A4(new_n654), .ZN(new_n655));
  NOR2_X1   g469(.A1(new_n242), .A2(new_n244), .ZN(new_n656));
  NAND3_X1  g470(.A1(new_n238), .A2(new_n239), .A3(new_n240), .ZN(new_n657));
  AOI21_X1  g471(.A(new_n246), .B1(new_n656), .B2(new_n657), .ZN(new_n658));
  INV_X1    g472(.A(new_n637), .ZN(new_n659));
  OAI21_X1  g473(.A(new_n655), .B1(new_n658), .B2(new_n659), .ZN(new_n660));
  INV_X1    g474(.A(new_n660), .ZN(new_n661));
  NAND2_X1  g475(.A1(new_n424), .A2(new_n433), .ZN(new_n662));
  INV_X1    g476(.A(new_n360), .ZN(new_n663));
  NAND2_X1  g477(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  NAND2_X1  g478(.A1(new_n664), .A2(KEYINPUT85), .ZN(new_n665));
  NAND3_X1  g479(.A1(new_n653), .A2(new_n661), .A3(new_n665), .ZN(new_n666));
  OAI21_X1  g480(.A(new_n646), .B1(new_n652), .B2(new_n666), .ZN(new_n667));
  AOI21_X1  g481(.A(new_n610), .B1(new_n354), .B2(new_n355), .ZN(new_n668));
  NOR3_X1   g482(.A1(new_n436), .A2(new_n437), .A3(new_n660), .ZN(new_n669));
  NAND3_X1  g483(.A1(new_n668), .A2(new_n669), .A3(KEYINPUT104), .ZN(new_n670));
  NAND2_X1  g484(.A1(new_n667), .A2(new_n670), .ZN(new_n671));
  XNOR2_X1  g485(.A(new_n671), .B(G128), .ZN(G30));
  NOR2_X1   g486(.A1(new_n436), .A2(new_n437), .ZN(new_n673));
  XNOR2_X1  g487(.A(new_n654), .B(KEYINPUT39), .ZN(new_n674));
  NAND2_X1  g488(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  OR2_X1    g489(.A1(new_n675), .A2(KEYINPUT40), .ZN(new_n676));
  NAND2_X1  g490(.A1(new_n675), .A2(KEYINPUT40), .ZN(new_n677));
  XOR2_X1   g491(.A(new_n487), .B(KEYINPUT38), .Z(new_n678));
  OAI21_X1  g492(.A(new_n316), .B1(new_n309), .B2(new_n340), .ZN(new_n679));
  NAND2_X1  g493(.A1(new_n341), .A2(new_n343), .ZN(new_n680));
  OAI211_X1 g494(.A(new_n679), .B(new_n234), .C1(new_n316), .C2(new_n680), .ZN(new_n681));
  AND2_X1   g495(.A1(new_n681), .A2(G472), .ZN(new_n682));
  NOR3_X1   g496(.A1(new_n682), .A2(new_n647), .A3(new_n648), .ZN(new_n683));
  NAND2_X1  g497(.A1(new_n238), .A2(new_n240), .ZN(new_n684));
  NAND2_X1  g498(.A1(new_n684), .A2(KEYINPUT79), .ZN(new_n685));
  OR2_X1    g499(.A1(new_n238), .A2(new_n243), .ZN(new_n686));
  NAND3_X1  g500(.A1(new_n685), .A2(new_n657), .A3(new_n686), .ZN(new_n687));
  AOI21_X1  g501(.A(new_n659), .B1(new_n687), .B2(new_n235), .ZN(new_n688));
  AND2_X1   g502(.A1(new_n544), .A2(new_n588), .ZN(new_n689));
  NAND3_X1  g503(.A1(new_n688), .A2(new_n689), .A3(new_n488), .ZN(new_n690));
  NOR3_X1   g504(.A1(new_n678), .A2(new_n683), .A3(new_n690), .ZN(new_n691));
  NAND3_X1  g505(.A1(new_n676), .A2(new_n677), .A3(new_n691), .ZN(new_n692));
  XOR2_X1   g506(.A(KEYINPUT105), .B(G143), .Z(new_n693));
  XNOR2_X1  g507(.A(new_n692), .B(new_n693), .ZN(G45));
  NOR3_X1   g508(.A1(new_n436), .A2(new_n437), .A3(new_n688), .ZN(new_n695));
  NAND3_X1  g509(.A1(new_n617), .A2(new_n544), .A3(new_n654), .ZN(new_n696));
  XNOR2_X1  g510(.A(new_n696), .B(KEYINPUT106), .ZN(new_n697));
  INV_X1    g511(.A(new_n697), .ZN(new_n698));
  NAND3_X1  g512(.A1(new_n668), .A2(new_n695), .A3(new_n698), .ZN(new_n699));
  XNOR2_X1  g513(.A(new_n699), .B(G146), .ZN(G48));
  NAND2_X1  g514(.A1(new_n422), .A2(new_n234), .ZN(new_n701));
  NAND2_X1  g515(.A1(new_n701), .A2(G469), .ZN(new_n702));
  NAND2_X1  g516(.A1(new_n702), .A2(new_n424), .ZN(new_n703));
  NOR2_X1   g517(.A1(new_n703), .A2(new_n360), .ZN(new_n704));
  NAND3_X1  g518(.A1(new_n356), .A2(new_n619), .A3(new_n704), .ZN(new_n705));
  NAND2_X1  g519(.A1(new_n705), .A2(KEYINPUT107), .ZN(new_n706));
  INV_X1    g520(.A(KEYINPUT107), .ZN(new_n707));
  NAND4_X1  g521(.A1(new_n356), .A2(new_n619), .A3(new_n707), .A4(new_n704), .ZN(new_n708));
  NAND2_X1  g522(.A1(new_n706), .A2(new_n708), .ZN(new_n709));
  XNOR2_X1  g523(.A(KEYINPUT41), .B(G113), .ZN(new_n710));
  XNOR2_X1  g524(.A(new_n709), .B(new_n710), .ZN(G15));
  NAND2_X1  g525(.A1(new_n354), .A2(new_n355), .ZN(new_n712));
  AOI21_X1  g526(.A(new_n236), .B1(new_n687), .B2(new_n235), .ZN(new_n713));
  NAND4_X1  g527(.A1(new_n712), .A2(new_n713), .A3(new_n630), .A4(new_n704), .ZN(new_n714));
  XNOR2_X1  g528(.A(new_n714), .B(G116), .ZN(G18));
  INV_X1    g529(.A(new_n639), .ZN(new_n716));
  NAND4_X1  g530(.A1(new_n712), .A2(new_n716), .A3(new_n611), .A4(new_n704), .ZN(new_n717));
  XNOR2_X1  g531(.A(new_n717), .B(G119), .ZN(G21));
  XNOR2_X1  g532(.A(new_n713), .B(KEYINPUT109), .ZN(new_n719));
  NAND2_X1  g533(.A1(new_n680), .A2(KEYINPUT28), .ZN(new_n720));
  AOI21_X1  g534(.A(new_n316), .B1(new_n720), .B2(new_n320), .ZN(new_n721));
  NAND2_X1  g535(.A1(new_n318), .A2(new_n332), .ZN(new_n722));
  OAI21_X1  g536(.A(new_n334), .B1(new_n721), .B2(new_n722), .ZN(new_n723));
  INV_X1    g537(.A(new_n723), .ZN(new_n724));
  NAND2_X1  g538(.A1(new_n602), .A2(KEYINPUT108), .ZN(new_n725));
  INV_X1    g539(.A(KEYINPUT108), .ZN(new_n726));
  NAND3_X1  g540(.A1(new_n601), .A2(new_n726), .A3(G472), .ZN(new_n727));
  AOI21_X1  g541(.A(new_n724), .B1(new_n725), .B2(new_n727), .ZN(new_n728));
  NAND3_X1  g542(.A1(new_n608), .A2(new_n689), .A3(new_n609), .ZN(new_n729));
  NAND4_X1  g543(.A1(new_n702), .A2(new_n663), .A3(new_n424), .A4(new_n597), .ZN(new_n730));
  NOR2_X1   g544(.A1(new_n729), .A2(new_n730), .ZN(new_n731));
  NAND3_X1  g545(.A1(new_n719), .A2(new_n728), .A3(new_n731), .ZN(new_n732));
  XNOR2_X1  g546(.A(new_n732), .B(G122), .ZN(G24));
  NAND2_X1  g547(.A1(new_n725), .A2(new_n727), .ZN(new_n734));
  INV_X1    g548(.A(KEYINPUT110), .ZN(new_n735));
  NAND4_X1  g549(.A1(new_n734), .A2(new_n735), .A3(new_n638), .A4(new_n723), .ZN(new_n736));
  AOI21_X1  g550(.A(new_n726), .B1(new_n601), .B2(G472), .ZN(new_n737));
  INV_X1    g551(.A(G472), .ZN(new_n738));
  AOI211_X1 g552(.A(KEYINPUT108), .B(new_n738), .C1(new_n333), .C2(new_n234), .ZN(new_n739));
  OAI211_X1 g553(.A(new_n638), .B(new_n723), .C1(new_n737), .C2(new_n739), .ZN(new_n740));
  NAND2_X1  g554(.A1(new_n740), .A2(KEYINPUT110), .ZN(new_n741));
  NAND2_X1  g555(.A1(new_n736), .A2(new_n741), .ZN(new_n742));
  NOR3_X1   g556(.A1(new_n610), .A2(new_n703), .A3(new_n360), .ZN(new_n743));
  NAND3_X1  g557(.A1(new_n742), .A2(new_n698), .A3(new_n743), .ZN(new_n744));
  XNOR2_X1  g558(.A(new_n744), .B(G125), .ZN(G27));
  NOR2_X1   g559(.A1(new_n487), .A2(new_n605), .ZN(new_n746));
  AND2_X1   g560(.A1(new_n746), .A2(new_n434), .ZN(new_n747));
  NAND3_X1  g561(.A1(new_n356), .A2(new_n698), .A3(new_n747), .ZN(new_n748));
  INV_X1    g562(.A(KEYINPUT42), .ZN(new_n749));
  NAND2_X1  g563(.A1(new_n748), .A2(new_n749), .ZN(new_n750));
  INV_X1    g564(.A(KEYINPUT32), .ZN(new_n751));
  NAND2_X1  g565(.A1(new_n335), .A2(new_n751), .ZN(new_n752));
  NAND3_X1  g566(.A1(new_n752), .A2(new_n350), .A3(new_n351), .ZN(new_n753));
  AND2_X1   g567(.A1(new_n719), .A2(new_n753), .ZN(new_n754));
  NAND4_X1  g568(.A1(new_n754), .A2(KEYINPUT42), .A3(new_n698), .A4(new_n747), .ZN(new_n755));
  NAND2_X1  g569(.A1(new_n750), .A2(new_n755), .ZN(new_n756));
  XNOR2_X1  g570(.A(new_n756), .B(G131), .ZN(G33));
  NAND3_X1  g571(.A1(new_n356), .A2(new_n655), .A3(new_n747), .ZN(new_n758));
  NAND2_X1  g572(.A1(new_n758), .A2(KEYINPUT111), .ZN(new_n759));
  INV_X1    g573(.A(KEYINPUT111), .ZN(new_n760));
  NAND4_X1  g574(.A1(new_n356), .A2(new_n760), .A3(new_n655), .A4(new_n747), .ZN(new_n761));
  NAND2_X1  g575(.A1(new_n759), .A2(new_n761), .ZN(new_n762));
  XNOR2_X1  g576(.A(new_n762), .B(G134), .ZN(G36));
  NAND2_X1  g577(.A1(new_n432), .A2(KEYINPUT45), .ZN(new_n764));
  INV_X1    g578(.A(new_n764), .ZN(new_n765));
  OAI21_X1  g579(.A(G469), .B1(new_n432), .B2(KEYINPUT45), .ZN(new_n766));
  NOR2_X1   g580(.A1(new_n765), .A2(new_n766), .ZN(new_n767));
  NOR2_X1   g581(.A1(new_n767), .A2(new_n425), .ZN(new_n768));
  AND2_X1   g582(.A1(new_n768), .A2(KEYINPUT46), .ZN(new_n769));
  OAI21_X1  g583(.A(new_n424), .B1(new_n768), .B2(KEYINPUT46), .ZN(new_n770));
  OAI21_X1  g584(.A(new_n663), .B1(new_n769), .B2(new_n770), .ZN(new_n771));
  INV_X1    g585(.A(new_n674), .ZN(new_n772));
  NOR2_X1   g586(.A1(new_n771), .A2(new_n772), .ZN(new_n773));
  AOI22_X1  g587(.A1(new_n612), .A2(new_n583), .B1(new_n614), .B2(new_n615), .ZN(new_n774));
  NOR2_X1   g588(.A1(new_n774), .A2(new_n544), .ZN(new_n775));
  XNOR2_X1  g589(.A(new_n775), .B(KEYINPUT43), .ZN(new_n776));
  NAND3_X1  g590(.A1(new_n776), .A2(new_n603), .A3(new_n638), .ZN(new_n777));
  INV_X1    g591(.A(KEYINPUT44), .ZN(new_n778));
  OR2_X1    g592(.A1(new_n777), .A2(new_n778), .ZN(new_n779));
  NAND2_X1  g593(.A1(new_n777), .A2(new_n778), .ZN(new_n780));
  NAND4_X1  g594(.A1(new_n773), .A2(new_n746), .A3(new_n779), .A4(new_n780), .ZN(new_n781));
  XOR2_X1   g595(.A(KEYINPUT112), .B(G137), .Z(new_n782));
  XNOR2_X1  g596(.A(new_n781), .B(new_n782), .ZN(G39));
  NOR2_X1   g597(.A1(new_n650), .A2(new_n651), .ZN(new_n784));
  NAND4_X1  g598(.A1(new_n784), .A2(new_n698), .A3(new_n247), .A4(new_n746), .ZN(new_n785));
  INV_X1    g599(.A(KEYINPUT113), .ZN(new_n786));
  XNOR2_X1  g600(.A(new_n785), .B(new_n786), .ZN(new_n787));
  INV_X1    g601(.A(KEYINPUT47), .ZN(new_n788));
  XNOR2_X1  g602(.A(new_n771), .B(new_n788), .ZN(new_n789));
  NAND2_X1  g603(.A1(new_n787), .A2(new_n789), .ZN(new_n790));
  XNOR2_X1  g604(.A(new_n790), .B(G140), .ZN(G42));
  NAND3_X1  g605(.A1(new_n719), .A2(new_n488), .A3(new_n663), .ZN(new_n792));
  XNOR2_X1  g606(.A(new_n792), .B(KEYINPUT114), .ZN(new_n793));
  NOR2_X1   g607(.A1(new_n703), .A2(KEYINPUT49), .ZN(new_n794));
  XNOR2_X1  g608(.A(new_n794), .B(KEYINPUT115), .ZN(new_n795));
  NAND3_X1  g609(.A1(new_n678), .A2(new_n683), .A3(new_n775), .ZN(new_n796));
  AOI21_X1  g610(.A(new_n796), .B1(KEYINPUT49), .B2(new_n703), .ZN(new_n797));
  NAND3_X1  g611(.A1(new_n793), .A2(new_n795), .A3(new_n797), .ZN(new_n798));
  AOI21_X1  g612(.A(new_n697), .B1(new_n736), .B2(new_n741), .ZN(new_n799));
  NAND2_X1  g613(.A1(new_n799), .A2(new_n747), .ZN(new_n800));
  INV_X1    g614(.A(KEYINPUT116), .ZN(new_n801));
  OAI21_X1  g615(.A(new_n801), .B1(new_n489), .B2(new_n629), .ZN(new_n802));
  INV_X1    g616(.A(new_n629), .ZN(new_n803));
  NAND4_X1  g617(.A1(new_n803), .A2(KEYINPUT116), .A3(new_n487), .A4(new_n488), .ZN(new_n804));
  NAND3_X1  g618(.A1(new_n618), .A2(new_n488), .A3(new_n487), .ZN(new_n805));
  NAND3_X1  g619(.A1(new_n802), .A2(new_n804), .A3(new_n805), .ZN(new_n806));
  AOI22_X1  g620(.A1(new_n604), .A2(new_n806), .B1(new_n640), .B2(new_n490), .ZN(new_n807));
  AND3_X1   g621(.A1(new_n746), .A2(new_n589), .A3(new_n654), .ZN(new_n808));
  NAND3_X1  g622(.A1(new_n695), .A2(new_n712), .A3(new_n808), .ZN(new_n809));
  AND4_X1   g623(.A1(new_n599), .A2(new_n800), .A3(new_n807), .A4(new_n809), .ZN(new_n810));
  NAND3_X1  g624(.A1(new_n717), .A2(new_n714), .A3(new_n732), .ZN(new_n811));
  AOI21_X1  g625(.A(new_n811), .B1(new_n708), .B2(new_n706), .ZN(new_n812));
  AOI22_X1  g626(.A1(new_n750), .A2(new_n755), .B1(new_n759), .B2(new_n761), .ZN(new_n813));
  AND3_X1   g627(.A1(new_n810), .A2(new_n812), .A3(new_n813), .ZN(new_n814));
  INV_X1    g628(.A(KEYINPUT52), .ZN(new_n815));
  NOR2_X1   g629(.A1(new_n683), .A2(new_n729), .ZN(new_n816));
  NAND2_X1  g630(.A1(new_n688), .A2(new_n654), .ZN(new_n817));
  OAI21_X1  g631(.A(KEYINPUT118), .B1(new_n817), .B2(new_n664), .ZN(new_n818));
  INV_X1    g632(.A(KEYINPUT118), .ZN(new_n819));
  NAND4_X1  g633(.A1(new_n434), .A2(new_n688), .A3(new_n819), .A4(new_n654), .ZN(new_n820));
  NAND3_X1  g634(.A1(new_n816), .A2(new_n818), .A3(new_n820), .ZN(new_n821));
  INV_X1    g635(.A(KEYINPUT119), .ZN(new_n822));
  NAND2_X1  g636(.A1(new_n821), .A2(new_n822), .ZN(new_n823));
  NAND4_X1  g637(.A1(new_n816), .A2(new_n818), .A3(KEYINPUT119), .A4(new_n820), .ZN(new_n824));
  NAND2_X1  g638(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  NAND2_X1  g639(.A1(new_n825), .A2(new_n699), .ZN(new_n826));
  AND3_X1   g640(.A1(new_n668), .A2(KEYINPUT104), .A3(new_n669), .ZN(new_n827));
  AOI21_X1  g641(.A(KEYINPUT104), .B1(new_n668), .B2(new_n669), .ZN(new_n828));
  OAI21_X1  g642(.A(new_n744), .B1(new_n827), .B2(new_n828), .ZN(new_n829));
  OAI21_X1  g643(.A(new_n815), .B1(new_n826), .B2(new_n829), .ZN(new_n830));
  AOI22_X1  g644(.A1(new_n667), .A2(new_n670), .B1(new_n799), .B2(new_n743), .ZN(new_n831));
  NAND4_X1  g645(.A1(new_n831), .A2(KEYINPUT52), .A3(new_n699), .A4(new_n825), .ZN(new_n832));
  NAND2_X1  g646(.A1(new_n830), .A2(new_n832), .ZN(new_n833));
  NAND2_X1  g647(.A1(new_n814), .A2(new_n833), .ZN(new_n834));
  NAND2_X1  g648(.A1(new_n834), .A2(KEYINPUT53), .ZN(new_n835));
  INV_X1    g649(.A(KEYINPUT53), .ZN(new_n836));
  NOR2_X1   g650(.A1(new_n652), .A2(new_n697), .ZN(new_n837));
  AOI22_X1  g651(.A1(new_n823), .A2(new_n824), .B1(new_n837), .B2(new_n695), .ZN(new_n838));
  AOI21_X1  g652(.A(KEYINPUT52), .B1(new_n838), .B2(new_n831), .ZN(new_n839));
  NAND3_X1  g653(.A1(new_n825), .A2(KEYINPUT52), .A3(new_n699), .ZN(new_n840));
  NAND2_X1  g654(.A1(new_n829), .A2(KEYINPUT117), .ZN(new_n841));
  INV_X1    g655(.A(KEYINPUT117), .ZN(new_n842));
  OAI211_X1 g656(.A(new_n744), .B(new_n842), .C1(new_n827), .C2(new_n828), .ZN(new_n843));
  AOI21_X1  g657(.A(new_n840), .B1(new_n841), .B2(new_n843), .ZN(new_n844));
  OAI211_X1 g658(.A(new_n814), .B(new_n836), .C1(new_n839), .C2(new_n844), .ZN(new_n845));
  AND3_X1   g659(.A1(new_n835), .A2(new_n845), .A3(KEYINPUT54), .ZN(new_n846));
  NAND2_X1  g660(.A1(new_n841), .A2(new_n843), .ZN(new_n847));
  INV_X1    g661(.A(new_n840), .ZN(new_n848));
  AOI21_X1  g662(.A(new_n839), .B1(new_n847), .B2(new_n848), .ZN(new_n849));
  NAND3_X1  g663(.A1(new_n810), .A2(new_n813), .A3(new_n812), .ZN(new_n850));
  OAI21_X1  g664(.A(KEYINPUT53), .B1(new_n849), .B2(new_n850), .ZN(new_n851));
  NAND3_X1  g665(.A1(new_n814), .A2(new_n836), .A3(new_n833), .ZN(new_n852));
  AOI21_X1  g666(.A(KEYINPUT54), .B1(new_n851), .B2(new_n852), .ZN(new_n853));
  NOR2_X1   g667(.A1(new_n846), .A2(new_n853), .ZN(new_n854));
  AND2_X1   g668(.A1(new_n719), .A2(new_n728), .ZN(new_n855));
  INV_X1    g669(.A(new_n593), .ZN(new_n856));
  AND2_X1   g670(.A1(new_n776), .A2(new_n856), .ZN(new_n857));
  NAND2_X1  g671(.A1(new_n855), .A2(new_n857), .ZN(new_n858));
  NAND3_X1  g672(.A1(new_n678), .A2(new_n605), .A3(new_n704), .ZN(new_n859));
  NOR2_X1   g673(.A1(new_n858), .A2(new_n859), .ZN(new_n860));
  XNOR2_X1  g674(.A(new_n860), .B(KEYINPUT50), .ZN(new_n861));
  INV_X1    g675(.A(new_n858), .ZN(new_n862));
  NOR2_X1   g676(.A1(new_n703), .A2(new_n663), .ZN(new_n863));
  OAI211_X1 g677(.A(new_n746), .B(new_n862), .C1(new_n789), .C2(new_n863), .ZN(new_n864));
  AND2_X1   g678(.A1(new_n704), .A2(new_n746), .ZN(new_n865));
  NAND4_X1  g679(.A1(new_n865), .A2(new_n713), .A3(new_n856), .A4(new_n683), .ZN(new_n866));
  NOR3_X1   g680(.A1(new_n866), .A2(new_n544), .A3(new_n617), .ZN(new_n867));
  NAND2_X1  g681(.A1(new_n857), .A2(new_n865), .ZN(new_n868));
  INV_X1    g682(.A(KEYINPUT120), .ZN(new_n869));
  NAND2_X1  g683(.A1(new_n868), .A2(new_n869), .ZN(new_n870));
  NAND3_X1  g684(.A1(new_n857), .A2(KEYINPUT120), .A3(new_n865), .ZN(new_n871));
  NAND2_X1  g685(.A1(new_n870), .A2(new_n871), .ZN(new_n872));
  AOI21_X1  g686(.A(new_n867), .B1(new_n872), .B2(new_n742), .ZN(new_n873));
  NAND3_X1  g687(.A1(new_n861), .A2(new_n864), .A3(new_n873), .ZN(new_n874));
  INV_X1    g688(.A(KEYINPUT51), .ZN(new_n875));
  NAND2_X1  g689(.A1(new_n874), .A2(new_n875), .ZN(new_n876));
  NAND2_X1  g690(.A1(new_n617), .A2(new_n544), .ZN(new_n877));
  INV_X1    g691(.A(new_n743), .ZN(new_n878));
  OAI221_X1 g692(.A(new_n591), .B1(new_n866), .B2(new_n877), .C1(new_n858), .C2(new_n878), .ZN(new_n879));
  NAND2_X1  g693(.A1(new_n872), .A2(new_n754), .ZN(new_n880));
  OR2_X1    g694(.A1(new_n880), .A2(KEYINPUT48), .ZN(new_n881));
  NAND2_X1  g695(.A1(new_n880), .A2(KEYINPUT48), .ZN(new_n882));
  AOI21_X1  g696(.A(new_n879), .B1(new_n881), .B2(new_n882), .ZN(new_n883));
  NAND4_X1  g697(.A1(new_n861), .A2(new_n864), .A3(KEYINPUT51), .A4(new_n873), .ZN(new_n884));
  AND3_X1   g698(.A1(new_n876), .A2(new_n883), .A3(new_n884), .ZN(new_n885));
  AOI21_X1  g699(.A(KEYINPUT121), .B1(new_n854), .B2(new_n885), .ZN(new_n886));
  INV_X1    g700(.A(new_n843), .ZN(new_n887));
  AOI21_X1  g701(.A(new_n842), .B1(new_n671), .B2(new_n744), .ZN(new_n888));
  OAI21_X1  g702(.A(new_n848), .B1(new_n887), .B2(new_n888), .ZN(new_n889));
  AOI21_X1  g703(.A(new_n850), .B1(new_n889), .B2(new_n830), .ZN(new_n890));
  OAI21_X1  g704(.A(new_n852), .B1(new_n890), .B2(new_n836), .ZN(new_n891));
  INV_X1    g705(.A(KEYINPUT54), .ZN(new_n892));
  NAND2_X1  g706(.A1(new_n891), .A2(new_n892), .ZN(new_n893));
  NAND3_X1  g707(.A1(new_n835), .A2(new_n845), .A3(KEYINPUT54), .ZN(new_n894));
  NAND4_X1  g708(.A1(new_n893), .A2(KEYINPUT121), .A3(new_n885), .A4(new_n894), .ZN(new_n895));
  NAND2_X1  g709(.A1(new_n590), .A2(new_n226), .ZN(new_n896));
  NAND2_X1  g710(.A1(new_n895), .A2(new_n896), .ZN(new_n897));
  OAI21_X1  g711(.A(new_n798), .B1(new_n886), .B2(new_n897), .ZN(G75));
  NOR2_X1   g712(.A1(new_n226), .A2(G952), .ZN(new_n899));
  INV_X1    g713(.A(new_n899), .ZN(new_n900));
  OAI211_X1 g714(.A(G902), .B(new_n852), .C1(new_n890), .C2(new_n836), .ZN(new_n901));
  NOR2_X1   g715(.A1(new_n901), .A2(new_n312), .ZN(new_n902));
  NAND2_X1  g716(.A1(new_n454), .A2(new_n456), .ZN(new_n903));
  XNOR2_X1  g717(.A(new_n903), .B(new_n462), .ZN(new_n904));
  XOR2_X1   g718(.A(new_n904), .B(KEYINPUT55), .Z(new_n905));
  OR2_X1    g719(.A1(new_n905), .A2(KEYINPUT56), .ZN(new_n906));
  OAI21_X1  g720(.A(new_n900), .B1(new_n902), .B2(new_n906), .ZN(new_n907));
  OR3_X1    g721(.A1(new_n901), .A2(KEYINPUT122), .A3(new_n312), .ZN(new_n908));
  INV_X1    g722(.A(KEYINPUT56), .ZN(new_n909));
  OAI21_X1  g723(.A(KEYINPUT122), .B1(new_n901), .B2(new_n312), .ZN(new_n910));
  NAND3_X1  g724(.A1(new_n908), .A2(new_n909), .A3(new_n910), .ZN(new_n911));
  AOI21_X1  g725(.A(new_n907), .B1(new_n911), .B2(new_n905), .ZN(G51));
  XNOR2_X1  g726(.A(new_n425), .B(KEYINPUT57), .ZN(new_n913));
  NAND3_X1  g727(.A1(new_n851), .A2(KEYINPUT54), .A3(new_n852), .ZN(new_n914));
  INV_X1    g728(.A(new_n914), .ZN(new_n915));
  OAI21_X1  g729(.A(new_n913), .B1(new_n915), .B2(new_n853), .ZN(new_n916));
  NAND2_X1  g730(.A1(new_n916), .A2(new_n422), .ZN(new_n917));
  NAND4_X1  g731(.A1(new_n851), .A2(G902), .A3(new_n767), .A4(new_n852), .ZN(new_n918));
  AOI21_X1  g732(.A(new_n899), .B1(new_n917), .B2(new_n918), .ZN(G54));
  INV_X1    g733(.A(new_n539), .ZN(new_n920));
  NAND2_X1  g734(.A1(KEYINPUT58), .A2(G475), .ZN(new_n921));
  OAI21_X1  g735(.A(new_n920), .B1(new_n901), .B2(new_n921), .ZN(new_n922));
  NAND2_X1  g736(.A1(new_n922), .A2(new_n900), .ZN(new_n923));
  NOR3_X1   g737(.A1(new_n901), .A2(new_n920), .A3(new_n921), .ZN(new_n924));
  NOR2_X1   g738(.A1(new_n923), .A2(new_n924), .ZN(G60));
  NOR2_X1   g739(.A1(new_n915), .A2(new_n853), .ZN(new_n926));
  NAND2_X1  g740(.A1(G478), .A2(G902), .ZN(new_n927));
  XNOR2_X1  g741(.A(new_n927), .B(KEYINPUT59), .ZN(new_n928));
  NAND2_X1  g742(.A1(new_n614), .A2(new_n928), .ZN(new_n929));
  OAI21_X1  g743(.A(new_n900), .B1(new_n926), .B2(new_n929), .ZN(new_n930));
  NAND2_X1  g744(.A1(new_n893), .A2(new_n894), .ZN(new_n931));
  AOI21_X1  g745(.A(new_n614), .B1(new_n931), .B2(new_n928), .ZN(new_n932));
  NOR2_X1   g746(.A1(new_n930), .A2(new_n932), .ZN(G63));
  NAND2_X1  g747(.A1(G217), .A2(G902), .ZN(new_n934));
  XOR2_X1   g748(.A(new_n934), .B(KEYINPUT60), .Z(new_n935));
  OAI211_X1 g749(.A(new_n852), .B(new_n935), .C1(new_n890), .C2(new_n836), .ZN(new_n936));
  NAND2_X1  g750(.A1(new_n936), .A2(new_n232), .ZN(new_n937));
  NAND4_X1  g751(.A1(new_n851), .A2(new_n635), .A3(new_n852), .A4(new_n935), .ZN(new_n938));
  NAND3_X1  g752(.A1(new_n937), .A2(new_n900), .A3(new_n938), .ZN(new_n939));
  INV_X1    g753(.A(KEYINPUT61), .ZN(new_n940));
  OR2_X1    g754(.A1(new_n940), .A2(KEYINPUT123), .ZN(new_n941));
  NAND2_X1  g755(.A1(new_n940), .A2(KEYINPUT123), .ZN(new_n942));
  NAND3_X1  g756(.A1(new_n939), .A2(new_n941), .A3(new_n942), .ZN(new_n943));
  AOI21_X1  g757(.A(new_n899), .B1(new_n936), .B2(new_n232), .ZN(new_n944));
  NAND4_X1  g758(.A1(new_n944), .A2(KEYINPUT123), .A3(new_n940), .A4(new_n938), .ZN(new_n945));
  AND2_X1   g759(.A1(new_n943), .A2(new_n945), .ZN(G66));
  NAND3_X1  g760(.A1(new_n594), .A2(G224), .A3(G953), .ZN(new_n947));
  NAND3_X1  g761(.A1(new_n812), .A2(new_n599), .A3(new_n807), .ZN(new_n948));
  OAI21_X1  g762(.A(new_n947), .B1(new_n948), .B2(G953), .ZN(new_n949));
  OAI21_X1  g763(.A(new_n903), .B1(G898), .B2(new_n226), .ZN(new_n950));
  XOR2_X1   g764(.A(new_n949), .B(new_n950), .Z(G69));
  AOI21_X1  g765(.A(new_n226), .B1(G227), .B2(G900), .ZN(new_n952));
  INV_X1    g766(.A(new_n952), .ZN(new_n953));
  AND3_X1   g767(.A1(new_n779), .A2(new_n746), .A3(new_n780), .ZN(new_n954));
  AND3_X1   g768(.A1(new_n754), .A2(new_n611), .A3(new_n689), .ZN(new_n955));
  OAI21_X1  g769(.A(new_n773), .B1(new_n954), .B2(new_n955), .ZN(new_n956));
  AND4_X1   g770(.A1(new_n756), .A2(new_n956), .A3(new_n790), .A4(new_n762), .ZN(new_n957));
  AND2_X1   g771(.A1(new_n847), .A2(new_n699), .ZN(new_n958));
  NAND3_X1  g772(.A1(new_n957), .A2(new_n226), .A3(new_n958), .ZN(new_n959));
  NAND2_X1  g773(.A1(new_n328), .A2(new_n289), .ZN(new_n960));
  OAI21_X1  g774(.A(new_n531), .B1(new_n532), .B2(new_n533), .ZN(new_n961));
  XNOR2_X1  g775(.A(new_n960), .B(new_n961), .ZN(new_n962));
  INV_X1    g776(.A(new_n962), .ZN(new_n963));
  AOI21_X1  g777(.A(new_n963), .B1(G900), .B2(G953), .ZN(new_n964));
  NAND2_X1  g778(.A1(new_n959), .A2(new_n964), .ZN(new_n965));
  NAND3_X1  g779(.A1(new_n847), .A2(new_n692), .A3(new_n699), .ZN(new_n966));
  OR2_X1    g780(.A1(new_n966), .A2(KEYINPUT62), .ZN(new_n967));
  NAND2_X1  g781(.A1(new_n966), .A2(KEYINPUT62), .ZN(new_n968));
  NAND3_X1  g782(.A1(new_n588), .A2(new_n628), .A3(new_n526), .ZN(new_n969));
  AND2_X1   g783(.A1(new_n877), .A2(new_n969), .ZN(new_n970));
  INV_X1    g784(.A(KEYINPUT125), .ZN(new_n971));
  OAI21_X1  g785(.A(new_n746), .B1(new_n970), .B2(new_n971), .ZN(new_n972));
  AOI21_X1  g786(.A(new_n972), .B1(new_n971), .B2(new_n970), .ZN(new_n973));
  NAND4_X1  g787(.A1(new_n973), .A2(new_n673), .A3(new_n356), .A4(new_n674), .ZN(new_n974));
  NAND2_X1  g788(.A1(new_n781), .A2(new_n974), .ZN(new_n975));
  XOR2_X1   g789(.A(new_n975), .B(KEYINPUT126), .Z(new_n976));
  NAND4_X1  g790(.A1(new_n967), .A2(new_n790), .A3(new_n968), .A4(new_n976), .ZN(new_n977));
  AND2_X1   g791(.A1(new_n977), .A2(new_n226), .ZN(new_n978));
  XOR2_X1   g792(.A(new_n962), .B(KEYINPUT124), .Z(new_n979));
  OAI211_X1 g793(.A(new_n953), .B(new_n965), .C1(new_n978), .C2(new_n979), .ZN(new_n980));
  AOI21_X1  g794(.A(new_n979), .B1(new_n977), .B2(new_n226), .ZN(new_n981));
  INV_X1    g795(.A(new_n965), .ZN(new_n982));
  OAI21_X1  g796(.A(new_n952), .B1(new_n981), .B2(new_n982), .ZN(new_n983));
  NAND2_X1  g797(.A1(new_n980), .A2(new_n983), .ZN(G72));
  NAND2_X1  g798(.A1(G472), .A2(G902), .ZN(new_n985));
  XOR2_X1   g799(.A(new_n985), .B(KEYINPUT63), .Z(new_n986));
  NAND2_X1  g800(.A1(new_n957), .A2(new_n958), .ZN(new_n987));
  OAI21_X1  g801(.A(new_n986), .B1(new_n987), .B2(new_n948), .ZN(new_n988));
  INV_X1    g802(.A(new_n348), .ZN(new_n989));
  NAND2_X1  g803(.A1(new_n988), .A2(new_n989), .ZN(new_n990));
  NAND2_X1  g804(.A1(new_n835), .A2(new_n845), .ZN(new_n991));
  NAND3_X1  g805(.A1(new_n679), .A2(new_n348), .A3(new_n986), .ZN(new_n992));
  OAI211_X1 g806(.A(new_n990), .B(new_n900), .C1(new_n991), .C2(new_n992), .ZN(new_n993));
  OAI21_X1  g807(.A(new_n986), .B1(new_n977), .B2(new_n948), .ZN(new_n994));
  INV_X1    g808(.A(KEYINPUT127), .ZN(new_n995));
  AOI21_X1  g809(.A(new_n679), .B1(new_n994), .B2(new_n995), .ZN(new_n996));
  OAI211_X1 g810(.A(KEYINPUT127), .B(new_n986), .C1(new_n977), .C2(new_n948), .ZN(new_n997));
  AOI21_X1  g811(.A(new_n993), .B1(new_n996), .B2(new_n997), .ZN(G57));
endmodule


