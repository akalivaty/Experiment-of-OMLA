

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300,
         n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311,
         n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322,
         n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333,
         n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344,
         n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355,
         n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
         n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
         n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
         n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
         n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410,
         n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421,
         n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432,
         n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443,
         n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454,
         n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465,
         n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
         n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487,
         n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
         n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
         n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586;

  XNOR2_X1 U322 ( .A(KEYINPUT93), .B(KEYINPUT25), .ZN(n449) );
  XOR2_X1 U323 ( .A(n340), .B(n339), .Z(n495) );
  AND2_X1 U324 ( .A1(G230GAT), .A2(G233GAT), .ZN(n290) );
  XNOR2_X1 U325 ( .A(KEYINPUT46), .B(KEYINPUT110), .ZN(n359) );
  XNOR2_X1 U326 ( .A(n360), .B(n359), .ZN(n377) );
  XNOR2_X1 U327 ( .A(n450), .B(n449), .ZN(n451) );
  INV_X1 U328 ( .A(KEYINPUT37), .ZN(n462) );
  XNOR2_X1 U329 ( .A(n334), .B(n290), .ZN(n292) );
  INV_X1 U330 ( .A(KEYINPUT55), .ZN(n424) );
  XNOR2_X1 U331 ( .A(n462), .B(KEYINPUT97), .ZN(n463) );
  XNOR2_X1 U332 ( .A(n329), .B(n328), .ZN(n330) );
  XNOR2_X1 U333 ( .A(n292), .B(n362), .ZN(n293) );
  XNOR2_X1 U334 ( .A(n464), .B(n463), .ZN(n504) );
  XNOR2_X1 U335 ( .A(n331), .B(n330), .ZN(n338) );
  XNOR2_X1 U336 ( .A(n303), .B(n302), .ZN(n304) );
  XNOR2_X1 U337 ( .A(n305), .B(n304), .ZN(n574) );
  INV_X1 U338 ( .A(G43GAT), .ZN(n468) );
  XNOR2_X1 U339 ( .A(n443), .B(n442), .ZN(n444) );
  XNOR2_X1 U340 ( .A(n468), .B(KEYINPUT40), .ZN(n469) );
  XNOR2_X1 U341 ( .A(n445), .B(n444), .ZN(G1349GAT) );
  XNOR2_X1 U342 ( .A(n470), .B(n469), .ZN(G1330GAT) );
  XOR2_X1 U343 ( .A(G176GAT), .B(G64GAT), .Z(n334) );
  XNOR2_X1 U344 ( .A(G71GAT), .B(G57GAT), .ZN(n291) );
  XNOR2_X1 U345 ( .A(n291), .B(KEYINPUT13), .ZN(n362) );
  XOR2_X1 U346 ( .A(n293), .B(KEYINPUT31), .Z(n305) );
  XOR2_X1 U347 ( .A(KEYINPUT71), .B(KEYINPUT72), .Z(n295) );
  XNOR2_X1 U348 ( .A(G99GAT), .B(G92GAT), .ZN(n294) );
  XNOR2_X1 U349 ( .A(n295), .B(n294), .ZN(n296) );
  XNOR2_X1 U350 ( .A(G85GAT), .B(n296), .ZN(n392) );
  XOR2_X1 U351 ( .A(KEYINPUT74), .B(KEYINPUT33), .Z(n298) );
  XNOR2_X1 U352 ( .A(G120GAT), .B(KEYINPUT73), .ZN(n297) );
  XNOR2_X1 U353 ( .A(n298), .B(n297), .ZN(n299) );
  XOR2_X1 U354 ( .A(n392), .B(n299), .Z(n303) );
  XOR2_X1 U355 ( .A(G78GAT), .B(G148GAT), .Z(n301) );
  XNOR2_X1 U356 ( .A(G106GAT), .B(G204GAT), .ZN(n300) );
  XNOR2_X1 U357 ( .A(n301), .B(n300), .ZN(n310) );
  XNOR2_X1 U358 ( .A(n310), .B(KEYINPUT32), .ZN(n302) );
  XNOR2_X1 U359 ( .A(n574), .B(KEYINPUT41), .ZN(n543) );
  XNOR2_X1 U360 ( .A(KEYINPUT100), .B(n543), .ZN(n525) );
  XOR2_X1 U361 ( .A(G211GAT), .B(KEYINPUT23), .Z(n312) );
  XNOR2_X1 U362 ( .A(KEYINPUT86), .B(KEYINPUT2), .ZN(n306) );
  XNOR2_X1 U363 ( .A(n306), .B(KEYINPUT85), .ZN(n307) );
  XOR2_X1 U364 ( .A(n307), .B(KEYINPUT3), .Z(n309) );
  XNOR2_X1 U365 ( .A(G155GAT), .B(G162GAT), .ZN(n308) );
  XNOR2_X1 U366 ( .A(n309), .B(n308), .ZN(n416) );
  XNOR2_X1 U367 ( .A(n416), .B(n310), .ZN(n311) );
  XNOR2_X1 U368 ( .A(n312), .B(n311), .ZN(n316) );
  XOR2_X1 U369 ( .A(KEYINPUT24), .B(KEYINPUT22), .Z(n314) );
  NAND2_X1 U370 ( .A1(G228GAT), .A2(G233GAT), .ZN(n313) );
  XNOR2_X1 U371 ( .A(n314), .B(n313), .ZN(n315) );
  XOR2_X1 U372 ( .A(n316), .B(n315), .Z(n323) );
  XNOR2_X1 U373 ( .A(G50GAT), .B(G22GAT), .ZN(n317) );
  XNOR2_X1 U374 ( .A(n317), .B(G141GAT), .ZN(n354) );
  XNOR2_X1 U375 ( .A(KEYINPUT82), .B(KEYINPUT21), .ZN(n318) );
  XNOR2_X1 U376 ( .A(n318), .B(KEYINPUT83), .ZN(n319) );
  XOR2_X1 U377 ( .A(n319), .B(KEYINPUT84), .Z(n321) );
  XNOR2_X1 U378 ( .A(G197GAT), .B(G218GAT), .ZN(n320) );
  XNOR2_X1 U379 ( .A(n321), .B(n320), .ZN(n340) );
  XNOR2_X1 U380 ( .A(n354), .B(n340), .ZN(n322) );
  XNOR2_X1 U381 ( .A(n323), .B(n322), .ZN(n455) );
  XOR2_X1 U382 ( .A(KEYINPUT19), .B(KEYINPUT17), .Z(n325) );
  XNOR2_X1 U383 ( .A(G169GAT), .B(KEYINPUT18), .ZN(n324) );
  XNOR2_X1 U384 ( .A(n325), .B(n324), .ZN(n427) );
  XOR2_X1 U385 ( .A(n427), .B(KEYINPUT89), .Z(n331) );
  XOR2_X1 U386 ( .A(KEYINPUT91), .B(KEYINPUT90), .Z(n327) );
  XNOR2_X1 U387 ( .A(G204GAT), .B(G92GAT), .ZN(n326) );
  XNOR2_X1 U388 ( .A(n327), .B(n326), .ZN(n329) );
  NAND2_X1 U389 ( .A1(G226GAT), .A2(G233GAT), .ZN(n328) );
  XOR2_X1 U390 ( .A(KEYINPUT77), .B(G211GAT), .Z(n333) );
  XNOR2_X1 U391 ( .A(G8GAT), .B(G183GAT), .ZN(n332) );
  XNOR2_X1 U392 ( .A(n333), .B(n332), .ZN(n366) );
  XOR2_X1 U393 ( .A(n334), .B(n366), .Z(n336) );
  XNOR2_X1 U394 ( .A(G36GAT), .B(G190GAT), .ZN(n335) );
  XNOR2_X1 U395 ( .A(n336), .B(n335), .ZN(n337) );
  XNOR2_X1 U396 ( .A(n338), .B(n337), .ZN(n339) );
  INV_X1 U397 ( .A(n495), .ZN(n510) );
  XNOR2_X1 U398 ( .A(G36GAT), .B(KEYINPUT8), .ZN(n341) );
  XNOR2_X1 U399 ( .A(n341), .B(G29GAT), .ZN(n342) );
  XOR2_X1 U400 ( .A(n342), .B(KEYINPUT7), .Z(n344) );
  XNOR2_X1 U401 ( .A(G43GAT), .B(KEYINPUT68), .ZN(n343) );
  XNOR2_X1 U402 ( .A(n344), .B(n343), .ZN(n391) );
  XOR2_X1 U403 ( .A(KEYINPUT69), .B(KEYINPUT66), .Z(n346) );
  XNOR2_X1 U404 ( .A(KEYINPUT30), .B(KEYINPUT65), .ZN(n345) );
  XNOR2_X1 U405 ( .A(n346), .B(n345), .ZN(n347) );
  XNOR2_X1 U406 ( .A(n391), .B(n347), .ZN(n358) );
  XOR2_X1 U407 ( .A(G15GAT), .B(G1GAT), .Z(n361) );
  XOR2_X1 U408 ( .A(G8GAT), .B(G197GAT), .Z(n349) );
  XNOR2_X1 U409 ( .A(G169GAT), .B(G113GAT), .ZN(n348) );
  XNOR2_X1 U410 ( .A(n349), .B(n348), .ZN(n350) );
  XOR2_X1 U411 ( .A(n361), .B(n350), .Z(n352) );
  NAND2_X1 U412 ( .A1(G229GAT), .A2(G233GAT), .ZN(n351) );
  XNOR2_X1 U413 ( .A(n352), .B(n351), .ZN(n353) );
  XOR2_X1 U414 ( .A(n353), .B(KEYINPUT29), .Z(n356) );
  XNOR2_X1 U415 ( .A(n354), .B(KEYINPUT67), .ZN(n355) );
  XNOR2_X1 U416 ( .A(n356), .B(n355), .ZN(n357) );
  XOR2_X1 U417 ( .A(n358), .B(n357), .Z(n540) );
  INV_X1 U418 ( .A(n540), .ZN(n569) );
  NAND2_X1 U419 ( .A1(n543), .A2(n569), .ZN(n360) );
  XOR2_X1 U420 ( .A(n362), .B(n361), .Z(n364) );
  NAND2_X1 U421 ( .A1(G231GAT), .A2(G233GAT), .ZN(n363) );
  XNOR2_X1 U422 ( .A(n364), .B(n363), .ZN(n365) );
  XOR2_X1 U423 ( .A(n365), .B(KEYINPUT12), .Z(n368) );
  XNOR2_X1 U424 ( .A(n366), .B(KEYINPUT14), .ZN(n367) );
  XNOR2_X1 U425 ( .A(n368), .B(n367), .ZN(n376) );
  XOR2_X1 U426 ( .A(G78GAT), .B(G155GAT), .Z(n370) );
  XNOR2_X1 U427 ( .A(G22GAT), .B(G127GAT), .ZN(n369) );
  XNOR2_X1 U428 ( .A(n370), .B(n369), .ZN(n374) );
  XOR2_X1 U429 ( .A(KEYINPUT15), .B(KEYINPUT78), .Z(n372) );
  XNOR2_X1 U430 ( .A(G64GAT), .B(KEYINPUT79), .ZN(n371) );
  XNOR2_X1 U431 ( .A(n372), .B(n371), .ZN(n373) );
  XOR2_X1 U432 ( .A(n374), .B(n373), .Z(n375) );
  XOR2_X1 U433 ( .A(n376), .B(n375), .Z(n471) );
  XOR2_X1 U434 ( .A(KEYINPUT109), .B(n471), .Z(n559) );
  NAND2_X1 U435 ( .A1(n377), .A2(n559), .ZN(n378) );
  XNOR2_X1 U436 ( .A(n378), .B(KEYINPUT111), .ZN(n395) );
  XOR2_X1 U437 ( .A(KEYINPUT75), .B(KEYINPUT64), .Z(n380) );
  XNOR2_X1 U438 ( .A(G218GAT), .B(KEYINPUT10), .ZN(n379) );
  XNOR2_X1 U439 ( .A(n380), .B(n379), .ZN(n384) );
  XOR2_X1 U440 ( .A(KEYINPUT11), .B(KEYINPUT9), .Z(n382) );
  XNOR2_X1 U441 ( .A(G162GAT), .B(KEYINPUT76), .ZN(n381) );
  XNOR2_X1 U442 ( .A(n382), .B(n381), .ZN(n383) );
  XOR2_X1 U443 ( .A(n384), .B(n383), .Z(n389) );
  XOR2_X1 U444 ( .A(G190GAT), .B(G134GAT), .Z(n426) );
  XOR2_X1 U445 ( .A(G106GAT), .B(n426), .Z(n386) );
  NAND2_X1 U446 ( .A1(G232GAT), .A2(G233GAT), .ZN(n385) );
  XNOR2_X1 U447 ( .A(n386), .B(n385), .ZN(n387) );
  XNOR2_X1 U448 ( .A(G50GAT), .B(n387), .ZN(n388) );
  XNOR2_X1 U449 ( .A(n389), .B(n388), .ZN(n390) );
  XNOR2_X1 U450 ( .A(n391), .B(n390), .ZN(n394) );
  INV_X1 U451 ( .A(n392), .ZN(n393) );
  XOR2_X1 U452 ( .A(n394), .B(n393), .Z(n561) );
  NAND2_X1 U453 ( .A1(n395), .A2(n561), .ZN(n396) );
  XNOR2_X1 U454 ( .A(n396), .B(KEYINPUT47), .ZN(n401) );
  XOR2_X1 U455 ( .A(n540), .B(KEYINPUT70), .Z(n555) );
  XNOR2_X1 U456 ( .A(KEYINPUT36), .B(n561), .ZN(n583) );
  NOR2_X1 U457 ( .A1(n583), .A2(n471), .ZN(n397) );
  XNOR2_X1 U458 ( .A(KEYINPUT45), .B(n397), .ZN(n398) );
  NAND2_X1 U459 ( .A1(n398), .A2(n574), .ZN(n399) );
  NOR2_X1 U460 ( .A1(n555), .A2(n399), .ZN(n400) );
  NOR2_X1 U461 ( .A1(n401), .A2(n400), .ZN(n402) );
  XNOR2_X1 U462 ( .A(KEYINPUT48), .B(n402), .ZN(n520) );
  NOR2_X1 U463 ( .A1(n510), .A2(n520), .ZN(n403) );
  XNOR2_X1 U464 ( .A(n403), .B(KEYINPUT54), .ZN(n423) );
  XOR2_X1 U465 ( .A(KEYINPUT6), .B(G57GAT), .Z(n405) );
  XNOR2_X1 U466 ( .A(G141GAT), .B(G1GAT), .ZN(n404) );
  XNOR2_X1 U467 ( .A(n405), .B(n404), .ZN(n409) );
  XOR2_X1 U468 ( .A(KEYINPUT4), .B(KEYINPUT87), .Z(n407) );
  XNOR2_X1 U469 ( .A(KEYINPUT5), .B(KEYINPUT88), .ZN(n406) );
  XNOR2_X1 U470 ( .A(n407), .B(n406), .ZN(n408) );
  XOR2_X1 U471 ( .A(n409), .B(n408), .Z(n418) );
  XOR2_X1 U472 ( .A(G85GAT), .B(G148GAT), .Z(n411) );
  XNOR2_X1 U473 ( .A(G29GAT), .B(G134GAT), .ZN(n410) );
  XNOR2_X1 U474 ( .A(n411), .B(n410), .ZN(n412) );
  XOR2_X1 U475 ( .A(KEYINPUT1), .B(n412), .Z(n414) );
  NAND2_X1 U476 ( .A1(G225GAT), .A2(G233GAT), .ZN(n413) );
  XNOR2_X1 U477 ( .A(n414), .B(n413), .ZN(n415) );
  XNOR2_X1 U478 ( .A(n416), .B(n415), .ZN(n417) );
  XNOR2_X1 U479 ( .A(n418), .B(n417), .ZN(n422) );
  XOR2_X1 U480 ( .A(KEYINPUT0), .B(G127GAT), .Z(n420) );
  XNOR2_X1 U481 ( .A(KEYINPUT80), .B(G120GAT), .ZN(n419) );
  XNOR2_X1 U482 ( .A(n420), .B(n419), .ZN(n421) );
  XNOR2_X1 U483 ( .A(G113GAT), .B(n421), .ZN(n437) );
  XOR2_X1 U484 ( .A(n422), .B(n437), .Z(n538) );
  INV_X1 U485 ( .A(n538), .ZN(n507) );
  NAND2_X1 U486 ( .A1(n423), .A2(n507), .ZN(n567) );
  NOR2_X1 U487 ( .A1(n455), .A2(n567), .ZN(n425) );
  XNOR2_X1 U488 ( .A(n425), .B(n424), .ZN(n440) );
  XOR2_X1 U489 ( .A(n427), .B(n426), .Z(n429) );
  NAND2_X1 U490 ( .A1(G227GAT), .A2(G233GAT), .ZN(n428) );
  XNOR2_X1 U491 ( .A(n429), .B(n428), .ZN(n433) );
  XOR2_X1 U492 ( .A(G176GAT), .B(G183GAT), .Z(n431) );
  XNOR2_X1 U493 ( .A(G15GAT), .B(KEYINPUT81), .ZN(n430) );
  XNOR2_X1 U494 ( .A(n431), .B(n430), .ZN(n432) );
  XOR2_X1 U495 ( .A(n433), .B(n432), .Z(n439) );
  XOR2_X1 U496 ( .A(KEYINPUT20), .B(G71GAT), .Z(n435) );
  XNOR2_X1 U497 ( .A(G43GAT), .B(G99GAT), .ZN(n434) );
  XNOR2_X1 U498 ( .A(n435), .B(n434), .ZN(n436) );
  XOR2_X1 U499 ( .A(n437), .B(n436), .Z(n438) );
  XOR2_X1 U500 ( .A(n439), .B(n438), .Z(n512) );
  INV_X1 U501 ( .A(n512), .ZN(n522) );
  NAND2_X1 U502 ( .A1(n440), .A2(n522), .ZN(n441) );
  XNOR2_X1 U503 ( .A(KEYINPUT120), .B(n441), .ZN(n562) );
  INV_X1 U504 ( .A(n562), .ZN(n556) );
  NAND2_X1 U505 ( .A1(n525), .A2(n556), .ZN(n445) );
  XOR2_X1 U506 ( .A(G176GAT), .B(KEYINPUT122), .Z(n443) );
  XNOR2_X1 U507 ( .A(KEYINPUT56), .B(KEYINPUT57), .ZN(n442) );
  INV_X1 U508 ( .A(KEYINPUT98), .ZN(n466) );
  NAND2_X1 U509 ( .A1(n512), .A2(n455), .ZN(n447) );
  INV_X1 U510 ( .A(KEYINPUT26), .ZN(n446) );
  XNOR2_X1 U511 ( .A(n447), .B(n446), .ZN(n566) );
  XNOR2_X1 U512 ( .A(KEYINPUT27), .B(n495), .ZN(n456) );
  NAND2_X1 U513 ( .A1(n566), .A2(n456), .ZN(n537) );
  XNOR2_X1 U514 ( .A(n537), .B(KEYINPUT92), .ZN(n452) );
  NOR2_X1 U515 ( .A1(n512), .A2(n510), .ZN(n448) );
  OR2_X1 U516 ( .A1(n455), .A2(n448), .ZN(n450) );
  NAND2_X1 U517 ( .A1(n452), .A2(n451), .ZN(n453) );
  XNOR2_X1 U518 ( .A(n453), .B(KEYINPUT94), .ZN(n454) );
  NAND2_X1 U519 ( .A1(n454), .A2(n507), .ZN(n459) );
  XNOR2_X1 U520 ( .A(n455), .B(KEYINPUT28), .ZN(n500) );
  INV_X1 U521 ( .A(n500), .ZN(n516) );
  NAND2_X1 U522 ( .A1(n516), .A2(n456), .ZN(n457) );
  NOR2_X1 U523 ( .A1(n507), .A2(n457), .ZN(n521) );
  NAND2_X1 U524 ( .A1(n521), .A2(n512), .ZN(n458) );
  NAND2_X1 U525 ( .A1(n459), .A2(n458), .ZN(n473) );
  NAND2_X1 U526 ( .A1(n473), .A2(n471), .ZN(n460) );
  XNOR2_X1 U527 ( .A(n460), .B(KEYINPUT96), .ZN(n461) );
  NOR2_X1 U528 ( .A1(n583), .A2(n461), .ZN(n464) );
  NAND2_X1 U529 ( .A1(n574), .A2(n555), .ZN(n475) );
  NOR2_X1 U530 ( .A1(n504), .A2(n475), .ZN(n465) );
  XNOR2_X1 U531 ( .A(n466), .B(n465), .ZN(n467) );
  XNOR2_X1 U532 ( .A(KEYINPUT38), .B(n467), .ZN(n487) );
  NOR2_X1 U533 ( .A1(n512), .A2(n487), .ZN(n470) );
  XOR2_X1 U534 ( .A(KEYINPUT95), .B(KEYINPUT34), .Z(n477) );
  INV_X1 U535 ( .A(n471), .ZN(n580) );
  NAND2_X1 U536 ( .A1(n561), .A2(n580), .ZN(n472) );
  XOR2_X1 U537 ( .A(KEYINPUT16), .B(n472), .Z(n474) );
  NAND2_X1 U538 ( .A1(n474), .A2(n473), .ZN(n489) );
  NOR2_X1 U539 ( .A1(n475), .A2(n489), .ZN(n482) );
  NAND2_X1 U540 ( .A1(n482), .A2(n538), .ZN(n476) );
  XNOR2_X1 U541 ( .A(n477), .B(n476), .ZN(n478) );
  XNOR2_X1 U542 ( .A(G1GAT), .B(n478), .ZN(G1324GAT) );
  NAND2_X1 U543 ( .A1(n495), .A2(n482), .ZN(n479) );
  XNOR2_X1 U544 ( .A(G8GAT), .B(n479), .ZN(G1325GAT) );
  XOR2_X1 U545 ( .A(G15GAT), .B(KEYINPUT35), .Z(n481) );
  NAND2_X1 U546 ( .A1(n482), .A2(n522), .ZN(n480) );
  XNOR2_X1 U547 ( .A(n481), .B(n480), .ZN(G1326GAT) );
  NAND2_X1 U548 ( .A1(n500), .A2(n482), .ZN(n483) );
  XNOR2_X1 U549 ( .A(n483), .B(G22GAT), .ZN(G1327GAT) );
  NOR2_X1 U550 ( .A1(n507), .A2(n487), .ZN(n484) );
  XNOR2_X1 U551 ( .A(n484), .B(KEYINPUT39), .ZN(n485) );
  XNOR2_X1 U552 ( .A(G29GAT), .B(n485), .ZN(G1328GAT) );
  NOR2_X1 U553 ( .A1(n510), .A2(n487), .ZN(n486) );
  XOR2_X1 U554 ( .A(G36GAT), .B(n486), .Z(G1329GAT) );
  NOR2_X1 U555 ( .A1(n516), .A2(n487), .ZN(n488) );
  XOR2_X1 U556 ( .A(G50GAT), .B(n488), .Z(G1331GAT) );
  XOR2_X1 U557 ( .A(KEYINPUT102), .B(KEYINPUT101), .Z(n491) );
  NAND2_X1 U558 ( .A1(n525), .A2(n540), .ZN(n505) );
  NOR2_X1 U559 ( .A1(n505), .A2(n489), .ZN(n501) );
  NAND2_X1 U560 ( .A1(n501), .A2(n538), .ZN(n490) );
  XNOR2_X1 U561 ( .A(n491), .B(n490), .ZN(n492) );
  XOR2_X1 U562 ( .A(n492), .B(KEYINPUT42), .Z(n494) );
  XNOR2_X1 U563 ( .A(G57GAT), .B(KEYINPUT99), .ZN(n493) );
  XNOR2_X1 U564 ( .A(n494), .B(n493), .ZN(G1332GAT) );
  XOR2_X1 U565 ( .A(G64GAT), .B(KEYINPUT103), .Z(n497) );
  NAND2_X1 U566 ( .A1(n501), .A2(n495), .ZN(n496) );
  XNOR2_X1 U567 ( .A(n497), .B(n496), .ZN(G1333GAT) );
  NAND2_X1 U568 ( .A1(n501), .A2(n522), .ZN(n498) );
  XNOR2_X1 U569 ( .A(n498), .B(KEYINPUT104), .ZN(n499) );
  XNOR2_X1 U570 ( .A(G71GAT), .B(n499), .ZN(G1334GAT) );
  XOR2_X1 U571 ( .A(G78GAT), .B(KEYINPUT43), .Z(n503) );
  NAND2_X1 U572 ( .A1(n501), .A2(n500), .ZN(n502) );
  XNOR2_X1 U573 ( .A(n503), .B(n502), .ZN(G1335GAT) );
  NOR2_X1 U574 ( .A1(n505), .A2(n504), .ZN(n506) );
  XNOR2_X1 U575 ( .A(n506), .B(KEYINPUT105), .ZN(n515) );
  NOR2_X1 U576 ( .A1(n507), .A2(n515), .ZN(n508) );
  XOR2_X1 U577 ( .A(n508), .B(KEYINPUT106), .Z(n509) );
  XNOR2_X1 U578 ( .A(G85GAT), .B(n509), .ZN(G1336GAT) );
  NOR2_X1 U579 ( .A1(n510), .A2(n515), .ZN(n511) );
  XOR2_X1 U580 ( .A(G92GAT), .B(n511), .Z(G1337GAT) );
  NOR2_X1 U581 ( .A1(n512), .A2(n515), .ZN(n514) );
  XNOR2_X1 U582 ( .A(G99GAT), .B(KEYINPUT107), .ZN(n513) );
  XNOR2_X1 U583 ( .A(n514), .B(n513), .ZN(G1338GAT) );
  NOR2_X1 U584 ( .A1(n516), .A2(n515), .ZN(n518) );
  XNOR2_X1 U585 ( .A(KEYINPUT44), .B(KEYINPUT108), .ZN(n517) );
  XNOR2_X1 U586 ( .A(n518), .B(n517), .ZN(n519) );
  XOR2_X1 U587 ( .A(G106GAT), .B(n519), .Z(G1339GAT) );
  NAND2_X1 U588 ( .A1(n522), .A2(n521), .ZN(n523) );
  NOR2_X1 U589 ( .A1(n520), .A2(n523), .ZN(n528) );
  NAND2_X1 U590 ( .A1(n555), .A2(n528), .ZN(n524) );
  XNOR2_X1 U591 ( .A(n524), .B(G113GAT), .ZN(G1340GAT) );
  XOR2_X1 U592 ( .A(G120GAT), .B(KEYINPUT49), .Z(n527) );
  NAND2_X1 U593 ( .A1(n528), .A2(n525), .ZN(n526) );
  XNOR2_X1 U594 ( .A(n527), .B(n526), .ZN(G1341GAT) );
  INV_X1 U595 ( .A(n528), .ZN(n532) );
  NOR2_X1 U596 ( .A1(n559), .A2(n532), .ZN(n530) );
  XNOR2_X1 U597 ( .A(KEYINPUT50), .B(KEYINPUT112), .ZN(n529) );
  XNOR2_X1 U598 ( .A(n530), .B(n529), .ZN(n531) );
  XOR2_X1 U599 ( .A(G127GAT), .B(n531), .Z(G1342GAT) );
  NOR2_X1 U600 ( .A1(n532), .A2(n561), .ZN(n536) );
  XOR2_X1 U601 ( .A(KEYINPUT113), .B(KEYINPUT51), .Z(n534) );
  XNOR2_X1 U602 ( .A(G134GAT), .B(KEYINPUT114), .ZN(n533) );
  XNOR2_X1 U603 ( .A(n534), .B(n533), .ZN(n535) );
  XNOR2_X1 U604 ( .A(n536), .B(n535), .ZN(G1343GAT) );
  NOR2_X1 U605 ( .A1(n520), .A2(n537), .ZN(n539) );
  NAND2_X1 U606 ( .A1(n539), .A2(n538), .ZN(n552) );
  NOR2_X1 U607 ( .A1(n540), .A2(n552), .ZN(n542) );
  XNOR2_X1 U608 ( .A(G141GAT), .B(KEYINPUT115), .ZN(n541) );
  XNOR2_X1 U609 ( .A(n542), .B(n541), .ZN(G1344GAT) );
  XOR2_X1 U610 ( .A(KEYINPUT53), .B(KEYINPUT117), .Z(n545) );
  INV_X1 U611 ( .A(n552), .ZN(n549) );
  NAND2_X1 U612 ( .A1(n549), .A2(n543), .ZN(n544) );
  XNOR2_X1 U613 ( .A(n545), .B(n544), .ZN(n546) );
  XOR2_X1 U614 ( .A(n546), .B(KEYINPUT116), .Z(n548) );
  XNOR2_X1 U615 ( .A(G148GAT), .B(KEYINPUT52), .ZN(n547) );
  XNOR2_X1 U616 ( .A(n548), .B(n547), .ZN(G1345GAT) );
  NAND2_X1 U617 ( .A1(n580), .A2(n549), .ZN(n550) );
  XNOR2_X1 U618 ( .A(n550), .B(KEYINPUT118), .ZN(n551) );
  XNOR2_X1 U619 ( .A(G155GAT), .B(n551), .ZN(G1346GAT) );
  NOR2_X1 U620 ( .A1(n561), .A2(n552), .ZN(n554) );
  XNOR2_X1 U621 ( .A(G162GAT), .B(KEYINPUT119), .ZN(n553) );
  XNOR2_X1 U622 ( .A(n554), .B(n553), .ZN(G1347GAT) );
  XOR2_X1 U623 ( .A(G169GAT), .B(KEYINPUT121), .Z(n558) );
  NAND2_X1 U624 ( .A1(n556), .A2(n555), .ZN(n557) );
  XNOR2_X1 U625 ( .A(n558), .B(n557), .ZN(G1348GAT) );
  NOR2_X1 U626 ( .A1(n559), .A2(n562), .ZN(n560) );
  XOR2_X1 U627 ( .A(G183GAT), .B(n560), .Z(G1350GAT) );
  NOR2_X1 U628 ( .A1(n562), .A2(n561), .ZN(n564) );
  XNOR2_X1 U629 ( .A(KEYINPUT58), .B(KEYINPUT123), .ZN(n563) );
  XNOR2_X1 U630 ( .A(n564), .B(n563), .ZN(n565) );
  XNOR2_X1 U631 ( .A(G190GAT), .B(n565), .ZN(G1351GAT) );
  INV_X1 U632 ( .A(n566), .ZN(n568) );
  NOR2_X1 U633 ( .A1(n568), .A2(n567), .ZN(n579) );
  NAND2_X1 U634 ( .A1(n579), .A2(n569), .ZN(n573) );
  XOR2_X1 U635 ( .A(KEYINPUT59), .B(KEYINPUT124), .Z(n571) );
  XNOR2_X1 U636 ( .A(G197GAT), .B(KEYINPUT60), .ZN(n570) );
  XNOR2_X1 U637 ( .A(n571), .B(n570), .ZN(n572) );
  XNOR2_X1 U638 ( .A(n573), .B(n572), .ZN(G1352GAT) );
  INV_X1 U639 ( .A(n579), .ZN(n582) );
  NOR2_X1 U640 ( .A1(n582), .A2(n574), .ZN(n578) );
  XOR2_X1 U641 ( .A(KEYINPUT125), .B(KEYINPUT61), .Z(n576) );
  XNOR2_X1 U642 ( .A(G204GAT), .B(KEYINPUT126), .ZN(n575) );
  XNOR2_X1 U643 ( .A(n576), .B(n575), .ZN(n577) );
  XNOR2_X1 U644 ( .A(n578), .B(n577), .ZN(G1353GAT) );
  NAND2_X1 U645 ( .A1(n580), .A2(n579), .ZN(n581) );
  XNOR2_X1 U646 ( .A(n581), .B(G211GAT), .ZN(G1354GAT) );
  NOR2_X1 U647 ( .A1(n583), .A2(n582), .ZN(n585) );
  XNOR2_X1 U648 ( .A(KEYINPUT127), .B(KEYINPUT62), .ZN(n584) );
  XNOR2_X1 U649 ( .A(n585), .B(n584), .ZN(n586) );
  XNOR2_X1 U650 ( .A(G218GAT), .B(n586), .ZN(G1355GAT) );
endmodule

