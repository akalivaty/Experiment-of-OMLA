//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 1 1 0 0 1 0 0 1 1 0 0 0 0 1 1 1 0 1 1 1 0 1 0 1 0 1 1 0 1 1 0 1 1 1 1 1 0 1 0 0 0 0 0 0 0 0 1 0 0 1 1 1 0 1 0 1 1 1 1 1 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:42:30 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n205, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1201, new_n1202, new_n1203, new_n1204, new_n1205,
    new_n1206, new_n1207, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1226, new_n1227, new_n1228, new_n1229, new_n1230,
    new_n1231, new_n1232, new_n1233, new_n1234, new_n1235, new_n1236,
    new_n1238, new_n1239, new_n1240, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1289, new_n1290, new_n1291, new_n1292, new_n1293,
    new_n1294, new_n1295, new_n1296, new_n1297, new_n1298;
  INV_X1    g0000(.A(G58), .ZN(new_n201));
  INV_X1    g0001(.A(G68), .ZN(new_n202));
  NAND3_X1  g0002(.A1(new_n201), .A2(new_n202), .A3(KEYINPUT64), .ZN(new_n203));
  INV_X1    g0003(.A(KEYINPUT64), .ZN(new_n204));
  OAI21_X1  g0004(.A(new_n204), .B1(G58), .B2(G68), .ZN(new_n205));
  AOI211_X1 g0005(.A(G50), .B(G77), .C1(new_n203), .C2(new_n205), .ZN(G353));
  OAI21_X1  g0006(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0007(.A(G1), .ZN(new_n208));
  INV_X1    g0008(.A(G20), .ZN(new_n209));
  NOR2_X1   g0009(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  INV_X1    g0010(.A(new_n210), .ZN(new_n211));
  NOR2_X1   g0011(.A1(new_n211), .A2(G13), .ZN(new_n212));
  OAI211_X1 g0012(.A(new_n212), .B(G250), .C1(G257), .C2(G264), .ZN(new_n213));
  XOR2_X1   g0013(.A(KEYINPUT65), .B(KEYINPUT0), .Z(new_n214));
  XNOR2_X1  g0014(.A(new_n213), .B(new_n214), .ZN(new_n215));
  AOI22_X1  g0015(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n216));
  INV_X1    g0016(.A(G238), .ZN(new_n217));
  INV_X1    g0017(.A(G87), .ZN(new_n218));
  INV_X1    g0018(.A(G250), .ZN(new_n219));
  OAI221_X1 g0019(.A(new_n216), .B1(new_n202), .B2(new_n217), .C1(new_n218), .C2(new_n219), .ZN(new_n220));
  AOI22_X1  g0020(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n221));
  AOI22_X1  g0021(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n222));
  NAND2_X1  g0022(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  OAI21_X1  g0023(.A(new_n211), .B1(new_n220), .B2(new_n223), .ZN(new_n224));
  XNOR2_X1  g0024(.A(new_n224), .B(KEYINPUT1), .ZN(new_n225));
  NAND2_X1  g0025(.A1(G1), .A2(G13), .ZN(new_n226));
  NOR2_X1   g0026(.A1(new_n226), .A2(new_n209), .ZN(new_n227));
  NAND2_X1  g0027(.A1(new_n203), .A2(new_n205), .ZN(new_n228));
  INV_X1    g0028(.A(G50), .ZN(new_n229));
  NOR2_X1   g0029(.A1(new_n228), .A2(new_n229), .ZN(new_n230));
  AOI211_X1 g0030(.A(new_n215), .B(new_n225), .C1(new_n227), .C2(new_n230), .ZN(G361));
  XNOR2_X1  g0031(.A(G238), .B(G244), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n232), .B(G232), .ZN(new_n233));
  XNOR2_X1  g0033(.A(KEYINPUT2), .B(G226), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n233), .B(new_n234), .ZN(new_n235));
  XOR2_X1   g0035(.A(G264), .B(G270), .Z(new_n236));
  XNOR2_X1  g0036(.A(G250), .B(G257), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n235), .B(new_n238), .ZN(G358));
  XNOR2_X1  g0039(.A(G68), .B(G77), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n240), .B(new_n201), .ZN(new_n241));
  XOR2_X1   g0041(.A(KEYINPUT66), .B(G50), .Z(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XNOR2_X1  g0043(.A(G87), .B(G97), .ZN(new_n244));
  XNOR2_X1  g0044(.A(G107), .B(G116), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n244), .B(new_n245), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n243), .B(new_n246), .ZN(G351));
  XNOR2_X1  g0047(.A(KEYINPUT8), .B(G58), .ZN(new_n248));
  INV_X1    g0048(.A(new_n248), .ZN(new_n249));
  OAI21_X1  g0049(.A(KEYINPUT68), .B1(new_n209), .B2(G1), .ZN(new_n250));
  INV_X1    g0050(.A(KEYINPUT68), .ZN(new_n251));
  NAND3_X1  g0051(.A1(new_n251), .A2(new_n208), .A3(G20), .ZN(new_n252));
  NAND2_X1  g0052(.A1(new_n250), .A2(new_n252), .ZN(new_n253));
  NAND3_X1  g0053(.A1(new_n208), .A2(G13), .A3(G20), .ZN(new_n254));
  NAND3_X1  g0054(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n255));
  NAND3_X1  g0055(.A1(new_n254), .A2(new_n226), .A3(new_n255), .ZN(new_n256));
  OAI21_X1  g0056(.A(new_n249), .B1(new_n253), .B2(new_n256), .ZN(new_n257));
  NAND2_X1  g0057(.A1(new_n248), .A2(new_n254), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n257), .A2(new_n258), .ZN(new_n259));
  XNOR2_X1  g0059(.A(new_n259), .B(KEYINPUT77), .ZN(new_n260));
  INV_X1    g0060(.A(KEYINPUT3), .ZN(new_n261));
  INV_X1    g0061(.A(G33), .ZN(new_n262));
  NAND2_X1  g0062(.A1(new_n261), .A2(new_n262), .ZN(new_n263));
  NAND2_X1  g0063(.A1(KEYINPUT3), .A2(G33), .ZN(new_n264));
  NAND3_X1  g0064(.A1(new_n263), .A2(new_n209), .A3(new_n264), .ZN(new_n265));
  INV_X1    g0065(.A(KEYINPUT76), .ZN(new_n266));
  XNOR2_X1  g0066(.A(KEYINPUT75), .B(KEYINPUT7), .ZN(new_n267));
  NAND3_X1  g0067(.A1(new_n265), .A2(new_n266), .A3(new_n267), .ZN(new_n268));
  AND2_X1   g0068(.A1(KEYINPUT3), .A2(G33), .ZN(new_n269));
  NOR2_X1   g0069(.A1(KEYINPUT3), .A2(G33), .ZN(new_n270));
  NOR2_X1   g0070(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  NAND3_X1  g0071(.A1(new_n271), .A2(KEYINPUT7), .A3(new_n209), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n268), .A2(new_n272), .ZN(new_n273));
  AOI21_X1  g0073(.A(new_n266), .B1(new_n265), .B2(new_n267), .ZN(new_n274));
  OAI21_X1  g0074(.A(G68), .B1(new_n273), .B2(new_n274), .ZN(new_n275));
  OAI211_X1 g0075(.A(new_n203), .B(new_n205), .C1(new_n201), .C2(new_n202), .ZN(new_n276));
  NOR2_X1   g0076(.A1(G20), .A2(G33), .ZN(new_n277));
  AOI22_X1  g0077(.A1(new_n276), .A2(G20), .B1(G159), .B2(new_n277), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n275), .A2(new_n278), .ZN(new_n279));
  INV_X1    g0079(.A(KEYINPUT16), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n279), .A2(new_n280), .ZN(new_n281));
  INV_X1    g0081(.A(KEYINPUT7), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n282), .A2(KEYINPUT75), .ZN(new_n283));
  INV_X1    g0083(.A(KEYINPUT75), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n284), .A2(KEYINPUT7), .ZN(new_n285));
  NAND2_X1  g0085(.A1(new_n283), .A2(new_n285), .ZN(new_n286));
  NOR2_X1   g0086(.A1(new_n265), .A2(new_n286), .ZN(new_n287));
  NOR3_X1   g0087(.A1(new_n269), .A2(new_n270), .A3(G20), .ZN(new_n288));
  OAI21_X1  g0088(.A(G68), .B1(new_n288), .B2(new_n282), .ZN(new_n289));
  OAI211_X1 g0089(.A(new_n278), .B(KEYINPUT16), .C1(new_n287), .C2(new_n289), .ZN(new_n290));
  NAND2_X1  g0090(.A1(new_n255), .A2(new_n226), .ZN(new_n291));
  AND2_X1   g0091(.A1(new_n290), .A2(new_n291), .ZN(new_n292));
  AOI21_X1  g0092(.A(new_n260), .B1(new_n281), .B2(new_n292), .ZN(new_n293));
  INV_X1    g0093(.A(KEYINPUT80), .ZN(new_n294));
  OAI211_X1 g0094(.A(G226), .B(G1698), .C1(new_n269), .C2(new_n270), .ZN(new_n295));
  INV_X1    g0095(.A(G1698), .ZN(new_n296));
  OAI211_X1 g0096(.A(G223), .B(new_n296), .C1(new_n269), .C2(new_n270), .ZN(new_n297));
  NAND2_X1  g0097(.A1(G33), .A2(G87), .ZN(new_n298));
  INV_X1    g0098(.A(KEYINPUT78), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n298), .A2(new_n299), .ZN(new_n300));
  NAND3_X1  g0100(.A1(KEYINPUT78), .A2(G33), .A3(G87), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n300), .A2(new_n301), .ZN(new_n302));
  NAND3_X1  g0102(.A1(new_n295), .A2(new_n297), .A3(new_n302), .ZN(new_n303));
  AOI21_X1  g0103(.A(new_n226), .B1(G33), .B2(G41), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n303), .A2(new_n304), .ZN(new_n305));
  INV_X1    g0105(.A(KEYINPUT79), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n305), .A2(new_n306), .ZN(new_n307));
  NAND3_X1  g0107(.A1(new_n303), .A2(KEYINPUT79), .A3(new_n304), .ZN(new_n308));
  NAND2_X1  g0108(.A1(G33), .A2(G41), .ZN(new_n309));
  NAND3_X1  g0109(.A1(new_n309), .A2(G1), .A3(G13), .ZN(new_n310));
  OAI21_X1  g0110(.A(new_n208), .B1(G41), .B2(G45), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n310), .A2(new_n311), .ZN(new_n312));
  INV_X1    g0112(.A(G232), .ZN(new_n313));
  INV_X1    g0113(.A(G274), .ZN(new_n314));
  OAI22_X1  g0114(.A1(new_n312), .A2(new_n313), .B1(new_n314), .B2(new_n311), .ZN(new_n315));
  NOR2_X1   g0115(.A1(new_n315), .A2(G190), .ZN(new_n316));
  NAND3_X1  g0116(.A1(new_n307), .A2(new_n308), .A3(new_n316), .ZN(new_n317));
  INV_X1    g0117(.A(new_n315), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n305), .A2(new_n318), .ZN(new_n319));
  INV_X1    g0119(.A(G200), .ZN(new_n320));
  NAND2_X1  g0120(.A1(new_n319), .A2(new_n320), .ZN(new_n321));
  AOI21_X1  g0121(.A(new_n294), .B1(new_n317), .B2(new_n321), .ZN(new_n322));
  AND3_X1   g0122(.A1(new_n317), .A2(new_n294), .A3(new_n321), .ZN(new_n323));
  OAI21_X1  g0123(.A(new_n293), .B1(new_n322), .B2(new_n323), .ZN(new_n324));
  INV_X1    g0124(.A(KEYINPUT17), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n324), .A2(new_n325), .ZN(new_n326));
  INV_X1    g0126(.A(G179), .ZN(new_n327));
  NAND4_X1  g0127(.A1(new_n307), .A2(new_n327), .A3(new_n318), .A4(new_n308), .ZN(new_n328));
  INV_X1    g0128(.A(G169), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n319), .A2(new_n329), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n328), .A2(new_n330), .ZN(new_n331));
  OAI21_X1  g0131(.A(KEYINPUT18), .B1(new_n293), .B2(new_n331), .ZN(new_n332));
  INV_X1    g0132(.A(new_n331), .ZN(new_n333));
  INV_X1    g0133(.A(KEYINPUT77), .ZN(new_n334));
  XNOR2_X1  g0134(.A(new_n259), .B(new_n334), .ZN(new_n335));
  AOI21_X1  g0135(.A(KEYINPUT16), .B1(new_n275), .B2(new_n278), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n290), .A2(new_n291), .ZN(new_n337));
  OAI21_X1  g0137(.A(new_n335), .B1(new_n336), .B2(new_n337), .ZN(new_n338));
  INV_X1    g0138(.A(KEYINPUT18), .ZN(new_n339));
  NAND3_X1  g0139(.A1(new_n333), .A2(new_n338), .A3(new_n339), .ZN(new_n340));
  OAI211_X1 g0140(.A(new_n293), .B(KEYINPUT17), .C1(new_n322), .C2(new_n323), .ZN(new_n341));
  NAND4_X1  g0141(.A1(new_n326), .A2(new_n332), .A3(new_n340), .A4(new_n341), .ZN(new_n342));
  INV_X1    g0142(.A(new_n342), .ZN(new_n343));
  NAND2_X1  g0143(.A1(new_n263), .A2(new_n264), .ZN(new_n344));
  NAND3_X1  g0144(.A1(new_n344), .A2(G222), .A3(new_n296), .ZN(new_n345));
  INV_X1    g0145(.A(G77), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n344), .A2(G1698), .ZN(new_n347));
  INV_X1    g0147(.A(G223), .ZN(new_n348));
  OAI221_X1 g0148(.A(new_n345), .B1(new_n346), .B2(new_n344), .C1(new_n347), .C2(new_n348), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n349), .A2(new_n304), .ZN(new_n350));
  NOR2_X1   g0150(.A1(new_n311), .A2(new_n314), .ZN(new_n351));
  INV_X1    g0151(.A(new_n312), .ZN(new_n352));
  XNOR2_X1  g0152(.A(KEYINPUT67), .B(G226), .ZN(new_n353));
  AOI21_X1  g0153(.A(new_n351), .B1(new_n352), .B2(new_n353), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n350), .A2(new_n354), .ZN(new_n355));
  INV_X1    g0155(.A(new_n355), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n356), .A2(new_n327), .ZN(new_n357));
  AOI21_X1  g0157(.A(new_n209), .B1(new_n228), .B2(new_n229), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n277), .A2(G150), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n209), .A2(G33), .ZN(new_n360));
  OAI21_X1  g0160(.A(new_n359), .B1(new_n248), .B2(new_n360), .ZN(new_n361));
  OAI21_X1  g0161(.A(new_n291), .B1(new_n358), .B2(new_n361), .ZN(new_n362));
  NOR2_X1   g0162(.A1(new_n253), .A2(new_n256), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n363), .A2(G50), .ZN(new_n364));
  OAI211_X1 g0164(.A(new_n362), .B(new_n364), .C1(G50), .C2(new_n254), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n355), .A2(new_n329), .ZN(new_n366));
  NAND3_X1  g0166(.A1(new_n357), .A2(new_n365), .A3(new_n366), .ZN(new_n367));
  INV_X1    g0167(.A(new_n367), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n356), .A2(G190), .ZN(new_n369));
  XNOR2_X1  g0169(.A(new_n369), .B(KEYINPUT73), .ZN(new_n370));
  INV_X1    g0170(.A(new_n370), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n355), .A2(G200), .ZN(new_n372));
  OR2_X1    g0172(.A1(new_n372), .A2(KEYINPUT72), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n372), .A2(KEYINPUT72), .ZN(new_n374));
  XNOR2_X1  g0174(.A(new_n365), .B(KEYINPUT9), .ZN(new_n375));
  NAND3_X1  g0175(.A1(new_n373), .A2(new_n374), .A3(new_n375), .ZN(new_n376));
  OAI21_X1  g0176(.A(KEYINPUT10), .B1(new_n371), .B2(new_n376), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n373), .A2(new_n374), .ZN(new_n378));
  NOR2_X1   g0178(.A1(new_n378), .A2(KEYINPUT10), .ZN(new_n379));
  OR2_X1    g0179(.A1(new_n375), .A2(KEYINPUT71), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n375), .A2(KEYINPUT71), .ZN(new_n381));
  NAND4_X1  g0181(.A1(new_n379), .A2(new_n370), .A3(new_n380), .A4(new_n381), .ZN(new_n382));
  AOI21_X1  g0182(.A(new_n368), .B1(new_n377), .B2(new_n382), .ZN(new_n383));
  OAI211_X1 g0183(.A(G232), .B(G1698), .C1(new_n269), .C2(new_n270), .ZN(new_n384));
  OAI211_X1 g0184(.A(G226), .B(new_n296), .C1(new_n269), .C2(new_n270), .ZN(new_n385));
  AND3_X1   g0185(.A1(KEYINPUT74), .A2(G33), .A3(G97), .ZN(new_n386));
  AOI21_X1  g0186(.A(KEYINPUT74), .B1(G33), .B2(G97), .ZN(new_n387));
  NOR2_X1   g0187(.A1(new_n386), .A2(new_n387), .ZN(new_n388));
  NAND3_X1  g0188(.A1(new_n384), .A2(new_n385), .A3(new_n388), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n389), .A2(new_n304), .ZN(new_n390));
  INV_X1    g0190(.A(KEYINPUT13), .ZN(new_n391));
  AOI21_X1  g0191(.A(new_n351), .B1(new_n352), .B2(G238), .ZN(new_n392));
  AND3_X1   g0192(.A1(new_n390), .A2(new_n391), .A3(new_n392), .ZN(new_n393));
  AOI21_X1  g0193(.A(new_n391), .B1(new_n390), .B2(new_n392), .ZN(new_n394));
  OAI21_X1  g0194(.A(G169), .B1(new_n393), .B2(new_n394), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n395), .A2(KEYINPUT14), .ZN(new_n396));
  INV_X1    g0196(.A(KEYINPUT14), .ZN(new_n397));
  OAI211_X1 g0197(.A(new_n397), .B(G169), .C1(new_n393), .C2(new_n394), .ZN(new_n398));
  NOR2_X1   g0198(.A1(new_n393), .A2(new_n394), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n399), .A2(G179), .ZN(new_n400));
  NAND3_X1  g0200(.A1(new_n396), .A2(new_n398), .A3(new_n400), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n277), .A2(G50), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n202), .A2(G20), .ZN(new_n403));
  OAI211_X1 g0203(.A(new_n402), .B(new_n403), .C1(new_n346), .C2(new_n360), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n404), .A2(new_n291), .ZN(new_n405));
  INV_X1    g0205(.A(KEYINPUT11), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n405), .A2(new_n406), .ZN(new_n407));
  NOR2_X1   g0207(.A1(new_n254), .A2(G68), .ZN(new_n408));
  INV_X1    g0208(.A(KEYINPUT12), .ZN(new_n409));
  XNOR2_X1  g0209(.A(new_n408), .B(new_n409), .ZN(new_n410));
  NAND3_X1  g0210(.A1(new_n404), .A2(KEYINPUT11), .A3(new_n291), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n363), .A2(G68), .ZN(new_n412));
  NAND4_X1  g0212(.A1(new_n407), .A2(new_n410), .A3(new_n411), .A4(new_n412), .ZN(new_n413));
  NAND2_X1  g0213(.A1(new_n401), .A2(new_n413), .ZN(new_n414));
  AOI21_X1  g0214(.A(new_n413), .B1(new_n399), .B2(G190), .ZN(new_n415));
  OAI21_X1  g0215(.A(G200), .B1(new_n393), .B2(new_n394), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n415), .A2(new_n416), .ZN(new_n417));
  AND2_X1   g0217(.A1(new_n414), .A2(new_n417), .ZN(new_n418));
  NAND3_X1  g0218(.A1(new_n344), .A2(G232), .A3(new_n296), .ZN(new_n419));
  INV_X1    g0219(.A(G107), .ZN(new_n420));
  OAI221_X1 g0220(.A(new_n419), .B1(new_n420), .B2(new_n344), .C1(new_n347), .C2(new_n217), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n421), .A2(new_n304), .ZN(new_n422));
  AOI21_X1  g0222(.A(new_n351), .B1(new_n352), .B2(G244), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n422), .A2(new_n423), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n424), .A2(G200), .ZN(new_n425));
  INV_X1    g0225(.A(new_n291), .ZN(new_n426));
  XNOR2_X1  g0226(.A(KEYINPUT15), .B(G87), .ZN(new_n427));
  INV_X1    g0227(.A(KEYINPUT69), .ZN(new_n428));
  OR2_X1    g0228(.A1(new_n427), .A2(new_n428), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n427), .A2(new_n428), .ZN(new_n430));
  NAND4_X1  g0230(.A1(new_n429), .A2(new_n209), .A3(G33), .A4(new_n430), .ZN(new_n431));
  AOI22_X1  g0231(.A1(new_n249), .A2(new_n277), .B1(G20), .B2(G77), .ZN(new_n432));
  AOI21_X1  g0232(.A(new_n426), .B1(new_n431), .B2(new_n432), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n363), .A2(G77), .ZN(new_n434));
  OAI21_X1  g0234(.A(new_n434), .B1(G77), .B2(new_n254), .ZN(new_n435));
  NOR2_X1   g0235(.A1(new_n433), .A2(new_n435), .ZN(new_n436));
  INV_X1    g0236(.A(G190), .ZN(new_n437));
  OAI211_X1 g0237(.A(new_n425), .B(new_n436), .C1(new_n437), .C2(new_n424), .ZN(new_n438));
  INV_X1    g0238(.A(new_n436), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n424), .A2(new_n329), .ZN(new_n440));
  NAND3_X1  g0240(.A1(new_n422), .A2(new_n327), .A3(new_n423), .ZN(new_n441));
  NAND3_X1  g0241(.A1(new_n439), .A2(new_n440), .A3(new_n441), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n438), .A2(new_n442), .ZN(new_n443));
  XOR2_X1   g0243(.A(new_n443), .B(KEYINPUT70), .Z(new_n444));
  AND4_X1   g0244(.A1(new_n343), .A2(new_n383), .A3(new_n418), .A4(new_n444), .ZN(new_n445));
  XNOR2_X1  g0245(.A(KEYINPUT5), .B(G41), .ZN(new_n446));
  NAND3_X1  g0246(.A1(new_n208), .A2(G45), .A3(G274), .ZN(new_n447));
  INV_X1    g0247(.A(new_n447), .ZN(new_n448));
  AND3_X1   g0248(.A1(new_n446), .A2(new_n448), .A3(new_n310), .ZN(new_n449));
  INV_X1    g0249(.A(G45), .ZN(new_n450));
  NOR2_X1   g0250(.A1(new_n450), .A2(G1), .ZN(new_n451));
  AOI21_X1  g0251(.A(new_n304), .B1(new_n451), .B2(new_n446), .ZN(new_n452));
  AOI21_X1  g0252(.A(new_n449), .B1(G270), .B2(new_n452), .ZN(new_n453));
  OAI211_X1 g0253(.A(G264), .B(G1698), .C1(new_n269), .C2(new_n270), .ZN(new_n454));
  OAI211_X1 g0254(.A(G257), .B(new_n296), .C1(new_n269), .C2(new_n270), .ZN(new_n455));
  INV_X1    g0255(.A(G303), .ZN(new_n456));
  OAI211_X1 g0256(.A(new_n454), .B(new_n455), .C1(new_n456), .C2(new_n344), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n457), .A2(new_n304), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n453), .A2(new_n458), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n459), .A2(G169), .ZN(new_n460));
  NOR2_X1   g0260(.A1(new_n262), .A2(G1), .ZN(new_n461));
  NOR2_X1   g0261(.A1(new_n256), .A2(new_n461), .ZN(new_n462));
  OR3_X1    g0262(.A1(new_n254), .A2(KEYINPUT85), .A3(G116), .ZN(new_n463));
  OAI21_X1  g0263(.A(KEYINPUT85), .B1(new_n254), .B2(G116), .ZN(new_n464));
  AOI22_X1  g0264(.A1(new_n462), .A2(G116), .B1(new_n463), .B2(new_n464), .ZN(new_n465));
  INV_X1    g0265(.A(G116), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n466), .A2(G20), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n291), .A2(new_n467), .ZN(new_n468));
  INV_X1    g0268(.A(KEYINPUT86), .ZN(new_n469));
  AOI21_X1  g0269(.A(G20), .B1(G33), .B2(G283), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n262), .A2(G97), .ZN(new_n471));
  AOI21_X1  g0271(.A(new_n469), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  NOR2_X1   g0272(.A1(new_n468), .A2(new_n472), .ZN(new_n473));
  NAND3_X1  g0273(.A1(new_n470), .A2(new_n471), .A3(new_n469), .ZN(new_n474));
  AOI21_X1  g0274(.A(KEYINPUT20), .B1(new_n473), .B2(new_n474), .ZN(new_n475));
  NAND2_X1  g0275(.A1(G33), .A2(G283), .ZN(new_n476));
  INV_X1    g0276(.A(G97), .ZN(new_n477));
  OAI211_X1 g0277(.A(new_n476), .B(new_n209), .C1(G33), .C2(new_n477), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n478), .A2(KEYINPUT86), .ZN(new_n479));
  AOI22_X1  g0279(.A1(new_n255), .A2(new_n226), .B1(G20), .B2(new_n466), .ZN(new_n480));
  NAND4_X1  g0280(.A1(new_n479), .A2(KEYINPUT20), .A3(new_n474), .A4(new_n480), .ZN(new_n481));
  INV_X1    g0281(.A(new_n481), .ZN(new_n482));
  OAI21_X1  g0282(.A(new_n465), .B1(new_n475), .B2(new_n482), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n483), .A2(KEYINPUT87), .ZN(new_n484));
  NAND3_X1  g0284(.A1(new_n479), .A2(new_n474), .A3(new_n480), .ZN(new_n485));
  INV_X1    g0285(.A(KEYINPUT20), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n485), .A2(new_n486), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n487), .A2(new_n481), .ZN(new_n488));
  INV_X1    g0288(.A(KEYINPUT87), .ZN(new_n489));
  NAND3_X1  g0289(.A1(new_n488), .A2(new_n489), .A3(new_n465), .ZN(new_n490));
  AOI21_X1  g0290(.A(new_n460), .B1(new_n484), .B2(new_n490), .ZN(new_n491));
  OAI21_X1  g0291(.A(KEYINPUT21), .B1(new_n491), .B2(KEYINPUT88), .ZN(new_n492));
  AND3_X1   g0292(.A1(new_n488), .A2(new_n489), .A3(new_n465), .ZN(new_n493));
  AOI21_X1  g0293(.A(new_n489), .B1(new_n488), .B2(new_n465), .ZN(new_n494));
  NOR2_X1   g0294(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n459), .A2(G200), .ZN(new_n496));
  OAI211_X1 g0296(.A(new_n495), .B(new_n496), .C1(new_n437), .C2(new_n459), .ZN(new_n497));
  AOI21_X1  g0297(.A(new_n329), .B1(new_n453), .B2(new_n458), .ZN(new_n498));
  OAI21_X1  g0298(.A(new_n498), .B1(new_n493), .B2(new_n494), .ZN(new_n499));
  INV_X1    g0299(.A(KEYINPUT88), .ZN(new_n500));
  INV_X1    g0300(.A(KEYINPUT21), .ZN(new_n501));
  NAND3_X1  g0301(.A1(new_n499), .A2(new_n500), .A3(new_n501), .ZN(new_n502));
  AND3_X1   g0302(.A1(new_n453), .A2(G179), .A3(new_n458), .ZN(new_n503));
  OAI21_X1  g0303(.A(new_n503), .B1(new_n493), .B2(new_n494), .ZN(new_n504));
  AND4_X1   g0304(.A1(new_n492), .A2(new_n497), .A3(new_n502), .A4(new_n504), .ZN(new_n505));
  OAI211_X1 g0305(.A(G244), .B(new_n296), .C1(new_n269), .C2(new_n270), .ZN(new_n506));
  INV_X1    g0306(.A(KEYINPUT4), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  NAND4_X1  g0308(.A1(new_n344), .A2(KEYINPUT4), .A3(G244), .A4(new_n296), .ZN(new_n509));
  NAND3_X1  g0309(.A1(new_n344), .A2(G250), .A3(G1698), .ZN(new_n510));
  NAND4_X1  g0310(.A1(new_n508), .A2(new_n509), .A3(new_n476), .A4(new_n510), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n511), .A2(new_n304), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n446), .A2(new_n451), .ZN(new_n513));
  NAND3_X1  g0313(.A1(new_n513), .A2(G257), .A3(new_n310), .ZN(new_n514));
  NAND3_X1  g0314(.A1(new_n446), .A2(new_n448), .A3(new_n310), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  INV_X1    g0316(.A(new_n516), .ZN(new_n517));
  NAND3_X1  g0317(.A1(new_n512), .A2(new_n437), .A3(new_n517), .ZN(new_n518));
  AOI21_X1  g0318(.A(new_n516), .B1(new_n304), .B2(new_n511), .ZN(new_n519));
  OAI21_X1  g0319(.A(new_n518), .B1(G200), .B2(new_n519), .ZN(new_n520));
  NOR2_X1   g0320(.A1(new_n254), .A2(G97), .ZN(new_n521));
  AOI21_X1  g0321(.A(new_n521), .B1(new_n462), .B2(G97), .ZN(new_n522));
  INV_X1    g0322(.A(new_n522), .ZN(new_n523));
  OAI21_X1  g0323(.A(G107), .B1(new_n273), .B2(new_n274), .ZN(new_n524));
  AND3_X1   g0324(.A1(new_n277), .A2(KEYINPUT81), .A3(G77), .ZN(new_n525));
  AOI21_X1  g0325(.A(KEYINPUT81), .B1(new_n277), .B2(G77), .ZN(new_n526));
  NOR2_X1   g0326(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  XNOR2_X1  g0327(.A(G97), .B(G107), .ZN(new_n528));
  INV_X1    g0328(.A(KEYINPUT6), .ZN(new_n529));
  NOR2_X1   g0329(.A1(new_n529), .A2(new_n477), .ZN(new_n530));
  AOI22_X1  g0330(.A1(new_n528), .A2(new_n529), .B1(new_n420), .B2(new_n530), .ZN(new_n531));
  OAI21_X1  g0331(.A(new_n527), .B1(new_n531), .B2(new_n209), .ZN(new_n532));
  INV_X1    g0332(.A(new_n532), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n524), .A2(new_n533), .ZN(new_n534));
  AOI21_X1  g0334(.A(new_n523), .B1(new_n534), .B2(new_n291), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n520), .A2(new_n535), .ZN(new_n536));
  OAI21_X1  g0336(.A(KEYINPUT76), .B1(new_n288), .B2(new_n286), .ZN(new_n537));
  NAND3_X1  g0337(.A1(new_n537), .A2(new_n268), .A3(new_n272), .ZN(new_n538));
  AOI21_X1  g0338(.A(new_n532), .B1(new_n538), .B2(G107), .ZN(new_n539));
  OAI21_X1  g0339(.A(new_n522), .B1(new_n539), .B2(new_n426), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n512), .A2(new_n517), .ZN(new_n541));
  NAND2_X1  g0341(.A1(new_n541), .A2(new_n329), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n519), .A2(new_n327), .ZN(new_n543));
  NAND3_X1  g0343(.A1(new_n540), .A2(new_n542), .A3(new_n543), .ZN(new_n544));
  INV_X1    g0344(.A(KEYINPUT83), .ZN(new_n545));
  NOR3_X1   g0345(.A1(G87), .A2(G97), .A3(G107), .ZN(new_n546));
  OAI21_X1  g0346(.A(KEYINPUT19), .B1(new_n386), .B2(new_n387), .ZN(new_n547));
  AOI21_X1  g0347(.A(new_n546), .B1(new_n547), .B2(new_n209), .ZN(new_n548));
  OAI211_X1 g0348(.A(new_n209), .B(G68), .C1(new_n269), .C2(new_n270), .ZN(new_n549));
  INV_X1    g0349(.A(KEYINPUT19), .ZN(new_n550));
  OAI21_X1  g0350(.A(new_n550), .B1(new_n360), .B2(new_n477), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n549), .A2(new_n551), .ZN(new_n552));
  OAI21_X1  g0352(.A(new_n545), .B1(new_n548), .B2(new_n552), .ZN(new_n553));
  INV_X1    g0353(.A(new_n546), .ZN(new_n554));
  NAND2_X1  g0354(.A1(G33), .A2(G97), .ZN(new_n555));
  INV_X1    g0355(.A(KEYINPUT74), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  NAND3_X1  g0357(.A1(KEYINPUT74), .A2(G33), .A3(G97), .ZN(new_n558));
  AOI21_X1  g0358(.A(new_n550), .B1(new_n557), .B2(new_n558), .ZN(new_n559));
  OAI21_X1  g0359(.A(new_n554), .B1(new_n559), .B2(G20), .ZN(new_n560));
  AND2_X1   g0360(.A1(new_n549), .A2(new_n551), .ZN(new_n561));
  NAND3_X1  g0361(.A1(new_n560), .A2(new_n561), .A3(KEYINPUT83), .ZN(new_n562));
  NAND3_X1  g0362(.A1(new_n553), .A2(new_n562), .A3(new_n291), .ZN(new_n563));
  AND2_X1   g0363(.A1(new_n429), .A2(new_n430), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n564), .A2(new_n462), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n429), .A2(new_n430), .ZN(new_n566));
  INV_X1    g0366(.A(new_n254), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  NAND3_X1  g0368(.A1(new_n563), .A2(new_n565), .A3(new_n568), .ZN(new_n569));
  OAI211_X1 g0369(.A(G244), .B(G1698), .C1(new_n269), .C2(new_n270), .ZN(new_n570));
  OAI211_X1 g0370(.A(G238), .B(new_n296), .C1(new_n269), .C2(new_n270), .ZN(new_n571));
  NAND2_X1  g0371(.A1(G33), .A2(G116), .ZN(new_n572));
  NAND3_X1  g0372(.A1(new_n570), .A2(new_n571), .A3(new_n572), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n573), .A2(new_n304), .ZN(new_n574));
  INV_X1    g0374(.A(KEYINPUT82), .ZN(new_n575));
  NOR2_X1   g0375(.A1(new_n447), .A2(new_n575), .ZN(new_n576));
  INV_X1    g0376(.A(new_n576), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n447), .A2(new_n575), .ZN(new_n578));
  NOR2_X1   g0378(.A1(new_n451), .A2(new_n219), .ZN(new_n579));
  AOI22_X1  g0379(.A1(new_n577), .A2(new_n578), .B1(new_n579), .B2(new_n310), .ZN(new_n580));
  AND3_X1   g0380(.A1(new_n574), .A2(new_n327), .A3(new_n580), .ZN(new_n581));
  AOI21_X1  g0381(.A(G169), .B1(new_n574), .B2(new_n580), .ZN(new_n582));
  NOR2_X1   g0382(.A1(new_n581), .A2(new_n582), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n569), .A2(new_n583), .ZN(new_n584));
  NAND3_X1  g0384(.A1(new_n574), .A2(new_n437), .A3(new_n580), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n208), .A2(G45), .ZN(new_n586));
  NAND3_X1  g0386(.A1(new_n310), .A2(G250), .A3(new_n586), .ZN(new_n587));
  INV_X1    g0387(.A(new_n578), .ZN(new_n588));
  OAI21_X1  g0388(.A(new_n587), .B1(new_n588), .B2(new_n576), .ZN(new_n589));
  AOI21_X1  g0389(.A(new_n589), .B1(new_n304), .B2(new_n573), .ZN(new_n590));
  OAI21_X1  g0390(.A(new_n585), .B1(new_n590), .B2(G200), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n462), .A2(G87), .ZN(new_n592));
  NAND4_X1  g0392(.A1(new_n591), .A2(new_n568), .A3(new_n563), .A4(new_n592), .ZN(new_n593));
  NAND4_X1  g0393(.A1(new_n536), .A2(new_n544), .A3(new_n584), .A4(new_n593), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n594), .A2(KEYINPUT84), .ZN(new_n595));
  OAI211_X1 g0395(.A(new_n209), .B(G87), .C1(new_n269), .C2(new_n270), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n596), .A2(KEYINPUT22), .ZN(new_n597));
  INV_X1    g0397(.A(KEYINPUT22), .ZN(new_n598));
  NAND4_X1  g0398(.A1(new_n344), .A2(new_n598), .A3(new_n209), .A4(G87), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n597), .A2(new_n599), .ZN(new_n600));
  INV_X1    g0400(.A(KEYINPUT24), .ZN(new_n601));
  NOR2_X1   g0401(.A1(new_n572), .A2(G20), .ZN(new_n602));
  INV_X1    g0402(.A(KEYINPUT23), .ZN(new_n603));
  OAI21_X1  g0403(.A(new_n603), .B1(new_n209), .B2(G107), .ZN(new_n604));
  NAND3_X1  g0404(.A1(new_n420), .A2(KEYINPUT23), .A3(G20), .ZN(new_n605));
  AOI21_X1  g0405(.A(new_n602), .B1(new_n604), .B2(new_n605), .ZN(new_n606));
  AND3_X1   g0406(.A1(new_n600), .A2(new_n601), .A3(new_n606), .ZN(new_n607));
  AOI21_X1  g0407(.A(new_n601), .B1(new_n600), .B2(new_n606), .ZN(new_n608));
  OAI21_X1  g0408(.A(new_n291), .B1(new_n607), .B2(new_n608), .ZN(new_n609));
  INV_X1    g0409(.A(KEYINPUT25), .ZN(new_n610));
  NOR3_X1   g0410(.A1(new_n254), .A2(new_n610), .A3(G107), .ZN(new_n611));
  INV_X1    g0411(.A(new_n611), .ZN(new_n612));
  OAI21_X1  g0412(.A(new_n610), .B1(new_n254), .B2(G107), .ZN(new_n613));
  AOI22_X1  g0413(.A1(new_n462), .A2(G107), .B1(new_n612), .B2(new_n613), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n609), .A2(new_n614), .ZN(new_n615));
  OAI211_X1 g0415(.A(G250), .B(new_n296), .C1(new_n269), .C2(new_n270), .ZN(new_n616));
  OAI211_X1 g0416(.A(G257), .B(G1698), .C1(new_n269), .C2(new_n270), .ZN(new_n617));
  NAND2_X1  g0417(.A1(G33), .A2(G294), .ZN(new_n618));
  NAND3_X1  g0418(.A1(new_n616), .A2(new_n617), .A3(new_n618), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n619), .A2(new_n304), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n452), .A2(G264), .ZN(new_n621));
  NAND3_X1  g0421(.A1(new_n620), .A2(new_n621), .A3(new_n515), .ZN(new_n622));
  INV_X1    g0422(.A(KEYINPUT89), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  AOI22_X1  g0424(.A1(new_n304), .A2(new_n619), .B1(new_n452), .B2(G264), .ZN(new_n625));
  NAND3_X1  g0425(.A1(new_n625), .A2(KEYINPUT89), .A3(new_n515), .ZN(new_n626));
  AND3_X1   g0426(.A1(new_n624), .A2(G169), .A3(new_n626), .ZN(new_n627));
  OAI21_X1  g0427(.A(KEYINPUT90), .B1(new_n622), .B2(new_n327), .ZN(new_n628));
  INV_X1    g0428(.A(KEYINPUT90), .ZN(new_n629));
  NAND4_X1  g0429(.A1(new_n625), .A2(new_n629), .A3(G179), .A4(new_n515), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n628), .A2(new_n630), .ZN(new_n631));
  OAI21_X1  g0431(.A(new_n615), .B1(new_n627), .B2(new_n631), .ZN(new_n632));
  AOI21_X1  g0432(.A(G190), .B1(new_n624), .B2(new_n626), .ZN(new_n633));
  INV_X1    g0433(.A(new_n622), .ZN(new_n634));
  NOR2_X1   g0434(.A1(new_n634), .A2(G200), .ZN(new_n635));
  OAI211_X1 g0435(.A(new_n609), .B(new_n614), .C1(new_n633), .C2(new_n635), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n632), .A2(new_n636), .ZN(new_n637));
  INV_X1    g0437(.A(new_n594), .ZN(new_n638));
  INV_X1    g0438(.A(KEYINPUT84), .ZN(new_n639));
  AOI21_X1  g0439(.A(new_n637), .B1(new_n638), .B2(new_n639), .ZN(new_n640));
  NAND4_X1  g0440(.A1(new_n445), .A2(new_n505), .A3(new_n595), .A4(new_n640), .ZN(new_n641));
  XOR2_X1   g0441(.A(new_n641), .B(KEYINPUT91), .Z(G372));
  INV_X1    g0442(.A(KEYINPUT94), .ZN(new_n643));
  XNOR2_X1  g0443(.A(new_n632), .B(KEYINPUT93), .ZN(new_n644));
  NAND3_X1  g0444(.A1(new_n492), .A2(new_n502), .A3(new_n504), .ZN(new_n645));
  OAI21_X1  g0445(.A(new_n643), .B1(new_n644), .B2(new_n645), .ZN(new_n646));
  INV_X1    g0446(.A(KEYINPUT93), .ZN(new_n647));
  XNOR2_X1  g0447(.A(new_n632), .B(new_n647), .ZN(new_n648));
  INV_X1    g0448(.A(new_n645), .ZN(new_n649));
  NAND3_X1  g0449(.A1(new_n648), .A2(new_n649), .A3(KEYINPUT94), .ZN(new_n650));
  INV_X1    g0450(.A(new_n633), .ZN(new_n651));
  INV_X1    g0451(.A(new_n635), .ZN(new_n652));
  AOI21_X1  g0452(.A(new_n615), .B1(new_n651), .B2(new_n652), .ZN(new_n653));
  OAI21_X1  g0453(.A(KEYINPUT92), .B1(new_n594), .B2(new_n653), .ZN(new_n654));
  NOR2_X1   g0454(.A1(new_n594), .A2(new_n653), .ZN(new_n655));
  INV_X1    g0455(.A(KEYINPUT92), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  NAND4_X1  g0457(.A1(new_n646), .A2(new_n650), .A3(new_n654), .A4(new_n657), .ZN(new_n658));
  INV_X1    g0458(.A(new_n584), .ZN(new_n659));
  INV_X1    g0459(.A(KEYINPUT26), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n584), .A2(new_n593), .ZN(new_n661));
  OAI21_X1  g0461(.A(new_n660), .B1(new_n661), .B2(new_n544), .ZN(new_n662));
  AND3_X1   g0462(.A1(new_n540), .A2(new_n543), .A3(new_n542), .ZN(new_n663));
  NAND4_X1  g0463(.A1(new_n663), .A2(KEYINPUT26), .A3(new_n584), .A4(new_n593), .ZN(new_n664));
  AOI21_X1  g0464(.A(new_n659), .B1(new_n662), .B2(new_n664), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n658), .A2(new_n665), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n445), .A2(new_n666), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n377), .A2(new_n382), .ZN(new_n668));
  AND2_X1   g0468(.A1(new_n332), .A2(new_n340), .ZN(new_n669));
  NAND3_X1  g0469(.A1(new_n326), .A2(new_n341), .A3(new_n417), .ZN(new_n670));
  INV_X1    g0470(.A(new_n442), .ZN(new_n671));
  AOI21_X1  g0471(.A(new_n671), .B1(new_n413), .B2(new_n401), .ZN(new_n672));
  OAI21_X1  g0472(.A(new_n669), .B1(new_n670), .B2(new_n672), .ZN(new_n673));
  AOI21_X1  g0473(.A(new_n368), .B1(new_n668), .B2(new_n673), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n667), .A2(new_n674), .ZN(G369));
  NAND3_X1  g0475(.A1(new_n208), .A2(new_n209), .A3(G13), .ZN(new_n676));
  OR2_X1    g0476(.A1(new_n676), .A2(KEYINPUT27), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n676), .A2(KEYINPUT27), .ZN(new_n678));
  NAND3_X1  g0478(.A1(new_n677), .A2(G213), .A3(new_n678), .ZN(new_n679));
  INV_X1    g0479(.A(G343), .ZN(new_n680));
  NOR2_X1   g0480(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  INV_X1    g0481(.A(new_n681), .ZN(new_n682));
  NOR2_X1   g0482(.A1(new_n495), .A2(new_n682), .ZN(new_n683));
  MUX2_X1   g0483(.A(new_n505), .B(new_n645), .S(new_n683), .Z(new_n684));
  AND2_X1   g0484(.A1(new_n684), .A2(G330), .ZN(new_n685));
  AOI21_X1  g0485(.A(new_n682), .B1(new_n609), .B2(new_n614), .ZN(new_n686));
  OAI22_X1  g0486(.A1(new_n637), .A2(new_n686), .B1(new_n632), .B2(new_n682), .ZN(new_n687));
  AND2_X1   g0487(.A1(new_n685), .A2(new_n687), .ZN(new_n688));
  NOR2_X1   g0488(.A1(new_n649), .A2(new_n681), .ZN(new_n689));
  INV_X1    g0489(.A(new_n637), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n644), .A2(new_n682), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  OR2_X1    g0493(.A1(new_n688), .A2(new_n693), .ZN(G399));
  INV_X1    g0494(.A(new_n212), .ZN(new_n695));
  NOR2_X1   g0495(.A1(new_n695), .A2(G41), .ZN(new_n696));
  INV_X1    g0496(.A(new_n696), .ZN(new_n697));
  NOR2_X1   g0497(.A1(new_n554), .A2(G116), .ZN(new_n698));
  NAND3_X1  g0498(.A1(new_n697), .A2(G1), .A3(new_n698), .ZN(new_n699));
  INV_X1    g0499(.A(new_n230), .ZN(new_n700));
  OAI21_X1  g0500(.A(new_n699), .B1(new_n700), .B2(new_n697), .ZN(new_n701));
  XNOR2_X1  g0501(.A(new_n701), .B(KEYINPUT95), .ZN(new_n702));
  XNOR2_X1  g0502(.A(new_n702), .B(KEYINPUT28), .ZN(new_n703));
  INV_X1    g0503(.A(KEYINPUT97), .ZN(new_n704));
  NAND4_X1  g0504(.A1(new_n640), .A2(new_n505), .A3(new_n595), .A4(new_n682), .ZN(new_n705));
  AND3_X1   g0505(.A1(new_n625), .A2(new_n574), .A3(new_n580), .ZN(new_n706));
  NAND3_X1  g0506(.A1(new_n706), .A2(new_n503), .A3(new_n519), .ZN(new_n707));
  INV_X1    g0507(.A(KEYINPUT30), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n707), .A2(new_n708), .ZN(new_n709));
  NAND4_X1  g0509(.A1(new_n706), .A2(new_n503), .A3(KEYINPUT30), .A4(new_n519), .ZN(new_n710));
  NAND2_X1  g0510(.A1(new_n709), .A2(new_n710), .ZN(new_n711));
  NAND2_X1  g0511(.A1(new_n574), .A2(new_n580), .ZN(new_n712));
  NAND3_X1  g0512(.A1(new_n459), .A2(new_n327), .A3(new_n712), .ZN(new_n713));
  OAI21_X1  g0513(.A(KEYINPUT96), .B1(new_n634), .B2(new_n519), .ZN(new_n714));
  INV_X1    g0514(.A(KEYINPUT96), .ZN(new_n715));
  NAND3_X1  g0515(.A1(new_n541), .A2(new_n715), .A3(new_n622), .ZN(new_n716));
  AOI21_X1  g0516(.A(new_n713), .B1(new_n714), .B2(new_n716), .ZN(new_n717));
  OAI211_X1 g0517(.A(KEYINPUT31), .B(new_n681), .C1(new_n711), .C2(new_n717), .ZN(new_n718));
  INV_X1    g0518(.A(new_n718), .ZN(new_n719));
  INV_X1    g0519(.A(new_n713), .ZN(new_n720));
  NOR3_X1   g0520(.A1(new_n634), .A2(new_n519), .A3(KEYINPUT96), .ZN(new_n721));
  AOI21_X1  g0521(.A(new_n715), .B1(new_n541), .B2(new_n622), .ZN(new_n722));
  OAI21_X1  g0522(.A(new_n720), .B1(new_n721), .B2(new_n722), .ZN(new_n723));
  NAND3_X1  g0523(.A1(new_n723), .A2(new_n709), .A3(new_n710), .ZN(new_n724));
  AOI21_X1  g0524(.A(KEYINPUT31), .B1(new_n724), .B2(new_n681), .ZN(new_n725));
  NOR2_X1   g0525(.A1(new_n719), .A2(new_n725), .ZN(new_n726));
  NAND2_X1  g0526(.A1(new_n705), .A2(new_n726), .ZN(new_n727));
  AOI21_X1  g0527(.A(new_n704), .B1(new_n727), .B2(G330), .ZN(new_n728));
  INV_X1    g0528(.A(G330), .ZN(new_n729));
  AOI211_X1 g0529(.A(KEYINPUT97), .B(new_n729), .C1(new_n705), .C2(new_n726), .ZN(new_n730));
  NOR2_X1   g0530(.A1(new_n728), .A2(new_n730), .ZN(new_n731));
  AOI21_X1  g0531(.A(new_n681), .B1(new_n658), .B2(new_n665), .ZN(new_n732));
  OR2_X1    g0532(.A1(new_n732), .A2(KEYINPUT29), .ZN(new_n733));
  NAND4_X1  g0533(.A1(new_n492), .A2(new_n502), .A3(new_n504), .A4(new_n632), .ZN(new_n734));
  NAND2_X1  g0534(.A1(new_n655), .A2(new_n734), .ZN(new_n735));
  NAND2_X1  g0535(.A1(new_n735), .A2(new_n665), .ZN(new_n736));
  AOI21_X1  g0536(.A(KEYINPUT98), .B1(new_n736), .B2(new_n682), .ZN(new_n737));
  INV_X1    g0537(.A(KEYINPUT98), .ZN(new_n738));
  AOI211_X1 g0538(.A(new_n738), .B(new_n681), .C1(new_n735), .C2(new_n665), .ZN(new_n739));
  OAI21_X1  g0539(.A(KEYINPUT29), .B1(new_n737), .B2(new_n739), .ZN(new_n740));
  AOI21_X1  g0540(.A(new_n731), .B1(new_n733), .B2(new_n740), .ZN(new_n741));
  OAI21_X1  g0541(.A(new_n703), .B1(new_n741), .B2(G1), .ZN(G364));
  INV_X1    g0542(.A(G13), .ZN(new_n743));
  NOR2_X1   g0543(.A1(new_n743), .A2(G20), .ZN(new_n744));
  AOI21_X1  g0544(.A(new_n208), .B1(new_n744), .B2(G45), .ZN(new_n745));
  INV_X1    g0545(.A(new_n745), .ZN(new_n746));
  NOR2_X1   g0546(.A1(new_n696), .A2(new_n746), .ZN(new_n747));
  NOR2_X1   g0547(.A1(new_n685), .A2(new_n747), .ZN(new_n748));
  OAI21_X1  g0548(.A(new_n748), .B1(G330), .B2(new_n684), .ZN(new_n749));
  XNOR2_X1  g0549(.A(new_n747), .B(KEYINPUT99), .ZN(new_n750));
  INV_X1    g0550(.A(new_n750), .ZN(new_n751));
  AOI21_X1  g0551(.A(new_n226), .B1(G20), .B2(new_n329), .ZN(new_n752));
  INV_X1    g0552(.A(new_n752), .ZN(new_n753));
  NOR2_X1   g0553(.A1(new_n327), .A2(new_n320), .ZN(new_n754));
  NOR2_X1   g0554(.A1(new_n209), .A2(G190), .ZN(new_n755));
  NAND2_X1  g0555(.A1(new_n754), .A2(new_n755), .ZN(new_n756));
  OAI21_X1  g0556(.A(new_n344), .B1(new_n756), .B2(new_n202), .ZN(new_n757));
  INV_X1    g0557(.A(new_n755), .ZN(new_n758));
  NOR3_X1   g0558(.A1(new_n758), .A2(G179), .A3(new_n320), .ZN(new_n759));
  INV_X1    g0559(.A(new_n759), .ZN(new_n760));
  NOR2_X1   g0560(.A1(new_n209), .A2(new_n437), .ZN(new_n761));
  NAND2_X1  g0561(.A1(new_n754), .A2(new_n761), .ZN(new_n762));
  OAI22_X1  g0562(.A1(new_n760), .A2(new_n420), .B1(new_n229), .B2(new_n762), .ZN(new_n763));
  INV_X1    g0563(.A(new_n761), .ZN(new_n764));
  NOR3_X1   g0564(.A1(new_n764), .A2(new_n320), .A3(G179), .ZN(new_n765));
  AOI211_X1 g0565(.A(new_n757), .B(new_n763), .C1(G87), .C2(new_n765), .ZN(new_n766));
  AND3_X1   g0566(.A1(new_n327), .A2(new_n320), .A3(KEYINPUT101), .ZN(new_n767));
  AOI21_X1  g0567(.A(KEYINPUT101), .B1(new_n327), .B2(new_n320), .ZN(new_n768));
  NOR2_X1   g0568(.A1(new_n767), .A2(new_n768), .ZN(new_n769));
  NOR2_X1   g0569(.A1(new_n769), .A2(new_n758), .ZN(new_n770));
  NAND2_X1  g0570(.A1(new_n770), .A2(G159), .ZN(new_n771));
  XOR2_X1   g0571(.A(new_n771), .B(KEYINPUT32), .Z(new_n772));
  INV_X1    g0572(.A(new_n769), .ZN(new_n773));
  AOI21_X1  g0573(.A(new_n209), .B1(new_n773), .B2(G190), .ZN(new_n774));
  INV_X1    g0574(.A(new_n774), .ZN(new_n775));
  NAND2_X1  g0575(.A1(new_n775), .A2(G97), .ZN(new_n776));
  NOR2_X1   g0576(.A1(new_n327), .A2(G200), .ZN(new_n777));
  NAND2_X1  g0577(.A1(new_n761), .A2(new_n777), .ZN(new_n778));
  NAND2_X1  g0578(.A1(new_n755), .A2(new_n777), .ZN(new_n779));
  OAI22_X1  g0579(.A1(new_n778), .A2(new_n201), .B1(new_n779), .B2(new_n346), .ZN(new_n780));
  XOR2_X1   g0580(.A(new_n780), .B(KEYINPUT100), .Z(new_n781));
  NAND4_X1  g0581(.A1(new_n766), .A2(new_n772), .A3(new_n776), .A4(new_n781), .ZN(new_n782));
  INV_X1    g0582(.A(new_n756), .ZN(new_n783));
  NOR2_X1   g0583(.A1(KEYINPUT33), .A2(G317), .ZN(new_n784));
  AND2_X1   g0584(.A1(KEYINPUT33), .A2(G317), .ZN(new_n785));
  OAI21_X1  g0585(.A(new_n783), .B1(new_n784), .B2(new_n785), .ZN(new_n786));
  INV_X1    g0586(.A(new_n765), .ZN(new_n787));
  OAI21_X1  g0587(.A(new_n786), .B1(new_n787), .B2(new_n456), .ZN(new_n788));
  AOI21_X1  g0588(.A(new_n788), .B1(G283), .B2(new_n759), .ZN(new_n789));
  INV_X1    g0589(.A(G311), .ZN(new_n790));
  OAI21_X1  g0590(.A(new_n271), .B1(new_n779), .B2(new_n790), .ZN(new_n791));
  INV_X1    g0591(.A(new_n778), .ZN(new_n792));
  AND2_X1   g0592(.A1(new_n792), .A2(G322), .ZN(new_n793));
  INV_X1    g0593(.A(new_n762), .ZN(new_n794));
  AOI211_X1 g0594(.A(new_n791), .B(new_n793), .C1(G326), .C2(new_n794), .ZN(new_n795));
  NAND2_X1  g0595(.A1(new_n775), .A2(G294), .ZN(new_n796));
  NAND2_X1  g0596(.A1(new_n770), .A2(G329), .ZN(new_n797));
  NAND4_X1  g0597(.A1(new_n789), .A2(new_n795), .A3(new_n796), .A4(new_n797), .ZN(new_n798));
  AOI21_X1  g0598(.A(new_n753), .B1(new_n782), .B2(new_n798), .ZN(new_n799));
  NOR2_X1   g0599(.A1(G13), .A2(G33), .ZN(new_n800));
  INV_X1    g0600(.A(new_n800), .ZN(new_n801));
  NOR2_X1   g0601(.A1(new_n801), .A2(G20), .ZN(new_n802));
  NOR2_X1   g0602(.A1(new_n802), .A2(new_n752), .ZN(new_n803));
  NOR2_X1   g0603(.A1(new_n695), .A2(new_n271), .ZN(new_n804));
  AOI22_X1  g0604(.A1(new_n804), .A2(G355), .B1(new_n466), .B2(new_n695), .ZN(new_n805));
  AND2_X1   g0605(.A1(new_n243), .A2(G45), .ZN(new_n806));
  NOR2_X1   g0606(.A1(new_n695), .A2(new_n344), .ZN(new_n807));
  OAI21_X1  g0607(.A(new_n807), .B1(new_n700), .B2(G45), .ZN(new_n808));
  OAI21_X1  g0608(.A(new_n805), .B1(new_n806), .B2(new_n808), .ZN(new_n809));
  AOI211_X1 g0609(.A(new_n751), .B(new_n799), .C1(new_n803), .C2(new_n809), .ZN(new_n810));
  XOR2_X1   g0610(.A(new_n810), .B(KEYINPUT102), .Z(new_n811));
  XOR2_X1   g0611(.A(new_n802), .B(KEYINPUT103), .Z(new_n812));
  OAI21_X1  g0612(.A(new_n811), .B1(new_n684), .B2(new_n812), .ZN(new_n813));
  AND2_X1   g0613(.A1(new_n749), .A2(new_n813), .ZN(new_n814));
  INV_X1    g0614(.A(new_n814), .ZN(G396));
  NOR2_X1   g0615(.A1(new_n752), .A2(new_n800), .ZN(new_n816));
  INV_X1    g0616(.A(new_n816), .ZN(new_n817));
  OAI21_X1  g0617(.A(new_n750), .B1(G77), .B2(new_n817), .ZN(new_n818));
  INV_X1    g0618(.A(new_n779), .ZN(new_n819));
  AOI22_X1  g0619(.A1(G143), .A2(new_n792), .B1(new_n819), .B2(G159), .ZN(new_n820));
  INV_X1    g0620(.A(G137), .ZN(new_n821));
  INV_X1    g0621(.A(G150), .ZN(new_n822));
  OAI221_X1 g0622(.A(new_n820), .B1(new_n821), .B2(new_n762), .C1(new_n822), .C2(new_n756), .ZN(new_n823));
  XOR2_X1   g0623(.A(new_n823), .B(KEYINPUT105), .Z(new_n824));
  XNOR2_X1  g0624(.A(new_n824), .B(KEYINPUT104), .ZN(new_n825));
  OR2_X1    g0625(.A1(new_n825), .A2(KEYINPUT34), .ZN(new_n826));
  NAND2_X1  g0626(.A1(new_n825), .A2(KEYINPUT34), .ZN(new_n827));
  NOR2_X1   g0627(.A1(new_n774), .A2(new_n201), .ZN(new_n828));
  OAI221_X1 g0628(.A(new_n344), .B1(new_n760), .B2(new_n202), .C1(new_n229), .C2(new_n787), .ZN(new_n829));
  AOI211_X1 g0629(.A(new_n828), .B(new_n829), .C1(G132), .C2(new_n770), .ZN(new_n830));
  NAND3_X1  g0630(.A1(new_n826), .A2(new_n827), .A3(new_n830), .ZN(new_n831));
  OAI22_X1  g0631(.A1(new_n760), .A2(new_n218), .B1(new_n779), .B2(new_n466), .ZN(new_n832));
  AOI211_X1 g0632(.A(new_n344), .B(new_n832), .C1(G294), .C2(new_n792), .ZN(new_n833));
  NAND2_X1  g0633(.A1(new_n770), .A2(G311), .ZN(new_n834));
  INV_X1    g0634(.A(G283), .ZN(new_n835));
  OAI22_X1  g0635(.A1(new_n762), .A2(new_n456), .B1(new_n756), .B2(new_n835), .ZN(new_n836));
  AOI21_X1  g0636(.A(new_n836), .B1(G107), .B2(new_n765), .ZN(new_n837));
  NAND4_X1  g0637(.A1(new_n833), .A2(new_n776), .A3(new_n834), .A4(new_n837), .ZN(new_n838));
  AOI21_X1  g0638(.A(new_n753), .B1(new_n831), .B2(new_n838), .ZN(new_n839));
  NOR2_X1   g0639(.A1(new_n442), .A2(new_n681), .ZN(new_n840));
  OAI21_X1  g0640(.A(new_n438), .B1(new_n436), .B2(new_n682), .ZN(new_n841));
  AOI21_X1  g0641(.A(new_n840), .B1(new_n841), .B2(new_n442), .ZN(new_n842));
  INV_X1    g0642(.A(new_n842), .ZN(new_n843));
  AOI211_X1 g0643(.A(new_n818), .B(new_n839), .C1(new_n800), .C2(new_n843), .ZN(new_n844));
  INV_X1    g0644(.A(new_n844), .ZN(new_n845));
  NOR2_X1   g0645(.A1(new_n732), .A2(new_n842), .ZN(new_n846));
  INV_X1    g0646(.A(new_n846), .ZN(new_n847));
  NAND3_X1  g0647(.A1(new_n666), .A2(new_n682), .A3(new_n842), .ZN(new_n848));
  NAND2_X1  g0648(.A1(new_n847), .A2(new_n848), .ZN(new_n849));
  INV_X1    g0649(.A(KEYINPUT106), .ZN(new_n850));
  INV_X1    g0650(.A(new_n731), .ZN(new_n851));
  NAND3_X1  g0651(.A1(new_n849), .A2(new_n850), .A3(new_n851), .ZN(new_n852));
  OAI221_X1 g0652(.A(new_n852), .B1(new_n851), .B2(new_n849), .C1(new_n696), .C2(new_n746), .ZN(new_n853));
  AOI21_X1  g0653(.A(new_n850), .B1(new_n849), .B2(new_n851), .ZN(new_n854));
  OAI21_X1  g0654(.A(new_n845), .B1(new_n853), .B2(new_n854), .ZN(G384));
  NAND2_X1  g0655(.A1(new_n227), .A2(G116), .ZN(new_n856));
  INV_X1    g0656(.A(new_n531), .ZN(new_n857));
  AOI21_X1  g0657(.A(new_n856), .B1(new_n857), .B2(KEYINPUT35), .ZN(new_n858));
  OAI21_X1  g0658(.A(new_n858), .B1(KEYINPUT35), .B2(new_n857), .ZN(new_n859));
  XNOR2_X1  g0659(.A(new_n859), .B(KEYINPUT36), .ZN(new_n860));
  OAI21_X1  g0660(.A(G77), .B1(new_n201), .B2(new_n202), .ZN(new_n861));
  OAI22_X1  g0661(.A1(new_n700), .A2(new_n861), .B1(G50), .B2(new_n202), .ZN(new_n862));
  NAND3_X1  g0662(.A1(new_n862), .A2(G1), .A3(new_n743), .ZN(new_n863));
  NAND2_X1  g0663(.A1(new_n860), .A2(new_n863), .ZN(new_n864));
  XNOR2_X1  g0664(.A(new_n864), .B(KEYINPUT107), .ZN(new_n865));
  OAI21_X1  g0665(.A(new_n278), .B1(new_n287), .B2(new_n289), .ZN(new_n866));
  NAND2_X1  g0666(.A1(new_n866), .A2(new_n280), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n292), .A2(new_n867), .ZN(new_n868));
  AOI21_X1  g0668(.A(new_n679), .B1(new_n868), .B2(new_n335), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n342), .A2(new_n869), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n317), .A2(new_n321), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n871), .A2(KEYINPUT80), .ZN(new_n872));
  NAND3_X1  g0672(.A1(new_n317), .A2(new_n294), .A3(new_n321), .ZN(new_n873));
  AOI21_X1  g0673(.A(new_n338), .B1(new_n872), .B2(new_n873), .ZN(new_n874));
  AOI22_X1  g0674(.A1(new_n868), .A2(new_n335), .B1(new_n331), .B2(new_n679), .ZN(new_n875));
  OAI21_X1  g0675(.A(KEYINPUT37), .B1(new_n874), .B2(new_n875), .ZN(new_n876));
  INV_X1    g0676(.A(new_n679), .ZN(new_n877));
  OAI21_X1  g0677(.A(new_n338), .B1(new_n333), .B2(new_n877), .ZN(new_n878));
  INV_X1    g0678(.A(KEYINPUT37), .ZN(new_n879));
  NAND3_X1  g0679(.A1(new_n324), .A2(new_n878), .A3(new_n879), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n876), .A2(new_n880), .ZN(new_n881));
  AOI21_X1  g0681(.A(KEYINPUT38), .B1(new_n870), .B2(new_n881), .ZN(new_n882));
  INV_X1    g0682(.A(new_n882), .ZN(new_n883));
  NAND3_X1  g0683(.A1(new_n870), .A2(KEYINPUT38), .A3(new_n881), .ZN(new_n884));
  NAND3_X1  g0684(.A1(new_n883), .A2(KEYINPUT39), .A3(new_n884), .ZN(new_n885));
  INV_X1    g0685(.A(KEYINPUT39), .ZN(new_n886));
  INV_X1    g0686(.A(KEYINPUT38), .ZN(new_n887));
  AOI221_X4 g0687(.A(new_n887), .B1(new_n876), .B2(new_n880), .C1(new_n342), .C2(new_n869), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n338), .A2(new_n877), .ZN(new_n889));
  INV_X1    g0689(.A(new_n889), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n342), .A2(new_n890), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n889), .A2(KEYINPUT109), .ZN(new_n892));
  NAND4_X1  g0692(.A1(new_n892), .A2(new_n324), .A3(new_n878), .A4(KEYINPUT37), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n281), .A2(new_n292), .ZN(new_n894));
  AOI22_X1  g0694(.A1(new_n894), .A2(new_n335), .B1(new_n331), .B2(new_n679), .ZN(new_n895));
  INV_X1    g0695(.A(KEYINPUT109), .ZN(new_n896));
  AOI21_X1  g0696(.A(new_n896), .B1(new_n338), .B2(new_n877), .ZN(new_n897));
  OAI22_X1  g0697(.A1(new_n874), .A2(new_n895), .B1(new_n897), .B2(new_n879), .ZN(new_n898));
  AND2_X1   g0698(.A1(new_n893), .A2(new_n898), .ZN(new_n899));
  AOI21_X1  g0699(.A(KEYINPUT38), .B1(new_n891), .B2(new_n899), .ZN(new_n900));
  OAI21_X1  g0700(.A(new_n886), .B1(new_n888), .B2(new_n900), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n885), .A2(new_n901), .ZN(new_n902));
  NOR2_X1   g0702(.A1(new_n414), .A2(new_n681), .ZN(new_n903));
  INV_X1    g0703(.A(new_n903), .ZN(new_n904));
  OAI22_X1  g0704(.A1(new_n902), .A2(new_n904), .B1(new_n669), .B2(new_n877), .ZN(new_n905));
  NOR2_X1   g0705(.A1(new_n888), .A2(new_n882), .ZN(new_n906));
  INV_X1    g0706(.A(new_n906), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n413), .A2(new_n681), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n908), .A2(KEYINPUT108), .ZN(new_n909));
  INV_X1    g0709(.A(KEYINPUT108), .ZN(new_n910));
  NAND3_X1  g0710(.A1(new_n413), .A2(new_n910), .A3(new_n681), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n909), .A2(new_n911), .ZN(new_n912));
  AOI221_X4 g0712(.A(new_n912), .B1(new_n416), .B2(new_n415), .C1(new_n401), .C2(new_n413), .ZN(new_n913));
  AND3_X1   g0713(.A1(new_n401), .A2(new_n413), .A3(new_n681), .ZN(new_n914));
  NOR2_X1   g0714(.A1(new_n913), .A2(new_n914), .ZN(new_n915));
  INV_X1    g0715(.A(new_n840), .ZN(new_n916));
  AOI21_X1  g0716(.A(new_n915), .B1(new_n848), .B2(new_n916), .ZN(new_n917));
  AOI21_X1  g0717(.A(new_n905), .B1(new_n907), .B2(new_n917), .ZN(new_n918));
  OAI211_X1 g0718(.A(new_n445), .B(new_n740), .C1(new_n732), .C2(KEYINPUT29), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n919), .A2(new_n674), .ZN(new_n920));
  XOR2_X1   g0720(.A(new_n918), .B(new_n920), .Z(new_n921));
  INV_X1    g0721(.A(KEYINPUT40), .ZN(new_n922));
  OAI21_X1  g0722(.A(new_n842), .B1(new_n913), .B2(new_n914), .ZN(new_n923));
  AOI211_X1 g0723(.A(new_n922), .B(new_n923), .C1(new_n705), .C2(new_n726), .ZN(new_n924));
  OAI21_X1  g0724(.A(KEYINPUT110), .B1(new_n888), .B2(new_n900), .ZN(new_n925));
  INV_X1    g0725(.A(KEYINPUT110), .ZN(new_n926));
  NAND2_X1  g0726(.A1(new_n893), .A2(new_n898), .ZN(new_n927));
  AOI21_X1  g0727(.A(new_n927), .B1(new_n342), .B2(new_n890), .ZN(new_n928));
  OAI211_X1 g0728(.A(new_n884), .B(new_n926), .C1(new_n928), .C2(KEYINPUT38), .ZN(new_n929));
  NAND3_X1  g0729(.A1(new_n924), .A2(new_n925), .A3(new_n929), .ZN(new_n930));
  INV_X1    g0730(.A(new_n923), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n727), .A2(new_n931), .ZN(new_n932));
  OAI21_X1  g0732(.A(new_n922), .B1(new_n906), .B2(new_n932), .ZN(new_n933));
  AND2_X1   g0733(.A1(new_n930), .A2(new_n933), .ZN(new_n934));
  NAND3_X1  g0734(.A1(new_n934), .A2(new_n445), .A3(new_n727), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n935), .A2(G330), .ZN(new_n936));
  AOI21_X1  g0736(.A(new_n934), .B1(new_n445), .B2(new_n727), .ZN(new_n937));
  OR2_X1    g0737(.A1(new_n936), .A2(new_n937), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n921), .A2(new_n938), .ZN(new_n939));
  OAI21_X1  g0739(.A(new_n939), .B1(new_n208), .B2(new_n744), .ZN(new_n940));
  NOR2_X1   g0740(.A1(new_n921), .A2(new_n938), .ZN(new_n941));
  OAI21_X1  g0741(.A(new_n865), .B1(new_n940), .B2(new_n941), .ZN(G367));
  INV_X1    g0742(.A(new_n807), .ZN(new_n943));
  OAI221_X1 g0743(.A(new_n803), .B1(new_n212), .B2(new_n566), .C1(new_n943), .C2(new_n238), .ZN(new_n944));
  AND2_X1   g0744(.A1(new_n750), .A2(new_n944), .ZN(new_n945));
  NAND3_X1  g0745(.A1(new_n563), .A2(new_n568), .A3(new_n592), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n946), .A2(new_n681), .ZN(new_n947));
  NAND3_X1  g0747(.A1(new_n584), .A2(new_n947), .A3(new_n593), .ZN(new_n948));
  OAI21_X1  g0748(.A(new_n948), .B1(new_n584), .B2(new_n947), .ZN(new_n949));
  OAI22_X1  g0749(.A1(new_n787), .A2(new_n201), .B1(new_n778), .B2(new_n822), .ZN(new_n950));
  AOI211_X1 g0750(.A(new_n271), .B(new_n950), .C1(G143), .C2(new_n794), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n775), .A2(G68), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n770), .A2(G137), .ZN(new_n953));
  OAI22_X1  g0753(.A1(new_n760), .A2(new_n346), .B1(new_n779), .B2(new_n229), .ZN(new_n954));
  AOI21_X1  g0754(.A(new_n954), .B1(G159), .B2(new_n783), .ZN(new_n955));
  NAND4_X1  g0755(.A1(new_n951), .A2(new_n952), .A3(new_n953), .A4(new_n955), .ZN(new_n956));
  AND3_X1   g0756(.A1(new_n765), .A2(KEYINPUT46), .A3(G116), .ZN(new_n957));
  NOR2_X1   g0757(.A1(new_n760), .A2(new_n477), .ZN(new_n958));
  AOI21_X1  g0758(.A(KEYINPUT46), .B1(new_n765), .B2(G116), .ZN(new_n959));
  NOR4_X1   g0759(.A1(new_n957), .A2(new_n958), .A3(new_n959), .A4(new_n344), .ZN(new_n960));
  INV_X1    g0760(.A(G294), .ZN(new_n961));
  OAI22_X1  g0761(.A1(new_n756), .A2(new_n961), .B1(new_n779), .B2(new_n835), .ZN(new_n962));
  OAI22_X1  g0762(.A1(new_n762), .A2(new_n790), .B1(new_n778), .B2(new_n456), .ZN(new_n963));
  AOI211_X1 g0763(.A(new_n962), .B(new_n963), .C1(G317), .C2(new_n770), .ZN(new_n964));
  OAI211_X1 g0764(.A(new_n960), .B(new_n964), .C1(new_n420), .C2(new_n774), .ZN(new_n965));
  NAND2_X1  g0765(.A1(new_n956), .A2(new_n965), .ZN(new_n966));
  XOR2_X1   g0766(.A(new_n966), .B(KEYINPUT47), .Z(new_n967));
  OAI221_X1 g0767(.A(new_n945), .B1(new_n812), .B2(new_n949), .C1(new_n967), .C2(new_n753), .ZN(new_n968));
  OAI211_X1 g0768(.A(new_n536), .B(new_n544), .C1(new_n535), .C2(new_n682), .ZN(new_n969));
  NAND2_X1  g0769(.A1(new_n663), .A2(new_n681), .ZN(new_n970));
  NAND2_X1  g0770(.A1(new_n969), .A2(new_n970), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n688), .A2(new_n971), .ZN(new_n972));
  XOR2_X1   g0772(.A(new_n972), .B(KEYINPUT111), .Z(new_n973));
  NAND3_X1  g0773(.A1(new_n689), .A2(new_n690), .A3(new_n971), .ZN(new_n974));
  OAI21_X1  g0774(.A(new_n544), .B1(new_n969), .B2(new_n632), .ZN(new_n975));
  AOI22_X1  g0775(.A1(new_n974), .A2(KEYINPUT42), .B1(new_n682), .B2(new_n975), .ZN(new_n976));
  OAI21_X1  g0776(.A(new_n976), .B1(KEYINPUT42), .B2(new_n974), .ZN(new_n977));
  NAND2_X1  g0777(.A1(new_n949), .A2(KEYINPUT43), .ZN(new_n978));
  NAND2_X1  g0778(.A1(new_n977), .A2(new_n978), .ZN(new_n979));
  INV_X1    g0779(.A(new_n979), .ZN(new_n980));
  NAND2_X1  g0780(.A1(new_n973), .A2(new_n980), .ZN(new_n981));
  INV_X1    g0781(.A(new_n981), .ZN(new_n982));
  NOR2_X1   g0782(.A1(new_n973), .A2(new_n980), .ZN(new_n983));
  OAI22_X1  g0783(.A1(new_n982), .A2(new_n983), .B1(KEYINPUT43), .B2(new_n949), .ZN(new_n984));
  INV_X1    g0784(.A(new_n983), .ZN(new_n985));
  NOR2_X1   g0785(.A1(new_n949), .A2(KEYINPUT43), .ZN(new_n986));
  NAND3_X1  g0786(.A1(new_n985), .A2(new_n981), .A3(new_n986), .ZN(new_n987));
  NAND2_X1  g0787(.A1(new_n984), .A2(new_n987), .ZN(new_n988));
  INV_X1    g0788(.A(new_n971), .ZN(new_n989));
  NAND2_X1  g0789(.A1(new_n693), .A2(new_n989), .ZN(new_n990));
  XOR2_X1   g0790(.A(new_n990), .B(KEYINPUT44), .Z(new_n991));
  NOR2_X1   g0791(.A1(new_n693), .A2(new_n989), .ZN(new_n992));
  XNOR2_X1  g0792(.A(new_n992), .B(KEYINPUT45), .ZN(new_n993));
  NAND2_X1  g0793(.A1(new_n991), .A2(new_n993), .ZN(new_n994));
  XNOR2_X1  g0794(.A(new_n994), .B(new_n688), .ZN(new_n995));
  OAI21_X1  g0795(.A(new_n691), .B1(new_n687), .B2(new_n689), .ZN(new_n996));
  XNOR2_X1  g0796(.A(new_n685), .B(new_n996), .ZN(new_n997));
  NAND2_X1  g0797(.A1(new_n741), .A2(new_n997), .ZN(new_n998));
  OAI21_X1  g0798(.A(new_n741), .B1(new_n995), .B2(new_n998), .ZN(new_n999));
  XOR2_X1   g0799(.A(new_n696), .B(KEYINPUT41), .Z(new_n1000));
  INV_X1    g0800(.A(new_n1000), .ZN(new_n1001));
  AOI21_X1  g0801(.A(new_n746), .B1(new_n999), .B2(new_n1001), .ZN(new_n1002));
  OAI21_X1  g0802(.A(new_n968), .B1(new_n988), .B2(new_n1002), .ZN(G387));
  INV_X1    g0803(.A(new_n998), .ZN(new_n1004));
  OAI21_X1  g0804(.A(KEYINPUT115), .B1(new_n1004), .B2(new_n697), .ZN(new_n1005));
  INV_X1    g0805(.A(KEYINPUT115), .ZN(new_n1006));
  NAND3_X1  g0806(.A1(new_n998), .A2(new_n1006), .A3(new_n696), .ZN(new_n1007));
  OAI211_X1 g0807(.A(new_n1005), .B(new_n1007), .C1(new_n741), .C2(new_n997), .ZN(new_n1008));
  NOR2_X1   g0808(.A1(new_n787), .A2(new_n346), .ZN(new_n1009));
  NOR2_X1   g0809(.A1(new_n779), .A2(new_n202), .ZN(new_n1010));
  NOR4_X1   g0810(.A1(new_n1009), .A2(new_n958), .A3(new_n271), .A4(new_n1010), .ZN(new_n1011));
  NAND2_X1  g0811(.A1(new_n775), .A2(new_n564), .ZN(new_n1012));
  AOI22_X1  g0812(.A1(new_n794), .A2(G159), .B1(new_n783), .B2(new_n249), .ZN(new_n1013));
  OAI21_X1  g0813(.A(new_n1013), .B1(new_n229), .B2(new_n778), .ZN(new_n1014));
  INV_X1    g0814(.A(new_n1014), .ZN(new_n1015));
  NAND2_X1  g0815(.A1(new_n770), .A2(G150), .ZN(new_n1016));
  NAND4_X1  g0816(.A1(new_n1011), .A2(new_n1012), .A3(new_n1015), .A4(new_n1016), .ZN(new_n1017));
  AOI22_X1  g0817(.A1(G322), .A2(new_n794), .B1(new_n783), .B2(G311), .ZN(new_n1018));
  INV_X1    g0818(.A(G317), .ZN(new_n1019));
  OAI221_X1 g0819(.A(new_n1018), .B1(new_n456), .B2(new_n779), .C1(new_n1019), .C2(new_n778), .ZN(new_n1020));
  XNOR2_X1  g0820(.A(new_n1020), .B(KEYINPUT48), .ZN(new_n1021));
  OAI221_X1 g0821(.A(new_n1021), .B1(new_n835), .B2(new_n774), .C1(new_n961), .C2(new_n787), .ZN(new_n1022));
  XOR2_X1   g0822(.A(new_n1022), .B(KEYINPUT49), .Z(new_n1023));
  NAND2_X1  g0823(.A1(new_n770), .A2(G326), .ZN(new_n1024));
  OAI211_X1 g0824(.A(new_n1024), .B(new_n271), .C1(new_n466), .C2(new_n760), .ZN(new_n1025));
  OAI21_X1  g0825(.A(new_n1017), .B1(new_n1023), .B2(new_n1025), .ZN(new_n1026));
  AOI21_X1  g0826(.A(new_n753), .B1(new_n1026), .B2(KEYINPUT114), .ZN(new_n1027));
  OAI21_X1  g0827(.A(new_n1027), .B1(KEYINPUT114), .B2(new_n1026), .ZN(new_n1028));
  INV_X1    g0828(.A(new_n698), .ZN(new_n1029));
  AOI22_X1  g0829(.A1(new_n804), .A2(new_n1029), .B1(new_n420), .B2(new_n695), .ZN(new_n1030));
  NOR2_X1   g0830(.A1(new_n235), .A2(new_n450), .ZN(new_n1031));
  XNOR2_X1  g0831(.A(KEYINPUT112), .B(KEYINPUT50), .ZN(new_n1032));
  OAI21_X1  g0832(.A(new_n1032), .B1(new_n248), .B2(G50), .ZN(new_n1033));
  AOI21_X1  g0833(.A(G45), .B1(G68), .B2(G77), .ZN(new_n1034));
  NAND3_X1  g0834(.A1(new_n1033), .A2(new_n698), .A3(new_n1034), .ZN(new_n1035));
  NOR3_X1   g0835(.A1(new_n248), .A2(new_n1032), .A3(G50), .ZN(new_n1036));
  OAI21_X1  g0836(.A(new_n807), .B1(new_n1035), .B2(new_n1036), .ZN(new_n1037));
  OAI21_X1  g0837(.A(new_n1030), .B1(new_n1031), .B2(new_n1037), .ZN(new_n1038));
  AOI21_X1  g0838(.A(new_n751), .B1(new_n1038), .B2(new_n803), .ZN(new_n1039));
  XOR2_X1   g0839(.A(new_n1039), .B(KEYINPUT113), .Z(new_n1040));
  OAI211_X1 g0840(.A(new_n1028), .B(new_n1040), .C1(new_n687), .C2(new_n812), .ZN(new_n1041));
  INV_X1    g0841(.A(new_n997), .ZN(new_n1042));
  OAI21_X1  g0842(.A(new_n1041), .B1(new_n1042), .B2(new_n745), .ZN(new_n1043));
  INV_X1    g0843(.A(new_n1043), .ZN(new_n1044));
  NAND2_X1  g0844(.A1(new_n1008), .A2(new_n1044), .ZN(G393));
  XOR2_X1   g0845(.A(new_n994), .B(new_n688), .Z(new_n1046));
  NAND2_X1  g0846(.A1(new_n1046), .A2(new_n1004), .ZN(new_n1047));
  NAND2_X1  g0847(.A1(new_n995), .A2(new_n998), .ZN(new_n1048));
  NAND3_X1  g0848(.A1(new_n1047), .A2(new_n1048), .A3(new_n696), .ZN(new_n1049));
  NAND2_X1  g0849(.A1(new_n1046), .A2(new_n746), .ZN(new_n1050));
  NAND2_X1  g0850(.A1(new_n807), .A2(new_n246), .ZN(new_n1051));
  OAI211_X1 g0851(.A(new_n1051), .B(new_n803), .C1(new_n477), .C2(new_n212), .ZN(new_n1052));
  INV_X1    g0852(.A(KEYINPUT116), .ZN(new_n1053));
  OR2_X1    g0853(.A1(new_n1052), .A2(new_n1053), .ZN(new_n1054));
  NAND2_X1  g0854(.A1(new_n1052), .A2(new_n1053), .ZN(new_n1055));
  NAND3_X1  g0855(.A1(new_n1054), .A2(new_n750), .A3(new_n1055), .ZN(new_n1056));
  OAI22_X1  g0856(.A1(new_n762), .A2(new_n1019), .B1(new_n778), .B2(new_n790), .ZN(new_n1057));
  XOR2_X1   g0857(.A(new_n1057), .B(KEYINPUT52), .Z(new_n1058));
  OAI21_X1  g0858(.A(new_n271), .B1(new_n760), .B2(new_n420), .ZN(new_n1059));
  OAI22_X1  g0859(.A1(new_n787), .A2(new_n835), .B1(new_n756), .B2(new_n456), .ZN(new_n1060));
  AOI211_X1 g0860(.A(new_n1059), .B(new_n1060), .C1(G294), .C2(new_n819), .ZN(new_n1061));
  NAND2_X1  g0861(.A1(new_n775), .A2(G116), .ZN(new_n1062));
  NAND2_X1  g0862(.A1(new_n1061), .A2(new_n1062), .ZN(new_n1063));
  AOI211_X1 g0863(.A(new_n1058), .B(new_n1063), .C1(G322), .C2(new_n770), .ZN(new_n1064));
  OR2_X1    g0864(.A1(new_n1064), .A2(KEYINPUT117), .ZN(new_n1065));
  NAND2_X1  g0865(.A1(new_n1064), .A2(KEYINPUT117), .ZN(new_n1066));
  OAI21_X1  g0866(.A(new_n344), .B1(new_n760), .B2(new_n218), .ZN(new_n1067));
  OAI22_X1  g0867(.A1(new_n787), .A2(new_n202), .B1(new_n756), .B2(new_n229), .ZN(new_n1068));
  AOI211_X1 g0868(.A(new_n1067), .B(new_n1068), .C1(new_n249), .C2(new_n819), .ZN(new_n1069));
  NAND2_X1  g0869(.A1(new_n770), .A2(G143), .ZN(new_n1070));
  INV_X1    g0870(.A(G159), .ZN(new_n1071));
  OAI22_X1  g0871(.A1(new_n762), .A2(new_n822), .B1(new_n778), .B2(new_n1071), .ZN(new_n1072));
  XNOR2_X1  g0872(.A(new_n1072), .B(KEYINPUT51), .ZN(new_n1073));
  NAND2_X1  g0873(.A1(new_n775), .A2(G77), .ZN(new_n1074));
  NAND4_X1  g0874(.A1(new_n1069), .A2(new_n1070), .A3(new_n1073), .A4(new_n1074), .ZN(new_n1075));
  NAND3_X1  g0875(.A1(new_n1065), .A2(new_n1066), .A3(new_n1075), .ZN(new_n1076));
  AOI21_X1  g0876(.A(new_n1056), .B1(new_n1076), .B2(new_n752), .ZN(new_n1077));
  INV_X1    g0877(.A(new_n802), .ZN(new_n1078));
  OAI21_X1  g0878(.A(new_n1077), .B1(new_n1078), .B2(new_n971), .ZN(new_n1079));
  NAND3_X1  g0879(.A1(new_n1049), .A2(new_n1050), .A3(new_n1079), .ZN(G390));
  NAND2_X1  g0880(.A1(new_n841), .A2(new_n442), .ZN(new_n1081));
  AOI21_X1  g0881(.A(new_n840), .B1(new_n732), .B2(new_n1081), .ZN(new_n1082));
  INV_X1    g0882(.A(new_n1082), .ZN(new_n1083));
  INV_X1    g0883(.A(new_n915), .ZN(new_n1084));
  AOI21_X1  g0884(.A(new_n1084), .B1(new_n731), .B2(new_n842), .ZN(new_n1085));
  NAND2_X1  g0885(.A1(new_n727), .A2(G330), .ZN(new_n1086));
  NOR2_X1   g0886(.A1(new_n1086), .A2(new_n923), .ZN(new_n1087));
  OAI21_X1  g0887(.A(new_n1083), .B1(new_n1085), .B2(new_n1087), .ZN(new_n1088));
  NAND2_X1  g0888(.A1(new_n731), .A2(new_n931), .ZN(new_n1089));
  OAI21_X1  g0889(.A(new_n915), .B1(new_n1086), .B2(new_n843), .ZN(new_n1090));
  NOR3_X1   g0890(.A1(new_n737), .A2(new_n739), .A3(new_n840), .ZN(new_n1091));
  INV_X1    g0891(.A(KEYINPUT118), .ZN(new_n1092));
  INV_X1    g0892(.A(new_n1081), .ZN(new_n1093));
  NOR3_X1   g0893(.A1(new_n1091), .A2(new_n1092), .A3(new_n1093), .ZN(new_n1094));
  NAND2_X1  g0894(.A1(new_n736), .A2(new_n682), .ZN(new_n1095));
  NAND2_X1  g0895(.A1(new_n1095), .A2(new_n738), .ZN(new_n1096));
  NAND3_X1  g0896(.A1(new_n736), .A2(KEYINPUT98), .A3(new_n682), .ZN(new_n1097));
  NAND3_X1  g0897(.A1(new_n1096), .A2(new_n1097), .A3(new_n916), .ZN(new_n1098));
  AOI21_X1  g0898(.A(KEYINPUT118), .B1(new_n1098), .B2(new_n1081), .ZN(new_n1099));
  OAI211_X1 g0899(.A(new_n1089), .B(new_n1090), .C1(new_n1094), .C2(new_n1099), .ZN(new_n1100));
  NAND2_X1  g0900(.A1(new_n1088), .A2(new_n1100), .ZN(new_n1101));
  NAND3_X1  g0901(.A1(new_n445), .A2(G330), .A3(new_n727), .ZN(new_n1102));
  NAND3_X1  g0902(.A1(new_n919), .A2(new_n674), .A3(new_n1102), .ZN(new_n1103));
  INV_X1    g0903(.A(new_n1103), .ZN(new_n1104));
  NAND2_X1  g0904(.A1(new_n1101), .A2(new_n1104), .ZN(new_n1105));
  OAI21_X1  g0905(.A(new_n1092), .B1(new_n1091), .B2(new_n1093), .ZN(new_n1106));
  NAND3_X1  g0906(.A1(new_n1098), .A2(KEYINPUT118), .A3(new_n1081), .ZN(new_n1107));
  NAND3_X1  g0907(.A1(new_n1106), .A2(new_n1084), .A3(new_n1107), .ZN(new_n1108));
  AND3_X1   g0908(.A1(new_n925), .A2(new_n904), .A3(new_n929), .ZN(new_n1109));
  NAND2_X1  g0909(.A1(new_n1108), .A2(new_n1109), .ZN(new_n1110));
  OAI21_X1  g0910(.A(new_n902), .B1(new_n917), .B2(new_n903), .ZN(new_n1111));
  AND3_X1   g0911(.A1(new_n1110), .A2(new_n1111), .A3(new_n1089), .ZN(new_n1112));
  INV_X1    g0912(.A(new_n1087), .ZN(new_n1113));
  AOI21_X1  g0913(.A(new_n1113), .B1(new_n1110), .B2(new_n1111), .ZN(new_n1114));
  OAI21_X1  g0914(.A(new_n1105), .B1(new_n1112), .B2(new_n1114), .ZN(new_n1115));
  AOI21_X1  g0915(.A(new_n1103), .B1(new_n1088), .B2(new_n1100), .ZN(new_n1116));
  NAND3_X1  g0916(.A1(new_n1110), .A2(new_n1111), .A3(new_n1089), .ZN(new_n1117));
  OAI21_X1  g0917(.A(new_n904), .B1(new_n1082), .B2(new_n915), .ZN(new_n1118));
  AOI22_X1  g0918(.A1(new_n1108), .A2(new_n1109), .B1(new_n1118), .B2(new_n902), .ZN(new_n1119));
  OAI211_X1 g0919(.A(new_n1116), .B(new_n1117), .C1(new_n1119), .C2(new_n1113), .ZN(new_n1120));
  NAND3_X1  g0920(.A1(new_n1115), .A2(new_n1120), .A3(new_n696), .ZN(new_n1121));
  OAI211_X1 g0921(.A(new_n1117), .B(new_n746), .C1(new_n1119), .C2(new_n1113), .ZN(new_n1122));
  NAND2_X1  g0922(.A1(new_n902), .A2(new_n800), .ZN(new_n1123));
  AOI21_X1  g0923(.A(new_n751), .B1(new_n248), .B2(new_n816), .ZN(new_n1124));
  OAI22_X1  g0924(.A1(new_n760), .A2(new_n202), .B1(new_n779), .B2(new_n477), .ZN(new_n1125));
  AOI211_X1 g0925(.A(new_n344), .B(new_n1125), .C1(G87), .C2(new_n765), .ZN(new_n1126));
  NAND2_X1  g0926(.A1(new_n770), .A2(G294), .ZN(new_n1127));
  OAI22_X1  g0927(.A1(new_n762), .A2(new_n835), .B1(new_n778), .B2(new_n466), .ZN(new_n1128));
  AOI21_X1  g0928(.A(new_n1128), .B1(G107), .B2(new_n783), .ZN(new_n1129));
  NAND4_X1  g0929(.A1(new_n1126), .A2(new_n1074), .A3(new_n1127), .A4(new_n1129), .ZN(new_n1130));
  XNOR2_X1  g0930(.A(KEYINPUT54), .B(G143), .ZN(new_n1131));
  NOR2_X1   g0931(.A1(new_n779), .A2(new_n1131), .ZN(new_n1132));
  INV_X1    g0932(.A(G132), .ZN(new_n1133));
  OAI22_X1  g0933(.A1(new_n760), .A2(new_n229), .B1(new_n1133), .B2(new_n778), .ZN(new_n1134));
  AOI211_X1 g0934(.A(new_n1132), .B(new_n1134), .C1(G128), .C2(new_n794), .ZN(new_n1135));
  NAND2_X1  g0935(.A1(new_n775), .A2(G159), .ZN(new_n1136));
  AOI21_X1  g0936(.A(new_n271), .B1(new_n783), .B2(G137), .ZN(new_n1137));
  INV_X1    g0937(.A(KEYINPUT53), .ZN(new_n1138));
  OAI21_X1  g0938(.A(new_n1138), .B1(new_n787), .B2(new_n822), .ZN(new_n1139));
  NAND3_X1  g0939(.A1(new_n765), .A2(KEYINPUT53), .A3(G150), .ZN(new_n1140));
  AOI22_X1  g0940(.A1(new_n1139), .A2(new_n1140), .B1(G125), .B2(new_n770), .ZN(new_n1141));
  NAND4_X1  g0941(.A1(new_n1135), .A2(new_n1136), .A3(new_n1137), .A4(new_n1141), .ZN(new_n1142));
  AND2_X1   g0942(.A1(new_n1130), .A2(new_n1142), .ZN(new_n1143));
  OAI211_X1 g0943(.A(new_n1123), .B(new_n1124), .C1(new_n753), .C2(new_n1143), .ZN(new_n1144));
  AND2_X1   g0944(.A1(new_n1122), .A2(new_n1144), .ZN(new_n1145));
  NAND2_X1  g0945(.A1(new_n1121), .A2(new_n1145), .ZN(G378));
  OAI21_X1  g0946(.A(new_n747), .B1(G50), .B2(new_n817), .ZN(new_n1147));
  XOR2_X1   g0947(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1148));
  INV_X1    g0948(.A(new_n1148), .ZN(new_n1149));
  NAND2_X1  g0949(.A1(new_n365), .A2(new_n877), .ZN(new_n1150));
  XOR2_X1   g0950(.A(new_n1150), .B(KEYINPUT120), .Z(new_n1151));
  INV_X1    g0951(.A(new_n1151), .ZN(new_n1152));
  NAND2_X1  g0952(.A1(new_n383), .A2(new_n1152), .ZN(new_n1153));
  INV_X1    g0953(.A(new_n1153), .ZN(new_n1154));
  NOR2_X1   g0954(.A1(new_n383), .A2(new_n1152), .ZN(new_n1155));
  OAI21_X1  g0955(.A(new_n1149), .B1(new_n1154), .B2(new_n1155), .ZN(new_n1156));
  INV_X1    g0956(.A(new_n1155), .ZN(new_n1157));
  NAND3_X1  g0957(.A1(new_n1157), .A2(new_n1148), .A3(new_n1153), .ZN(new_n1158));
  NAND2_X1  g0958(.A1(new_n1156), .A2(new_n1158), .ZN(new_n1159));
  NOR2_X1   g0959(.A1(new_n1159), .A2(new_n801), .ZN(new_n1160));
  INV_X1    g0960(.A(G41), .ZN(new_n1161));
  AOI21_X1  g0961(.A(G50), .B1(new_n264), .B2(new_n1161), .ZN(new_n1162));
  AOI22_X1  g0962(.A1(G116), .A2(new_n794), .B1(new_n792), .B2(G107), .ZN(new_n1163));
  OAI221_X1 g0963(.A(new_n1163), .B1(new_n477), .B2(new_n756), .C1(new_n201), .C2(new_n760), .ZN(new_n1164));
  NOR4_X1   g0964(.A1(new_n1164), .A2(G41), .A3(new_n344), .A4(new_n1009), .ZN(new_n1165));
  AOI22_X1  g0965(.A1(new_n564), .A2(new_n819), .B1(G283), .B2(new_n770), .ZN(new_n1166));
  NAND3_X1  g0966(.A1(new_n1165), .A2(new_n952), .A3(new_n1166), .ZN(new_n1167));
  INV_X1    g0967(.A(KEYINPUT58), .ZN(new_n1168));
  AOI21_X1  g0968(.A(new_n1162), .B1(new_n1167), .B2(new_n1168), .ZN(new_n1169));
  OAI22_X1  g0969(.A1(new_n756), .A2(new_n1133), .B1(new_n779), .B2(new_n821), .ZN(new_n1170));
  XNOR2_X1  g0970(.A(new_n1170), .B(KEYINPUT119), .ZN(new_n1171));
  NAND2_X1  g0971(.A1(new_n792), .A2(G128), .ZN(new_n1172));
  NAND2_X1  g0972(.A1(new_n794), .A2(G125), .ZN(new_n1173));
  OAI211_X1 g0973(.A(new_n1172), .B(new_n1173), .C1(new_n787), .C2(new_n1131), .ZN(new_n1174));
  AOI211_X1 g0974(.A(new_n1171), .B(new_n1174), .C1(G150), .C2(new_n775), .ZN(new_n1175));
  INV_X1    g0975(.A(new_n1175), .ZN(new_n1176));
  NOR2_X1   g0976(.A1(new_n1176), .A2(KEYINPUT59), .ZN(new_n1177));
  OAI211_X1 g0977(.A(new_n262), .B(new_n1161), .C1(new_n760), .C2(new_n1071), .ZN(new_n1178));
  AOI21_X1  g0978(.A(new_n1178), .B1(new_n770), .B2(G124), .ZN(new_n1179));
  INV_X1    g0979(.A(KEYINPUT59), .ZN(new_n1180));
  OAI21_X1  g0980(.A(new_n1179), .B1(new_n1175), .B2(new_n1180), .ZN(new_n1181));
  OAI221_X1 g0981(.A(new_n1169), .B1(new_n1168), .B2(new_n1167), .C1(new_n1177), .C2(new_n1181), .ZN(new_n1182));
  AOI211_X1 g0982(.A(new_n1147), .B(new_n1160), .C1(new_n752), .C2(new_n1182), .ZN(new_n1183));
  NAND3_X1  g0983(.A1(new_n930), .A2(G330), .A3(new_n933), .ZN(new_n1184));
  INV_X1    g0984(.A(KEYINPUT121), .ZN(new_n1185));
  NAND2_X1  g0985(.A1(new_n1184), .A2(new_n1185), .ZN(new_n1186));
  NAND4_X1  g0986(.A1(new_n930), .A2(new_n933), .A3(KEYINPUT121), .A4(G330), .ZN(new_n1187));
  NAND3_X1  g0987(.A1(new_n1186), .A2(new_n1187), .A3(new_n1159), .ZN(new_n1188));
  AND2_X1   g0988(.A1(new_n1156), .A2(new_n1158), .ZN(new_n1189));
  NAND4_X1  g0989(.A1(new_n934), .A2(new_n1189), .A3(KEYINPUT121), .A4(G330), .ZN(new_n1190));
  AND3_X1   g0990(.A1(new_n1188), .A2(new_n918), .A3(new_n1190), .ZN(new_n1191));
  AOI21_X1  g0991(.A(new_n918), .B1(new_n1188), .B2(new_n1190), .ZN(new_n1192));
  NOR2_X1   g0992(.A1(new_n1191), .A2(new_n1192), .ZN(new_n1193));
  AOI21_X1  g0993(.A(new_n1183), .B1(new_n1193), .B2(new_n746), .ZN(new_n1194));
  OAI21_X1  g0994(.A(new_n1117), .B1(new_n1119), .B2(new_n1113), .ZN(new_n1195));
  OAI21_X1  g0995(.A(new_n1104), .B1(new_n1195), .B2(new_n1105), .ZN(new_n1196));
  NAND3_X1  g0996(.A1(new_n1196), .A2(KEYINPUT57), .A3(new_n1193), .ZN(new_n1197));
  NAND2_X1  g0997(.A1(new_n1197), .A2(new_n696), .ZN(new_n1198));
  AOI21_X1  g0998(.A(KEYINPUT57), .B1(new_n1196), .B2(new_n1193), .ZN(new_n1199));
  OAI21_X1  g0999(.A(new_n1194), .B1(new_n1198), .B2(new_n1199), .ZN(G375));
  OAI22_X1  g1000(.A1(new_n756), .A2(new_n466), .B1(new_n779), .B2(new_n420), .ZN(new_n1201));
  XNOR2_X1  g1001(.A(new_n1201), .B(KEYINPUT122), .ZN(new_n1202));
  OAI21_X1  g1002(.A(new_n271), .B1(new_n760), .B2(new_n346), .ZN(new_n1203));
  OAI22_X1  g1003(.A1(new_n787), .A2(new_n477), .B1(new_n778), .B2(new_n835), .ZN(new_n1204));
  AOI211_X1 g1004(.A(new_n1203), .B(new_n1204), .C1(G294), .C2(new_n794), .ZN(new_n1205));
  NAND2_X1  g1005(.A1(new_n1205), .A2(new_n1012), .ZN(new_n1206));
  AOI211_X1 g1006(.A(new_n1202), .B(new_n1206), .C1(G303), .C2(new_n770), .ZN(new_n1207));
  OR2_X1    g1007(.A1(new_n1207), .A2(KEYINPUT123), .ZN(new_n1208));
  NOR2_X1   g1008(.A1(new_n756), .A2(new_n1131), .ZN(new_n1209));
  OAI22_X1  g1009(.A1(new_n778), .A2(new_n821), .B1(new_n779), .B2(new_n822), .ZN(new_n1210));
  AOI211_X1 g1010(.A(new_n1209), .B(new_n1210), .C1(G159), .C2(new_n765), .ZN(new_n1211));
  NAND2_X1  g1011(.A1(new_n775), .A2(G50), .ZN(new_n1212));
  AOI21_X1  g1012(.A(new_n271), .B1(new_n759), .B2(G58), .ZN(new_n1213));
  OR3_X1    g1013(.A1(new_n762), .A2(KEYINPUT124), .A3(new_n1133), .ZN(new_n1214));
  OAI21_X1  g1014(.A(KEYINPUT124), .B1(new_n762), .B2(new_n1133), .ZN(new_n1215));
  AOI22_X1  g1015(.A1(new_n1214), .A2(new_n1215), .B1(new_n770), .B2(G128), .ZN(new_n1216));
  NAND4_X1  g1016(.A1(new_n1211), .A2(new_n1212), .A3(new_n1213), .A4(new_n1216), .ZN(new_n1217));
  NAND2_X1  g1017(.A1(new_n1208), .A2(new_n1217), .ZN(new_n1218));
  AOI21_X1  g1018(.A(new_n1218), .B1(KEYINPUT123), .B2(new_n1207), .ZN(new_n1219));
  OAI221_X1 g1019(.A(new_n750), .B1(G68), .B2(new_n817), .C1(new_n1219), .C2(new_n753), .ZN(new_n1220));
  AOI21_X1  g1020(.A(new_n1220), .B1(new_n800), .B2(new_n915), .ZN(new_n1221));
  AOI21_X1  g1021(.A(new_n1221), .B1(new_n1101), .B2(new_n746), .ZN(new_n1222));
  NAND2_X1  g1022(.A1(new_n1105), .A2(new_n1001), .ZN(new_n1223));
  NOR2_X1   g1023(.A1(new_n1101), .A2(new_n1104), .ZN(new_n1224));
  OAI21_X1  g1024(.A(new_n1222), .B1(new_n1223), .B2(new_n1224), .ZN(G381));
  INV_X1    g1025(.A(G390), .ZN(new_n1226));
  INV_X1    g1026(.A(G384), .ZN(new_n1227));
  NAND2_X1  g1027(.A1(new_n1226), .A2(new_n1227), .ZN(new_n1228));
  NOR2_X1   g1028(.A1(G393), .A2(G396), .ZN(new_n1229));
  INV_X1    g1029(.A(new_n1229), .ZN(new_n1230));
  NOR4_X1   g1030(.A1(new_n1228), .A2(G387), .A3(new_n1230), .A4(G381), .ZN(new_n1231));
  OR2_X1    g1031(.A1(new_n1198), .A2(new_n1199), .ZN(new_n1232));
  NAND2_X1  g1032(.A1(G378), .A2(KEYINPUT125), .ZN(new_n1233));
  INV_X1    g1033(.A(KEYINPUT125), .ZN(new_n1234));
  NAND3_X1  g1034(.A1(new_n1121), .A2(new_n1145), .A3(new_n1234), .ZN(new_n1235));
  AND2_X1   g1035(.A1(new_n1233), .A2(new_n1235), .ZN(new_n1236));
  NAND4_X1  g1036(.A1(new_n1231), .A2(new_n1194), .A3(new_n1232), .A4(new_n1236), .ZN(G407));
  NAND2_X1  g1037(.A1(new_n680), .A2(G213), .ZN(new_n1238));
  INV_X1    g1038(.A(new_n1238), .ZN(new_n1239));
  NAND4_X1  g1039(.A1(new_n1236), .A2(new_n1232), .A3(new_n1194), .A4(new_n1239), .ZN(new_n1240));
  NAND3_X1  g1040(.A1(G407), .A2(new_n1240), .A3(G213), .ZN(G409));
  NAND2_X1  g1041(.A1(G393), .A2(G396), .ZN(new_n1242));
  AOI21_X1  g1042(.A(G390), .B1(new_n1230), .B2(new_n1242), .ZN(new_n1243));
  INV_X1    g1043(.A(new_n1243), .ZN(new_n1244));
  NAND2_X1  g1044(.A1(G387), .A2(KEYINPUT126), .ZN(new_n1245));
  INV_X1    g1045(.A(KEYINPUT126), .ZN(new_n1246));
  OAI211_X1 g1046(.A(new_n1246), .B(new_n968), .C1(new_n988), .C2(new_n1002), .ZN(new_n1247));
  NAND3_X1  g1047(.A1(new_n1230), .A2(G390), .A3(new_n1242), .ZN(new_n1248));
  NAND4_X1  g1048(.A1(new_n1244), .A2(new_n1245), .A3(new_n1247), .A4(new_n1248), .ZN(new_n1249));
  NAND2_X1  g1049(.A1(new_n1245), .A2(new_n1247), .ZN(new_n1250));
  INV_X1    g1050(.A(new_n1248), .ZN(new_n1251));
  OAI21_X1  g1051(.A(new_n1250), .B1(new_n1251), .B2(new_n1243), .ZN(new_n1252));
  NAND2_X1  g1052(.A1(new_n1249), .A2(new_n1252), .ZN(new_n1253));
  OAI211_X1 g1053(.A(G378), .B(new_n1194), .C1(new_n1198), .C2(new_n1199), .ZN(new_n1254));
  NAND3_X1  g1054(.A1(new_n1196), .A2(new_n1001), .A3(new_n1193), .ZN(new_n1255));
  NAND2_X1  g1055(.A1(new_n1255), .A2(new_n1194), .ZN(new_n1256));
  NAND3_X1  g1056(.A1(new_n1233), .A2(new_n1256), .A3(new_n1235), .ZN(new_n1257));
  NAND2_X1  g1057(.A1(new_n1254), .A2(new_n1257), .ZN(new_n1258));
  NAND2_X1  g1058(.A1(new_n1258), .A2(new_n1238), .ZN(new_n1259));
  NAND4_X1  g1059(.A1(new_n1088), .A2(KEYINPUT60), .A3(new_n1100), .A4(new_n1103), .ZN(new_n1260));
  AND2_X1   g1060(.A1(new_n1260), .A2(new_n696), .ZN(new_n1261));
  INV_X1    g1061(.A(KEYINPUT60), .ZN(new_n1262));
  NOR2_X1   g1062(.A1(new_n1116), .A2(new_n1262), .ZN(new_n1263));
  OAI21_X1  g1063(.A(new_n1261), .B1(new_n1263), .B2(new_n1224), .ZN(new_n1264));
  NAND3_X1  g1064(.A1(new_n1264), .A2(G384), .A3(new_n1222), .ZN(new_n1265));
  INV_X1    g1065(.A(new_n1265), .ZN(new_n1266));
  AOI21_X1  g1066(.A(G384), .B1(new_n1264), .B2(new_n1222), .ZN(new_n1267));
  OAI211_X1 g1067(.A(G2897), .B(new_n1239), .C1(new_n1266), .C2(new_n1267), .ZN(new_n1268));
  INV_X1    g1068(.A(new_n1267), .ZN(new_n1269));
  NAND2_X1  g1069(.A1(new_n1239), .A2(G2897), .ZN(new_n1270));
  NAND3_X1  g1070(.A1(new_n1269), .A2(new_n1265), .A3(new_n1270), .ZN(new_n1271));
  NAND2_X1  g1071(.A1(new_n1268), .A2(new_n1271), .ZN(new_n1272));
  INV_X1    g1072(.A(new_n1272), .ZN(new_n1273));
  AOI21_X1  g1073(.A(KEYINPUT61), .B1(new_n1259), .B2(new_n1273), .ZN(new_n1274));
  AOI21_X1  g1074(.A(new_n1239), .B1(new_n1254), .B2(new_n1257), .ZN(new_n1275));
  NOR2_X1   g1075(.A1(new_n1266), .A2(new_n1267), .ZN(new_n1276));
  NAND2_X1  g1076(.A1(new_n1275), .A2(new_n1276), .ZN(new_n1277));
  INV_X1    g1077(.A(KEYINPUT63), .ZN(new_n1278));
  NAND2_X1  g1078(.A1(new_n1277), .A2(new_n1278), .ZN(new_n1279));
  NAND3_X1  g1079(.A1(new_n1275), .A2(KEYINPUT63), .A3(new_n1276), .ZN(new_n1280));
  NAND4_X1  g1080(.A1(new_n1253), .A2(new_n1274), .A3(new_n1279), .A4(new_n1280), .ZN(new_n1281));
  INV_X1    g1081(.A(KEYINPUT62), .ZN(new_n1282));
  AND3_X1   g1082(.A1(new_n1275), .A2(new_n1282), .A3(new_n1276), .ZN(new_n1283));
  INV_X1    g1083(.A(KEYINPUT61), .ZN(new_n1284));
  OAI21_X1  g1084(.A(new_n1284), .B1(new_n1275), .B2(new_n1272), .ZN(new_n1285));
  AOI21_X1  g1085(.A(new_n1282), .B1(new_n1275), .B2(new_n1276), .ZN(new_n1286));
  NOR3_X1   g1086(.A1(new_n1283), .A2(new_n1285), .A3(new_n1286), .ZN(new_n1287));
  OAI21_X1  g1087(.A(new_n1281), .B1(new_n1287), .B2(new_n1253), .ZN(G405));
  NAND2_X1  g1088(.A1(new_n1236), .A2(G375), .ZN(new_n1289));
  NAND2_X1  g1089(.A1(new_n1289), .A2(new_n1254), .ZN(new_n1290));
  INV_X1    g1090(.A(KEYINPUT127), .ZN(new_n1291));
  NAND2_X1  g1091(.A1(new_n1276), .A2(new_n1291), .ZN(new_n1292));
  OAI21_X1  g1092(.A(KEYINPUT127), .B1(new_n1266), .B2(new_n1267), .ZN(new_n1293));
  NAND3_X1  g1093(.A1(new_n1290), .A2(new_n1292), .A3(new_n1293), .ZN(new_n1294));
  NAND4_X1  g1094(.A1(new_n1289), .A2(new_n1291), .A3(new_n1276), .A4(new_n1254), .ZN(new_n1295));
  NAND2_X1  g1095(.A1(new_n1294), .A2(new_n1295), .ZN(new_n1296));
  NAND2_X1  g1096(.A1(new_n1296), .A2(new_n1253), .ZN(new_n1297));
  NAND4_X1  g1097(.A1(new_n1294), .A2(new_n1249), .A3(new_n1252), .A4(new_n1295), .ZN(new_n1298));
  NAND2_X1  g1098(.A1(new_n1297), .A2(new_n1298), .ZN(G402));
endmodule


