//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 1 0 0 0 0 0 0 1 0 1 1 1 0 0 0 0 1 0 1 0 1 0 0 0 0 0 0 1 0 0 1 1 1 1 0 0 0 0 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 0 0 1 0 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:31:18 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n443, new_n447, new_n451, new_n452, new_n453, new_n456, new_n457,
    new_n458, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n520, new_n521, new_n522, new_n523, new_n524, new_n525,
    new_n526, new_n527, new_n528, new_n529, new_n531, new_n532, new_n533,
    new_n534, new_n535, new_n536, new_n537, new_n538, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n548, new_n549, new_n550,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n560, new_n561, new_n562, new_n563, new_n566, new_n567, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n575, new_n576, new_n577,
    new_n578, new_n579, new_n580, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n604, new_n607, new_n608, new_n610, new_n611, new_n612,
    new_n613, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1155, new_n1156, new_n1157, new_n1158, new_n1159, new_n1160,
    new_n1161, new_n1162, new_n1163;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  XNOR2_X1  g004(.A(KEYINPUT64), .B(G1083), .ZN(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(new_n443));
  XNOR2_X1  g018(.A(new_n443), .B(KEYINPUT65), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g025(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n451));
  XNOR2_X1  g026(.A(new_n451), .B(KEYINPUT2), .ZN(new_n452));
  NOR4_X1   g027(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n453));
  NAND2_X1  g028(.A1(new_n452), .A2(new_n453), .ZN(G261));
  INV_X1    g029(.A(G261), .ZN(G325));
  INV_X1    g030(.A(G2106), .ZN(new_n456));
  INV_X1    g031(.A(G567), .ZN(new_n457));
  OAI22_X1  g032(.A1(new_n452), .A2(new_n456), .B1(new_n457), .B2(new_n453), .ZN(new_n458));
  XOR2_X1   g033(.A(new_n458), .B(KEYINPUT66), .Z(G319));
  INV_X1    g034(.A(KEYINPUT67), .ZN(new_n460));
  INV_X1    g035(.A(G2104), .ZN(new_n461));
  NAND3_X1  g036(.A1(new_n460), .A2(new_n461), .A3(KEYINPUT3), .ZN(new_n462));
  INV_X1    g037(.A(KEYINPUT3), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n463), .A2(G2104), .ZN(new_n464));
  AND2_X1   g039(.A1(new_n462), .A2(new_n464), .ZN(new_n465));
  INV_X1    g040(.A(G2105), .ZN(new_n466));
  OAI21_X1  g041(.A(KEYINPUT67), .B1(new_n463), .B2(G2104), .ZN(new_n467));
  NAND4_X1  g042(.A1(new_n465), .A2(G137), .A3(new_n466), .A4(new_n467), .ZN(new_n468));
  INV_X1    g043(.A(KEYINPUT68), .ZN(new_n469));
  AOI21_X1  g044(.A(new_n469), .B1(G2104), .B2(new_n466), .ZN(new_n470));
  NOR3_X1   g045(.A1(new_n461), .A2(KEYINPUT68), .A3(G2105), .ZN(new_n471));
  OAI21_X1  g046(.A(G101), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n468), .A2(new_n472), .ZN(new_n473));
  INV_X1    g048(.A(new_n473), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n461), .A2(KEYINPUT3), .ZN(new_n475));
  NAND3_X1  g050(.A1(new_n475), .A2(new_n464), .A3(G125), .ZN(new_n476));
  NAND2_X1  g051(.A1(G113), .A2(G2104), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n478), .A2(G2105), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n474), .A2(new_n479), .ZN(new_n480));
  INV_X1    g055(.A(new_n480), .ZN(G160));
  NAND4_X1  g056(.A1(new_n467), .A2(new_n462), .A3(G2105), .A4(new_n464), .ZN(new_n482));
  INV_X1    g057(.A(G124), .ZN(new_n483));
  NOR2_X1   g058(.A1(new_n466), .A2(G112), .ZN(new_n484));
  OAI21_X1  g059(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n485));
  OAI22_X1  g060(.A1(new_n482), .A2(new_n483), .B1(new_n484), .B2(new_n485), .ZN(new_n486));
  NAND4_X1  g061(.A1(new_n467), .A2(new_n462), .A3(new_n466), .A4(new_n464), .ZN(new_n487));
  INV_X1    g062(.A(new_n487), .ZN(new_n488));
  AOI21_X1  g063(.A(new_n486), .B1(new_n488), .B2(G136), .ZN(G162));
  NOR2_X1   g064(.A1(new_n466), .A2(G114), .ZN(new_n490));
  OAI21_X1  g065(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n491));
  NOR2_X1   g066(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  INV_X1    g067(.A(new_n482), .ZN(new_n493));
  AOI21_X1  g068(.A(new_n492), .B1(new_n493), .B2(G126), .ZN(new_n494));
  INV_X1    g069(.A(G138), .ZN(new_n495));
  NOR2_X1   g070(.A1(new_n495), .A2(G2105), .ZN(new_n496));
  NAND4_X1  g071(.A1(new_n467), .A2(new_n462), .A3(new_n464), .A4(new_n496), .ZN(new_n497));
  NAND2_X1  g072(.A1(new_n497), .A2(KEYINPUT4), .ZN(new_n498));
  INV_X1    g073(.A(KEYINPUT4), .ZN(new_n499));
  OAI211_X1 g074(.A(G138), .B(new_n466), .C1(new_n499), .C2(KEYINPUT69), .ZN(new_n500));
  INV_X1    g075(.A(KEYINPUT69), .ZN(new_n501));
  NOR2_X1   g076(.A1(new_n501), .A2(KEYINPUT4), .ZN(new_n502));
  NOR2_X1   g077(.A1(new_n500), .A2(new_n502), .ZN(new_n503));
  AND2_X1   g078(.A1(new_n475), .A2(new_n464), .ZN(new_n504));
  NAND2_X1  g079(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  NAND2_X1  g080(.A1(new_n498), .A2(new_n505), .ZN(new_n506));
  NAND2_X1  g081(.A1(new_n494), .A2(new_n506), .ZN(new_n507));
  INV_X1    g082(.A(new_n507), .ZN(G164));
  XNOR2_X1  g083(.A(KEYINPUT5), .B(G543), .ZN(new_n509));
  XNOR2_X1  g084(.A(KEYINPUT6), .B(G651), .ZN(new_n510));
  NAND3_X1  g085(.A1(new_n509), .A2(new_n510), .A3(G88), .ZN(new_n511));
  NAND3_X1  g086(.A1(new_n510), .A2(G50), .A3(G543), .ZN(new_n512));
  INV_X1    g087(.A(KEYINPUT70), .ZN(new_n513));
  AND3_X1   g088(.A1(new_n511), .A2(new_n512), .A3(new_n513), .ZN(new_n514));
  AOI21_X1  g089(.A(new_n513), .B1(new_n511), .B2(new_n512), .ZN(new_n515));
  INV_X1    g090(.A(G651), .ZN(new_n516));
  AOI22_X1  g091(.A1(new_n509), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n517));
  OAI22_X1  g092(.A1(new_n514), .A2(new_n515), .B1(new_n516), .B2(new_n517), .ZN(new_n518));
  INV_X1    g093(.A(new_n518), .ZN(G166));
  XOR2_X1   g094(.A(KEYINPUT71), .B(KEYINPUT7), .Z(new_n520));
  NAND3_X1  g095(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n521));
  XNOR2_X1  g096(.A(new_n520), .B(new_n521), .ZN(new_n522));
  NAND3_X1  g097(.A1(new_n509), .A2(G63), .A3(G651), .ZN(new_n523));
  NAND2_X1  g098(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  NAND2_X1  g099(.A1(new_n510), .A2(new_n509), .ZN(new_n525));
  XNOR2_X1  g100(.A(KEYINPUT72), .B(G89), .ZN(new_n526));
  NAND2_X1  g101(.A1(new_n510), .A2(G543), .ZN(new_n527));
  INV_X1    g102(.A(G51), .ZN(new_n528));
  OAI22_X1  g103(.A1(new_n525), .A2(new_n526), .B1(new_n527), .B2(new_n528), .ZN(new_n529));
  NOR2_X1   g104(.A1(new_n524), .A2(new_n529), .ZN(G168));
  INV_X1    g105(.A(G90), .ZN(new_n531));
  INV_X1    g106(.A(G52), .ZN(new_n532));
  OAI22_X1  g107(.A1(new_n525), .A2(new_n531), .B1(new_n527), .B2(new_n532), .ZN(new_n533));
  INV_X1    g108(.A(KEYINPUT73), .ZN(new_n534));
  XNOR2_X1  g109(.A(new_n533), .B(new_n534), .ZN(new_n535));
  AOI22_X1  g110(.A1(new_n509), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n536));
  OR2_X1    g111(.A1(new_n536), .A2(new_n516), .ZN(new_n537));
  NAND2_X1  g112(.A1(new_n535), .A2(new_n537), .ZN(new_n538));
  INV_X1    g113(.A(new_n538), .ZN(G171));
  INV_X1    g114(.A(G81), .ZN(new_n540));
  XNOR2_X1  g115(.A(KEYINPUT74), .B(G43), .ZN(new_n541));
  OAI22_X1  g116(.A1(new_n525), .A2(new_n540), .B1(new_n527), .B2(new_n541), .ZN(new_n542));
  AOI22_X1  g117(.A1(new_n509), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n543));
  NOR2_X1   g118(.A1(new_n543), .A2(new_n516), .ZN(new_n544));
  NOR2_X1   g119(.A1(new_n542), .A2(new_n544), .ZN(new_n545));
  NAND2_X1  g120(.A1(new_n545), .A2(G860), .ZN(G153));
  NAND4_X1  g121(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g122(.A1(G1), .A2(G3), .ZN(new_n548));
  XNOR2_X1  g123(.A(new_n548), .B(KEYINPUT8), .ZN(new_n549));
  NAND4_X1  g124(.A1(G319), .A2(G483), .A3(G661), .A4(new_n549), .ZN(new_n550));
  XNOR2_X1  g125(.A(new_n550), .B(KEYINPUT75), .ZN(G188));
  NAND3_X1  g126(.A1(new_n510), .A2(G53), .A3(G543), .ZN(new_n552));
  XOR2_X1   g127(.A(new_n552), .B(KEYINPUT9), .Z(new_n553));
  XNOR2_X1  g128(.A(KEYINPUT76), .B(G65), .ZN(new_n554));
  AOI22_X1  g129(.A1(new_n509), .A2(new_n554), .B1(G78), .B2(G543), .ZN(new_n555));
  INV_X1    g130(.A(G91), .ZN(new_n556));
  OAI22_X1  g131(.A1(new_n555), .A2(new_n516), .B1(new_n556), .B2(new_n525), .ZN(new_n557));
  NOR2_X1   g132(.A1(new_n553), .A2(new_n557), .ZN(new_n558));
  INV_X1    g133(.A(new_n558), .ZN(G299));
  NAND2_X1  g134(.A1(G171), .A2(KEYINPUT77), .ZN(new_n560));
  INV_X1    g135(.A(KEYINPUT77), .ZN(new_n561));
  NAND2_X1  g136(.A1(new_n538), .A2(new_n561), .ZN(new_n562));
  NAND2_X1  g137(.A1(new_n560), .A2(new_n562), .ZN(new_n563));
  INV_X1    g138(.A(new_n563), .ZN(G301));
  INV_X1    g139(.A(G168), .ZN(G286));
  OR2_X1    g140(.A1(new_n518), .A2(KEYINPUT78), .ZN(new_n566));
  NAND2_X1  g141(.A1(new_n518), .A2(KEYINPUT78), .ZN(new_n567));
  AND2_X1   g142(.A1(new_n566), .A2(new_n567), .ZN(G303));
  AND2_X1   g143(.A1(new_n510), .A2(new_n509), .ZN(new_n569));
  NAND2_X1  g144(.A1(new_n569), .A2(G87), .ZN(new_n570));
  AND2_X1   g145(.A1(new_n510), .A2(G543), .ZN(new_n571));
  NAND2_X1  g146(.A1(new_n571), .A2(G49), .ZN(new_n572));
  OAI21_X1  g147(.A(G651), .B1(new_n509), .B2(G74), .ZN(new_n573));
  NAND3_X1  g148(.A1(new_n570), .A2(new_n572), .A3(new_n573), .ZN(G288));
  INV_X1    g149(.A(G86), .ZN(new_n575));
  INV_X1    g150(.A(G48), .ZN(new_n576));
  OAI22_X1  g151(.A1(new_n525), .A2(new_n575), .B1(new_n527), .B2(new_n576), .ZN(new_n577));
  AOI22_X1  g152(.A1(new_n509), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n578));
  NOR2_X1   g153(.A1(new_n578), .A2(new_n516), .ZN(new_n579));
  NOR2_X1   g154(.A1(new_n577), .A2(new_n579), .ZN(new_n580));
  INV_X1    g155(.A(new_n580), .ZN(G305));
  INV_X1    g156(.A(G85), .ZN(new_n582));
  INV_X1    g157(.A(G47), .ZN(new_n583));
  OAI22_X1  g158(.A1(new_n525), .A2(new_n582), .B1(new_n527), .B2(new_n583), .ZN(new_n584));
  OR2_X1    g159(.A1(new_n584), .A2(KEYINPUT80), .ZN(new_n585));
  NAND2_X1  g160(.A1(new_n584), .A2(KEYINPUT80), .ZN(new_n586));
  NAND2_X1  g161(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  AOI22_X1  g162(.A1(new_n509), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n588));
  NOR2_X1   g163(.A1(new_n588), .A2(new_n516), .ZN(new_n589));
  OR2_X1    g164(.A1(new_n589), .A2(KEYINPUT79), .ZN(new_n590));
  NAND2_X1  g165(.A1(new_n589), .A2(KEYINPUT79), .ZN(new_n591));
  NAND2_X1  g166(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  NAND2_X1  g167(.A1(new_n587), .A2(new_n592), .ZN(G290));
  AOI22_X1  g168(.A1(new_n509), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n594));
  INV_X1    g169(.A(G54), .ZN(new_n595));
  OAI22_X1  g170(.A1(new_n594), .A2(new_n516), .B1(new_n595), .B2(new_n527), .ZN(new_n596));
  XNOR2_X1  g171(.A(new_n596), .B(KEYINPUT81), .ZN(new_n597));
  NAND2_X1  g172(.A1(new_n569), .A2(G92), .ZN(new_n598));
  XOR2_X1   g173(.A(new_n598), .B(KEYINPUT10), .Z(new_n599));
  NAND2_X1  g174(.A1(new_n597), .A2(new_n599), .ZN(new_n600));
  NOR2_X1   g175(.A1(new_n600), .A2(G868), .ZN(new_n601));
  AOI21_X1  g176(.A(new_n601), .B1(new_n563), .B2(G868), .ZN(G284));
  AOI21_X1  g177(.A(new_n601), .B1(new_n563), .B2(G868), .ZN(G321));
  NAND2_X1  g178(.A1(G286), .A2(G868), .ZN(new_n604));
  OAI21_X1  g179(.A(new_n604), .B1(G868), .B2(new_n558), .ZN(G297));
  OAI21_X1  g180(.A(new_n604), .B1(G868), .B2(new_n558), .ZN(G280));
  INV_X1    g181(.A(new_n600), .ZN(new_n607));
  INV_X1    g182(.A(G559), .ZN(new_n608));
  OAI21_X1  g183(.A(new_n607), .B1(new_n608), .B2(G860), .ZN(G148));
  INV_X1    g184(.A(new_n545), .ZN(new_n610));
  INV_X1    g185(.A(G868), .ZN(new_n611));
  NAND2_X1  g186(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  NOR2_X1   g187(.A1(new_n600), .A2(G559), .ZN(new_n613));
  OAI21_X1  g188(.A(new_n612), .B1(new_n613), .B2(new_n611), .ZN(G323));
  XNOR2_X1  g189(.A(G323), .B(KEYINPUT11), .ZN(G282));
  OR2_X1    g190(.A1(new_n470), .A2(new_n471), .ZN(new_n616));
  NAND2_X1  g191(.A1(new_n616), .A2(new_n504), .ZN(new_n617));
  XOR2_X1   g192(.A(KEYINPUT82), .B(KEYINPUT12), .Z(new_n618));
  XNOR2_X1  g193(.A(new_n617), .B(new_n618), .ZN(new_n619));
  XOR2_X1   g194(.A(KEYINPUT13), .B(G2100), .Z(new_n620));
  XNOR2_X1  g195(.A(new_n619), .B(new_n620), .ZN(new_n621));
  OAI21_X1  g196(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n622));
  INV_X1    g197(.A(KEYINPUT83), .ZN(new_n623));
  INV_X1    g198(.A(G111), .ZN(new_n624));
  AOI22_X1  g199(.A1(new_n622), .A2(new_n623), .B1(new_n624), .B2(G2105), .ZN(new_n625));
  OAI21_X1  g200(.A(new_n625), .B1(new_n623), .B2(new_n622), .ZN(new_n626));
  INV_X1    g201(.A(G123), .ZN(new_n627));
  OAI21_X1  g202(.A(new_n626), .B1(new_n627), .B2(new_n482), .ZN(new_n628));
  AOI21_X1  g203(.A(new_n628), .B1(new_n488), .B2(G135), .ZN(new_n629));
  INV_X1    g204(.A(G2096), .ZN(new_n630));
  NAND2_X1  g205(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  OR2_X1    g206(.A1(new_n629), .A2(new_n630), .ZN(new_n632));
  NAND3_X1  g207(.A1(new_n621), .A2(new_n631), .A3(new_n632), .ZN(G156));
  XNOR2_X1  g208(.A(G2427), .B(G2430), .ZN(new_n634));
  XNOR2_X1  g209(.A(new_n634), .B(KEYINPUT85), .ZN(new_n635));
  XNOR2_X1  g210(.A(KEYINPUT84), .B(G2438), .ZN(new_n636));
  XNOR2_X1  g211(.A(new_n635), .B(new_n636), .ZN(new_n637));
  XNOR2_X1  g212(.A(KEYINPUT15), .B(G2435), .ZN(new_n638));
  INV_X1    g213(.A(new_n638), .ZN(new_n639));
  OR2_X1    g214(.A1(new_n637), .A2(new_n639), .ZN(new_n640));
  NAND2_X1  g215(.A1(new_n637), .A2(new_n639), .ZN(new_n641));
  NAND3_X1  g216(.A1(new_n640), .A2(KEYINPUT14), .A3(new_n641), .ZN(new_n642));
  XOR2_X1   g217(.A(G2443), .B(G2446), .Z(new_n643));
  XNOR2_X1  g218(.A(new_n642), .B(new_n643), .ZN(new_n644));
  XOR2_X1   g219(.A(G2451), .B(G2454), .Z(new_n645));
  XNOR2_X1  g220(.A(new_n645), .B(KEYINPUT16), .ZN(new_n646));
  XNOR2_X1  g221(.A(new_n646), .B(KEYINPUT86), .ZN(new_n647));
  XNOR2_X1  g222(.A(new_n644), .B(new_n647), .ZN(new_n648));
  XNOR2_X1  g223(.A(G1341), .B(G1348), .ZN(new_n649));
  NOR2_X1   g224(.A1(new_n648), .A2(new_n649), .ZN(new_n650));
  XNOR2_X1  g225(.A(new_n650), .B(KEYINPUT87), .ZN(new_n651));
  NAND2_X1  g226(.A1(new_n648), .A2(new_n649), .ZN(new_n652));
  NAND3_X1  g227(.A1(new_n651), .A2(G14), .A3(new_n652), .ZN(new_n653));
  XNOR2_X1  g228(.A(new_n653), .B(KEYINPUT88), .ZN(G401));
  INV_X1    g229(.A(KEYINPUT18), .ZN(new_n655));
  XOR2_X1   g230(.A(G2084), .B(G2090), .Z(new_n656));
  XNOR2_X1  g231(.A(G2067), .B(G2678), .ZN(new_n657));
  NAND2_X1  g232(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  NAND2_X1  g233(.A1(new_n658), .A2(KEYINPUT17), .ZN(new_n659));
  NOR2_X1   g234(.A1(new_n656), .A2(new_n657), .ZN(new_n660));
  OAI21_X1  g235(.A(new_n655), .B1(new_n659), .B2(new_n660), .ZN(new_n661));
  XNOR2_X1  g236(.A(new_n661), .B(G2100), .ZN(new_n662));
  XOR2_X1   g237(.A(G2072), .B(G2078), .Z(new_n663));
  AOI21_X1  g238(.A(new_n663), .B1(new_n658), .B2(KEYINPUT18), .ZN(new_n664));
  XNOR2_X1  g239(.A(new_n664), .B(G2096), .ZN(new_n665));
  XNOR2_X1  g240(.A(new_n662), .B(new_n665), .ZN(G227));
  XOR2_X1   g241(.A(G1971), .B(G1976), .Z(new_n667));
  XNOR2_X1  g242(.A(new_n667), .B(KEYINPUT19), .ZN(new_n668));
  XOR2_X1   g243(.A(G1956), .B(G2474), .Z(new_n669));
  XOR2_X1   g244(.A(G1961), .B(G1966), .Z(new_n670));
  AND2_X1   g245(.A1(new_n669), .A2(new_n670), .ZN(new_n671));
  NAND2_X1  g246(.A1(new_n668), .A2(new_n671), .ZN(new_n672));
  XNOR2_X1  g247(.A(new_n672), .B(KEYINPUT20), .ZN(new_n673));
  NOR2_X1   g248(.A1(new_n669), .A2(new_n670), .ZN(new_n674));
  NOR3_X1   g249(.A1(new_n668), .A2(new_n671), .A3(new_n674), .ZN(new_n675));
  AOI21_X1  g250(.A(new_n675), .B1(new_n668), .B2(new_n674), .ZN(new_n676));
  NAND2_X1  g251(.A1(new_n673), .A2(new_n676), .ZN(new_n677));
  XNOR2_X1  g252(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n678));
  XNOR2_X1  g253(.A(new_n677), .B(new_n678), .ZN(new_n679));
  XNOR2_X1  g254(.A(G1991), .B(G1996), .ZN(new_n680));
  XNOR2_X1  g255(.A(new_n679), .B(new_n680), .ZN(new_n681));
  XNOR2_X1  g256(.A(G1981), .B(G1986), .ZN(new_n682));
  XNOR2_X1  g257(.A(new_n681), .B(new_n682), .ZN(G229));
  NOR2_X1   g258(.A1(G6), .A2(G16), .ZN(new_n684));
  AOI21_X1  g259(.A(new_n684), .B1(new_n580), .B2(G16), .ZN(new_n685));
  XNOR2_X1  g260(.A(new_n685), .B(KEYINPUT32), .ZN(new_n686));
  INV_X1    g261(.A(G1981), .ZN(new_n687));
  XNOR2_X1  g262(.A(new_n686), .B(new_n687), .ZN(new_n688));
  NAND2_X1  g263(.A1(G166), .A2(G16), .ZN(new_n689));
  OAI21_X1  g264(.A(new_n689), .B1(G16), .B2(G22), .ZN(new_n690));
  INV_X1    g265(.A(G1971), .ZN(new_n691));
  NAND2_X1  g266(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  OR2_X1    g267(.A1(new_n690), .A2(new_n691), .ZN(new_n693));
  INV_X1    g268(.A(G16), .ZN(new_n694));
  NAND2_X1  g269(.A1(new_n694), .A2(G23), .ZN(new_n695));
  INV_X1    g270(.A(G288), .ZN(new_n696));
  OAI21_X1  g271(.A(new_n695), .B1(new_n696), .B2(new_n694), .ZN(new_n697));
  XOR2_X1   g272(.A(KEYINPUT33), .B(G1976), .Z(new_n698));
  XOR2_X1   g273(.A(new_n697), .B(new_n698), .Z(new_n699));
  NAND4_X1  g274(.A1(new_n688), .A2(new_n692), .A3(new_n693), .A4(new_n699), .ZN(new_n700));
  OR2_X1    g275(.A1(new_n700), .A2(KEYINPUT34), .ZN(new_n701));
  NAND2_X1  g276(.A1(new_n700), .A2(KEYINPUT34), .ZN(new_n702));
  NAND2_X1  g277(.A1(new_n694), .A2(G24), .ZN(new_n703));
  INV_X1    g278(.A(G290), .ZN(new_n704));
  OAI21_X1  g279(.A(new_n703), .B1(new_n704), .B2(new_n694), .ZN(new_n705));
  XNOR2_X1  g280(.A(new_n705), .B(G1986), .ZN(new_n706));
  OR2_X1    g281(.A1(G25), .A2(G29), .ZN(new_n707));
  AND2_X1   g282(.A1(new_n493), .A2(G119), .ZN(new_n708));
  XNOR2_X1  g283(.A(new_n708), .B(KEYINPUT89), .ZN(new_n709));
  OAI21_X1  g284(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n710));
  INV_X1    g285(.A(G107), .ZN(new_n711));
  AOI21_X1  g286(.A(new_n710), .B1(new_n711), .B2(G2105), .ZN(new_n712));
  AOI21_X1  g287(.A(new_n712), .B1(new_n488), .B2(G131), .ZN(new_n713));
  NAND2_X1  g288(.A1(new_n709), .A2(new_n713), .ZN(new_n714));
  INV_X1    g289(.A(G29), .ZN(new_n715));
  OAI21_X1  g290(.A(new_n707), .B1(new_n714), .B2(new_n715), .ZN(new_n716));
  XOR2_X1   g291(.A(KEYINPUT35), .B(G1991), .Z(new_n717));
  NOR2_X1   g292(.A1(new_n716), .A2(new_n717), .ZN(new_n718));
  AND2_X1   g293(.A1(new_n716), .A2(new_n717), .ZN(new_n719));
  NOR3_X1   g294(.A1(new_n706), .A2(new_n718), .A3(new_n719), .ZN(new_n720));
  NAND3_X1  g295(.A1(new_n701), .A2(new_n702), .A3(new_n720), .ZN(new_n721));
  XNOR2_X1  g296(.A(new_n721), .B(KEYINPUT36), .ZN(new_n722));
  NOR2_X1   g297(.A1(new_n607), .A2(new_n694), .ZN(new_n723));
  AOI21_X1  g298(.A(new_n723), .B1(G4), .B2(new_n694), .ZN(new_n724));
  INV_X1    g299(.A(new_n724), .ZN(new_n725));
  AND2_X1   g300(.A1(new_n725), .A2(G1348), .ZN(new_n726));
  NOR2_X1   g301(.A1(new_n725), .A2(G1348), .ZN(new_n727));
  INV_X1    g302(.A(KEYINPUT24), .ZN(new_n728));
  OAI21_X1  g303(.A(new_n715), .B1(new_n728), .B2(G34), .ZN(new_n729));
  OR2_X1    g304(.A1(new_n729), .A2(KEYINPUT93), .ZN(new_n730));
  NAND2_X1  g305(.A1(new_n729), .A2(KEYINPUT93), .ZN(new_n731));
  NAND2_X1  g306(.A1(new_n728), .A2(G34), .ZN(new_n732));
  NAND3_X1  g307(.A1(new_n730), .A2(new_n731), .A3(new_n732), .ZN(new_n733));
  OAI21_X1  g308(.A(new_n733), .B1(new_n480), .B2(new_n715), .ZN(new_n734));
  INV_X1    g309(.A(G2084), .ZN(new_n735));
  NOR2_X1   g310(.A1(new_n734), .A2(new_n735), .ZN(new_n736));
  INV_X1    g311(.A(new_n736), .ZN(new_n737));
  NOR2_X1   g312(.A1(new_n737), .A2(KEYINPUT94), .ZN(new_n738));
  NOR3_X1   g313(.A1(new_n726), .A2(new_n727), .A3(new_n738), .ZN(new_n739));
  NAND3_X1  g314(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n740));
  INV_X1    g315(.A(KEYINPUT26), .ZN(new_n741));
  NAND2_X1  g316(.A1(new_n740), .A2(new_n741), .ZN(new_n742));
  OR2_X1    g317(.A1(new_n740), .A2(new_n741), .ZN(new_n743));
  AOI22_X1  g318(.A1(new_n616), .A2(G105), .B1(new_n742), .B2(new_n743), .ZN(new_n744));
  INV_X1    g319(.A(G129), .ZN(new_n745));
  OAI21_X1  g320(.A(new_n744), .B1(new_n745), .B2(new_n482), .ZN(new_n746));
  AND2_X1   g321(.A1(new_n488), .A2(G141), .ZN(new_n747));
  NOR2_X1   g322(.A1(new_n746), .A2(new_n747), .ZN(new_n748));
  XNOR2_X1  g323(.A(new_n748), .B(KEYINPUT95), .ZN(new_n749));
  INV_X1    g324(.A(new_n749), .ZN(new_n750));
  NAND2_X1  g325(.A1(new_n750), .A2(G29), .ZN(new_n751));
  OAI21_X1  g326(.A(new_n751), .B1(G29), .B2(G32), .ZN(new_n752));
  XNOR2_X1  g327(.A(KEYINPUT27), .B(G1996), .ZN(new_n753));
  NOR2_X1   g328(.A1(new_n752), .A2(new_n753), .ZN(new_n754));
  NOR2_X1   g329(.A1(G16), .A2(G19), .ZN(new_n755));
  AOI21_X1  g330(.A(new_n755), .B1(new_n545), .B2(G16), .ZN(new_n756));
  NOR2_X1   g331(.A1(new_n756), .A2(G1341), .ZN(new_n757));
  NOR2_X1   g332(.A1(G168), .A2(new_n694), .ZN(new_n758));
  AOI21_X1  g333(.A(new_n758), .B1(new_n694), .B2(G21), .ZN(new_n759));
  INV_X1    g334(.A(new_n759), .ZN(new_n760));
  AOI21_X1  g335(.A(new_n757), .B1(new_n760), .B2(G1966), .ZN(new_n761));
  NAND2_X1  g336(.A1(new_n737), .A2(KEYINPUT94), .ZN(new_n762));
  INV_X1    g337(.A(KEYINPUT30), .ZN(new_n763));
  AND2_X1   g338(.A1(new_n763), .A2(G28), .ZN(new_n764));
  OAI21_X1  g339(.A(new_n715), .B1(new_n763), .B2(G28), .ZN(new_n765));
  AND2_X1   g340(.A1(KEYINPUT31), .A2(G11), .ZN(new_n766));
  NOR2_X1   g341(.A1(KEYINPUT31), .A2(G11), .ZN(new_n767));
  OAI22_X1  g342(.A1(new_n764), .A2(new_n765), .B1(new_n766), .B2(new_n767), .ZN(new_n768));
  INV_X1    g343(.A(G1966), .ZN(new_n769));
  AOI21_X1  g344(.A(new_n768), .B1(new_n759), .B2(new_n769), .ZN(new_n770));
  AOI22_X1  g345(.A1(new_n756), .A2(G1341), .B1(G29), .B2(new_n629), .ZN(new_n771));
  NAND4_X1  g346(.A1(new_n761), .A2(new_n762), .A3(new_n770), .A4(new_n771), .ZN(new_n772));
  NAND2_X1  g347(.A1(new_n694), .A2(G20), .ZN(new_n773));
  XOR2_X1   g348(.A(new_n773), .B(KEYINPUT23), .Z(new_n774));
  AOI21_X1  g349(.A(new_n774), .B1(G299), .B2(G16), .ZN(new_n775));
  XNOR2_X1  g350(.A(new_n775), .B(G1956), .ZN(new_n776));
  NAND2_X1  g351(.A1(new_n715), .A2(G27), .ZN(new_n777));
  OAI21_X1  g352(.A(new_n777), .B1(G164), .B2(new_n715), .ZN(new_n778));
  INV_X1    g353(.A(G2078), .ZN(new_n779));
  XNOR2_X1  g354(.A(new_n778), .B(new_n779), .ZN(new_n780));
  NAND2_X1  g355(.A1(new_n734), .A2(new_n735), .ZN(new_n781));
  NAND3_X1  g356(.A1(new_n776), .A2(new_n780), .A3(new_n781), .ZN(new_n782));
  AND2_X1   g357(.A1(new_n715), .A2(G33), .ZN(new_n783));
  NAND3_X1  g358(.A1(new_n466), .A2(G103), .A3(G2104), .ZN(new_n784));
  XNOR2_X1  g359(.A(new_n784), .B(KEYINPUT92), .ZN(new_n785));
  XNOR2_X1  g360(.A(new_n785), .B(KEYINPUT25), .ZN(new_n786));
  NAND2_X1  g361(.A1(new_n488), .A2(G139), .ZN(new_n787));
  AOI22_X1  g362(.A1(new_n504), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n788));
  OAI211_X1 g363(.A(new_n786), .B(new_n787), .C1(new_n466), .C2(new_n788), .ZN(new_n789));
  AOI21_X1  g364(.A(new_n783), .B1(new_n789), .B2(G29), .ZN(new_n790));
  INV_X1    g365(.A(new_n790), .ZN(new_n791));
  OR2_X1    g366(.A1(new_n791), .A2(G2072), .ZN(new_n792));
  NOR2_X1   g367(.A1(G5), .A2(G16), .ZN(new_n793));
  XOR2_X1   g368(.A(new_n793), .B(KEYINPUT97), .Z(new_n794));
  OAI21_X1  g369(.A(new_n794), .B1(new_n538), .B2(new_n694), .ZN(new_n795));
  INV_X1    g370(.A(G1961), .ZN(new_n796));
  OR2_X1    g371(.A1(new_n795), .A2(new_n796), .ZN(new_n797));
  NAND2_X1  g372(.A1(new_n795), .A2(new_n796), .ZN(new_n798));
  NAND2_X1  g373(.A1(new_n791), .A2(G2072), .ZN(new_n799));
  NAND4_X1  g374(.A1(new_n792), .A2(new_n797), .A3(new_n798), .A4(new_n799), .ZN(new_n800));
  NOR4_X1   g375(.A1(new_n754), .A2(new_n772), .A3(new_n782), .A4(new_n800), .ZN(new_n801));
  NAND2_X1  g376(.A1(new_n752), .A2(new_n753), .ZN(new_n802));
  XOR2_X1   g377(.A(new_n802), .B(KEYINPUT96), .Z(new_n803));
  XOR2_X1   g378(.A(KEYINPUT91), .B(KEYINPUT28), .Z(new_n804));
  NAND2_X1  g379(.A1(new_n715), .A2(G26), .ZN(new_n805));
  XNOR2_X1  g380(.A(new_n804), .B(new_n805), .ZN(new_n806));
  INV_X1    g381(.A(G140), .ZN(new_n807));
  NOR2_X1   g382(.A1(new_n487), .A2(new_n807), .ZN(new_n808));
  XNOR2_X1  g383(.A(new_n808), .B(KEYINPUT90), .ZN(new_n809));
  OAI21_X1  g384(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n810));
  INV_X1    g385(.A(G116), .ZN(new_n811));
  AOI21_X1  g386(.A(new_n810), .B1(new_n811), .B2(G2105), .ZN(new_n812));
  AOI21_X1  g387(.A(new_n812), .B1(new_n493), .B2(G128), .ZN(new_n813));
  AND2_X1   g388(.A1(new_n809), .A2(new_n813), .ZN(new_n814));
  OAI21_X1  g389(.A(new_n806), .B1(new_n814), .B2(new_n715), .ZN(new_n815));
  XNOR2_X1  g390(.A(new_n815), .B(G2067), .ZN(new_n816));
  NAND2_X1  g391(.A1(new_n715), .A2(G35), .ZN(new_n817));
  OAI21_X1  g392(.A(new_n817), .B1(G162), .B2(new_n715), .ZN(new_n818));
  XNOR2_X1  g393(.A(new_n818), .B(KEYINPUT29), .ZN(new_n819));
  XNOR2_X1  g394(.A(new_n819), .B(G2090), .ZN(new_n820));
  NOR3_X1   g395(.A1(new_n803), .A2(new_n816), .A3(new_n820), .ZN(new_n821));
  NAND4_X1  g396(.A1(new_n722), .A2(new_n739), .A3(new_n801), .A4(new_n821), .ZN(G150));
  INV_X1    g397(.A(G150), .ZN(G311));
  XNOR2_X1  g398(.A(KEYINPUT98), .B(G93), .ZN(new_n824));
  AOI22_X1  g399(.A1(new_n569), .A2(new_n824), .B1(new_n571), .B2(G55), .ZN(new_n825));
  AOI22_X1  g400(.A1(new_n509), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n826));
  OR2_X1    g401(.A1(new_n826), .A2(new_n516), .ZN(new_n827));
  NAND2_X1  g402(.A1(new_n825), .A2(new_n827), .ZN(new_n828));
  NAND2_X1  g403(.A1(new_n828), .A2(KEYINPUT99), .ZN(new_n829));
  INV_X1    g404(.A(KEYINPUT99), .ZN(new_n830));
  NAND3_X1  g405(.A1(new_n825), .A2(new_n830), .A3(new_n827), .ZN(new_n831));
  AOI21_X1  g406(.A(new_n545), .B1(new_n829), .B2(new_n831), .ZN(new_n832));
  NOR2_X1   g407(.A1(new_n610), .A2(new_n828), .ZN(new_n833));
  NOR2_X1   g408(.A1(new_n832), .A2(new_n833), .ZN(new_n834));
  XNOR2_X1  g409(.A(new_n834), .B(KEYINPUT38), .ZN(new_n835));
  NAND2_X1  g410(.A1(new_n607), .A2(G559), .ZN(new_n836));
  XNOR2_X1  g411(.A(new_n835), .B(new_n836), .ZN(new_n837));
  AND2_X1   g412(.A1(new_n837), .A2(KEYINPUT39), .ZN(new_n838));
  NOR2_X1   g413(.A1(new_n837), .A2(KEYINPUT39), .ZN(new_n839));
  NOR3_X1   g414(.A1(new_n838), .A2(new_n839), .A3(G860), .ZN(new_n840));
  NAND2_X1  g415(.A1(new_n829), .A2(new_n831), .ZN(new_n841));
  NAND2_X1  g416(.A1(new_n841), .A2(G860), .ZN(new_n842));
  XNOR2_X1  g417(.A(new_n842), .B(KEYINPUT101), .ZN(new_n843));
  XNOR2_X1  g418(.A(new_n843), .B(KEYINPUT100), .ZN(new_n844));
  XNOR2_X1  g419(.A(new_n844), .B(KEYINPUT37), .ZN(new_n845));
  OR2_X1    g420(.A1(new_n840), .A2(new_n845), .ZN(G145));
  XNOR2_X1  g421(.A(new_n480), .B(new_n629), .ZN(new_n847));
  XNOR2_X1  g422(.A(new_n847), .B(G162), .ZN(new_n848));
  XNOR2_X1  g423(.A(new_n814), .B(new_n507), .ZN(new_n849));
  XNOR2_X1  g424(.A(new_n849), .B(new_n619), .ZN(new_n850));
  OAI21_X1  g425(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n851));
  INV_X1    g426(.A(G118), .ZN(new_n852));
  AOI21_X1  g427(.A(new_n851), .B1(new_n852), .B2(G2105), .ZN(new_n853));
  NAND2_X1  g428(.A1(new_n488), .A2(G142), .ZN(new_n854));
  XNOR2_X1  g429(.A(new_n854), .B(KEYINPUT102), .ZN(new_n855));
  AOI211_X1 g430(.A(new_n853), .B(new_n855), .C1(G130), .C2(new_n493), .ZN(new_n856));
  XOR2_X1   g431(.A(new_n856), .B(new_n714), .Z(new_n857));
  XNOR2_X1  g432(.A(new_n850), .B(new_n857), .ZN(new_n858));
  NAND2_X1  g433(.A1(new_n789), .A2(new_n748), .ZN(new_n859));
  OAI21_X1  g434(.A(new_n859), .B1(new_n750), .B2(new_n789), .ZN(new_n860));
  INV_X1    g435(.A(new_n860), .ZN(new_n861));
  NAND2_X1  g436(.A1(new_n858), .A2(new_n861), .ZN(new_n862));
  INV_X1    g437(.A(new_n862), .ZN(new_n863));
  NOR2_X1   g438(.A1(new_n858), .A2(new_n861), .ZN(new_n864));
  OAI21_X1  g439(.A(new_n848), .B1(new_n863), .B2(new_n864), .ZN(new_n865));
  INV_X1    g440(.A(G37), .ZN(new_n866));
  OR2_X1    g441(.A1(new_n858), .A2(new_n861), .ZN(new_n867));
  INV_X1    g442(.A(new_n848), .ZN(new_n868));
  NAND3_X1  g443(.A1(new_n867), .A2(new_n868), .A3(new_n862), .ZN(new_n869));
  NAND3_X1  g444(.A1(new_n865), .A2(new_n866), .A3(new_n869), .ZN(new_n870));
  XNOR2_X1  g445(.A(new_n870), .B(KEYINPUT40), .ZN(G395));
  NAND2_X1  g446(.A1(new_n841), .A2(new_n611), .ZN(new_n872));
  NAND2_X1  g447(.A1(new_n600), .A2(new_n558), .ZN(new_n873));
  INV_X1    g448(.A(new_n873), .ZN(new_n874));
  NOR2_X1   g449(.A1(new_n600), .A2(new_n558), .ZN(new_n875));
  NOR2_X1   g450(.A1(new_n874), .A2(new_n875), .ZN(new_n876));
  INV_X1    g451(.A(KEYINPUT41), .ZN(new_n877));
  NOR3_X1   g452(.A1(new_n874), .A2(new_n877), .A3(new_n875), .ZN(new_n878));
  AOI21_X1  g453(.A(new_n875), .B1(KEYINPUT103), .B2(new_n873), .ZN(new_n879));
  INV_X1    g454(.A(KEYINPUT103), .ZN(new_n880));
  NAND3_X1  g455(.A1(new_n600), .A2(new_n880), .A3(new_n558), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n879), .A2(new_n881), .ZN(new_n882));
  AOI21_X1  g457(.A(new_n878), .B1(new_n882), .B2(new_n877), .ZN(new_n883));
  XOR2_X1   g458(.A(new_n834), .B(new_n613), .Z(new_n884));
  MUX2_X1   g459(.A(new_n876), .B(new_n883), .S(new_n884), .Z(new_n885));
  NAND2_X1  g460(.A1(new_n704), .A2(new_n518), .ZN(new_n886));
  NAND2_X1  g461(.A1(G290), .A2(G166), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n886), .A2(new_n887), .ZN(new_n888));
  XNOR2_X1  g463(.A(new_n696), .B(new_n580), .ZN(new_n889));
  INV_X1    g464(.A(new_n889), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n888), .A2(new_n890), .ZN(new_n891));
  NAND3_X1  g466(.A1(new_n886), .A2(new_n889), .A3(new_n887), .ZN(new_n892));
  NAND2_X1  g467(.A1(new_n891), .A2(new_n892), .ZN(new_n893));
  XOR2_X1   g468(.A(new_n893), .B(KEYINPUT42), .Z(new_n894));
  XNOR2_X1  g469(.A(new_n885), .B(new_n894), .ZN(new_n895));
  OAI21_X1  g470(.A(new_n872), .B1(new_n895), .B2(new_n611), .ZN(G295));
  OAI21_X1  g471(.A(new_n872), .B1(new_n895), .B2(new_n611), .ZN(G331));
  NAND2_X1  g472(.A1(new_n834), .A2(KEYINPUT104), .ZN(new_n898));
  INV_X1    g473(.A(KEYINPUT104), .ZN(new_n899));
  OAI21_X1  g474(.A(new_n899), .B1(new_n832), .B2(new_n833), .ZN(new_n900));
  NAND2_X1  g475(.A1(new_n898), .A2(new_n900), .ZN(new_n901));
  NAND2_X1  g476(.A1(new_n563), .A2(G168), .ZN(new_n902));
  NOR2_X1   g477(.A1(G171), .A2(G168), .ZN(new_n903));
  INV_X1    g478(.A(new_n903), .ZN(new_n904));
  NAND3_X1  g479(.A1(new_n901), .A2(new_n902), .A3(new_n904), .ZN(new_n905));
  AOI21_X1  g480(.A(G286), .B1(new_n560), .B2(new_n562), .ZN(new_n906));
  OAI211_X1 g481(.A(new_n898), .B(new_n900), .C1(new_n906), .C2(new_n903), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n905), .A2(new_n907), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n908), .A2(new_n883), .ZN(new_n909));
  AND3_X1   g484(.A1(new_n891), .A2(KEYINPUT105), .A3(new_n892), .ZN(new_n910));
  AOI21_X1  g485(.A(KEYINPUT105), .B1(new_n891), .B2(new_n892), .ZN(new_n911));
  NOR2_X1   g486(.A1(new_n910), .A2(new_n911), .ZN(new_n912));
  NAND3_X1  g487(.A1(new_n905), .A2(new_n907), .A3(new_n876), .ZN(new_n913));
  AND3_X1   g488(.A1(new_n909), .A2(new_n912), .A3(new_n913), .ZN(new_n914));
  AOI22_X1  g489(.A1(new_n909), .A2(new_n913), .B1(new_n892), .B2(new_n891), .ZN(new_n915));
  NOR3_X1   g490(.A1(new_n914), .A2(new_n915), .A3(G37), .ZN(new_n916));
  NOR2_X1   g491(.A1(new_n916), .A2(KEYINPUT43), .ZN(new_n917));
  NOR2_X1   g492(.A1(new_n915), .A2(G37), .ZN(new_n918));
  NAND3_X1  g493(.A1(new_n908), .A2(KEYINPUT41), .A3(new_n882), .ZN(new_n919));
  INV_X1    g494(.A(new_n876), .ZN(new_n920));
  AOI21_X1  g495(.A(new_n877), .B1(new_n905), .B2(new_n907), .ZN(new_n921));
  OAI211_X1 g496(.A(new_n919), .B(new_n912), .C1(new_n920), .C2(new_n921), .ZN(new_n922));
  AND3_X1   g497(.A1(new_n918), .A2(KEYINPUT43), .A3(new_n922), .ZN(new_n923));
  OAI21_X1  g498(.A(KEYINPUT44), .B1(new_n917), .B2(new_n923), .ZN(new_n924));
  INV_X1    g499(.A(KEYINPUT43), .ZN(new_n925));
  OAI21_X1  g500(.A(KEYINPUT106), .B1(new_n916), .B2(new_n925), .ZN(new_n926));
  INV_X1    g501(.A(KEYINPUT106), .ZN(new_n927));
  NAND2_X1  g502(.A1(new_n909), .A2(new_n913), .ZN(new_n928));
  NAND2_X1  g503(.A1(new_n928), .A2(new_n893), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n929), .A2(new_n866), .ZN(new_n930));
  OAI211_X1 g505(.A(new_n927), .B(KEYINPUT43), .C1(new_n930), .C2(new_n914), .ZN(new_n931));
  NAND4_X1  g506(.A1(new_n929), .A2(new_n922), .A3(new_n925), .A4(new_n866), .ZN(new_n932));
  NAND2_X1  g507(.A1(new_n932), .A2(KEYINPUT107), .ZN(new_n933));
  INV_X1    g508(.A(KEYINPUT107), .ZN(new_n934));
  NAND4_X1  g509(.A1(new_n918), .A2(new_n934), .A3(new_n925), .A4(new_n922), .ZN(new_n935));
  AOI22_X1  g510(.A1(new_n926), .A2(new_n931), .B1(new_n933), .B2(new_n935), .ZN(new_n936));
  OAI21_X1  g511(.A(new_n924), .B1(new_n936), .B2(KEYINPUT44), .ZN(G397));
  INV_X1    g512(.A(G1384), .ZN(new_n938));
  AOI22_X1  g513(.A1(KEYINPUT4), .A2(new_n497), .B1(new_n503), .B2(new_n504), .ZN(new_n939));
  INV_X1    g514(.A(G126), .ZN(new_n940));
  OAI22_X1  g515(.A1(new_n482), .A2(new_n940), .B1(new_n490), .B2(new_n491), .ZN(new_n941));
  OAI21_X1  g516(.A(new_n938), .B1(new_n939), .B2(new_n941), .ZN(new_n942));
  INV_X1    g517(.A(KEYINPUT45), .ZN(new_n943));
  NAND2_X1  g518(.A1(new_n942), .A2(new_n943), .ZN(new_n944));
  NAND4_X1  g519(.A1(new_n468), .A2(new_n479), .A3(G40), .A4(new_n472), .ZN(new_n945));
  NOR2_X1   g520(.A1(new_n944), .A2(new_n945), .ZN(new_n946));
  XOR2_X1   g521(.A(new_n946), .B(KEYINPUT109), .Z(new_n947));
  INV_X1    g522(.A(G2067), .ZN(new_n948));
  XNOR2_X1  g523(.A(new_n814), .B(new_n948), .ZN(new_n949));
  INV_X1    g524(.A(new_n748), .ZN(new_n950));
  OAI21_X1  g525(.A(new_n947), .B1(new_n949), .B2(new_n950), .ZN(new_n951));
  INV_X1    g526(.A(G1996), .ZN(new_n952));
  NAND2_X1  g527(.A1(new_n946), .A2(new_n952), .ZN(new_n953));
  XNOR2_X1  g528(.A(new_n953), .B(KEYINPUT46), .ZN(new_n954));
  NAND2_X1  g529(.A1(new_n951), .A2(new_n954), .ZN(new_n955));
  XOR2_X1   g530(.A(new_n955), .B(KEYINPUT47), .Z(new_n956));
  INV_X1    g531(.A(new_n947), .ZN(new_n957));
  NOR2_X1   g532(.A1(new_n749), .A2(new_n953), .ZN(new_n958));
  XNOR2_X1  g533(.A(new_n958), .B(KEYINPUT108), .ZN(new_n959));
  NOR2_X1   g534(.A1(new_n748), .A2(new_n952), .ZN(new_n960));
  OAI21_X1  g535(.A(new_n947), .B1(new_n949), .B2(new_n960), .ZN(new_n961));
  AND2_X1   g536(.A1(new_n959), .A2(new_n961), .ZN(new_n962));
  NAND4_X1  g537(.A1(new_n962), .A2(new_n709), .A3(new_n713), .A4(new_n717), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n814), .A2(new_n948), .ZN(new_n964));
  AOI21_X1  g539(.A(new_n957), .B1(new_n963), .B2(new_n964), .ZN(new_n965));
  XNOR2_X1  g540(.A(new_n714), .B(new_n717), .ZN(new_n966));
  XOR2_X1   g541(.A(new_n966), .B(KEYINPUT110), .Z(new_n967));
  NAND2_X1  g542(.A1(new_n967), .A2(new_n947), .ZN(new_n968));
  NAND2_X1  g543(.A1(new_n962), .A2(new_n968), .ZN(new_n969));
  INV_X1    g544(.A(new_n969), .ZN(new_n970));
  INV_X1    g545(.A(new_n946), .ZN(new_n971));
  NOR3_X1   g546(.A1(new_n971), .A2(G1986), .A3(G290), .ZN(new_n972));
  XOR2_X1   g547(.A(new_n972), .B(KEYINPUT48), .Z(new_n973));
  AOI211_X1 g548(.A(new_n956), .B(new_n965), .C1(new_n970), .C2(new_n973), .ZN(new_n974));
  AOI21_X1  g549(.A(G1384), .B1(new_n494), .B2(new_n506), .ZN(new_n975));
  AND4_X1   g550(.A1(G40), .A2(new_n468), .A3(new_n479), .A4(new_n472), .ZN(new_n976));
  NAND2_X1  g551(.A1(new_n975), .A2(new_n976), .ZN(new_n977));
  NAND2_X1  g552(.A1(new_n977), .A2(G8), .ZN(new_n978));
  INV_X1    g553(.A(new_n978), .ZN(new_n979));
  INV_X1    g554(.A(KEYINPUT49), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n580), .A2(new_n687), .ZN(new_n981));
  INV_X1    g556(.A(new_n981), .ZN(new_n982));
  NOR2_X1   g557(.A1(new_n580), .A2(new_n687), .ZN(new_n983));
  OAI21_X1  g558(.A(new_n980), .B1(new_n982), .B2(new_n983), .ZN(new_n984));
  NAND2_X1  g559(.A1(G305), .A2(G1981), .ZN(new_n985));
  NAND3_X1  g560(.A1(new_n985), .A2(KEYINPUT49), .A3(new_n981), .ZN(new_n986));
  NAND3_X1  g561(.A1(new_n979), .A2(new_n984), .A3(new_n986), .ZN(new_n987));
  INV_X1    g562(.A(G1976), .ZN(new_n988));
  NAND3_X1  g563(.A1(new_n987), .A2(new_n988), .A3(new_n696), .ZN(new_n989));
  NAND2_X1  g564(.A1(new_n989), .A2(new_n981), .ZN(new_n990));
  INV_X1    g565(.A(KEYINPUT115), .ZN(new_n991));
  NAND2_X1  g566(.A1(new_n990), .A2(new_n991), .ZN(new_n992));
  NAND2_X1  g567(.A1(new_n992), .A2(new_n979), .ZN(new_n993));
  NOR2_X1   g568(.A1(new_n990), .A2(new_n991), .ZN(new_n994));
  NAND2_X1  g569(.A1(new_n696), .A2(G1976), .ZN(new_n995));
  AOI21_X1  g570(.A(KEYINPUT52), .B1(G288), .B2(new_n988), .ZN(new_n996));
  NAND3_X1  g571(.A1(new_n979), .A2(new_n995), .A3(new_n996), .ZN(new_n997));
  NAND3_X1  g572(.A1(new_n977), .A2(new_n995), .A3(G8), .ZN(new_n998));
  NAND2_X1  g573(.A1(new_n998), .A2(KEYINPUT52), .ZN(new_n999));
  NAND3_X1  g574(.A1(new_n987), .A2(new_n997), .A3(new_n999), .ZN(new_n1000));
  INV_X1    g575(.A(KEYINPUT114), .ZN(new_n1001));
  NAND2_X1  g576(.A1(new_n1000), .A2(new_n1001), .ZN(new_n1002));
  NAND4_X1  g577(.A1(new_n987), .A2(new_n997), .A3(KEYINPUT114), .A4(new_n999), .ZN(new_n1003));
  AND2_X1   g578(.A1(new_n1002), .A2(new_n1003), .ZN(new_n1004));
  OAI211_X1 g579(.A(KEYINPUT45), .B(new_n938), .C1(new_n939), .C2(new_n941), .ZN(new_n1005));
  NAND3_X1  g580(.A1(new_n944), .A2(new_n976), .A3(new_n1005), .ZN(new_n1006));
  NAND2_X1  g581(.A1(new_n1006), .A2(KEYINPUT111), .ZN(new_n1007));
  INV_X1    g582(.A(KEYINPUT111), .ZN(new_n1008));
  NAND4_X1  g583(.A1(new_n944), .A2(new_n1008), .A3(new_n976), .A4(new_n1005), .ZN(new_n1009));
  NAND3_X1  g584(.A1(new_n1007), .A2(new_n691), .A3(new_n1009), .ZN(new_n1010));
  OAI21_X1  g585(.A(new_n976), .B1(new_n942), .B2(KEYINPUT50), .ZN(new_n1011));
  INV_X1    g586(.A(KEYINPUT112), .ZN(new_n1012));
  INV_X1    g587(.A(KEYINPUT50), .ZN(new_n1013));
  OAI21_X1  g588(.A(new_n1012), .B1(new_n975), .B2(new_n1013), .ZN(new_n1014));
  NAND3_X1  g589(.A1(new_n942), .A2(KEYINPUT112), .A3(KEYINPUT50), .ZN(new_n1015));
  AOI21_X1  g590(.A(new_n1011), .B1(new_n1014), .B2(new_n1015), .ZN(new_n1016));
  INV_X1    g591(.A(G2090), .ZN(new_n1017));
  NAND2_X1  g592(.A1(new_n1016), .A2(new_n1017), .ZN(new_n1018));
  NAND2_X1  g593(.A1(new_n1010), .A2(new_n1018), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n1019), .A2(KEYINPUT113), .ZN(new_n1020));
  NAND3_X1  g595(.A1(new_n566), .A2(G8), .A3(new_n567), .ZN(new_n1021));
  INV_X1    g596(.A(KEYINPUT55), .ZN(new_n1022));
  XNOR2_X1  g597(.A(new_n1021), .B(new_n1022), .ZN(new_n1023));
  INV_X1    g598(.A(KEYINPUT113), .ZN(new_n1024));
  NAND3_X1  g599(.A1(new_n1010), .A2(new_n1018), .A3(new_n1024), .ZN(new_n1025));
  NAND4_X1  g600(.A1(new_n1020), .A2(G8), .A3(new_n1023), .A4(new_n1025), .ZN(new_n1026));
  OAI22_X1  g601(.A1(new_n993), .A2(new_n994), .B1(new_n1004), .B2(new_n1026), .ZN(new_n1027));
  INV_X1    g602(.A(KEYINPUT63), .ZN(new_n1028));
  AOI21_X1  g603(.A(new_n945), .B1(new_n975), .B2(new_n1013), .ZN(new_n1029));
  OAI211_X1 g604(.A(new_n1029), .B(new_n1017), .C1(new_n1013), .C2(new_n975), .ZN(new_n1030));
  NAND2_X1  g605(.A1(new_n1010), .A2(new_n1030), .ZN(new_n1031));
  NAND2_X1  g606(.A1(new_n1031), .A2(G8), .ZN(new_n1032));
  XNOR2_X1  g607(.A(new_n1021), .B(KEYINPUT55), .ZN(new_n1033));
  AOI21_X1  g608(.A(new_n1000), .B1(new_n1032), .B2(new_n1033), .ZN(new_n1034));
  NAND2_X1  g609(.A1(new_n1034), .A2(new_n1026), .ZN(new_n1035));
  INV_X1    g610(.A(G8), .ZN(new_n1036));
  NOR2_X1   g611(.A1(G286), .A2(new_n1036), .ZN(new_n1037));
  NAND2_X1  g612(.A1(new_n1006), .A2(new_n769), .ZN(new_n1038));
  AND3_X1   g613(.A1(new_n942), .A2(KEYINPUT112), .A3(KEYINPUT50), .ZN(new_n1039));
  AOI21_X1  g614(.A(KEYINPUT112), .B1(new_n942), .B2(KEYINPUT50), .ZN(new_n1040));
  OAI211_X1 g615(.A(new_n735), .B(new_n1029), .C1(new_n1039), .C2(new_n1040), .ZN(new_n1041));
  INV_X1    g616(.A(KEYINPUT116), .ZN(new_n1042));
  OAI21_X1  g617(.A(new_n1038), .B1(new_n1041), .B2(new_n1042), .ZN(new_n1043));
  AOI21_X1  g618(.A(KEYINPUT116), .B1(new_n1016), .B2(new_n735), .ZN(new_n1044));
  OAI211_X1 g619(.A(KEYINPUT117), .B(new_n1037), .C1(new_n1043), .C2(new_n1044), .ZN(new_n1045));
  INV_X1    g620(.A(new_n1045), .ZN(new_n1046));
  NAND2_X1  g621(.A1(new_n1041), .A2(new_n1042), .ZN(new_n1047));
  NAND2_X1  g622(.A1(new_n1014), .A2(new_n1015), .ZN(new_n1048));
  NAND4_X1  g623(.A1(new_n1048), .A2(KEYINPUT116), .A3(new_n735), .A4(new_n1029), .ZN(new_n1049));
  NAND3_X1  g624(.A1(new_n1047), .A2(new_n1038), .A3(new_n1049), .ZN(new_n1050));
  AOI21_X1  g625(.A(KEYINPUT117), .B1(new_n1050), .B2(new_n1037), .ZN(new_n1051));
  NOR2_X1   g626(.A1(new_n1046), .A2(new_n1051), .ZN(new_n1052));
  OAI21_X1  g627(.A(new_n1028), .B1(new_n1035), .B2(new_n1052), .ZN(new_n1053));
  NAND2_X1  g628(.A1(new_n1050), .A2(new_n1037), .ZN(new_n1054));
  INV_X1    g629(.A(KEYINPUT117), .ZN(new_n1055));
  NAND2_X1  g630(.A1(new_n1054), .A2(new_n1055), .ZN(new_n1056));
  NAND2_X1  g631(.A1(new_n1056), .A2(new_n1045), .ZN(new_n1057));
  AOI21_X1  g632(.A(new_n1028), .B1(new_n1002), .B2(new_n1003), .ZN(new_n1058));
  NAND2_X1  g633(.A1(new_n1025), .A2(G8), .ZN(new_n1059));
  AOI21_X1  g634(.A(new_n1024), .B1(new_n1010), .B2(new_n1018), .ZN(new_n1060));
  OAI21_X1  g635(.A(new_n1033), .B1(new_n1059), .B2(new_n1060), .ZN(new_n1061));
  NAND4_X1  g636(.A1(new_n1057), .A2(new_n1058), .A3(new_n1061), .A4(new_n1026), .ZN(new_n1062));
  AOI21_X1  g637(.A(new_n1027), .B1(new_n1053), .B2(new_n1062), .ZN(new_n1063));
  INV_X1    g638(.A(KEYINPUT51), .ZN(new_n1064));
  NOR2_X1   g639(.A1(new_n1043), .A2(new_n1044), .ZN(new_n1065));
  AOI21_X1  g640(.A(new_n1036), .B1(new_n1065), .B2(G168), .ZN(new_n1066));
  NAND2_X1  g641(.A1(new_n1050), .A2(G286), .ZN(new_n1067));
  AOI21_X1  g642(.A(new_n1064), .B1(new_n1066), .B2(new_n1067), .ZN(new_n1068));
  OAI21_X1  g643(.A(G8), .B1(new_n1050), .B2(G286), .ZN(new_n1069));
  NOR2_X1   g644(.A1(new_n1069), .A2(KEYINPUT51), .ZN(new_n1070));
  OAI21_X1  g645(.A(KEYINPUT62), .B1(new_n1068), .B2(new_n1070), .ZN(new_n1071));
  INV_X1    g646(.A(new_n1067), .ZN(new_n1072));
  OAI21_X1  g647(.A(KEYINPUT51), .B1(new_n1072), .B2(new_n1069), .ZN(new_n1073));
  INV_X1    g648(.A(KEYINPUT62), .ZN(new_n1074));
  NAND2_X1  g649(.A1(new_n1066), .A2(new_n1064), .ZN(new_n1075));
  NAND3_X1  g650(.A1(new_n1073), .A2(new_n1074), .A3(new_n1075), .ZN(new_n1076));
  OR2_X1    g651(.A1(new_n1016), .A2(G1961), .ZN(new_n1077));
  AND2_X1   g652(.A1(new_n944), .A2(new_n1005), .ZN(new_n1078));
  NAND4_X1  g653(.A1(new_n1078), .A2(KEYINPUT53), .A3(new_n779), .A4(new_n976), .ZN(new_n1079));
  AOI21_X1  g654(.A(G2078), .B1(new_n1007), .B2(new_n1009), .ZN(new_n1080));
  OAI211_X1 g655(.A(new_n1077), .B(new_n1079), .C1(new_n1080), .C2(KEYINPUT53), .ZN(new_n1081));
  AND2_X1   g656(.A1(new_n1081), .A2(new_n563), .ZN(new_n1082));
  AND3_X1   g657(.A1(new_n1082), .A2(new_n1026), .A3(new_n1034), .ZN(new_n1083));
  NAND3_X1  g658(.A1(new_n1071), .A2(new_n1076), .A3(new_n1083), .ZN(new_n1084));
  XNOR2_X1  g659(.A(KEYINPUT56), .B(G2072), .ZN(new_n1085));
  NAND3_X1  g660(.A1(new_n1078), .A2(new_n976), .A3(new_n1085), .ZN(new_n1086));
  OR2_X1    g661(.A1(G299), .A2(KEYINPUT57), .ZN(new_n1087));
  NAND2_X1  g662(.A1(G299), .A2(KEYINPUT57), .ZN(new_n1088));
  INV_X1    g663(.A(G1956), .ZN(new_n1089));
  NOR2_X1   g664(.A1(new_n975), .A2(new_n1013), .ZN(new_n1090));
  OAI21_X1  g665(.A(new_n1089), .B1(new_n1011), .B2(new_n1090), .ZN(new_n1091));
  NAND4_X1  g666(.A1(new_n1086), .A2(new_n1087), .A3(new_n1088), .A4(new_n1091), .ZN(new_n1092));
  INV_X1    g667(.A(new_n1092), .ZN(new_n1093));
  OAI22_X1  g668(.A1(new_n1016), .A2(G1348), .B1(G2067), .B2(new_n977), .ZN(new_n1094));
  XNOR2_X1  g669(.A(new_n1094), .B(KEYINPUT118), .ZN(new_n1095));
  NAND2_X1  g670(.A1(new_n1095), .A2(new_n607), .ZN(new_n1096));
  NAND2_X1  g671(.A1(new_n1086), .A2(new_n1091), .ZN(new_n1097));
  NAND2_X1  g672(.A1(new_n1087), .A2(new_n1088), .ZN(new_n1098));
  NAND2_X1  g673(.A1(new_n1097), .A2(new_n1098), .ZN(new_n1099));
  NAND2_X1  g674(.A1(new_n1099), .A2(KEYINPUT119), .ZN(new_n1100));
  INV_X1    g675(.A(KEYINPUT119), .ZN(new_n1101));
  NAND3_X1  g676(.A1(new_n1097), .A2(new_n1098), .A3(new_n1101), .ZN(new_n1102));
  AND2_X1   g677(.A1(new_n1100), .A2(new_n1102), .ZN(new_n1103));
  AOI21_X1  g678(.A(new_n1093), .B1(new_n1096), .B2(new_n1103), .ZN(new_n1104));
  NAND4_X1  g679(.A1(new_n1100), .A2(KEYINPUT61), .A3(new_n1102), .A4(new_n1092), .ZN(new_n1105));
  NAND2_X1  g680(.A1(new_n1099), .A2(new_n1092), .ZN(new_n1106));
  XOR2_X1   g681(.A(KEYINPUT121), .B(KEYINPUT61), .Z(new_n1107));
  NAND2_X1  g682(.A1(new_n1106), .A2(new_n1107), .ZN(new_n1108));
  NAND2_X1  g683(.A1(new_n1105), .A2(new_n1108), .ZN(new_n1109));
  NAND4_X1  g684(.A1(new_n944), .A2(new_n952), .A3(new_n976), .A4(new_n1005), .ZN(new_n1110));
  INV_X1    g685(.A(KEYINPUT120), .ZN(new_n1111));
  OR2_X1    g686(.A1(new_n1110), .A2(new_n1111), .ZN(new_n1112));
  XOR2_X1   g687(.A(KEYINPUT58), .B(G1341), .Z(new_n1113));
  AOI22_X1  g688(.A1(new_n1110), .A2(new_n1111), .B1(new_n977), .B2(new_n1113), .ZN(new_n1114));
  AOI21_X1  g689(.A(new_n610), .B1(new_n1112), .B2(new_n1114), .ZN(new_n1115));
  XNOR2_X1  g690(.A(new_n1115), .B(KEYINPUT59), .ZN(new_n1116));
  NOR2_X1   g691(.A1(new_n1109), .A2(new_n1116), .ZN(new_n1117));
  INV_X1    g692(.A(KEYINPUT60), .ZN(new_n1118));
  NAND2_X1  g693(.A1(new_n1095), .A2(new_n1118), .ZN(new_n1119));
  XNOR2_X1  g694(.A(new_n600), .B(KEYINPUT122), .ZN(new_n1120));
  INV_X1    g695(.A(KEYINPUT118), .ZN(new_n1121));
  NAND2_X1  g696(.A1(new_n1094), .A2(new_n1121), .ZN(new_n1122));
  INV_X1    g697(.A(new_n1122), .ZN(new_n1123));
  NOR2_X1   g698(.A1(new_n1094), .A2(new_n1121), .ZN(new_n1124));
  OAI211_X1 g699(.A(KEYINPUT60), .B(new_n1120), .C1(new_n1123), .C2(new_n1124), .ZN(new_n1125));
  INV_X1    g700(.A(new_n1124), .ZN(new_n1126));
  AOI21_X1  g701(.A(new_n1118), .B1(new_n1126), .B2(new_n1122), .ZN(new_n1127));
  OR2_X1    g702(.A1(new_n607), .A2(KEYINPUT122), .ZN(new_n1128));
  OAI211_X1 g703(.A(new_n1119), .B(new_n1125), .C1(new_n1127), .C2(new_n1128), .ZN(new_n1129));
  AOI21_X1  g704(.A(new_n1104), .B1(new_n1117), .B2(new_n1129), .ZN(new_n1130));
  NAND2_X1  g705(.A1(new_n1073), .A2(new_n1075), .ZN(new_n1131));
  INV_X1    g706(.A(new_n1035), .ZN(new_n1132));
  XNOR2_X1  g707(.A(KEYINPUT123), .B(KEYINPUT54), .ZN(new_n1133));
  OR2_X1    g708(.A1(new_n473), .A2(KEYINPUT124), .ZN(new_n1134));
  NAND2_X1  g709(.A1(new_n473), .A2(KEYINPUT124), .ZN(new_n1135));
  AND4_X1   g710(.A1(KEYINPUT53), .A2(new_n479), .A3(G40), .A4(new_n779), .ZN(new_n1136));
  NAND4_X1  g711(.A1(new_n1078), .A2(new_n1134), .A3(new_n1135), .A4(new_n1136), .ZN(new_n1137));
  OAI211_X1 g712(.A(new_n1077), .B(new_n1137), .C1(new_n1080), .C2(KEYINPUT53), .ZN(new_n1138));
  NOR2_X1   g713(.A1(new_n1138), .A2(new_n563), .ZN(new_n1139));
  OAI21_X1  g714(.A(new_n1133), .B1(new_n1082), .B2(new_n1139), .ZN(new_n1140));
  NAND2_X1  g715(.A1(new_n1138), .A2(G171), .ZN(new_n1141));
  OAI211_X1 g716(.A(new_n1141), .B(KEYINPUT54), .C1(new_n563), .C2(new_n1081), .ZN(new_n1142));
  NAND4_X1  g717(.A1(new_n1131), .A2(new_n1132), .A3(new_n1140), .A4(new_n1142), .ZN(new_n1143));
  OAI211_X1 g718(.A(new_n1063), .B(new_n1084), .C1(new_n1130), .C2(new_n1143), .ZN(new_n1144));
  XNOR2_X1  g719(.A(G290), .B(G1986), .ZN(new_n1145));
  AOI21_X1  g720(.A(new_n969), .B1(new_n946), .B2(new_n1145), .ZN(new_n1146));
  AND3_X1   g721(.A1(new_n1144), .A2(KEYINPUT125), .A3(new_n1146), .ZN(new_n1147));
  AOI21_X1  g722(.A(KEYINPUT125), .B1(new_n1144), .B2(new_n1146), .ZN(new_n1148));
  OAI21_X1  g723(.A(new_n974), .B1(new_n1147), .B2(new_n1148), .ZN(new_n1149));
  NAND2_X1  g724(.A1(new_n1149), .A2(KEYINPUT126), .ZN(new_n1150));
  INV_X1    g725(.A(KEYINPUT126), .ZN(new_n1151));
  OAI211_X1 g726(.A(new_n1151), .B(new_n974), .C1(new_n1147), .C2(new_n1148), .ZN(new_n1152));
  NAND2_X1  g727(.A1(new_n1150), .A2(new_n1152), .ZN(G329));
  assign    G231 = 1'b0;
  NAND2_X1  g728(.A1(new_n926), .A2(new_n931), .ZN(new_n1155));
  NAND2_X1  g729(.A1(new_n933), .A2(new_n935), .ZN(new_n1156));
  NAND2_X1  g730(.A1(new_n1155), .A2(new_n1156), .ZN(new_n1157));
  NOR3_X1   g731(.A1(G229), .A2(new_n458), .A3(G227), .ZN(new_n1158));
  AND3_X1   g732(.A1(new_n870), .A2(new_n653), .A3(new_n1158), .ZN(new_n1159));
  AOI21_X1  g733(.A(KEYINPUT127), .B1(new_n1157), .B2(new_n1159), .ZN(new_n1160));
  NAND3_X1  g734(.A1(new_n870), .A2(new_n653), .A3(new_n1158), .ZN(new_n1161));
  INV_X1    g735(.A(KEYINPUT127), .ZN(new_n1162));
  NOR3_X1   g736(.A1(new_n936), .A2(new_n1161), .A3(new_n1162), .ZN(new_n1163));
  NOR2_X1   g737(.A1(new_n1160), .A2(new_n1163), .ZN(G308));
  NAND2_X1  g738(.A1(new_n1157), .A2(new_n1159), .ZN(G225));
endmodule


