//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 1 0 0 0 0 1 1 0 0 1 0 1 0 1 1 1 0 1 1 1 0 0 0 0 0 0 1 0 0 0 1 0 0 0 0 1 0 0 1 0 0 0 0 1 0 0 0 1 0 0 0 0 1 1 0 1 1 1 0 1 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:22:57 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n705, new_n706, new_n707, new_n708, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n723, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n731, new_n732, new_n733, new_n734, new_n735,
    new_n736, new_n737, new_n738, new_n739, new_n740, new_n741, new_n743,
    new_n744, new_n745, new_n746, new_n747, new_n748, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n763, new_n764, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n785, new_n786, new_n787, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n906, new_n907, new_n908, new_n909, new_n910,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n936, new_n937, new_n938, new_n939, new_n940, new_n942,
    new_n943, new_n944, new_n945, new_n946, new_n947, new_n948, new_n949,
    new_n950, new_n951, new_n953, new_n954, new_n955, new_n956, new_n957,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n988, new_n989, new_n990, new_n991, new_n992, new_n993, new_n994,
    new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004;
  INV_X1    g000(.A(G472), .ZN(new_n187));
  XNOR2_X1  g001(.A(KEYINPUT69), .B(G902), .ZN(new_n188));
  INV_X1    g002(.A(new_n188), .ZN(new_n189));
  INV_X1    g003(.A(G134), .ZN(new_n190));
  NAND2_X1  g004(.A1(new_n190), .A2(KEYINPUT65), .ZN(new_n191));
  INV_X1    g005(.A(KEYINPUT65), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n192), .A2(G134), .ZN(new_n193));
  AOI21_X1  g007(.A(G137), .B1(new_n191), .B2(new_n193), .ZN(new_n194));
  INV_X1    g008(.A(G137), .ZN(new_n195));
  NOR2_X1   g009(.A1(new_n195), .A2(G134), .ZN(new_n196));
  OAI211_X1 g010(.A(KEYINPUT66), .B(G131), .C1(new_n194), .C2(new_n196), .ZN(new_n197));
  INV_X1    g011(.A(new_n197), .ZN(new_n198));
  INV_X1    g012(.A(new_n196), .ZN(new_n199));
  XNOR2_X1  g013(.A(KEYINPUT65), .B(G134), .ZN(new_n200));
  OAI21_X1  g014(.A(new_n199), .B1(new_n200), .B2(G137), .ZN(new_n201));
  AOI21_X1  g015(.A(KEYINPUT66), .B1(new_n201), .B2(G131), .ZN(new_n202));
  NOR2_X1   g016(.A1(new_n198), .A2(new_n202), .ZN(new_n203));
  INV_X1    g017(.A(G143), .ZN(new_n204));
  OAI21_X1  g018(.A(KEYINPUT1), .B1(new_n204), .B2(G146), .ZN(new_n205));
  NOR2_X1   g019(.A1(new_n204), .A2(G146), .ZN(new_n206));
  INV_X1    g020(.A(G146), .ZN(new_n207));
  NOR2_X1   g021(.A1(new_n207), .A2(G143), .ZN(new_n208));
  OAI211_X1 g022(.A(G128), .B(new_n205), .C1(new_n206), .C2(new_n208), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n207), .A2(G143), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n204), .A2(G146), .ZN(new_n211));
  INV_X1    g025(.A(G128), .ZN(new_n212));
  OAI211_X1 g026(.A(new_n210), .B(new_n211), .C1(KEYINPUT1), .C2(new_n212), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n209), .A2(new_n213), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n191), .A2(new_n193), .ZN(new_n215));
  AOI21_X1  g029(.A(KEYINPUT11), .B1(new_n215), .B2(new_n195), .ZN(new_n216));
  NAND3_X1  g030(.A1(new_n191), .A2(new_n193), .A3(G137), .ZN(new_n217));
  NAND3_X1  g031(.A1(new_n195), .A2(KEYINPUT11), .A3(G134), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n217), .A2(new_n218), .ZN(new_n219));
  NOR2_X1   g033(.A1(new_n216), .A2(new_n219), .ZN(new_n220));
  INV_X1    g034(.A(G131), .ZN(new_n221));
  AOI21_X1  g035(.A(new_n214), .B1(new_n220), .B2(new_n221), .ZN(new_n222));
  OAI21_X1  g036(.A(G131), .B1(new_n216), .B2(new_n219), .ZN(new_n223));
  INV_X1    g037(.A(KEYINPUT11), .ZN(new_n224));
  OAI21_X1  g038(.A(new_n224), .B1(new_n200), .B2(G137), .ZN(new_n225));
  NAND2_X1  g039(.A1(KEYINPUT11), .A2(G134), .ZN(new_n226));
  NOR2_X1   g040(.A1(new_n226), .A2(G137), .ZN(new_n227));
  AOI21_X1  g041(.A(new_n227), .B1(new_n200), .B2(G137), .ZN(new_n228));
  NAND3_X1  g042(.A1(new_n225), .A2(new_n228), .A3(new_n221), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n223), .A2(new_n229), .ZN(new_n230));
  NAND2_X1  g044(.A1(KEYINPUT0), .A2(G128), .ZN(new_n231));
  NAND3_X1  g045(.A1(new_n210), .A2(new_n211), .A3(new_n231), .ZN(new_n232));
  NOR2_X1   g046(.A1(new_n206), .A2(new_n208), .ZN(new_n233));
  XOR2_X1   g047(.A(KEYINPUT0), .B(G128), .Z(new_n234));
  OAI21_X1  g048(.A(new_n232), .B1(new_n233), .B2(new_n234), .ZN(new_n235));
  AOI22_X1  g049(.A1(new_n203), .A2(new_n222), .B1(new_n230), .B2(new_n235), .ZN(new_n236));
  INV_X1    g050(.A(KEYINPUT67), .ZN(new_n237));
  INV_X1    g051(.A(G119), .ZN(new_n238));
  OAI21_X1  g052(.A(new_n237), .B1(new_n238), .B2(G116), .ZN(new_n239));
  INV_X1    g053(.A(G116), .ZN(new_n240));
  NAND3_X1  g054(.A1(new_n240), .A2(KEYINPUT67), .A3(G119), .ZN(new_n241));
  AOI22_X1  g055(.A1(new_n239), .A2(new_n241), .B1(G116), .B2(new_n238), .ZN(new_n242));
  XOR2_X1   g056(.A(KEYINPUT2), .B(G113), .Z(new_n243));
  NAND2_X1  g057(.A1(new_n242), .A2(new_n243), .ZN(new_n244));
  INV_X1    g058(.A(new_n244), .ZN(new_n245));
  NOR2_X1   g059(.A1(new_n242), .A2(new_n243), .ZN(new_n246));
  NOR2_X1   g060(.A1(new_n245), .A2(new_n246), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n236), .A2(new_n247), .ZN(new_n248));
  NOR3_X1   g062(.A1(new_n216), .A2(new_n219), .A3(G131), .ZN(new_n249));
  AOI21_X1  g063(.A(new_n221), .B1(new_n225), .B2(new_n228), .ZN(new_n250));
  OAI21_X1  g064(.A(new_n235), .B1(new_n249), .B2(new_n250), .ZN(new_n251));
  OAI21_X1  g065(.A(G131), .B1(new_n194), .B2(new_n196), .ZN(new_n252));
  INV_X1    g066(.A(KEYINPUT66), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n252), .A2(new_n253), .ZN(new_n254));
  AND2_X1   g068(.A1(new_n209), .A2(new_n213), .ZN(new_n255));
  NAND4_X1  g069(.A1(new_n254), .A2(new_n229), .A3(new_n255), .A4(new_n197), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n251), .A2(new_n256), .ZN(new_n257));
  INV_X1    g071(.A(new_n247), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n257), .A2(new_n258), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n248), .A2(new_n259), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n260), .A2(KEYINPUT28), .ZN(new_n261));
  INV_X1    g075(.A(KEYINPUT28), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n248), .A2(new_n262), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n261), .A2(new_n263), .ZN(new_n264));
  INV_X1    g078(.A(new_n264), .ZN(new_n265));
  NOR2_X1   g079(.A1(G237), .A2(G953), .ZN(new_n266));
  NAND2_X1  g080(.A1(new_n266), .A2(G210), .ZN(new_n267));
  XOR2_X1   g081(.A(new_n267), .B(KEYINPUT27), .Z(new_n268));
  XNOR2_X1  g082(.A(KEYINPUT26), .B(G101), .ZN(new_n269));
  XOR2_X1   g083(.A(new_n268), .B(new_n269), .Z(new_n270));
  INV_X1    g084(.A(new_n270), .ZN(new_n271));
  INV_X1    g085(.A(KEYINPUT29), .ZN(new_n272));
  NOR2_X1   g086(.A1(new_n271), .A2(new_n272), .ZN(new_n273));
  AOI21_X1  g087(.A(new_n189), .B1(new_n265), .B2(new_n273), .ZN(new_n274));
  XOR2_X1   g088(.A(KEYINPUT68), .B(KEYINPUT28), .Z(new_n275));
  NAND2_X1  g089(.A1(new_n260), .A2(new_n275), .ZN(new_n276));
  NAND3_X1  g090(.A1(new_n276), .A2(new_n270), .A3(new_n263), .ZN(new_n277));
  INV_X1    g091(.A(new_n248), .ZN(new_n278));
  INV_X1    g092(.A(KEYINPUT30), .ZN(new_n279));
  OAI21_X1  g093(.A(new_n279), .B1(new_n236), .B2(KEYINPUT64), .ZN(new_n280));
  INV_X1    g094(.A(KEYINPUT64), .ZN(new_n281));
  NAND3_X1  g095(.A1(new_n257), .A2(new_n281), .A3(KEYINPUT30), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n280), .A2(new_n282), .ZN(new_n283));
  AOI21_X1  g097(.A(new_n278), .B1(new_n283), .B2(new_n258), .ZN(new_n284));
  OAI211_X1 g098(.A(new_n277), .B(new_n272), .C1(new_n284), .C2(new_n270), .ZN(new_n285));
  AOI21_X1  g099(.A(new_n187), .B1(new_n274), .B2(new_n285), .ZN(new_n286));
  INV_X1    g100(.A(new_n286), .ZN(new_n287));
  INV_X1    g101(.A(KEYINPUT32), .ZN(new_n288));
  AOI21_X1  g102(.A(new_n270), .B1(new_n276), .B2(new_n263), .ZN(new_n289));
  INV_X1    g103(.A(new_n289), .ZN(new_n290));
  AOI21_X1  g104(.A(KEYINPUT31), .B1(new_n284), .B2(new_n270), .ZN(new_n291));
  AOI21_X1  g105(.A(KEYINPUT30), .B1(new_n257), .B2(new_n281), .ZN(new_n292));
  AOI211_X1 g106(.A(KEYINPUT64), .B(new_n279), .C1(new_n251), .C2(new_n256), .ZN(new_n293));
  OAI21_X1  g107(.A(new_n258), .B1(new_n292), .B2(new_n293), .ZN(new_n294));
  NAND4_X1  g108(.A1(new_n294), .A2(KEYINPUT31), .A3(new_n270), .A4(new_n248), .ZN(new_n295));
  INV_X1    g109(.A(new_n295), .ZN(new_n296));
  OAI21_X1  g110(.A(new_n290), .B1(new_n291), .B2(new_n296), .ZN(new_n297));
  NOR2_X1   g111(.A1(G472), .A2(G902), .ZN(new_n298));
  AOI21_X1  g112(.A(new_n288), .B1(new_n297), .B2(new_n298), .ZN(new_n299));
  NAND3_X1  g113(.A1(new_n294), .A2(new_n270), .A3(new_n248), .ZN(new_n300));
  INV_X1    g114(.A(KEYINPUT31), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n300), .A2(new_n301), .ZN(new_n302));
  AOI21_X1  g116(.A(new_n289), .B1(new_n302), .B2(new_n295), .ZN(new_n303));
  INV_X1    g117(.A(new_n298), .ZN(new_n304));
  NOR3_X1   g118(.A1(new_n303), .A2(KEYINPUT32), .A3(new_n304), .ZN(new_n305));
  OAI21_X1  g119(.A(new_n287), .B1(new_n299), .B2(new_n305), .ZN(new_n306));
  INV_X1    g120(.A(G478), .ZN(new_n307));
  NOR2_X1   g121(.A1(KEYINPUT91), .A2(KEYINPUT15), .ZN(new_n308));
  INV_X1    g122(.A(new_n308), .ZN(new_n309));
  NAND2_X1  g123(.A1(KEYINPUT91), .A2(KEYINPUT15), .ZN(new_n310));
  AOI21_X1  g124(.A(new_n307), .B1(new_n309), .B2(new_n310), .ZN(new_n311));
  INV_X1    g125(.A(new_n311), .ZN(new_n312));
  INV_X1    g126(.A(KEYINPUT88), .ZN(new_n313));
  OAI21_X1  g127(.A(new_n313), .B1(new_n204), .B2(G128), .ZN(new_n314));
  NAND3_X1  g128(.A1(new_n212), .A2(KEYINPUT88), .A3(G143), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n314), .A2(new_n315), .ZN(new_n316));
  INV_X1    g130(.A(KEYINPUT87), .ZN(new_n317));
  OAI21_X1  g131(.A(new_n317), .B1(new_n212), .B2(G143), .ZN(new_n318));
  NAND3_X1  g132(.A1(new_n204), .A2(KEYINPUT87), .A3(G128), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n318), .A2(new_n319), .ZN(new_n320));
  INV_X1    g134(.A(KEYINPUT13), .ZN(new_n321));
  OAI21_X1  g135(.A(new_n316), .B1(new_n320), .B2(new_n321), .ZN(new_n322));
  AOI21_X1  g136(.A(KEYINPUT13), .B1(new_n318), .B2(new_n319), .ZN(new_n323));
  OAI21_X1  g137(.A(G134), .B1(new_n322), .B2(new_n323), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n324), .A2(KEYINPUT89), .ZN(new_n325));
  INV_X1    g139(.A(KEYINPUT89), .ZN(new_n326));
  OAI211_X1 g140(.A(new_n326), .B(G134), .C1(new_n322), .C2(new_n323), .ZN(new_n327));
  NAND3_X1  g141(.A1(new_n320), .A2(new_n316), .A3(new_n200), .ZN(new_n328));
  INV_X1    g142(.A(new_n328), .ZN(new_n329));
  XNOR2_X1  g143(.A(G116), .B(G122), .ZN(new_n330));
  XNOR2_X1  g144(.A(new_n330), .B(G107), .ZN(new_n331));
  NOR2_X1   g145(.A1(new_n329), .A2(new_n331), .ZN(new_n332));
  NAND3_X1  g146(.A1(new_n325), .A2(new_n327), .A3(new_n332), .ZN(new_n333));
  INV_X1    g147(.A(G107), .ZN(new_n334));
  INV_X1    g148(.A(G122), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n335), .A2(G116), .ZN(new_n336));
  AOI21_X1  g150(.A(new_n334), .B1(new_n336), .B2(KEYINPUT14), .ZN(new_n337));
  XNOR2_X1  g151(.A(new_n337), .B(new_n330), .ZN(new_n338));
  AOI21_X1  g152(.A(new_n200), .B1(new_n320), .B2(new_n316), .ZN(new_n339));
  OAI21_X1  g153(.A(new_n338), .B1(new_n329), .B2(new_n339), .ZN(new_n340));
  INV_X1    g154(.A(KEYINPUT90), .ZN(new_n341));
  NOR2_X1   g155(.A1(new_n340), .A2(new_n341), .ZN(new_n342));
  INV_X1    g156(.A(new_n339), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n343), .A2(new_n328), .ZN(new_n344));
  AOI21_X1  g158(.A(KEYINPUT90), .B1(new_n344), .B2(new_n338), .ZN(new_n345));
  OAI21_X1  g159(.A(new_n333), .B1(new_n342), .B2(new_n345), .ZN(new_n346));
  XNOR2_X1  g160(.A(KEYINPUT9), .B(G234), .ZN(new_n347));
  INV_X1    g161(.A(G217), .ZN(new_n348));
  NOR3_X1   g162(.A1(new_n347), .A2(new_n348), .A3(G953), .ZN(new_n349));
  INV_X1    g163(.A(new_n349), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n346), .A2(new_n350), .ZN(new_n351));
  OAI211_X1 g165(.A(new_n333), .B(new_n349), .C1(new_n342), .C2(new_n345), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n351), .A2(new_n352), .ZN(new_n353));
  AOI21_X1  g167(.A(new_n312), .B1(new_n353), .B2(new_n188), .ZN(new_n354));
  AOI211_X1 g168(.A(new_n189), .B(new_n311), .C1(new_n351), .C2(new_n352), .ZN(new_n355));
  NOR2_X1   g169(.A1(new_n354), .A2(new_n355), .ZN(new_n356));
  NOR2_X1   g170(.A1(G475), .A2(G902), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n266), .A2(G214), .ZN(new_n358));
  NAND2_X1  g172(.A1(new_n358), .A2(new_n204), .ZN(new_n359));
  INV_X1    g173(.A(G237), .ZN(new_n360));
  INV_X1    g174(.A(G953), .ZN(new_n361));
  NAND4_X1  g175(.A1(new_n360), .A2(new_n361), .A3(G143), .A4(G214), .ZN(new_n362));
  AND2_X1   g176(.A1(new_n362), .A2(KEYINPUT83), .ZN(new_n363));
  INV_X1    g177(.A(KEYINPUT83), .ZN(new_n364));
  NAND4_X1  g178(.A1(new_n266), .A2(new_n364), .A3(G143), .A4(G214), .ZN(new_n365));
  INV_X1    g179(.A(new_n365), .ZN(new_n366));
  OAI211_X1 g180(.A(new_n221), .B(new_n359), .C1(new_n363), .C2(new_n366), .ZN(new_n367));
  INV_X1    g181(.A(KEYINPUT85), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n367), .A2(new_n368), .ZN(new_n369));
  OAI21_X1  g183(.A(new_n359), .B1(new_n363), .B2(new_n366), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n370), .A2(G131), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n362), .A2(KEYINPUT83), .ZN(new_n372));
  AOI22_X1  g186(.A1(new_n372), .A2(new_n365), .B1(new_n204), .B2(new_n358), .ZN(new_n373));
  NAND3_X1  g187(.A1(new_n373), .A2(KEYINPUT85), .A3(new_n221), .ZN(new_n374));
  INV_X1    g188(.A(KEYINPUT17), .ZN(new_n375));
  NAND4_X1  g189(.A1(new_n369), .A2(new_n371), .A3(new_n374), .A4(new_n375), .ZN(new_n376));
  NOR3_X1   g190(.A1(new_n373), .A2(new_n375), .A3(new_n221), .ZN(new_n377));
  INV_X1    g191(.A(G140), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n378), .A2(G125), .ZN(new_n379));
  INV_X1    g193(.A(G125), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n380), .A2(G140), .ZN(new_n381));
  NAND3_X1  g195(.A1(new_n379), .A2(new_n381), .A3(KEYINPUT16), .ZN(new_n382));
  OR3_X1    g196(.A1(new_n380), .A2(KEYINPUT16), .A3(G140), .ZN(new_n383));
  NAND3_X1  g197(.A1(new_n382), .A2(new_n383), .A3(G146), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n384), .A2(KEYINPUT70), .ZN(new_n385));
  INV_X1    g199(.A(KEYINPUT70), .ZN(new_n386));
  NAND4_X1  g200(.A1(new_n382), .A2(new_n383), .A3(new_n386), .A4(G146), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n382), .A2(new_n383), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n388), .A2(new_n207), .ZN(new_n389));
  NAND3_X1  g203(.A1(new_n385), .A2(new_n387), .A3(new_n389), .ZN(new_n390));
  NOR2_X1   g204(.A1(new_n377), .A2(new_n390), .ZN(new_n391));
  NAND2_X1  g205(.A1(new_n376), .A2(new_n391), .ZN(new_n392));
  XNOR2_X1  g206(.A(G113), .B(G122), .ZN(new_n393));
  INV_X1    g207(.A(G104), .ZN(new_n394));
  XNOR2_X1  g208(.A(new_n393), .B(new_n394), .ZN(new_n395));
  INV_X1    g209(.A(KEYINPUT18), .ZN(new_n396));
  NOR2_X1   g210(.A1(new_n396), .A2(new_n221), .ZN(new_n397));
  INV_X1    g211(.A(new_n397), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n373), .A2(new_n398), .ZN(new_n399));
  AND2_X1   g213(.A1(new_n379), .A2(new_n381), .ZN(new_n400));
  XNOR2_X1  g214(.A(new_n400), .B(new_n207), .ZN(new_n401));
  INV_X1    g215(.A(KEYINPUT84), .ZN(new_n402));
  AOI21_X1  g216(.A(new_n402), .B1(new_n370), .B2(new_n397), .ZN(new_n403));
  NOR3_X1   g217(.A1(new_n373), .A2(KEYINPUT84), .A3(new_n398), .ZN(new_n404));
  OAI211_X1 g218(.A(new_n399), .B(new_n401), .C1(new_n403), .C2(new_n404), .ZN(new_n405));
  AND3_X1   g219(.A1(new_n392), .A2(new_n395), .A3(new_n405), .ZN(new_n406));
  NAND3_X1  g220(.A1(new_n369), .A2(new_n374), .A3(new_n371), .ZN(new_n407));
  INV_X1    g221(.A(new_n384), .ZN(new_n408));
  XNOR2_X1  g222(.A(new_n400), .B(KEYINPUT19), .ZN(new_n409));
  AOI21_X1  g223(.A(new_n408), .B1(new_n409), .B2(new_n207), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n407), .A2(new_n410), .ZN(new_n411));
  AOI21_X1  g225(.A(new_n395), .B1(new_n411), .B2(new_n405), .ZN(new_n412));
  OAI21_X1  g226(.A(new_n357), .B1(new_n406), .B2(new_n412), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n413), .A2(KEYINPUT20), .ZN(new_n414));
  INV_X1    g228(.A(new_n412), .ZN(new_n415));
  NAND3_X1  g229(.A1(new_n392), .A2(new_n395), .A3(new_n405), .ZN(new_n416));
  NAND2_X1  g230(.A1(new_n415), .A2(new_n416), .ZN(new_n417));
  INV_X1    g231(.A(KEYINPUT20), .ZN(new_n418));
  NAND3_X1  g232(.A1(new_n417), .A2(new_n418), .A3(new_n357), .ZN(new_n419));
  NAND2_X1  g233(.A1(new_n414), .A2(new_n419), .ZN(new_n420));
  AND2_X1   g234(.A1(new_n356), .A2(new_n420), .ZN(new_n421));
  INV_X1    g235(.A(G902), .ZN(new_n422));
  AOI21_X1  g236(.A(new_n395), .B1(new_n392), .B2(new_n405), .ZN(new_n423));
  OAI21_X1  g237(.A(new_n422), .B1(new_n406), .B2(new_n423), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n424), .A2(KEYINPUT86), .ZN(new_n425));
  INV_X1    g239(.A(KEYINPUT86), .ZN(new_n426));
  OAI211_X1 g240(.A(new_n426), .B(new_n422), .C1(new_n406), .C2(new_n423), .ZN(new_n427));
  NAND3_X1  g241(.A1(new_n425), .A2(G475), .A3(new_n427), .ZN(new_n428));
  INV_X1    g242(.A(G952), .ZN(new_n429));
  AOI211_X1 g243(.A(G953), .B(new_n429), .C1(G234), .C2(G237), .ZN(new_n430));
  AOI211_X1 g244(.A(new_n361), .B(new_n188), .C1(G234), .C2(G237), .ZN(new_n431));
  XNOR2_X1  g245(.A(KEYINPUT21), .B(G898), .ZN(new_n432));
  AOI21_X1  g246(.A(new_n430), .B1(new_n431), .B2(new_n432), .ZN(new_n433));
  INV_X1    g247(.A(new_n433), .ZN(new_n434));
  NAND3_X1  g248(.A1(new_n421), .A2(new_n428), .A3(new_n434), .ZN(new_n435));
  XNOR2_X1  g249(.A(G110), .B(G140), .ZN(new_n436));
  INV_X1    g250(.A(G227), .ZN(new_n437));
  NOR2_X1   g251(.A1(new_n437), .A2(G953), .ZN(new_n438));
  XOR2_X1   g252(.A(new_n436), .B(new_n438), .Z(new_n439));
  INV_X1    g253(.A(new_n439), .ZN(new_n440));
  INV_X1    g254(.A(KEYINPUT10), .ZN(new_n441));
  NOR2_X1   g255(.A1(new_n334), .A2(G104), .ZN(new_n442));
  INV_X1    g256(.A(new_n442), .ZN(new_n443));
  INV_X1    g257(.A(G101), .ZN(new_n444));
  AND3_X1   g258(.A1(new_n334), .A2(KEYINPUT3), .A3(G104), .ZN(new_n445));
  AOI21_X1  g259(.A(KEYINPUT3), .B1(new_n334), .B2(G104), .ZN(new_n446));
  OAI211_X1 g260(.A(new_n443), .B(new_n444), .C1(new_n445), .C2(new_n446), .ZN(new_n447));
  INV_X1    g261(.A(KEYINPUT74), .ZN(new_n448));
  OAI21_X1  g262(.A(new_n448), .B1(new_n334), .B2(G104), .ZN(new_n449));
  NAND3_X1  g263(.A1(new_n394), .A2(KEYINPUT74), .A3(G107), .ZN(new_n450));
  AOI22_X1  g264(.A1(new_n449), .A2(new_n450), .B1(G104), .B2(new_n334), .ZN(new_n451));
  OAI21_X1  g265(.A(new_n447), .B1(new_n444), .B2(new_n451), .ZN(new_n452));
  OAI21_X1  g266(.A(new_n441), .B1(new_n452), .B2(new_n214), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n334), .A2(G104), .ZN(new_n454));
  AND3_X1   g268(.A1(new_n394), .A2(KEYINPUT74), .A3(G107), .ZN(new_n455));
  AOI21_X1  g269(.A(KEYINPUT74), .B1(new_n394), .B2(G107), .ZN(new_n456));
  OAI21_X1  g270(.A(new_n454), .B1(new_n455), .B2(new_n456), .ZN(new_n457));
  NAND2_X1  g271(.A1(new_n457), .A2(G101), .ZN(new_n458));
  NAND4_X1  g272(.A1(new_n255), .A2(KEYINPUT10), .A3(new_n447), .A4(new_n458), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n453), .A2(new_n459), .ZN(new_n460));
  OAI21_X1  g274(.A(new_n443), .B1(new_n445), .B2(new_n446), .ZN(new_n461));
  NAND3_X1  g275(.A1(new_n461), .A2(KEYINPUT72), .A3(G101), .ZN(new_n462));
  INV_X1    g276(.A(KEYINPUT72), .ZN(new_n463));
  INV_X1    g277(.A(KEYINPUT3), .ZN(new_n464));
  OAI21_X1  g278(.A(new_n464), .B1(new_n394), .B2(G107), .ZN(new_n465));
  NAND3_X1  g279(.A1(new_n334), .A2(KEYINPUT3), .A3(G104), .ZN(new_n466));
  AOI21_X1  g280(.A(new_n442), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  OAI21_X1  g281(.A(new_n463), .B1(new_n467), .B2(new_n444), .ZN(new_n468));
  INV_X1    g282(.A(KEYINPUT4), .ZN(new_n469));
  AOI21_X1  g283(.A(new_n469), .B1(new_n467), .B2(new_n444), .ZN(new_n470));
  NAND3_X1  g284(.A1(new_n462), .A2(new_n468), .A3(new_n470), .ZN(new_n471));
  INV_X1    g285(.A(KEYINPUT73), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n471), .A2(new_n472), .ZN(new_n473));
  NAND4_X1  g287(.A1(new_n462), .A2(new_n468), .A3(new_n470), .A4(KEYINPUT73), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n473), .A2(new_n474), .ZN(new_n475));
  NOR3_X1   g289(.A1(new_n467), .A2(KEYINPUT4), .A3(new_n444), .ZN(new_n476));
  INV_X1    g290(.A(new_n476), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n477), .A2(new_n235), .ZN(new_n478));
  INV_X1    g292(.A(new_n478), .ZN(new_n479));
  AOI21_X1  g293(.A(new_n460), .B1(new_n475), .B2(new_n479), .ZN(new_n480));
  INV_X1    g294(.A(new_n230), .ZN(new_n481));
  AOI21_X1  g295(.A(new_n440), .B1(new_n480), .B2(new_n481), .ZN(new_n482));
  AOI21_X1  g296(.A(new_n478), .B1(new_n473), .B2(new_n474), .ZN(new_n483));
  OAI21_X1  g297(.A(new_n230), .B1(new_n483), .B2(new_n460), .ZN(new_n484));
  NAND2_X1  g298(.A1(new_n482), .A2(new_n484), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n475), .A2(new_n479), .ZN(new_n486));
  NAND4_X1  g300(.A1(new_n486), .A2(new_n481), .A3(new_n453), .A4(new_n459), .ZN(new_n487));
  XNOR2_X1  g301(.A(KEYINPUT75), .B(KEYINPUT12), .ZN(new_n488));
  NOR2_X1   g302(.A1(new_n452), .A2(new_n214), .ZN(new_n489));
  AOI22_X1  g303(.A1(new_n458), .A2(new_n447), .B1(new_n213), .B2(new_n209), .ZN(new_n490));
  OAI211_X1 g304(.A(new_n230), .B(new_n488), .C1(new_n489), .C2(new_n490), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n491), .A2(KEYINPUT76), .ZN(new_n492));
  NAND3_X1  g306(.A1(new_n255), .A2(new_n447), .A3(new_n458), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n452), .A2(new_n214), .ZN(new_n494));
  NAND2_X1  g308(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  INV_X1    g309(.A(KEYINPUT76), .ZN(new_n496));
  NAND4_X1  g310(.A1(new_n495), .A2(new_n496), .A3(new_n230), .A4(new_n488), .ZN(new_n497));
  OAI21_X1  g311(.A(new_n230), .B1(new_n489), .B2(new_n490), .ZN(new_n498));
  INV_X1    g312(.A(KEYINPUT12), .ZN(new_n499));
  NAND2_X1  g313(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  NAND3_X1  g314(.A1(new_n492), .A2(new_n497), .A3(new_n500), .ZN(new_n501));
  NAND3_X1  g315(.A1(new_n487), .A2(new_n501), .A3(KEYINPUT77), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n502), .A2(new_n440), .ZN(new_n503));
  AOI21_X1  g317(.A(KEYINPUT77), .B1(new_n487), .B2(new_n501), .ZN(new_n504));
  OAI211_X1 g318(.A(G469), .B(new_n485), .C1(new_n503), .C2(new_n504), .ZN(new_n505));
  INV_X1    g319(.A(G469), .ZN(new_n506));
  AND2_X1   g320(.A1(new_n482), .A2(new_n501), .ZN(new_n507));
  AOI21_X1  g321(.A(new_n439), .B1(new_n487), .B2(new_n484), .ZN(new_n508));
  OAI211_X1 g322(.A(new_n506), .B(new_n188), .C1(new_n507), .C2(new_n508), .ZN(new_n509));
  NOR2_X1   g323(.A1(new_n506), .A2(new_n422), .ZN(new_n510));
  INV_X1    g324(.A(new_n510), .ZN(new_n511));
  NAND3_X1  g325(.A1(new_n505), .A2(new_n509), .A3(new_n511), .ZN(new_n512));
  INV_X1    g326(.A(G221), .ZN(new_n513));
  INV_X1    g327(.A(new_n347), .ZN(new_n514));
  AOI21_X1  g328(.A(new_n513), .B1(new_n514), .B2(new_n422), .ZN(new_n515));
  INV_X1    g329(.A(new_n515), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n512), .A2(new_n516), .ZN(new_n517));
  NOR2_X1   g331(.A1(new_n435), .A2(new_n517), .ZN(new_n518));
  XNOR2_X1  g332(.A(KEYINPUT22), .B(G137), .ZN(new_n519));
  AND3_X1   g333(.A1(new_n361), .A2(G221), .A3(G234), .ZN(new_n520));
  XNOR2_X1  g334(.A(new_n519), .B(new_n520), .ZN(new_n521));
  INV_X1    g335(.A(KEYINPUT23), .ZN(new_n522));
  OAI21_X1  g336(.A(new_n522), .B1(new_n238), .B2(G128), .ZN(new_n523));
  NAND3_X1  g337(.A1(new_n212), .A2(KEYINPUT23), .A3(G119), .ZN(new_n524));
  OAI211_X1 g338(.A(new_n523), .B(new_n524), .C1(G119), .C2(new_n212), .ZN(new_n525));
  XNOR2_X1  g339(.A(G119), .B(G128), .ZN(new_n526));
  XOR2_X1   g340(.A(KEYINPUT24), .B(G110), .Z(new_n527));
  AOI22_X1  g341(.A1(new_n525), .A2(G110), .B1(new_n526), .B2(new_n527), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n390), .A2(new_n528), .ZN(new_n529));
  OAI22_X1  g343(.A1(new_n525), .A2(G110), .B1(new_n526), .B2(new_n527), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n400), .A2(new_n207), .ZN(new_n531));
  NAND3_X1  g345(.A1(new_n530), .A2(new_n384), .A3(new_n531), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n529), .A2(new_n532), .ZN(new_n533));
  INV_X1    g347(.A(KEYINPUT71), .ZN(new_n534));
  AOI21_X1  g348(.A(new_n521), .B1(new_n533), .B2(new_n534), .ZN(new_n535));
  NAND3_X1  g349(.A1(new_n529), .A2(KEYINPUT71), .A3(new_n532), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  NAND4_X1  g351(.A1(new_n529), .A2(KEYINPUT71), .A3(new_n521), .A4(new_n532), .ZN(new_n538));
  AOI21_X1  g352(.A(new_n189), .B1(new_n537), .B2(new_n538), .ZN(new_n539));
  INV_X1    g353(.A(KEYINPUT25), .ZN(new_n540));
  OR2_X1    g354(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  AOI21_X1  g355(.A(new_n348), .B1(new_n188), .B2(G234), .ZN(new_n542));
  INV_X1    g356(.A(new_n542), .ZN(new_n543));
  AOI21_X1  g357(.A(new_n543), .B1(new_n539), .B2(new_n540), .ZN(new_n544));
  NAND2_X1  g358(.A1(new_n541), .A2(new_n544), .ZN(new_n545));
  NAND2_X1  g359(.A1(new_n537), .A2(new_n538), .ZN(new_n546));
  NOR2_X1   g360(.A1(new_n542), .A2(G902), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n546), .A2(new_n547), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n545), .A2(new_n548), .ZN(new_n549));
  INV_X1    g363(.A(new_n549), .ZN(new_n550));
  OAI21_X1  g364(.A(G214), .B1(G237), .B2(G902), .ZN(new_n551));
  INV_X1    g365(.A(new_n551), .ZN(new_n552));
  OAI21_X1  g366(.A(G210), .B1(G237), .B2(G902), .ZN(new_n553));
  INV_X1    g367(.A(new_n553), .ZN(new_n554));
  OAI21_X1  g368(.A(new_n477), .B1(new_n245), .B2(new_n246), .ZN(new_n555));
  INV_X1    g369(.A(new_n555), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n475), .A2(new_n556), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n238), .A2(G116), .ZN(new_n558));
  OAI21_X1  g372(.A(G113), .B1(new_n558), .B2(KEYINPUT5), .ZN(new_n559));
  AOI21_X1  g373(.A(new_n559), .B1(new_n242), .B2(KEYINPUT5), .ZN(new_n560));
  NOR3_X1   g374(.A1(new_n452), .A2(new_n245), .A3(new_n560), .ZN(new_n561));
  INV_X1    g375(.A(new_n561), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n557), .A2(new_n562), .ZN(new_n563));
  INV_X1    g377(.A(KEYINPUT6), .ZN(new_n564));
  XNOR2_X1  g378(.A(G110), .B(G122), .ZN(new_n565));
  INV_X1    g379(.A(new_n565), .ZN(new_n566));
  NAND4_X1  g380(.A1(new_n563), .A2(KEYINPUT78), .A3(new_n564), .A4(new_n566), .ZN(new_n567));
  AOI21_X1  g381(.A(new_n555), .B1(new_n473), .B2(new_n474), .ZN(new_n568));
  OAI211_X1 g382(.A(new_n564), .B(new_n566), .C1(new_n568), .C2(new_n561), .ZN(new_n569));
  INV_X1    g383(.A(KEYINPUT78), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n569), .A2(new_n570), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n567), .A2(new_n571), .ZN(new_n572));
  AOI21_X1  g386(.A(G125), .B1(new_n209), .B2(new_n213), .ZN(new_n573));
  INV_X1    g387(.A(KEYINPUT79), .ZN(new_n574));
  OAI211_X1 g388(.A(G125), .B(new_n232), .C1(new_n233), .C2(new_n234), .ZN(new_n575));
  AOI21_X1  g389(.A(new_n573), .B1(new_n574), .B2(new_n575), .ZN(new_n576));
  INV_X1    g390(.A(new_n575), .ZN(new_n577));
  NAND2_X1  g391(.A1(new_n577), .A2(KEYINPUT79), .ZN(new_n578));
  NAND2_X1  g392(.A1(new_n576), .A2(new_n578), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n361), .A2(G224), .ZN(new_n580));
  XOR2_X1   g394(.A(new_n579), .B(new_n580), .Z(new_n581));
  NOR3_X1   g395(.A1(new_n568), .A2(new_n561), .A3(new_n566), .ZN(new_n582));
  INV_X1    g396(.A(new_n582), .ZN(new_n583));
  OAI21_X1  g397(.A(new_n566), .B1(new_n568), .B2(new_n561), .ZN(new_n584));
  NAND3_X1  g398(.A1(new_n583), .A2(KEYINPUT6), .A3(new_n584), .ZN(new_n585));
  AND3_X1   g399(.A1(new_n572), .A2(new_n581), .A3(new_n585), .ZN(new_n586));
  AND2_X1   g400(.A1(KEYINPUT80), .A2(KEYINPUT7), .ZN(new_n587));
  NOR2_X1   g401(.A1(KEYINPUT80), .A2(KEYINPUT7), .ZN(new_n588));
  OAI21_X1  g402(.A(new_n580), .B1(new_n587), .B2(new_n588), .ZN(new_n589));
  OAI21_X1  g403(.A(new_n589), .B1(new_n577), .B2(new_n573), .ZN(new_n590));
  NAND2_X1  g404(.A1(new_n590), .A2(KEYINPUT81), .ZN(new_n591));
  INV_X1    g405(.A(KEYINPUT81), .ZN(new_n592));
  OAI211_X1 g406(.A(new_n592), .B(new_n589), .C1(new_n577), .C2(new_n573), .ZN(new_n593));
  NAND2_X1  g407(.A1(new_n591), .A2(new_n593), .ZN(new_n594));
  XNOR2_X1  g408(.A(new_n565), .B(KEYINPUT8), .ZN(new_n595));
  INV_X1    g409(.A(new_n560), .ZN(new_n596));
  AOI22_X1  g410(.A1(new_n596), .A2(new_n244), .B1(new_n447), .B2(new_n458), .ZN(new_n597));
  OAI21_X1  g411(.A(new_n595), .B1(new_n597), .B2(new_n561), .ZN(new_n598));
  NAND4_X1  g412(.A1(new_n576), .A2(new_n578), .A3(KEYINPUT7), .A4(new_n580), .ZN(new_n599));
  NAND3_X1  g413(.A1(new_n594), .A2(new_n598), .A3(new_n599), .ZN(new_n600));
  OAI21_X1  g414(.A(new_n422), .B1(new_n582), .B2(new_n600), .ZN(new_n601));
  INV_X1    g415(.A(KEYINPUT82), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n601), .A2(new_n602), .ZN(new_n603));
  OAI211_X1 g417(.A(KEYINPUT82), .B(new_n422), .C1(new_n582), .C2(new_n600), .ZN(new_n604));
  NAND2_X1  g418(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  OAI21_X1  g419(.A(new_n554), .B1(new_n586), .B2(new_n605), .ZN(new_n606));
  NAND3_X1  g420(.A1(new_n572), .A2(new_n581), .A3(new_n585), .ZN(new_n607));
  NAND4_X1  g421(.A1(new_n607), .A2(new_n553), .A3(new_n603), .A4(new_n604), .ZN(new_n608));
  AOI21_X1  g422(.A(new_n552), .B1(new_n606), .B2(new_n608), .ZN(new_n609));
  NAND4_X1  g423(.A1(new_n306), .A2(new_n518), .A3(new_n550), .A4(new_n609), .ZN(new_n610));
  XNOR2_X1  g424(.A(new_n610), .B(G101), .ZN(G3));
  NAND2_X1  g425(.A1(new_n609), .A2(new_n434), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n428), .A2(new_n420), .ZN(new_n613));
  INV_X1    g427(.A(KEYINPUT33), .ZN(new_n614));
  OR2_X1    g428(.A1(new_n614), .A2(KEYINPUT92), .ZN(new_n615));
  NAND2_X1  g429(.A1(new_n614), .A2(KEYINPUT92), .ZN(new_n616));
  INV_X1    g430(.A(new_n352), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n340), .A2(new_n341), .ZN(new_n618));
  NAND3_X1  g432(.A1(new_n344), .A2(KEYINPUT90), .A3(new_n338), .ZN(new_n619));
  NAND2_X1  g433(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  AOI21_X1  g434(.A(new_n349), .B1(new_n620), .B2(new_n333), .ZN(new_n621));
  OAI211_X1 g435(.A(new_n615), .B(new_n616), .C1(new_n617), .C2(new_n621), .ZN(new_n622));
  NAND4_X1  g436(.A1(new_n351), .A2(KEYINPUT92), .A3(new_n614), .A4(new_n352), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  NOR2_X1   g438(.A1(new_n189), .A2(new_n307), .ZN(new_n625));
  NAND2_X1  g439(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  AOI21_X1  g440(.A(G478), .B1(new_n353), .B2(new_n188), .ZN(new_n627));
  INV_X1    g441(.A(new_n627), .ZN(new_n628));
  NAND2_X1  g442(.A1(new_n626), .A2(new_n628), .ZN(new_n629));
  NAND2_X1  g443(.A1(new_n613), .A2(new_n629), .ZN(new_n630));
  NOR2_X1   g444(.A1(new_n612), .A2(new_n630), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n297), .A2(new_n188), .ZN(new_n632));
  AOI22_X1  g446(.A1(new_n632), .A2(G472), .B1(new_n298), .B2(new_n297), .ZN(new_n633));
  NOR2_X1   g447(.A1(new_n517), .A2(new_n549), .ZN(new_n634));
  NAND3_X1  g448(.A1(new_n631), .A2(new_n633), .A3(new_n634), .ZN(new_n635));
  XOR2_X1   g449(.A(KEYINPUT34), .B(G104), .Z(new_n636));
  XNOR2_X1  g450(.A(new_n635), .B(new_n636), .ZN(G6));
  NAND2_X1  g451(.A1(new_n428), .A2(KEYINPUT93), .ZN(new_n638));
  INV_X1    g452(.A(G475), .ZN(new_n639));
  AOI21_X1  g453(.A(new_n639), .B1(new_n424), .B2(KEYINPUT86), .ZN(new_n640));
  INV_X1    g454(.A(KEYINPUT93), .ZN(new_n641));
  NAND3_X1  g455(.A1(new_n640), .A2(new_n641), .A3(new_n427), .ZN(new_n642));
  NAND2_X1  g456(.A1(new_n638), .A2(new_n642), .ZN(new_n643));
  INV_X1    g457(.A(new_n643), .ZN(new_n644));
  NOR2_X1   g458(.A1(new_n617), .A2(new_n621), .ZN(new_n645));
  OAI21_X1  g459(.A(new_n311), .B1(new_n645), .B2(new_n189), .ZN(new_n646));
  NAND3_X1  g460(.A1(new_n353), .A2(new_n188), .A3(new_n312), .ZN(new_n647));
  NAND2_X1  g461(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  AND2_X1   g462(.A1(new_n648), .A2(new_n420), .ZN(new_n649));
  AND4_X1   g463(.A1(new_n609), .A2(new_n434), .A3(new_n644), .A4(new_n649), .ZN(new_n650));
  NAND3_X1  g464(.A1(new_n650), .A2(new_n633), .A3(new_n634), .ZN(new_n651));
  XOR2_X1   g465(.A(KEYINPUT35), .B(G107), .Z(new_n652));
  XNOR2_X1  g466(.A(new_n651), .B(new_n652), .ZN(G9));
  NOR2_X1   g467(.A1(new_n521), .A2(KEYINPUT36), .ZN(new_n654));
  XNOR2_X1  g468(.A(new_n533), .B(new_n654), .ZN(new_n655));
  NAND2_X1  g469(.A1(new_n655), .A2(new_n547), .ZN(new_n656));
  INV_X1    g470(.A(new_n656), .ZN(new_n657));
  AOI21_X1  g471(.A(new_n657), .B1(new_n541), .B2(new_n544), .ZN(new_n658));
  INV_X1    g472(.A(new_n658), .ZN(new_n659));
  NAND4_X1  g473(.A1(new_n518), .A2(new_n633), .A3(new_n609), .A4(new_n659), .ZN(new_n660));
  XNOR2_X1  g474(.A(new_n660), .B(KEYINPUT94), .ZN(new_n661));
  XNOR2_X1  g475(.A(KEYINPUT37), .B(G110), .ZN(new_n662));
  XNOR2_X1  g476(.A(new_n661), .B(new_n662), .ZN(G12));
  AOI211_X1 g477(.A(new_n552), .B(new_n658), .C1(new_n606), .C2(new_n608), .ZN(new_n664));
  INV_X1    g478(.A(new_n517), .ZN(new_n665));
  INV_X1    g479(.A(G900), .ZN(new_n666));
  AOI21_X1  g480(.A(new_n430), .B1(new_n431), .B2(new_n666), .ZN(new_n667));
  INV_X1    g481(.A(new_n667), .ZN(new_n668));
  AND4_X1   g482(.A1(new_n638), .A2(new_n649), .A3(new_n642), .A4(new_n668), .ZN(new_n669));
  NAND4_X1  g483(.A1(new_n306), .A2(new_n664), .A3(new_n665), .A4(new_n669), .ZN(new_n670));
  INV_X1    g484(.A(KEYINPUT95), .ZN(new_n671));
  NAND2_X1  g485(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  NAND3_X1  g486(.A1(new_n297), .A2(new_n288), .A3(new_n298), .ZN(new_n673));
  OAI21_X1  g487(.A(KEYINPUT32), .B1(new_n303), .B2(new_n304), .ZN(new_n674));
  NAND2_X1  g488(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  AOI21_X1  g489(.A(new_n517), .B1(new_n675), .B2(new_n287), .ZN(new_n676));
  NAND4_X1  g490(.A1(new_n676), .A2(KEYINPUT95), .A3(new_n669), .A4(new_n664), .ZN(new_n677));
  NAND2_X1  g491(.A1(new_n672), .A2(new_n677), .ZN(new_n678));
  XNOR2_X1  g492(.A(new_n678), .B(G128), .ZN(G30));
  XOR2_X1   g493(.A(new_n667), .B(KEYINPUT39), .Z(new_n680));
  NAND2_X1  g494(.A1(new_n665), .A2(new_n680), .ZN(new_n681));
  XOR2_X1   g495(.A(new_n681), .B(KEYINPUT100), .Z(new_n682));
  NAND2_X1  g496(.A1(new_n682), .A2(KEYINPUT40), .ZN(new_n683));
  XNOR2_X1  g497(.A(new_n681), .B(KEYINPUT100), .ZN(new_n684));
  INV_X1    g498(.A(KEYINPUT40), .ZN(new_n685));
  NAND2_X1  g499(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  NAND2_X1  g500(.A1(new_n606), .A2(new_n608), .ZN(new_n687));
  XOR2_X1   g501(.A(KEYINPUT97), .B(KEYINPUT38), .Z(new_n688));
  XNOR2_X1  g502(.A(new_n688), .B(KEYINPUT96), .ZN(new_n689));
  XOR2_X1   g503(.A(new_n687), .B(new_n689), .Z(new_n690));
  AOI22_X1  g504(.A1(new_n640), .A2(new_n427), .B1(new_n414), .B2(new_n419), .ZN(new_n691));
  NOR4_X1   g505(.A1(new_n659), .A2(new_n691), .A3(new_n552), .A4(new_n356), .ZN(new_n692));
  AND2_X1   g506(.A1(new_n692), .A2(KEYINPUT99), .ZN(new_n693));
  INV_X1    g507(.A(new_n675), .ZN(new_n694));
  NAND2_X1  g508(.A1(new_n260), .A2(new_n271), .ZN(new_n695));
  XNOR2_X1  g509(.A(new_n695), .B(KEYINPUT98), .ZN(new_n696));
  INV_X1    g510(.A(new_n300), .ZN(new_n697));
  OAI21_X1  g511(.A(new_n422), .B1(new_n696), .B2(new_n697), .ZN(new_n698));
  AND2_X1   g512(.A1(new_n698), .A2(G472), .ZN(new_n699));
  NOR2_X1   g513(.A1(new_n694), .A2(new_n699), .ZN(new_n700));
  NOR2_X1   g514(.A1(new_n692), .A2(KEYINPUT99), .ZN(new_n701));
  NOR4_X1   g515(.A1(new_n690), .A2(new_n693), .A3(new_n700), .A4(new_n701), .ZN(new_n702));
  NAND3_X1  g516(.A1(new_n683), .A2(new_n686), .A3(new_n702), .ZN(new_n703));
  XNOR2_X1  g517(.A(new_n703), .B(G143), .ZN(G45));
  AOI21_X1  g518(.A(new_n627), .B1(new_n624), .B2(new_n625), .ZN(new_n705));
  NOR3_X1   g519(.A1(new_n691), .A2(new_n705), .A3(new_n667), .ZN(new_n706));
  AND4_X1   g520(.A1(new_n306), .A2(new_n664), .A3(new_n665), .A4(new_n706), .ZN(new_n707));
  XOR2_X1   g521(.A(KEYINPUT101), .B(G146), .Z(new_n708));
  XNOR2_X1  g522(.A(new_n707), .B(new_n708), .ZN(G48));
  AOI21_X1  g523(.A(new_n286), .B1(new_n673), .B2(new_n674), .ZN(new_n710));
  NAND2_X1  g524(.A1(new_n487), .A2(new_n484), .ZN(new_n711));
  AOI22_X1  g525(.A1(new_n711), .A2(new_n440), .B1(new_n482), .B2(new_n501), .ZN(new_n712));
  OAI21_X1  g526(.A(G469), .B1(new_n712), .B2(new_n189), .ZN(new_n713));
  NAND3_X1  g527(.A1(new_n713), .A2(new_n516), .A3(new_n509), .ZN(new_n714));
  INV_X1    g528(.A(KEYINPUT102), .ZN(new_n715));
  NAND2_X1  g529(.A1(new_n714), .A2(new_n715), .ZN(new_n716));
  NAND4_X1  g530(.A1(new_n713), .A2(KEYINPUT102), .A3(new_n509), .A4(new_n516), .ZN(new_n717));
  NAND2_X1  g531(.A1(new_n716), .A2(new_n717), .ZN(new_n718));
  NOR3_X1   g532(.A1(new_n710), .A2(new_n718), .A3(new_n549), .ZN(new_n719));
  NAND2_X1  g533(.A1(new_n719), .A2(new_n631), .ZN(new_n720));
  XNOR2_X1  g534(.A(KEYINPUT41), .B(G113), .ZN(new_n721));
  XNOR2_X1  g535(.A(new_n720), .B(new_n721), .ZN(G15));
  NAND2_X1  g536(.A1(new_n719), .A2(new_n650), .ZN(new_n723));
  XNOR2_X1  g537(.A(new_n723), .B(G116), .ZN(G18));
  NAND4_X1  g538(.A1(new_n659), .A2(new_n421), .A3(new_n428), .A4(new_n434), .ZN(new_n725));
  NOR2_X1   g539(.A1(new_n710), .A2(new_n725), .ZN(new_n726));
  AND3_X1   g540(.A1(new_n713), .A2(new_n516), .A3(new_n509), .ZN(new_n727));
  AND2_X1   g541(.A1(new_n609), .A2(new_n727), .ZN(new_n728));
  NAND2_X1  g542(.A1(new_n726), .A2(new_n728), .ZN(new_n729));
  XNOR2_X1  g543(.A(new_n729), .B(G119), .ZN(G21));
  NAND3_X1  g544(.A1(new_n716), .A2(new_n434), .A3(new_n717), .ZN(new_n731));
  XOR2_X1   g545(.A(KEYINPUT103), .B(G472), .Z(new_n732));
  OAI21_X1  g546(.A(new_n732), .B1(new_n303), .B2(new_n189), .ZN(new_n733));
  NAND2_X1  g547(.A1(new_n264), .A2(new_n271), .ZN(new_n734));
  OAI21_X1  g548(.A(new_n734), .B1(new_n291), .B2(new_n296), .ZN(new_n735));
  NAND2_X1  g549(.A1(new_n735), .A2(new_n298), .ZN(new_n736));
  NAND3_X1  g550(.A1(new_n550), .A2(new_n733), .A3(new_n736), .ZN(new_n737));
  NOR2_X1   g551(.A1(new_n731), .A2(new_n737), .ZN(new_n738));
  NAND3_X1  g552(.A1(new_n609), .A2(new_n648), .A3(new_n613), .ZN(new_n739));
  INV_X1    g553(.A(new_n739), .ZN(new_n740));
  NAND2_X1  g554(.A1(new_n738), .A2(new_n740), .ZN(new_n741));
  XNOR2_X1  g555(.A(new_n741), .B(G122), .ZN(G24));
  NAND4_X1  g556(.A1(new_n687), .A2(new_n706), .A3(new_n551), .A4(new_n727), .ZN(new_n743));
  NAND3_X1  g557(.A1(new_n733), .A2(new_n736), .A3(new_n659), .ZN(new_n744));
  INV_X1    g558(.A(KEYINPUT104), .ZN(new_n745));
  NAND2_X1  g559(.A1(new_n744), .A2(new_n745), .ZN(new_n746));
  NAND4_X1  g560(.A1(new_n733), .A2(new_n736), .A3(KEYINPUT104), .A4(new_n659), .ZN(new_n747));
  AOI21_X1  g561(.A(new_n743), .B1(new_n746), .B2(new_n747), .ZN(new_n748));
  XNOR2_X1  g562(.A(new_n748), .B(new_n380), .ZN(G27));
  NAND3_X1  g563(.A1(new_n606), .A2(new_n551), .A3(new_n608), .ZN(new_n750));
  NOR2_X1   g564(.A1(new_n750), .A2(new_n517), .ZN(new_n751));
  NAND4_X1  g565(.A1(new_n751), .A2(new_n306), .A3(new_n550), .A4(new_n706), .ZN(new_n752));
  INV_X1    g566(.A(KEYINPUT42), .ZN(new_n753));
  NAND2_X1  g567(.A1(new_n752), .A2(new_n753), .ZN(new_n754));
  NAND3_X1  g568(.A1(new_n306), .A2(KEYINPUT105), .A3(new_n550), .ZN(new_n755));
  INV_X1    g569(.A(KEYINPUT105), .ZN(new_n756));
  OAI21_X1  g570(.A(new_n756), .B1(new_n710), .B2(new_n549), .ZN(new_n757));
  NAND3_X1  g571(.A1(new_n613), .A2(new_n629), .A3(new_n668), .ZN(new_n758));
  NOR4_X1   g572(.A1(new_n750), .A2(new_n517), .A3(new_n758), .A4(new_n753), .ZN(new_n759));
  NAND3_X1  g573(.A1(new_n755), .A2(new_n757), .A3(new_n759), .ZN(new_n760));
  NAND2_X1  g574(.A1(new_n754), .A2(new_n760), .ZN(new_n761));
  XNOR2_X1  g575(.A(new_n761), .B(G131), .ZN(G33));
  NOR2_X1   g576(.A1(new_n710), .A2(new_n549), .ZN(new_n763));
  NAND3_X1  g577(.A1(new_n763), .A2(new_n669), .A3(new_n751), .ZN(new_n764));
  XNOR2_X1  g578(.A(new_n764), .B(G134), .ZN(G36));
  NAND2_X1  g579(.A1(new_n691), .A2(new_n629), .ZN(new_n766));
  NAND2_X1  g580(.A1(KEYINPUT106), .A2(KEYINPUT43), .ZN(new_n767));
  NOR2_X1   g581(.A1(KEYINPUT106), .A2(KEYINPUT43), .ZN(new_n768));
  INV_X1    g582(.A(new_n768), .ZN(new_n769));
  NAND3_X1  g583(.A1(new_n766), .A2(new_n767), .A3(new_n769), .ZN(new_n770));
  OAI21_X1  g584(.A(new_n770), .B1(new_n766), .B2(new_n769), .ZN(new_n771));
  NOR3_X1   g585(.A1(new_n771), .A2(new_n633), .A3(new_n658), .ZN(new_n772));
  AOI21_X1  g586(.A(new_n750), .B1(new_n772), .B2(KEYINPUT44), .ZN(new_n773));
  OAI21_X1  g587(.A(new_n773), .B1(KEYINPUT44), .B2(new_n772), .ZN(new_n774));
  OAI21_X1  g588(.A(new_n485), .B1(new_n503), .B2(new_n504), .ZN(new_n775));
  XNOR2_X1  g589(.A(new_n775), .B(KEYINPUT45), .ZN(new_n776));
  AOI21_X1  g590(.A(new_n510), .B1(new_n776), .B2(G469), .ZN(new_n777));
  OR2_X1    g591(.A1(new_n777), .A2(KEYINPUT46), .ZN(new_n778));
  INV_X1    g592(.A(new_n509), .ZN(new_n779));
  AOI21_X1  g593(.A(new_n779), .B1(new_n777), .B2(KEYINPUT46), .ZN(new_n780));
  AOI21_X1  g594(.A(new_n515), .B1(new_n778), .B2(new_n780), .ZN(new_n781));
  NAND2_X1  g595(.A1(new_n781), .A2(new_n680), .ZN(new_n782));
  NOR2_X1   g596(.A1(new_n774), .A2(new_n782), .ZN(new_n783));
  XNOR2_X1  g597(.A(new_n783), .B(new_n195), .ZN(G39));
  XNOR2_X1  g598(.A(new_n781), .B(KEYINPUT47), .ZN(new_n785));
  NOR4_X1   g599(.A1(new_n306), .A2(new_n550), .A3(new_n758), .A4(new_n750), .ZN(new_n786));
  NAND2_X1  g600(.A1(new_n785), .A2(new_n786), .ZN(new_n787));
  XNOR2_X1  g601(.A(new_n787), .B(G140), .ZN(G42));
  INV_X1    g602(.A(new_n430), .ZN(new_n789));
  NOR3_X1   g603(.A1(new_n771), .A2(new_n789), .A3(new_n737), .ZN(new_n790));
  NAND4_X1  g604(.A1(new_n790), .A2(new_n690), .A3(new_n552), .A4(new_n727), .ZN(new_n791));
  INV_X1    g605(.A(KEYINPUT112), .ZN(new_n792));
  INV_X1    g606(.A(KEYINPUT50), .ZN(new_n793));
  NAND2_X1  g607(.A1(new_n792), .A2(new_n793), .ZN(new_n794));
  AND2_X1   g608(.A1(new_n791), .A2(new_n794), .ZN(new_n795));
  NOR2_X1   g609(.A1(new_n791), .A2(new_n794), .ZN(new_n796));
  OAI22_X1  g610(.A1(new_n795), .A2(new_n796), .B1(new_n792), .B2(new_n793), .ZN(new_n797));
  NOR2_X1   g611(.A1(new_n771), .A2(new_n789), .ZN(new_n798));
  NOR2_X1   g612(.A1(new_n750), .A2(new_n714), .ZN(new_n799));
  NAND2_X1  g613(.A1(new_n798), .A2(new_n799), .ZN(new_n800));
  XOR2_X1   g614(.A(new_n800), .B(KEYINPUT113), .Z(new_n801));
  NAND2_X1  g615(.A1(new_n746), .A2(new_n747), .ZN(new_n802));
  NAND2_X1  g616(.A1(new_n801), .A2(new_n802), .ZN(new_n803));
  NOR2_X1   g617(.A1(new_n549), .A2(new_n789), .ZN(new_n804));
  AND3_X1   g618(.A1(new_n700), .A2(new_n799), .A3(new_n804), .ZN(new_n805));
  NAND3_X1  g619(.A1(new_n805), .A2(new_n691), .A3(new_n705), .ZN(new_n806));
  XOR2_X1   g620(.A(new_n806), .B(KEYINPUT114), .Z(new_n807));
  NAND3_X1  g621(.A1(new_n797), .A2(new_n803), .A3(new_n807), .ZN(new_n808));
  NAND2_X1  g622(.A1(new_n713), .A2(new_n509), .ZN(new_n809));
  INV_X1    g623(.A(new_n809), .ZN(new_n810));
  AOI21_X1  g624(.A(new_n785), .B1(new_n515), .B2(new_n810), .ZN(new_n811));
  INV_X1    g625(.A(new_n750), .ZN(new_n812));
  NAND2_X1  g626(.A1(new_n790), .A2(new_n812), .ZN(new_n813));
  NOR2_X1   g627(.A1(new_n811), .A2(new_n813), .ZN(new_n814));
  INV_X1    g628(.A(KEYINPUT115), .ZN(new_n815));
  INV_X1    g629(.A(KEYINPUT51), .ZN(new_n816));
  OAI22_X1  g630(.A1(new_n808), .A2(new_n814), .B1(new_n815), .B2(new_n816), .ZN(new_n817));
  OAI21_X1  g631(.A(new_n817), .B1(KEYINPUT115), .B2(KEYINPUT51), .ZN(new_n818));
  INV_X1    g632(.A(KEYINPUT116), .ZN(new_n819));
  INV_X1    g633(.A(new_n801), .ZN(new_n820));
  NAND2_X1  g634(.A1(new_n755), .A2(new_n757), .ZN(new_n821));
  OAI21_X1  g635(.A(new_n819), .B1(new_n820), .B2(new_n821), .ZN(new_n822));
  INV_X1    g636(.A(new_n821), .ZN(new_n823));
  NAND3_X1  g637(.A1(new_n801), .A2(KEYINPUT116), .A3(new_n823), .ZN(new_n824));
  AND3_X1   g638(.A1(new_n822), .A2(KEYINPUT48), .A3(new_n824), .ZN(new_n825));
  AOI21_X1  g639(.A(new_n822), .B1(KEYINPUT48), .B2(new_n824), .ZN(new_n826));
  NAND3_X1  g640(.A1(new_n805), .A2(new_n613), .A3(new_n629), .ZN(new_n827));
  NAND2_X1  g641(.A1(new_n790), .A2(new_n728), .ZN(new_n828));
  NAND4_X1  g642(.A1(new_n827), .A2(G952), .A3(new_n361), .A4(new_n828), .ZN(new_n829));
  NOR3_X1   g643(.A1(new_n825), .A2(new_n826), .A3(new_n829), .ZN(new_n830));
  OAI211_X1 g644(.A(new_n815), .B(new_n816), .C1(new_n808), .C2(new_n814), .ZN(new_n831));
  NAND3_X1  g645(.A1(new_n818), .A2(new_n830), .A3(new_n831), .ZN(new_n832));
  NOR2_X1   g646(.A1(new_n659), .A2(new_n667), .ZN(new_n833));
  AND3_X1   g647(.A1(new_n665), .A2(KEYINPUT109), .A3(new_n833), .ZN(new_n834));
  AOI21_X1  g648(.A(KEYINPUT109), .B1(new_n665), .B2(new_n833), .ZN(new_n835));
  OAI221_X1 g649(.A(new_n740), .B1(new_n694), .B2(new_n699), .C1(new_n834), .C2(new_n835), .ZN(new_n836));
  NOR2_X1   g650(.A1(new_n707), .A2(new_n748), .ZN(new_n837));
  NAND3_X1  g651(.A1(new_n678), .A2(new_n836), .A3(new_n837), .ZN(new_n838));
  INV_X1    g652(.A(KEYINPUT52), .ZN(new_n839));
  NAND2_X1  g653(.A1(new_n838), .A2(new_n839), .ZN(new_n840));
  NAND4_X1  g654(.A1(new_n678), .A2(new_n836), .A3(new_n837), .A4(KEYINPUT52), .ZN(new_n841));
  NAND2_X1  g655(.A1(new_n840), .A2(new_n841), .ZN(new_n842));
  NOR3_X1   g656(.A1(new_n750), .A2(new_n517), .A3(new_n758), .ZN(new_n843));
  NAND2_X1  g657(.A1(new_n802), .A2(new_n843), .ZN(new_n844));
  NOR2_X1   g658(.A1(new_n750), .A2(new_n658), .ZN(new_n845));
  NAND4_X1  g659(.A1(new_n644), .A2(KEYINPUT108), .A3(new_n421), .A4(new_n668), .ZN(new_n846));
  INV_X1    g660(.A(KEYINPUT108), .ZN(new_n847));
  NAND2_X1  g661(.A1(new_n421), .A2(new_n668), .ZN(new_n848));
  OAI21_X1  g662(.A(new_n847), .B1(new_n848), .B2(new_n643), .ZN(new_n849));
  NAND4_X1  g663(.A1(new_n676), .A2(new_n845), .A3(new_n846), .A4(new_n849), .ZN(new_n850));
  AND3_X1   g664(.A1(new_n844), .A2(new_n764), .A3(new_n850), .ZN(new_n851));
  AOI211_X1 g665(.A(new_n552), .B(new_n433), .C1(new_n606), .C2(new_n608), .ZN(new_n852));
  OAI21_X1  g666(.A(new_n630), .B1(new_n356), .B2(new_n613), .ZN(new_n853));
  NAND4_X1  g667(.A1(new_n852), .A2(new_n634), .A3(new_n633), .A4(new_n853), .ZN(new_n854));
  NAND3_X1  g668(.A1(new_n610), .A2(new_n660), .A3(new_n854), .ZN(new_n855));
  INV_X1    g669(.A(new_n855), .ZN(new_n856));
  NAND2_X1  g670(.A1(new_n851), .A2(new_n856), .ZN(new_n857));
  AOI22_X1  g671(.A1(new_n719), .A2(new_n631), .B1(new_n728), .B2(new_n726), .ZN(new_n858));
  AOI22_X1  g672(.A1(new_n719), .A2(new_n650), .B1(new_n738), .B2(new_n740), .ZN(new_n859));
  NAND3_X1  g673(.A1(new_n761), .A2(new_n858), .A3(new_n859), .ZN(new_n860));
  NOR2_X1   g674(.A1(new_n857), .A2(new_n860), .ZN(new_n861));
  AOI21_X1  g675(.A(KEYINPUT53), .B1(new_n842), .B2(new_n861), .ZN(new_n862));
  INV_X1    g676(.A(KEYINPUT111), .ZN(new_n863));
  AND2_X1   g677(.A1(new_n840), .A2(new_n841), .ZN(new_n864));
  AND3_X1   g678(.A1(new_n761), .A2(new_n858), .A3(new_n859), .ZN(new_n865));
  INV_X1    g679(.A(KEYINPUT110), .ZN(new_n866));
  NAND3_X1  g680(.A1(new_n844), .A2(new_n764), .A3(new_n850), .ZN(new_n867));
  OAI21_X1  g681(.A(new_n866), .B1(new_n867), .B2(new_n855), .ZN(new_n868));
  NOR4_X1   g682(.A1(new_n710), .A2(new_n549), .A3(new_n750), .A4(new_n517), .ZN(new_n869));
  AOI22_X1  g683(.A1(new_n869), .A2(new_n669), .B1(new_n802), .B2(new_n843), .ZN(new_n870));
  NAND4_X1  g684(.A1(new_n856), .A2(new_n870), .A3(KEYINPUT110), .A4(new_n850), .ZN(new_n871));
  NAND4_X1  g685(.A1(new_n865), .A2(new_n868), .A3(new_n871), .A4(KEYINPUT53), .ZN(new_n872));
  OAI21_X1  g686(.A(new_n863), .B1(new_n864), .B2(new_n872), .ZN(new_n873));
  AOI21_X1  g687(.A(KEYINPUT110), .B1(new_n851), .B2(new_n856), .ZN(new_n874));
  NOR3_X1   g688(.A1(new_n867), .A2(new_n866), .A3(new_n855), .ZN(new_n875));
  NAND4_X1  g689(.A1(new_n761), .A2(KEYINPUT53), .A3(new_n858), .A4(new_n859), .ZN(new_n876));
  NOR3_X1   g690(.A1(new_n874), .A2(new_n875), .A3(new_n876), .ZN(new_n877));
  NAND3_X1  g691(.A1(new_n877), .A2(KEYINPUT111), .A3(new_n842), .ZN(new_n878));
  AOI21_X1  g692(.A(new_n862), .B1(new_n873), .B2(new_n878), .ZN(new_n879));
  INV_X1    g693(.A(KEYINPUT54), .ZN(new_n880));
  NAND2_X1  g694(.A1(new_n879), .A2(new_n880), .ZN(new_n881));
  INV_X1    g695(.A(new_n862), .ZN(new_n882));
  NAND3_X1  g696(.A1(new_n842), .A2(KEYINPUT53), .A3(new_n861), .ZN(new_n883));
  NAND2_X1  g697(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  NAND2_X1  g698(.A1(new_n884), .A2(KEYINPUT54), .ZN(new_n885));
  NAND2_X1  g699(.A1(new_n881), .A2(new_n885), .ZN(new_n886));
  OAI22_X1  g700(.A1(new_n832), .A2(new_n886), .B1(G952), .B2(G953), .ZN(new_n887));
  XOR2_X1   g701(.A(new_n809), .B(KEYINPUT49), .Z(new_n888));
  NAND3_X1  g702(.A1(new_n690), .A2(new_n700), .A3(new_n888), .ZN(new_n889));
  NOR4_X1   g703(.A1(new_n766), .A2(new_n549), .A3(new_n552), .A4(new_n515), .ZN(new_n890));
  XNOR2_X1  g704(.A(new_n890), .B(KEYINPUT107), .ZN(new_n891));
  OAI21_X1  g705(.A(new_n887), .B1(new_n889), .B2(new_n891), .ZN(G75));
  NAND2_X1  g706(.A1(new_n572), .A2(new_n585), .ZN(new_n893));
  XNOR2_X1  g707(.A(new_n893), .B(new_n581), .ZN(new_n894));
  XNOR2_X1  g708(.A(new_n894), .B(KEYINPUT55), .ZN(new_n895));
  INV_X1    g709(.A(new_n895), .ZN(new_n896));
  NOR3_X1   g710(.A1(new_n879), .A2(new_n188), .A3(new_n553), .ZN(new_n897));
  OAI21_X1  g711(.A(new_n896), .B1(new_n897), .B2(KEYINPUT56), .ZN(new_n898));
  NOR3_X1   g712(.A1(new_n864), .A2(new_n872), .A3(new_n863), .ZN(new_n899));
  AOI21_X1  g713(.A(KEYINPUT111), .B1(new_n877), .B2(new_n842), .ZN(new_n900));
  OAI21_X1  g714(.A(new_n882), .B1(new_n899), .B2(new_n900), .ZN(new_n901));
  NAND3_X1  g715(.A1(new_n901), .A2(new_n189), .A3(new_n554), .ZN(new_n902));
  INV_X1    g716(.A(KEYINPUT56), .ZN(new_n903));
  NAND3_X1  g717(.A1(new_n902), .A2(new_n903), .A3(new_n895), .ZN(new_n904));
  NOR2_X1   g718(.A1(new_n361), .A2(G952), .ZN(new_n905));
  INV_X1    g719(.A(new_n905), .ZN(new_n906));
  NAND3_X1  g720(.A1(new_n898), .A2(new_n904), .A3(new_n906), .ZN(new_n907));
  NAND2_X1  g721(.A1(new_n907), .A2(KEYINPUT117), .ZN(new_n908));
  INV_X1    g722(.A(KEYINPUT117), .ZN(new_n909));
  NAND4_X1  g723(.A1(new_n898), .A2(new_n909), .A3(new_n904), .A4(new_n906), .ZN(new_n910));
  NAND2_X1  g724(.A1(new_n908), .A2(new_n910), .ZN(G51));
  INV_X1    g725(.A(KEYINPUT118), .ZN(new_n912));
  NAND2_X1  g726(.A1(new_n776), .A2(G469), .ZN(new_n913));
  NOR3_X1   g727(.A1(new_n879), .A2(new_n188), .A3(new_n913), .ZN(new_n914));
  XNOR2_X1  g728(.A(new_n510), .B(KEYINPUT57), .ZN(new_n915));
  NAND2_X1  g729(.A1(new_n873), .A2(new_n878), .ZN(new_n916));
  AOI21_X1  g730(.A(new_n880), .B1(new_n916), .B2(new_n882), .ZN(new_n917));
  AOI211_X1 g731(.A(KEYINPUT54), .B(new_n862), .C1(new_n873), .C2(new_n878), .ZN(new_n918));
  OAI21_X1  g732(.A(new_n915), .B1(new_n917), .B2(new_n918), .ZN(new_n919));
  INV_X1    g733(.A(new_n712), .ZN(new_n920));
  AOI21_X1  g734(.A(new_n914), .B1(new_n919), .B2(new_n920), .ZN(new_n921));
  OAI21_X1  g735(.A(new_n912), .B1(new_n921), .B2(new_n905), .ZN(new_n922));
  NAND2_X1  g736(.A1(new_n901), .A2(KEYINPUT54), .ZN(new_n923));
  NAND2_X1  g737(.A1(new_n923), .A2(new_n881), .ZN(new_n924));
  AOI21_X1  g738(.A(new_n712), .B1(new_n924), .B2(new_n915), .ZN(new_n925));
  OAI211_X1 g739(.A(KEYINPUT118), .B(new_n906), .C1(new_n925), .C2(new_n914), .ZN(new_n926));
  NAND2_X1  g740(.A1(new_n922), .A2(new_n926), .ZN(G54));
  INV_X1    g741(.A(KEYINPUT58), .ZN(new_n928));
  OAI21_X1  g742(.A(KEYINPUT119), .B1(new_n928), .B2(new_n639), .ZN(new_n929));
  OR3_X1    g743(.A1(new_n928), .A2(new_n639), .A3(KEYINPUT119), .ZN(new_n930));
  NAND4_X1  g744(.A1(new_n901), .A2(new_n189), .A3(new_n929), .A4(new_n930), .ZN(new_n931));
  INV_X1    g745(.A(new_n417), .ZN(new_n932));
  AND2_X1   g746(.A1(new_n931), .A2(new_n932), .ZN(new_n933));
  NOR2_X1   g747(.A1(new_n931), .A2(new_n932), .ZN(new_n934));
  NOR3_X1   g748(.A1(new_n933), .A2(new_n934), .A3(new_n905), .ZN(G60));
  NAND2_X1  g749(.A1(G478), .A2(G902), .ZN(new_n936));
  XOR2_X1   g750(.A(new_n936), .B(KEYINPUT59), .Z(new_n937));
  INV_X1    g751(.A(new_n937), .ZN(new_n938));
  AND3_X1   g752(.A1(new_n924), .A2(new_n624), .A3(new_n938), .ZN(new_n939));
  AOI21_X1  g753(.A(new_n624), .B1(new_n886), .B2(new_n938), .ZN(new_n940));
  NOR3_X1   g754(.A1(new_n939), .A2(new_n940), .A3(new_n905), .ZN(G63));
  XNOR2_X1  g755(.A(KEYINPUT121), .B(KEYINPUT60), .ZN(new_n942));
  NAND2_X1  g756(.A1(G217), .A2(G902), .ZN(new_n943));
  XNOR2_X1  g757(.A(new_n942), .B(new_n943), .ZN(new_n944));
  NOR2_X1   g758(.A1(new_n879), .A2(new_n944), .ZN(new_n945));
  NAND2_X1  g759(.A1(new_n945), .A2(new_n655), .ZN(new_n946));
  OAI211_X1 g760(.A(new_n538), .B(new_n537), .C1(new_n879), .C2(new_n944), .ZN(new_n947));
  NAND3_X1  g761(.A1(new_n946), .A2(new_n906), .A3(new_n947), .ZN(new_n948));
  INV_X1    g762(.A(KEYINPUT120), .ZN(new_n949));
  AND3_X1   g763(.A1(new_n948), .A2(new_n949), .A3(KEYINPUT61), .ZN(new_n950));
  AOI21_X1  g764(.A(KEYINPUT61), .B1(new_n948), .B2(new_n949), .ZN(new_n951));
  NOR2_X1   g765(.A1(new_n950), .A2(new_n951), .ZN(G66));
  NAND2_X1  g766(.A1(G224), .A2(G953), .ZN(new_n953));
  NOR2_X1   g767(.A1(new_n432), .A2(new_n953), .ZN(new_n954));
  AND3_X1   g768(.A1(new_n856), .A2(new_n858), .A3(new_n859), .ZN(new_n955));
  AOI21_X1  g769(.A(new_n954), .B1(new_n955), .B2(new_n361), .ZN(new_n956));
  OAI21_X1  g770(.A(new_n893), .B1(G898), .B2(new_n361), .ZN(new_n957));
  XNOR2_X1  g771(.A(new_n956), .B(new_n957), .ZN(G69));
  NAND2_X1  g772(.A1(new_n678), .A2(new_n837), .ZN(new_n959));
  NOR2_X1   g773(.A1(new_n783), .A2(new_n959), .ZN(new_n960));
  INV_X1    g774(.A(KEYINPUT125), .ZN(new_n961));
  XNOR2_X1  g775(.A(new_n960), .B(new_n961), .ZN(new_n962));
  NAND4_X1  g776(.A1(new_n781), .A2(new_n823), .A3(new_n680), .A4(new_n740), .ZN(new_n963));
  NAND4_X1  g777(.A1(new_n787), .A2(new_n761), .A3(new_n764), .A4(new_n963), .ZN(new_n964));
  NOR3_X1   g778(.A1(new_n962), .A2(G953), .A3(new_n964), .ZN(new_n965));
  XOR2_X1   g779(.A(new_n283), .B(new_n409), .Z(new_n966));
  AOI21_X1  g780(.A(new_n966), .B1(G900), .B2(G953), .ZN(new_n967));
  INV_X1    g781(.A(new_n967), .ZN(new_n968));
  OAI21_X1  g782(.A(KEYINPUT124), .B1(new_n965), .B2(new_n968), .ZN(new_n969));
  OAI21_X1  g783(.A(G953), .B1(new_n437), .B2(new_n666), .ZN(new_n970));
  NAND2_X1  g784(.A1(new_n969), .A2(new_n970), .ZN(new_n971));
  INV_X1    g785(.A(new_n783), .ZN(new_n972));
  NAND4_X1  g786(.A1(new_n684), .A2(new_n763), .A3(new_n812), .A4(new_n853), .ZN(new_n973));
  XNOR2_X1  g787(.A(new_n973), .B(KEYINPUT123), .ZN(new_n974));
  NAND3_X1  g788(.A1(new_n972), .A2(new_n974), .A3(new_n787), .ZN(new_n975));
  INV_X1    g789(.A(KEYINPUT62), .ZN(new_n976));
  OR2_X1    g790(.A1(new_n976), .A2(KEYINPUT122), .ZN(new_n977));
  AND2_X1   g791(.A1(new_n703), .A2(new_n977), .ZN(new_n978));
  INV_X1    g792(.A(new_n959), .ZN(new_n979));
  NAND2_X1  g793(.A1(new_n978), .A2(new_n979), .ZN(new_n980));
  NAND3_X1  g794(.A1(new_n980), .A2(KEYINPUT122), .A3(new_n976), .ZN(new_n981));
  NAND2_X1  g795(.A1(new_n976), .A2(KEYINPUT122), .ZN(new_n982));
  NAND3_X1  g796(.A1(new_n978), .A2(new_n979), .A3(new_n982), .ZN(new_n983));
  AOI21_X1  g797(.A(new_n975), .B1(new_n981), .B2(new_n983), .ZN(new_n984));
  OAI21_X1  g798(.A(new_n966), .B1(new_n984), .B2(G953), .ZN(new_n985));
  OAI21_X1  g799(.A(new_n985), .B1(new_n965), .B2(new_n968), .ZN(new_n986));
  XNOR2_X1  g800(.A(new_n971), .B(new_n986), .ZN(G72));
  XNOR2_X1  g801(.A(KEYINPUT126), .B(KEYINPUT63), .ZN(new_n988));
  NOR2_X1   g802(.A1(new_n187), .A2(new_n422), .ZN(new_n989));
  XOR2_X1   g803(.A(new_n988), .B(new_n989), .Z(new_n990));
  INV_X1    g804(.A(new_n990), .ZN(new_n991));
  NOR2_X1   g805(.A1(new_n284), .A2(new_n270), .ZN(new_n992));
  OAI211_X1 g806(.A(new_n884), .B(new_n991), .C1(new_n992), .C2(new_n697), .ZN(new_n993));
  NOR2_X1   g807(.A1(new_n962), .A2(new_n964), .ZN(new_n994));
  AOI21_X1  g808(.A(new_n990), .B1(new_n994), .B2(new_n955), .ZN(new_n995));
  NAND2_X1  g809(.A1(new_n284), .A2(new_n271), .ZN(new_n996));
  OAI211_X1 g810(.A(new_n906), .B(new_n993), .C1(new_n995), .C2(new_n996), .ZN(new_n997));
  NAND2_X1  g811(.A1(new_n984), .A2(new_n955), .ZN(new_n998));
  NAND2_X1  g812(.A1(new_n998), .A2(new_n991), .ZN(new_n999));
  NOR2_X1   g813(.A1(new_n284), .A2(new_n271), .ZN(new_n1000));
  NAND2_X1  g814(.A1(new_n999), .A2(new_n1000), .ZN(new_n1001));
  NAND2_X1  g815(.A1(new_n1001), .A2(KEYINPUT127), .ZN(new_n1002));
  INV_X1    g816(.A(KEYINPUT127), .ZN(new_n1003));
  NAND3_X1  g817(.A1(new_n999), .A2(new_n1003), .A3(new_n1000), .ZN(new_n1004));
  AOI21_X1  g818(.A(new_n997), .B1(new_n1002), .B2(new_n1004), .ZN(G57));
endmodule


