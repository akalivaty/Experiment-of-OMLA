//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 0 0 0 0 0 1 1 1 1 0 0 0 1 0 1 1 1 1 1 0 1 1 0 0 0 1 1 1 1 1 0 0 1 0 0 1 1 1 0 1 1 0 0 1 1 1 0 1 1 1 1 1 1 0 0 1 1 1 1 0 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:40:43 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n244, new_n245,
    new_n247, new_n248, new_n249, new_n250, new_n251, new_n252, new_n253,
    new_n254, new_n255, new_n256, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1184, new_n1185, new_n1186, new_n1187,
    new_n1188, new_n1189, new_n1190, new_n1191, new_n1192, new_n1193,
    new_n1194, new_n1195, new_n1196, new_n1197, new_n1198, new_n1199,
    new_n1200, new_n1201, new_n1202, new_n1203, new_n1204, new_n1205,
    new_n1206, new_n1207, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1215, new_n1217, new_n1219, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1278, new_n1279, new_n1280, new_n1281,
    new_n1282, new_n1283, new_n1284, new_n1285, new_n1286, new_n1287,
    new_n1288, new_n1289;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0005(.A1(G1), .A2(G20), .ZN(new_n206));
  XNOR2_X1  g0006(.A(KEYINPUT65), .B(G68), .ZN(new_n207));
  INV_X1    g0007(.A(new_n207), .ZN(new_n208));
  INV_X1    g0008(.A(G58), .ZN(new_n209));
  INV_X1    g0009(.A(G232), .ZN(new_n210));
  INV_X1    g0010(.A(G107), .ZN(new_n211));
  INV_X1    g0011(.A(G264), .ZN(new_n212));
  OAI22_X1  g0012(.A1(new_n209), .A2(new_n210), .B1(new_n211), .B2(new_n212), .ZN(new_n213));
  INV_X1    g0013(.A(KEYINPUT66), .ZN(new_n214));
  AOI22_X1  g0014(.A1(new_n208), .A2(G238), .B1(new_n213), .B2(new_n214), .ZN(new_n215));
  OAI21_X1  g0015(.A(new_n215), .B1(new_n214), .B2(new_n213), .ZN(new_n216));
  AOI22_X1  g0016(.A1(G97), .A2(G257), .B1(G116), .B2(G270), .ZN(new_n217));
  AOI22_X1  g0017(.A1(G50), .A2(G226), .B1(G87), .B2(G250), .ZN(new_n218));
  INV_X1    g0018(.A(G77), .ZN(new_n219));
  INV_X1    g0019(.A(G244), .ZN(new_n220));
  OAI211_X1 g0020(.A(new_n217), .B(new_n218), .C1(new_n219), .C2(new_n220), .ZN(new_n221));
  OAI21_X1  g0021(.A(new_n206), .B1(new_n216), .B2(new_n221), .ZN(new_n222));
  XOR2_X1   g0022(.A(new_n222), .B(KEYINPUT1), .Z(new_n223));
  NOR2_X1   g0023(.A1(new_n206), .A2(G13), .ZN(new_n224));
  OAI211_X1 g0024(.A(new_n224), .B(G250), .C1(G257), .C2(G264), .ZN(new_n225));
  XOR2_X1   g0025(.A(new_n225), .B(KEYINPUT0), .Z(new_n226));
  NAND2_X1  g0026(.A1(G1), .A2(G13), .ZN(new_n227));
  INV_X1    g0027(.A(G20), .ZN(new_n228));
  NOR2_X1   g0028(.A1(new_n227), .A2(new_n228), .ZN(new_n229));
  XNOR2_X1  g0029(.A(new_n229), .B(KEYINPUT64), .ZN(new_n230));
  INV_X1    g0030(.A(new_n201), .ZN(new_n231));
  NAND2_X1  g0031(.A1(new_n231), .A2(G50), .ZN(new_n232));
  INV_X1    g0032(.A(new_n232), .ZN(new_n233));
  AOI21_X1  g0033(.A(new_n226), .B1(new_n230), .B2(new_n233), .ZN(new_n234));
  NAND2_X1  g0034(.A1(new_n223), .A2(new_n234), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n235), .B(KEYINPUT67), .ZN(G361));
  XOR2_X1   g0036(.A(G264), .B(G270), .Z(new_n237));
  XNOR2_X1  g0037(.A(G250), .B(G257), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XNOR2_X1  g0039(.A(KEYINPUT68), .B(KEYINPUT69), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XNOR2_X1  g0041(.A(G238), .B(G244), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n242), .B(G232), .ZN(new_n243));
  XOR2_X1   g0043(.A(KEYINPUT2), .B(G226), .Z(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XOR2_X1   g0045(.A(new_n241), .B(new_n245), .Z(G358));
  XNOR2_X1  g0046(.A(G107), .B(G116), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n247), .B(KEYINPUT70), .ZN(new_n248));
  XNOR2_X1  g0048(.A(G87), .B(G97), .ZN(new_n249));
  XNOR2_X1  g0049(.A(new_n248), .B(new_n249), .ZN(new_n250));
  NAND2_X1  g0050(.A1(new_n202), .A2(G68), .ZN(new_n251));
  INV_X1    g0051(.A(G68), .ZN(new_n252));
  NAND2_X1  g0052(.A1(new_n252), .A2(G50), .ZN(new_n253));
  NAND2_X1  g0053(.A1(new_n251), .A2(new_n253), .ZN(new_n254));
  XNOR2_X1  g0054(.A(G58), .B(G77), .ZN(new_n255));
  XNOR2_X1  g0055(.A(new_n254), .B(new_n255), .ZN(new_n256));
  XNOR2_X1  g0056(.A(new_n250), .B(new_n256), .ZN(G351));
  INV_X1    g0057(.A(G1), .ZN(new_n258));
  OAI211_X1 g0058(.A(new_n258), .B(G274), .C1(G41), .C2(G45), .ZN(new_n259));
  XNOR2_X1  g0059(.A(new_n259), .B(KEYINPUT71), .ZN(new_n260));
  INV_X1    g0060(.A(G226), .ZN(new_n261));
  INV_X1    g0061(.A(G33), .ZN(new_n262));
  INV_X1    g0062(.A(G41), .ZN(new_n263));
  OAI211_X1 g0063(.A(G1), .B(G13), .C1(new_n262), .C2(new_n263), .ZN(new_n264));
  OAI21_X1  g0064(.A(new_n258), .B1(G41), .B2(G45), .ZN(new_n265));
  NAND2_X1  g0065(.A1(new_n264), .A2(new_n265), .ZN(new_n266));
  OAI21_X1  g0066(.A(new_n260), .B1(new_n261), .B2(new_n266), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n262), .A2(KEYINPUT3), .ZN(new_n268));
  INV_X1    g0068(.A(KEYINPUT3), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n269), .A2(G33), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n268), .A2(new_n270), .ZN(new_n271));
  INV_X1    g0071(.A(KEYINPUT72), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n271), .A2(new_n272), .ZN(new_n273));
  NAND3_X1  g0073(.A1(new_n268), .A2(new_n270), .A3(KEYINPUT72), .ZN(new_n274));
  AOI21_X1  g0074(.A(G1698), .B1(new_n273), .B2(new_n274), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n275), .A2(G222), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n273), .A2(new_n274), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n277), .A2(G1698), .ZN(new_n278));
  INV_X1    g0078(.A(G223), .ZN(new_n279));
  OAI221_X1 g0079(.A(new_n276), .B1(new_n219), .B2(new_n277), .C1(new_n278), .C2(new_n279), .ZN(new_n280));
  INV_X1    g0080(.A(new_n264), .ZN(new_n281));
  AOI21_X1  g0081(.A(new_n267), .B1(new_n280), .B2(new_n281), .ZN(new_n282));
  INV_X1    g0082(.A(new_n282), .ZN(new_n283));
  NOR2_X1   g0083(.A1(new_n283), .A2(G179), .ZN(new_n284));
  NAND3_X1  g0084(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n285));
  INV_X1    g0085(.A(KEYINPUT73), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n285), .A2(new_n286), .ZN(new_n287));
  NAND4_X1  g0087(.A1(KEYINPUT73), .A2(G1), .A3(G20), .A4(G33), .ZN(new_n288));
  NAND3_X1  g0088(.A1(new_n287), .A2(new_n227), .A3(new_n288), .ZN(new_n289));
  AOI21_X1  g0089(.A(new_n289), .B1(new_n258), .B2(G20), .ZN(new_n290));
  NAND2_X1  g0090(.A1(new_n290), .A2(G50), .ZN(new_n291));
  NAND3_X1  g0091(.A1(new_n258), .A2(G13), .A3(G20), .ZN(new_n292));
  INV_X1    g0092(.A(new_n292), .ZN(new_n293));
  NAND2_X1  g0093(.A1(new_n293), .A2(new_n202), .ZN(new_n294));
  XNOR2_X1  g0094(.A(KEYINPUT8), .B(G58), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n228), .A2(G33), .ZN(new_n296));
  INV_X1    g0096(.A(G150), .ZN(new_n297));
  NOR2_X1   g0097(.A1(G20), .A2(G33), .ZN(new_n298));
  INV_X1    g0098(.A(new_n298), .ZN(new_n299));
  OAI22_X1  g0099(.A1(new_n295), .A2(new_n296), .B1(new_n297), .B2(new_n299), .ZN(new_n300));
  AOI21_X1  g0100(.A(new_n300), .B1(G20), .B2(new_n203), .ZN(new_n301));
  INV_X1    g0101(.A(new_n289), .ZN(new_n302));
  OAI211_X1 g0102(.A(new_n291), .B(new_n294), .C1(new_n301), .C2(new_n302), .ZN(new_n303));
  OAI21_X1  g0103(.A(new_n303), .B1(new_n282), .B2(G169), .ZN(new_n304));
  NOR2_X1   g0104(.A1(new_n284), .A2(new_n304), .ZN(new_n305));
  XNOR2_X1  g0105(.A(new_n303), .B(KEYINPUT9), .ZN(new_n306));
  INV_X1    g0106(.A(G200), .ZN(new_n307));
  OAI21_X1  g0107(.A(new_n306), .B1(new_n307), .B2(new_n282), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n282), .A2(G190), .ZN(new_n309));
  INV_X1    g0109(.A(new_n309), .ZN(new_n310));
  OAI21_X1  g0110(.A(KEYINPUT10), .B1(new_n308), .B2(new_n310), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n283), .A2(G200), .ZN(new_n312));
  INV_X1    g0112(.A(KEYINPUT10), .ZN(new_n313));
  NAND4_X1  g0113(.A1(new_n312), .A2(new_n313), .A3(new_n309), .A4(new_n306), .ZN(new_n314));
  AOI21_X1  g0114(.A(new_n305), .B1(new_n311), .B2(new_n314), .ZN(new_n315));
  OAI21_X1  g0115(.A(new_n260), .B1(new_n220), .B2(new_n266), .ZN(new_n316));
  XOR2_X1   g0116(.A(new_n316), .B(KEYINPUT74), .Z(new_n317));
  INV_X1    g0117(.A(G238), .ZN(new_n318));
  OAI22_X1  g0118(.A1(new_n278), .A2(new_n318), .B1(new_n211), .B2(new_n277), .ZN(new_n319));
  AND3_X1   g0119(.A1(new_n268), .A2(new_n270), .A3(KEYINPUT72), .ZN(new_n320));
  AOI21_X1  g0120(.A(KEYINPUT72), .B1(new_n268), .B2(new_n270), .ZN(new_n321));
  NOR2_X1   g0121(.A1(new_n320), .A2(new_n321), .ZN(new_n322));
  NOR3_X1   g0122(.A1(new_n322), .A2(new_n210), .A3(G1698), .ZN(new_n323));
  OAI21_X1  g0123(.A(new_n281), .B1(new_n319), .B2(new_n323), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n317), .A2(new_n324), .ZN(new_n325));
  INV_X1    g0125(.A(G169), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n325), .A2(new_n326), .ZN(new_n327));
  INV_X1    g0127(.A(new_n295), .ZN(new_n328));
  AOI22_X1  g0128(.A1(new_n328), .A2(new_n298), .B1(G20), .B2(G77), .ZN(new_n329));
  XOR2_X1   g0129(.A(KEYINPUT15), .B(G87), .Z(new_n330));
  INV_X1    g0130(.A(new_n330), .ZN(new_n331));
  OAI21_X1  g0131(.A(new_n329), .B1(new_n331), .B2(new_n296), .ZN(new_n332));
  AOI22_X1  g0132(.A1(new_n332), .A2(new_n289), .B1(new_n219), .B2(new_n293), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n290), .A2(G77), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n333), .A2(new_n334), .ZN(new_n335));
  INV_X1    g0135(.A(KEYINPUT75), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n335), .A2(new_n336), .ZN(new_n337));
  NAND3_X1  g0137(.A1(new_n333), .A2(KEYINPUT75), .A3(new_n334), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n337), .A2(new_n338), .ZN(new_n339));
  OAI211_X1 g0139(.A(new_n327), .B(new_n339), .C1(G179), .C2(new_n325), .ZN(new_n340));
  INV_X1    g0140(.A(KEYINPUT76), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n325), .A2(G200), .ZN(new_n342));
  NAND3_X1  g0142(.A1(new_n317), .A2(G190), .A3(new_n324), .ZN(new_n343));
  NAND4_X1  g0143(.A1(new_n342), .A2(new_n337), .A3(new_n338), .A4(new_n343), .ZN(new_n344));
  AND3_X1   g0144(.A1(new_n340), .A2(new_n341), .A3(new_n344), .ZN(new_n345));
  AOI21_X1  g0145(.A(new_n341), .B1(new_n340), .B2(new_n344), .ZN(new_n346));
  OAI21_X1  g0146(.A(new_n315), .B1(new_n345), .B2(new_n346), .ZN(new_n347));
  OAI21_X1  g0147(.A(new_n231), .B1(new_n207), .B2(new_n209), .ZN(new_n348));
  AOI22_X1  g0148(.A1(new_n348), .A2(G20), .B1(G159), .B2(new_n298), .ZN(new_n349));
  OAI21_X1  g0149(.A(KEYINPUT82), .B1(new_n262), .B2(KEYINPUT3), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n350), .A2(new_n268), .ZN(new_n351));
  NAND3_X1  g0151(.A1(new_n262), .A2(KEYINPUT82), .A3(KEYINPUT3), .ZN(new_n352));
  AOI21_X1  g0152(.A(G20), .B1(new_n351), .B2(new_n352), .ZN(new_n353));
  INV_X1    g0153(.A(KEYINPUT7), .ZN(new_n354));
  OAI21_X1  g0154(.A(G68), .B1(new_n353), .B2(new_n354), .ZN(new_n355));
  AOI211_X1 g0155(.A(KEYINPUT7), .B(G20), .C1(new_n351), .C2(new_n352), .ZN(new_n356));
  OAI211_X1 g0156(.A(KEYINPUT16), .B(new_n349), .C1(new_n355), .C2(new_n356), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n348), .A2(G20), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n298), .A2(G159), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n358), .A2(new_n359), .ZN(new_n360));
  NAND3_X1  g0160(.A1(new_n271), .A2(KEYINPUT7), .A3(new_n228), .ZN(new_n361));
  NOR3_X1   g0161(.A1(new_n320), .A2(new_n321), .A3(G20), .ZN(new_n362));
  OAI21_X1  g0162(.A(new_n361), .B1(new_n362), .B2(KEYINPUT7), .ZN(new_n363));
  AOI21_X1  g0163(.A(new_n360), .B1(new_n363), .B2(new_n208), .ZN(new_n364));
  XNOR2_X1  g0164(.A(KEYINPUT83), .B(KEYINPUT16), .ZN(new_n365));
  OAI211_X1 g0165(.A(new_n289), .B(new_n357), .C1(new_n364), .C2(new_n365), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n295), .A2(new_n292), .ZN(new_n367));
  OAI21_X1  g0167(.A(new_n367), .B1(new_n290), .B2(new_n295), .ZN(new_n368));
  OAI21_X1  g0168(.A(new_n260), .B1(new_n210), .B2(new_n266), .ZN(new_n369));
  INV_X1    g0169(.A(G1698), .ZN(new_n370));
  NOR2_X1   g0170(.A1(new_n261), .A2(new_n370), .ZN(new_n371));
  INV_X1    g0171(.A(KEYINPUT82), .ZN(new_n372));
  AOI21_X1  g0172(.A(new_n372), .B1(new_n269), .B2(G33), .ZN(new_n373));
  NOR2_X1   g0173(.A1(new_n269), .A2(G33), .ZN(new_n374));
  OAI211_X1 g0174(.A(new_n352), .B(new_n371), .C1(new_n373), .C2(new_n374), .ZN(new_n375));
  INV_X1    g0175(.A(KEYINPUT84), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n375), .A2(new_n376), .ZN(new_n377));
  NAND2_X1  g0177(.A1(G33), .A2(G87), .ZN(new_n378));
  NAND4_X1  g0178(.A1(new_n351), .A2(G223), .A3(new_n370), .A4(new_n352), .ZN(new_n379));
  NAND4_X1  g0179(.A1(new_n351), .A2(KEYINPUT84), .A3(new_n352), .A4(new_n371), .ZN(new_n380));
  NAND4_X1  g0180(.A1(new_n377), .A2(new_n378), .A3(new_n379), .A4(new_n380), .ZN(new_n381));
  AOI21_X1  g0181(.A(new_n369), .B1(new_n381), .B2(new_n281), .ZN(new_n382));
  XNOR2_X1  g0182(.A(KEYINPUT86), .B(G190), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n382), .A2(new_n383), .ZN(new_n384));
  NAND2_X1  g0184(.A1(new_n381), .A2(new_n281), .ZN(new_n385));
  INV_X1    g0185(.A(new_n369), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n385), .A2(new_n386), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n387), .A2(G200), .ZN(new_n388));
  NAND4_X1  g0188(.A1(new_n366), .A2(new_n368), .A3(new_n384), .A4(new_n388), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n389), .A2(KEYINPUT17), .ZN(new_n390));
  INV_X1    g0190(.A(new_n368), .ZN(new_n391));
  OAI21_X1  g0191(.A(new_n352), .B1(new_n373), .B2(new_n374), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n392), .A2(new_n228), .ZN(new_n393));
  AOI21_X1  g0193(.A(new_n252), .B1(new_n393), .B2(KEYINPUT7), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n353), .A2(new_n354), .ZN(new_n395));
  AOI21_X1  g0195(.A(new_n360), .B1(new_n394), .B2(new_n395), .ZN(new_n396));
  AOI21_X1  g0196(.A(new_n302), .B1(new_n396), .B2(KEYINPUT16), .ZN(new_n397));
  INV_X1    g0197(.A(new_n361), .ZN(new_n398));
  NAND3_X1  g0198(.A1(new_n273), .A2(new_n228), .A3(new_n274), .ZN(new_n399));
  AOI21_X1  g0199(.A(new_n398), .B1(new_n399), .B2(new_n354), .ZN(new_n400));
  OAI21_X1  g0200(.A(new_n349), .B1(new_n400), .B2(new_n207), .ZN(new_n401));
  INV_X1    g0201(.A(new_n365), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n401), .A2(new_n402), .ZN(new_n403));
  AOI21_X1  g0203(.A(new_n391), .B1(new_n397), .B2(new_n403), .ZN(new_n404));
  INV_X1    g0204(.A(KEYINPUT17), .ZN(new_n405));
  NAND4_X1  g0205(.A1(new_n404), .A2(new_n405), .A3(new_n384), .A4(new_n388), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n390), .A2(new_n406), .ZN(new_n407));
  INV_X1    g0207(.A(KEYINPUT18), .ZN(new_n408));
  NOR2_X1   g0208(.A1(new_n382), .A2(new_n326), .ZN(new_n409));
  INV_X1    g0209(.A(G179), .ZN(new_n410));
  AOI211_X1 g0210(.A(new_n410), .B(new_n369), .C1(new_n381), .C2(new_n281), .ZN(new_n411));
  NOR2_X1   g0211(.A1(new_n409), .A2(new_n411), .ZN(new_n412));
  OAI21_X1  g0212(.A(new_n408), .B1(new_n404), .B2(new_n412), .ZN(new_n413));
  AOI21_X1  g0213(.A(KEYINPUT7), .B1(new_n322), .B2(new_n228), .ZN(new_n414));
  OAI21_X1  g0214(.A(new_n208), .B1(new_n414), .B2(new_n398), .ZN(new_n415));
  AOI21_X1  g0215(.A(new_n365), .B1(new_n415), .B2(new_n349), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n357), .A2(new_n289), .ZN(new_n417));
  OAI21_X1  g0217(.A(new_n368), .B1(new_n416), .B2(new_n417), .ZN(new_n418));
  INV_X1    g0218(.A(KEYINPUT85), .ZN(new_n419));
  NAND3_X1  g0219(.A1(new_n385), .A2(G179), .A3(new_n386), .ZN(new_n420));
  OAI21_X1  g0220(.A(new_n420), .B1(new_n326), .B2(new_n382), .ZN(new_n421));
  NAND4_X1  g0221(.A1(new_n418), .A2(new_n419), .A3(KEYINPUT18), .A4(new_n421), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n413), .A2(new_n422), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n387), .A2(G169), .ZN(new_n424));
  AOI22_X1  g0224(.A1(new_n366), .A2(new_n368), .B1(new_n424), .B2(new_n420), .ZN(new_n425));
  AOI21_X1  g0225(.A(new_n419), .B1(new_n425), .B2(KEYINPUT18), .ZN(new_n426));
  OAI21_X1  g0226(.A(new_n407), .B1(new_n423), .B2(new_n426), .ZN(new_n427));
  NOR2_X1   g0227(.A1(new_n208), .A2(new_n228), .ZN(new_n428));
  OAI22_X1  g0228(.A1(new_n299), .A2(new_n202), .B1(new_n296), .B2(new_n219), .ZN(new_n429));
  OAI21_X1  g0229(.A(new_n289), .B1(new_n428), .B2(new_n429), .ZN(new_n430));
  XNOR2_X1  g0230(.A(new_n430), .B(KEYINPUT11), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n290), .A2(G68), .ZN(new_n432));
  OAI21_X1  g0232(.A(KEYINPUT12), .B1(new_n208), .B2(new_n292), .ZN(new_n433));
  OR2_X1    g0233(.A1(KEYINPUT12), .A2(G68), .ZN(new_n434));
  OR3_X1    g0234(.A1(new_n292), .A2(new_n434), .A3(KEYINPUT79), .ZN(new_n435));
  OAI21_X1  g0235(.A(KEYINPUT79), .B1(new_n292), .B2(new_n434), .ZN(new_n436));
  NAND3_X1  g0236(.A1(new_n433), .A2(new_n435), .A3(new_n436), .ZN(new_n437));
  AND3_X1   g0237(.A1(new_n432), .A2(KEYINPUT80), .A3(new_n437), .ZN(new_n438));
  AOI21_X1  g0238(.A(KEYINPUT80), .B1(new_n432), .B2(new_n437), .ZN(new_n439));
  OAI21_X1  g0239(.A(new_n431), .B1(new_n438), .B2(new_n439), .ZN(new_n440));
  XNOR2_X1  g0240(.A(new_n440), .B(KEYINPUT81), .ZN(new_n441));
  AOI22_X1  g0241(.A1(new_n275), .A2(G226), .B1(G33), .B2(G97), .ZN(new_n442));
  NAND3_X1  g0242(.A1(new_n277), .A2(G232), .A3(G1698), .ZN(new_n443));
  AOI21_X1  g0243(.A(new_n264), .B1(new_n442), .B2(new_n443), .ZN(new_n444));
  INV_X1    g0244(.A(KEYINPUT77), .ZN(new_n445));
  OAI21_X1  g0245(.A(G238), .B1(new_n266), .B2(new_n445), .ZN(new_n446));
  AOI21_X1  g0246(.A(KEYINPUT77), .B1(new_n264), .B2(new_n265), .ZN(new_n447));
  OAI21_X1  g0247(.A(new_n260), .B1(new_n446), .B2(new_n447), .ZN(new_n448));
  OAI21_X1  g0248(.A(KEYINPUT13), .B1(new_n444), .B2(new_n448), .ZN(new_n449));
  NAND3_X1  g0249(.A1(new_n277), .A2(G226), .A3(new_n370), .ZN(new_n450));
  NAND2_X1  g0250(.A1(G33), .A2(G97), .ZN(new_n451));
  NAND3_X1  g0251(.A1(new_n443), .A2(new_n450), .A3(new_n451), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n452), .A2(new_n281), .ZN(new_n453));
  INV_X1    g0253(.A(KEYINPUT13), .ZN(new_n454));
  INV_X1    g0254(.A(new_n448), .ZN(new_n455));
  NAND3_X1  g0255(.A1(new_n453), .A2(new_n454), .A3(new_n455), .ZN(new_n456));
  NAND3_X1  g0256(.A1(new_n449), .A2(new_n456), .A3(G179), .ZN(new_n457));
  AOI21_X1  g0257(.A(new_n326), .B1(new_n449), .B2(new_n456), .ZN(new_n458));
  INV_X1    g0258(.A(KEYINPUT14), .ZN(new_n459));
  OAI21_X1  g0259(.A(new_n457), .B1(new_n458), .B2(new_n459), .ZN(new_n460));
  NOR3_X1   g0260(.A1(new_n444), .A2(KEYINPUT13), .A3(new_n448), .ZN(new_n461));
  AOI21_X1  g0261(.A(new_n454), .B1(new_n453), .B2(new_n455), .ZN(new_n462));
  OAI211_X1 g0262(.A(new_n459), .B(G169), .C1(new_n461), .C2(new_n462), .ZN(new_n463));
  INV_X1    g0263(.A(new_n463), .ZN(new_n464));
  OAI21_X1  g0264(.A(new_n441), .B1(new_n460), .B2(new_n464), .ZN(new_n465));
  INV_X1    g0265(.A(new_n465), .ZN(new_n466));
  NAND3_X1  g0266(.A1(new_n449), .A2(new_n456), .A3(G190), .ZN(new_n467));
  INV_X1    g0267(.A(KEYINPUT78), .ZN(new_n468));
  OR2_X1    g0268(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  INV_X1    g0269(.A(KEYINPUT81), .ZN(new_n470));
  XNOR2_X1  g0270(.A(new_n440), .B(new_n470), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n467), .A2(new_n468), .ZN(new_n472));
  OAI21_X1  g0272(.A(G200), .B1(new_n461), .B2(new_n462), .ZN(new_n473));
  NAND4_X1  g0273(.A1(new_n469), .A2(new_n471), .A3(new_n472), .A4(new_n473), .ZN(new_n474));
  INV_X1    g0274(.A(new_n474), .ZN(new_n475));
  NOR4_X1   g0275(.A1(new_n347), .A2(new_n427), .A3(new_n466), .A4(new_n475), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n293), .A2(new_n211), .ZN(new_n477));
  INV_X1    g0277(.A(KEYINPUT25), .ZN(new_n478));
  XNOR2_X1  g0278(.A(new_n477), .B(new_n478), .ZN(new_n479));
  OAI21_X1  g0279(.A(new_n292), .B1(G1), .B2(new_n262), .ZN(new_n480));
  NOR2_X1   g0280(.A1(new_n289), .A2(new_n480), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n481), .A2(G107), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n479), .A2(new_n482), .ZN(new_n483));
  NAND2_X1  g0283(.A1(KEYINPUT22), .A2(G87), .ZN(new_n484));
  INV_X1    g0284(.A(G116), .ZN(new_n485));
  OAI22_X1  g0285(.A1(new_n392), .A2(new_n484), .B1(new_n262), .B2(new_n485), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n486), .A2(new_n228), .ZN(new_n487));
  INV_X1    g0287(.A(KEYINPUT22), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n228), .A2(G87), .ZN(new_n489));
  OAI21_X1  g0289(.A(new_n488), .B1(new_n322), .B2(new_n489), .ZN(new_n490));
  NOR2_X1   g0290(.A1(new_n228), .A2(G107), .ZN(new_n491));
  XNOR2_X1  g0291(.A(new_n491), .B(KEYINPUT23), .ZN(new_n492));
  NAND3_X1  g0292(.A1(new_n487), .A2(new_n490), .A3(new_n492), .ZN(new_n493));
  INV_X1    g0293(.A(KEYINPUT24), .ZN(new_n494));
  AOI21_X1  g0294(.A(new_n302), .B1(new_n493), .B2(new_n494), .ZN(new_n495));
  NAND4_X1  g0295(.A1(new_n487), .A2(new_n490), .A3(KEYINPUT24), .A4(new_n492), .ZN(new_n496));
  AOI21_X1  g0296(.A(new_n483), .B1(new_n495), .B2(new_n496), .ZN(new_n497));
  INV_X1    g0297(.A(new_n352), .ZN(new_n498));
  AOI21_X1  g0298(.A(new_n498), .B1(new_n268), .B2(new_n350), .ZN(new_n499));
  INV_X1    g0299(.A(G257), .ZN(new_n500));
  NOR2_X1   g0300(.A1(new_n500), .A2(new_n370), .ZN(new_n501));
  AOI22_X1  g0301(.A1(new_n499), .A2(new_n501), .B1(G33), .B2(G294), .ZN(new_n502));
  NAND4_X1  g0302(.A1(new_n499), .A2(KEYINPUT92), .A3(G250), .A4(new_n370), .ZN(new_n503));
  NAND4_X1  g0303(.A1(new_n351), .A2(G250), .A3(new_n370), .A4(new_n352), .ZN(new_n504));
  INV_X1    g0304(.A(KEYINPUT92), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  NAND3_X1  g0306(.A1(new_n502), .A2(new_n503), .A3(new_n506), .ZN(new_n507));
  XNOR2_X1  g0307(.A(KEYINPUT5), .B(G41), .ZN(new_n508));
  INV_X1    g0308(.A(G45), .ZN(new_n509));
  NOR2_X1   g0309(.A1(new_n509), .A2(G1), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n508), .A2(new_n510), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n511), .A2(new_n264), .ZN(new_n512));
  INV_X1    g0312(.A(new_n512), .ZN(new_n513));
  AOI22_X1  g0313(.A1(new_n507), .A2(new_n281), .B1(G264), .B2(new_n513), .ZN(new_n514));
  INV_X1    g0314(.A(G190), .ZN(new_n515));
  NAND3_X1  g0315(.A1(new_n508), .A2(G274), .A3(new_n510), .ZN(new_n516));
  AND3_X1   g0316(.A1(new_n514), .A2(new_n515), .A3(new_n516), .ZN(new_n517));
  AOI21_X1  g0317(.A(G200), .B1(new_n514), .B2(new_n516), .ZN(new_n518));
  OAI21_X1  g0318(.A(new_n497), .B1(new_n517), .B2(new_n518), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n519), .A2(KEYINPUT94), .ZN(new_n520));
  INV_X1    g0320(.A(KEYINPUT94), .ZN(new_n521));
  OAI211_X1 g0321(.A(new_n521), .B(new_n497), .C1(new_n517), .C2(new_n518), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n520), .A2(new_n522), .ZN(new_n523));
  INV_X1    g0323(.A(KEYINPUT93), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n514), .A2(new_n516), .ZN(new_n525));
  NOR2_X1   g0325(.A1(new_n525), .A2(new_n410), .ZN(new_n526));
  AOI21_X1  g0326(.A(new_n326), .B1(new_n514), .B2(new_n516), .ZN(new_n527));
  OAI21_X1  g0327(.A(new_n524), .B1(new_n526), .B2(new_n527), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n525), .A2(G169), .ZN(new_n529));
  OAI211_X1 g0329(.A(new_n529), .B(KEYINPUT93), .C1(new_n410), .C2(new_n525), .ZN(new_n530));
  INV_X1    g0330(.A(new_n497), .ZN(new_n531));
  NAND3_X1  g0331(.A1(new_n528), .A2(new_n530), .A3(new_n531), .ZN(new_n532));
  AND2_X1   g0332(.A1(new_n523), .A2(new_n532), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n481), .A2(G97), .ZN(new_n534));
  INV_X1    g0334(.A(G97), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n293), .A2(new_n535), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n534), .A2(new_n536), .ZN(new_n537));
  NAND3_X1  g0337(.A1(new_n211), .A2(KEYINPUT6), .A3(G97), .ZN(new_n538));
  NOR2_X1   g0338(.A1(new_n535), .A2(new_n211), .ZN(new_n539));
  NOR2_X1   g0339(.A1(G97), .A2(G107), .ZN(new_n540));
  NOR2_X1   g0340(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  OAI21_X1  g0341(.A(new_n538), .B1(new_n541), .B2(KEYINPUT6), .ZN(new_n542));
  AOI22_X1  g0342(.A1(new_n542), .A2(G20), .B1(G77), .B2(new_n298), .ZN(new_n543));
  OAI21_X1  g0343(.A(new_n543), .B1(new_n400), .B2(new_n211), .ZN(new_n544));
  AOI21_X1  g0344(.A(new_n537), .B1(new_n544), .B2(new_n289), .ZN(new_n545));
  INV_X1    g0345(.A(new_n545), .ZN(new_n546));
  OAI21_X1  g0346(.A(new_n516), .B1(new_n512), .B2(new_n500), .ZN(new_n547));
  INV_X1    g0347(.A(KEYINPUT87), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  OAI211_X1 g0349(.A(KEYINPUT87), .B(new_n516), .C1(new_n512), .C2(new_n500), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  NAND4_X1  g0351(.A1(new_n351), .A2(G244), .A3(new_n370), .A4(new_n352), .ZN(new_n552));
  INV_X1    g0352(.A(KEYINPUT4), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n552), .A2(new_n553), .ZN(new_n554));
  NOR2_X1   g0354(.A1(new_n553), .A2(new_n220), .ZN(new_n555));
  OAI211_X1 g0355(.A(new_n370), .B(new_n555), .C1(new_n320), .C2(new_n321), .ZN(new_n556));
  OAI211_X1 g0356(.A(G250), .B(G1698), .C1(new_n320), .C2(new_n321), .ZN(new_n557));
  NAND2_X1  g0357(.A1(G33), .A2(G283), .ZN(new_n558));
  NAND4_X1  g0358(.A1(new_n554), .A2(new_n556), .A3(new_n557), .A4(new_n558), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n559), .A2(new_n281), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n551), .A2(new_n560), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n561), .A2(new_n326), .ZN(new_n562));
  AOI22_X1  g0362(.A1(new_n549), .A2(new_n550), .B1(new_n559), .B2(new_n281), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n563), .A2(new_n410), .ZN(new_n564));
  NAND3_X1  g0364(.A1(new_n546), .A2(new_n562), .A3(new_n564), .ZN(new_n565));
  NAND3_X1  g0365(.A1(new_n551), .A2(new_n560), .A3(G190), .ZN(new_n566));
  OAI211_X1 g0366(.A(new_n545), .B(new_n566), .C1(new_n307), .C2(new_n563), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n565), .A2(new_n567), .ZN(new_n568));
  INV_X1    g0368(.A(KEYINPUT21), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n481), .A2(G116), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n293), .A2(new_n485), .ZN(new_n571));
  INV_X1    g0371(.A(KEYINPUT90), .ZN(new_n572));
  XNOR2_X1  g0372(.A(new_n571), .B(new_n572), .ZN(new_n573));
  AOI21_X1  g0373(.A(G20), .B1(G33), .B2(G283), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n262), .A2(G97), .ZN(new_n575));
  AOI22_X1  g0375(.A1(new_n574), .A2(new_n575), .B1(G20), .B2(new_n485), .ZN(new_n576));
  AOI21_X1  g0376(.A(KEYINPUT20), .B1(new_n289), .B2(new_n576), .ZN(new_n577));
  AND2_X1   g0377(.A1(new_n577), .A2(KEYINPUT91), .ZN(new_n578));
  NAND3_X1  g0378(.A1(new_n289), .A2(new_n576), .A3(KEYINPUT20), .ZN(new_n579));
  OAI21_X1  g0379(.A(new_n579), .B1(new_n577), .B2(KEYINPUT91), .ZN(new_n580));
  OAI211_X1 g0380(.A(new_n570), .B(new_n573), .C1(new_n578), .C2(new_n580), .ZN(new_n581));
  INV_X1    g0381(.A(new_n581), .ZN(new_n582));
  NAND3_X1  g0382(.A1(new_n273), .A2(G303), .A3(new_n274), .ZN(new_n583));
  NOR2_X1   g0383(.A1(G257), .A2(G1698), .ZN(new_n584));
  AOI21_X1  g0384(.A(new_n584), .B1(new_n212), .B2(G1698), .ZN(new_n585));
  NAND3_X1  g0385(.A1(new_n351), .A2(new_n585), .A3(new_n352), .ZN(new_n586));
  AOI21_X1  g0386(.A(new_n264), .B1(new_n583), .B2(new_n586), .ZN(new_n587));
  INV_X1    g0387(.A(G270), .ZN(new_n588));
  OAI21_X1  g0388(.A(new_n516), .B1(new_n512), .B2(new_n588), .ZN(new_n589));
  OAI21_X1  g0389(.A(G169), .B1(new_n587), .B2(new_n589), .ZN(new_n590));
  OAI21_X1  g0390(.A(new_n569), .B1(new_n582), .B2(new_n590), .ZN(new_n591));
  OAI21_X1  g0391(.A(G200), .B1(new_n587), .B2(new_n589), .ZN(new_n592));
  NOR2_X1   g0392(.A1(new_n587), .A2(new_n589), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n593), .A2(new_n383), .ZN(new_n594));
  NAND3_X1  g0394(.A1(new_n582), .A2(new_n592), .A3(new_n594), .ZN(new_n595));
  INV_X1    g0395(.A(new_n590), .ZN(new_n596));
  NAND3_X1  g0396(.A1(new_n596), .A2(new_n581), .A3(KEYINPUT21), .ZN(new_n597));
  NOR3_X1   g0397(.A1(new_n587), .A2(new_n589), .A3(new_n410), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n581), .A2(new_n598), .ZN(new_n599));
  NAND4_X1  g0399(.A1(new_n591), .A2(new_n595), .A3(new_n597), .A4(new_n599), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n510), .A2(G274), .ZN(new_n601));
  OAI21_X1  g0401(.A(G250), .B1(new_n509), .B2(G1), .ZN(new_n602));
  OAI21_X1  g0402(.A(new_n601), .B1(new_n281), .B2(new_n602), .ZN(new_n603));
  NAND4_X1  g0403(.A1(new_n351), .A2(G238), .A3(new_n370), .A4(new_n352), .ZN(new_n604));
  NAND4_X1  g0404(.A1(new_n351), .A2(G244), .A3(G1698), .A4(new_n352), .ZN(new_n605));
  OAI211_X1 g0405(.A(new_n604), .B(new_n605), .C1(new_n262), .C2(new_n485), .ZN(new_n606));
  AOI21_X1  g0406(.A(new_n603), .B1(new_n606), .B2(new_n281), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n607), .A2(G190), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n608), .A2(KEYINPUT89), .ZN(new_n609));
  NOR2_X1   g0409(.A1(new_n330), .A2(new_n292), .ZN(new_n610));
  INV_X1    g0410(.A(G87), .ZN(new_n611));
  NOR3_X1   g0411(.A1(new_n289), .A2(new_n480), .A3(new_n611), .ZN(new_n612));
  INV_X1    g0412(.A(KEYINPUT19), .ZN(new_n613));
  OAI21_X1  g0413(.A(new_n228), .B1(new_n451), .B2(new_n613), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n540), .A2(new_n611), .ZN(new_n615));
  NAND3_X1  g0415(.A1(new_n228), .A2(G33), .A3(G97), .ZN(new_n616));
  AOI22_X1  g0416(.A1(new_n614), .A2(new_n615), .B1(new_n613), .B2(new_n616), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n228), .A2(G68), .ZN(new_n618));
  OAI21_X1  g0418(.A(new_n617), .B1(new_n392), .B2(new_n618), .ZN(new_n619));
  AOI21_X1  g0419(.A(new_n302), .B1(new_n619), .B2(KEYINPUT88), .ZN(new_n620));
  INV_X1    g0420(.A(KEYINPUT88), .ZN(new_n621));
  OAI211_X1 g0421(.A(new_n617), .B(new_n621), .C1(new_n392), .C2(new_n618), .ZN(new_n622));
  AOI211_X1 g0422(.A(new_n610), .B(new_n612), .C1(new_n620), .C2(new_n622), .ZN(new_n623));
  INV_X1    g0423(.A(KEYINPUT89), .ZN(new_n624));
  NAND3_X1  g0424(.A1(new_n607), .A2(new_n624), .A3(G190), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n606), .A2(new_n281), .ZN(new_n626));
  INV_X1    g0426(.A(new_n603), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n628), .A2(G200), .ZN(new_n629));
  NAND4_X1  g0429(.A1(new_n609), .A2(new_n623), .A3(new_n625), .A4(new_n629), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n628), .A2(new_n326), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n620), .A2(new_n622), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n481), .A2(new_n330), .ZN(new_n633));
  INV_X1    g0433(.A(new_n610), .ZN(new_n634));
  NAND3_X1  g0434(.A1(new_n632), .A2(new_n633), .A3(new_n634), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n607), .A2(new_n410), .ZN(new_n636));
  NAND3_X1  g0436(.A1(new_n631), .A2(new_n635), .A3(new_n636), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n630), .A2(new_n637), .ZN(new_n638));
  NOR3_X1   g0438(.A1(new_n568), .A2(new_n600), .A3(new_n638), .ZN(new_n639));
  AND3_X1   g0439(.A1(new_n476), .A2(new_n533), .A3(new_n639), .ZN(G372));
  INV_X1    g0440(.A(new_n565), .ZN(new_n641));
  INV_X1    g0441(.A(KEYINPUT26), .ZN(new_n642));
  NAND3_X1  g0442(.A1(new_n623), .A2(new_n629), .A3(new_n608), .ZN(new_n643));
  NAND3_X1  g0443(.A1(new_n643), .A2(new_n637), .A3(KEYINPUT95), .ZN(new_n644));
  INV_X1    g0444(.A(new_n644), .ZN(new_n645));
  AOI21_X1  g0445(.A(KEYINPUT95), .B1(new_n643), .B2(new_n637), .ZN(new_n646));
  OAI211_X1 g0446(.A(new_n641), .B(new_n642), .C1(new_n645), .C2(new_n646), .ZN(new_n647));
  INV_X1    g0447(.A(new_n637), .ZN(new_n648));
  AOI21_X1  g0448(.A(new_n545), .B1(new_n326), .B2(new_n561), .ZN(new_n649));
  NAND4_X1  g0449(.A1(new_n630), .A2(new_n649), .A3(new_n564), .A4(new_n637), .ZN(new_n650));
  AOI21_X1  g0450(.A(new_n648), .B1(new_n650), .B2(KEYINPUT26), .ZN(new_n651));
  AND2_X1   g0451(.A1(new_n647), .A2(new_n651), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n643), .A2(new_n637), .ZN(new_n653));
  INV_X1    g0453(.A(KEYINPUT95), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  AOI21_X1  g0455(.A(new_n568), .B1(new_n655), .B2(new_n644), .ZN(new_n656));
  NAND3_X1  g0456(.A1(new_n591), .A2(new_n597), .A3(new_n599), .ZN(new_n657));
  INV_X1    g0457(.A(KEYINPUT96), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  NAND4_X1  g0459(.A1(new_n591), .A2(new_n597), .A3(new_n599), .A4(KEYINPUT96), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  OAI21_X1  g0461(.A(new_n531), .B1(new_n526), .B2(new_n527), .ZN(new_n662));
  INV_X1    g0462(.A(new_n662), .ZN(new_n663));
  OAI211_X1 g0463(.A(new_n656), .B(new_n523), .C1(new_n661), .C2(new_n663), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n652), .A2(new_n664), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n476), .A2(new_n665), .ZN(new_n666));
  NAND3_X1  g0466(.A1(new_n418), .A2(KEYINPUT18), .A3(new_n421), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n413), .A2(new_n667), .ZN(new_n668));
  AND2_X1   g0468(.A1(new_n465), .A2(new_n340), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n474), .A2(new_n407), .ZN(new_n670));
  OAI21_X1  g0470(.A(new_n668), .B1(new_n669), .B2(new_n670), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n311), .A2(new_n314), .ZN(new_n672));
  AOI21_X1  g0472(.A(new_n305), .B1(new_n671), .B2(new_n672), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n666), .A2(new_n673), .ZN(G369));
  INV_X1    g0474(.A(G13), .ZN(new_n675));
  NOR2_X1   g0475(.A1(new_n675), .A2(G20), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n676), .A2(new_n258), .ZN(new_n677));
  OR2_X1    g0477(.A1(new_n677), .A2(KEYINPUT27), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n677), .A2(KEYINPUT27), .ZN(new_n679));
  NAND3_X1  g0479(.A1(new_n678), .A2(G213), .A3(new_n679), .ZN(new_n680));
  INV_X1    g0480(.A(G343), .ZN(new_n681));
  NOR2_X1   g0481(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n531), .A2(new_n682), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n533), .A2(new_n683), .ZN(new_n684));
  INV_X1    g0484(.A(KEYINPUT97), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  NAND3_X1  g0486(.A1(new_n533), .A2(KEYINPUT97), .A3(new_n683), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  INV_X1    g0488(.A(new_n682), .ZN(new_n689));
  OR2_X1    g0489(.A1(new_n532), .A2(new_n689), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n688), .A2(new_n690), .ZN(new_n691));
  INV_X1    g0491(.A(new_n691), .ZN(new_n692));
  NOR2_X1   g0492(.A1(new_n582), .A2(new_n689), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n661), .A2(new_n693), .ZN(new_n694));
  OAI21_X1  g0494(.A(new_n694), .B1(new_n600), .B2(new_n693), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n695), .A2(G330), .ZN(new_n696));
  NOR2_X1   g0496(.A1(new_n692), .A2(new_n696), .ZN(new_n697));
  INV_X1    g0497(.A(new_n657), .ZN(new_n698));
  NOR2_X1   g0498(.A1(new_n698), .A2(new_n682), .ZN(new_n699));
  NAND3_X1  g0499(.A1(new_n686), .A2(new_n687), .A3(new_n699), .ZN(new_n700));
  NAND2_X1  g0500(.A1(new_n663), .A2(new_n689), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  OR2_X1    g0502(.A1(new_n697), .A2(new_n702), .ZN(G399));
  INV_X1    g0503(.A(new_n224), .ZN(new_n704));
  OR3_X1    g0504(.A1(new_n704), .A2(KEYINPUT98), .A3(G41), .ZN(new_n705));
  OAI21_X1  g0505(.A(KEYINPUT98), .B1(new_n704), .B2(G41), .ZN(new_n706));
  NAND2_X1  g0506(.A1(new_n705), .A2(new_n706), .ZN(new_n707));
  INV_X1    g0507(.A(new_n707), .ZN(new_n708));
  NOR2_X1   g0508(.A1(new_n615), .A2(G116), .ZN(new_n709));
  INV_X1    g0509(.A(new_n709), .ZN(new_n710));
  NOR3_X1   g0510(.A1(new_n708), .A2(new_n258), .A3(new_n710), .ZN(new_n711));
  AOI21_X1  g0511(.A(new_n711), .B1(new_n233), .B2(new_n708), .ZN(new_n712));
  XOR2_X1   g0512(.A(new_n712), .B(KEYINPUT28), .Z(new_n713));
  AOI21_X1  g0513(.A(new_n682), .B1(new_n652), .B2(new_n664), .ZN(new_n714));
  NOR2_X1   g0514(.A1(new_n714), .A2(KEYINPUT29), .ZN(new_n715));
  AOI21_X1  g0515(.A(new_n565), .B1(new_n655), .B2(new_n644), .ZN(new_n716));
  NOR2_X1   g0516(.A1(new_n716), .A2(new_n642), .ZN(new_n717));
  OAI21_X1  g0517(.A(new_n637), .B1(new_n650), .B2(KEYINPUT26), .ZN(new_n718));
  NOR2_X1   g0518(.A1(new_n717), .A2(new_n718), .ZN(new_n719));
  NAND2_X1  g0519(.A1(new_n532), .A2(new_n698), .ZN(new_n720));
  NAND3_X1  g0520(.A1(new_n720), .A2(new_n523), .A3(new_n656), .ZN(new_n721));
  AOI21_X1  g0521(.A(new_n682), .B1(new_n719), .B2(new_n721), .ZN(new_n722));
  AOI21_X1  g0522(.A(new_n715), .B1(KEYINPUT29), .B2(new_n722), .ZN(new_n723));
  INV_X1    g0523(.A(G330), .ZN(new_n724));
  NAND4_X1  g0524(.A1(new_n639), .A2(new_n523), .A3(new_n532), .A4(new_n689), .ZN(new_n725));
  INV_X1    g0525(.A(KEYINPUT30), .ZN(new_n726));
  NAND2_X1  g0526(.A1(new_n507), .A2(new_n281), .ZN(new_n727));
  NAND2_X1  g0527(.A1(new_n513), .A2(G264), .ZN(new_n728));
  NAND4_X1  g0528(.A1(new_n727), .A2(new_n598), .A3(new_n728), .A4(new_n607), .ZN(new_n729));
  OAI21_X1  g0529(.A(new_n726), .B1(new_n729), .B2(new_n561), .ZN(new_n730));
  AND2_X1   g0530(.A1(new_n598), .A2(new_n607), .ZN(new_n731));
  NAND4_X1  g0531(.A1(new_n731), .A2(KEYINPUT30), .A3(new_n514), .A4(new_n563), .ZN(new_n732));
  NOR3_X1   g0532(.A1(new_n607), .A2(new_n593), .A3(G179), .ZN(new_n733));
  NAND3_X1  g0533(.A1(new_n525), .A2(new_n733), .A3(new_n561), .ZN(new_n734));
  NAND3_X1  g0534(.A1(new_n730), .A2(new_n732), .A3(new_n734), .ZN(new_n735));
  NAND2_X1  g0535(.A1(new_n735), .A2(new_n682), .ZN(new_n736));
  NAND2_X1  g0536(.A1(new_n736), .A2(KEYINPUT31), .ZN(new_n737));
  INV_X1    g0537(.A(KEYINPUT31), .ZN(new_n738));
  NAND3_X1  g0538(.A1(new_n735), .A2(new_n738), .A3(new_n682), .ZN(new_n739));
  NAND2_X1  g0539(.A1(new_n737), .A2(new_n739), .ZN(new_n740));
  AOI21_X1  g0540(.A(new_n724), .B1(new_n725), .B2(new_n740), .ZN(new_n741));
  NOR2_X1   g0541(.A1(new_n723), .A2(new_n741), .ZN(new_n742));
  OAI21_X1  g0542(.A(new_n713), .B1(new_n742), .B2(G1), .ZN(G364));
  INV_X1    g0543(.A(new_n696), .ZN(new_n744));
  AOI21_X1  g0544(.A(new_n258), .B1(new_n676), .B2(G45), .ZN(new_n745));
  INV_X1    g0545(.A(new_n745), .ZN(new_n746));
  NOR2_X1   g0546(.A1(new_n708), .A2(new_n746), .ZN(new_n747));
  NOR2_X1   g0547(.A1(new_n744), .A2(new_n747), .ZN(new_n748));
  OAI21_X1  g0548(.A(new_n748), .B1(G330), .B2(new_n695), .ZN(new_n749));
  INV_X1    g0549(.A(new_n747), .ZN(new_n750));
  NAND3_X1  g0550(.A1(new_n277), .A2(G355), .A3(new_n224), .ZN(new_n751));
  NOR2_X1   g0551(.A1(new_n499), .A2(new_n704), .ZN(new_n752));
  OAI21_X1  g0552(.A(new_n752), .B1(G45), .B2(new_n232), .ZN(new_n753));
  NOR2_X1   g0553(.A1(new_n256), .A2(new_n509), .ZN(new_n754));
  OAI221_X1 g0554(.A(new_n751), .B1(G116), .B2(new_n224), .C1(new_n753), .C2(new_n754), .ZN(new_n755));
  NOR2_X1   g0555(.A1(G13), .A2(G33), .ZN(new_n756));
  INV_X1    g0556(.A(new_n756), .ZN(new_n757));
  NOR2_X1   g0557(.A1(new_n757), .A2(G20), .ZN(new_n758));
  AOI21_X1  g0558(.A(new_n227), .B1(G20), .B2(new_n326), .ZN(new_n759));
  NOR2_X1   g0559(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  AOI21_X1  g0560(.A(new_n750), .B1(new_n755), .B2(new_n760), .ZN(new_n761));
  INV_X1    g0561(.A(new_n759), .ZN(new_n762));
  NOR3_X1   g0562(.A1(new_n515), .A2(G179), .A3(G200), .ZN(new_n763));
  NOR2_X1   g0563(.A1(new_n763), .A2(new_n228), .ZN(new_n764));
  INV_X1    g0564(.A(new_n764), .ZN(new_n765));
  NAND2_X1  g0565(.A1(new_n765), .A2(G97), .ZN(new_n766));
  NOR3_X1   g0566(.A1(new_n228), .A2(new_n410), .A3(G200), .ZN(new_n767));
  AND2_X1   g0567(.A1(new_n383), .A2(new_n767), .ZN(new_n768));
  INV_X1    g0568(.A(new_n768), .ZN(new_n769));
  OAI211_X1 g0569(.A(new_n766), .B(new_n277), .C1(new_n769), .C2(new_n209), .ZN(new_n770));
  NOR2_X1   g0570(.A1(new_n228), .A2(G190), .ZN(new_n771));
  NOR2_X1   g0571(.A1(new_n307), .A2(G179), .ZN(new_n772));
  NAND2_X1  g0572(.A1(new_n771), .A2(new_n772), .ZN(new_n773));
  INV_X1    g0573(.A(new_n773), .ZN(new_n774));
  NOR4_X1   g0574(.A1(new_n228), .A2(new_n410), .A3(new_n307), .A4(G190), .ZN(new_n775));
  AOI22_X1  g0575(.A1(new_n774), .A2(G107), .B1(new_n775), .B2(G68), .ZN(new_n776));
  NAND3_X1  g0576(.A1(new_n772), .A2(G20), .A3(G190), .ZN(new_n777));
  OAI21_X1  g0577(.A(new_n776), .B1(new_n611), .B2(new_n777), .ZN(new_n778));
  INV_X1    g0578(.A(KEYINPUT32), .ZN(new_n779));
  NAND3_X1  g0579(.A1(new_n771), .A2(new_n410), .A3(new_n307), .ZN(new_n780));
  INV_X1    g0580(.A(G159), .ZN(new_n781));
  OAI21_X1  g0581(.A(new_n779), .B1(new_n780), .B2(new_n781), .ZN(new_n782));
  INV_X1    g0582(.A(new_n780), .ZN(new_n783));
  NAND3_X1  g0583(.A1(new_n783), .A2(KEYINPUT32), .A3(G159), .ZN(new_n784));
  AOI211_X1 g0584(.A(new_n770), .B(new_n778), .C1(new_n782), .C2(new_n784), .ZN(new_n785));
  NAND2_X1  g0585(.A1(new_n767), .A2(new_n515), .ZN(new_n786));
  INV_X1    g0586(.A(new_n786), .ZN(new_n787));
  OR2_X1    g0587(.A1(new_n787), .A2(KEYINPUT99), .ZN(new_n788));
  NAND2_X1  g0588(.A1(new_n787), .A2(KEYINPUT99), .ZN(new_n789));
  NAND2_X1  g0589(.A1(new_n788), .A2(new_n789), .ZN(new_n790));
  INV_X1    g0590(.A(new_n790), .ZN(new_n791));
  NAND4_X1  g0591(.A1(new_n383), .A2(G20), .A3(G179), .A4(G200), .ZN(new_n792));
  AND2_X1   g0592(.A1(new_n792), .A2(KEYINPUT100), .ZN(new_n793));
  NOR2_X1   g0593(.A1(new_n792), .A2(KEYINPUT100), .ZN(new_n794));
  NOR2_X1   g0594(.A1(new_n793), .A2(new_n794), .ZN(new_n795));
  INV_X1    g0595(.A(new_n795), .ZN(new_n796));
  AOI22_X1  g0596(.A1(G77), .A2(new_n791), .B1(new_n796), .B2(G50), .ZN(new_n797));
  XNOR2_X1  g0597(.A(KEYINPUT101), .B(G326), .ZN(new_n798));
  NAND2_X1  g0598(.A1(new_n796), .A2(new_n798), .ZN(new_n799));
  INV_X1    g0599(.A(G322), .ZN(new_n800));
  OAI21_X1  g0600(.A(new_n322), .B1(new_n769), .B2(new_n800), .ZN(new_n801));
  INV_X1    g0601(.A(new_n775), .ZN(new_n802));
  XOR2_X1   g0602(.A(KEYINPUT33), .B(G317), .Z(new_n803));
  INV_X1    g0603(.A(G329), .ZN(new_n804));
  OAI22_X1  g0604(.A1(new_n802), .A2(new_n803), .B1(new_n804), .B2(new_n780), .ZN(new_n805));
  INV_X1    g0605(.A(G303), .ZN(new_n806));
  INV_X1    g0606(.A(G283), .ZN(new_n807));
  OAI22_X1  g0607(.A1(new_n777), .A2(new_n806), .B1(new_n773), .B2(new_n807), .ZN(new_n808));
  INV_X1    g0608(.A(G311), .ZN(new_n809));
  INV_X1    g0609(.A(G294), .ZN(new_n810));
  OAI22_X1  g0610(.A1(new_n786), .A2(new_n809), .B1(new_n764), .B2(new_n810), .ZN(new_n811));
  NOR4_X1   g0611(.A1(new_n801), .A2(new_n805), .A3(new_n808), .A4(new_n811), .ZN(new_n812));
  AOI22_X1  g0612(.A1(new_n785), .A2(new_n797), .B1(new_n799), .B2(new_n812), .ZN(new_n813));
  INV_X1    g0613(.A(new_n758), .ZN(new_n814));
  OAI221_X1 g0614(.A(new_n761), .B1(new_n762), .B2(new_n813), .C1(new_n695), .C2(new_n814), .ZN(new_n815));
  NAND2_X1  g0615(.A1(new_n749), .A2(new_n815), .ZN(G396));
  NAND2_X1  g0616(.A1(new_n339), .A2(new_n682), .ZN(new_n817));
  NAND2_X1  g0617(.A1(new_n344), .A2(new_n817), .ZN(new_n818));
  NAND2_X1  g0618(.A1(new_n818), .A2(new_n340), .ZN(new_n819));
  OR2_X1    g0619(.A1(new_n340), .A2(new_n682), .ZN(new_n820));
  AND2_X1   g0620(.A1(new_n819), .A2(new_n820), .ZN(new_n821));
  XNOR2_X1  g0621(.A(new_n714), .B(new_n821), .ZN(new_n822));
  INV_X1    g0622(.A(new_n741), .ZN(new_n823));
  AOI21_X1  g0623(.A(new_n747), .B1(new_n822), .B2(new_n823), .ZN(new_n824));
  OAI21_X1  g0624(.A(new_n824), .B1(new_n823), .B2(new_n822), .ZN(new_n825));
  NOR2_X1   g0625(.A1(new_n759), .A2(new_n756), .ZN(new_n826));
  AOI21_X1  g0626(.A(new_n750), .B1(new_n219), .B2(new_n826), .ZN(new_n827));
  OAI22_X1  g0627(.A1(new_n790), .A2(new_n485), .B1(new_n795), .B2(new_n806), .ZN(new_n828));
  OAI22_X1  g0628(.A1(new_n777), .A2(new_n211), .B1(new_n780), .B2(new_n809), .ZN(new_n829));
  OAI22_X1  g0629(.A1(new_n802), .A2(new_n807), .B1(new_n773), .B2(new_n611), .ZN(new_n830));
  OAI211_X1 g0630(.A(new_n766), .B(new_n322), .C1(new_n769), .C2(new_n810), .ZN(new_n831));
  NOR4_X1   g0631(.A1(new_n828), .A2(new_n829), .A3(new_n830), .A4(new_n831), .ZN(new_n832));
  NAND2_X1  g0632(.A1(new_n783), .A2(G132), .ZN(new_n833));
  OAI221_X1 g0633(.A(new_n833), .B1(new_n202), .B2(new_n777), .C1(new_n252), .C2(new_n773), .ZN(new_n834));
  OAI21_X1  g0634(.A(new_n499), .B1(new_n209), .B2(new_n764), .ZN(new_n835));
  AOI22_X1  g0635(.A1(new_n768), .A2(G143), .B1(G150), .B2(new_n775), .ZN(new_n836));
  INV_X1    g0636(.A(G137), .ZN(new_n837));
  OAI221_X1 g0637(.A(new_n836), .B1(new_n795), .B2(new_n837), .C1(new_n781), .C2(new_n790), .ZN(new_n838));
  INV_X1    g0638(.A(KEYINPUT34), .ZN(new_n839));
  AOI211_X1 g0639(.A(new_n834), .B(new_n835), .C1(new_n838), .C2(new_n839), .ZN(new_n840));
  OR2_X1    g0640(.A1(new_n838), .A2(new_n839), .ZN(new_n841));
  AOI21_X1  g0641(.A(new_n832), .B1(new_n840), .B2(new_n841), .ZN(new_n842));
  OAI221_X1 g0642(.A(new_n827), .B1(new_n762), .B2(new_n842), .C1(new_n821), .C2(new_n757), .ZN(new_n843));
  NAND2_X1  g0643(.A1(new_n825), .A2(new_n843), .ZN(G384));
  AOI211_X1 g0644(.A(new_n219), .B(new_n232), .C1(new_n208), .C2(G58), .ZN(new_n845));
  XOR2_X1   g0645(.A(new_n251), .B(KEYINPUT103), .Z(new_n846));
  OAI211_X1 g0646(.A(G1), .B(new_n675), .C1(new_n845), .C2(new_n846), .ZN(new_n847));
  OAI211_X1 g0647(.A(new_n230), .B(G116), .C1(new_n542), .C2(KEYINPUT35), .ZN(new_n848));
  AOI21_X1  g0648(.A(new_n848), .B1(KEYINPUT35), .B2(new_n542), .ZN(new_n849));
  XOR2_X1   g0649(.A(new_n849), .B(KEYINPUT102), .Z(new_n850));
  INV_X1    g0650(.A(KEYINPUT36), .ZN(new_n851));
  OAI21_X1  g0651(.A(new_n847), .B1(new_n850), .B2(new_n851), .ZN(new_n852));
  AOI21_X1  g0652(.A(new_n852), .B1(new_n851), .B2(new_n850), .ZN(new_n853));
  NAND2_X1  g0653(.A1(new_n725), .A2(new_n740), .ZN(new_n854));
  NAND2_X1  g0654(.A1(new_n441), .A2(new_n682), .ZN(new_n855));
  NAND3_X1  g0655(.A1(new_n465), .A2(new_n474), .A3(new_n855), .ZN(new_n856));
  OAI211_X1 g0656(.A(new_n441), .B(new_n682), .C1(new_n460), .C2(new_n464), .ZN(new_n857));
  NAND2_X1  g0657(.A1(new_n856), .A2(new_n857), .ZN(new_n858));
  AND3_X1   g0658(.A1(new_n854), .A2(new_n821), .A3(new_n858), .ZN(new_n859));
  INV_X1    g0659(.A(KEYINPUT38), .ZN(new_n860));
  NAND2_X1  g0660(.A1(new_n393), .A2(KEYINPUT7), .ZN(new_n861));
  NAND3_X1  g0661(.A1(new_n861), .A2(G68), .A3(new_n395), .ZN(new_n862));
  AOI21_X1  g0662(.A(new_n365), .B1(new_n862), .B2(new_n349), .ZN(new_n863));
  OAI21_X1  g0663(.A(new_n368), .B1(new_n417), .B2(new_n863), .ZN(new_n864));
  NAND2_X1  g0664(.A1(new_n864), .A2(KEYINPUT104), .ZN(new_n865));
  INV_X1    g0665(.A(new_n680), .ZN(new_n866));
  INV_X1    g0666(.A(KEYINPUT104), .ZN(new_n867));
  OAI211_X1 g0667(.A(new_n368), .B(new_n867), .C1(new_n417), .C2(new_n863), .ZN(new_n868));
  NAND3_X1  g0668(.A1(new_n865), .A2(new_n866), .A3(new_n868), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n667), .A2(KEYINPUT85), .ZN(new_n870));
  NAND3_X1  g0670(.A1(new_n870), .A2(new_n422), .A3(new_n413), .ZN(new_n871));
  AOI21_X1  g0671(.A(new_n869), .B1(new_n871), .B2(new_n407), .ZN(new_n872));
  OAI211_X1 g0672(.A(new_n420), .B(new_n680), .C1(new_n326), .C2(new_n382), .ZN(new_n873));
  NAND2_X1  g0673(.A1(new_n418), .A2(new_n873), .ZN(new_n874));
  INV_X1    g0674(.A(KEYINPUT37), .ZN(new_n875));
  NAND3_X1  g0675(.A1(new_n874), .A2(new_n875), .A3(new_n389), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n876), .A2(KEYINPUT105), .ZN(new_n877));
  INV_X1    g0677(.A(KEYINPUT105), .ZN(new_n878));
  NAND4_X1  g0678(.A1(new_n874), .A2(new_n389), .A3(new_n878), .A4(new_n875), .ZN(new_n879));
  NAND3_X1  g0679(.A1(new_n865), .A2(new_n873), .A3(new_n868), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n880), .A2(new_n389), .ZN(new_n881));
  AOI22_X1  g0681(.A1(new_n877), .A2(new_n879), .B1(new_n881), .B2(KEYINPUT37), .ZN(new_n882));
  OAI21_X1  g0682(.A(new_n860), .B1(new_n872), .B2(new_n882), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n877), .A2(new_n879), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n881), .A2(KEYINPUT37), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n884), .A2(new_n885), .ZN(new_n886));
  INV_X1    g0686(.A(new_n869), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n427), .A2(new_n887), .ZN(new_n888));
  NAND3_X1  g0688(.A1(new_n886), .A2(new_n888), .A3(KEYINPUT38), .ZN(new_n889));
  NAND3_X1  g0689(.A1(new_n883), .A2(new_n889), .A3(KEYINPUT106), .ZN(new_n890));
  INV_X1    g0690(.A(KEYINPUT106), .ZN(new_n891));
  OAI211_X1 g0691(.A(new_n891), .B(new_n860), .C1(new_n872), .C2(new_n882), .ZN(new_n892));
  NAND3_X1  g0692(.A1(new_n859), .A2(new_n890), .A3(new_n892), .ZN(new_n893));
  INV_X1    g0693(.A(KEYINPUT40), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  AOI21_X1  g0695(.A(new_n875), .B1(new_n874), .B2(new_n389), .ZN(new_n896));
  AOI21_X1  g0696(.A(new_n896), .B1(new_n877), .B2(new_n879), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n418), .A2(new_n866), .ZN(new_n898));
  AOI21_X1  g0698(.A(new_n898), .B1(new_n407), .B2(new_n668), .ZN(new_n899));
  OAI21_X1  g0699(.A(new_n860), .B1(new_n897), .B2(new_n899), .ZN(new_n900));
  AOI21_X1  g0700(.A(new_n894), .B1(new_n889), .B2(new_n900), .ZN(new_n901));
  NAND3_X1  g0701(.A1(new_n901), .A2(new_n859), .A3(KEYINPUT107), .ZN(new_n902));
  INV_X1    g0702(.A(new_n902), .ZN(new_n903));
  AOI21_X1  g0703(.A(KEYINPUT107), .B1(new_n901), .B2(new_n859), .ZN(new_n904));
  OAI211_X1 g0704(.A(new_n895), .B(G330), .C1(new_n903), .C2(new_n904), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n476), .A2(new_n741), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n905), .A2(new_n906), .ZN(new_n907));
  INV_X1    g0707(.A(new_n904), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n908), .A2(new_n902), .ZN(new_n909));
  NAND4_X1  g0709(.A1(new_n909), .A2(new_n476), .A3(new_n854), .A4(new_n895), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n907), .A2(new_n910), .ZN(new_n911));
  INV_X1    g0711(.A(new_n721), .ZN(new_n912));
  OR2_X1    g0712(.A1(new_n650), .A2(KEYINPUT26), .ZN(new_n913));
  OAI211_X1 g0713(.A(new_n913), .B(new_n637), .C1(new_n642), .C2(new_n716), .ZN(new_n914));
  OAI211_X1 g0714(.A(KEYINPUT29), .B(new_n689), .C1(new_n912), .C2(new_n914), .ZN(new_n915));
  OAI211_X1 g0715(.A(new_n915), .B(new_n476), .C1(KEYINPUT29), .C2(new_n714), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n916), .A2(new_n673), .ZN(new_n917));
  XOR2_X1   g0717(.A(new_n911), .B(new_n917), .Z(new_n918));
  NAND3_X1  g0718(.A1(new_n413), .A2(new_n667), .A3(new_n680), .ZN(new_n919));
  NAND3_X1  g0719(.A1(new_n665), .A2(new_n689), .A3(new_n821), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n920), .A2(new_n820), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n921), .A2(new_n858), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n890), .A2(new_n892), .ZN(new_n923));
  OAI21_X1  g0723(.A(new_n919), .B1(new_n922), .B2(new_n923), .ZN(new_n924));
  NOR2_X1   g0724(.A1(new_n465), .A2(new_n682), .ZN(new_n925));
  AOI21_X1  g0725(.A(KEYINPUT39), .B1(new_n889), .B2(new_n900), .ZN(new_n926));
  AOI21_X1  g0726(.A(new_n926), .B1(new_n923), .B2(KEYINPUT39), .ZN(new_n927));
  AOI21_X1  g0727(.A(new_n924), .B1(new_n925), .B2(new_n927), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n918), .A2(new_n928), .ZN(new_n929));
  OAI21_X1  g0729(.A(new_n929), .B1(new_n258), .B2(new_n676), .ZN(new_n930));
  NOR2_X1   g0730(.A1(new_n918), .A2(new_n928), .ZN(new_n931));
  OAI21_X1  g0731(.A(new_n853), .B1(new_n930), .B2(new_n931), .ZN(G367));
  OR2_X1    g0732(.A1(new_n623), .A2(new_n689), .ZN(new_n933));
  OAI21_X1  g0733(.A(new_n933), .B1(new_n645), .B2(new_n646), .ZN(new_n934));
  OR2_X1    g0734(.A1(new_n933), .A2(new_n637), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n934), .A2(new_n935), .ZN(new_n936));
  NOR2_X1   g0736(.A1(new_n936), .A2(KEYINPUT43), .ZN(new_n937));
  INV_X1    g0737(.A(KEYINPUT108), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n641), .A2(new_n682), .ZN(new_n939));
  OAI211_X1 g0739(.A(new_n565), .B(new_n567), .C1(new_n545), .C2(new_n689), .ZN(new_n940));
  NAND2_X1  g0740(.A1(new_n939), .A2(new_n940), .ZN(new_n941));
  AOI21_X1  g0741(.A(new_n938), .B1(new_n697), .B2(new_n941), .ZN(new_n942));
  INV_X1    g0742(.A(new_n942), .ZN(new_n943));
  NAND3_X1  g0743(.A1(new_n697), .A2(new_n938), .A3(new_n941), .ZN(new_n944));
  AOI21_X1  g0744(.A(new_n937), .B1(new_n943), .B2(new_n944), .ZN(new_n945));
  INV_X1    g0745(.A(new_n945), .ZN(new_n946));
  INV_X1    g0746(.A(new_n941), .ZN(new_n947));
  NOR2_X1   g0747(.A1(new_n700), .A2(new_n947), .ZN(new_n948));
  INV_X1    g0748(.A(KEYINPUT42), .ZN(new_n949));
  NOR2_X1   g0749(.A1(new_n948), .A2(new_n949), .ZN(new_n950));
  OAI21_X1  g0750(.A(new_n565), .B1(new_n532), .B2(new_n940), .ZN(new_n951));
  AOI21_X1  g0751(.A(new_n950), .B1(new_n689), .B2(new_n951), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n948), .A2(new_n949), .ZN(new_n953));
  NAND2_X1  g0753(.A1(new_n952), .A2(new_n953), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n936), .A2(KEYINPUT43), .ZN(new_n955));
  NAND2_X1  g0755(.A1(new_n954), .A2(new_n955), .ZN(new_n956));
  INV_X1    g0756(.A(new_n956), .ZN(new_n957));
  NAND3_X1  g0757(.A1(new_n943), .A2(new_n937), .A3(new_n944), .ZN(new_n958));
  NAND3_X1  g0758(.A1(new_n946), .A2(new_n957), .A3(new_n958), .ZN(new_n959));
  INV_X1    g0759(.A(new_n958), .ZN(new_n960));
  OAI21_X1  g0760(.A(new_n956), .B1(new_n960), .B2(new_n945), .ZN(new_n961));
  XNOR2_X1  g0761(.A(new_n707), .B(KEYINPUT41), .ZN(new_n962));
  NAND3_X1  g0762(.A1(new_n700), .A2(new_n701), .A3(new_n941), .ZN(new_n963));
  INV_X1    g0763(.A(KEYINPUT45), .ZN(new_n964));
  XNOR2_X1  g0764(.A(new_n963), .B(new_n964), .ZN(new_n965));
  AOI21_X1  g0765(.A(KEYINPUT44), .B1(new_n702), .B2(new_n947), .ZN(new_n966));
  NAND2_X1  g0766(.A1(new_n702), .A2(new_n947), .ZN(new_n967));
  INV_X1    g0767(.A(KEYINPUT44), .ZN(new_n968));
  NOR2_X1   g0768(.A1(new_n967), .A2(new_n968), .ZN(new_n969));
  OAI21_X1  g0769(.A(new_n965), .B1(new_n966), .B2(new_n969), .ZN(new_n970));
  NAND2_X1  g0770(.A1(new_n970), .A2(new_n697), .ZN(new_n971));
  INV_X1    g0771(.A(new_n699), .ZN(new_n972));
  NAND3_X1  g0772(.A1(new_n688), .A2(new_n690), .A3(new_n972), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n973), .A2(new_n700), .ZN(new_n974));
  NAND2_X1  g0774(.A1(new_n974), .A2(new_n744), .ZN(new_n975));
  NAND3_X1  g0775(.A1(new_n973), .A2(new_n696), .A3(new_n700), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n975), .A2(new_n976), .ZN(new_n977));
  NAND2_X1  g0777(.A1(new_n977), .A2(new_n742), .ZN(new_n978));
  NAND2_X1  g0778(.A1(new_n978), .A2(KEYINPUT109), .ZN(new_n979));
  XNOR2_X1  g0779(.A(new_n967), .B(new_n968), .ZN(new_n980));
  INV_X1    g0780(.A(new_n697), .ZN(new_n981));
  NAND3_X1  g0781(.A1(new_n980), .A2(new_n981), .A3(new_n965), .ZN(new_n982));
  INV_X1    g0782(.A(KEYINPUT109), .ZN(new_n983));
  NAND3_X1  g0783(.A1(new_n977), .A2(new_n983), .A3(new_n742), .ZN(new_n984));
  NAND4_X1  g0784(.A1(new_n971), .A2(new_n979), .A3(new_n982), .A4(new_n984), .ZN(new_n985));
  AOI21_X1  g0785(.A(new_n962), .B1(new_n985), .B2(new_n742), .ZN(new_n986));
  OAI211_X1 g0786(.A(new_n959), .B(new_n961), .C1(new_n986), .C2(new_n746), .ZN(new_n987));
  INV_X1    g0787(.A(new_n752), .ZN(new_n988));
  NOR2_X1   g0788(.A1(new_n241), .A2(new_n988), .ZN(new_n989));
  OAI21_X1  g0789(.A(new_n760), .B1(new_n224), .B2(new_n331), .ZN(new_n990));
  OAI21_X1  g0790(.A(new_n747), .B1(new_n989), .B2(new_n990), .ZN(new_n991));
  XOR2_X1   g0791(.A(new_n991), .B(KEYINPUT110), .Z(new_n992));
  OAI221_X1 g0792(.A(new_n277), .B1(new_n252), .B2(new_n764), .C1(new_n769), .C2(new_n297), .ZN(new_n993));
  NAND2_X1  g0793(.A1(new_n774), .A2(G77), .ZN(new_n994));
  OAI21_X1  g0794(.A(new_n994), .B1(new_n837), .B2(new_n780), .ZN(new_n995));
  OAI22_X1  g0795(.A1(new_n802), .A2(new_n781), .B1(new_n209), .B2(new_n777), .ZN(new_n996));
  NOR3_X1   g0796(.A1(new_n993), .A2(new_n995), .A3(new_n996), .ZN(new_n997));
  INV_X1    g0797(.A(G143), .ZN(new_n998));
  OAI221_X1 g0798(.A(new_n997), .B1(new_n202), .B2(new_n790), .C1(new_n998), .C2(new_n795), .ZN(new_n999));
  XNOR2_X1  g0799(.A(KEYINPUT111), .B(G317), .ZN(new_n1000));
  AOI22_X1  g0800(.A1(new_n783), .A2(new_n1000), .B1(new_n775), .B2(G294), .ZN(new_n1001));
  OAI21_X1  g0801(.A(new_n1001), .B1(new_n535), .B2(new_n773), .ZN(new_n1002));
  INV_X1    g0802(.A(new_n777), .ZN(new_n1003));
  NAND3_X1  g0803(.A1(new_n1003), .A2(KEYINPUT46), .A3(G116), .ZN(new_n1004));
  INV_X1    g0804(.A(KEYINPUT46), .ZN(new_n1005));
  OAI21_X1  g0805(.A(new_n1005), .B1(new_n777), .B2(new_n485), .ZN(new_n1006));
  OAI211_X1 g0806(.A(new_n1004), .B(new_n1006), .C1(new_n211), .C2(new_n764), .ZN(new_n1007));
  OAI21_X1  g0807(.A(new_n392), .B1(new_n769), .B2(new_n806), .ZN(new_n1008));
  NOR3_X1   g0808(.A1(new_n1002), .A2(new_n1007), .A3(new_n1008), .ZN(new_n1009));
  OAI221_X1 g0809(.A(new_n1009), .B1(new_n807), .B2(new_n790), .C1(new_n809), .C2(new_n795), .ZN(new_n1010));
  NAND2_X1  g0810(.A1(new_n999), .A2(new_n1010), .ZN(new_n1011));
  INV_X1    g0811(.A(new_n1011), .ZN(new_n1012));
  AND2_X1   g0812(.A1(new_n1012), .A2(KEYINPUT47), .ZN(new_n1013));
  OAI21_X1  g0813(.A(new_n759), .B1(new_n1012), .B2(KEYINPUT47), .ZN(new_n1014));
  OAI221_X1 g0814(.A(new_n992), .B1(new_n1013), .B2(new_n1014), .C1(new_n936), .C2(new_n814), .ZN(new_n1015));
  NAND2_X1  g0815(.A1(new_n987), .A2(new_n1015), .ZN(new_n1016));
  XNOR2_X1  g0816(.A(new_n1016), .B(KEYINPUT112), .ZN(new_n1017));
  INV_X1    g0817(.A(new_n1017), .ZN(G387));
  OAI211_X1 g0818(.A(new_n975), .B(new_n976), .C1(new_n741), .C2(new_n723), .ZN(new_n1019));
  NAND3_X1  g0819(.A1(new_n978), .A2(new_n708), .A3(new_n1019), .ZN(new_n1020));
  NOR2_X1   g0820(.A1(new_n691), .A2(new_n814), .ZN(new_n1021));
  NAND2_X1  g0821(.A1(new_n245), .A2(G45), .ZN(new_n1022));
  NOR2_X1   g0822(.A1(new_n295), .A2(G50), .ZN(new_n1023));
  XNOR2_X1  g0823(.A(new_n1023), .B(KEYINPUT50), .ZN(new_n1024));
  OAI21_X1  g0824(.A(new_n509), .B1(new_n252), .B2(new_n219), .ZN(new_n1025));
  AOI21_X1  g0825(.A(new_n1025), .B1(new_n710), .B2(KEYINPUT113), .ZN(new_n1026));
  OAI211_X1 g0826(.A(new_n1024), .B(new_n1026), .C1(KEYINPUT113), .C2(new_n710), .ZN(new_n1027));
  NAND3_X1  g0827(.A1(new_n1022), .A2(new_n752), .A3(new_n1027), .ZN(new_n1028));
  NAND3_X1  g0828(.A1(new_n277), .A2(new_n224), .A3(new_n710), .ZN(new_n1029));
  OAI211_X1 g0829(.A(new_n1028), .B(new_n1029), .C1(G107), .C2(new_n224), .ZN(new_n1030));
  AOI21_X1  g0830(.A(new_n750), .B1(new_n1030), .B2(new_n760), .ZN(new_n1031));
  NOR2_X1   g0831(.A1(new_n795), .A2(new_n781), .ZN(new_n1032));
  AOI21_X1  g0832(.A(new_n392), .B1(new_n787), .B2(G68), .ZN(new_n1033));
  NAND2_X1  g0833(.A1(new_n765), .A2(new_n330), .ZN(new_n1034));
  OAI211_X1 g0834(.A(new_n1033), .B(new_n1034), .C1(new_n769), .C2(new_n202), .ZN(new_n1035));
  OAI22_X1  g0835(.A1(new_n777), .A2(new_n219), .B1(new_n773), .B2(new_n535), .ZN(new_n1036));
  OAI22_X1  g0836(.A1(new_n802), .A2(new_n295), .B1(new_n780), .B2(new_n297), .ZN(new_n1037));
  NOR4_X1   g0837(.A1(new_n1032), .A2(new_n1035), .A3(new_n1036), .A4(new_n1037), .ZN(new_n1038));
  AOI22_X1  g0838(.A1(new_n768), .A2(new_n1000), .B1(G311), .B2(new_n775), .ZN(new_n1039));
  OAI221_X1 g0839(.A(new_n1039), .B1(new_n795), .B2(new_n800), .C1(new_n806), .C2(new_n790), .ZN(new_n1040));
  XNOR2_X1  g0840(.A(new_n1040), .B(KEYINPUT48), .ZN(new_n1041));
  OAI221_X1 g0841(.A(new_n1041), .B1(new_n807), .B2(new_n764), .C1(new_n810), .C2(new_n777), .ZN(new_n1042));
  XNOR2_X1  g0842(.A(new_n1042), .B(KEYINPUT49), .ZN(new_n1043));
  NOR2_X1   g0843(.A1(new_n773), .A2(new_n485), .ZN(new_n1044));
  AOI211_X1 g0844(.A(new_n1044), .B(new_n499), .C1(new_n783), .C2(new_n798), .ZN(new_n1045));
  AOI21_X1  g0845(.A(new_n1038), .B1(new_n1043), .B2(new_n1045), .ZN(new_n1046));
  OAI21_X1  g0846(.A(new_n1031), .B1(new_n1046), .B2(new_n762), .ZN(new_n1047));
  OR3_X1    g0847(.A1(new_n1021), .A2(KEYINPUT114), .A3(new_n1047), .ZN(new_n1048));
  OAI21_X1  g0848(.A(KEYINPUT114), .B1(new_n1021), .B2(new_n1047), .ZN(new_n1049));
  AOI22_X1  g0849(.A1(new_n1048), .A2(new_n1049), .B1(new_n977), .B2(new_n746), .ZN(new_n1050));
  NAND2_X1  g0850(.A1(new_n1020), .A2(new_n1050), .ZN(G393));
  INV_X1    g0851(.A(new_n982), .ZN(new_n1052));
  AOI21_X1  g0852(.A(new_n981), .B1(new_n980), .B2(new_n965), .ZN(new_n1053));
  OAI21_X1  g0853(.A(new_n978), .B1(new_n1052), .B2(new_n1053), .ZN(new_n1054));
  NAND3_X1  g0854(.A1(new_n1054), .A2(new_n708), .A3(new_n985), .ZN(new_n1055));
  NAND3_X1  g0855(.A1(new_n971), .A2(new_n746), .A3(new_n982), .ZN(new_n1056));
  OAI221_X1 g0856(.A(new_n760), .B1(new_n535), .B2(new_n224), .C1(new_n250), .C2(new_n988), .ZN(new_n1057));
  NAND2_X1  g0857(.A1(new_n1057), .A2(new_n747), .ZN(new_n1058));
  AOI22_X1  g0858(.A1(new_n796), .A2(G317), .B1(G311), .B2(new_n768), .ZN(new_n1059));
  XNOR2_X1  g0859(.A(new_n1059), .B(KEYINPUT52), .ZN(new_n1060));
  OAI221_X1 g0860(.A(new_n322), .B1(new_n485), .B2(new_n764), .C1(new_n810), .C2(new_n786), .ZN(new_n1061));
  OAI22_X1  g0861(.A1(new_n777), .A2(new_n807), .B1(new_n773), .B2(new_n211), .ZN(new_n1062));
  OAI22_X1  g0862(.A1(new_n802), .A2(new_n806), .B1(new_n780), .B2(new_n800), .ZN(new_n1063));
  OR3_X1    g0863(.A1(new_n1061), .A2(new_n1062), .A3(new_n1063), .ZN(new_n1064));
  OAI22_X1  g0864(.A1(new_n795), .A2(new_n297), .B1(new_n781), .B2(new_n769), .ZN(new_n1065));
  INV_X1    g0865(.A(KEYINPUT51), .ZN(new_n1066));
  NAND2_X1  g0866(.A1(new_n1065), .A2(new_n1066), .ZN(new_n1067));
  OAI22_X1  g0867(.A1(new_n777), .A2(new_n207), .B1(new_n780), .B2(new_n998), .ZN(new_n1068));
  XNOR2_X1  g0868(.A(new_n1068), .B(KEYINPUT115), .ZN(new_n1069));
  NOR2_X1   g0869(.A1(new_n764), .A2(new_n219), .ZN(new_n1070));
  OAI22_X1  g0870(.A1(new_n802), .A2(new_n202), .B1(new_n773), .B2(new_n611), .ZN(new_n1071));
  NOR4_X1   g0871(.A1(new_n1069), .A2(new_n392), .A3(new_n1070), .A4(new_n1071), .ZN(new_n1072));
  OAI211_X1 g0872(.A(new_n1067), .B(new_n1072), .C1(new_n295), .C2(new_n790), .ZN(new_n1073));
  NOR2_X1   g0873(.A1(new_n1065), .A2(new_n1066), .ZN(new_n1074));
  OAI22_X1  g0874(.A1(new_n1060), .A2(new_n1064), .B1(new_n1073), .B2(new_n1074), .ZN(new_n1075));
  INV_X1    g0875(.A(KEYINPUT116), .ZN(new_n1076));
  OR2_X1    g0876(.A1(new_n1075), .A2(new_n1076), .ZN(new_n1077));
  AOI21_X1  g0877(.A(new_n762), .B1(new_n1075), .B2(new_n1076), .ZN(new_n1078));
  AOI21_X1  g0878(.A(new_n1058), .B1(new_n1077), .B2(new_n1078), .ZN(new_n1079));
  OAI21_X1  g0879(.A(new_n1079), .B1(new_n814), .B2(new_n941), .ZN(new_n1080));
  AND2_X1   g0880(.A1(new_n1056), .A2(new_n1080), .ZN(new_n1081));
  NAND2_X1  g0881(.A1(new_n1055), .A2(new_n1081), .ZN(G390));
  XNOR2_X1  g0882(.A(new_n925), .B(KEYINPUT117), .ZN(new_n1083));
  AOI21_X1  g0883(.A(new_n1083), .B1(new_n889), .B2(new_n900), .ZN(new_n1084));
  INV_X1    g0884(.A(new_n820), .ZN(new_n1085));
  AOI21_X1  g0885(.A(new_n1085), .B1(new_n722), .B2(new_n819), .ZN(new_n1086));
  INV_X1    g0886(.A(new_n858), .ZN(new_n1087));
  OAI21_X1  g0887(.A(new_n1084), .B1(new_n1086), .B2(new_n1087), .ZN(new_n1088));
  AOI21_X1  g0888(.A(new_n925), .B1(new_n921), .B2(new_n858), .ZN(new_n1089));
  OAI21_X1  g0889(.A(new_n1088), .B1(new_n927), .B2(new_n1089), .ZN(new_n1090));
  AND2_X1   g0890(.A1(new_n859), .A2(G330), .ZN(new_n1091));
  NAND2_X1  g0891(.A1(new_n1090), .A2(new_n1091), .ZN(new_n1092));
  NAND2_X1  g0892(.A1(new_n859), .A2(G330), .ZN(new_n1093));
  OAI211_X1 g0893(.A(new_n1088), .B(new_n1093), .C1(new_n927), .C2(new_n1089), .ZN(new_n1094));
  NAND2_X1  g0894(.A1(new_n1092), .A2(new_n1094), .ZN(new_n1095));
  NAND3_X1  g0895(.A1(new_n916), .A2(new_n673), .A3(new_n906), .ZN(new_n1096));
  AND3_X1   g0896(.A1(new_n854), .A2(G330), .A3(new_n821), .ZN(new_n1097));
  NOR2_X1   g0897(.A1(new_n1097), .A2(new_n858), .ZN(new_n1098));
  OAI21_X1  g0898(.A(new_n921), .B1(new_n1091), .B2(new_n1098), .ZN(new_n1099));
  INV_X1    g0899(.A(KEYINPUT118), .ZN(new_n1100));
  OAI21_X1  g0900(.A(new_n1100), .B1(new_n1097), .B2(new_n858), .ZN(new_n1101));
  NAND3_X1  g0901(.A1(new_n854), .A2(G330), .A3(new_n821), .ZN(new_n1102));
  NAND3_X1  g0902(.A1(new_n1102), .A2(KEYINPUT118), .A3(new_n1087), .ZN(new_n1103));
  NAND4_X1  g0903(.A1(new_n1101), .A2(new_n1093), .A3(new_n1103), .A4(new_n1086), .ZN(new_n1104));
  AOI21_X1  g0904(.A(new_n1096), .B1(new_n1099), .B2(new_n1104), .ZN(new_n1105));
  INV_X1    g0905(.A(new_n1105), .ZN(new_n1106));
  NAND2_X1  g0906(.A1(new_n1095), .A2(new_n1106), .ZN(new_n1107));
  NAND3_X1  g0907(.A1(new_n1092), .A2(new_n1105), .A3(new_n1094), .ZN(new_n1108));
  NAND3_X1  g0908(.A1(new_n1107), .A2(new_n708), .A3(new_n1108), .ZN(new_n1109));
  NAND3_X1  g0909(.A1(new_n1092), .A2(new_n746), .A3(new_n1094), .ZN(new_n1110));
  INV_X1    g0910(.A(KEYINPUT120), .ZN(new_n1111));
  INV_X1    g0911(.A(new_n826), .ZN(new_n1112));
  OAI21_X1  g0912(.A(new_n747), .B1(new_n328), .B2(new_n1112), .ZN(new_n1113));
  AOI22_X1  g0913(.A1(G97), .A2(new_n791), .B1(new_n796), .B2(G283), .ZN(new_n1114));
  NOR2_X1   g0914(.A1(new_n780), .A2(new_n810), .ZN(new_n1115));
  OAI22_X1  g0915(.A1(new_n777), .A2(new_n611), .B1(new_n773), .B2(new_n252), .ZN(new_n1116));
  AOI211_X1 g0916(.A(new_n1115), .B(new_n1116), .C1(G107), .C2(new_n775), .ZN(new_n1117));
  AOI211_X1 g0917(.A(new_n277), .B(new_n1070), .C1(G116), .C2(new_n768), .ZN(new_n1118));
  NAND3_X1  g0918(.A1(new_n1114), .A2(new_n1117), .A3(new_n1118), .ZN(new_n1119));
  AOI21_X1  g0919(.A(new_n322), .B1(G50), .B2(new_n774), .ZN(new_n1120));
  AOI22_X1  g0920(.A1(new_n796), .A2(G128), .B1(new_n1120), .B2(KEYINPUT119), .ZN(new_n1121));
  XOR2_X1   g0921(.A(KEYINPUT54), .B(G143), .Z(new_n1122));
  INV_X1    g0922(.A(new_n1122), .ZN(new_n1123));
  OAI221_X1 g0923(.A(new_n1121), .B1(KEYINPUT119), .B2(new_n1120), .C1(new_n790), .C2(new_n1123), .ZN(new_n1124));
  NOR3_X1   g0924(.A1(new_n777), .A2(KEYINPUT53), .A3(new_n297), .ZN(new_n1125));
  INV_X1    g0925(.A(KEYINPUT53), .ZN(new_n1126));
  AOI21_X1  g0926(.A(new_n1126), .B1(new_n1003), .B2(G150), .ZN(new_n1127));
  AOI211_X1 g0927(.A(new_n1125), .B(new_n1127), .C1(G132), .C2(new_n768), .ZN(new_n1128));
  AOI22_X1  g0928(.A1(new_n783), .A2(G125), .B1(new_n775), .B2(G137), .ZN(new_n1129));
  OAI211_X1 g0929(.A(new_n1128), .B(new_n1129), .C1(new_n781), .C2(new_n764), .ZN(new_n1130));
  OAI21_X1  g0930(.A(new_n1119), .B1(new_n1124), .B2(new_n1130), .ZN(new_n1131));
  AOI21_X1  g0931(.A(new_n1113), .B1(new_n1131), .B2(new_n759), .ZN(new_n1132));
  OAI21_X1  g0932(.A(new_n1132), .B1(new_n927), .B2(new_n757), .ZN(new_n1133));
  AND3_X1   g0933(.A1(new_n1110), .A2(new_n1111), .A3(new_n1133), .ZN(new_n1134));
  AOI21_X1  g0934(.A(new_n1111), .B1(new_n1110), .B2(new_n1133), .ZN(new_n1135));
  OAI21_X1  g0935(.A(new_n1109), .B1(new_n1134), .B2(new_n1135), .ZN(G378));
  NAND2_X1  g0936(.A1(new_n303), .A2(new_n866), .ZN(new_n1137));
  INV_X1    g0937(.A(new_n1137), .ZN(new_n1138));
  XNOR2_X1  g0938(.A(new_n315), .B(new_n1138), .ZN(new_n1139));
  XNOR2_X1  g0939(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1140));
  XOR2_X1   g0940(.A(new_n1139), .B(new_n1140), .Z(new_n1141));
  NAND2_X1  g0941(.A1(new_n905), .A2(new_n1141), .ZN(new_n1142));
  INV_X1    g0942(.A(new_n1141), .ZN(new_n1143));
  NAND4_X1  g0943(.A1(new_n909), .A2(G330), .A3(new_n895), .A4(new_n1143), .ZN(new_n1144));
  NAND2_X1  g0944(.A1(new_n1142), .A2(new_n1144), .ZN(new_n1145));
  INV_X1    g0945(.A(new_n928), .ZN(new_n1146));
  NAND2_X1  g0946(.A1(new_n1145), .A2(new_n1146), .ZN(new_n1147));
  NAND3_X1  g0947(.A1(new_n1142), .A2(new_n928), .A3(new_n1144), .ZN(new_n1148));
  NAND2_X1  g0948(.A1(new_n1147), .A2(new_n1148), .ZN(new_n1149));
  NAND2_X1  g0949(.A1(new_n1141), .A2(new_n756), .ZN(new_n1150));
  OAI21_X1  g0950(.A(new_n747), .B1(G50), .B2(new_n1112), .ZN(new_n1151));
  NOR2_X1   g0951(.A1(G33), .A2(G41), .ZN(new_n1152));
  AOI211_X1 g0952(.A(G50), .B(new_n1152), .C1(new_n392), .C2(new_n263), .ZN(new_n1153));
  AOI22_X1  g0953(.A1(new_n1003), .A2(G77), .B1(new_n774), .B2(G58), .ZN(new_n1154));
  OAI21_X1  g0954(.A(new_n1154), .B1(new_n807), .B2(new_n780), .ZN(new_n1155));
  OAI22_X1  g0955(.A1(new_n769), .A2(new_n211), .B1(new_n252), .B2(new_n764), .ZN(new_n1156));
  NOR4_X1   g0956(.A1(new_n1155), .A2(new_n1156), .A3(G41), .A4(new_n499), .ZN(new_n1157));
  AOI22_X1  g0957(.A1(new_n787), .A2(new_n330), .B1(G97), .B2(new_n775), .ZN(new_n1158));
  XNOR2_X1  g0958(.A(new_n1158), .B(KEYINPUT121), .ZN(new_n1159));
  OAI211_X1 g0959(.A(new_n1157), .B(new_n1159), .C1(new_n485), .C2(new_n795), .ZN(new_n1160));
  INV_X1    g0960(.A(KEYINPUT58), .ZN(new_n1161));
  AOI21_X1  g0961(.A(new_n1153), .B1(new_n1160), .B2(new_n1161), .ZN(new_n1162));
  AOI22_X1  g0962(.A1(new_n765), .A2(G150), .B1(new_n1003), .B2(new_n1122), .ZN(new_n1163));
  INV_X1    g0963(.A(G128), .ZN(new_n1164));
  OAI21_X1  g0964(.A(new_n1163), .B1(new_n769), .B2(new_n1164), .ZN(new_n1165));
  AOI21_X1  g0965(.A(new_n1165), .B1(new_n796), .B2(G125), .ZN(new_n1166));
  AOI22_X1  g0966(.A1(new_n787), .A2(G137), .B1(G132), .B2(new_n775), .ZN(new_n1167));
  XNOR2_X1  g0967(.A(new_n1167), .B(KEYINPUT122), .ZN(new_n1168));
  NAND2_X1  g0968(.A1(new_n1166), .A2(new_n1168), .ZN(new_n1169));
  XNOR2_X1  g0969(.A(new_n1169), .B(KEYINPUT59), .ZN(new_n1170));
  INV_X1    g0970(.A(G124), .ZN(new_n1171));
  OAI221_X1 g0971(.A(new_n1152), .B1(new_n773), .B2(new_n781), .C1(new_n1171), .C2(new_n780), .ZN(new_n1172));
  OAI221_X1 g0972(.A(new_n1162), .B1(new_n1161), .B2(new_n1160), .C1(new_n1170), .C2(new_n1172), .ZN(new_n1173));
  AOI21_X1  g0973(.A(new_n1151), .B1(new_n1173), .B2(new_n759), .ZN(new_n1174));
  AOI22_X1  g0974(.A1(new_n1149), .A2(new_n746), .B1(new_n1150), .B2(new_n1174), .ZN(new_n1175));
  INV_X1    g0975(.A(new_n1096), .ZN(new_n1176));
  NAND2_X1  g0976(.A1(new_n1108), .A2(new_n1176), .ZN(new_n1177));
  AND3_X1   g0977(.A1(new_n1142), .A2(new_n928), .A3(new_n1144), .ZN(new_n1178));
  AOI21_X1  g0978(.A(new_n928), .B1(new_n1142), .B2(new_n1144), .ZN(new_n1179));
  OAI211_X1 g0979(.A(new_n1177), .B(KEYINPUT57), .C1(new_n1178), .C2(new_n1179), .ZN(new_n1180));
  NAND2_X1  g0980(.A1(new_n1180), .A2(new_n708), .ZN(new_n1181));
  AOI21_X1  g0981(.A(KEYINPUT57), .B1(new_n1149), .B2(new_n1177), .ZN(new_n1182));
  OAI21_X1  g0982(.A(new_n1175), .B1(new_n1181), .B2(new_n1182), .ZN(G375));
  AOI21_X1  g0983(.A(new_n750), .B1(new_n252), .B2(new_n826), .ZN(new_n1184));
  AOI22_X1  g0984(.A1(G107), .A2(new_n791), .B1(new_n796), .B2(G294), .ZN(new_n1185));
  OAI211_X1 g0985(.A(new_n1034), .B(new_n322), .C1(new_n769), .C2(new_n807), .ZN(new_n1186));
  OAI21_X1  g0986(.A(new_n994), .B1(new_n802), .B2(new_n485), .ZN(new_n1187));
  OAI22_X1  g0987(.A1(new_n777), .A2(new_n535), .B1(new_n780), .B2(new_n806), .ZN(new_n1188));
  NOR3_X1   g0988(.A1(new_n1186), .A2(new_n1187), .A3(new_n1188), .ZN(new_n1189));
  NAND2_X1  g0989(.A1(new_n796), .A2(G132), .ZN(new_n1190));
  OAI21_X1  g0990(.A(new_n499), .B1(new_n769), .B2(new_n837), .ZN(new_n1191));
  OAI22_X1  g0991(.A1(new_n802), .A2(new_n1123), .B1(new_n780), .B2(new_n1164), .ZN(new_n1192));
  OAI22_X1  g0992(.A1(new_n777), .A2(new_n781), .B1(new_n773), .B2(new_n209), .ZN(new_n1193));
  OAI22_X1  g0993(.A1(new_n786), .A2(new_n297), .B1(new_n764), .B2(new_n202), .ZN(new_n1194));
  NOR4_X1   g0994(.A1(new_n1191), .A2(new_n1192), .A3(new_n1193), .A4(new_n1194), .ZN(new_n1195));
  AOI22_X1  g0995(.A1(new_n1185), .A2(new_n1189), .B1(new_n1190), .B2(new_n1195), .ZN(new_n1196));
  OAI221_X1 g0996(.A(new_n1184), .B1(new_n762), .B2(new_n1196), .C1(new_n858), .C2(new_n757), .ZN(new_n1197));
  AND2_X1   g0997(.A1(new_n1099), .A2(new_n1104), .ZN(new_n1198));
  OAI211_X1 g0998(.A(KEYINPUT123), .B(new_n1197), .C1(new_n1198), .C2(new_n745), .ZN(new_n1199));
  INV_X1    g0999(.A(KEYINPUT123), .ZN(new_n1200));
  AOI21_X1  g1000(.A(new_n745), .B1(new_n1099), .B2(new_n1104), .ZN(new_n1201));
  INV_X1    g1001(.A(new_n1197), .ZN(new_n1202));
  OAI21_X1  g1002(.A(new_n1200), .B1(new_n1201), .B2(new_n1202), .ZN(new_n1203));
  NAND2_X1  g1003(.A1(new_n1199), .A2(new_n1203), .ZN(new_n1204));
  INV_X1    g1004(.A(new_n962), .ZN(new_n1205));
  NAND3_X1  g1005(.A1(new_n1099), .A2(new_n1104), .A3(new_n1096), .ZN(new_n1206));
  NAND3_X1  g1006(.A1(new_n1106), .A2(new_n1205), .A3(new_n1206), .ZN(new_n1207));
  NAND2_X1  g1007(.A1(new_n1204), .A2(new_n1207), .ZN(G381));
  INV_X1    g1008(.A(G396), .ZN(new_n1209));
  NAND3_X1  g1009(.A1(new_n1020), .A2(new_n1209), .A3(new_n1050), .ZN(new_n1210));
  NOR4_X1   g1010(.A1(G390), .A2(G384), .A3(G381), .A4(new_n1210), .ZN(new_n1211));
  NAND2_X1  g1011(.A1(new_n1017), .A2(new_n1211), .ZN(new_n1212));
  INV_X1    g1012(.A(G375), .ZN(new_n1213));
  AND3_X1   g1013(.A1(new_n1109), .A2(new_n1110), .A3(new_n1133), .ZN(new_n1214));
  NAND2_X1  g1014(.A1(new_n1213), .A2(new_n1214), .ZN(new_n1215));
  OR2_X1    g1015(.A1(new_n1212), .A2(new_n1215), .ZN(G407));
  NAND3_X1  g1016(.A1(new_n1213), .A2(new_n681), .A3(new_n1214), .ZN(new_n1217));
  OAI211_X1 g1017(.A(G213), .B(new_n1217), .C1(new_n1212), .C2(new_n1215), .ZN(G409));
  AOI21_X1  g1018(.A(new_n1209), .B1(new_n1020), .B2(new_n1050), .ZN(new_n1219));
  INV_X1    g1019(.A(new_n1219), .ZN(new_n1220));
  AOI21_X1  g1020(.A(KEYINPUT112), .B1(new_n1220), .B2(new_n1210), .ZN(new_n1221));
  NOR2_X1   g1021(.A1(G390), .A2(new_n1221), .ZN(new_n1222));
  INV_X1    g1022(.A(new_n1210), .ZN(new_n1223));
  NOR2_X1   g1023(.A1(new_n1223), .A2(new_n1219), .ZN(new_n1224));
  AOI21_X1  g1024(.A(new_n1224), .B1(new_n1055), .B2(new_n1081), .ZN(new_n1225));
  OAI211_X1 g1025(.A(new_n987), .B(new_n1015), .C1(new_n1222), .C2(new_n1225), .ZN(new_n1226));
  OAI211_X1 g1026(.A(new_n1055), .B(new_n1081), .C1(new_n1224), .C2(KEYINPUT112), .ZN(new_n1227));
  NAND2_X1  g1027(.A1(new_n1220), .A2(new_n1210), .ZN(new_n1228));
  NAND2_X1  g1028(.A1(G390), .A2(new_n1228), .ZN(new_n1229));
  NAND3_X1  g1029(.A1(new_n1016), .A2(new_n1227), .A3(new_n1229), .ZN(new_n1230));
  INV_X1    g1030(.A(KEYINPUT61), .ZN(new_n1231));
  AND3_X1   g1031(.A1(new_n1226), .A2(new_n1230), .A3(new_n1231), .ZN(new_n1232));
  OAI211_X1 g1032(.A(G378), .B(new_n1175), .C1(new_n1181), .C2(new_n1182), .ZN(new_n1233));
  AND3_X1   g1033(.A1(new_n1149), .A2(new_n1205), .A3(new_n1177), .ZN(new_n1234));
  NAND2_X1  g1034(.A1(new_n1150), .A2(new_n1174), .ZN(new_n1235));
  NOR2_X1   g1035(.A1(new_n1178), .A2(new_n1179), .ZN(new_n1236));
  OAI21_X1  g1036(.A(new_n1235), .B1(new_n1236), .B2(new_n745), .ZN(new_n1237));
  OAI21_X1  g1037(.A(new_n1214), .B1(new_n1234), .B2(new_n1237), .ZN(new_n1238));
  NAND2_X1  g1038(.A1(new_n1233), .A2(new_n1238), .ZN(new_n1239));
  INV_X1    g1039(.A(G213), .ZN(new_n1240));
  NOR2_X1   g1040(.A1(new_n1240), .A2(G343), .ZN(new_n1241));
  INV_X1    g1041(.A(new_n1241), .ZN(new_n1242));
  NAND2_X1  g1042(.A1(new_n1239), .A2(new_n1242), .ZN(new_n1243));
  NAND3_X1  g1043(.A1(new_n1198), .A2(KEYINPUT60), .A3(new_n1096), .ZN(new_n1244));
  INV_X1    g1044(.A(KEYINPUT60), .ZN(new_n1245));
  NAND2_X1  g1045(.A1(new_n1206), .A2(new_n1245), .ZN(new_n1246));
  NAND4_X1  g1046(.A1(new_n1244), .A2(new_n708), .A3(new_n1106), .A4(new_n1246), .ZN(new_n1247));
  AOI21_X1  g1047(.A(G384), .B1(new_n1204), .B2(new_n1247), .ZN(new_n1248));
  INV_X1    g1048(.A(new_n1248), .ZN(new_n1249));
  NAND3_X1  g1049(.A1(new_n1204), .A2(new_n1247), .A3(G384), .ZN(new_n1250));
  NAND3_X1  g1050(.A1(new_n1249), .A2(KEYINPUT124), .A3(new_n1250), .ZN(new_n1251));
  INV_X1    g1051(.A(KEYINPUT124), .ZN(new_n1252));
  INV_X1    g1052(.A(new_n1250), .ZN(new_n1253));
  OAI21_X1  g1053(.A(new_n1252), .B1(new_n1253), .B2(new_n1248), .ZN(new_n1254));
  NAND2_X1  g1054(.A1(new_n1241), .A2(G2897), .ZN(new_n1255));
  NAND3_X1  g1055(.A1(new_n1251), .A2(new_n1254), .A3(new_n1255), .ZN(new_n1256));
  INV_X1    g1056(.A(new_n1256), .ZN(new_n1257));
  INV_X1    g1057(.A(new_n1255), .ZN(new_n1258));
  NOR2_X1   g1058(.A1(new_n1253), .A2(new_n1248), .ZN(new_n1259));
  AOI22_X1  g1059(.A1(new_n1243), .A2(new_n1257), .B1(new_n1258), .B2(new_n1259), .ZN(new_n1260));
  INV_X1    g1060(.A(KEYINPUT63), .ZN(new_n1261));
  NAND2_X1  g1061(.A1(new_n1251), .A2(new_n1254), .ZN(new_n1262));
  INV_X1    g1062(.A(new_n1262), .ZN(new_n1263));
  OAI21_X1  g1063(.A(new_n1261), .B1(new_n1243), .B2(new_n1263), .ZN(new_n1264));
  AOI21_X1  g1064(.A(new_n1241), .B1(new_n1233), .B2(new_n1238), .ZN(new_n1265));
  NAND3_X1  g1065(.A1(new_n1265), .A2(KEYINPUT63), .A3(new_n1262), .ZN(new_n1266));
  NAND4_X1  g1066(.A1(new_n1232), .A2(new_n1260), .A3(new_n1264), .A4(new_n1266), .ZN(new_n1267));
  NAND2_X1  g1067(.A1(new_n1259), .A2(new_n1258), .ZN(new_n1268));
  XNOR2_X1  g1068(.A(KEYINPUT125), .B(KEYINPUT61), .ZN(new_n1269));
  OAI211_X1 g1069(.A(new_n1268), .B(new_n1269), .C1(new_n1265), .C2(new_n1256), .ZN(new_n1270));
  INV_X1    g1070(.A(KEYINPUT62), .ZN(new_n1271));
  AND4_X1   g1071(.A1(new_n1271), .A2(new_n1239), .A3(new_n1242), .A4(new_n1262), .ZN(new_n1272));
  AOI21_X1  g1072(.A(new_n1271), .B1(new_n1265), .B2(new_n1262), .ZN(new_n1273));
  NOR3_X1   g1073(.A1(new_n1270), .A2(new_n1272), .A3(new_n1273), .ZN(new_n1274));
  NAND2_X1  g1074(.A1(new_n1226), .A2(new_n1230), .ZN(new_n1275));
  INV_X1    g1075(.A(new_n1275), .ZN(new_n1276));
  OAI21_X1  g1076(.A(new_n1267), .B1(new_n1274), .B2(new_n1276), .ZN(G405));
  INV_X1    g1077(.A(KEYINPUT127), .ZN(new_n1278));
  NAND2_X1  g1078(.A1(new_n1275), .A2(new_n1278), .ZN(new_n1279));
  NAND3_X1  g1079(.A1(new_n1226), .A2(new_n1230), .A3(KEYINPUT127), .ZN(new_n1280));
  NAND2_X1  g1080(.A1(G375), .A2(new_n1214), .ZN(new_n1281));
  AOI22_X1  g1081(.A1(new_n1233), .A2(new_n1281), .B1(new_n1262), .B2(KEYINPUT126), .ZN(new_n1282));
  INV_X1    g1082(.A(KEYINPUT126), .ZN(new_n1283));
  NAND2_X1  g1083(.A1(new_n1283), .A2(KEYINPUT124), .ZN(new_n1284));
  NAND4_X1  g1084(.A1(new_n1281), .A2(new_n1259), .A3(new_n1233), .A4(new_n1284), .ZN(new_n1285));
  INV_X1    g1085(.A(new_n1285), .ZN(new_n1286));
  OAI211_X1 g1086(.A(new_n1279), .B(new_n1280), .C1(new_n1282), .C2(new_n1286), .ZN(new_n1287));
  NOR2_X1   g1087(.A1(new_n1286), .A2(new_n1282), .ZN(new_n1288));
  NAND3_X1  g1088(.A1(new_n1288), .A2(new_n1278), .A3(new_n1275), .ZN(new_n1289));
  NAND2_X1  g1089(.A1(new_n1287), .A2(new_n1289), .ZN(G402));
endmodule


