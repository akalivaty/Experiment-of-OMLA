//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 1 0 0 1 0 1 1 1 0 1 1 0 0 1 0 0 0 0 1 0 0 1 1 0 1 0 1 0 0 1 1 0 1 0 0 0 1 0 0 1 0 1 0 1 0 1 1 0 1 0 1 1 0 1 1 1 0 1 1 0 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:41:21 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n236, new_n237,
    new_n238, new_n240, new_n241, new_n242, new_n243, new_n244, new_n245,
    new_n246, new_n247, new_n248, new_n250, new_n251, new_n252, new_n253,
    new_n254, new_n255, new_n256, new_n257, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1246, new_n1247,
    new_n1248, new_n1250, new_n1251, new_n1252, new_n1253, new_n1254,
    new_n1255, new_n1256, new_n1257, new_n1258, new_n1259, new_n1260,
    new_n1261, new_n1263, new_n1264, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1315, new_n1316, new_n1317,
    new_n1318, new_n1319, new_n1320;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0005(.A1(G1), .A2(G20), .ZN(new_n206));
  AOI22_X1  g0006(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n207));
  INV_X1    g0007(.A(G68), .ZN(new_n208));
  INV_X1    g0008(.A(G238), .ZN(new_n209));
  INV_X1    g0009(.A(G87), .ZN(new_n210));
  INV_X1    g0010(.A(G250), .ZN(new_n211));
  OAI221_X1 g0011(.A(new_n207), .B1(new_n208), .B2(new_n209), .C1(new_n210), .C2(new_n211), .ZN(new_n212));
  AOI22_X1  g0012(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n213));
  INV_X1    g0013(.A(G77), .ZN(new_n214));
  INV_X1    g0014(.A(G244), .ZN(new_n215));
  INV_X1    g0015(.A(G107), .ZN(new_n216));
  INV_X1    g0016(.A(G264), .ZN(new_n217));
  OAI221_X1 g0017(.A(new_n213), .B1(new_n214), .B2(new_n215), .C1(new_n216), .C2(new_n217), .ZN(new_n218));
  OAI21_X1  g0018(.A(new_n206), .B1(new_n212), .B2(new_n218), .ZN(new_n219));
  OR2_X1    g0019(.A1(new_n219), .A2(KEYINPUT1), .ZN(new_n220));
  NOR2_X1   g0020(.A1(new_n206), .A2(G13), .ZN(new_n221));
  INV_X1    g0021(.A(new_n221), .ZN(new_n222));
  INV_X1    g0022(.A(G257), .ZN(new_n223));
  AOI211_X1 g0023(.A(new_n211), .B(new_n222), .C1(new_n223), .C2(new_n217), .ZN(new_n224));
  OR2_X1    g0024(.A1(new_n224), .A2(KEYINPUT0), .ZN(new_n225));
  INV_X1    g0025(.A(G20), .ZN(new_n226));
  NAND2_X1  g0026(.A1(new_n226), .A2(KEYINPUT64), .ZN(new_n227));
  INV_X1    g0027(.A(KEYINPUT64), .ZN(new_n228));
  NAND2_X1  g0028(.A1(new_n228), .A2(G20), .ZN(new_n229));
  NAND2_X1  g0029(.A1(new_n227), .A2(new_n229), .ZN(new_n230));
  NAND2_X1  g0030(.A1(G1), .A2(G13), .ZN(new_n231));
  INV_X1    g0031(.A(new_n231), .ZN(new_n232));
  NAND2_X1  g0032(.A1(new_n230), .A2(new_n232), .ZN(new_n233));
  INV_X1    g0033(.A(new_n201), .ZN(new_n234));
  NAND2_X1  g0034(.A1(new_n234), .A2(G50), .ZN(new_n235));
  NOR2_X1   g0035(.A1(new_n233), .A2(new_n235), .ZN(new_n236));
  AOI21_X1  g0036(.A(new_n236), .B1(new_n224), .B2(KEYINPUT0), .ZN(new_n237));
  NAND3_X1  g0037(.A1(new_n220), .A2(new_n225), .A3(new_n237), .ZN(new_n238));
  AOI21_X1  g0038(.A(new_n238), .B1(KEYINPUT1), .B2(new_n219), .ZN(G361));
  XNOR2_X1  g0039(.A(G250), .B(G257), .ZN(new_n240));
  XNOR2_X1  g0040(.A(G264), .B(G270), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n242), .B(KEYINPUT65), .ZN(new_n243));
  XNOR2_X1  g0043(.A(G238), .B(G244), .ZN(new_n244));
  INV_X1    g0044(.A(G232), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n244), .B(new_n245), .ZN(new_n246));
  XNOR2_X1  g0046(.A(KEYINPUT2), .B(G226), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n246), .B(new_n247), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n243), .B(new_n248), .ZN(G358));
  NAND2_X1  g0049(.A1(new_n202), .A2(G68), .ZN(new_n250));
  NAND2_X1  g0050(.A1(new_n208), .A2(G50), .ZN(new_n251));
  NAND2_X1  g0051(.A1(new_n250), .A2(new_n251), .ZN(new_n252));
  XNOR2_X1  g0052(.A(G58), .B(G77), .ZN(new_n253));
  XNOR2_X1  g0053(.A(new_n252), .B(new_n253), .ZN(new_n254));
  XNOR2_X1  g0054(.A(G87), .B(G116), .ZN(new_n255));
  XNOR2_X1  g0055(.A(G97), .B(G107), .ZN(new_n256));
  XNOR2_X1  g0056(.A(new_n255), .B(new_n256), .ZN(new_n257));
  XOR2_X1   g0057(.A(new_n254), .B(new_n257), .Z(G351));
  INV_X1    g0058(.A(G1), .ZN(new_n259));
  OAI21_X1  g0059(.A(new_n259), .B1(G41), .B2(G45), .ZN(new_n260));
  INV_X1    g0060(.A(G274), .ZN(new_n261));
  NOR2_X1   g0061(.A1(new_n260), .A2(new_n261), .ZN(new_n262));
  AOI21_X1  g0062(.A(new_n231), .B1(G33), .B2(G41), .ZN(new_n263));
  INV_X1    g0063(.A(new_n260), .ZN(new_n264));
  NOR2_X1   g0064(.A1(new_n263), .A2(new_n264), .ZN(new_n265));
  AND2_X1   g0065(.A1(new_n265), .A2(G226), .ZN(new_n266));
  INV_X1    g0066(.A(KEYINPUT3), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n267), .A2(G33), .ZN(new_n268));
  INV_X1    g0068(.A(G33), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n269), .A2(KEYINPUT3), .ZN(new_n270));
  INV_X1    g0070(.A(KEYINPUT66), .ZN(new_n271));
  AND3_X1   g0071(.A1(new_n268), .A2(new_n270), .A3(new_n271), .ZN(new_n272));
  AOI21_X1  g0072(.A(new_n271), .B1(new_n268), .B2(new_n270), .ZN(new_n273));
  NOR2_X1   g0073(.A1(new_n272), .A2(new_n273), .ZN(new_n274));
  INV_X1    g0074(.A(G1698), .ZN(new_n275));
  NAND3_X1  g0075(.A1(new_n274), .A2(G222), .A3(new_n275), .ZN(new_n276));
  NAND3_X1  g0076(.A1(new_n274), .A2(G223), .A3(G1698), .ZN(new_n277));
  OAI211_X1 g0077(.A(new_n276), .B(new_n277), .C1(new_n214), .C2(new_n274), .ZN(new_n278));
  AOI211_X1 g0078(.A(new_n262), .B(new_n266), .C1(new_n278), .C2(new_n263), .ZN(new_n279));
  INV_X1    g0079(.A(KEYINPUT9), .ZN(new_n280));
  NOR2_X1   g0080(.A1(G20), .A2(G33), .ZN(new_n281));
  AOI22_X1  g0081(.A1(new_n203), .A2(G20), .B1(G150), .B2(new_n281), .ZN(new_n282));
  INV_X1    g0082(.A(KEYINPUT67), .ZN(new_n283));
  OAI21_X1  g0083(.A(new_n283), .B1(new_n230), .B2(new_n269), .ZN(new_n284));
  XNOR2_X1  g0084(.A(KEYINPUT64), .B(G20), .ZN(new_n285));
  NAND3_X1  g0085(.A1(new_n285), .A2(KEYINPUT67), .A3(G33), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n284), .A2(new_n286), .ZN(new_n287));
  XNOR2_X1  g0087(.A(KEYINPUT8), .B(G58), .ZN(new_n288));
  OAI21_X1  g0088(.A(new_n282), .B1(new_n287), .B2(new_n288), .ZN(new_n289));
  NAND3_X1  g0089(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n290));
  AND2_X1   g0090(.A1(new_n290), .A2(new_n231), .ZN(new_n291));
  INV_X1    g0091(.A(new_n291), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n289), .A2(new_n292), .ZN(new_n293));
  INV_X1    g0093(.A(G13), .ZN(new_n294));
  NOR2_X1   g0094(.A1(new_n294), .A2(G1), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n295), .A2(G20), .ZN(new_n296));
  INV_X1    g0096(.A(new_n296), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n297), .A2(new_n202), .ZN(new_n298));
  INV_X1    g0098(.A(KEYINPUT68), .ZN(new_n299));
  OAI21_X1  g0099(.A(new_n299), .B1(new_n292), .B2(new_n297), .ZN(new_n300));
  NAND3_X1  g0100(.A1(new_n291), .A2(new_n296), .A3(KEYINPUT68), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n259), .A2(G20), .ZN(new_n302));
  NAND3_X1  g0102(.A1(new_n300), .A2(new_n301), .A3(new_n302), .ZN(new_n303));
  OAI211_X1 g0103(.A(new_n293), .B(new_n298), .C1(new_n202), .C2(new_n303), .ZN(new_n304));
  AOI22_X1  g0104(.A1(new_n279), .A2(G190), .B1(new_n280), .B2(new_n304), .ZN(new_n305));
  INV_X1    g0105(.A(G200), .ZN(new_n306));
  OAI221_X1 g0106(.A(new_n305), .B1(new_n280), .B2(new_n304), .C1(new_n306), .C2(new_n279), .ZN(new_n307));
  XNOR2_X1  g0107(.A(new_n307), .B(KEYINPUT10), .ZN(new_n308));
  INV_X1    g0108(.A(G179), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n279), .A2(new_n309), .ZN(new_n310));
  OAI211_X1 g0110(.A(new_n310), .B(new_n304), .C1(G169), .C2(new_n279), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n308), .A2(new_n311), .ZN(new_n312));
  INV_X1    g0112(.A(new_n312), .ZN(new_n313));
  INV_X1    g0113(.A(new_n288), .ZN(new_n314));
  NOR2_X1   g0114(.A1(new_n297), .A2(new_n314), .ZN(new_n315));
  AOI21_X1  g0115(.A(new_n315), .B1(new_n303), .B2(new_n314), .ZN(new_n316));
  NOR2_X1   g0116(.A1(KEYINPUT7), .A2(G20), .ZN(new_n317));
  OAI21_X1  g0117(.A(new_n317), .B1(new_n272), .B2(new_n273), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n268), .A2(new_n270), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n319), .A2(new_n285), .ZN(new_n320));
  NAND2_X1  g0120(.A1(new_n320), .A2(KEYINPUT7), .ZN(new_n321));
  NAND3_X1  g0121(.A1(new_n318), .A2(G68), .A3(new_n321), .ZN(new_n322));
  INV_X1    g0122(.A(G58), .ZN(new_n323));
  NOR2_X1   g0123(.A1(new_n323), .A2(new_n208), .ZN(new_n324));
  OAI21_X1  g0124(.A(G20), .B1(new_n324), .B2(new_n201), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n281), .A2(G159), .ZN(new_n326));
  NAND3_X1  g0126(.A1(new_n322), .A2(new_n325), .A3(new_n326), .ZN(new_n327));
  INV_X1    g0127(.A(KEYINPUT16), .ZN(new_n328));
  AOI21_X1  g0128(.A(new_n291), .B1(new_n327), .B2(new_n328), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n325), .A2(new_n326), .ZN(new_n330));
  OAI21_X1  g0130(.A(KEYINPUT74), .B1(new_n269), .B2(KEYINPUT3), .ZN(new_n331));
  INV_X1    g0131(.A(KEYINPUT74), .ZN(new_n332));
  NAND3_X1  g0132(.A1(new_n332), .A2(new_n267), .A3(G33), .ZN(new_n333));
  NAND3_X1  g0133(.A1(new_n331), .A2(new_n333), .A3(new_n270), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n334), .A2(new_n226), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n335), .A2(KEYINPUT7), .ZN(new_n336));
  INV_X1    g0136(.A(KEYINPUT7), .ZN(new_n337));
  AND3_X1   g0137(.A1(new_n227), .A2(new_n229), .A3(new_n337), .ZN(new_n338));
  AOI21_X1  g0138(.A(new_n208), .B1(new_n338), .B2(new_n334), .ZN(new_n339));
  AOI21_X1  g0139(.A(new_n330), .B1(new_n336), .B2(new_n339), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n340), .A2(KEYINPUT16), .ZN(new_n341));
  AOI21_X1  g0141(.A(new_n316), .B1(new_n329), .B2(new_n341), .ZN(new_n342));
  OR2_X1    g0142(.A1(G223), .A2(G1698), .ZN(new_n343));
  OAI21_X1  g0143(.A(new_n343), .B1(G226), .B2(new_n275), .ZN(new_n344));
  OAI22_X1  g0144(.A1(new_n334), .A2(new_n344), .B1(new_n269), .B2(new_n210), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n345), .A2(new_n263), .ZN(new_n346));
  INV_X1    g0146(.A(KEYINPUT75), .ZN(new_n347));
  AOI21_X1  g0147(.A(new_n262), .B1(new_n265), .B2(G232), .ZN(new_n348));
  NAND4_X1  g0148(.A1(new_n346), .A2(new_n347), .A3(new_n309), .A4(new_n348), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n346), .A2(new_n348), .ZN(new_n350));
  OAI21_X1  g0150(.A(KEYINPUT75), .B1(new_n350), .B2(G179), .ZN(new_n351));
  AOI21_X1  g0151(.A(G169), .B1(new_n346), .B2(new_n348), .ZN(new_n352));
  OAI21_X1  g0152(.A(new_n349), .B1(new_n351), .B2(new_n352), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n353), .A2(KEYINPUT76), .ZN(new_n354));
  INV_X1    g0154(.A(KEYINPUT76), .ZN(new_n355));
  OAI211_X1 g0155(.A(new_n355), .B(new_n349), .C1(new_n351), .C2(new_n352), .ZN(new_n356));
  AOI21_X1  g0156(.A(new_n342), .B1(new_n354), .B2(new_n356), .ZN(new_n357));
  INV_X1    g0157(.A(new_n357), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n358), .A2(KEYINPUT18), .ZN(new_n359));
  INV_X1    g0159(.A(KEYINPUT18), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n357), .A2(new_n360), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n319), .A2(KEYINPUT66), .ZN(new_n362));
  NAND3_X1  g0162(.A1(new_n268), .A2(new_n270), .A3(new_n271), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n362), .A2(new_n363), .ZN(new_n364));
  AOI22_X1  g0164(.A1(new_n364), .A2(new_n317), .B1(KEYINPUT7), .B2(new_n320), .ZN(new_n365));
  AOI21_X1  g0165(.A(new_n330), .B1(new_n365), .B2(G68), .ZN(new_n366));
  OAI211_X1 g0166(.A(new_n341), .B(new_n292), .C1(new_n366), .C2(KEYINPUT16), .ZN(new_n367));
  INV_X1    g0167(.A(new_n316), .ZN(new_n368));
  AOI21_X1  g0168(.A(new_n306), .B1(new_n346), .B2(new_n348), .ZN(new_n369));
  INV_X1    g0169(.A(new_n350), .ZN(new_n370));
  AOI21_X1  g0170(.A(new_n369), .B1(new_n370), .B2(G190), .ZN(new_n371));
  NAND3_X1  g0171(.A1(new_n367), .A2(new_n368), .A3(new_n371), .ZN(new_n372));
  XNOR2_X1  g0172(.A(new_n372), .B(KEYINPUT17), .ZN(new_n373));
  NAND3_X1  g0173(.A1(new_n359), .A2(new_n361), .A3(new_n373), .ZN(new_n374));
  INV_X1    g0174(.A(new_n374), .ZN(new_n375));
  NOR2_X1   g0175(.A1(G226), .A2(G1698), .ZN(new_n376));
  AOI21_X1  g0176(.A(new_n376), .B1(new_n245), .B2(G1698), .ZN(new_n377));
  NAND3_X1  g0177(.A1(new_n362), .A2(new_n363), .A3(new_n377), .ZN(new_n378));
  NAND2_X1  g0178(.A1(G33), .A2(G97), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n378), .A2(new_n379), .ZN(new_n380));
  INV_X1    g0180(.A(KEYINPUT72), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n380), .A2(new_n381), .ZN(new_n382));
  NAND3_X1  g0182(.A1(new_n378), .A2(KEYINPUT72), .A3(new_n379), .ZN(new_n383));
  NAND3_X1  g0183(.A1(new_n382), .A2(new_n263), .A3(new_n383), .ZN(new_n384));
  INV_X1    g0184(.A(KEYINPUT13), .ZN(new_n385));
  AOI21_X1  g0185(.A(new_n262), .B1(new_n265), .B2(G238), .ZN(new_n386));
  NAND3_X1  g0186(.A1(new_n384), .A2(new_n385), .A3(new_n386), .ZN(new_n387));
  INV_X1    g0187(.A(new_n387), .ZN(new_n388));
  AOI21_X1  g0188(.A(new_n385), .B1(new_n384), .B2(new_n386), .ZN(new_n389));
  NOR2_X1   g0189(.A1(new_n388), .A2(new_n389), .ZN(new_n390));
  NAND2_X1  g0190(.A1(new_n390), .A2(G190), .ZN(new_n391));
  INV_X1    g0191(.A(new_n389), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n392), .A2(new_n387), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n393), .A2(G200), .ZN(new_n394));
  NAND3_X1  g0194(.A1(new_n284), .A2(G77), .A3(new_n286), .ZN(new_n395));
  AOI22_X1  g0195(.A1(new_n281), .A2(G50), .B1(G20), .B2(new_n208), .ZN(new_n396));
  AOI21_X1  g0196(.A(new_n291), .B1(new_n395), .B2(new_n396), .ZN(new_n397));
  OR2_X1    g0197(.A1(new_n397), .A2(KEYINPUT11), .ZN(new_n398));
  NAND3_X1  g0198(.A1(new_n291), .A2(G68), .A3(new_n302), .ZN(new_n399));
  INV_X1    g0199(.A(KEYINPUT12), .ZN(new_n400));
  AOI21_X1  g0200(.A(new_n400), .B1(new_n297), .B2(new_n208), .ZN(new_n401));
  NOR3_X1   g0201(.A1(new_n296), .A2(KEYINPUT12), .A3(G68), .ZN(new_n402));
  OAI21_X1  g0202(.A(new_n399), .B1(new_n401), .B2(new_n402), .ZN(new_n403));
  AOI21_X1  g0203(.A(new_n403), .B1(new_n397), .B2(KEYINPUT11), .ZN(new_n404));
  AND2_X1   g0204(.A1(new_n398), .A2(new_n404), .ZN(new_n405));
  NAND3_X1  g0205(.A1(new_n391), .A2(new_n394), .A3(new_n405), .ZN(new_n406));
  INV_X1    g0206(.A(new_n406), .ZN(new_n407));
  OAI22_X1  g0207(.A1(new_n393), .A2(new_n309), .B1(KEYINPUT73), .B2(KEYINPUT14), .ZN(new_n408));
  NAND2_X1  g0208(.A1(KEYINPUT73), .A2(KEYINPUT14), .ZN(new_n409));
  INV_X1    g0209(.A(G169), .ZN(new_n410));
  OAI21_X1  g0210(.A(new_n409), .B1(new_n390), .B2(new_n410), .ZN(new_n411));
  NAND4_X1  g0211(.A1(new_n393), .A2(KEYINPUT73), .A3(KEYINPUT14), .A4(G169), .ZN(new_n412));
  AOI21_X1  g0212(.A(new_n408), .B1(new_n411), .B2(new_n412), .ZN(new_n413));
  INV_X1    g0213(.A(new_n413), .ZN(new_n414));
  INV_X1    g0214(.A(new_n405), .ZN(new_n415));
  AOI21_X1  g0215(.A(new_n407), .B1(new_n414), .B2(new_n415), .ZN(new_n416));
  XNOR2_X1  g0216(.A(KEYINPUT15), .B(G87), .ZN(new_n417));
  XNOR2_X1  g0217(.A(new_n417), .B(KEYINPUT70), .ZN(new_n418));
  NAND3_X1  g0218(.A1(new_n418), .A2(new_n284), .A3(new_n286), .ZN(new_n419));
  AOI22_X1  g0219(.A1(new_n314), .A2(new_n281), .B1(new_n230), .B2(G77), .ZN(new_n420));
  AOI21_X1  g0220(.A(new_n291), .B1(new_n419), .B2(new_n420), .ZN(new_n421));
  NAND3_X1  g0221(.A1(new_n291), .A2(G77), .A3(new_n302), .ZN(new_n422));
  OAI21_X1  g0222(.A(new_n422), .B1(G77), .B2(new_n296), .ZN(new_n423));
  NOR2_X1   g0223(.A1(new_n421), .A2(new_n423), .ZN(new_n424));
  INV_X1    g0224(.A(new_n424), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n425), .A2(KEYINPUT71), .ZN(new_n426));
  INV_X1    g0226(.A(KEYINPUT71), .ZN(new_n427));
  INV_X1    g0227(.A(G41), .ZN(new_n428));
  OAI21_X1  g0228(.A(new_n232), .B1(new_n269), .B2(new_n428), .ZN(new_n429));
  AOI21_X1  g0229(.A(new_n429), .B1(new_n364), .B2(new_n216), .ZN(new_n430));
  NOR2_X1   g0230(.A1(G232), .A2(G1698), .ZN(new_n431));
  AOI21_X1  g0231(.A(new_n431), .B1(new_n209), .B2(G1698), .ZN(new_n432));
  OAI21_X1  g0232(.A(new_n430), .B1(new_n364), .B2(new_n432), .ZN(new_n433));
  AOI21_X1  g0233(.A(new_n262), .B1(new_n265), .B2(G244), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n433), .A2(new_n434), .ZN(new_n435));
  AOI22_X1  g0235(.A1(new_n424), .A2(new_n427), .B1(G200), .B2(new_n435), .ZN(new_n436));
  NAND4_X1  g0236(.A1(new_n433), .A2(KEYINPUT69), .A3(G190), .A4(new_n434), .ZN(new_n437));
  INV_X1    g0237(.A(KEYINPUT69), .ZN(new_n438));
  INV_X1    g0238(.A(G190), .ZN(new_n439));
  OAI21_X1  g0239(.A(new_n438), .B1(new_n435), .B2(new_n439), .ZN(new_n440));
  NAND4_X1  g0240(.A1(new_n426), .A2(new_n436), .A3(new_n437), .A4(new_n440), .ZN(new_n441));
  NAND2_X1  g0241(.A1(new_n435), .A2(new_n410), .ZN(new_n442));
  OAI211_X1 g0242(.A(new_n425), .B(new_n442), .C1(G179), .C2(new_n435), .ZN(new_n443));
  AND2_X1   g0243(.A1(new_n441), .A2(new_n443), .ZN(new_n444));
  NAND4_X1  g0244(.A1(new_n313), .A2(new_n375), .A3(new_n416), .A4(new_n444), .ZN(new_n445));
  INV_X1    g0245(.A(new_n445), .ZN(new_n446));
  INV_X1    g0246(.A(G303), .ZN(new_n447));
  AOI21_X1  g0247(.A(new_n447), .B1(new_n362), .B2(new_n363), .ZN(new_n448));
  NAND4_X1  g0248(.A1(new_n331), .A2(new_n333), .A3(new_n275), .A4(new_n270), .ZN(new_n449));
  NOR2_X1   g0249(.A1(new_n449), .A2(new_n223), .ZN(new_n450));
  NOR2_X1   g0250(.A1(new_n448), .A2(new_n450), .ZN(new_n451));
  AND2_X1   g0251(.A1(G264), .A2(G1698), .ZN(new_n452));
  NAND4_X1  g0252(.A1(new_n331), .A2(new_n333), .A3(new_n270), .A4(new_n452), .ZN(new_n453));
  INV_X1    g0253(.A(KEYINPUT81), .ZN(new_n454));
  XNOR2_X1  g0254(.A(new_n453), .B(new_n454), .ZN(new_n455));
  AOI21_X1  g0255(.A(new_n429), .B1(new_n451), .B2(new_n455), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n428), .A2(KEYINPUT5), .ZN(new_n457));
  OR2_X1    g0257(.A1(new_n457), .A2(KEYINPUT77), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n457), .A2(KEYINPUT77), .ZN(new_n459));
  INV_X1    g0259(.A(G45), .ZN(new_n460));
  NOR2_X1   g0260(.A1(new_n460), .A2(G1), .ZN(new_n461));
  INV_X1    g0261(.A(KEYINPUT5), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n462), .A2(G41), .ZN(new_n463));
  NAND4_X1  g0263(.A1(new_n458), .A2(new_n459), .A3(new_n461), .A4(new_n463), .ZN(new_n464));
  NAND2_X1  g0264(.A1(new_n429), .A2(G274), .ZN(new_n465));
  NAND3_X1  g0265(.A1(new_n461), .A2(new_n457), .A3(new_n463), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n466), .A2(new_n429), .ZN(new_n467));
  INV_X1    g0267(.A(G270), .ZN(new_n468));
  OAI22_X1  g0268(.A1(new_n464), .A2(new_n465), .B1(new_n467), .B2(new_n468), .ZN(new_n469));
  OAI21_X1  g0269(.A(KEYINPUT82), .B1(new_n456), .B2(new_n469), .ZN(new_n470));
  OAI22_X1  g0270(.A1(new_n274), .A2(new_n447), .B1(new_n223), .B2(new_n449), .ZN(new_n471));
  XNOR2_X1  g0271(.A(new_n453), .B(KEYINPUT81), .ZN(new_n472));
  OAI21_X1  g0272(.A(new_n263), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  INV_X1    g0273(.A(KEYINPUT82), .ZN(new_n474));
  INV_X1    g0274(.A(new_n469), .ZN(new_n475));
  NAND3_X1  g0275(.A1(new_n473), .A2(new_n474), .A3(new_n475), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n470), .A2(new_n476), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n477), .A2(G190), .ZN(new_n478));
  INV_X1    g0278(.A(G116), .ZN(new_n479));
  AOI21_X1  g0279(.A(new_n291), .B1(G20), .B2(new_n479), .ZN(new_n480));
  INV_X1    g0280(.A(KEYINPUT84), .ZN(new_n481));
  NAND2_X1  g0281(.A1(G33), .A2(G283), .ZN(new_n482));
  INV_X1    g0282(.A(G97), .ZN(new_n483));
  OAI21_X1  g0283(.A(new_n482), .B1(new_n483), .B2(G33), .ZN(new_n484));
  INV_X1    g0284(.A(new_n484), .ZN(new_n485));
  AOI21_X1  g0285(.A(new_n481), .B1(new_n485), .B2(new_n285), .ZN(new_n486));
  NOR3_X1   g0286(.A1(new_n230), .A2(new_n484), .A3(KEYINPUT84), .ZN(new_n487));
  OAI21_X1  g0287(.A(new_n480), .B1(new_n486), .B2(new_n487), .ZN(new_n488));
  INV_X1    g0288(.A(KEYINPUT20), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  OAI211_X1 g0290(.A(KEYINPUT20), .B(new_n480), .C1(new_n486), .C2(new_n487), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n259), .A2(G33), .ZN(new_n493));
  NAND3_X1  g0293(.A1(new_n291), .A2(new_n296), .A3(new_n493), .ZN(new_n494));
  INV_X1    g0294(.A(new_n494), .ZN(new_n495));
  NAND3_X1  g0295(.A1(new_n297), .A2(KEYINPUT83), .A3(new_n479), .ZN(new_n496));
  INV_X1    g0296(.A(KEYINPUT83), .ZN(new_n497));
  OAI21_X1  g0297(.A(new_n497), .B1(new_n296), .B2(G116), .ZN(new_n498));
  AOI22_X1  g0298(.A1(G116), .A2(new_n495), .B1(new_n496), .B2(new_n498), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n492), .A2(new_n499), .ZN(new_n500));
  INV_X1    g0300(.A(new_n500), .ZN(new_n501));
  OAI211_X1 g0301(.A(new_n478), .B(new_n501), .C1(new_n306), .C2(new_n477), .ZN(new_n502));
  AOI21_X1  g0302(.A(new_n410), .B1(new_n492), .B2(new_n499), .ZN(new_n503));
  NAND3_X1  g0303(.A1(new_n503), .A2(new_n470), .A3(new_n476), .ZN(new_n504));
  INV_X1    g0304(.A(KEYINPUT21), .ZN(new_n505));
  NOR3_X1   g0305(.A1(new_n456), .A2(new_n309), .A3(new_n469), .ZN(new_n506));
  AOI22_X1  g0306(.A1(new_n504), .A2(new_n505), .B1(new_n500), .B2(new_n506), .ZN(new_n507));
  NAND4_X1  g0307(.A1(new_n503), .A2(new_n470), .A3(KEYINPUT21), .A4(new_n476), .ZN(new_n508));
  AND3_X1   g0308(.A1(new_n502), .A2(new_n507), .A3(new_n508), .ZN(new_n509));
  NOR2_X1   g0309(.A1(new_n418), .A2(new_n296), .ZN(new_n510));
  INV_X1    g0310(.A(new_n510), .ZN(new_n511));
  INV_X1    g0311(.A(KEYINPUT70), .ZN(new_n512));
  XNOR2_X1  g0312(.A(new_n417), .B(new_n512), .ZN(new_n513));
  NOR3_X1   g0313(.A1(new_n513), .A2(KEYINPUT80), .A3(new_n494), .ZN(new_n514));
  INV_X1    g0314(.A(KEYINPUT80), .ZN(new_n515));
  AOI21_X1  g0315(.A(new_n515), .B1(new_n418), .B2(new_n495), .ZN(new_n516));
  NOR2_X1   g0316(.A1(new_n514), .A2(new_n516), .ZN(new_n517));
  INV_X1    g0317(.A(KEYINPUT19), .ZN(new_n518));
  OAI21_X1  g0318(.A(new_n518), .B1(new_n287), .B2(new_n483), .ZN(new_n519));
  NOR2_X1   g0319(.A1(new_n334), .A2(new_n230), .ZN(new_n520));
  XOR2_X1   g0320(.A(KEYINPUT79), .B(G87), .Z(new_n521));
  NOR2_X1   g0321(.A1(G97), .A2(G107), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  OAI21_X1  g0323(.A(new_n285), .B1(new_n518), .B2(new_n379), .ZN(new_n524));
  AOI22_X1  g0324(.A1(new_n520), .A2(G68), .B1(new_n523), .B2(new_n524), .ZN(new_n525));
  AND2_X1   g0325(.A1(new_n519), .A2(new_n525), .ZN(new_n526));
  OAI211_X1 g0326(.A(new_n511), .B(new_n517), .C1(new_n526), .C2(new_n291), .ZN(new_n527));
  NAND2_X1  g0327(.A1(G33), .A2(G116), .ZN(new_n528));
  OAI21_X1  g0328(.A(new_n528), .B1(new_n449), .B2(new_n209), .ZN(new_n529));
  NAND4_X1  g0329(.A1(new_n331), .A2(new_n333), .A3(G244), .A4(new_n270), .ZN(new_n530));
  NOR2_X1   g0330(.A1(new_n530), .A2(new_n275), .ZN(new_n531));
  OAI21_X1  g0331(.A(new_n263), .B1(new_n529), .B2(new_n531), .ZN(new_n532));
  NOR3_X1   g0332(.A1(new_n263), .A2(new_n211), .A3(new_n461), .ZN(new_n533));
  AOI21_X1  g0333(.A(new_n533), .B1(G274), .B2(new_n461), .ZN(new_n534));
  NAND2_X1  g0334(.A1(new_n532), .A2(new_n534), .ZN(new_n535));
  INV_X1    g0335(.A(KEYINPUT78), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  NAND3_X1  g0337(.A1(new_n532), .A2(KEYINPUT78), .A3(new_n534), .ZN(new_n538));
  NAND3_X1  g0338(.A1(new_n537), .A2(new_n309), .A3(new_n538), .ZN(new_n539));
  INV_X1    g0339(.A(new_n538), .ZN(new_n540));
  AOI21_X1  g0340(.A(KEYINPUT78), .B1(new_n532), .B2(new_n534), .ZN(new_n541));
  NOR2_X1   g0341(.A1(new_n540), .A2(new_n541), .ZN(new_n542));
  OAI211_X1 g0342(.A(new_n527), .B(new_n539), .C1(new_n542), .C2(G169), .ZN(new_n543));
  OAI21_X1  g0343(.A(G200), .B1(new_n540), .B2(new_n541), .ZN(new_n544));
  NAND3_X1  g0344(.A1(new_n537), .A2(G190), .A3(new_n538), .ZN(new_n545));
  AOI21_X1  g0345(.A(new_n291), .B1(new_n519), .B2(new_n525), .ZN(new_n546));
  NOR2_X1   g0346(.A1(new_n494), .A2(new_n210), .ZN(new_n547));
  NOR3_X1   g0347(.A1(new_n546), .A2(new_n510), .A3(new_n547), .ZN(new_n548));
  NAND3_X1  g0348(.A1(new_n544), .A2(new_n545), .A3(new_n548), .ZN(new_n549));
  AND2_X1   g0349(.A1(new_n543), .A2(new_n549), .ZN(new_n550));
  OAI22_X1  g0350(.A1(new_n464), .A2(new_n465), .B1(new_n467), .B2(new_n223), .ZN(new_n551));
  NAND4_X1  g0351(.A1(new_n362), .A2(G250), .A3(G1698), .A4(new_n363), .ZN(new_n552));
  INV_X1    g0352(.A(KEYINPUT4), .ZN(new_n553));
  NOR2_X1   g0353(.A1(new_n553), .A2(new_n215), .ZN(new_n554));
  NAND4_X1  g0354(.A1(new_n362), .A2(new_n275), .A3(new_n363), .A4(new_n554), .ZN(new_n555));
  OAI21_X1  g0355(.A(new_n553), .B1(new_n530), .B2(G1698), .ZN(new_n556));
  NAND4_X1  g0356(.A1(new_n552), .A2(new_n555), .A3(new_n556), .A4(new_n482), .ZN(new_n557));
  AOI21_X1  g0357(.A(new_n551), .B1(new_n557), .B2(new_n263), .ZN(new_n558));
  NOR2_X1   g0358(.A1(new_n558), .A2(G169), .ZN(new_n559));
  AOI211_X1 g0359(.A(G179), .B(new_n551), .C1(new_n557), .C2(new_n263), .ZN(new_n560));
  NOR2_X1   g0360(.A1(new_n296), .A2(G97), .ZN(new_n561));
  AOI21_X1  g0361(.A(new_n561), .B1(new_n495), .B2(G97), .ZN(new_n562));
  INV_X1    g0362(.A(new_n562), .ZN(new_n563));
  NAND3_X1  g0363(.A1(new_n318), .A2(G107), .A3(new_n321), .ZN(new_n564));
  INV_X1    g0364(.A(KEYINPUT6), .ZN(new_n565));
  NOR3_X1   g0365(.A1(new_n565), .A2(new_n483), .A3(G107), .ZN(new_n566));
  AOI21_X1  g0366(.A(new_n566), .B1(new_n565), .B2(new_n256), .ZN(new_n567));
  INV_X1    g0367(.A(new_n567), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n568), .A2(new_n230), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n281), .A2(G77), .ZN(new_n570));
  NAND3_X1  g0370(.A1(new_n564), .A2(new_n569), .A3(new_n570), .ZN(new_n571));
  AOI21_X1  g0371(.A(new_n563), .B1(new_n571), .B2(new_n292), .ZN(new_n572));
  NOR3_X1   g0372(.A1(new_n559), .A2(new_n560), .A3(new_n572), .ZN(new_n573));
  INV_X1    g0373(.A(new_n573), .ZN(new_n574));
  OAI21_X1  g0374(.A(new_n570), .B1(new_n567), .B2(new_n285), .ZN(new_n575));
  AOI21_X1  g0375(.A(new_n575), .B1(new_n365), .B2(G107), .ZN(new_n576));
  OAI21_X1  g0376(.A(new_n562), .B1(new_n576), .B2(new_n291), .ZN(new_n577));
  INV_X1    g0377(.A(new_n558), .ZN(new_n578));
  AOI21_X1  g0378(.A(new_n577), .B1(G200), .B2(new_n578), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n558), .A2(G190), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n574), .A2(new_n581), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n223), .A2(G1698), .ZN(new_n583));
  OAI21_X1  g0383(.A(new_n583), .B1(G250), .B2(G1698), .ZN(new_n584));
  INV_X1    g0384(.A(G294), .ZN(new_n585));
  OAI22_X1  g0385(.A1(new_n334), .A2(new_n584), .B1(new_n269), .B2(new_n585), .ZN(new_n586));
  INV_X1    g0386(.A(KEYINPUT87), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n586), .A2(new_n587), .ZN(new_n588));
  OAI221_X1 g0388(.A(KEYINPUT87), .B1(new_n269), .B2(new_n585), .C1(new_n334), .C2(new_n584), .ZN(new_n589));
  NAND3_X1  g0389(.A1(new_n588), .A2(new_n263), .A3(new_n589), .ZN(new_n590));
  NAND3_X1  g0390(.A1(new_n466), .A2(new_n429), .A3(G264), .ZN(new_n591));
  AND2_X1   g0391(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  OR2_X1    g0392(.A1(new_n464), .A2(new_n465), .ZN(new_n593));
  NAND3_X1  g0393(.A1(new_n592), .A2(new_n309), .A3(new_n593), .ZN(new_n594));
  NAND3_X1  g0394(.A1(new_n590), .A2(new_n593), .A3(new_n591), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n595), .A2(new_n410), .ZN(new_n596));
  NOR2_X1   g0396(.A1(KEYINPUT23), .A2(G107), .ZN(new_n597));
  INV_X1    g0397(.A(new_n597), .ZN(new_n598));
  INV_X1    g0398(.A(KEYINPUT23), .ZN(new_n599));
  AOI21_X1  g0399(.A(new_n599), .B1(G20), .B2(new_n216), .ZN(new_n600));
  INV_X1    g0400(.A(KEYINPUT85), .ZN(new_n601));
  OAI22_X1  g0401(.A1(new_n285), .A2(new_n598), .B1(new_n600), .B2(new_n601), .ZN(new_n602));
  OAI21_X1  g0402(.A(KEYINPUT23), .B1(new_n226), .B2(G107), .ZN(new_n603));
  OAI22_X1  g0403(.A1(new_n603), .A2(KEYINPUT85), .B1(G20), .B2(new_n528), .ZN(new_n604));
  OAI21_X1  g0404(.A(KEYINPUT86), .B1(new_n602), .B2(new_n604), .ZN(new_n605));
  AOI22_X1  g0405(.A1(new_n230), .A2(new_n597), .B1(KEYINPUT85), .B2(new_n603), .ZN(new_n606));
  INV_X1    g0406(.A(KEYINPUT86), .ZN(new_n607));
  NOR2_X1   g0407(.A1(new_n528), .A2(G20), .ZN(new_n608));
  AOI21_X1  g0408(.A(new_n608), .B1(new_n600), .B2(new_n601), .ZN(new_n609));
  NAND3_X1  g0409(.A1(new_n606), .A2(new_n607), .A3(new_n609), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n605), .A2(new_n610), .ZN(new_n611));
  AND3_X1   g0411(.A1(new_n227), .A2(new_n229), .A3(G87), .ZN(new_n612));
  NAND3_X1  g0412(.A1(new_n362), .A2(new_n612), .A3(new_n363), .ZN(new_n613));
  INV_X1    g0413(.A(KEYINPUT22), .ZN(new_n614));
  NOR2_X1   g0414(.A1(new_n614), .A2(new_n210), .ZN(new_n615));
  AOI22_X1  g0415(.A1(new_n613), .A2(new_n614), .B1(new_n520), .B2(new_n615), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n611), .A2(new_n616), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n617), .A2(KEYINPUT24), .ZN(new_n618));
  INV_X1    g0418(.A(KEYINPUT24), .ZN(new_n619));
  NAND3_X1  g0419(.A1(new_n611), .A2(new_n616), .A3(new_n619), .ZN(new_n620));
  AOI21_X1  g0420(.A(new_n291), .B1(new_n618), .B2(new_n620), .ZN(new_n621));
  AOI21_X1  g0421(.A(KEYINPUT25), .B1(new_n297), .B2(new_n216), .ZN(new_n622));
  INV_X1    g0422(.A(new_n622), .ZN(new_n623));
  NAND3_X1  g0423(.A1(new_n297), .A2(KEYINPUT25), .A3(new_n216), .ZN(new_n624));
  AOI22_X1  g0424(.A1(new_n623), .A2(new_n624), .B1(new_n495), .B2(G107), .ZN(new_n625));
  INV_X1    g0425(.A(new_n625), .ZN(new_n626));
  OAI211_X1 g0426(.A(new_n594), .B(new_n596), .C1(new_n621), .C2(new_n626), .ZN(new_n627));
  INV_X1    g0427(.A(new_n627), .ZN(new_n628));
  AND3_X1   g0428(.A1(new_n611), .A2(new_n616), .A3(new_n619), .ZN(new_n629));
  AOI21_X1  g0429(.A(new_n619), .B1(new_n611), .B2(new_n616), .ZN(new_n630));
  OAI21_X1  g0430(.A(new_n292), .B1(new_n629), .B2(new_n630), .ZN(new_n631));
  NAND4_X1  g0431(.A1(new_n590), .A2(G190), .A3(new_n593), .A4(new_n591), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n595), .A2(G200), .ZN(new_n633));
  NAND4_X1  g0433(.A1(new_n631), .A2(new_n632), .A3(new_n625), .A4(new_n633), .ZN(new_n634));
  INV_X1    g0434(.A(new_n634), .ZN(new_n635));
  NOR3_X1   g0435(.A1(new_n582), .A2(new_n628), .A3(new_n635), .ZN(new_n636));
  AND4_X1   g0436(.A1(new_n446), .A2(new_n509), .A3(new_n550), .A4(new_n636), .ZN(G372));
  NAND2_X1  g0437(.A1(new_n406), .A2(new_n373), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n414), .A2(new_n415), .ZN(new_n639));
  AOI21_X1  g0439(.A(new_n638), .B1(new_n639), .B2(new_n443), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n359), .A2(new_n361), .ZN(new_n641));
  OAI21_X1  g0441(.A(new_n308), .B1(new_n640), .B2(new_n641), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n642), .A2(new_n311), .ZN(new_n643));
  INV_X1    g0443(.A(new_n643), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n504), .A2(new_n505), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n506), .A2(new_n500), .ZN(new_n646));
  NAND4_X1  g0446(.A1(new_n627), .A2(new_n645), .A3(new_n508), .A4(new_n646), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n535), .A2(new_n410), .ZN(new_n648));
  NAND3_X1  g0448(.A1(new_n527), .A2(new_n539), .A3(new_n648), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n535), .A2(G200), .ZN(new_n650));
  NAND3_X1  g0450(.A1(new_n545), .A2(new_n548), .A3(new_n650), .ZN(new_n651));
  AND3_X1   g0451(.A1(new_n634), .A2(new_n649), .A3(new_n651), .ZN(new_n652));
  AOI21_X1  g0452(.A(new_n573), .B1(new_n580), .B2(new_n579), .ZN(new_n653));
  NAND3_X1  g0453(.A1(new_n647), .A2(new_n652), .A3(new_n653), .ZN(new_n654));
  AND2_X1   g0454(.A1(new_n649), .A2(new_n651), .ZN(new_n655));
  INV_X1    g0455(.A(KEYINPUT26), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n558), .A2(new_n309), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n657), .A2(new_n577), .ZN(new_n658));
  OAI21_X1  g0458(.A(KEYINPUT88), .B1(new_n658), .B2(new_n559), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n578), .A2(new_n410), .ZN(new_n660));
  INV_X1    g0460(.A(KEYINPUT88), .ZN(new_n661));
  NAND4_X1  g0461(.A1(new_n660), .A2(new_n661), .A3(new_n657), .A4(new_n577), .ZN(new_n662));
  NAND4_X1  g0462(.A1(new_n655), .A2(new_n656), .A3(new_n659), .A4(new_n662), .ZN(new_n663));
  NAND3_X1  g0463(.A1(new_n543), .A2(new_n549), .A3(new_n573), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n664), .A2(KEYINPUT26), .ZN(new_n665));
  NAND4_X1  g0465(.A1(new_n654), .A2(new_n649), .A3(new_n663), .A4(new_n665), .ZN(new_n666));
  INV_X1    g0466(.A(new_n666), .ZN(new_n667));
  OAI21_X1  g0467(.A(new_n644), .B1(new_n445), .B2(new_n667), .ZN(G369));
  NAND2_X1  g0468(.A1(new_n507), .A2(new_n508), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n285), .A2(new_n295), .ZN(new_n670));
  OAI21_X1  g0470(.A(G213), .B1(new_n670), .B2(KEYINPUT27), .ZN(new_n671));
  AOI21_X1  g0471(.A(new_n671), .B1(KEYINPUT27), .B2(new_n670), .ZN(new_n672));
  XNOR2_X1  g0472(.A(new_n672), .B(KEYINPUT89), .ZN(new_n673));
  INV_X1    g0473(.A(G343), .ZN(new_n674));
  NOR2_X1   g0474(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  INV_X1    g0475(.A(new_n675), .ZN(new_n676));
  NOR2_X1   g0476(.A1(new_n676), .A2(new_n501), .ZN(new_n677));
  MUX2_X1   g0477(.A(new_n509), .B(new_n669), .S(new_n677), .Z(new_n678));
  NAND2_X1  g0478(.A1(new_n678), .A2(G330), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n631), .A2(new_n625), .ZN(new_n680));
  AND2_X1   g0480(.A1(new_n680), .A2(new_n675), .ZN(new_n681));
  OAI21_X1  g0481(.A(new_n627), .B1(new_n681), .B2(new_n635), .ZN(new_n682));
  NOR2_X1   g0482(.A1(new_n627), .A2(new_n675), .ZN(new_n683));
  INV_X1    g0483(.A(new_n683), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n682), .A2(new_n684), .ZN(new_n685));
  NOR2_X1   g0485(.A1(new_n679), .A2(new_n685), .ZN(new_n686));
  INV_X1    g0486(.A(new_n686), .ZN(new_n687));
  AOI21_X1  g0487(.A(new_n675), .B1(new_n507), .B2(new_n508), .ZN(new_n688));
  NAND3_X1  g0488(.A1(new_n682), .A2(new_n684), .A3(new_n688), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n689), .A2(new_n684), .ZN(new_n690));
  INV_X1    g0490(.A(KEYINPUT90), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  INV_X1    g0492(.A(new_n692), .ZN(new_n693));
  NOR2_X1   g0493(.A1(new_n690), .A2(new_n691), .ZN(new_n694));
  OAI21_X1  g0494(.A(new_n687), .B1(new_n693), .B2(new_n694), .ZN(G399));
  NOR2_X1   g0495(.A1(new_n222), .A2(G41), .ZN(new_n696));
  INV_X1    g0496(.A(new_n696), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n697), .A2(G1), .ZN(new_n698));
  NAND3_X1  g0498(.A1(new_n521), .A2(new_n479), .A3(new_n522), .ZN(new_n699));
  OAI22_X1  g0499(.A1(new_n698), .A2(new_n699), .B1(new_n235), .B2(new_n697), .ZN(new_n700));
  XOR2_X1   g0500(.A(KEYINPUT91), .B(KEYINPUT28), .Z(new_n701));
  XNOR2_X1  g0501(.A(new_n700), .B(new_n701), .ZN(new_n702));
  NAND3_X1  g0502(.A1(new_n550), .A2(new_n656), .A3(new_n573), .ZN(new_n703));
  NAND4_X1  g0503(.A1(new_n659), .A2(new_n662), .A3(new_n649), .A4(new_n651), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n704), .A2(KEYINPUT26), .ZN(new_n705));
  NAND3_X1  g0505(.A1(new_n703), .A2(new_n705), .A3(new_n649), .ZN(new_n706));
  NAND2_X1  g0506(.A1(new_n647), .A2(new_n652), .ZN(new_n707));
  INV_X1    g0507(.A(new_n707), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n582), .A2(KEYINPUT92), .ZN(new_n709));
  INV_X1    g0509(.A(KEYINPUT92), .ZN(new_n710));
  NAND3_X1  g0510(.A1(new_n574), .A2(new_n581), .A3(new_n710), .ZN(new_n711));
  NAND4_X1  g0511(.A1(new_n708), .A2(KEYINPUT93), .A3(new_n709), .A4(new_n711), .ZN(new_n712));
  INV_X1    g0512(.A(KEYINPUT93), .ZN(new_n713));
  NAND2_X1  g0513(.A1(new_n709), .A2(new_n711), .ZN(new_n714));
  OAI21_X1  g0514(.A(new_n713), .B1(new_n714), .B2(new_n707), .ZN(new_n715));
  AOI21_X1  g0515(.A(new_n706), .B1(new_n712), .B2(new_n715), .ZN(new_n716));
  OAI21_X1  g0516(.A(KEYINPUT29), .B1(new_n716), .B2(new_n675), .ZN(new_n717));
  NOR2_X1   g0517(.A1(new_n667), .A2(new_n675), .ZN(new_n718));
  INV_X1    g0518(.A(KEYINPUT29), .ZN(new_n719));
  NAND2_X1  g0519(.A1(new_n718), .A2(new_n719), .ZN(new_n720));
  NAND4_X1  g0520(.A1(new_n509), .A2(new_n636), .A3(new_n550), .A4(new_n676), .ZN(new_n721));
  AND2_X1   g0521(.A1(new_n506), .A2(new_n592), .ZN(new_n722));
  NAND4_X1  g0522(.A1(new_n722), .A2(KEYINPUT30), .A3(new_n542), .A4(new_n558), .ZN(new_n723));
  INV_X1    g0523(.A(KEYINPUT30), .ZN(new_n724));
  NAND3_X1  g0524(.A1(new_n506), .A2(new_n558), .A3(new_n592), .ZN(new_n725));
  INV_X1    g0525(.A(new_n542), .ZN(new_n726));
  OAI21_X1  g0526(.A(new_n724), .B1(new_n725), .B2(new_n726), .ZN(new_n727));
  NAND4_X1  g0527(.A1(new_n578), .A2(new_n309), .A3(new_n535), .A4(new_n595), .ZN(new_n728));
  OAI211_X1 g0528(.A(new_n723), .B(new_n727), .C1(new_n477), .C2(new_n728), .ZN(new_n729));
  NAND2_X1  g0529(.A1(new_n729), .A2(new_n675), .ZN(new_n730));
  INV_X1    g0530(.A(KEYINPUT31), .ZN(new_n731));
  NAND2_X1  g0531(.A1(new_n730), .A2(new_n731), .ZN(new_n732));
  NAND3_X1  g0532(.A1(new_n729), .A2(KEYINPUT31), .A3(new_n675), .ZN(new_n733));
  NAND3_X1  g0533(.A1(new_n721), .A2(new_n732), .A3(new_n733), .ZN(new_n734));
  NAND2_X1  g0534(.A1(new_n734), .A2(G330), .ZN(new_n735));
  NAND3_X1  g0535(.A1(new_n717), .A2(new_n720), .A3(new_n735), .ZN(new_n736));
  OR2_X1    g0536(.A1(new_n736), .A2(KEYINPUT94), .ZN(new_n737));
  NAND2_X1  g0537(.A1(new_n736), .A2(KEYINPUT94), .ZN(new_n738));
  NAND2_X1  g0538(.A1(new_n737), .A2(new_n738), .ZN(new_n739));
  OAI21_X1  g0539(.A(new_n702), .B1(new_n739), .B2(G1), .ZN(G364));
  NOR2_X1   g0540(.A1(new_n230), .A2(new_n294), .ZN(new_n741));
  NAND2_X1  g0541(.A1(new_n741), .A2(G45), .ZN(new_n742));
  NAND2_X1  g0542(.A1(new_n742), .A2(G1), .ZN(new_n743));
  NOR2_X1   g0543(.A1(new_n743), .A2(new_n696), .ZN(new_n744));
  INV_X1    g0544(.A(new_n744), .ZN(new_n745));
  NOR2_X1   g0545(.A1(G13), .A2(G33), .ZN(new_n746));
  INV_X1    g0546(.A(new_n746), .ZN(new_n747));
  NOR2_X1   g0547(.A1(new_n747), .A2(G20), .ZN(new_n748));
  INV_X1    g0548(.A(new_n748), .ZN(new_n749));
  OR2_X1    g0549(.A1(new_n678), .A2(new_n749), .ZN(new_n750));
  AOI21_X1  g0550(.A(new_n231), .B1(G20), .B2(new_n410), .ZN(new_n751));
  NOR2_X1   g0551(.A1(new_n748), .A2(new_n751), .ZN(new_n752));
  INV_X1    g0552(.A(new_n752), .ZN(new_n753));
  OR2_X1    g0553(.A1(new_n254), .A2(new_n460), .ZN(new_n754));
  AND3_X1   g0554(.A1(new_n331), .A2(new_n333), .A3(new_n270), .ZN(new_n755));
  NOR2_X1   g0555(.A1(new_n755), .A2(new_n222), .ZN(new_n756));
  OAI211_X1 g0556(.A(new_n754), .B(new_n756), .C1(G45), .C2(new_n235), .ZN(new_n757));
  NOR2_X1   g0557(.A1(new_n364), .A2(new_n222), .ZN(new_n758));
  AOI22_X1  g0558(.A1(new_n758), .A2(G355), .B1(new_n479), .B2(new_n222), .ZN(new_n759));
  AOI21_X1  g0559(.A(new_n753), .B1(new_n757), .B2(new_n759), .ZN(new_n760));
  NOR2_X1   g0560(.A1(new_n306), .A2(G179), .ZN(new_n761));
  INV_X1    g0561(.A(new_n761), .ZN(new_n762));
  NOR3_X1   g0562(.A1(new_n285), .A2(new_n762), .A3(G190), .ZN(new_n763));
  INV_X1    g0563(.A(new_n763), .ZN(new_n764));
  INV_X1    g0564(.A(G283), .ZN(new_n765));
  NOR2_X1   g0565(.A1(new_n764), .A2(new_n765), .ZN(new_n766));
  NOR2_X1   g0566(.A1(G179), .A2(G200), .ZN(new_n767));
  AOI21_X1  g0567(.A(new_n285), .B1(G190), .B2(new_n767), .ZN(new_n768));
  NOR3_X1   g0568(.A1(new_n762), .A2(new_n226), .A3(new_n439), .ZN(new_n769));
  INV_X1    g0569(.A(new_n769), .ZN(new_n770));
  OAI221_X1 g0570(.A(new_n364), .B1(new_n768), .B2(new_n585), .C1(new_n770), .C2(new_n447), .ZN(new_n771));
  NAND3_X1  g0571(.A1(new_n230), .A2(new_n439), .A3(new_n767), .ZN(new_n772));
  INV_X1    g0572(.A(new_n772), .ZN(new_n773));
  AOI211_X1 g0573(.A(new_n766), .B(new_n771), .C1(G329), .C2(new_n773), .ZN(new_n774));
  NOR2_X1   g0574(.A1(new_n285), .A2(new_n309), .ZN(new_n775));
  NAND2_X1  g0575(.A1(new_n775), .A2(G190), .ZN(new_n776));
  NOR2_X1   g0576(.A1(new_n776), .A2(new_n306), .ZN(new_n777));
  INV_X1    g0577(.A(new_n777), .ZN(new_n778));
  INV_X1    g0578(.A(G326), .ZN(new_n779));
  NAND3_X1  g0579(.A1(new_n775), .A2(new_n439), .A3(G200), .ZN(new_n780));
  XOR2_X1   g0580(.A(KEYINPUT33), .B(G317), .Z(new_n781));
  OAI22_X1  g0581(.A1(new_n778), .A2(new_n779), .B1(new_n780), .B2(new_n781), .ZN(new_n782));
  NOR2_X1   g0582(.A1(new_n776), .A2(G200), .ZN(new_n783));
  AOI21_X1  g0583(.A(new_n782), .B1(G322), .B2(new_n783), .ZN(new_n784));
  INV_X1    g0584(.A(G311), .ZN(new_n785));
  NAND3_X1  g0585(.A1(new_n775), .A2(new_n439), .A3(new_n306), .ZN(new_n786));
  INV_X1    g0586(.A(KEYINPUT95), .ZN(new_n787));
  NAND2_X1  g0587(.A1(new_n786), .A2(new_n787), .ZN(new_n788));
  INV_X1    g0588(.A(new_n788), .ZN(new_n789));
  NOR2_X1   g0589(.A1(new_n786), .A2(new_n787), .ZN(new_n790));
  NOR2_X1   g0590(.A1(new_n789), .A2(new_n790), .ZN(new_n791));
  OAI211_X1 g0591(.A(new_n774), .B(new_n784), .C1(new_n785), .C2(new_n791), .ZN(new_n792));
  OAI22_X1  g0592(.A1(new_n778), .A2(new_n202), .B1(new_n208), .B2(new_n780), .ZN(new_n793));
  INV_X1    g0593(.A(KEYINPUT32), .ZN(new_n794));
  INV_X1    g0594(.A(G159), .ZN(new_n795));
  NOR2_X1   g0595(.A1(new_n772), .A2(new_n795), .ZN(new_n796));
  AOI21_X1  g0596(.A(new_n793), .B1(new_n794), .B2(new_n796), .ZN(new_n797));
  INV_X1    g0597(.A(new_n768), .ZN(new_n798));
  NAND2_X1  g0598(.A1(new_n798), .A2(G97), .ZN(new_n799));
  NOR2_X1   g0599(.A1(new_n764), .A2(new_n216), .ZN(new_n800));
  OAI21_X1  g0600(.A(new_n274), .B1(new_n770), .B2(new_n521), .ZN(new_n801));
  NOR2_X1   g0601(.A1(new_n800), .A2(new_n801), .ZN(new_n802));
  INV_X1    g0602(.A(new_n796), .ZN(new_n803));
  AOI22_X1  g0603(.A1(new_n783), .A2(G58), .B1(new_n803), .B2(KEYINPUT32), .ZN(new_n804));
  NAND4_X1  g0604(.A1(new_n797), .A2(new_n799), .A3(new_n802), .A4(new_n804), .ZN(new_n805));
  NOR2_X1   g0605(.A1(new_n791), .A2(new_n214), .ZN(new_n806));
  OAI21_X1  g0606(.A(new_n792), .B1(new_n805), .B2(new_n806), .ZN(new_n807));
  AOI21_X1  g0607(.A(new_n760), .B1(new_n807), .B2(new_n751), .ZN(new_n808));
  AOI21_X1  g0608(.A(new_n745), .B1(new_n750), .B2(new_n808), .ZN(new_n809));
  INV_X1    g0609(.A(new_n809), .ZN(new_n810));
  INV_X1    g0610(.A(KEYINPUT96), .ZN(new_n811));
  INV_X1    g0611(.A(new_n679), .ZN(new_n812));
  NOR2_X1   g0612(.A1(new_n678), .A2(G330), .ZN(new_n813));
  OAI21_X1  g0613(.A(new_n745), .B1(new_n812), .B2(new_n813), .ZN(new_n814));
  AND3_X1   g0614(.A1(new_n810), .A2(new_n811), .A3(new_n814), .ZN(new_n815));
  AOI21_X1  g0615(.A(new_n811), .B1(new_n810), .B2(new_n814), .ZN(new_n816));
  OR2_X1    g0616(.A1(new_n815), .A2(new_n816), .ZN(new_n817));
  INV_X1    g0617(.A(new_n817), .ZN(G396));
  NOR2_X1   g0618(.A1(new_n443), .A2(new_n675), .ZN(new_n819));
  NAND2_X1  g0619(.A1(new_n675), .A2(new_n425), .ZN(new_n820));
  NAND2_X1  g0620(.A1(new_n441), .A2(new_n820), .ZN(new_n821));
  AOI21_X1  g0621(.A(new_n819), .B1(new_n821), .B2(new_n443), .ZN(new_n822));
  INV_X1    g0622(.A(KEYINPUT99), .ZN(new_n823));
  XNOR2_X1  g0623(.A(new_n822), .B(new_n823), .ZN(new_n824));
  OR2_X1    g0624(.A1(new_n718), .A2(new_n824), .ZN(new_n825));
  OAI211_X1 g0625(.A(new_n665), .B(new_n649), .C1(KEYINPUT26), .C2(new_n704), .ZN(new_n826));
  AND3_X1   g0626(.A1(new_n647), .A2(new_n652), .A3(new_n653), .ZN(new_n827));
  OAI211_X1 g0627(.A(new_n676), .B(new_n822), .C1(new_n826), .C2(new_n827), .ZN(new_n828));
  INV_X1    g0628(.A(KEYINPUT100), .ZN(new_n829));
  NAND2_X1  g0629(.A1(new_n828), .A2(new_n829), .ZN(new_n830));
  NAND4_X1  g0630(.A1(new_n666), .A2(KEYINPUT100), .A3(new_n676), .A4(new_n822), .ZN(new_n831));
  NAND2_X1  g0631(.A1(new_n830), .A2(new_n831), .ZN(new_n832));
  AND2_X1   g0632(.A1(new_n825), .A2(new_n832), .ZN(new_n833));
  INV_X1    g0633(.A(new_n735), .ZN(new_n834));
  AND2_X1   g0634(.A1(new_n833), .A2(new_n834), .ZN(new_n835));
  OAI21_X1  g0635(.A(new_n745), .B1(new_n833), .B2(new_n834), .ZN(new_n836));
  NOR2_X1   g0636(.A1(new_n822), .A2(new_n747), .ZN(new_n837));
  INV_X1    g0637(.A(new_n751), .ZN(new_n838));
  AOI21_X1  g0638(.A(new_n274), .B1(G107), .B2(new_n769), .ZN(new_n839));
  NAND2_X1  g0639(.A1(new_n773), .A2(G311), .ZN(new_n840));
  NAND2_X1  g0640(.A1(new_n763), .A2(G87), .ZN(new_n841));
  NAND4_X1  g0641(.A1(new_n839), .A2(new_n799), .A3(new_n840), .A4(new_n841), .ZN(new_n842));
  INV_X1    g0642(.A(new_n780), .ZN(new_n843));
  AOI22_X1  g0643(.A1(G294), .A2(new_n783), .B1(new_n843), .B2(G283), .ZN(new_n844));
  OAI21_X1  g0644(.A(new_n844), .B1(new_n447), .B2(new_n778), .ZN(new_n845));
  INV_X1    g0645(.A(new_n791), .ZN(new_n846));
  AOI211_X1 g0646(.A(new_n842), .B(new_n845), .C1(G116), .C2(new_n846), .ZN(new_n847));
  XNOR2_X1  g0647(.A(new_n847), .B(KEYINPUT97), .ZN(new_n848));
  AOI22_X1  g0648(.A1(G137), .A2(new_n777), .B1(new_n783), .B2(G143), .ZN(new_n849));
  INV_X1    g0649(.A(G150), .ZN(new_n850));
  OAI221_X1 g0650(.A(new_n849), .B1(new_n850), .B2(new_n780), .C1(new_n791), .C2(new_n795), .ZN(new_n851));
  INV_X1    g0651(.A(KEYINPUT34), .ZN(new_n852));
  NOR2_X1   g0652(.A1(new_n851), .A2(new_n852), .ZN(new_n853));
  OAI21_X1  g0653(.A(new_n755), .B1(new_n770), .B2(new_n202), .ZN(new_n854));
  OAI22_X1  g0654(.A1(new_n764), .A2(new_n208), .B1(new_n323), .B2(new_n768), .ZN(new_n855));
  AOI211_X1 g0655(.A(new_n854), .B(new_n855), .C1(G132), .C2(new_n773), .ZN(new_n856));
  INV_X1    g0656(.A(new_n851), .ZN(new_n857));
  OAI21_X1  g0657(.A(new_n856), .B1(new_n857), .B2(KEYINPUT34), .ZN(new_n858));
  OAI21_X1  g0658(.A(new_n848), .B1(new_n853), .B2(new_n858), .ZN(new_n859));
  INV_X1    g0659(.A(KEYINPUT98), .ZN(new_n860));
  AOI21_X1  g0660(.A(new_n838), .B1(new_n859), .B2(new_n860), .ZN(new_n861));
  OAI21_X1  g0661(.A(new_n861), .B1(new_n860), .B2(new_n859), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n838), .A2(new_n747), .ZN(new_n863));
  OAI211_X1 g0663(.A(new_n862), .B(new_n744), .C1(G77), .C2(new_n863), .ZN(new_n864));
  OAI22_X1  g0664(.A1(new_n835), .A2(new_n836), .B1(new_n837), .B2(new_n864), .ZN(G384));
  NOR2_X1   g0665(.A1(new_n233), .A2(new_n479), .ZN(new_n866));
  OAI21_X1  g0666(.A(new_n866), .B1(new_n568), .B2(KEYINPUT35), .ZN(new_n867));
  INV_X1    g0667(.A(KEYINPUT101), .ZN(new_n868));
  AOI22_X1  g0668(.A1(new_n867), .A2(new_n868), .B1(KEYINPUT35), .B2(new_n568), .ZN(new_n869));
  OAI21_X1  g0669(.A(new_n869), .B1(new_n868), .B2(new_n867), .ZN(new_n870));
  XOR2_X1   g0670(.A(new_n870), .B(KEYINPUT36), .Z(new_n871));
  OR3_X1    g0671(.A1(new_n235), .A2(new_n214), .A3(new_n324), .ZN(new_n872));
  AOI211_X1 g0672(.A(new_n259), .B(G13), .C1(new_n872), .C2(new_n250), .ZN(new_n873));
  NOR2_X1   g0673(.A1(new_n871), .A2(new_n873), .ZN(new_n874));
  AOI21_X1  g0674(.A(new_n819), .B1(new_n830), .B2(new_n831), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n415), .A2(new_n675), .ZN(new_n876));
  OAI211_X1 g0676(.A(new_n406), .B(new_n876), .C1(new_n413), .C2(new_n405), .ZN(new_n877));
  OAI21_X1  g0677(.A(new_n877), .B1(new_n413), .B2(new_n876), .ZN(new_n878));
  INV_X1    g0678(.A(new_n878), .ZN(new_n879));
  NOR2_X1   g0679(.A1(new_n875), .A2(new_n879), .ZN(new_n880));
  INV_X1    g0680(.A(KEYINPUT38), .ZN(new_n881));
  AOI211_X1 g0681(.A(new_n328), .B(new_n330), .C1(new_n336), .C2(new_n339), .ZN(new_n882));
  OAI21_X1  g0682(.A(new_n292), .B1(new_n340), .B2(KEYINPUT16), .ZN(new_n883));
  AOI21_X1  g0683(.A(new_n882), .B1(new_n883), .B2(KEYINPUT102), .ZN(new_n884));
  INV_X1    g0684(.A(KEYINPUT102), .ZN(new_n885));
  OAI211_X1 g0685(.A(new_n885), .B(new_n292), .C1(new_n340), .C2(KEYINPUT16), .ZN(new_n886));
  AOI21_X1  g0686(.A(new_n316), .B1(new_n884), .B2(new_n886), .ZN(new_n887));
  OAI21_X1  g0687(.A(new_n372), .B1(new_n887), .B2(new_n673), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n883), .A2(KEYINPUT102), .ZN(new_n889));
  NAND3_X1  g0689(.A1(new_n889), .A2(new_n341), .A3(new_n886), .ZN(new_n890));
  AOI22_X1  g0690(.A1(new_n354), .A2(new_n356), .B1(new_n890), .B2(new_n368), .ZN(new_n891));
  OAI21_X1  g0691(.A(KEYINPUT37), .B1(new_n888), .B2(new_n891), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n892), .A2(KEYINPUT103), .ZN(new_n893));
  INV_X1    g0693(.A(KEYINPUT104), .ZN(new_n894));
  INV_X1    g0694(.A(KEYINPUT103), .ZN(new_n895));
  OAI211_X1 g0695(.A(new_n895), .B(KEYINPUT37), .C1(new_n888), .C2(new_n891), .ZN(new_n896));
  OAI21_X1  g0696(.A(new_n372), .B1(new_n342), .B2(new_n673), .ZN(new_n897));
  OR3_X1    g0697(.A1(new_n357), .A2(new_n897), .A3(KEYINPUT37), .ZN(new_n898));
  NAND4_X1  g0698(.A1(new_n893), .A2(new_n894), .A3(new_n896), .A4(new_n898), .ZN(new_n899));
  INV_X1    g0699(.A(new_n673), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n890), .A2(new_n368), .ZN(new_n901));
  NAND3_X1  g0701(.A1(new_n374), .A2(new_n900), .A3(new_n901), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n899), .A2(new_n902), .ZN(new_n903));
  NOR3_X1   g0703(.A1(new_n357), .A2(new_n897), .A3(KEYINPUT37), .ZN(new_n904));
  INV_X1    g0704(.A(KEYINPUT37), .ZN(new_n905));
  AND3_X1   g0705(.A1(new_n367), .A2(new_n368), .A3(new_n371), .ZN(new_n906));
  AOI21_X1  g0706(.A(new_n906), .B1(new_n901), .B2(new_n900), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n354), .A2(new_n356), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n908), .A2(new_n901), .ZN(new_n909));
  AOI21_X1  g0709(.A(new_n905), .B1(new_n907), .B2(new_n909), .ZN(new_n910));
  AOI21_X1  g0710(.A(new_n904), .B1(new_n910), .B2(new_n895), .ZN(new_n911));
  AOI21_X1  g0711(.A(new_n894), .B1(new_n911), .B2(new_n893), .ZN(new_n912));
  OAI21_X1  g0712(.A(new_n881), .B1(new_n903), .B2(new_n912), .ZN(new_n913));
  NOR2_X1   g0713(.A1(new_n910), .A2(new_n895), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n898), .A2(new_n896), .ZN(new_n915));
  OAI21_X1  g0715(.A(KEYINPUT104), .B1(new_n914), .B2(new_n915), .ZN(new_n916));
  NAND4_X1  g0716(.A1(new_n916), .A2(KEYINPUT38), .A3(new_n899), .A4(new_n902), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n913), .A2(new_n917), .ZN(new_n918));
  AOI22_X1  g0718(.A1(new_n880), .A2(new_n918), .B1(new_n641), .B2(new_n673), .ZN(new_n919));
  OR2_X1    g0719(.A1(new_n342), .A2(new_n673), .ZN(new_n920));
  NOR2_X1   g0720(.A1(new_n357), .A2(new_n897), .ZN(new_n921));
  NOR2_X1   g0721(.A1(new_n921), .A2(new_n905), .ZN(new_n922));
  OAI22_X1  g0722(.A1(new_n375), .A2(new_n920), .B1(new_n922), .B2(new_n904), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n923), .A2(new_n881), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n917), .A2(new_n924), .ZN(new_n925));
  INV_X1    g0725(.A(KEYINPUT39), .ZN(new_n926));
  NAND2_X1  g0726(.A1(new_n925), .A2(new_n926), .ZN(new_n927));
  NAND3_X1  g0727(.A1(new_n414), .A2(new_n415), .A3(new_n676), .ZN(new_n928));
  INV_X1    g0728(.A(new_n928), .ZN(new_n929));
  NAND3_X1  g0729(.A1(new_n913), .A2(KEYINPUT39), .A3(new_n917), .ZN(new_n930));
  NAND3_X1  g0730(.A1(new_n927), .A2(new_n929), .A3(new_n930), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n919), .A2(new_n931), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n717), .A2(new_n720), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n933), .A2(new_n446), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n934), .A2(new_n644), .ZN(new_n935));
  XNOR2_X1  g0735(.A(new_n932), .B(new_n935), .ZN(new_n936));
  INV_X1    g0736(.A(KEYINPUT105), .ZN(new_n937));
  NOR2_X1   g0737(.A1(new_n937), .A2(KEYINPUT31), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n730), .A2(new_n938), .ZN(new_n939));
  OAI211_X1 g0739(.A(new_n729), .B(new_n675), .C1(new_n937), .C2(KEYINPUT31), .ZN(new_n940));
  NAND3_X1  g0740(.A1(new_n721), .A2(new_n939), .A3(new_n940), .ZN(new_n941));
  AND3_X1   g0741(.A1(new_n878), .A2(new_n941), .A3(new_n822), .ZN(new_n942));
  NAND3_X1  g0742(.A1(new_n925), .A2(new_n942), .A3(KEYINPUT40), .ZN(new_n943));
  NAND3_X1  g0743(.A1(new_n878), .A2(new_n941), .A3(new_n822), .ZN(new_n944));
  AOI21_X1  g0744(.A(new_n944), .B1(new_n913), .B2(new_n917), .ZN(new_n945));
  OAI21_X1  g0745(.A(new_n943), .B1(new_n945), .B2(KEYINPUT40), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n446), .A2(new_n941), .ZN(new_n947));
  OR2_X1    g0747(.A1(new_n946), .A2(new_n947), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n946), .A2(new_n947), .ZN(new_n949));
  NAND3_X1  g0749(.A1(new_n948), .A2(G330), .A3(new_n949), .ZN(new_n950));
  AND2_X1   g0750(.A1(new_n936), .A2(new_n950), .ZN(new_n951));
  INV_X1    g0751(.A(KEYINPUT106), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n951), .A2(new_n952), .ZN(new_n953));
  OAI221_X1 g0753(.A(new_n953), .B1(new_n259), .B2(new_n741), .C1(new_n936), .C2(new_n950), .ZN(new_n954));
  NOR2_X1   g0754(.A1(new_n951), .A2(new_n952), .ZN(new_n955));
  OAI21_X1  g0755(.A(new_n874), .B1(new_n954), .B2(new_n955), .ZN(G367));
  OAI21_X1  g0756(.A(new_n752), .B1(new_n513), .B2(new_n221), .ZN(new_n957));
  AOI21_X1  g0757(.A(new_n957), .B1(new_n242), .B2(new_n756), .ZN(new_n958));
  NAND2_X1  g0758(.A1(new_n763), .A2(G97), .ZN(new_n959));
  OAI21_X1  g0759(.A(new_n959), .B1(new_n216), .B2(new_n768), .ZN(new_n960));
  AOI21_X1  g0760(.A(KEYINPUT46), .B1(new_n769), .B2(G116), .ZN(new_n961));
  NAND3_X1  g0761(.A1(new_n769), .A2(KEYINPUT46), .A3(G116), .ZN(new_n962));
  NAND2_X1  g0762(.A1(new_n962), .A2(new_n334), .ZN(new_n963));
  AOI211_X1 g0763(.A(new_n961), .B(new_n963), .C1(G303), .C2(new_n783), .ZN(new_n964));
  OAI221_X1 g0764(.A(new_n964), .B1(new_n585), .B2(new_n780), .C1(new_n785), .C2(new_n778), .ZN(new_n965));
  AOI211_X1 g0765(.A(new_n960), .B(new_n965), .C1(G317), .C2(new_n773), .ZN(new_n966));
  OAI21_X1  g0766(.A(new_n966), .B1(new_n765), .B2(new_n791), .ZN(new_n967));
  AOI22_X1  g0767(.A1(G143), .A2(new_n777), .B1(new_n783), .B2(G150), .ZN(new_n968));
  OAI21_X1  g0768(.A(new_n968), .B1(new_n795), .B2(new_n780), .ZN(new_n969));
  NAND2_X1  g0769(.A1(new_n763), .A2(G77), .ZN(new_n970));
  OAI211_X1 g0770(.A(new_n970), .B(new_n274), .C1(new_n323), .C2(new_n770), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n798), .A2(G68), .ZN(new_n972));
  INV_X1    g0772(.A(G137), .ZN(new_n973));
  OAI21_X1  g0773(.A(new_n972), .B1(new_n973), .B2(new_n772), .ZN(new_n974));
  NOR3_X1   g0774(.A1(new_n969), .A2(new_n971), .A3(new_n974), .ZN(new_n975));
  OAI21_X1  g0775(.A(new_n975), .B1(new_n202), .B2(new_n791), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n967), .A2(new_n976), .ZN(new_n977));
  XNOR2_X1  g0777(.A(new_n977), .B(KEYINPUT47), .ZN(new_n978));
  AOI211_X1 g0778(.A(new_n745), .B(new_n958), .C1(new_n978), .C2(new_n751), .ZN(new_n979));
  OR2_X1    g0779(.A1(new_n676), .A2(new_n548), .ZN(new_n980));
  OR2_X1    g0780(.A1(new_n980), .A2(new_n649), .ZN(new_n981));
  NAND2_X1  g0781(.A1(new_n980), .A2(new_n655), .ZN(new_n982));
  NAND3_X1  g0782(.A1(new_n981), .A2(new_n982), .A3(KEYINPUT107), .ZN(new_n983));
  OAI21_X1  g0783(.A(new_n983), .B1(KEYINPUT107), .B2(new_n981), .ZN(new_n984));
  INV_X1    g0784(.A(new_n984), .ZN(new_n985));
  OAI21_X1  g0785(.A(new_n979), .B1(new_n985), .B2(new_n749), .ZN(new_n986));
  NOR2_X1   g0786(.A1(new_n985), .A2(KEYINPUT43), .ZN(new_n987));
  INV_X1    g0787(.A(new_n987), .ZN(new_n988));
  OAI211_X1 g0788(.A(new_n709), .B(new_n711), .C1(new_n572), .C2(new_n676), .ZN(new_n989));
  NAND2_X1  g0789(.A1(new_n573), .A2(new_n675), .ZN(new_n990));
  NAND2_X1  g0790(.A1(new_n989), .A2(new_n990), .ZN(new_n991));
  INV_X1    g0791(.A(new_n991), .ZN(new_n992));
  NOR2_X1   g0792(.A1(new_n992), .A2(new_n689), .ZN(new_n993));
  XNOR2_X1  g0793(.A(new_n993), .B(KEYINPUT42), .ZN(new_n994));
  XNOR2_X1  g0794(.A(new_n991), .B(KEYINPUT108), .ZN(new_n995));
  INV_X1    g0795(.A(new_n995), .ZN(new_n996));
  AOI21_X1  g0796(.A(new_n573), .B1(new_n996), .B2(new_n628), .ZN(new_n997));
  OAI21_X1  g0797(.A(new_n994), .B1(new_n997), .B2(new_n675), .ZN(new_n998));
  INV_X1    g0798(.A(KEYINPUT43), .ZN(new_n999));
  OAI21_X1  g0799(.A(new_n998), .B1(new_n999), .B2(new_n984), .ZN(new_n1000));
  NOR2_X1   g0800(.A1(new_n687), .A2(new_n995), .ZN(new_n1001));
  XNOR2_X1  g0801(.A(new_n1001), .B(KEYINPUT109), .ZN(new_n1002));
  NAND2_X1  g0802(.A1(new_n1000), .A2(new_n1002), .ZN(new_n1003));
  INV_X1    g0803(.A(new_n1003), .ZN(new_n1004));
  NOR2_X1   g0804(.A1(new_n1000), .A2(new_n1002), .ZN(new_n1005));
  OAI21_X1  g0805(.A(new_n988), .B1(new_n1004), .B2(new_n1005), .ZN(new_n1006));
  INV_X1    g0806(.A(new_n1005), .ZN(new_n1007));
  NAND3_X1  g0807(.A1(new_n1007), .A2(new_n987), .A3(new_n1003), .ZN(new_n1008));
  NAND2_X1  g0808(.A1(new_n1006), .A2(new_n1008), .ZN(new_n1009));
  INV_X1    g0809(.A(new_n694), .ZN(new_n1010));
  AOI21_X1  g0810(.A(new_n992), .B1(new_n1010), .B2(new_n692), .ZN(new_n1011));
  XNOR2_X1  g0811(.A(new_n1011), .B(KEYINPUT45), .ZN(new_n1012));
  NOR3_X1   g0812(.A1(new_n693), .A2(new_n694), .A3(new_n991), .ZN(new_n1013));
  XNOR2_X1  g0813(.A(new_n1013), .B(KEYINPUT44), .ZN(new_n1014));
  NAND2_X1  g0814(.A1(new_n1012), .A2(new_n1014), .ZN(new_n1015));
  NAND2_X1  g0815(.A1(new_n1015), .A2(new_n686), .ZN(new_n1016));
  NAND3_X1  g0816(.A1(new_n1012), .A2(new_n1014), .A3(new_n687), .ZN(new_n1017));
  XOR2_X1   g0817(.A(new_n685), .B(new_n688), .Z(new_n1018));
  XNOR2_X1  g0818(.A(new_n1018), .B(new_n679), .ZN(new_n1019));
  INV_X1    g0819(.A(new_n1019), .ZN(new_n1020));
  NAND4_X1  g0820(.A1(new_n1016), .A2(new_n739), .A3(new_n1017), .A4(new_n1020), .ZN(new_n1021));
  NAND2_X1  g0821(.A1(new_n1021), .A2(new_n739), .ZN(new_n1022));
  XOR2_X1   g0822(.A(KEYINPUT110), .B(KEYINPUT41), .Z(new_n1023));
  XNOR2_X1  g0823(.A(new_n696), .B(new_n1023), .ZN(new_n1024));
  AOI21_X1  g0824(.A(new_n743), .B1(new_n1022), .B2(new_n1024), .ZN(new_n1025));
  OAI21_X1  g0825(.A(new_n986), .B1(new_n1009), .B2(new_n1025), .ZN(new_n1026));
  INV_X1    g0826(.A(KEYINPUT111), .ZN(new_n1027));
  NAND2_X1  g0827(.A1(new_n1026), .A2(new_n1027), .ZN(new_n1028));
  OAI211_X1 g0828(.A(KEYINPUT111), .B(new_n986), .C1(new_n1009), .C2(new_n1025), .ZN(new_n1029));
  AND2_X1   g0829(.A1(new_n1028), .A2(new_n1029), .ZN(G387));
  NAND2_X1  g0830(.A1(new_n739), .A2(new_n1020), .ZN(new_n1031));
  NAND3_X1  g0831(.A1(new_n737), .A2(new_n738), .A3(new_n1019), .ZN(new_n1032));
  NAND3_X1  g0832(.A1(new_n1031), .A2(new_n696), .A3(new_n1032), .ZN(new_n1033));
  NAND2_X1  g0833(.A1(new_n758), .A2(new_n699), .ZN(new_n1034));
  OAI21_X1  g0834(.A(new_n1034), .B1(G107), .B2(new_n221), .ZN(new_n1035));
  AOI211_X1 g0835(.A(new_n222), .B(new_n755), .C1(new_n248), .C2(G45), .ZN(new_n1036));
  XOR2_X1   g0836(.A(new_n699), .B(KEYINPUT112), .Z(new_n1037));
  OAI21_X1  g0837(.A(new_n460), .B1(new_n208), .B2(new_n214), .ZN(new_n1038));
  NAND2_X1  g0838(.A1(new_n314), .A2(new_n202), .ZN(new_n1039));
  AOI21_X1  g0839(.A(new_n1038), .B1(new_n1039), .B2(KEYINPUT50), .ZN(new_n1040));
  OAI211_X1 g0840(.A(new_n1037), .B(new_n1040), .C1(KEYINPUT50), .C2(new_n1039), .ZN(new_n1041));
  AOI21_X1  g0841(.A(new_n1035), .B1(new_n1036), .B2(new_n1041), .ZN(new_n1042));
  NAND2_X1  g0842(.A1(new_n777), .A2(G159), .ZN(new_n1043));
  XNOR2_X1  g0843(.A(new_n1043), .B(KEYINPUT113), .ZN(new_n1044));
  NOR2_X1   g0844(.A1(new_n791), .A2(new_n208), .ZN(new_n1045));
  NAND2_X1  g0845(.A1(new_n418), .A2(new_n798), .ZN(new_n1046));
  AOI21_X1  g0846(.A(new_n334), .B1(new_n769), .B2(G77), .ZN(new_n1047));
  NAND2_X1  g0847(.A1(new_n773), .A2(G150), .ZN(new_n1048));
  NAND4_X1  g0848(.A1(new_n1046), .A2(new_n959), .A3(new_n1047), .A4(new_n1048), .ZN(new_n1049));
  INV_X1    g0849(.A(new_n783), .ZN(new_n1050));
  OAI22_X1  g0850(.A1(new_n1050), .A2(new_n202), .B1(new_n288), .B2(new_n780), .ZN(new_n1051));
  NOR4_X1   g0851(.A1(new_n1044), .A2(new_n1045), .A3(new_n1049), .A4(new_n1051), .ZN(new_n1052));
  AOI22_X1  g0852(.A1(G317), .A2(new_n783), .B1(new_n777), .B2(G322), .ZN(new_n1053));
  OAI21_X1  g0853(.A(new_n1053), .B1(new_n785), .B2(new_n780), .ZN(new_n1054));
  AOI21_X1  g0854(.A(new_n1054), .B1(G303), .B2(new_n846), .ZN(new_n1055));
  OR2_X1    g0855(.A1(new_n1055), .A2(KEYINPUT48), .ZN(new_n1056));
  NAND2_X1  g0856(.A1(new_n1055), .A2(KEYINPUT48), .ZN(new_n1057));
  AOI22_X1  g0857(.A1(new_n798), .A2(G283), .B1(G294), .B2(new_n769), .ZN(new_n1058));
  XNOR2_X1  g0858(.A(new_n1058), .B(KEYINPUT114), .ZN(new_n1059));
  NAND3_X1  g0859(.A1(new_n1056), .A2(new_n1057), .A3(new_n1059), .ZN(new_n1060));
  INV_X1    g0860(.A(KEYINPUT49), .ZN(new_n1061));
  NOR2_X1   g0861(.A1(new_n1060), .A2(new_n1061), .ZN(new_n1062));
  OAI221_X1 g0862(.A(new_n334), .B1(new_n779), .B2(new_n772), .C1(new_n764), .C2(new_n479), .ZN(new_n1063));
  XOR2_X1   g0863(.A(new_n1063), .B(KEYINPUT115), .Z(new_n1064));
  NOR2_X1   g0864(.A1(new_n1062), .A2(new_n1064), .ZN(new_n1065));
  NAND2_X1  g0865(.A1(new_n1060), .A2(new_n1061), .ZN(new_n1066));
  AOI21_X1  g0866(.A(new_n1052), .B1(new_n1065), .B2(new_n1066), .ZN(new_n1067));
  OAI221_X1 g0867(.A(new_n744), .B1(new_n753), .B2(new_n1042), .C1(new_n1067), .C2(new_n838), .ZN(new_n1068));
  AOI21_X1  g0868(.A(new_n1068), .B1(new_n685), .B2(new_n748), .ZN(new_n1069));
  AOI21_X1  g0869(.A(new_n1069), .B1(new_n1020), .B2(new_n743), .ZN(new_n1070));
  NAND2_X1  g0870(.A1(new_n1033), .A2(new_n1070), .ZN(G393));
  NAND2_X1  g0871(.A1(new_n1016), .A2(new_n1017), .ZN(new_n1072));
  AND2_X1   g0872(.A1(new_n1072), .A2(new_n1031), .ZN(new_n1073));
  NAND2_X1  g0873(.A1(new_n1021), .A2(new_n696), .ZN(new_n1074));
  NOR2_X1   g0874(.A1(new_n1073), .A2(new_n1074), .ZN(new_n1075));
  NOR2_X1   g0875(.A1(new_n768), .A2(new_n214), .ZN(new_n1076));
  AOI21_X1  g0876(.A(new_n1076), .B1(new_n843), .B2(G50), .ZN(new_n1077));
  OAI21_X1  g0877(.A(new_n1077), .B1(new_n791), .B2(new_n288), .ZN(new_n1078));
  XNOR2_X1  g0878(.A(new_n1078), .B(KEYINPUT116), .ZN(new_n1079));
  AOI22_X1  g0879(.A1(G150), .A2(new_n777), .B1(new_n783), .B2(G159), .ZN(new_n1080));
  XNOR2_X1  g0880(.A(new_n1080), .B(KEYINPUT51), .ZN(new_n1081));
  AOI21_X1  g0881(.A(new_n334), .B1(new_n769), .B2(G68), .ZN(new_n1082));
  NAND2_X1  g0882(.A1(new_n773), .A2(G143), .ZN(new_n1083));
  NAND3_X1  g0883(.A1(new_n1082), .A2(new_n1083), .A3(new_n841), .ZN(new_n1084));
  NOR3_X1   g0884(.A1(new_n1079), .A2(new_n1081), .A3(new_n1084), .ZN(new_n1085));
  INV_X1    g0885(.A(new_n800), .ZN(new_n1086));
  NAND2_X1  g0886(.A1(new_n843), .A2(G303), .ZN(new_n1087));
  AOI21_X1  g0887(.A(new_n274), .B1(G283), .B2(new_n769), .ZN(new_n1088));
  AOI22_X1  g0888(.A1(new_n798), .A2(G116), .B1(new_n773), .B2(G322), .ZN(new_n1089));
  NAND4_X1  g0889(.A1(new_n1086), .A2(new_n1087), .A3(new_n1088), .A4(new_n1089), .ZN(new_n1090));
  AOI22_X1  g0890(.A1(G311), .A2(new_n783), .B1(new_n777), .B2(G317), .ZN(new_n1091));
  XNOR2_X1  g0891(.A(new_n1091), .B(KEYINPUT52), .ZN(new_n1092));
  AOI211_X1 g0892(.A(new_n1090), .B(new_n1092), .C1(G294), .C2(new_n846), .ZN(new_n1093));
  OAI21_X1  g0893(.A(new_n751), .B1(new_n1085), .B2(new_n1093), .ZN(new_n1094));
  AND2_X1   g0894(.A1(new_n257), .A2(new_n756), .ZN(new_n1095));
  OAI21_X1  g0895(.A(new_n752), .B1(new_n483), .B2(new_n221), .ZN(new_n1096));
  OAI211_X1 g0896(.A(new_n1094), .B(new_n744), .C1(new_n1095), .C2(new_n1096), .ZN(new_n1097));
  XOR2_X1   g0897(.A(new_n1097), .B(KEYINPUT117), .Z(new_n1098));
  OAI21_X1  g0898(.A(new_n1098), .B1(new_n996), .B2(new_n749), .ZN(new_n1099));
  INV_X1    g0899(.A(new_n743), .ZN(new_n1100));
  OAI21_X1  g0900(.A(new_n1099), .B1(new_n1072), .B2(new_n1100), .ZN(new_n1101));
  NOR2_X1   g0901(.A1(new_n1075), .A2(new_n1101), .ZN(new_n1102));
  INV_X1    g0902(.A(new_n1102), .ZN(G390));
  OAI21_X1  g0903(.A(new_n928), .B1(new_n875), .B2(new_n879), .ZN(new_n1104));
  AND3_X1   g0904(.A1(new_n913), .A2(KEYINPUT39), .A3(new_n917), .ZN(new_n1105));
  AOI21_X1  g0905(.A(KEYINPUT39), .B1(new_n917), .B2(new_n924), .ZN(new_n1106));
  OAI21_X1  g0906(.A(new_n1104), .B1(new_n1105), .B2(new_n1106), .ZN(new_n1107));
  NAND2_X1  g0907(.A1(new_n712), .A2(new_n715), .ZN(new_n1108));
  INV_X1    g0908(.A(new_n706), .ZN(new_n1109));
  AOI21_X1  g0909(.A(new_n675), .B1(new_n1108), .B2(new_n1109), .ZN(new_n1110));
  NAND2_X1  g0910(.A1(new_n821), .A2(new_n443), .ZN(new_n1111));
  AOI21_X1  g0911(.A(new_n819), .B1(new_n1110), .B2(new_n1111), .ZN(new_n1112));
  OAI211_X1 g0912(.A(new_n928), .B(new_n925), .C1(new_n1112), .C2(new_n879), .ZN(new_n1113));
  NAND4_X1  g0913(.A1(new_n878), .A2(new_n734), .A3(G330), .A4(new_n822), .ZN(new_n1114));
  NAND3_X1  g0914(.A1(new_n1107), .A2(new_n1113), .A3(new_n1114), .ZN(new_n1115));
  NAND2_X1  g0915(.A1(new_n1115), .A2(KEYINPUT118), .ZN(new_n1116));
  INV_X1    g0916(.A(KEYINPUT118), .ZN(new_n1117));
  NAND4_X1  g0917(.A1(new_n1107), .A2(new_n1113), .A3(new_n1117), .A4(new_n1114), .ZN(new_n1118));
  NAND4_X1  g0918(.A1(new_n878), .A2(new_n941), .A3(G330), .A4(new_n822), .ZN(new_n1119));
  INV_X1    g0919(.A(new_n1119), .ZN(new_n1120));
  INV_X1    g0920(.A(new_n819), .ZN(new_n1121));
  NAND2_X1  g0921(.A1(new_n832), .A2(new_n1121), .ZN(new_n1122));
  NAND2_X1  g0922(.A1(new_n1122), .A2(new_n878), .ZN(new_n1123));
  AOI22_X1  g0923(.A1(new_n1123), .A2(new_n928), .B1(new_n927), .B2(new_n930), .ZN(new_n1124));
  NAND2_X1  g0924(.A1(new_n925), .A2(new_n928), .ZN(new_n1125));
  NAND2_X1  g0925(.A1(new_n1110), .A2(new_n1111), .ZN(new_n1126));
  NAND2_X1  g0926(.A1(new_n1126), .A2(new_n1121), .ZN(new_n1127));
  AOI21_X1  g0927(.A(new_n1125), .B1(new_n1127), .B2(new_n878), .ZN(new_n1128));
  OAI21_X1  g0928(.A(new_n1120), .B1(new_n1124), .B2(new_n1128), .ZN(new_n1129));
  NAND3_X1  g0929(.A1(new_n1116), .A2(new_n1118), .A3(new_n1129), .ZN(new_n1130));
  NAND3_X1  g0930(.A1(new_n941), .A2(G330), .A3(new_n824), .ZN(new_n1131));
  NAND2_X1  g0931(.A1(new_n1131), .A2(new_n879), .ZN(new_n1132));
  AND2_X1   g0932(.A1(new_n1132), .A2(new_n1114), .ZN(new_n1133));
  NAND3_X1  g0933(.A1(new_n734), .A2(G330), .A3(new_n822), .ZN(new_n1134));
  NAND2_X1  g0934(.A1(new_n1134), .A2(new_n879), .ZN(new_n1135));
  NAND2_X1  g0935(.A1(new_n1135), .A2(new_n1119), .ZN(new_n1136));
  AOI22_X1  g0936(.A1(new_n1133), .A2(new_n1112), .B1(new_n1136), .B2(new_n1122), .ZN(new_n1137));
  NAND2_X1  g0937(.A1(new_n941), .A2(G330), .ZN(new_n1138));
  NOR2_X1   g0938(.A1(new_n445), .A2(new_n1138), .ZN(new_n1139));
  INV_X1    g0939(.A(new_n1139), .ZN(new_n1140));
  NAND3_X1  g0940(.A1(new_n934), .A2(new_n1140), .A3(new_n644), .ZN(new_n1141));
  NOR2_X1   g0941(.A1(new_n1137), .A2(new_n1141), .ZN(new_n1142));
  INV_X1    g0942(.A(new_n1142), .ZN(new_n1143));
  NAND2_X1  g0943(.A1(new_n1130), .A2(new_n1143), .ZN(new_n1144));
  NAND4_X1  g0944(.A1(new_n1116), .A2(new_n1118), .A3(new_n1129), .A4(new_n1142), .ZN(new_n1145));
  NAND3_X1  g0945(.A1(new_n1144), .A2(new_n696), .A3(new_n1145), .ZN(new_n1146));
  AND3_X1   g0946(.A1(new_n1116), .A2(new_n1118), .A3(new_n1129), .ZN(new_n1147));
  OAI21_X1  g0947(.A(new_n746), .B1(new_n1105), .B2(new_n1106), .ZN(new_n1148));
  OAI21_X1  g0948(.A(new_n744), .B1(new_n314), .B2(new_n863), .ZN(new_n1149));
  OAI221_X1 g0949(.A(new_n364), .B1(new_n770), .B2(new_n210), .C1(new_n764), .C2(new_n208), .ZN(new_n1150));
  AOI211_X1 g0950(.A(new_n1076), .B(new_n1150), .C1(G294), .C2(new_n773), .ZN(new_n1151));
  OAI22_X1  g0951(.A1(new_n778), .A2(new_n765), .B1(new_n216), .B2(new_n780), .ZN(new_n1152));
  AOI21_X1  g0952(.A(new_n1152), .B1(G116), .B2(new_n783), .ZN(new_n1153));
  OAI211_X1 g0953(.A(new_n1151), .B(new_n1153), .C1(new_n483), .C2(new_n791), .ZN(new_n1154));
  XNOR2_X1  g0954(.A(KEYINPUT54), .B(G143), .ZN(new_n1155));
  NOR2_X1   g0955(.A1(new_n791), .A2(new_n1155), .ZN(new_n1156));
  NOR3_X1   g0956(.A1(new_n770), .A2(KEYINPUT53), .A3(new_n850), .ZN(new_n1157));
  OAI21_X1  g0957(.A(KEYINPUT53), .B1(new_n770), .B2(new_n850), .ZN(new_n1158));
  NAND2_X1  g0958(.A1(new_n1158), .A2(new_n274), .ZN(new_n1159));
  AOI211_X1 g0959(.A(new_n1157), .B(new_n1159), .C1(G137), .C2(new_n843), .ZN(new_n1160));
  AOI22_X1  g0960(.A1(G128), .A2(new_n777), .B1(new_n783), .B2(G132), .ZN(new_n1161));
  OAI22_X1  g0961(.A1(new_n764), .A2(new_n202), .B1(new_n795), .B2(new_n768), .ZN(new_n1162));
  AOI21_X1  g0962(.A(new_n1162), .B1(G125), .B2(new_n773), .ZN(new_n1163));
  NAND3_X1  g0963(.A1(new_n1160), .A2(new_n1161), .A3(new_n1163), .ZN(new_n1164));
  OAI21_X1  g0964(.A(new_n1154), .B1(new_n1156), .B2(new_n1164), .ZN(new_n1165));
  AOI21_X1  g0965(.A(new_n1149), .B1(new_n1165), .B2(new_n751), .ZN(new_n1166));
  AOI22_X1  g0966(.A1(new_n1147), .A2(new_n743), .B1(new_n1148), .B2(new_n1166), .ZN(new_n1167));
  NAND2_X1  g0967(.A1(new_n1146), .A2(new_n1167), .ZN(G378));
  AOI21_X1  g0968(.A(new_n445), .B1(new_n717), .B2(new_n720), .ZN(new_n1169));
  NOR3_X1   g0969(.A1(new_n1169), .A2(new_n643), .A3(new_n1139), .ZN(new_n1170));
  NAND2_X1  g0970(.A1(new_n1145), .A2(new_n1170), .ZN(new_n1171));
  OAI211_X1 g0971(.A(new_n943), .B(G330), .C1(new_n945), .C2(KEYINPUT40), .ZN(new_n1172));
  NAND2_X1  g0972(.A1(new_n900), .A2(new_n304), .ZN(new_n1173));
  XNOR2_X1  g0973(.A(new_n312), .B(new_n1173), .ZN(new_n1174));
  XNOR2_X1  g0974(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1175));
  INV_X1    g0975(.A(new_n1175), .ZN(new_n1176));
  XNOR2_X1  g0976(.A(new_n1174), .B(new_n1176), .ZN(new_n1177));
  AND2_X1   g0977(.A1(new_n1172), .A2(new_n1177), .ZN(new_n1178));
  NOR2_X1   g0978(.A1(new_n1172), .A2(new_n1177), .ZN(new_n1179));
  OAI21_X1  g0979(.A(new_n932), .B1(new_n1178), .B2(new_n1179), .ZN(new_n1180));
  OR2_X1    g0980(.A1(new_n1172), .A2(new_n1177), .ZN(new_n1181));
  INV_X1    g0981(.A(new_n932), .ZN(new_n1182));
  NAND2_X1  g0982(.A1(new_n1172), .A2(new_n1177), .ZN(new_n1183));
  NAND3_X1  g0983(.A1(new_n1181), .A2(new_n1182), .A3(new_n1183), .ZN(new_n1184));
  NAND2_X1  g0984(.A1(new_n1180), .A2(new_n1184), .ZN(new_n1185));
  NAND2_X1  g0985(.A1(new_n1171), .A2(new_n1185), .ZN(new_n1186));
  INV_X1    g0986(.A(KEYINPUT57), .ZN(new_n1187));
  NAND2_X1  g0987(.A1(new_n1186), .A2(new_n1187), .ZN(new_n1188));
  AOI21_X1  g0988(.A(new_n1187), .B1(new_n1180), .B2(new_n1184), .ZN(new_n1189));
  AOI21_X1  g0989(.A(new_n697), .B1(new_n1189), .B2(new_n1171), .ZN(new_n1190));
  NAND2_X1  g0990(.A1(new_n1188), .A2(new_n1190), .ZN(new_n1191));
  NAND2_X1  g0991(.A1(new_n1177), .A2(new_n746), .ZN(new_n1192));
  OAI21_X1  g0992(.A(new_n744), .B1(G50), .B2(new_n863), .ZN(new_n1193));
  NAND2_X1  g0993(.A1(new_n763), .A2(G58), .ZN(new_n1194));
  XNOR2_X1  g0994(.A(new_n1194), .B(KEYINPUT119), .ZN(new_n1195));
  AOI211_X1 g0995(.A(G41), .B(new_n755), .C1(G77), .C2(new_n769), .ZN(new_n1196));
  OAI211_X1 g0996(.A(new_n1195), .B(new_n1196), .C1(new_n765), .C2(new_n772), .ZN(new_n1197));
  XOR2_X1   g0997(.A(new_n1197), .B(KEYINPUT120), .Z(new_n1198));
  NAND2_X1  g0998(.A1(new_n783), .A2(G107), .ZN(new_n1199));
  XNOR2_X1  g0999(.A(new_n1199), .B(KEYINPUT121), .ZN(new_n1200));
  OAI221_X1 g1000(.A(new_n972), .B1(new_n483), .B2(new_n780), .C1(new_n778), .C2(new_n479), .ZN(new_n1201));
  AOI21_X1  g1001(.A(new_n1201), .B1(new_n418), .B2(new_n846), .ZN(new_n1202));
  NAND3_X1  g1002(.A1(new_n1198), .A2(new_n1200), .A3(new_n1202), .ZN(new_n1203));
  XNOR2_X1  g1003(.A(new_n1203), .B(KEYINPUT58), .ZN(new_n1204));
  NAND2_X1  g1004(.A1(new_n798), .A2(G150), .ZN(new_n1205));
  INV_X1    g1005(.A(G132), .ZN(new_n1206));
  OAI221_X1 g1006(.A(new_n1205), .B1(new_n1206), .B2(new_n780), .C1(new_n770), .C2(new_n1155), .ZN(new_n1207));
  NAND2_X1  g1007(.A1(new_n777), .A2(G125), .ZN(new_n1208));
  INV_X1    g1008(.A(G128), .ZN(new_n1209));
  OAI21_X1  g1009(.A(new_n1208), .B1(new_n1050), .B2(new_n1209), .ZN(new_n1210));
  AOI211_X1 g1010(.A(new_n1207), .B(new_n1210), .C1(new_n846), .C2(G137), .ZN(new_n1211));
  INV_X1    g1011(.A(KEYINPUT59), .ZN(new_n1212));
  OR2_X1    g1012(.A1(new_n1211), .A2(new_n1212), .ZN(new_n1213));
  NAND2_X1  g1013(.A1(new_n1211), .A2(new_n1212), .ZN(new_n1214));
  NAND2_X1  g1014(.A1(new_n763), .A2(G159), .ZN(new_n1215));
  AOI211_X1 g1015(.A(G33), .B(G41), .C1(new_n773), .C2(G124), .ZN(new_n1216));
  NAND4_X1  g1016(.A1(new_n1213), .A2(new_n1214), .A3(new_n1215), .A4(new_n1216), .ZN(new_n1217));
  AOI21_X1  g1017(.A(G50), .B1(new_n269), .B2(new_n428), .ZN(new_n1218));
  OAI21_X1  g1018(.A(new_n1218), .B1(new_n755), .B2(G41), .ZN(new_n1219));
  NAND3_X1  g1019(.A1(new_n1204), .A2(new_n1217), .A3(new_n1219), .ZN(new_n1220));
  AOI21_X1  g1020(.A(new_n1193), .B1(new_n1220), .B2(new_n751), .ZN(new_n1221));
  AOI22_X1  g1021(.A1(new_n1185), .A2(new_n743), .B1(new_n1192), .B2(new_n1221), .ZN(new_n1222));
  NAND2_X1  g1022(.A1(new_n1191), .A2(new_n1222), .ZN(G375));
  NAND2_X1  g1023(.A1(new_n1137), .A2(new_n1141), .ZN(new_n1224));
  NAND3_X1  g1024(.A1(new_n1143), .A2(new_n1024), .A3(new_n1224), .ZN(new_n1225));
  AOI21_X1  g1025(.A(new_n274), .B1(G97), .B2(new_n769), .ZN(new_n1226));
  NAND2_X1  g1026(.A1(new_n773), .A2(G303), .ZN(new_n1227));
  NAND4_X1  g1027(.A1(new_n1226), .A2(new_n1046), .A3(new_n970), .A4(new_n1227), .ZN(new_n1228));
  AOI22_X1  g1028(.A1(G283), .A2(new_n783), .B1(new_n777), .B2(G294), .ZN(new_n1229));
  OAI21_X1  g1029(.A(new_n1229), .B1(new_n479), .B2(new_n780), .ZN(new_n1230));
  AOI211_X1 g1030(.A(new_n1228), .B(new_n1230), .C1(G107), .C2(new_n846), .ZN(new_n1231));
  AOI21_X1  g1031(.A(new_n334), .B1(new_n769), .B2(G159), .ZN(new_n1232));
  OAI221_X1 g1032(.A(new_n1232), .B1(new_n1209), .B2(new_n772), .C1(new_n780), .C2(new_n1155), .ZN(new_n1233));
  OR3_X1    g1033(.A1(new_n778), .A2(KEYINPUT122), .A3(new_n1206), .ZN(new_n1234));
  OAI21_X1  g1034(.A(KEYINPUT122), .B1(new_n778), .B2(new_n1206), .ZN(new_n1235));
  NAND3_X1  g1035(.A1(new_n1234), .A2(new_n1195), .A3(new_n1235), .ZN(new_n1236));
  AOI211_X1 g1036(.A(new_n1233), .B(new_n1236), .C1(G137), .C2(new_n783), .ZN(new_n1237));
  OAI22_X1  g1037(.A1(new_n791), .A2(new_n850), .B1(new_n202), .B2(new_n768), .ZN(new_n1238));
  XOR2_X1   g1038(.A(new_n1238), .B(KEYINPUT123), .Z(new_n1239));
  AOI21_X1  g1039(.A(new_n1231), .B1(new_n1237), .B2(new_n1239), .ZN(new_n1240));
  OAI221_X1 g1040(.A(new_n744), .B1(G68), .B2(new_n863), .C1(new_n1240), .C2(new_n838), .ZN(new_n1241));
  AOI21_X1  g1041(.A(new_n1241), .B1(new_n879), .B2(new_n746), .ZN(new_n1242));
  AOI22_X1  g1042(.A1(new_n942), .A2(G330), .B1(new_n1134), .B2(new_n879), .ZN(new_n1243));
  NAND2_X1  g1043(.A1(new_n1132), .A2(new_n1114), .ZN(new_n1244));
  OAI22_X1  g1044(.A1(new_n875), .A2(new_n1243), .B1(new_n1127), .B2(new_n1244), .ZN(new_n1245));
  AOI21_X1  g1045(.A(new_n1242), .B1(new_n1245), .B2(new_n743), .ZN(new_n1246));
  NAND2_X1  g1046(.A1(new_n1225), .A2(new_n1246), .ZN(new_n1247));
  XOR2_X1   g1047(.A(new_n1247), .B(KEYINPUT124), .Z(new_n1248));
  INV_X1    g1048(.A(new_n1248), .ZN(G381));
  NOR2_X1   g1049(.A1(G393), .A2(G396), .ZN(new_n1250));
  INV_X1    g1050(.A(G384), .ZN(new_n1251));
  AOI21_X1  g1051(.A(KEYINPUT125), .B1(new_n1250), .B2(new_n1251), .ZN(new_n1252));
  NAND3_X1  g1052(.A1(new_n1250), .A2(KEYINPUT125), .A3(new_n1251), .ZN(new_n1253));
  NAND3_X1  g1053(.A1(new_n1248), .A2(new_n1102), .A3(new_n1253), .ZN(new_n1254));
  OR3_X1    g1054(.A1(G387), .A2(new_n1252), .A3(new_n1254), .ZN(new_n1255));
  NAND2_X1  g1055(.A1(new_n1185), .A2(new_n743), .ZN(new_n1256));
  NAND2_X1  g1056(.A1(new_n1192), .A2(new_n1221), .ZN(new_n1257));
  NAND2_X1  g1057(.A1(new_n1256), .A2(new_n1257), .ZN(new_n1258));
  AOI21_X1  g1058(.A(new_n1258), .B1(new_n1188), .B2(new_n1190), .ZN(new_n1259));
  INV_X1    g1059(.A(G378), .ZN(new_n1260));
  NAND2_X1  g1060(.A1(new_n1259), .A2(new_n1260), .ZN(new_n1261));
  OR2_X1    g1061(.A1(new_n1255), .A2(new_n1261), .ZN(G407));
  NAND2_X1  g1062(.A1(new_n674), .A2(G213), .ZN(new_n1263));
  OR2_X1    g1063(.A1(new_n1261), .A2(new_n1263), .ZN(new_n1264));
  OAI211_X1 g1064(.A(new_n1264), .B(G213), .C1(new_n1255), .C2(new_n1261), .ZN(G409));
  NAND3_X1  g1065(.A1(new_n1171), .A2(new_n1024), .A3(new_n1185), .ZN(new_n1266));
  NAND4_X1  g1066(.A1(new_n1222), .A2(new_n1266), .A3(new_n1146), .A4(new_n1167), .ZN(new_n1267));
  OAI211_X1 g1067(.A(new_n1263), .B(new_n1267), .C1(new_n1259), .C2(new_n1260), .ZN(new_n1268));
  INV_X1    g1068(.A(KEYINPUT126), .ZN(new_n1269));
  INV_X1    g1069(.A(KEYINPUT60), .ZN(new_n1270));
  AOI21_X1  g1070(.A(new_n1270), .B1(new_n1245), .B2(new_n1170), .ZN(new_n1271));
  NOR2_X1   g1071(.A1(new_n1245), .A2(new_n1170), .ZN(new_n1272));
  OAI21_X1  g1072(.A(new_n1269), .B1(new_n1271), .B2(new_n1272), .ZN(new_n1273));
  OAI21_X1  g1073(.A(KEYINPUT60), .B1(new_n1137), .B2(new_n1141), .ZN(new_n1274));
  NAND3_X1  g1074(.A1(new_n1274), .A2(KEYINPUT126), .A3(new_n1224), .ZN(new_n1275));
  AOI21_X1  g1075(.A(new_n697), .B1(new_n1272), .B2(KEYINPUT60), .ZN(new_n1276));
  NAND3_X1  g1076(.A1(new_n1273), .A2(new_n1275), .A3(new_n1276), .ZN(new_n1277));
  AND3_X1   g1077(.A1(new_n1277), .A2(G384), .A3(new_n1246), .ZN(new_n1278));
  AOI21_X1  g1078(.A(G384), .B1(new_n1277), .B2(new_n1246), .ZN(new_n1279));
  NOR2_X1   g1079(.A1(new_n1278), .A2(new_n1279), .ZN(new_n1280));
  INV_X1    g1080(.A(new_n1280), .ZN(new_n1281));
  OAI21_X1  g1081(.A(KEYINPUT62), .B1(new_n1268), .B2(new_n1281), .ZN(new_n1282));
  NAND3_X1  g1082(.A1(new_n674), .A2(G213), .A3(G2897), .ZN(new_n1283));
  INV_X1    g1083(.A(new_n1283), .ZN(new_n1284));
  OAI21_X1  g1084(.A(new_n1284), .B1(new_n1278), .B2(new_n1279), .ZN(new_n1285));
  NAND2_X1  g1085(.A1(new_n1277), .A2(new_n1246), .ZN(new_n1286));
  NAND2_X1  g1086(.A1(new_n1286), .A2(new_n1251), .ZN(new_n1287));
  NAND3_X1  g1087(.A1(new_n1277), .A2(G384), .A3(new_n1246), .ZN(new_n1288));
  NAND3_X1  g1088(.A1(new_n1287), .A2(new_n1288), .A3(new_n1283), .ZN(new_n1289));
  AND2_X1   g1089(.A1(new_n1285), .A2(new_n1289), .ZN(new_n1290));
  AOI21_X1  g1090(.A(KEYINPUT61), .B1(new_n1268), .B2(new_n1290), .ZN(new_n1291));
  NAND2_X1  g1091(.A1(G375), .A2(G378), .ZN(new_n1292));
  AND2_X1   g1092(.A1(new_n1267), .A2(new_n1263), .ZN(new_n1293));
  INV_X1    g1093(.A(KEYINPUT62), .ZN(new_n1294));
  NAND4_X1  g1094(.A1(new_n1292), .A2(new_n1293), .A3(new_n1294), .A4(new_n1280), .ZN(new_n1295));
  NAND3_X1  g1095(.A1(new_n1282), .A2(new_n1291), .A3(new_n1295), .ZN(new_n1296));
  XNOR2_X1  g1096(.A(new_n1026), .B(new_n1102), .ZN(new_n1297));
  XNOR2_X1  g1097(.A(G393), .B(new_n817), .ZN(new_n1298));
  INV_X1    g1098(.A(KEYINPUT127), .ZN(new_n1299));
  XNOR2_X1  g1099(.A(new_n1298), .B(new_n1299), .ZN(new_n1300));
  NOR2_X1   g1100(.A1(new_n1026), .A2(new_n1102), .ZN(new_n1301));
  NOR2_X1   g1101(.A1(new_n1301), .A2(new_n1298), .ZN(new_n1302));
  NAND3_X1  g1102(.A1(new_n1028), .A2(new_n1029), .A3(new_n1102), .ZN(new_n1303));
  AOI22_X1  g1103(.A1(new_n1297), .A2(new_n1300), .B1(new_n1302), .B2(new_n1303), .ZN(new_n1304));
  NAND2_X1  g1104(.A1(new_n1296), .A2(new_n1304), .ZN(new_n1305));
  NAND2_X1  g1105(.A1(new_n1302), .A2(new_n1303), .ZN(new_n1306));
  AND2_X1   g1106(.A1(new_n1026), .A2(new_n1102), .ZN(new_n1307));
  OAI21_X1  g1107(.A(new_n1300), .B1(new_n1307), .B2(new_n1301), .ZN(new_n1308));
  NAND2_X1  g1108(.A1(new_n1306), .A2(new_n1308), .ZN(new_n1309));
  INV_X1    g1109(.A(KEYINPUT63), .ZN(new_n1310));
  OAI21_X1  g1110(.A(new_n1310), .B1(new_n1268), .B2(new_n1281), .ZN(new_n1311));
  NAND4_X1  g1111(.A1(new_n1292), .A2(new_n1293), .A3(KEYINPUT63), .A4(new_n1280), .ZN(new_n1312));
  NAND4_X1  g1112(.A1(new_n1309), .A2(new_n1291), .A3(new_n1311), .A4(new_n1312), .ZN(new_n1313));
  NAND2_X1  g1113(.A1(new_n1305), .A2(new_n1313), .ZN(G405));
  NAND2_X1  g1114(.A1(new_n1292), .A2(new_n1261), .ZN(new_n1315));
  NAND2_X1  g1115(.A1(new_n1315), .A2(new_n1280), .ZN(new_n1316));
  NAND3_X1  g1116(.A1(new_n1292), .A2(new_n1261), .A3(new_n1281), .ZN(new_n1317));
  NAND2_X1  g1117(.A1(new_n1316), .A2(new_n1317), .ZN(new_n1318));
  NAND2_X1  g1118(.A1(new_n1318), .A2(new_n1309), .ZN(new_n1319));
  NAND3_X1  g1119(.A1(new_n1304), .A2(new_n1316), .A3(new_n1317), .ZN(new_n1320));
  NAND2_X1  g1120(.A1(new_n1319), .A2(new_n1320), .ZN(G402));
endmodule


