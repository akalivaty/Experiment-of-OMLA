//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 1 1 0 1 0 0 1 1 0 1 0 1 0 1 0 1 0 0 0 1 1 1 0 1 0 0 1 0 1 0 0 1 0 1 0 0 0 1 1 0 1 1 0 1 1 0 0 0 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:16:51 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n664, new_n665,
    new_n667, new_n668, new_n669, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n692, new_n693, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n709, new_n710, new_n711, new_n713, new_n714,
    new_n715, new_n716, new_n717, new_n718, new_n719, new_n720, new_n722,
    new_n723, new_n724, new_n725, new_n726, new_n727, new_n728, new_n729,
    new_n731, new_n732, new_n734, new_n735, new_n736, new_n737, new_n738,
    new_n739, new_n740, new_n741, new_n742, new_n743, new_n744, new_n745,
    new_n746, new_n747, new_n748, new_n749, new_n750, new_n751, new_n752,
    new_n753, new_n754, new_n755, new_n756, new_n757, new_n758, new_n759,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n769, new_n770, new_n771, new_n772, new_n773, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n841,
    new_n842, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n851, new_n852, new_n854, new_n855, new_n856, new_n857,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n917, new_n918, new_n920, new_n921, new_n922, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n935, new_n936, new_n937, new_n939, new_n940, new_n941,
    new_n943, new_n944, new_n945, new_n946, new_n947, new_n949, new_n950,
    new_n951, new_n952, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n960, new_n961, new_n962, new_n963, new_n964, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972;
  XNOR2_X1  g000(.A(G78gat), .B(G106gat), .ZN(new_n202));
  INV_X1    g001(.A(new_n202), .ZN(new_n203));
  XNOR2_X1  g002(.A(KEYINPUT75), .B(KEYINPUT31), .ZN(new_n204));
  XNOR2_X1  g003(.A(new_n204), .B(G50gat), .ZN(new_n205));
  INV_X1    g004(.A(new_n205), .ZN(new_n206));
  XOR2_X1   g005(.A(G211gat), .B(G218gat), .Z(new_n207));
  INV_X1    g006(.A(new_n207), .ZN(new_n208));
  INV_X1    g007(.A(KEYINPUT69), .ZN(new_n209));
  NOR2_X1   g008(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  XOR2_X1   g009(.A(G197gat), .B(G204gat), .Z(new_n211));
  XNOR2_X1  g010(.A(KEYINPUT68), .B(G211gat), .ZN(new_n212));
  NAND2_X1  g011(.A1(new_n212), .A2(G218gat), .ZN(new_n213));
  INV_X1    g012(.A(KEYINPUT22), .ZN(new_n214));
  AOI21_X1  g013(.A(new_n211), .B1(new_n213), .B2(new_n214), .ZN(new_n215));
  XNOR2_X1  g014(.A(new_n210), .B(new_n215), .ZN(new_n216));
  NAND2_X1  g015(.A1(new_n216), .A2(KEYINPUT70), .ZN(new_n217));
  NAND2_X1  g016(.A1(new_n213), .A2(new_n214), .ZN(new_n218));
  INV_X1    g017(.A(new_n211), .ZN(new_n219));
  NAND2_X1  g018(.A1(new_n218), .A2(new_n219), .ZN(new_n220));
  NAND2_X1  g019(.A1(new_n220), .A2(new_n210), .ZN(new_n221));
  OAI21_X1  g020(.A(new_n215), .B1(new_n209), .B2(new_n208), .ZN(new_n222));
  NAND2_X1  g021(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  INV_X1    g022(.A(KEYINPUT70), .ZN(new_n224));
  NAND2_X1  g023(.A1(new_n223), .A2(new_n224), .ZN(new_n225));
  XNOR2_X1  g024(.A(G141gat), .B(G148gat), .ZN(new_n226));
  INV_X1    g025(.A(new_n226), .ZN(new_n227));
  OR2_X1    g026(.A1(G155gat), .A2(G162gat), .ZN(new_n228));
  NAND2_X1  g027(.A1(G155gat), .A2(G162gat), .ZN(new_n229));
  NAND2_X1  g028(.A1(new_n228), .A2(new_n229), .ZN(new_n230));
  NAND2_X1  g029(.A1(new_n229), .A2(KEYINPUT2), .ZN(new_n231));
  NAND3_X1  g030(.A1(new_n227), .A2(new_n230), .A3(new_n231), .ZN(new_n232));
  OAI211_X1 g031(.A(new_n229), .B(new_n228), .C1(new_n226), .C2(KEYINPUT2), .ZN(new_n233));
  XOR2_X1   g032(.A(KEYINPUT71), .B(KEYINPUT3), .Z(new_n234));
  NAND3_X1  g033(.A1(new_n232), .A2(new_n233), .A3(new_n234), .ZN(new_n235));
  INV_X1    g034(.A(KEYINPUT29), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n235), .A2(new_n236), .ZN(new_n237));
  NAND3_X1  g036(.A1(new_n217), .A2(new_n225), .A3(new_n237), .ZN(new_n238));
  INV_X1    g037(.A(G228gat), .ZN(new_n239));
  INV_X1    g038(.A(G233gat), .ZN(new_n240));
  NOR2_X1   g039(.A1(new_n239), .A2(new_n240), .ZN(new_n241));
  NAND2_X1  g040(.A1(new_n232), .A2(new_n233), .ZN(new_n242));
  INV_X1    g041(.A(new_n242), .ZN(new_n243));
  AOI21_X1  g042(.A(KEYINPUT3), .B1(new_n223), .B2(new_n236), .ZN(new_n244));
  OAI211_X1 g043(.A(new_n238), .B(new_n241), .C1(new_n243), .C2(new_n244), .ZN(new_n245));
  NAND3_X1  g044(.A1(new_n218), .A2(new_n207), .A3(new_n219), .ZN(new_n246));
  NAND2_X1  g045(.A1(new_n246), .A2(new_n236), .ZN(new_n247));
  NOR2_X1   g046(.A1(new_n215), .A2(new_n207), .ZN(new_n248));
  OAI21_X1  g047(.A(new_n234), .B1(new_n247), .B2(new_n248), .ZN(new_n249));
  AOI22_X1  g048(.A1(new_n249), .A2(new_n242), .B1(new_n216), .B2(new_n237), .ZN(new_n250));
  NOR3_X1   g049(.A1(new_n250), .A2(KEYINPUT77), .A3(new_n241), .ZN(new_n251));
  INV_X1    g050(.A(KEYINPUT77), .ZN(new_n252));
  NAND3_X1  g051(.A1(new_n237), .A2(new_n221), .A3(new_n222), .ZN(new_n253));
  INV_X1    g052(.A(new_n234), .ZN(new_n254));
  NAND2_X1  g053(.A1(new_n220), .A2(new_n208), .ZN(new_n255));
  AOI21_X1  g054(.A(KEYINPUT29), .B1(new_n215), .B2(new_n207), .ZN(new_n256));
  AOI21_X1  g055(.A(new_n254), .B1(new_n255), .B2(new_n256), .ZN(new_n257));
  OAI21_X1  g056(.A(new_n253), .B1(new_n257), .B2(new_n243), .ZN(new_n258));
  INV_X1    g057(.A(new_n241), .ZN(new_n259));
  AOI21_X1  g058(.A(new_n252), .B1(new_n258), .B2(new_n259), .ZN(new_n260));
  OAI21_X1  g059(.A(new_n245), .B1(new_n251), .B2(new_n260), .ZN(new_n261));
  NAND2_X1  g060(.A1(new_n261), .A2(G22gat), .ZN(new_n262));
  INV_X1    g061(.A(G22gat), .ZN(new_n263));
  OAI211_X1 g062(.A(new_n245), .B(new_n263), .C1(new_n251), .C2(new_n260), .ZN(new_n264));
  NAND2_X1  g063(.A1(new_n262), .A2(new_n264), .ZN(new_n265));
  INV_X1    g064(.A(KEYINPUT76), .ZN(new_n266));
  AOI21_X1  g065(.A(new_n206), .B1(new_n265), .B2(new_n266), .ZN(new_n267));
  AOI211_X1 g066(.A(KEYINPUT76), .B(new_n205), .C1(new_n262), .C2(new_n264), .ZN(new_n268));
  OAI21_X1  g067(.A(new_n203), .B1(new_n267), .B2(new_n268), .ZN(new_n269));
  INV_X1    g068(.A(new_n264), .ZN(new_n270));
  OAI21_X1  g069(.A(KEYINPUT77), .B1(new_n250), .B2(new_n241), .ZN(new_n271));
  NAND3_X1  g070(.A1(new_n258), .A2(new_n252), .A3(new_n259), .ZN(new_n272));
  NAND2_X1  g071(.A1(new_n271), .A2(new_n272), .ZN(new_n273));
  AOI21_X1  g072(.A(new_n263), .B1(new_n273), .B2(new_n245), .ZN(new_n274));
  OAI21_X1  g073(.A(new_n266), .B1(new_n270), .B2(new_n274), .ZN(new_n275));
  NAND2_X1  g074(.A1(new_n275), .A2(new_n205), .ZN(new_n276));
  NAND3_X1  g075(.A1(new_n265), .A2(new_n266), .A3(new_n206), .ZN(new_n277));
  NAND3_X1  g076(.A1(new_n276), .A2(new_n277), .A3(new_n202), .ZN(new_n278));
  NAND2_X1  g077(.A1(new_n269), .A2(new_n278), .ZN(new_n279));
  NAND2_X1  g078(.A1(G225gat), .A2(G233gat), .ZN(new_n280));
  NAND2_X1  g079(.A1(new_n242), .A2(KEYINPUT3), .ZN(new_n281));
  XOR2_X1   g080(.A(G127gat), .B(G134gat), .Z(new_n282));
  INV_X1    g081(.A(new_n282), .ZN(new_n283));
  XNOR2_X1  g082(.A(G113gat), .B(G120gat), .ZN(new_n284));
  NOR2_X1   g083(.A1(new_n284), .A2(KEYINPUT1), .ZN(new_n285));
  NAND2_X1  g084(.A1(new_n283), .A2(new_n285), .ZN(new_n286));
  OAI21_X1  g085(.A(new_n282), .B1(KEYINPUT1), .B2(new_n284), .ZN(new_n287));
  NAND2_X1  g086(.A1(new_n286), .A2(new_n287), .ZN(new_n288));
  NAND3_X1  g087(.A1(new_n281), .A2(new_n288), .A3(new_n235), .ZN(new_n289));
  NAND4_X1  g088(.A1(new_n286), .A2(new_n232), .A3(new_n233), .A4(new_n287), .ZN(new_n290));
  NOR2_X1   g089(.A1(new_n290), .A2(KEYINPUT4), .ZN(new_n291));
  NAND2_X1  g090(.A1(new_n290), .A2(KEYINPUT4), .ZN(new_n292));
  AOI21_X1  g091(.A(new_n291), .B1(KEYINPUT72), .B2(new_n292), .ZN(new_n293));
  INV_X1    g092(.A(KEYINPUT72), .ZN(new_n294));
  NOR3_X1   g093(.A1(new_n290), .A2(new_n294), .A3(KEYINPUT4), .ZN(new_n295));
  OAI211_X1 g094(.A(new_n280), .B(new_n289), .C1(new_n293), .C2(new_n295), .ZN(new_n296));
  INV_X1    g095(.A(KEYINPUT5), .ZN(new_n297));
  NAND2_X1  g096(.A1(new_n288), .A2(new_n242), .ZN(new_n298));
  NAND2_X1  g097(.A1(new_n298), .A2(new_n290), .ZN(new_n299));
  INV_X1    g098(.A(new_n280), .ZN(new_n300));
  AOI21_X1  g099(.A(new_n297), .B1(new_n299), .B2(new_n300), .ZN(new_n301));
  NAND2_X1  g100(.A1(new_n296), .A2(new_n301), .ZN(new_n302));
  NOR2_X1   g101(.A1(new_n300), .A2(KEYINPUT5), .ZN(new_n303));
  INV_X1    g102(.A(new_n292), .ZN(new_n304));
  OAI211_X1 g103(.A(new_n289), .B(new_n303), .C1(new_n304), .C2(new_n291), .ZN(new_n305));
  NAND2_X1  g104(.A1(new_n302), .A2(new_n305), .ZN(new_n306));
  XNOR2_X1  g105(.A(G1gat), .B(G29gat), .ZN(new_n307));
  XNOR2_X1  g106(.A(new_n307), .B(KEYINPUT74), .ZN(new_n308));
  XNOR2_X1  g107(.A(G57gat), .B(G85gat), .ZN(new_n309));
  XNOR2_X1  g108(.A(new_n308), .B(new_n309), .ZN(new_n310));
  XNOR2_X1  g109(.A(KEYINPUT73), .B(KEYINPUT0), .ZN(new_n311));
  XOR2_X1   g110(.A(new_n310), .B(new_n311), .Z(new_n312));
  INV_X1    g111(.A(new_n312), .ZN(new_n313));
  NAND2_X1  g112(.A1(new_n306), .A2(new_n313), .ZN(new_n314));
  INV_X1    g113(.A(new_n305), .ZN(new_n315));
  AOI21_X1  g114(.A(new_n315), .B1(new_n296), .B2(new_n301), .ZN(new_n316));
  AOI21_X1  g115(.A(KEYINPUT6), .B1(new_n316), .B2(new_n312), .ZN(new_n317));
  NAND2_X1  g116(.A1(new_n314), .A2(new_n317), .ZN(new_n318));
  NAND3_X1  g117(.A1(new_n306), .A2(KEYINPUT6), .A3(new_n313), .ZN(new_n319));
  NAND2_X1  g118(.A1(new_n318), .A2(new_n319), .ZN(new_n320));
  INV_X1    g119(.A(new_n320), .ZN(new_n321));
  XNOR2_X1  g120(.A(KEYINPUT27), .B(G183gat), .ZN(new_n322));
  INV_X1    g121(.A(G190gat), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n322), .A2(new_n323), .ZN(new_n324));
  XNOR2_X1  g123(.A(new_n324), .B(KEYINPUT28), .ZN(new_n325));
  NOR2_X1   g124(.A1(G169gat), .A2(G176gat), .ZN(new_n326));
  NAND2_X1  g125(.A1(new_n326), .A2(KEYINPUT26), .ZN(new_n327));
  NAND2_X1  g126(.A1(G183gat), .A2(G190gat), .ZN(new_n328));
  NAND2_X1  g127(.A1(new_n327), .A2(new_n328), .ZN(new_n329));
  NAND2_X1  g128(.A1(G169gat), .A2(G176gat), .ZN(new_n330));
  INV_X1    g129(.A(KEYINPUT26), .ZN(new_n331));
  NAND2_X1  g130(.A1(new_n330), .A2(new_n331), .ZN(new_n332));
  NOR2_X1   g131(.A1(new_n332), .A2(new_n326), .ZN(new_n333));
  NOR2_X1   g132(.A1(new_n329), .A2(new_n333), .ZN(new_n334));
  INV_X1    g133(.A(new_n334), .ZN(new_n335));
  OR3_X1    g134(.A1(new_n326), .A2(KEYINPUT64), .A3(KEYINPUT23), .ZN(new_n336));
  OAI21_X1  g135(.A(KEYINPUT64), .B1(new_n326), .B2(KEYINPUT23), .ZN(new_n337));
  NAND2_X1  g136(.A1(new_n326), .A2(KEYINPUT23), .ZN(new_n338));
  NAND4_X1  g137(.A1(new_n336), .A2(new_n337), .A3(new_n338), .A4(new_n330), .ZN(new_n339));
  NOR2_X1   g138(.A1(G183gat), .A2(G190gat), .ZN(new_n340));
  INV_X1    g139(.A(new_n328), .ZN(new_n341));
  AOI21_X1  g140(.A(new_n340), .B1(new_n341), .B2(KEYINPUT24), .ZN(new_n342));
  INV_X1    g141(.A(KEYINPUT24), .ZN(new_n343));
  NAND2_X1  g142(.A1(new_n328), .A2(new_n343), .ZN(new_n344));
  AOI21_X1  g143(.A(KEYINPUT25), .B1(new_n342), .B2(new_n344), .ZN(new_n345));
  INV_X1    g144(.A(new_n345), .ZN(new_n346));
  OAI22_X1  g145(.A1(new_n325), .A2(new_n335), .B1(new_n339), .B2(new_n346), .ZN(new_n347));
  INV_X1    g146(.A(KEYINPUT25), .ZN(new_n348));
  AND2_X1   g147(.A1(new_n343), .A2(KEYINPUT65), .ZN(new_n349));
  NOR2_X1   g148(.A1(new_n343), .A2(KEYINPUT65), .ZN(new_n350));
  OAI21_X1  g149(.A(new_n328), .B1(new_n349), .B2(new_n350), .ZN(new_n351));
  INV_X1    g150(.A(KEYINPUT66), .ZN(new_n352));
  NAND2_X1  g151(.A1(new_n351), .A2(new_n352), .ZN(new_n353));
  OAI211_X1 g152(.A(KEYINPUT66), .B(new_n328), .C1(new_n349), .C2(new_n350), .ZN(new_n354));
  NAND3_X1  g153(.A1(new_n353), .A2(new_n342), .A3(new_n354), .ZN(new_n355));
  INV_X1    g154(.A(new_n339), .ZN(new_n356));
  AOI21_X1  g155(.A(new_n348), .B1(new_n355), .B2(new_n356), .ZN(new_n357));
  INV_X1    g156(.A(G226gat), .ZN(new_n358));
  NOR2_X1   g157(.A1(new_n358), .A2(new_n240), .ZN(new_n359));
  OAI22_X1  g158(.A1(new_n347), .A2(new_n357), .B1(KEYINPUT29), .B2(new_n359), .ZN(new_n360));
  INV_X1    g159(.A(new_n357), .ZN(new_n361));
  INV_X1    g160(.A(KEYINPUT28), .ZN(new_n362));
  XNOR2_X1  g161(.A(new_n324), .B(new_n362), .ZN(new_n363));
  AOI22_X1  g162(.A1(new_n363), .A2(new_n334), .B1(new_n356), .B2(new_n345), .ZN(new_n364));
  INV_X1    g163(.A(new_n359), .ZN(new_n365));
  NAND3_X1  g164(.A1(new_n361), .A2(new_n364), .A3(new_n365), .ZN(new_n366));
  AND3_X1   g165(.A1(new_n360), .A2(new_n366), .A3(new_n216), .ZN(new_n367));
  AOI22_X1  g166(.A1(new_n360), .A2(new_n366), .B1(new_n217), .B2(new_n225), .ZN(new_n368));
  OR2_X1    g167(.A1(new_n367), .A2(new_n368), .ZN(new_n369));
  XNOR2_X1  g168(.A(G8gat), .B(G36gat), .ZN(new_n370));
  XNOR2_X1  g169(.A(G64gat), .B(G92gat), .ZN(new_n371));
  XNOR2_X1  g170(.A(new_n370), .B(new_n371), .ZN(new_n372));
  INV_X1    g171(.A(new_n372), .ZN(new_n373));
  NAND2_X1  g172(.A1(new_n369), .A2(new_n373), .ZN(new_n374));
  OR3_X1    g173(.A1(new_n367), .A2(new_n368), .A3(new_n373), .ZN(new_n375));
  NAND3_X1  g174(.A1(new_n374), .A2(KEYINPUT30), .A3(new_n375), .ZN(new_n376));
  INV_X1    g175(.A(KEYINPUT30), .ZN(new_n377));
  NAND3_X1  g176(.A1(new_n369), .A2(new_n377), .A3(new_n373), .ZN(new_n378));
  NAND2_X1  g177(.A1(new_n376), .A2(new_n378), .ZN(new_n379));
  INV_X1    g178(.A(new_n379), .ZN(new_n380));
  OAI21_X1  g179(.A(new_n279), .B1(new_n321), .B2(new_n380), .ZN(new_n381));
  NAND4_X1  g180(.A1(new_n361), .A2(new_n364), .A3(new_n286), .A4(new_n287), .ZN(new_n382));
  INV_X1    g181(.A(G227gat), .ZN(new_n383));
  NOR2_X1   g182(.A1(new_n383), .A2(new_n240), .ZN(new_n384));
  INV_X1    g183(.A(new_n384), .ZN(new_n385));
  OAI21_X1  g184(.A(new_n288), .B1(new_n347), .B2(new_n357), .ZN(new_n386));
  NAND3_X1  g185(.A1(new_n382), .A2(new_n385), .A3(new_n386), .ZN(new_n387));
  XOR2_X1   g186(.A(new_n387), .B(KEYINPUT34), .Z(new_n388));
  INV_X1    g187(.A(new_n388), .ZN(new_n389));
  XNOR2_X1  g188(.A(G15gat), .B(G43gat), .ZN(new_n390));
  XNOR2_X1  g189(.A(G71gat), .B(G99gat), .ZN(new_n391));
  XOR2_X1   g190(.A(new_n390), .B(new_n391), .Z(new_n392));
  AOI21_X1  g191(.A(new_n385), .B1(new_n382), .B2(new_n386), .ZN(new_n393));
  OAI21_X1  g192(.A(new_n392), .B1(new_n393), .B2(KEYINPUT33), .ZN(new_n394));
  INV_X1    g193(.A(KEYINPUT32), .ZN(new_n395));
  NOR2_X1   g194(.A1(new_n393), .A2(new_n395), .ZN(new_n396));
  NOR2_X1   g195(.A1(new_n394), .A2(new_n396), .ZN(new_n397));
  INV_X1    g196(.A(new_n397), .ZN(new_n398));
  NAND2_X1  g197(.A1(new_n394), .A2(new_n396), .ZN(new_n399));
  NAND3_X1  g198(.A1(new_n389), .A2(new_n398), .A3(new_n399), .ZN(new_n400));
  INV_X1    g199(.A(new_n399), .ZN(new_n401));
  OAI21_X1  g200(.A(new_n388), .B1(new_n401), .B2(new_n397), .ZN(new_n402));
  NAND2_X1  g201(.A1(new_n400), .A2(new_n402), .ZN(new_n403));
  OR2_X1    g202(.A1(new_n403), .A2(KEYINPUT36), .ZN(new_n404));
  INV_X1    g203(.A(KEYINPUT67), .ZN(new_n405));
  NAND2_X1  g204(.A1(new_n389), .A2(new_n405), .ZN(new_n406));
  OAI211_X1 g205(.A(new_n400), .B(new_n406), .C1(new_n402), .C2(new_n405), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n407), .A2(KEYINPUT36), .ZN(new_n408));
  NAND2_X1  g207(.A1(new_n404), .A2(new_n408), .ZN(new_n409));
  XNOR2_X1  g208(.A(KEYINPUT79), .B(KEYINPUT37), .ZN(new_n410));
  OAI21_X1  g209(.A(new_n410), .B1(new_n367), .B2(new_n368), .ZN(new_n411));
  NAND2_X1  g210(.A1(new_n360), .A2(new_n366), .ZN(new_n412));
  NAND2_X1  g211(.A1(new_n412), .A2(new_n223), .ZN(new_n413));
  NAND4_X1  g212(.A1(new_n360), .A2(new_n366), .A3(new_n217), .A4(new_n225), .ZN(new_n414));
  NAND3_X1  g213(.A1(new_n413), .A2(new_n414), .A3(KEYINPUT37), .ZN(new_n415));
  INV_X1    g214(.A(KEYINPUT38), .ZN(new_n416));
  NAND4_X1  g215(.A1(new_n411), .A2(new_n415), .A3(new_n416), .A4(new_n372), .ZN(new_n417));
  INV_X1    g216(.A(KEYINPUT80), .ZN(new_n418));
  NAND2_X1  g217(.A1(new_n417), .A2(new_n418), .ZN(new_n419));
  AND3_X1   g218(.A1(new_n419), .A2(new_n318), .A3(new_n319), .ZN(new_n420));
  NOR2_X1   g219(.A1(new_n417), .A2(new_n418), .ZN(new_n421));
  INV_X1    g220(.A(new_n421), .ZN(new_n422));
  NAND4_X1  g221(.A1(new_n420), .A2(KEYINPUT81), .A3(new_n374), .A4(new_n422), .ZN(new_n423));
  INV_X1    g222(.A(KEYINPUT37), .ZN(new_n424));
  OAI21_X1  g223(.A(new_n411), .B1(new_n369), .B2(new_n424), .ZN(new_n425));
  OAI21_X1  g224(.A(KEYINPUT38), .B1(new_n425), .B2(new_n373), .ZN(new_n426));
  INV_X1    g225(.A(KEYINPUT81), .ZN(new_n427));
  NAND4_X1  g226(.A1(new_n419), .A2(new_n318), .A3(new_n319), .A4(new_n374), .ZN(new_n428));
  OAI21_X1  g227(.A(new_n427), .B1(new_n428), .B2(new_n421), .ZN(new_n429));
  AND3_X1   g228(.A1(new_n423), .A2(new_n426), .A3(new_n429), .ZN(new_n430));
  OAI21_X1  g229(.A(new_n289), .B1(new_n304), .B2(new_n291), .ZN(new_n431));
  NAND2_X1  g230(.A1(new_n431), .A2(new_n300), .ZN(new_n432));
  OAI211_X1 g231(.A(new_n432), .B(KEYINPUT39), .C1(new_n300), .C2(new_n299), .ZN(new_n433));
  OAI211_X1 g232(.A(new_n433), .B(new_n312), .C1(KEYINPUT39), .C2(new_n432), .ZN(new_n434));
  NAND2_X1  g233(.A1(new_n434), .A2(KEYINPUT78), .ZN(new_n435));
  OR2_X1    g234(.A1(new_n435), .A2(KEYINPUT40), .ZN(new_n436));
  NAND2_X1  g235(.A1(new_n435), .A2(KEYINPUT40), .ZN(new_n437));
  NAND4_X1  g236(.A1(new_n380), .A2(new_n314), .A3(new_n436), .A4(new_n437), .ZN(new_n438));
  NAND3_X1  g237(.A1(new_n438), .A2(new_n269), .A3(new_n278), .ZN(new_n439));
  OAI211_X1 g238(.A(new_n381), .B(new_n409), .C1(new_n430), .C2(new_n439), .ZN(new_n440));
  AND4_X1   g239(.A1(KEYINPUT35), .A2(new_n269), .A3(new_n278), .A4(new_n407), .ZN(new_n441));
  AND2_X1   g240(.A1(new_n379), .A2(new_n320), .ZN(new_n442));
  INV_X1    g241(.A(KEYINPUT35), .ZN(new_n443));
  NAND4_X1  g242(.A1(new_n269), .A2(new_n278), .A3(new_n442), .A4(new_n403), .ZN(new_n444));
  AOI22_X1  g243(.A1(new_n441), .A2(new_n442), .B1(new_n443), .B2(new_n444), .ZN(new_n445));
  NAND2_X1  g244(.A1(new_n440), .A2(new_n445), .ZN(new_n446));
  NAND3_X1  g245(.A1(KEYINPUT96), .A2(G85gat), .A3(G92gat), .ZN(new_n447));
  INV_X1    g246(.A(KEYINPUT95), .ZN(new_n448));
  NAND2_X1  g247(.A1(new_n447), .A2(new_n448), .ZN(new_n449));
  NAND3_X1  g248(.A1(KEYINPUT95), .A2(G85gat), .A3(G92gat), .ZN(new_n450));
  NAND3_X1  g249(.A1(new_n449), .A2(KEYINPUT7), .A3(new_n450), .ZN(new_n451));
  XNOR2_X1  g250(.A(G99gat), .B(G106gat), .ZN(new_n452));
  INV_X1    g251(.A(KEYINPUT7), .ZN(new_n453));
  NAND3_X1  g252(.A1(new_n447), .A2(new_n448), .A3(new_n453), .ZN(new_n454));
  NAND2_X1  g253(.A1(G99gat), .A2(G106gat), .ZN(new_n455));
  INV_X1    g254(.A(G85gat), .ZN(new_n456));
  INV_X1    g255(.A(G92gat), .ZN(new_n457));
  AOI22_X1  g256(.A1(KEYINPUT8), .A2(new_n455), .B1(new_n456), .B2(new_n457), .ZN(new_n458));
  NAND4_X1  g257(.A1(new_n451), .A2(new_n452), .A3(new_n454), .A4(new_n458), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n459), .A2(KEYINPUT97), .ZN(new_n460));
  AND2_X1   g259(.A1(new_n458), .A2(new_n454), .ZN(new_n461));
  INV_X1    g260(.A(KEYINPUT97), .ZN(new_n462));
  NAND4_X1  g261(.A1(new_n461), .A2(new_n462), .A3(new_n452), .A4(new_n451), .ZN(new_n463));
  NAND2_X1  g262(.A1(new_n460), .A2(new_n463), .ZN(new_n464));
  INV_X1    g263(.A(new_n452), .ZN(new_n465));
  AND3_X1   g264(.A1(new_n449), .A2(KEYINPUT7), .A3(new_n450), .ZN(new_n466));
  NAND2_X1  g265(.A1(new_n458), .A2(new_n454), .ZN(new_n467));
  OAI21_X1  g266(.A(new_n465), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  INV_X1    g267(.A(KEYINPUT98), .ZN(new_n469));
  NAND2_X1  g268(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  OAI211_X1 g269(.A(KEYINPUT98), .B(new_n465), .C1(new_n466), .C2(new_n467), .ZN(new_n471));
  NAND3_X1  g270(.A1(new_n464), .A2(new_n470), .A3(new_n471), .ZN(new_n472));
  INV_X1    g271(.A(new_n472), .ZN(new_n473));
  OR2_X1    g272(.A1(KEYINPUT83), .A2(KEYINPUT14), .ZN(new_n474));
  NAND2_X1  g273(.A1(KEYINPUT83), .A2(KEYINPUT14), .ZN(new_n475));
  OAI211_X1 g274(.A(new_n474), .B(new_n475), .C1(G29gat), .C2(G36gat), .ZN(new_n476));
  INV_X1    g275(.A(G29gat), .ZN(new_n477));
  INV_X1    g276(.A(G36gat), .ZN(new_n478));
  NAND4_X1  g277(.A1(new_n477), .A2(new_n478), .A3(KEYINPUT83), .A4(KEYINPUT14), .ZN(new_n479));
  OAI211_X1 g278(.A(new_n476), .B(new_n479), .C1(new_n477), .C2(new_n478), .ZN(new_n480));
  XNOR2_X1  g279(.A(G43gat), .B(G50gat), .ZN(new_n481));
  OR2_X1    g280(.A1(new_n481), .A2(KEYINPUT15), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n481), .A2(KEYINPUT82), .ZN(new_n483));
  INV_X1    g282(.A(KEYINPUT82), .ZN(new_n484));
  INV_X1    g283(.A(G43gat), .ZN(new_n485));
  NOR2_X1   g284(.A1(new_n485), .A2(G50gat), .ZN(new_n486));
  INV_X1    g285(.A(G50gat), .ZN(new_n487));
  NOR2_X1   g286(.A1(new_n487), .A2(G43gat), .ZN(new_n488));
  OAI21_X1  g287(.A(new_n484), .B1(new_n486), .B2(new_n488), .ZN(new_n489));
  NAND3_X1  g288(.A1(new_n483), .A2(new_n489), .A3(KEYINPUT15), .ZN(new_n490));
  AOI21_X1  g289(.A(new_n480), .B1(new_n482), .B2(new_n490), .ZN(new_n491));
  AND2_X1   g290(.A1(new_n480), .A2(new_n490), .ZN(new_n492));
  NOR2_X1   g291(.A1(new_n491), .A2(new_n492), .ZN(new_n493));
  AND2_X1   g292(.A1(G232gat), .A2(G233gat), .ZN(new_n494));
  AOI22_X1  g293(.A1(new_n473), .A2(new_n493), .B1(KEYINPUT41), .B2(new_n494), .ZN(new_n495));
  OAI21_X1  g294(.A(KEYINPUT17), .B1(new_n491), .B2(new_n492), .ZN(new_n496));
  INV_X1    g295(.A(KEYINPUT17), .ZN(new_n497));
  NAND2_X1  g296(.A1(new_n480), .A2(new_n490), .ZN(new_n498));
  AND2_X1   g297(.A1(new_n490), .A2(new_n482), .ZN(new_n499));
  OAI211_X1 g298(.A(new_n497), .B(new_n498), .C1(new_n499), .C2(new_n480), .ZN(new_n500));
  NAND3_X1  g299(.A1(new_n496), .A2(new_n472), .A3(new_n500), .ZN(new_n501));
  XNOR2_X1  g300(.A(G190gat), .B(G218gat), .ZN(new_n502));
  INV_X1    g301(.A(new_n502), .ZN(new_n503));
  NAND3_X1  g302(.A1(new_n495), .A2(new_n501), .A3(new_n503), .ZN(new_n504));
  INV_X1    g303(.A(new_n504), .ZN(new_n505));
  NOR2_X1   g304(.A1(new_n494), .A2(KEYINPUT41), .ZN(new_n506));
  XNOR2_X1  g305(.A(G134gat), .B(G162gat), .ZN(new_n507));
  XOR2_X1   g306(.A(new_n506), .B(new_n507), .Z(new_n508));
  INV_X1    g307(.A(new_n508), .ZN(new_n509));
  AOI21_X1  g308(.A(new_n503), .B1(new_n495), .B2(new_n501), .ZN(new_n510));
  OR3_X1    g309(.A1(new_n505), .A2(new_n509), .A3(new_n510), .ZN(new_n511));
  OAI21_X1  g310(.A(new_n509), .B1(new_n505), .B2(new_n510), .ZN(new_n512));
  NAND2_X1  g311(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  NAND2_X1  g312(.A1(G71gat), .A2(G78gat), .ZN(new_n514));
  INV_X1    g313(.A(G71gat), .ZN(new_n515));
  INV_X1    g314(.A(G78gat), .ZN(new_n516));
  NAND2_X1  g315(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  XNOR2_X1  g316(.A(G57gat), .B(G64gat), .ZN(new_n518));
  INV_X1    g317(.A(KEYINPUT9), .ZN(new_n519));
  OAI211_X1 g318(.A(new_n514), .B(new_n517), .C1(new_n518), .C2(new_n519), .ZN(new_n520));
  NAND3_X1  g319(.A1(new_n515), .A2(new_n516), .A3(KEYINPUT9), .ZN(new_n521));
  NAND2_X1  g320(.A1(new_n521), .A2(new_n514), .ZN(new_n522));
  INV_X1    g321(.A(KEYINPUT89), .ZN(new_n523));
  NAND2_X1  g322(.A1(new_n523), .A2(G57gat), .ZN(new_n524));
  INV_X1    g323(.A(G64gat), .ZN(new_n525));
  NAND2_X1  g324(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  NAND2_X1  g325(.A1(new_n522), .A2(new_n526), .ZN(new_n527));
  NAND3_X1  g326(.A1(new_n523), .A2(KEYINPUT88), .A3(G57gat), .ZN(new_n528));
  OR2_X1    g327(.A1(KEYINPUT88), .A2(G57gat), .ZN(new_n529));
  AOI21_X1  g328(.A(new_n525), .B1(new_n528), .B2(new_n529), .ZN(new_n530));
  OAI21_X1  g329(.A(new_n520), .B1(new_n527), .B2(new_n530), .ZN(new_n531));
  XOR2_X1   g330(.A(KEYINPUT90), .B(KEYINPUT21), .Z(new_n532));
  NAND2_X1  g331(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  NAND2_X1  g332(.A1(new_n531), .A2(KEYINPUT93), .ZN(new_n534));
  AOI22_X1  g333(.A1(new_n521), .A2(new_n514), .B1(new_n524), .B2(new_n525), .ZN(new_n535));
  NAND2_X1  g334(.A1(new_n528), .A2(new_n529), .ZN(new_n536));
  NAND2_X1  g335(.A1(new_n536), .A2(G64gat), .ZN(new_n537));
  AND2_X1   g336(.A1(new_n525), .A2(G57gat), .ZN(new_n538));
  NOR2_X1   g337(.A1(new_n525), .A2(G57gat), .ZN(new_n539));
  OAI21_X1  g338(.A(KEYINPUT9), .B1(new_n538), .B2(new_n539), .ZN(new_n540));
  AND2_X1   g339(.A1(new_n517), .A2(new_n514), .ZN(new_n541));
  AOI22_X1  g340(.A1(new_n535), .A2(new_n537), .B1(new_n540), .B2(new_n541), .ZN(new_n542));
  INV_X1    g341(.A(KEYINPUT93), .ZN(new_n543));
  NAND2_X1  g342(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  NAND2_X1  g343(.A1(new_n534), .A2(new_n544), .ZN(new_n545));
  NAND2_X1  g344(.A1(new_n545), .A2(KEYINPUT21), .ZN(new_n546));
  INV_X1    g345(.A(KEYINPUT94), .ZN(new_n547));
  INV_X1    g346(.A(G15gat), .ZN(new_n548));
  NAND2_X1  g347(.A1(new_n548), .A2(new_n263), .ZN(new_n549));
  NAND2_X1  g348(.A1(G15gat), .A2(G22gat), .ZN(new_n550));
  NAND2_X1  g349(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  NAND2_X1  g350(.A1(new_n551), .A2(KEYINPUT84), .ZN(new_n552));
  AOI21_X1  g351(.A(KEYINPUT16), .B1(new_n549), .B2(new_n550), .ZN(new_n553));
  OAI21_X1  g352(.A(new_n552), .B1(G1gat), .B2(new_n553), .ZN(new_n554));
  XOR2_X1   g353(.A(KEYINPUT85), .B(G8gat), .Z(new_n555));
  INV_X1    g354(.A(G1gat), .ZN(new_n556));
  NAND4_X1  g355(.A1(new_n551), .A2(KEYINPUT84), .A3(KEYINPUT16), .A4(new_n556), .ZN(new_n557));
  AND3_X1   g356(.A1(new_n554), .A2(new_n555), .A3(new_n557), .ZN(new_n558));
  INV_X1    g357(.A(G8gat), .ZN(new_n559));
  NOR2_X1   g358(.A1(new_n559), .A2(KEYINPUT85), .ZN(new_n560));
  AOI21_X1  g359(.A(new_n560), .B1(new_n554), .B2(new_n557), .ZN(new_n561));
  NOR2_X1   g360(.A1(new_n558), .A2(new_n561), .ZN(new_n562));
  NAND3_X1  g361(.A1(new_n546), .A2(new_n547), .A3(new_n562), .ZN(new_n563));
  INV_X1    g362(.A(KEYINPUT21), .ZN(new_n564));
  AOI21_X1  g363(.A(new_n564), .B1(new_n534), .B2(new_n544), .ZN(new_n565));
  NAND3_X1  g364(.A1(new_n554), .A2(new_n555), .A3(new_n557), .ZN(new_n566));
  AND2_X1   g365(.A1(new_n554), .A2(new_n557), .ZN(new_n567));
  OAI21_X1  g366(.A(new_n566), .B1(new_n567), .B2(new_n560), .ZN(new_n568));
  OAI21_X1  g367(.A(KEYINPUT94), .B1(new_n565), .B2(new_n568), .ZN(new_n569));
  XOR2_X1   g368(.A(KEYINPUT92), .B(KEYINPUT19), .Z(new_n570));
  INV_X1    g369(.A(new_n570), .ZN(new_n571));
  AND3_X1   g370(.A1(new_n563), .A2(new_n569), .A3(new_n571), .ZN(new_n572));
  AOI21_X1  g371(.A(new_n571), .B1(new_n563), .B2(new_n569), .ZN(new_n573));
  OAI21_X1  g372(.A(new_n533), .B1(new_n572), .B2(new_n573), .ZN(new_n574));
  NAND2_X1  g373(.A1(new_n563), .A2(new_n569), .ZN(new_n575));
  NAND2_X1  g374(.A1(new_n575), .A2(new_n570), .ZN(new_n576));
  INV_X1    g375(.A(new_n533), .ZN(new_n577));
  NAND3_X1  g376(.A1(new_n563), .A2(new_n569), .A3(new_n571), .ZN(new_n578));
  NAND3_X1  g377(.A1(new_n576), .A2(new_n577), .A3(new_n578), .ZN(new_n579));
  XOR2_X1   g378(.A(G127gat), .B(G155gat), .Z(new_n580));
  INV_X1    g379(.A(new_n580), .ZN(new_n581));
  AND3_X1   g380(.A1(new_n574), .A2(new_n579), .A3(new_n581), .ZN(new_n582));
  AOI21_X1  g381(.A(new_n581), .B1(new_n574), .B2(new_n579), .ZN(new_n583));
  XOR2_X1   g382(.A(G183gat), .B(G211gat), .Z(new_n584));
  NAND2_X1  g383(.A1(G231gat), .A2(G233gat), .ZN(new_n585));
  XNOR2_X1  g384(.A(new_n584), .B(new_n585), .ZN(new_n586));
  XNOR2_X1  g385(.A(KEYINPUT91), .B(KEYINPUT20), .ZN(new_n587));
  XOR2_X1   g386(.A(new_n586), .B(new_n587), .Z(new_n588));
  INV_X1    g387(.A(new_n588), .ZN(new_n589));
  NOR3_X1   g388(.A1(new_n582), .A2(new_n583), .A3(new_n589), .ZN(new_n590));
  NOR3_X1   g389(.A1(new_n572), .A2(new_n573), .A3(new_n533), .ZN(new_n591));
  AOI21_X1  g390(.A(new_n577), .B1(new_n576), .B2(new_n578), .ZN(new_n592));
  OAI21_X1  g391(.A(new_n580), .B1(new_n591), .B2(new_n592), .ZN(new_n593));
  NAND3_X1  g392(.A1(new_n574), .A2(new_n579), .A3(new_n581), .ZN(new_n594));
  AOI21_X1  g393(.A(new_n588), .B1(new_n593), .B2(new_n594), .ZN(new_n595));
  OAI21_X1  g394(.A(new_n513), .B1(new_n590), .B2(new_n595), .ZN(new_n596));
  INV_X1    g395(.A(KEYINPUT99), .ZN(new_n597));
  NAND2_X1  g396(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  OAI21_X1  g397(.A(new_n589), .B1(new_n582), .B2(new_n583), .ZN(new_n599));
  NAND3_X1  g398(.A1(new_n593), .A2(new_n594), .A3(new_n588), .ZN(new_n600));
  NAND2_X1  g399(.A1(new_n599), .A2(new_n600), .ZN(new_n601));
  NAND3_X1  g400(.A1(new_n601), .A2(KEYINPUT99), .A3(new_n513), .ZN(new_n602));
  AND2_X1   g401(.A1(new_n598), .A2(new_n602), .ZN(new_n603));
  AND2_X1   g402(.A1(new_n446), .A2(new_n603), .ZN(new_n604));
  XNOR2_X1  g403(.A(G113gat), .B(G141gat), .ZN(new_n605));
  INV_X1    g404(.A(G197gat), .ZN(new_n606));
  XNOR2_X1  g405(.A(new_n605), .B(new_n606), .ZN(new_n607));
  XNOR2_X1  g406(.A(KEYINPUT11), .B(G169gat), .ZN(new_n608));
  XNOR2_X1  g407(.A(new_n607), .B(new_n608), .ZN(new_n609));
  XNOR2_X1  g408(.A(new_n609), .B(KEYINPUT12), .ZN(new_n610));
  NAND3_X1  g409(.A1(new_n496), .A2(new_n500), .A3(new_n562), .ZN(new_n611));
  NAND2_X1  g410(.A1(G229gat), .A2(G233gat), .ZN(new_n612));
  NAND2_X1  g411(.A1(new_n568), .A2(new_n493), .ZN(new_n613));
  NAND3_X1  g412(.A1(new_n611), .A2(new_n612), .A3(new_n613), .ZN(new_n614));
  XOR2_X1   g413(.A(KEYINPUT86), .B(KEYINPUT18), .Z(new_n615));
  NAND2_X1  g414(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  AOI21_X1  g415(.A(new_n610), .B1(new_n616), .B2(KEYINPUT87), .ZN(new_n617));
  OAI21_X1  g416(.A(new_n498), .B1(new_n499), .B2(new_n480), .ZN(new_n618));
  NAND2_X1  g417(.A1(new_n562), .A2(new_n618), .ZN(new_n619));
  NAND2_X1  g418(.A1(new_n613), .A2(new_n619), .ZN(new_n620));
  XNOR2_X1  g419(.A(new_n612), .B(KEYINPUT13), .ZN(new_n621));
  INV_X1    g420(.A(new_n621), .ZN(new_n622));
  NAND2_X1  g421(.A1(new_n620), .A2(new_n622), .ZN(new_n623));
  NAND4_X1  g422(.A1(new_n611), .A2(KEYINPUT18), .A3(new_n612), .A4(new_n613), .ZN(new_n624));
  NAND3_X1  g423(.A1(new_n616), .A2(new_n623), .A3(new_n624), .ZN(new_n625));
  XNOR2_X1  g424(.A(new_n617), .B(new_n625), .ZN(new_n626));
  INV_X1    g425(.A(new_n626), .ZN(new_n627));
  XNOR2_X1  g426(.A(G120gat), .B(G148gat), .ZN(new_n628));
  XNOR2_X1  g427(.A(G176gat), .B(G204gat), .ZN(new_n629));
  XNOR2_X1  g428(.A(new_n628), .B(new_n629), .ZN(new_n630));
  NAND2_X1  g429(.A1(G230gat), .A2(G233gat), .ZN(new_n631));
  INV_X1    g430(.A(new_n631), .ZN(new_n632));
  NAND2_X1  g431(.A1(new_n472), .A2(new_n531), .ZN(new_n633));
  INV_X1    g432(.A(KEYINPUT100), .ZN(new_n634));
  NAND2_X1  g433(.A1(new_n468), .A2(new_n634), .ZN(new_n635));
  OAI211_X1 g434(.A(KEYINPUT100), .B(new_n465), .C1(new_n466), .C2(new_n467), .ZN(new_n636));
  NAND4_X1  g435(.A1(new_n464), .A2(new_n542), .A3(new_n635), .A4(new_n636), .ZN(new_n637));
  XNOR2_X1  g436(.A(KEYINPUT101), .B(KEYINPUT10), .ZN(new_n638));
  NAND3_X1  g437(.A1(new_n633), .A2(new_n637), .A3(new_n638), .ZN(new_n639));
  NAND3_X1  g438(.A1(new_n473), .A2(KEYINPUT10), .A3(new_n545), .ZN(new_n640));
  AOI21_X1  g439(.A(new_n632), .B1(new_n639), .B2(new_n640), .ZN(new_n641));
  AOI21_X1  g440(.A(new_n631), .B1(new_n633), .B2(new_n637), .ZN(new_n642));
  OAI21_X1  g441(.A(new_n630), .B1(new_n641), .B2(new_n642), .ZN(new_n643));
  NAND2_X1  g442(.A1(new_n639), .A2(new_n640), .ZN(new_n644));
  AOI21_X1  g443(.A(new_n642), .B1(new_n644), .B2(new_n631), .ZN(new_n645));
  INV_X1    g444(.A(new_n630), .ZN(new_n646));
  AOI21_X1  g445(.A(KEYINPUT102), .B1(new_n645), .B2(new_n646), .ZN(new_n647));
  INV_X1    g446(.A(KEYINPUT102), .ZN(new_n648));
  NOR4_X1   g447(.A1(new_n641), .A2(new_n648), .A3(new_n642), .A4(new_n630), .ZN(new_n649));
  OAI21_X1  g448(.A(new_n643), .B1(new_n647), .B2(new_n649), .ZN(new_n650));
  NOR2_X1   g449(.A1(new_n627), .A2(new_n650), .ZN(new_n651));
  NAND2_X1  g450(.A1(new_n604), .A2(new_n651), .ZN(new_n652));
  NOR2_X1   g451(.A1(new_n652), .A2(new_n320), .ZN(new_n653));
  XNOR2_X1  g452(.A(new_n653), .B(new_n556), .ZN(G1324gat));
  INV_X1    g453(.A(new_n652), .ZN(new_n655));
  NAND2_X1  g454(.A1(new_n655), .A2(new_n380), .ZN(new_n656));
  XNOR2_X1  g455(.A(KEYINPUT103), .B(KEYINPUT16), .ZN(new_n657));
  XNOR2_X1  g456(.A(new_n657), .B(G8gat), .ZN(new_n658));
  NOR3_X1   g457(.A1(new_n656), .A2(KEYINPUT42), .A3(new_n658), .ZN(new_n659));
  INV_X1    g458(.A(KEYINPUT42), .ZN(new_n660));
  AOI21_X1  g459(.A(new_n660), .B1(new_n656), .B2(G8gat), .ZN(new_n661));
  OR2_X1    g460(.A1(new_n656), .A2(new_n658), .ZN(new_n662));
  AOI21_X1  g461(.A(new_n659), .B1(new_n661), .B2(new_n662), .ZN(G1325gat));
  NOR3_X1   g462(.A1(new_n652), .A2(new_n548), .A3(new_n409), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n655), .A2(new_n403), .ZN(new_n665));
  AOI21_X1  g464(.A(new_n664), .B1(new_n548), .B2(new_n665), .ZN(G1326gat));
  INV_X1    g465(.A(new_n279), .ZN(new_n667));
  NOR2_X1   g466(.A1(new_n652), .A2(new_n667), .ZN(new_n668));
  XOR2_X1   g467(.A(KEYINPUT43), .B(G22gat), .Z(new_n669));
  XNOR2_X1  g468(.A(new_n668), .B(new_n669), .ZN(G1327gat));
  AOI21_X1  g469(.A(new_n513), .B1(new_n440), .B2(new_n445), .ZN(new_n671));
  INV_X1    g470(.A(new_n601), .ZN(new_n672));
  NAND2_X1  g471(.A1(new_n672), .A2(new_n651), .ZN(new_n673));
  INV_X1    g472(.A(new_n673), .ZN(new_n674));
  NAND2_X1  g473(.A1(new_n671), .A2(new_n674), .ZN(new_n675));
  NOR3_X1   g474(.A1(new_n675), .A2(G29gat), .A3(new_n320), .ZN(new_n676));
  XNOR2_X1  g475(.A(KEYINPUT104), .B(KEYINPUT45), .ZN(new_n677));
  XNOR2_X1  g476(.A(new_n676), .B(new_n677), .ZN(new_n678));
  INV_X1    g477(.A(KEYINPUT44), .ZN(new_n679));
  INV_X1    g478(.A(new_n513), .ZN(new_n680));
  AOI21_X1  g479(.A(new_n679), .B1(new_n446), .B2(new_n680), .ZN(new_n681));
  AOI211_X1 g480(.A(KEYINPUT44), .B(new_n513), .C1(new_n440), .C2(new_n445), .ZN(new_n682));
  OR2_X1    g481(.A1(new_n681), .A2(new_n682), .ZN(new_n683));
  NAND3_X1  g482(.A1(new_n683), .A2(new_n321), .A3(new_n674), .ZN(new_n684));
  INV_X1    g483(.A(new_n684), .ZN(new_n685));
  OAI21_X1  g484(.A(new_n678), .B1(new_n685), .B2(new_n477), .ZN(G1328gat));
  NAND3_X1  g485(.A1(new_n683), .A2(new_n380), .A3(new_n674), .ZN(new_n687));
  INV_X1    g486(.A(KEYINPUT105), .ZN(new_n688));
  NAND2_X1  g487(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  NAND4_X1  g488(.A1(new_n683), .A2(KEYINPUT105), .A3(new_n380), .A4(new_n674), .ZN(new_n690));
  NAND3_X1  g489(.A1(new_n689), .A2(G36gat), .A3(new_n690), .ZN(new_n691));
  NOR3_X1   g490(.A1(new_n675), .A2(G36gat), .A3(new_n379), .ZN(new_n692));
  XNOR2_X1  g491(.A(new_n692), .B(KEYINPUT46), .ZN(new_n693));
  NAND2_X1  g492(.A1(new_n691), .A2(new_n693), .ZN(G1329gat));
  INV_X1    g493(.A(new_n403), .ZN(new_n695));
  OAI21_X1  g494(.A(new_n485), .B1(new_n675), .B2(new_n695), .ZN(new_n696));
  NAND3_X1  g495(.A1(new_n683), .A2(G43gat), .A3(new_n674), .ZN(new_n697));
  OAI21_X1  g496(.A(new_n696), .B1(new_n697), .B2(new_n409), .ZN(new_n698));
  NAND2_X1  g497(.A1(new_n698), .A2(KEYINPUT47), .ZN(new_n699));
  INV_X1    g498(.A(KEYINPUT47), .ZN(new_n700));
  OAI211_X1 g499(.A(new_n700), .B(new_n696), .C1(new_n697), .C2(new_n409), .ZN(new_n701));
  NAND2_X1  g500(.A1(new_n699), .A2(new_n701), .ZN(G1330gat));
  OAI211_X1 g501(.A(new_n279), .B(new_n674), .C1(new_n681), .C2(new_n682), .ZN(new_n703));
  NAND2_X1  g502(.A1(new_n703), .A2(G50gat), .ZN(new_n704));
  NAND4_X1  g503(.A1(new_n671), .A2(new_n487), .A3(new_n279), .A4(new_n674), .ZN(new_n705));
  AOI21_X1  g504(.A(KEYINPUT106), .B1(new_n704), .B2(new_n705), .ZN(new_n706));
  INV_X1    g505(.A(KEYINPUT48), .ZN(new_n707));
  XNOR2_X1  g506(.A(new_n706), .B(new_n707), .ZN(G1331gat));
  NAND4_X1  g507(.A1(new_n446), .A2(new_n627), .A3(new_n650), .A4(new_n603), .ZN(new_n709));
  NOR2_X1   g508(.A1(new_n709), .A2(new_n320), .ZN(new_n710));
  XOR2_X1   g509(.A(KEYINPUT88), .B(G57gat), .Z(new_n711));
  XNOR2_X1  g510(.A(new_n710), .B(new_n711), .ZN(G1332gat));
  XNOR2_X1  g511(.A(new_n379), .B(KEYINPUT108), .ZN(new_n713));
  NOR2_X1   g512(.A1(new_n709), .A2(KEYINPUT107), .ZN(new_n714));
  INV_X1    g513(.A(new_n714), .ZN(new_n715));
  NAND2_X1  g514(.A1(new_n709), .A2(KEYINPUT107), .ZN(new_n716));
  AOI21_X1  g515(.A(new_n713), .B1(new_n715), .B2(new_n716), .ZN(new_n717));
  NOR2_X1   g516(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n718));
  AND2_X1   g517(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n719));
  OAI21_X1  g518(.A(new_n717), .B1(new_n718), .B2(new_n719), .ZN(new_n720));
  OAI21_X1  g519(.A(new_n720), .B1(new_n717), .B2(new_n718), .ZN(G1333gat));
  INV_X1    g520(.A(new_n409), .ZN(new_n722));
  INV_X1    g521(.A(new_n716), .ZN(new_n723));
  OAI211_X1 g522(.A(G71gat), .B(new_n722), .C1(new_n723), .C2(new_n714), .ZN(new_n724));
  NOR2_X1   g523(.A1(new_n709), .A2(new_n695), .ZN(new_n725));
  OAI21_X1  g524(.A(new_n724), .B1(G71gat), .B2(new_n725), .ZN(new_n726));
  NAND2_X1  g525(.A1(new_n726), .A2(KEYINPUT50), .ZN(new_n727));
  INV_X1    g526(.A(KEYINPUT50), .ZN(new_n728));
  OAI211_X1 g527(.A(new_n724), .B(new_n728), .C1(G71gat), .C2(new_n725), .ZN(new_n729));
  NAND2_X1  g528(.A1(new_n727), .A2(new_n729), .ZN(G1334gat));
  OAI21_X1  g529(.A(new_n279), .B1(new_n723), .B2(new_n714), .ZN(new_n731));
  XOR2_X1   g530(.A(KEYINPUT109), .B(G78gat), .Z(new_n732));
  XNOR2_X1  g531(.A(new_n731), .B(new_n732), .ZN(G1335gat));
  NOR2_X1   g532(.A1(new_n601), .A2(new_n626), .ZN(new_n734));
  OAI211_X1 g533(.A(new_n650), .B(new_n734), .C1(new_n681), .C2(new_n682), .ZN(new_n735));
  INV_X1    g534(.A(KEYINPUT110), .ZN(new_n736));
  OR3_X1    g535(.A1(new_n735), .A2(new_n736), .A3(new_n320), .ZN(new_n737));
  OAI21_X1  g536(.A(new_n736), .B1(new_n735), .B2(new_n320), .ZN(new_n738));
  NAND3_X1  g537(.A1(new_n737), .A2(G85gat), .A3(new_n738), .ZN(new_n739));
  INV_X1    g538(.A(new_n643), .ZN(new_n740));
  INV_X1    g539(.A(new_n642), .ZN(new_n741));
  NAND2_X1  g540(.A1(new_n545), .A2(KEYINPUT10), .ZN(new_n742));
  NOR2_X1   g541(.A1(new_n742), .A2(new_n472), .ZN(new_n743));
  NAND2_X1  g542(.A1(new_n636), .A2(new_n542), .ZN(new_n744));
  AOI21_X1  g543(.A(new_n744), .B1(new_n460), .B2(new_n463), .ZN(new_n745));
  AOI22_X1  g544(.A1(new_n745), .A2(new_n635), .B1(new_n472), .B2(new_n531), .ZN(new_n746));
  AOI21_X1  g545(.A(new_n743), .B1(new_n746), .B2(new_n638), .ZN(new_n747));
  OAI211_X1 g546(.A(new_n741), .B(new_n646), .C1(new_n747), .C2(new_n632), .ZN(new_n748));
  NAND2_X1  g547(.A1(new_n748), .A2(new_n648), .ZN(new_n749));
  NAND3_X1  g548(.A1(new_n645), .A2(KEYINPUT102), .A3(new_n646), .ZN(new_n750));
  AOI21_X1  g549(.A(new_n740), .B1(new_n749), .B2(new_n750), .ZN(new_n751));
  NAND2_X1  g550(.A1(new_n671), .A2(new_n734), .ZN(new_n752));
  INV_X1    g551(.A(KEYINPUT51), .ZN(new_n753));
  NOR2_X1   g552(.A1(new_n753), .A2(KEYINPUT111), .ZN(new_n754));
  AOI21_X1  g553(.A(new_n751), .B1(new_n752), .B2(new_n754), .ZN(new_n755));
  INV_X1    g554(.A(new_n754), .ZN(new_n756));
  NAND2_X1  g555(.A1(new_n753), .A2(KEYINPUT111), .ZN(new_n757));
  NAND4_X1  g556(.A1(new_n671), .A2(new_n734), .A3(new_n756), .A4(new_n757), .ZN(new_n758));
  NAND3_X1  g557(.A1(new_n755), .A2(new_n456), .A3(new_n758), .ZN(new_n759));
  OAI21_X1  g558(.A(new_n739), .B1(new_n320), .B2(new_n759), .ZN(G1336gat));
  OAI21_X1  g559(.A(G92gat), .B1(new_n735), .B2(new_n713), .ZN(new_n761));
  INV_X1    g560(.A(KEYINPUT52), .ZN(new_n762));
  INV_X1    g561(.A(new_n713), .ZN(new_n763));
  NAND4_X1  g562(.A1(new_n755), .A2(new_n457), .A3(new_n763), .A4(new_n758), .ZN(new_n764));
  NAND3_X1  g563(.A1(new_n761), .A2(new_n762), .A3(new_n764), .ZN(new_n765));
  OAI21_X1  g564(.A(G92gat), .B1(new_n735), .B2(new_n379), .ZN(new_n766));
  AND2_X1   g565(.A1(new_n766), .A2(new_n764), .ZN(new_n767));
  OAI21_X1  g566(.A(new_n765), .B1(new_n767), .B2(new_n762), .ZN(G1337gat));
  OAI21_X1  g567(.A(G99gat), .B1(new_n735), .B2(new_n409), .ZN(new_n769));
  INV_X1    g568(.A(G99gat), .ZN(new_n770));
  NAND4_X1  g569(.A1(new_n755), .A2(new_n770), .A3(new_n403), .A4(new_n758), .ZN(new_n771));
  NAND2_X1  g570(.A1(new_n769), .A2(new_n771), .ZN(new_n772));
  INV_X1    g571(.A(KEYINPUT112), .ZN(new_n773));
  XNOR2_X1  g572(.A(new_n772), .B(new_n773), .ZN(G1338gat));
  OAI21_X1  g573(.A(G106gat), .B1(new_n735), .B2(new_n667), .ZN(new_n775));
  INV_X1    g574(.A(G106gat), .ZN(new_n776));
  NAND4_X1  g575(.A1(new_n755), .A2(new_n776), .A3(new_n279), .A4(new_n758), .ZN(new_n777));
  AOI211_X1 g576(.A(KEYINPUT113), .B(KEYINPUT53), .C1(new_n775), .C2(new_n777), .ZN(new_n778));
  OR2_X1    g577(.A1(KEYINPUT113), .A2(KEYINPUT53), .ZN(new_n779));
  NAND2_X1  g578(.A1(KEYINPUT113), .A2(KEYINPUT53), .ZN(new_n780));
  AND4_X1   g579(.A1(new_n779), .A2(new_n775), .A3(new_n780), .A4(new_n777), .ZN(new_n781));
  NOR2_X1   g580(.A1(new_n778), .A2(new_n781), .ZN(G1339gat));
  NOR2_X1   g581(.A1(new_n650), .A2(new_n626), .ZN(new_n783));
  NAND3_X1  g582(.A1(new_n598), .A2(new_n602), .A3(new_n783), .ZN(new_n784));
  INV_X1    g583(.A(new_n784), .ZN(new_n785));
  AOI21_X1  g584(.A(new_n612), .B1(new_n611), .B2(new_n613), .ZN(new_n786));
  AND3_X1   g585(.A1(new_n613), .A2(new_n619), .A3(new_n621), .ZN(new_n787));
  OAI21_X1  g586(.A(new_n609), .B1(new_n786), .B2(new_n787), .ZN(new_n788));
  NAND2_X1  g587(.A1(new_n788), .A2(KEYINPUT116), .ZN(new_n789));
  NAND4_X1  g588(.A1(new_n616), .A2(new_n623), .A3(new_n610), .A4(new_n624), .ZN(new_n790));
  INV_X1    g589(.A(KEYINPUT116), .ZN(new_n791));
  OAI211_X1 g590(.A(new_n791), .B(new_n609), .C1(new_n786), .C2(new_n787), .ZN(new_n792));
  NAND3_X1  g591(.A1(new_n789), .A2(new_n790), .A3(new_n792), .ZN(new_n793));
  INV_X1    g592(.A(KEYINPUT118), .ZN(new_n794));
  NOR3_X1   g593(.A1(new_n751), .A2(new_n793), .A3(new_n794), .ZN(new_n795));
  INV_X1    g594(.A(new_n793), .ZN(new_n796));
  AOI21_X1  g595(.A(KEYINPUT118), .B1(new_n650), .B2(new_n796), .ZN(new_n797));
  NOR2_X1   g596(.A1(new_n795), .A2(new_n797), .ZN(new_n798));
  INV_X1    g597(.A(KEYINPUT54), .ZN(new_n799));
  NAND3_X1  g598(.A1(new_n644), .A2(new_n799), .A3(new_n631), .ZN(new_n800));
  NAND2_X1  g599(.A1(new_n800), .A2(new_n630), .ZN(new_n801));
  NAND3_X1  g600(.A1(new_n639), .A2(new_n632), .A3(new_n640), .ZN(new_n802));
  INV_X1    g601(.A(KEYINPUT114), .ZN(new_n803));
  AOI21_X1  g602(.A(new_n799), .B1(new_n802), .B2(new_n803), .ZN(new_n804));
  AND3_X1   g603(.A1(new_n639), .A2(new_n632), .A3(new_n640), .ZN(new_n805));
  AOI21_X1  g604(.A(new_n641), .B1(new_n805), .B2(KEYINPUT114), .ZN(new_n806));
  AOI21_X1  g605(.A(new_n801), .B1(new_n804), .B2(new_n806), .ZN(new_n807));
  AOI22_X1  g606(.A1(new_n807), .A2(KEYINPUT55), .B1(new_n749), .B2(new_n750), .ZN(new_n808));
  INV_X1    g607(.A(KEYINPUT115), .ZN(new_n809));
  NAND2_X1  g608(.A1(new_n802), .A2(new_n803), .ZN(new_n810));
  NAND2_X1  g609(.A1(new_n644), .A2(new_n631), .ZN(new_n811));
  NAND4_X1  g610(.A1(new_n639), .A2(new_n640), .A3(KEYINPUT114), .A4(new_n632), .ZN(new_n812));
  NAND4_X1  g611(.A1(new_n810), .A2(new_n811), .A3(KEYINPUT54), .A4(new_n812), .ZN(new_n813));
  AOI21_X1  g612(.A(new_n646), .B1(new_n641), .B2(new_n799), .ZN(new_n814));
  NAND2_X1  g613(.A1(new_n813), .A2(new_n814), .ZN(new_n815));
  INV_X1    g614(.A(KEYINPUT55), .ZN(new_n816));
  AOI21_X1  g615(.A(new_n809), .B1(new_n815), .B2(new_n816), .ZN(new_n817));
  AOI211_X1 g616(.A(KEYINPUT115), .B(KEYINPUT55), .C1(new_n813), .C2(new_n814), .ZN(new_n818));
  OAI211_X1 g617(.A(new_n808), .B(new_n626), .C1(new_n817), .C2(new_n818), .ZN(new_n819));
  NAND2_X1  g618(.A1(new_n798), .A2(new_n819), .ZN(new_n820));
  NAND2_X1  g619(.A1(new_n820), .A2(new_n513), .ZN(new_n821));
  NOR2_X1   g620(.A1(new_n513), .A2(new_n793), .ZN(new_n822));
  OAI211_X1 g621(.A(new_n808), .B(new_n822), .C1(new_n817), .C2(new_n818), .ZN(new_n823));
  NAND2_X1  g622(.A1(new_n823), .A2(KEYINPUT117), .ZN(new_n824));
  OAI21_X1  g623(.A(KEYINPUT115), .B1(new_n807), .B2(KEYINPUT55), .ZN(new_n825));
  NAND3_X1  g624(.A1(new_n815), .A2(new_n809), .A3(new_n816), .ZN(new_n826));
  NAND2_X1  g625(.A1(new_n825), .A2(new_n826), .ZN(new_n827));
  INV_X1    g626(.A(KEYINPUT117), .ZN(new_n828));
  NAND4_X1  g627(.A1(new_n827), .A2(new_n828), .A3(new_n808), .A4(new_n822), .ZN(new_n829));
  NAND2_X1  g628(.A1(new_n824), .A2(new_n829), .ZN(new_n830));
  NAND2_X1  g629(.A1(new_n821), .A2(new_n830), .ZN(new_n831));
  AOI21_X1  g630(.A(new_n785), .B1(new_n831), .B2(new_n672), .ZN(new_n832));
  NOR2_X1   g631(.A1(new_n832), .A2(new_n320), .ZN(new_n833));
  NOR2_X1   g632(.A1(new_n279), .A2(new_n695), .ZN(new_n834));
  NAND3_X1  g633(.A1(new_n833), .A2(new_n834), .A3(new_n713), .ZN(new_n835));
  OAI21_X1  g634(.A(G113gat), .B1(new_n835), .B2(new_n627), .ZN(new_n836));
  AND2_X1   g635(.A1(new_n667), .A2(new_n407), .ZN(new_n837));
  NAND3_X1  g636(.A1(new_n833), .A2(new_n837), .A3(new_n713), .ZN(new_n838));
  OR2_X1    g637(.A1(new_n838), .A2(G113gat), .ZN(new_n839));
  OAI21_X1  g638(.A(new_n836), .B1(new_n839), .B2(new_n627), .ZN(G1340gat));
  OAI21_X1  g639(.A(G120gat), .B1(new_n835), .B2(new_n751), .ZN(new_n841));
  OR2_X1    g640(.A1(new_n838), .A2(G120gat), .ZN(new_n842));
  OAI21_X1  g641(.A(new_n841), .B1(new_n842), .B2(new_n751), .ZN(G1341gat));
  INV_X1    g642(.A(KEYINPUT120), .ZN(new_n844));
  OR3_X1    g643(.A1(new_n838), .A2(new_n844), .A3(new_n672), .ZN(new_n845));
  INV_X1    g644(.A(G127gat), .ZN(new_n846));
  OAI21_X1  g645(.A(new_n844), .B1(new_n838), .B2(new_n672), .ZN(new_n847));
  NAND3_X1  g646(.A1(new_n845), .A2(new_n846), .A3(new_n847), .ZN(new_n848));
  NOR3_X1   g647(.A1(new_n835), .A2(new_n846), .A3(new_n672), .ZN(new_n849));
  INV_X1    g648(.A(KEYINPUT119), .ZN(new_n850));
  OR2_X1    g649(.A1(new_n849), .A2(new_n850), .ZN(new_n851));
  NAND2_X1  g650(.A1(new_n849), .A2(new_n850), .ZN(new_n852));
  AND3_X1   g651(.A1(new_n848), .A2(new_n851), .A3(new_n852), .ZN(G1342gat));
  NAND2_X1  g652(.A1(new_n833), .A2(new_n837), .ZN(new_n854));
  NOR4_X1   g653(.A1(new_n854), .A2(G134gat), .A3(new_n380), .A4(new_n513), .ZN(new_n855));
  XNOR2_X1  g654(.A(new_n855), .B(KEYINPUT56), .ZN(new_n856));
  OAI21_X1  g655(.A(G134gat), .B1(new_n835), .B2(new_n513), .ZN(new_n857));
  NAND2_X1  g656(.A1(new_n856), .A2(new_n857), .ZN(G1343gat));
  NAND2_X1  g657(.A1(new_n650), .A2(new_n796), .ZN(new_n859));
  NAND3_X1  g658(.A1(new_n815), .A2(KEYINPUT121), .A3(new_n816), .ZN(new_n860));
  NAND2_X1  g659(.A1(new_n749), .A2(new_n750), .ZN(new_n861));
  NAND2_X1  g660(.A1(new_n860), .A2(new_n861), .ZN(new_n862));
  INV_X1    g661(.A(KEYINPUT121), .ZN(new_n863));
  AOI21_X1  g662(.A(new_n863), .B1(new_n813), .B2(new_n814), .ZN(new_n864));
  OAI21_X1  g663(.A(new_n626), .B1(new_n864), .B2(new_n816), .ZN(new_n865));
  OAI21_X1  g664(.A(new_n859), .B1(new_n862), .B2(new_n865), .ZN(new_n866));
  NAND2_X1  g665(.A1(new_n866), .A2(new_n513), .ZN(new_n867));
  AOI21_X1  g666(.A(new_n601), .B1(new_n830), .B2(new_n867), .ZN(new_n868));
  OAI21_X1  g667(.A(new_n279), .B1(new_n868), .B2(new_n785), .ZN(new_n869));
  NAND2_X1  g668(.A1(new_n869), .A2(KEYINPUT57), .ZN(new_n870));
  NOR3_X1   g669(.A1(new_n722), .A2(new_n320), .A3(new_n763), .ZN(new_n871));
  INV_X1    g670(.A(KEYINPUT57), .ZN(new_n872));
  AOI21_X1  g671(.A(new_n601), .B1(new_n821), .B2(new_n830), .ZN(new_n873));
  OAI211_X1 g672(.A(new_n872), .B(new_n279), .C1(new_n873), .C2(new_n785), .ZN(new_n874));
  NAND4_X1  g673(.A1(new_n870), .A2(new_n626), .A3(new_n871), .A4(new_n874), .ZN(new_n875));
  NAND2_X1  g674(.A1(new_n875), .A2(G141gat), .ZN(new_n876));
  AOI21_X1  g675(.A(KEYINPUT58), .B1(new_n876), .B2(KEYINPUT122), .ZN(new_n877));
  OAI21_X1  g676(.A(new_n279), .B1(new_n873), .B2(new_n785), .ZN(new_n878));
  INV_X1    g677(.A(new_n878), .ZN(new_n879));
  NAND2_X1  g678(.A1(new_n879), .A2(new_n871), .ZN(new_n880));
  INV_X1    g679(.A(new_n880), .ZN(new_n881));
  NOR2_X1   g680(.A1(new_n627), .A2(G141gat), .ZN(new_n882));
  AOI22_X1  g681(.A1(new_n881), .A2(new_n882), .B1(new_n875), .B2(G141gat), .ZN(new_n883));
  XNOR2_X1  g682(.A(new_n877), .B(new_n883), .ZN(G1344gat));
  INV_X1    g683(.A(KEYINPUT124), .ZN(new_n885));
  OAI21_X1  g684(.A(new_n861), .B1(new_n815), .B2(new_n816), .ZN(new_n886));
  AOI21_X1  g685(.A(new_n886), .B1(new_n825), .B2(new_n826), .ZN(new_n887));
  AOI22_X1  g686(.A1(new_n866), .A2(new_n513), .B1(new_n887), .B2(new_n822), .ZN(new_n888));
  OAI211_X1 g687(.A(new_n885), .B(new_n784), .C1(new_n888), .C2(new_n601), .ZN(new_n889));
  INV_X1    g688(.A(new_n889), .ZN(new_n890));
  OAI21_X1  g689(.A(KEYINPUT55), .B1(new_n807), .B2(new_n863), .ZN(new_n891));
  NAND4_X1  g690(.A1(new_n891), .A2(new_n626), .A3(new_n861), .A4(new_n860), .ZN(new_n892));
  AOI21_X1  g691(.A(new_n680), .B1(new_n892), .B2(new_n859), .ZN(new_n893));
  INV_X1    g692(.A(new_n823), .ZN(new_n894));
  OAI21_X1  g693(.A(new_n672), .B1(new_n893), .B2(new_n894), .ZN(new_n895));
  AOI21_X1  g694(.A(new_n885), .B1(new_n895), .B2(new_n784), .ZN(new_n896));
  NOR2_X1   g695(.A1(new_n890), .A2(new_n896), .ZN(new_n897));
  NOR2_X1   g696(.A1(new_n667), .A2(KEYINPUT57), .ZN(new_n898));
  AOI22_X1  g697(.A1(new_n897), .A2(new_n898), .B1(new_n878), .B2(KEYINPUT57), .ZN(new_n899));
  NAND4_X1  g698(.A1(new_n899), .A2(KEYINPUT125), .A3(new_n650), .A4(new_n871), .ZN(new_n900));
  OAI21_X1  g699(.A(KEYINPUT57), .B1(new_n832), .B2(new_n667), .ZN(new_n901));
  AOI21_X1  g700(.A(new_n601), .B1(new_n867), .B2(new_n823), .ZN(new_n902));
  OAI21_X1  g701(.A(KEYINPUT124), .B1(new_n902), .B2(new_n785), .ZN(new_n903));
  NAND3_X1  g702(.A1(new_n903), .A2(new_n898), .A3(new_n889), .ZN(new_n904));
  NAND4_X1  g703(.A1(new_n901), .A2(new_n650), .A3(new_n871), .A4(new_n904), .ZN(new_n905));
  INV_X1    g704(.A(KEYINPUT125), .ZN(new_n906));
  NAND2_X1  g705(.A1(new_n905), .A2(new_n906), .ZN(new_n907));
  NAND3_X1  g706(.A1(new_n900), .A2(new_n907), .A3(G148gat), .ZN(new_n908));
  XOR2_X1   g707(.A(KEYINPUT123), .B(KEYINPUT59), .Z(new_n909));
  NAND2_X1  g708(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  INV_X1    g709(.A(KEYINPUT59), .ZN(new_n911));
  NAND3_X1  g710(.A1(new_n870), .A2(new_n871), .A3(new_n874), .ZN(new_n912));
  OAI211_X1 g711(.A(new_n911), .B(G148gat), .C1(new_n912), .C2(new_n751), .ZN(new_n913));
  NAND2_X1  g712(.A1(new_n910), .A2(new_n913), .ZN(new_n914));
  OR3_X1    g713(.A1(new_n880), .A2(G148gat), .A3(new_n751), .ZN(new_n915));
  NAND2_X1  g714(.A1(new_n914), .A2(new_n915), .ZN(G1345gat));
  AOI21_X1  g715(.A(G155gat), .B1(new_n881), .B2(new_n601), .ZN(new_n917));
  NOR2_X1   g716(.A1(new_n912), .A2(new_n672), .ZN(new_n918));
  AOI21_X1  g717(.A(new_n917), .B1(G155gat), .B2(new_n918), .ZN(G1346gat));
  OAI21_X1  g718(.A(G162gat), .B1(new_n912), .B2(new_n513), .ZN(new_n920));
  NOR3_X1   g719(.A1(new_n380), .A2(G162gat), .A3(new_n513), .ZN(new_n921));
  NAND4_X1  g720(.A1(new_n879), .A2(new_n321), .A3(new_n409), .A4(new_n921), .ZN(new_n922));
  NAND2_X1  g721(.A1(new_n920), .A2(new_n922), .ZN(G1347gat));
  INV_X1    g722(.A(new_n832), .ZN(new_n924));
  NAND4_X1  g723(.A1(new_n924), .A2(new_n320), .A3(new_n380), .A4(new_n834), .ZN(new_n925));
  OAI21_X1  g724(.A(G169gat), .B1(new_n925), .B2(new_n627), .ZN(new_n926));
  NAND3_X1  g725(.A1(new_n924), .A2(new_n320), .A3(new_n763), .ZN(new_n927));
  INV_X1    g726(.A(new_n927), .ZN(new_n928));
  NAND2_X1  g727(.A1(new_n928), .A2(new_n837), .ZN(new_n929));
  OR2_X1    g728(.A1(new_n929), .A2(KEYINPUT126), .ZN(new_n930));
  INV_X1    g729(.A(G169gat), .ZN(new_n931));
  NAND2_X1  g730(.A1(new_n929), .A2(KEYINPUT126), .ZN(new_n932));
  NAND3_X1  g731(.A1(new_n930), .A2(new_n931), .A3(new_n932), .ZN(new_n933));
  OAI21_X1  g732(.A(new_n926), .B1(new_n933), .B2(new_n627), .ZN(G1348gat));
  INV_X1    g733(.A(G176gat), .ZN(new_n935));
  NOR3_X1   g734(.A1(new_n925), .A2(new_n935), .A3(new_n751), .ZN(new_n936));
  NAND3_X1  g735(.A1(new_n930), .A2(new_n650), .A3(new_n932), .ZN(new_n937));
  AOI21_X1  g736(.A(new_n936), .B1(new_n937), .B2(new_n935), .ZN(G1349gat));
  OAI21_X1  g737(.A(G183gat), .B1(new_n925), .B2(new_n672), .ZN(new_n939));
  NAND2_X1  g738(.A1(new_n601), .A2(new_n322), .ZN(new_n940));
  OAI21_X1  g739(.A(new_n939), .B1(new_n929), .B2(new_n940), .ZN(new_n941));
  XNOR2_X1  g740(.A(new_n941), .B(KEYINPUT60), .ZN(G1350gat));
  NAND4_X1  g741(.A1(new_n930), .A2(new_n323), .A3(new_n680), .A4(new_n932), .ZN(new_n943));
  OAI21_X1  g742(.A(G190gat), .B1(new_n925), .B2(new_n513), .ZN(new_n944));
  AND2_X1   g743(.A1(new_n944), .A2(KEYINPUT61), .ZN(new_n945));
  OR2_X1    g744(.A1(new_n944), .A2(KEYINPUT61), .ZN(new_n946));
  INV_X1    g745(.A(new_n946), .ZN(new_n947));
  OAI21_X1  g746(.A(new_n943), .B1(new_n945), .B2(new_n947), .ZN(G1351gat));
  NOR3_X1   g747(.A1(new_n927), .A2(new_n667), .A3(new_n722), .ZN(new_n949));
  NAND3_X1  g748(.A1(new_n949), .A2(new_n606), .A3(new_n626), .ZN(new_n950));
  NOR3_X1   g749(.A1(new_n722), .A2(new_n321), .A3(new_n379), .ZN(new_n951));
  AND3_X1   g750(.A1(new_n899), .A2(new_n626), .A3(new_n951), .ZN(new_n952));
  OAI21_X1  g751(.A(new_n950), .B1(new_n606), .B2(new_n952), .ZN(G1352gat));
  INV_X1    g752(.A(G204gat), .ZN(new_n954));
  NAND3_X1  g753(.A1(new_n949), .A2(new_n954), .A3(new_n650), .ZN(new_n955));
  OR2_X1    g754(.A1(new_n955), .A2(KEYINPUT62), .ZN(new_n956));
  NAND2_X1  g755(.A1(new_n955), .A2(KEYINPUT62), .ZN(new_n957));
  AND3_X1   g756(.A1(new_n899), .A2(new_n650), .A3(new_n951), .ZN(new_n958));
  OAI211_X1 g757(.A(new_n956), .B(new_n957), .C1(new_n954), .C2(new_n958), .ZN(G1353gat));
  INV_X1    g758(.A(new_n212), .ZN(new_n960));
  NAND3_X1  g759(.A1(new_n949), .A2(new_n960), .A3(new_n601), .ZN(new_n961));
  NAND3_X1  g760(.A1(new_n899), .A2(new_n601), .A3(new_n951), .ZN(new_n962));
  AND3_X1   g761(.A1(new_n962), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n963));
  AOI21_X1  g762(.A(KEYINPUT63), .B1(new_n962), .B2(G211gat), .ZN(new_n964));
  OAI21_X1  g763(.A(new_n961), .B1(new_n963), .B2(new_n964), .ZN(G1354gat));
  NOR2_X1   g764(.A1(new_n927), .A2(new_n722), .ZN(new_n966));
  INV_X1    g765(.A(G218gat), .ZN(new_n967));
  NAND4_X1  g766(.A1(new_n966), .A2(new_n967), .A3(new_n279), .A4(new_n680), .ZN(new_n968));
  NAND4_X1  g767(.A1(new_n901), .A2(new_n680), .A3(new_n904), .A4(new_n951), .ZN(new_n969));
  NAND2_X1  g768(.A1(new_n969), .A2(G218gat), .ZN(new_n970));
  NAND2_X1  g769(.A1(new_n968), .A2(new_n970), .ZN(new_n971));
  INV_X1    g770(.A(KEYINPUT127), .ZN(new_n972));
  XNOR2_X1  g771(.A(new_n971), .B(new_n972), .ZN(G1355gat));
endmodule


