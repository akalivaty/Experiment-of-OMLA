//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 1 1 0 0 0 0 0 0 0 1 0 1 0 0 1 1 1 1 0 0 1 1 0 0 1 0 0 0 1 0 1 1 0 0 1 0 0 0 0 1 0 0 0 0 1 1 0 1 0 0 1 1 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:18:14 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n701, new_n702, new_n703, new_n704, new_n705, new_n706,
    new_n708, new_n709, new_n710, new_n711, new_n712, new_n714, new_n715,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n772, new_n773,
    new_n774, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n797, new_n798, new_n799, new_n800, new_n801, new_n802, new_n803,
    new_n804, new_n805, new_n807, new_n808, new_n809, new_n811, new_n812,
    new_n813, new_n814, new_n816, new_n817, new_n818, new_n819, new_n821,
    new_n822, new_n824, new_n825, new_n826, new_n827, new_n828, new_n829,
    new_n830, new_n831, new_n832, new_n833, new_n834, new_n835, new_n836,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n845,
    new_n846, new_n847, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n891, new_n892, new_n894, new_n895, new_n897, new_n898, new_n899,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n948, new_n949, new_n950,
    new_n951, new_n953, new_n954, new_n955, new_n957, new_n958, new_n959,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n970, new_n971, new_n973, new_n974, new_n975, new_n976,
    new_n978, new_n979, new_n980, new_n982, new_n983, new_n984, new_n985,
    new_n986, new_n987, new_n988, new_n989, new_n990, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1003, new_n1004, new_n1005, new_n1006, new_n1008,
    new_n1009;
  INV_X1    g000(.A(G113gat), .ZN(new_n202));
  NAND2_X1  g001(.A1(new_n202), .A2(KEYINPUT70), .ZN(new_n203));
  INV_X1    g002(.A(KEYINPUT70), .ZN(new_n204));
  NAND2_X1  g003(.A1(new_n204), .A2(G113gat), .ZN(new_n205));
  NAND3_X1  g004(.A1(new_n203), .A2(new_n205), .A3(G120gat), .ZN(new_n206));
  INV_X1    g005(.A(KEYINPUT69), .ZN(new_n207));
  OAI21_X1  g006(.A(new_n207), .B1(new_n202), .B2(G120gat), .ZN(new_n208));
  INV_X1    g007(.A(G120gat), .ZN(new_n209));
  NAND3_X1  g008(.A1(new_n209), .A2(KEYINPUT69), .A3(G113gat), .ZN(new_n210));
  NAND3_X1  g009(.A1(new_n206), .A2(new_n208), .A3(new_n210), .ZN(new_n211));
  INV_X1    g010(.A(G134gat), .ZN(new_n212));
  NAND2_X1  g011(.A1(new_n212), .A2(G127gat), .ZN(new_n213));
  INV_X1    g012(.A(G127gat), .ZN(new_n214));
  NAND2_X1  g013(.A1(new_n214), .A2(G134gat), .ZN(new_n215));
  INV_X1    g014(.A(KEYINPUT1), .ZN(new_n216));
  AND3_X1   g015(.A1(new_n213), .A2(new_n215), .A3(new_n216), .ZN(new_n217));
  NOR2_X1   g016(.A1(new_n202), .A2(G120gat), .ZN(new_n218));
  NOR2_X1   g017(.A1(new_n209), .A2(G113gat), .ZN(new_n219));
  OAI21_X1  g018(.A(new_n216), .B1(new_n218), .B2(new_n219), .ZN(new_n220));
  NAND2_X1  g019(.A1(new_n213), .A2(new_n215), .ZN(new_n221));
  AOI22_X1  g020(.A1(new_n211), .A2(new_n217), .B1(new_n220), .B2(new_n221), .ZN(new_n222));
  NAND2_X1  g021(.A1(G169gat), .A2(G176gat), .ZN(new_n223));
  INV_X1    g022(.A(KEYINPUT26), .ZN(new_n224));
  NAND2_X1  g023(.A1(new_n223), .A2(new_n224), .ZN(new_n225));
  INV_X1    g024(.A(KEYINPUT67), .ZN(new_n226));
  INV_X1    g025(.A(G169gat), .ZN(new_n227));
  INV_X1    g026(.A(G176gat), .ZN(new_n228));
  NAND2_X1  g027(.A1(new_n227), .A2(new_n228), .ZN(new_n229));
  NAND3_X1  g028(.A1(new_n225), .A2(new_n226), .A3(new_n229), .ZN(new_n230));
  INV_X1    g029(.A(KEYINPUT68), .ZN(new_n231));
  OAI21_X1  g030(.A(new_n231), .B1(new_n229), .B2(KEYINPUT26), .ZN(new_n232));
  AOI21_X1  g031(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n233));
  NOR2_X1   g032(.A1(G169gat), .A2(G176gat), .ZN(new_n234));
  OAI21_X1  g033(.A(KEYINPUT67), .B1(new_n233), .B2(new_n234), .ZN(new_n235));
  NAND3_X1  g034(.A1(new_n234), .A2(KEYINPUT68), .A3(new_n224), .ZN(new_n236));
  NAND4_X1  g035(.A1(new_n230), .A2(new_n232), .A3(new_n235), .A4(new_n236), .ZN(new_n237));
  INV_X1    g036(.A(new_n237), .ZN(new_n238));
  NAND2_X1  g037(.A1(G183gat), .A2(G190gat), .ZN(new_n239));
  NAND2_X1  g038(.A1(KEYINPUT66), .A2(G183gat), .ZN(new_n240));
  AOI21_X1  g039(.A(G190gat), .B1(new_n240), .B2(KEYINPUT27), .ZN(new_n241));
  INV_X1    g040(.A(KEYINPUT27), .ZN(new_n242));
  NAND3_X1  g041(.A1(new_n242), .A2(KEYINPUT66), .A3(G183gat), .ZN(new_n243));
  AOI21_X1  g042(.A(KEYINPUT28), .B1(new_n241), .B2(new_n243), .ZN(new_n244));
  NAND2_X1  g043(.A1(new_n242), .A2(G183gat), .ZN(new_n245));
  INV_X1    g044(.A(G183gat), .ZN(new_n246));
  NAND2_X1  g045(.A1(new_n246), .A2(KEYINPUT27), .ZN(new_n247));
  INV_X1    g046(.A(G190gat), .ZN(new_n248));
  AND4_X1   g047(.A1(KEYINPUT28), .A2(new_n245), .A3(new_n247), .A4(new_n248), .ZN(new_n249));
  OAI21_X1  g048(.A(new_n239), .B1(new_n244), .B2(new_n249), .ZN(new_n250));
  NOR2_X1   g049(.A1(new_n238), .A2(new_n250), .ZN(new_n251));
  NAND2_X1  g050(.A1(KEYINPUT24), .A2(G183gat), .ZN(new_n252));
  OAI21_X1  g051(.A(new_n223), .B1(new_n252), .B2(G190gat), .ZN(new_n253));
  AOI21_X1  g052(.A(KEYINPUT23), .B1(new_n227), .B2(new_n228), .ZN(new_n254));
  NOR2_X1   g053(.A1(new_n253), .A2(new_n254), .ZN(new_n255));
  OR2_X1    g054(.A1(KEYINPUT24), .A2(G183gat), .ZN(new_n256));
  NAND3_X1  g055(.A1(new_n256), .A2(G190gat), .A3(new_n252), .ZN(new_n257));
  INV_X1    g056(.A(KEYINPUT65), .ZN(new_n258));
  INV_X1    g057(.A(KEYINPUT23), .ZN(new_n259));
  OAI21_X1  g058(.A(new_n258), .B1(new_n229), .B2(new_n259), .ZN(new_n260));
  NAND3_X1  g059(.A1(new_n234), .A2(KEYINPUT65), .A3(KEYINPUT23), .ZN(new_n261));
  NAND4_X1  g060(.A1(new_n255), .A2(new_n257), .A3(new_n260), .A4(new_n261), .ZN(new_n262));
  INV_X1    g061(.A(KEYINPUT25), .ZN(new_n263));
  NAND3_X1  g062(.A1(new_n248), .A2(KEYINPUT24), .A3(G183gat), .ZN(new_n264));
  OAI211_X1 g063(.A(new_n264), .B(new_n223), .C1(KEYINPUT23), .C2(new_n234), .ZN(new_n265));
  NAND2_X1  g064(.A1(new_n252), .A2(G190gat), .ZN(new_n266));
  NOR2_X1   g065(.A1(KEYINPUT24), .A2(G183gat), .ZN(new_n267));
  NOR2_X1   g066(.A1(new_n266), .A2(new_n267), .ZN(new_n268));
  NOR2_X1   g067(.A1(new_n265), .A2(new_n268), .ZN(new_n269));
  AOI21_X1  g068(.A(new_n263), .B1(new_n234), .B2(KEYINPUT23), .ZN(new_n270));
  AOI22_X1  g069(.A1(new_n262), .A2(new_n263), .B1(new_n269), .B2(new_n270), .ZN(new_n271));
  OAI21_X1  g070(.A(new_n222), .B1(new_n251), .B2(new_n271), .ZN(new_n272));
  NAND2_X1  g071(.A1(new_n262), .A2(new_n263), .ZN(new_n273));
  NAND2_X1  g072(.A1(new_n269), .A2(new_n270), .ZN(new_n274));
  NAND2_X1  g073(.A1(new_n273), .A2(new_n274), .ZN(new_n275));
  AND3_X1   g074(.A1(new_n203), .A2(new_n205), .A3(G120gat), .ZN(new_n276));
  NAND2_X1  g075(.A1(new_n208), .A2(new_n210), .ZN(new_n277));
  OAI21_X1  g076(.A(new_n217), .B1(new_n276), .B2(new_n277), .ZN(new_n278));
  NAND2_X1  g077(.A1(new_n220), .A2(new_n221), .ZN(new_n279));
  NAND2_X1  g078(.A1(new_n278), .A2(new_n279), .ZN(new_n280));
  OAI211_X1 g079(.A(new_n237), .B(new_n239), .C1(new_n244), .C2(new_n249), .ZN(new_n281));
  NAND3_X1  g080(.A1(new_n275), .A2(new_n280), .A3(new_n281), .ZN(new_n282));
  NAND2_X1  g081(.A1(G227gat), .A2(G233gat), .ZN(new_n283));
  XNOR2_X1  g082(.A(new_n283), .B(KEYINPUT64), .ZN(new_n284));
  NAND3_X1  g083(.A1(new_n272), .A2(new_n282), .A3(new_n284), .ZN(new_n285));
  NAND2_X1  g084(.A1(new_n285), .A2(KEYINPUT32), .ZN(new_n286));
  INV_X1    g085(.A(KEYINPUT33), .ZN(new_n287));
  NAND2_X1  g086(.A1(new_n285), .A2(new_n287), .ZN(new_n288));
  XOR2_X1   g087(.A(G15gat), .B(G43gat), .Z(new_n289));
  XNOR2_X1  g088(.A(G71gat), .B(G99gat), .ZN(new_n290));
  XNOR2_X1  g089(.A(new_n289), .B(new_n290), .ZN(new_n291));
  NAND3_X1  g090(.A1(new_n286), .A2(new_n288), .A3(new_n291), .ZN(new_n292));
  INV_X1    g091(.A(new_n291), .ZN(new_n293));
  OAI211_X1 g092(.A(new_n285), .B(KEYINPUT32), .C1(new_n287), .C2(new_n293), .ZN(new_n294));
  NAND2_X1  g093(.A1(new_n292), .A2(new_n294), .ZN(new_n295));
  NOR3_X1   g094(.A1(new_n251), .A2(new_n271), .A3(new_n222), .ZN(new_n296));
  AOI21_X1  g095(.A(new_n280), .B1(new_n275), .B2(new_n281), .ZN(new_n297));
  OAI21_X1  g096(.A(new_n283), .B1(new_n296), .B2(new_n297), .ZN(new_n298));
  NAND2_X1  g097(.A1(new_n298), .A2(KEYINPUT34), .ZN(new_n299));
  NOR2_X1   g098(.A1(new_n284), .A2(KEYINPUT34), .ZN(new_n300));
  OAI21_X1  g099(.A(new_n300), .B1(new_n296), .B2(new_n297), .ZN(new_n301));
  INV_X1    g100(.A(KEYINPUT71), .ZN(new_n302));
  NAND2_X1  g101(.A1(new_n301), .A2(new_n302), .ZN(new_n303));
  OAI211_X1 g102(.A(KEYINPUT71), .B(new_n300), .C1(new_n296), .C2(new_n297), .ZN(new_n304));
  NAND3_X1  g103(.A1(new_n299), .A2(new_n303), .A3(new_n304), .ZN(new_n305));
  NOR2_X1   g104(.A1(new_n295), .A2(new_n305), .ZN(new_n306));
  AOI22_X1  g105(.A1(new_n302), .A2(new_n301), .B1(new_n298), .B2(KEYINPUT34), .ZN(new_n307));
  AOI22_X1  g106(.A1(new_n304), .A2(new_n307), .B1(new_n292), .B2(new_n294), .ZN(new_n308));
  NOR2_X1   g107(.A1(new_n306), .A2(new_n308), .ZN(new_n309));
  INV_X1    g108(.A(KEYINPUT35), .ZN(new_n310));
  XNOR2_X1  g109(.A(G78gat), .B(G106gat), .ZN(new_n311));
  XNOR2_X1  g110(.A(KEYINPUT31), .B(G50gat), .ZN(new_n312));
  XNOR2_X1  g111(.A(new_n311), .B(new_n312), .ZN(new_n313));
  INV_X1    g112(.A(G22gat), .ZN(new_n314));
  NAND2_X1  g113(.A1(G228gat), .A2(G233gat), .ZN(new_n315));
  NAND2_X1  g114(.A1(G155gat), .A2(G162gat), .ZN(new_n316));
  NAND2_X1  g115(.A1(new_n316), .A2(KEYINPUT2), .ZN(new_n317));
  INV_X1    g116(.A(G141gat), .ZN(new_n318));
  INV_X1    g117(.A(G148gat), .ZN(new_n319));
  NAND2_X1  g118(.A1(new_n318), .A2(new_n319), .ZN(new_n320));
  NAND2_X1  g119(.A1(G141gat), .A2(G148gat), .ZN(new_n321));
  NAND3_X1  g120(.A1(new_n317), .A2(new_n320), .A3(new_n321), .ZN(new_n322));
  NAND2_X1  g121(.A1(new_n316), .A2(KEYINPUT77), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n322), .A2(new_n323), .ZN(new_n324));
  XNOR2_X1  g123(.A(G155gat), .B(G162gat), .ZN(new_n325));
  INV_X1    g124(.A(new_n325), .ZN(new_n326));
  NAND2_X1  g125(.A1(new_n324), .A2(new_n326), .ZN(new_n327));
  NAND3_X1  g126(.A1(new_n322), .A2(new_n325), .A3(new_n323), .ZN(new_n328));
  NAND2_X1  g127(.A1(new_n327), .A2(new_n328), .ZN(new_n329));
  INV_X1    g128(.A(KEYINPUT29), .ZN(new_n330));
  INV_X1    g129(.A(G204gat), .ZN(new_n331));
  AND2_X1   g130(.A1(KEYINPUT72), .A2(G197gat), .ZN(new_n332));
  NOR2_X1   g131(.A1(KEYINPUT72), .A2(G197gat), .ZN(new_n333));
  OAI21_X1  g132(.A(new_n331), .B1(new_n332), .B2(new_n333), .ZN(new_n334));
  INV_X1    g133(.A(KEYINPUT72), .ZN(new_n335));
  INV_X1    g134(.A(G197gat), .ZN(new_n336));
  NAND2_X1  g135(.A1(new_n335), .A2(new_n336), .ZN(new_n337));
  NAND2_X1  g136(.A1(KEYINPUT72), .A2(G197gat), .ZN(new_n338));
  NAND3_X1  g137(.A1(new_n337), .A2(G204gat), .A3(new_n338), .ZN(new_n339));
  NAND2_X1  g138(.A1(new_n334), .A2(new_n339), .ZN(new_n340));
  AND2_X1   g139(.A1(G211gat), .A2(G218gat), .ZN(new_n341));
  NOR2_X1   g140(.A1(G211gat), .A2(G218gat), .ZN(new_n342));
  NOR2_X1   g141(.A1(new_n341), .A2(new_n342), .ZN(new_n343));
  INV_X1    g142(.A(new_n343), .ZN(new_n344));
  OR2_X1    g143(.A1(new_n341), .A2(KEYINPUT22), .ZN(new_n345));
  AND3_X1   g144(.A1(new_n340), .A2(new_n344), .A3(new_n345), .ZN(new_n346));
  AOI21_X1  g145(.A(new_n344), .B1(new_n340), .B2(new_n345), .ZN(new_n347));
  OAI21_X1  g146(.A(new_n330), .B1(new_n346), .B2(new_n347), .ZN(new_n348));
  INV_X1    g147(.A(KEYINPUT3), .ZN(new_n349));
  AOI21_X1  g148(.A(new_n329), .B1(new_n348), .B2(new_n349), .ZN(new_n350));
  NOR3_X1   g149(.A1(new_n332), .A2(new_n333), .A3(new_n331), .ZN(new_n351));
  AOI21_X1  g150(.A(G204gat), .B1(new_n337), .B2(new_n338), .ZN(new_n352));
  OAI21_X1  g151(.A(new_n345), .B1(new_n351), .B2(new_n352), .ZN(new_n353));
  NAND2_X1  g152(.A1(new_n353), .A2(new_n343), .ZN(new_n354));
  NAND3_X1  g153(.A1(new_n340), .A2(new_n344), .A3(new_n345), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n354), .A2(new_n355), .ZN(new_n356));
  AND3_X1   g155(.A1(new_n322), .A2(new_n325), .A3(new_n323), .ZN(new_n357));
  AOI21_X1  g156(.A(new_n325), .B1(new_n322), .B2(new_n323), .ZN(new_n358));
  OAI21_X1  g157(.A(new_n349), .B1(new_n357), .B2(new_n358), .ZN(new_n359));
  AOI21_X1  g158(.A(new_n356), .B1(new_n330), .B2(new_n359), .ZN(new_n360));
  OAI21_X1  g159(.A(new_n315), .B1(new_n350), .B2(new_n360), .ZN(new_n361));
  NOR2_X1   g160(.A1(new_n357), .A2(new_n358), .ZN(new_n362));
  AOI21_X1  g161(.A(KEYINPUT29), .B1(new_n354), .B2(new_n355), .ZN(new_n363));
  OAI21_X1  g162(.A(new_n362), .B1(new_n363), .B2(KEYINPUT3), .ZN(new_n364));
  INV_X1    g163(.A(new_n315), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n359), .A2(new_n330), .ZN(new_n366));
  NOR2_X1   g165(.A1(new_n346), .A2(new_n347), .ZN(new_n367));
  NAND2_X1  g166(.A1(new_n366), .A2(new_n367), .ZN(new_n368));
  NAND3_X1  g167(.A1(new_n364), .A2(new_n365), .A3(new_n368), .ZN(new_n369));
  AOI21_X1  g168(.A(new_n314), .B1(new_n361), .B2(new_n369), .ZN(new_n370));
  INV_X1    g169(.A(KEYINPUT81), .ZN(new_n371));
  OAI21_X1  g170(.A(new_n313), .B1(new_n370), .B2(new_n371), .ZN(new_n372));
  NOR3_X1   g171(.A1(new_n350), .A2(new_n360), .A3(new_n315), .ZN(new_n373));
  AOI21_X1  g172(.A(new_n365), .B1(new_n364), .B2(new_n368), .ZN(new_n374));
  OAI21_X1  g173(.A(G22gat), .B1(new_n373), .B2(new_n374), .ZN(new_n375));
  NAND3_X1  g174(.A1(new_n361), .A2(new_n314), .A3(new_n369), .ZN(new_n376));
  NAND2_X1  g175(.A1(new_n375), .A2(new_n376), .ZN(new_n377));
  NAND2_X1  g176(.A1(new_n372), .A2(new_n377), .ZN(new_n378));
  NAND4_X1  g177(.A1(new_n375), .A2(new_n371), .A3(new_n376), .A4(new_n313), .ZN(new_n379));
  NAND2_X1  g178(.A1(new_n378), .A2(new_n379), .ZN(new_n380));
  NAND3_X1  g179(.A1(new_n309), .A2(new_n310), .A3(new_n380), .ZN(new_n381));
  OAI211_X1 g180(.A(new_n279), .B(new_n278), .C1(new_n357), .C2(new_n358), .ZN(new_n382));
  INV_X1    g181(.A(KEYINPUT4), .ZN(new_n383));
  NAND2_X1  g182(.A1(new_n382), .A2(new_n383), .ZN(new_n384));
  INV_X1    g183(.A(KEYINPUT5), .ZN(new_n385));
  XNOR2_X1  g184(.A(KEYINPUT78), .B(KEYINPUT4), .ZN(new_n386));
  INV_X1    g185(.A(new_n386), .ZN(new_n387));
  NAND3_X1  g186(.A1(new_n329), .A2(new_n222), .A3(new_n387), .ZN(new_n388));
  NAND3_X1  g187(.A1(new_n384), .A2(new_n385), .A3(new_n388), .ZN(new_n389));
  NAND3_X1  g188(.A1(new_n327), .A2(KEYINPUT3), .A3(new_n328), .ZN(new_n390));
  NAND3_X1  g189(.A1(new_n359), .A2(new_n390), .A3(new_n280), .ZN(new_n391));
  NAND2_X1  g190(.A1(G225gat), .A2(G233gat), .ZN(new_n392));
  NAND2_X1  g191(.A1(new_n391), .A2(new_n392), .ZN(new_n393));
  NOR2_X1   g192(.A1(new_n389), .A2(new_n393), .ZN(new_n394));
  INV_X1    g193(.A(new_n392), .ZN(new_n395));
  AOI21_X1  g194(.A(new_n222), .B1(new_n362), .B2(KEYINPUT3), .ZN(new_n396));
  AOI21_X1  g195(.A(new_n395), .B1(new_n396), .B2(new_n359), .ZN(new_n397));
  NAND3_X1  g196(.A1(new_n329), .A2(new_n383), .A3(new_n222), .ZN(new_n398));
  AOI21_X1  g197(.A(new_n386), .B1(new_n329), .B2(new_n222), .ZN(new_n399));
  INV_X1    g198(.A(KEYINPUT79), .ZN(new_n400));
  OAI21_X1  g199(.A(new_n398), .B1(new_n399), .B2(new_n400), .ZN(new_n401));
  OAI21_X1  g200(.A(new_n387), .B1(new_n362), .B2(new_n280), .ZN(new_n402));
  NOR2_X1   g201(.A1(new_n402), .A2(KEYINPUT79), .ZN(new_n403));
  OAI21_X1  g202(.A(new_n397), .B1(new_n401), .B2(new_n403), .ZN(new_n404));
  NAND3_X1  g203(.A1(new_n213), .A2(new_n215), .A3(new_n216), .ZN(new_n405));
  INV_X1    g204(.A(new_n277), .ZN(new_n406));
  AOI21_X1  g205(.A(new_n405), .B1(new_n406), .B2(new_n206), .ZN(new_n407));
  AND2_X1   g206(.A1(new_n220), .A2(new_n221), .ZN(new_n408));
  OAI211_X1 g207(.A(new_n327), .B(new_n328), .C1(new_n407), .C2(new_n408), .ZN(new_n409));
  NAND2_X1  g208(.A1(new_n409), .A2(new_n382), .ZN(new_n410));
  AOI21_X1  g209(.A(new_n385), .B1(new_n410), .B2(new_n395), .ZN(new_n411));
  AOI21_X1  g210(.A(new_n394), .B1(new_n404), .B2(new_n411), .ZN(new_n412));
  INV_X1    g211(.A(KEYINPUT6), .ZN(new_n413));
  XNOR2_X1  g212(.A(G1gat), .B(G29gat), .ZN(new_n414));
  XNOR2_X1  g213(.A(new_n414), .B(KEYINPUT0), .ZN(new_n415));
  XNOR2_X1  g214(.A(G57gat), .B(G85gat), .ZN(new_n416));
  XNOR2_X1  g215(.A(new_n415), .B(new_n416), .ZN(new_n417));
  INV_X1    g216(.A(new_n417), .ZN(new_n418));
  NOR3_X1   g217(.A1(new_n412), .A2(new_n413), .A3(new_n418), .ZN(new_n419));
  INV_X1    g218(.A(KEYINPUT85), .ZN(new_n420));
  INV_X1    g219(.A(new_n394), .ZN(new_n421));
  INV_X1    g220(.A(new_n382), .ZN(new_n422));
  AOI22_X1  g221(.A1(new_n402), .A2(KEYINPUT79), .B1(new_n422), .B2(new_n383), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n399), .A2(new_n400), .ZN(new_n424));
  AOI21_X1  g223(.A(new_n393), .B1(new_n423), .B2(new_n424), .ZN(new_n425));
  NAND2_X1  g224(.A1(new_n410), .A2(new_n395), .ZN(new_n426));
  NAND2_X1  g225(.A1(new_n426), .A2(KEYINPUT5), .ZN(new_n427));
  OAI21_X1  g226(.A(new_n421), .B1(new_n425), .B2(new_n427), .ZN(new_n428));
  AOI21_X1  g227(.A(new_n420), .B1(new_n428), .B2(new_n417), .ZN(new_n429));
  NOR3_X1   g228(.A1(new_n412), .A2(KEYINPUT85), .A3(new_n418), .ZN(new_n430));
  NOR2_X1   g229(.A1(new_n429), .A2(new_n430), .ZN(new_n431));
  OAI211_X1 g230(.A(new_n418), .B(new_n421), .C1(new_n425), .C2(new_n427), .ZN(new_n432));
  INV_X1    g231(.A(KEYINPUT80), .ZN(new_n433));
  NAND2_X1  g232(.A1(new_n432), .A2(new_n433), .ZN(new_n434));
  NAND3_X1  g233(.A1(new_n412), .A2(KEYINPUT80), .A3(new_n418), .ZN(new_n435));
  AOI21_X1  g234(.A(KEYINPUT6), .B1(new_n434), .B2(new_n435), .ZN(new_n436));
  AOI21_X1  g235(.A(new_n419), .B1(new_n431), .B2(new_n436), .ZN(new_n437));
  NAND2_X1  g236(.A1(G226gat), .A2(G233gat), .ZN(new_n438));
  OAI21_X1  g237(.A(KEYINPUT74), .B1(new_n251), .B2(new_n271), .ZN(new_n439));
  INV_X1    g238(.A(KEYINPUT74), .ZN(new_n440));
  NAND3_X1  g239(.A1(new_n275), .A2(new_n440), .A3(new_n281), .ZN(new_n441));
  AOI21_X1  g240(.A(new_n438), .B1(new_n439), .B2(new_n441), .ZN(new_n442));
  XOR2_X1   g241(.A(new_n438), .B(KEYINPUT73), .Z(new_n443));
  NAND2_X1  g242(.A1(new_n275), .A2(new_n281), .ZN(new_n444));
  AOI21_X1  g243(.A(new_n443), .B1(new_n444), .B2(new_n330), .ZN(new_n445));
  OAI21_X1  g244(.A(new_n367), .B1(new_n442), .B2(new_n445), .ZN(new_n446));
  AOI21_X1  g245(.A(new_n367), .B1(new_n444), .B2(new_n443), .ZN(new_n447));
  AOI21_X1  g246(.A(KEYINPUT29), .B1(new_n439), .B2(new_n441), .ZN(new_n448));
  INV_X1    g247(.A(new_n438), .ZN(new_n449));
  OAI21_X1  g248(.A(new_n447), .B1(new_n448), .B2(new_n449), .ZN(new_n450));
  XNOR2_X1  g249(.A(G8gat), .B(G36gat), .ZN(new_n451));
  XNOR2_X1  g250(.A(G64gat), .B(G92gat), .ZN(new_n452));
  XOR2_X1   g251(.A(new_n451), .B(new_n452), .Z(new_n453));
  AND4_X1   g252(.A1(KEYINPUT30), .A2(new_n446), .A3(new_n450), .A4(new_n453), .ZN(new_n454));
  AOI21_X1  g253(.A(new_n453), .B1(new_n446), .B2(new_n450), .ZN(new_n455));
  NOR2_X1   g254(.A1(new_n454), .A2(new_n455), .ZN(new_n456));
  NAND3_X1  g255(.A1(new_n446), .A2(new_n450), .A3(new_n453), .ZN(new_n457));
  INV_X1    g256(.A(KEYINPUT30), .ZN(new_n458));
  AND3_X1   g257(.A1(new_n457), .A2(KEYINPUT76), .A3(new_n458), .ZN(new_n459));
  AOI21_X1  g258(.A(KEYINPUT76), .B1(new_n457), .B2(new_n458), .ZN(new_n460));
  OAI21_X1  g259(.A(new_n456), .B1(new_n459), .B2(new_n460), .ZN(new_n461));
  NOR3_X1   g260(.A1(new_n381), .A2(new_n437), .A3(new_n461), .ZN(new_n462));
  OAI21_X1  g261(.A(KEYINPUT75), .B1(new_n454), .B2(new_n455), .ZN(new_n463));
  NAND2_X1  g262(.A1(new_n446), .A2(new_n450), .ZN(new_n464));
  INV_X1    g263(.A(new_n453), .ZN(new_n465));
  NAND2_X1  g264(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  INV_X1    g265(.A(KEYINPUT75), .ZN(new_n467));
  NAND4_X1  g266(.A1(new_n446), .A2(new_n450), .A3(KEYINPUT30), .A4(new_n453), .ZN(new_n468));
  NAND3_X1  g267(.A1(new_n466), .A2(new_n467), .A3(new_n468), .ZN(new_n469));
  NAND2_X1  g268(.A1(new_n463), .A2(new_n469), .ZN(new_n470));
  AOI21_X1  g269(.A(KEYINPUT6), .B1(new_n428), .B2(new_n417), .ZN(new_n471));
  NOR2_X1   g270(.A1(new_n432), .A2(new_n433), .ZN(new_n472));
  AOI21_X1  g271(.A(KEYINPUT80), .B1(new_n412), .B2(new_n418), .ZN(new_n473));
  OAI21_X1  g272(.A(new_n471), .B1(new_n472), .B2(new_n473), .ZN(new_n474));
  INV_X1    g273(.A(new_n419), .ZN(new_n475));
  NAND2_X1  g274(.A1(new_n457), .A2(new_n458), .ZN(new_n476));
  INV_X1    g275(.A(KEYINPUT76), .ZN(new_n477));
  NAND2_X1  g276(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  NAND3_X1  g277(.A1(new_n457), .A2(KEYINPUT76), .A3(new_n458), .ZN(new_n479));
  AOI22_X1  g278(.A1(new_n474), .A2(new_n475), .B1(new_n478), .B2(new_n479), .ZN(new_n480));
  INV_X1    g279(.A(KEYINPUT86), .ZN(new_n481));
  AND3_X1   g280(.A1(new_n309), .A2(new_n481), .A3(new_n380), .ZN(new_n482));
  AOI21_X1  g281(.A(new_n481), .B1(new_n309), .B2(new_n380), .ZN(new_n483));
  OAI211_X1 g282(.A(new_n470), .B(new_n480), .C1(new_n482), .C2(new_n483), .ZN(new_n484));
  AOI21_X1  g283(.A(new_n462), .B1(new_n484), .B2(KEYINPUT35), .ZN(new_n485));
  AND2_X1   g284(.A1(new_n378), .A2(new_n379), .ZN(new_n486));
  OAI21_X1  g285(.A(new_n413), .B1(new_n412), .B2(new_n418), .ZN(new_n487));
  AOI21_X1  g286(.A(new_n487), .B1(new_n434), .B2(new_n435), .ZN(new_n488));
  OAI22_X1  g287(.A1(new_n488), .A2(new_n419), .B1(new_n460), .B2(new_n459), .ZN(new_n489));
  NOR3_X1   g288(.A1(new_n454), .A2(KEYINPUT75), .A3(new_n455), .ZN(new_n490));
  AOI21_X1  g289(.A(new_n467), .B1(new_n466), .B2(new_n468), .ZN(new_n491));
  NOR2_X1   g290(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  OAI21_X1  g291(.A(new_n486), .B1(new_n489), .B2(new_n492), .ZN(new_n493));
  XNOR2_X1  g292(.A(new_n309), .B(KEYINPUT36), .ZN(new_n494));
  NAND2_X1  g293(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  NAND3_X1  g294(.A1(new_n391), .A2(new_n384), .A3(new_n388), .ZN(new_n496));
  NAND2_X1  g295(.A1(new_n496), .A2(new_n395), .ZN(new_n497));
  NAND2_X1  g296(.A1(new_n497), .A2(KEYINPUT83), .ZN(new_n498));
  INV_X1    g297(.A(KEYINPUT83), .ZN(new_n499));
  NAND3_X1  g298(.A1(new_n496), .A2(new_n499), .A3(new_n395), .ZN(new_n500));
  NAND2_X1  g299(.A1(new_n498), .A2(new_n500), .ZN(new_n501));
  OAI21_X1  g300(.A(KEYINPUT39), .B1(new_n410), .B2(new_n395), .ZN(new_n502));
  OR2_X1    g301(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  INV_X1    g302(.A(KEYINPUT39), .ZN(new_n504));
  NAND2_X1  g303(.A1(new_n501), .A2(new_n504), .ZN(new_n505));
  NAND4_X1  g304(.A1(new_n503), .A2(new_n505), .A3(KEYINPUT40), .A4(new_n418), .ZN(new_n506));
  AND2_X1   g305(.A1(new_n506), .A2(new_n431), .ZN(new_n507));
  NAND3_X1  g306(.A1(new_n503), .A2(new_n418), .A3(new_n505), .ZN(new_n508));
  INV_X1    g307(.A(KEYINPUT84), .ZN(new_n509));
  INV_X1    g308(.A(KEYINPUT40), .ZN(new_n510));
  AND3_X1   g309(.A1(new_n508), .A2(new_n509), .A3(new_n510), .ZN(new_n511));
  AOI21_X1  g310(.A(new_n509), .B1(new_n508), .B2(new_n510), .ZN(new_n512));
  OAI211_X1 g311(.A(new_n507), .B(new_n461), .C1(new_n511), .C2(new_n512), .ZN(new_n513));
  OAI21_X1  g312(.A(new_n465), .B1(new_n464), .B2(KEYINPUT37), .ZN(new_n514));
  AOI21_X1  g313(.A(new_n356), .B1(new_n444), .B2(new_n443), .ZN(new_n515));
  OAI21_X1  g314(.A(new_n515), .B1(new_n448), .B2(new_n449), .ZN(new_n516));
  OAI21_X1  g315(.A(new_n356), .B1(new_n442), .B2(new_n445), .ZN(new_n517));
  NAND3_X1  g316(.A1(new_n516), .A2(new_n517), .A3(KEYINPUT37), .ZN(new_n518));
  INV_X1    g317(.A(KEYINPUT38), .ZN(new_n519));
  NAND2_X1  g318(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  OAI21_X1  g319(.A(new_n457), .B1(new_n514), .B2(new_n520), .ZN(new_n521));
  NAND2_X1  g320(.A1(new_n464), .A2(KEYINPUT37), .ZN(new_n522));
  AND2_X1   g321(.A1(new_n465), .A2(KEYINPUT37), .ZN(new_n523));
  OAI21_X1  g322(.A(new_n522), .B1(new_n455), .B2(new_n523), .ZN(new_n524));
  AOI21_X1  g323(.A(new_n521), .B1(KEYINPUT38), .B2(new_n524), .ZN(new_n525));
  AOI21_X1  g324(.A(new_n486), .B1(new_n525), .B2(new_n437), .ZN(new_n526));
  AOI22_X1  g325(.A1(new_n495), .A2(KEYINPUT82), .B1(new_n513), .B2(new_n526), .ZN(new_n527));
  INV_X1    g326(.A(KEYINPUT82), .ZN(new_n528));
  NAND3_X1  g327(.A1(new_n493), .A2(new_n528), .A3(new_n494), .ZN(new_n529));
  AOI21_X1  g328(.A(new_n485), .B1(new_n527), .B2(new_n529), .ZN(new_n530));
  XNOR2_X1  g329(.A(G15gat), .B(G22gat), .ZN(new_n531));
  INV_X1    g330(.A(KEYINPUT16), .ZN(new_n532));
  OAI21_X1  g331(.A(new_n531), .B1(new_n532), .B2(G1gat), .ZN(new_n533));
  OAI21_X1  g332(.A(new_n533), .B1(G1gat), .B2(new_n531), .ZN(new_n534));
  INV_X1    g333(.A(G8gat), .ZN(new_n535));
  XNOR2_X1  g334(.A(new_n534), .B(new_n535), .ZN(new_n536));
  INV_X1    g335(.A(new_n536), .ZN(new_n537));
  INV_X1    g336(.A(G29gat), .ZN(new_n538));
  INV_X1    g337(.A(G36gat), .ZN(new_n539));
  NAND3_X1  g338(.A1(new_n538), .A2(new_n539), .A3(KEYINPUT14), .ZN(new_n540));
  INV_X1    g339(.A(KEYINPUT14), .ZN(new_n541));
  OAI21_X1  g340(.A(new_n541), .B1(G29gat), .B2(G36gat), .ZN(new_n542));
  NAND2_X1  g341(.A1(new_n540), .A2(new_n542), .ZN(new_n543));
  INV_X1    g342(.A(KEYINPUT89), .ZN(new_n544));
  XNOR2_X1  g343(.A(new_n543), .B(new_n544), .ZN(new_n545));
  XNOR2_X1  g344(.A(KEYINPUT90), .B(G36gat), .ZN(new_n546));
  INV_X1    g345(.A(KEYINPUT91), .ZN(new_n547));
  NAND3_X1  g346(.A1(new_n546), .A2(new_n547), .A3(G29gat), .ZN(new_n548));
  INV_X1    g347(.A(new_n546), .ZN(new_n549));
  OAI21_X1  g348(.A(KEYINPUT91), .B1(new_n549), .B2(new_n538), .ZN(new_n550));
  NAND3_X1  g349(.A1(new_n545), .A2(new_n548), .A3(new_n550), .ZN(new_n551));
  XNOR2_X1  g350(.A(G43gat), .B(G50gat), .ZN(new_n552));
  NAND2_X1  g351(.A1(new_n552), .A2(KEYINPUT15), .ZN(new_n553));
  INV_X1    g352(.A(new_n553), .ZN(new_n554));
  AND2_X1   g353(.A1(new_n550), .A2(new_n548), .ZN(new_n555));
  NOR2_X1   g354(.A1(new_n552), .A2(KEYINPUT15), .ZN(new_n556));
  NOR3_X1   g355(.A1(new_n554), .A2(new_n543), .A3(new_n556), .ZN(new_n557));
  AOI22_X1  g356(.A1(new_n551), .A2(new_n554), .B1(new_n555), .B2(new_n557), .ZN(new_n558));
  AOI21_X1  g357(.A(new_n537), .B1(new_n558), .B2(KEYINPUT17), .ZN(new_n559));
  NAND2_X1  g358(.A1(new_n551), .A2(new_n554), .ZN(new_n560));
  NAND2_X1  g359(.A1(new_n555), .A2(new_n557), .ZN(new_n561));
  NAND2_X1  g360(.A1(new_n560), .A2(new_n561), .ZN(new_n562));
  INV_X1    g361(.A(KEYINPUT17), .ZN(new_n563));
  AOI21_X1  g362(.A(KEYINPUT92), .B1(new_n562), .B2(new_n563), .ZN(new_n564));
  INV_X1    g363(.A(KEYINPUT92), .ZN(new_n565));
  NOR3_X1   g364(.A1(new_n558), .A2(new_n565), .A3(KEYINPUT17), .ZN(new_n566));
  OAI21_X1  g365(.A(new_n559), .B1(new_n564), .B2(new_n566), .ZN(new_n567));
  NAND2_X1  g366(.A1(G229gat), .A2(G233gat), .ZN(new_n568));
  INV_X1    g367(.A(KEYINPUT93), .ZN(new_n569));
  NAND3_X1  g368(.A1(new_n562), .A2(new_n569), .A3(new_n537), .ZN(new_n570));
  OAI21_X1  g369(.A(KEYINPUT93), .B1(new_n558), .B2(new_n536), .ZN(new_n571));
  NAND2_X1  g370(.A1(new_n570), .A2(new_n571), .ZN(new_n572));
  NAND3_X1  g371(.A1(new_n567), .A2(new_n568), .A3(new_n572), .ZN(new_n573));
  INV_X1    g372(.A(KEYINPUT18), .ZN(new_n574));
  NAND2_X1  g373(.A1(new_n573), .A2(new_n574), .ZN(new_n575));
  NAND4_X1  g374(.A1(new_n567), .A2(KEYINPUT18), .A3(new_n568), .A4(new_n572), .ZN(new_n576));
  XOR2_X1   g375(.A(new_n568), .B(KEYINPUT13), .Z(new_n577));
  INV_X1    g376(.A(new_n577), .ZN(new_n578));
  NAND2_X1  g377(.A1(new_n558), .A2(new_n536), .ZN(new_n579));
  AOI21_X1  g378(.A(new_n578), .B1(new_n572), .B2(new_n579), .ZN(new_n580));
  INV_X1    g379(.A(new_n580), .ZN(new_n581));
  NAND3_X1  g380(.A1(new_n575), .A2(new_n576), .A3(new_n581), .ZN(new_n582));
  XNOR2_X1  g381(.A(G113gat), .B(G141gat), .ZN(new_n583));
  XNOR2_X1  g382(.A(KEYINPUT87), .B(G197gat), .ZN(new_n584));
  XNOR2_X1  g383(.A(new_n583), .B(new_n584), .ZN(new_n585));
  XOR2_X1   g384(.A(KEYINPUT11), .B(G169gat), .Z(new_n586));
  XNOR2_X1  g385(.A(new_n585), .B(new_n586), .ZN(new_n587));
  XOR2_X1   g386(.A(KEYINPUT88), .B(KEYINPUT12), .Z(new_n588));
  XNOR2_X1  g387(.A(new_n587), .B(new_n588), .ZN(new_n589));
  NAND2_X1  g388(.A1(new_n582), .A2(new_n589), .ZN(new_n590));
  AOI21_X1  g389(.A(new_n580), .B1(new_n573), .B2(new_n574), .ZN(new_n591));
  INV_X1    g390(.A(new_n589), .ZN(new_n592));
  NAND3_X1  g391(.A1(new_n591), .A2(new_n592), .A3(new_n576), .ZN(new_n593));
  NAND2_X1  g392(.A1(new_n590), .A2(new_n593), .ZN(new_n594));
  INV_X1    g393(.A(new_n594), .ZN(new_n595));
  NOR2_X1   g394(.A1(new_n530), .A2(new_n595), .ZN(new_n596));
  NAND2_X1  g395(.A1(G85gat), .A2(G92gat), .ZN(new_n597));
  XNOR2_X1  g396(.A(new_n597), .B(KEYINPUT7), .ZN(new_n598));
  XOR2_X1   g397(.A(G99gat), .B(G106gat), .Z(new_n599));
  INV_X1    g398(.A(new_n599), .ZN(new_n600));
  NAND2_X1  g399(.A1(G99gat), .A2(G106gat), .ZN(new_n601));
  INV_X1    g400(.A(G85gat), .ZN(new_n602));
  INV_X1    g401(.A(G92gat), .ZN(new_n603));
  AOI22_X1  g402(.A1(KEYINPUT8), .A2(new_n601), .B1(new_n602), .B2(new_n603), .ZN(new_n604));
  AND3_X1   g403(.A1(new_n598), .A2(new_n600), .A3(new_n604), .ZN(new_n605));
  AOI21_X1  g404(.A(new_n600), .B1(new_n598), .B2(new_n604), .ZN(new_n606));
  NOR2_X1   g405(.A1(new_n605), .A2(new_n606), .ZN(new_n607));
  AND2_X1   g406(.A1(G232gat), .A2(G233gat), .ZN(new_n608));
  AOI22_X1  g407(.A1(new_n562), .A2(new_n607), .B1(KEYINPUT41), .B2(new_n608), .ZN(new_n609));
  NAND3_X1  g408(.A1(new_n562), .A2(KEYINPUT92), .A3(new_n563), .ZN(new_n610));
  OAI21_X1  g409(.A(new_n565), .B1(new_n558), .B2(KEYINPUT17), .ZN(new_n611));
  NAND2_X1  g410(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  AOI21_X1  g411(.A(new_n607), .B1(new_n558), .B2(KEYINPUT17), .ZN(new_n613));
  NAND3_X1  g412(.A1(new_n612), .A2(KEYINPUT99), .A3(new_n613), .ZN(new_n614));
  INV_X1    g413(.A(new_n614), .ZN(new_n615));
  AOI21_X1  g414(.A(KEYINPUT99), .B1(new_n612), .B2(new_n613), .ZN(new_n616));
  OAI21_X1  g415(.A(new_n609), .B1(new_n615), .B2(new_n616), .ZN(new_n617));
  XOR2_X1   g416(.A(G190gat), .B(G218gat), .Z(new_n618));
  NAND2_X1  g417(.A1(new_n617), .A2(new_n618), .ZN(new_n619));
  NOR2_X1   g418(.A1(new_n608), .A2(KEYINPUT41), .ZN(new_n620));
  XNOR2_X1  g419(.A(G134gat), .B(G162gat), .ZN(new_n621));
  XNOR2_X1  g420(.A(new_n620), .B(new_n621), .ZN(new_n622));
  INV_X1    g421(.A(new_n618), .ZN(new_n623));
  OAI211_X1 g422(.A(new_n623), .B(new_n609), .C1(new_n615), .C2(new_n616), .ZN(new_n624));
  NAND3_X1  g423(.A1(new_n619), .A2(new_n622), .A3(new_n624), .ZN(new_n625));
  INV_X1    g424(.A(new_n625), .ZN(new_n626));
  AOI21_X1  g425(.A(new_n622), .B1(new_n619), .B2(new_n624), .ZN(new_n627));
  NOR2_X1   g426(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  NAND2_X1  g427(.A1(G71gat), .A2(G78gat), .ZN(new_n629));
  INV_X1    g428(.A(KEYINPUT9), .ZN(new_n630));
  AOI21_X1  g429(.A(KEYINPUT94), .B1(new_n629), .B2(new_n630), .ZN(new_n631));
  XOR2_X1   g430(.A(G71gat), .B(G78gat), .Z(new_n632));
  AOI21_X1  g431(.A(new_n631), .B1(new_n632), .B2(KEYINPUT95), .ZN(new_n633));
  XNOR2_X1  g432(.A(G71gat), .B(G78gat), .ZN(new_n634));
  INV_X1    g433(.A(KEYINPUT95), .ZN(new_n635));
  NAND2_X1  g434(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  NAND3_X1  g435(.A1(new_n629), .A2(KEYINPUT94), .A3(new_n630), .ZN(new_n637));
  NAND2_X1  g436(.A1(G57gat), .A2(G64gat), .ZN(new_n638));
  OR2_X1    g437(.A1(G57gat), .A2(G64gat), .ZN(new_n639));
  NAND3_X1  g438(.A1(new_n637), .A2(new_n638), .A3(new_n639), .ZN(new_n640));
  INV_X1    g439(.A(new_n640), .ZN(new_n641));
  NAND3_X1  g440(.A1(new_n633), .A2(new_n636), .A3(new_n641), .ZN(new_n642));
  OAI211_X1 g441(.A(new_n635), .B(new_n634), .C1(new_n640), .C2(new_n631), .ZN(new_n643));
  NAND2_X1  g442(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  NOR2_X1   g443(.A1(new_n644), .A2(KEYINPUT21), .ZN(new_n645));
  XNOR2_X1  g444(.A(G127gat), .B(G155gat), .ZN(new_n646));
  XNOR2_X1  g445(.A(new_n646), .B(KEYINPUT20), .ZN(new_n647));
  XNOR2_X1  g446(.A(new_n645), .B(new_n647), .ZN(new_n648));
  AOI21_X1  g447(.A(new_n537), .B1(KEYINPUT21), .B2(new_n644), .ZN(new_n649));
  XNOR2_X1  g448(.A(new_n648), .B(new_n649), .ZN(new_n650));
  XNOR2_X1  g449(.A(KEYINPUT97), .B(KEYINPUT19), .ZN(new_n651));
  XNOR2_X1  g450(.A(new_n651), .B(KEYINPUT98), .ZN(new_n652));
  NAND2_X1  g451(.A1(G231gat), .A2(G233gat), .ZN(new_n653));
  XNOR2_X1  g452(.A(new_n653), .B(KEYINPUT96), .ZN(new_n654));
  XNOR2_X1  g453(.A(new_n652), .B(new_n654), .ZN(new_n655));
  XNOR2_X1  g454(.A(G183gat), .B(G211gat), .ZN(new_n656));
  XNOR2_X1  g455(.A(new_n655), .B(new_n656), .ZN(new_n657));
  XNOR2_X1  g456(.A(new_n650), .B(new_n657), .ZN(new_n658));
  NOR2_X1   g457(.A1(new_n628), .A2(new_n658), .ZN(new_n659));
  INV_X1    g458(.A(KEYINPUT100), .ZN(new_n660));
  OR3_X1    g459(.A1(new_n607), .A2(new_n644), .A3(new_n660), .ZN(new_n661));
  NAND2_X1  g460(.A1(new_n607), .A2(new_n644), .ZN(new_n662));
  OAI211_X1 g461(.A(new_n642), .B(new_n643), .C1(new_n605), .C2(new_n606), .ZN(new_n663));
  NAND3_X1  g462(.A1(new_n662), .A2(new_n660), .A3(new_n663), .ZN(new_n664));
  AOI21_X1  g463(.A(KEYINPUT10), .B1(new_n661), .B2(new_n664), .ZN(new_n665));
  INV_X1    g464(.A(new_n665), .ZN(new_n666));
  INV_X1    g465(.A(KEYINPUT102), .ZN(new_n667));
  NAND3_X1  g466(.A1(new_n607), .A2(new_n644), .A3(KEYINPUT10), .ZN(new_n668));
  XNOR2_X1  g467(.A(new_n668), .B(KEYINPUT101), .ZN(new_n669));
  NAND3_X1  g468(.A1(new_n666), .A2(new_n667), .A3(new_n669), .ZN(new_n670));
  INV_X1    g469(.A(KEYINPUT101), .ZN(new_n671));
  XNOR2_X1  g470(.A(new_n668), .B(new_n671), .ZN(new_n672));
  OAI21_X1  g471(.A(KEYINPUT102), .B1(new_n665), .B2(new_n672), .ZN(new_n673));
  NAND2_X1  g472(.A1(G230gat), .A2(G233gat), .ZN(new_n674));
  NAND3_X1  g473(.A1(new_n670), .A2(new_n673), .A3(new_n674), .ZN(new_n675));
  INV_X1    g474(.A(new_n674), .ZN(new_n676));
  NAND3_X1  g475(.A1(new_n661), .A2(new_n664), .A3(new_n676), .ZN(new_n677));
  XOR2_X1   g476(.A(G120gat), .B(G148gat), .Z(new_n678));
  XNOR2_X1  g477(.A(new_n678), .B(KEYINPUT103), .ZN(new_n679));
  XNOR2_X1  g478(.A(G176gat), .B(G204gat), .ZN(new_n680));
  XOR2_X1   g479(.A(new_n679), .B(new_n680), .Z(new_n681));
  INV_X1    g480(.A(new_n681), .ZN(new_n682));
  AND2_X1   g481(.A1(new_n677), .A2(new_n682), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n675), .A2(new_n683), .ZN(new_n684));
  NOR2_X1   g483(.A1(new_n665), .A2(new_n672), .ZN(new_n685));
  OAI21_X1  g484(.A(new_n677), .B1(new_n685), .B2(new_n676), .ZN(new_n686));
  NAND2_X1  g485(.A1(new_n686), .A2(new_n681), .ZN(new_n687));
  NAND2_X1  g486(.A1(new_n684), .A2(new_n687), .ZN(new_n688));
  INV_X1    g487(.A(new_n688), .ZN(new_n689));
  NAND2_X1  g488(.A1(new_n659), .A2(new_n689), .ZN(new_n690));
  NAND2_X1  g489(.A1(new_n690), .A2(KEYINPUT104), .ZN(new_n691));
  INV_X1    g490(.A(KEYINPUT104), .ZN(new_n692));
  NAND3_X1  g491(.A1(new_n659), .A2(new_n692), .A3(new_n689), .ZN(new_n693));
  AND2_X1   g492(.A1(new_n691), .A2(new_n693), .ZN(new_n694));
  NAND2_X1  g493(.A1(new_n596), .A2(new_n694), .ZN(new_n695));
  NAND2_X1  g494(.A1(new_n474), .A2(new_n475), .ZN(new_n696));
  NOR2_X1   g495(.A1(new_n695), .A2(new_n696), .ZN(new_n697));
  XNOR2_X1  g496(.A(new_n697), .B(KEYINPUT106), .ZN(new_n698));
  XOR2_X1   g497(.A(KEYINPUT105), .B(G1gat), .Z(new_n699));
  XNOR2_X1  g498(.A(new_n698), .B(new_n699), .ZN(G1324gat));
  INV_X1    g499(.A(new_n695), .ZN(new_n701));
  AOI21_X1  g500(.A(new_n535), .B1(new_n701), .B2(new_n461), .ZN(new_n702));
  INV_X1    g501(.A(new_n461), .ZN(new_n703));
  XNOR2_X1  g502(.A(KEYINPUT16), .B(G8gat), .ZN(new_n704));
  NOR3_X1   g503(.A1(new_n695), .A2(new_n703), .A3(new_n704), .ZN(new_n705));
  OAI21_X1  g504(.A(KEYINPUT42), .B1(new_n702), .B2(new_n705), .ZN(new_n706));
  OAI21_X1  g505(.A(new_n706), .B1(KEYINPUT42), .B2(new_n705), .ZN(G1325gat));
  OAI21_X1  g506(.A(G15gat), .B1(new_n695), .B2(new_n494), .ZN(new_n708));
  NAND2_X1  g507(.A1(new_n295), .A2(new_n305), .ZN(new_n709));
  NAND4_X1  g508(.A1(new_n307), .A2(new_n292), .A3(new_n294), .A4(new_n304), .ZN(new_n710));
  NAND2_X1  g509(.A1(new_n709), .A2(new_n710), .ZN(new_n711));
  OR2_X1    g510(.A1(new_n711), .A2(G15gat), .ZN(new_n712));
  OAI21_X1  g511(.A(new_n708), .B1(new_n695), .B2(new_n712), .ZN(G1326gat));
  NOR2_X1   g512(.A1(new_n695), .A2(new_n380), .ZN(new_n714));
  XOR2_X1   g513(.A(KEYINPUT43), .B(G22gat), .Z(new_n715));
  XNOR2_X1  g514(.A(new_n714), .B(new_n715), .ZN(G1327gat));
  INV_X1    g515(.A(new_n628), .ZN(new_n717));
  INV_X1    g516(.A(new_n658), .ZN(new_n718));
  NOR2_X1   g517(.A1(new_n718), .A2(new_n688), .ZN(new_n719));
  INV_X1    g518(.A(new_n719), .ZN(new_n720));
  NOR4_X1   g519(.A1(new_n530), .A2(new_n595), .A3(new_n717), .A4(new_n720), .ZN(new_n721));
  INV_X1    g520(.A(new_n696), .ZN(new_n722));
  NAND3_X1  g521(.A1(new_n721), .A2(new_n538), .A3(new_n722), .ZN(new_n723));
  XNOR2_X1  g522(.A(new_n723), .B(KEYINPUT45), .ZN(new_n724));
  INV_X1    g523(.A(KEYINPUT107), .ZN(new_n725));
  AND4_X1   g524(.A1(new_n592), .A2(new_n575), .A3(new_n576), .A4(new_n581), .ZN(new_n726));
  AOI21_X1  g525(.A(new_n592), .B1(new_n591), .B2(new_n576), .ZN(new_n727));
  OAI21_X1  g526(.A(new_n725), .B1(new_n726), .B2(new_n727), .ZN(new_n728));
  NAND3_X1  g527(.A1(new_n590), .A2(KEYINPUT107), .A3(new_n593), .ZN(new_n729));
  NAND2_X1  g528(.A1(new_n728), .A2(new_n729), .ZN(new_n730));
  NOR2_X1   g529(.A1(new_n730), .A2(new_n720), .ZN(new_n731));
  INV_X1    g530(.A(new_n731), .ZN(new_n732));
  OAI211_X1 g531(.A(KEYINPUT108), .B(KEYINPUT44), .C1(new_n530), .C2(new_n717), .ZN(new_n733));
  INV_X1    g532(.A(KEYINPUT108), .ZN(new_n734));
  AOI21_X1  g533(.A(new_n380), .B1(new_n480), .B2(new_n470), .ZN(new_n735));
  XNOR2_X1  g534(.A(new_n711), .B(KEYINPUT36), .ZN(new_n736));
  OAI21_X1  g535(.A(KEYINPUT82), .B1(new_n735), .B2(new_n736), .ZN(new_n737));
  NAND2_X1  g536(.A1(new_n526), .A2(new_n513), .ZN(new_n738));
  NAND3_X1  g537(.A1(new_n737), .A2(new_n738), .A3(new_n529), .ZN(new_n739));
  OR3_X1    g538(.A1(new_n381), .A2(new_n437), .A3(new_n461), .ZN(new_n740));
  NAND2_X1  g539(.A1(new_n478), .A2(new_n479), .ZN(new_n741));
  NAND3_X1  g540(.A1(new_n696), .A2(new_n470), .A3(new_n741), .ZN(new_n742));
  OAI21_X1  g541(.A(KEYINPUT86), .B1(new_n486), .B2(new_n711), .ZN(new_n743));
  NAND3_X1  g542(.A1(new_n309), .A2(new_n481), .A3(new_n380), .ZN(new_n744));
  AOI21_X1  g543(.A(new_n742), .B1(new_n743), .B2(new_n744), .ZN(new_n745));
  OAI21_X1  g544(.A(new_n740), .B1(new_n745), .B2(new_n310), .ZN(new_n746));
  AOI21_X1  g545(.A(new_n717), .B1(new_n739), .B2(new_n746), .ZN(new_n747));
  INV_X1    g546(.A(KEYINPUT44), .ZN(new_n748));
  OAI21_X1  g547(.A(new_n734), .B1(new_n747), .B2(new_n748), .ZN(new_n749));
  NAND2_X1  g548(.A1(new_n733), .A2(new_n749), .ZN(new_n750));
  NAND2_X1  g549(.A1(new_n743), .A2(new_n744), .ZN(new_n751));
  NOR2_X1   g550(.A1(new_n489), .A2(new_n492), .ZN(new_n752));
  AOI21_X1  g551(.A(new_n310), .B1(new_n751), .B2(new_n752), .ZN(new_n753));
  OAI21_X1  g552(.A(KEYINPUT109), .B1(new_n753), .B2(new_n462), .ZN(new_n754));
  INV_X1    g553(.A(KEYINPUT109), .ZN(new_n755));
  OAI211_X1 g554(.A(new_n755), .B(new_n740), .C1(new_n745), .C2(new_n310), .ZN(new_n756));
  NOR2_X1   g555(.A1(new_n735), .A2(new_n736), .ZN(new_n757));
  NAND2_X1  g556(.A1(new_n738), .A2(new_n757), .ZN(new_n758));
  NAND3_X1  g557(.A1(new_n754), .A2(new_n756), .A3(new_n758), .ZN(new_n759));
  NAND2_X1  g558(.A1(new_n759), .A2(KEYINPUT110), .ZN(new_n760));
  AOI22_X1  g559(.A1(new_n485), .A2(new_n755), .B1(new_n757), .B2(new_n738), .ZN(new_n761));
  INV_X1    g560(.A(KEYINPUT110), .ZN(new_n762));
  NAND3_X1  g561(.A1(new_n761), .A2(new_n762), .A3(new_n754), .ZN(new_n763));
  NOR2_X1   g562(.A1(new_n717), .A2(KEYINPUT44), .ZN(new_n764));
  NAND3_X1  g563(.A1(new_n760), .A2(new_n763), .A3(new_n764), .ZN(new_n765));
  AOI21_X1  g564(.A(new_n732), .B1(new_n750), .B2(new_n765), .ZN(new_n766));
  NAND2_X1  g565(.A1(new_n766), .A2(KEYINPUT111), .ZN(new_n767));
  INV_X1    g566(.A(new_n767), .ZN(new_n768));
  NOR2_X1   g567(.A1(new_n766), .A2(KEYINPUT111), .ZN(new_n769));
  NOR3_X1   g568(.A1(new_n768), .A2(new_n769), .A3(new_n696), .ZN(new_n770));
  OAI21_X1  g569(.A(new_n724), .B1(new_n770), .B2(new_n538), .ZN(G1328gat));
  NAND3_X1  g570(.A1(new_n721), .A2(new_n549), .A3(new_n461), .ZN(new_n772));
  XOR2_X1   g571(.A(new_n772), .B(KEYINPUT46), .Z(new_n773));
  NOR3_X1   g572(.A1(new_n768), .A2(new_n769), .A3(new_n703), .ZN(new_n774));
  OAI21_X1  g573(.A(new_n773), .B1(new_n774), .B2(new_n549), .ZN(G1329gat));
  INV_X1    g574(.A(G43gat), .ZN(new_n776));
  AOI21_X1  g575(.A(new_n776), .B1(new_n766), .B2(new_n736), .ZN(new_n777));
  NOR2_X1   g576(.A1(new_n711), .A2(G43gat), .ZN(new_n778));
  NAND2_X1  g577(.A1(new_n721), .A2(new_n778), .ZN(new_n779));
  NAND2_X1  g578(.A1(new_n779), .A2(KEYINPUT47), .ZN(new_n780));
  OAI21_X1  g579(.A(KEYINPUT112), .B1(new_n777), .B2(new_n780), .ZN(new_n781));
  INV_X1    g580(.A(new_n780), .ZN(new_n782));
  INV_X1    g581(.A(KEYINPUT112), .ZN(new_n783));
  AOI211_X1 g582(.A(new_n494), .B(new_n732), .C1(new_n750), .C2(new_n765), .ZN(new_n784));
  OAI211_X1 g583(.A(new_n782), .B(new_n783), .C1(new_n784), .C2(new_n776), .ZN(new_n785));
  NAND2_X1  g584(.A1(new_n781), .A2(new_n785), .ZN(new_n786));
  INV_X1    g585(.A(new_n779), .ZN(new_n787));
  INV_X1    g586(.A(KEYINPUT111), .ZN(new_n788));
  AOI21_X1  g587(.A(new_n762), .B1(new_n761), .B2(new_n754), .ZN(new_n789));
  AND4_X1   g588(.A1(new_n762), .A2(new_n754), .A3(new_n756), .A4(new_n758), .ZN(new_n790));
  NOR2_X1   g589(.A1(new_n789), .A2(new_n790), .ZN(new_n791));
  AOI22_X1  g590(.A1(new_n791), .A2(new_n764), .B1(new_n749), .B2(new_n733), .ZN(new_n792));
  OAI21_X1  g591(.A(new_n788), .B1(new_n792), .B2(new_n732), .ZN(new_n793));
  NAND3_X1  g592(.A1(new_n793), .A2(new_n736), .A3(new_n767), .ZN(new_n794));
  AOI21_X1  g593(.A(new_n787), .B1(new_n794), .B2(G43gat), .ZN(new_n795));
  OAI21_X1  g594(.A(new_n786), .B1(new_n795), .B2(KEYINPUT47), .ZN(G1330gat));
  INV_X1    g595(.A(new_n766), .ZN(new_n797));
  OAI21_X1  g596(.A(G50gat), .B1(new_n797), .B2(new_n380), .ZN(new_n798));
  NOR2_X1   g597(.A1(new_n380), .A2(G50gat), .ZN(new_n799));
  XOR2_X1   g598(.A(new_n799), .B(KEYINPUT113), .Z(new_n800));
  NAND2_X1  g599(.A1(new_n721), .A2(new_n800), .ZN(new_n801));
  NAND3_X1  g600(.A1(new_n798), .A2(KEYINPUT48), .A3(new_n801), .ZN(new_n802));
  INV_X1    g601(.A(new_n801), .ZN(new_n803));
  NAND3_X1  g602(.A1(new_n793), .A2(new_n486), .A3(new_n767), .ZN(new_n804));
  AOI21_X1  g603(.A(new_n803), .B1(new_n804), .B2(G50gat), .ZN(new_n805));
  OAI21_X1  g604(.A(new_n802), .B1(new_n805), .B2(KEYINPUT48), .ZN(G1331gat));
  NAND4_X1  g605(.A1(new_n791), .A2(new_n659), .A3(new_n688), .A4(new_n730), .ZN(new_n807));
  INV_X1    g606(.A(new_n807), .ZN(new_n808));
  NAND2_X1  g607(.A1(new_n808), .A2(new_n722), .ZN(new_n809));
  XNOR2_X1  g608(.A(new_n809), .B(G57gat), .ZN(G1332gat));
  NOR2_X1   g609(.A1(new_n807), .A2(new_n703), .ZN(new_n811));
  NOR2_X1   g610(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n812));
  AND2_X1   g611(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n813));
  OAI21_X1  g612(.A(new_n811), .B1(new_n812), .B2(new_n813), .ZN(new_n814));
  OAI21_X1  g613(.A(new_n814), .B1(new_n811), .B2(new_n812), .ZN(G1333gat));
  OAI21_X1  g614(.A(G71gat), .B1(new_n807), .B2(new_n494), .ZN(new_n816));
  OR2_X1    g615(.A1(new_n711), .A2(G71gat), .ZN(new_n817));
  OAI21_X1  g616(.A(new_n816), .B1(new_n807), .B2(new_n817), .ZN(new_n818));
  INV_X1    g617(.A(KEYINPUT50), .ZN(new_n819));
  XNOR2_X1  g618(.A(new_n818), .B(new_n819), .ZN(G1334gat));
  NOR2_X1   g619(.A1(new_n807), .A2(new_n380), .ZN(new_n821));
  XNOR2_X1  g620(.A(KEYINPUT114), .B(G78gat), .ZN(new_n822));
  XNOR2_X1  g621(.A(new_n821), .B(new_n822), .ZN(G1335gat));
  NAND2_X1  g622(.A1(new_n750), .A2(new_n765), .ZN(new_n824));
  NAND2_X1  g623(.A1(new_n730), .A2(new_n658), .ZN(new_n825));
  NOR2_X1   g624(.A1(new_n825), .A2(new_n689), .ZN(new_n826));
  NAND2_X1  g625(.A1(new_n824), .A2(new_n826), .ZN(new_n827));
  OAI21_X1  g626(.A(G85gat), .B1(new_n827), .B2(new_n696), .ZN(new_n828));
  NOR2_X1   g627(.A1(new_n825), .A2(new_n717), .ZN(new_n829));
  NAND2_X1  g628(.A1(new_n759), .A2(new_n829), .ZN(new_n830));
  INV_X1    g629(.A(KEYINPUT51), .ZN(new_n831));
  NOR2_X1   g630(.A1(new_n830), .A2(new_n831), .ZN(new_n832));
  AOI21_X1  g631(.A(KEYINPUT51), .B1(new_n759), .B2(new_n829), .ZN(new_n833));
  NOR2_X1   g632(.A1(new_n832), .A2(new_n833), .ZN(new_n834));
  NOR2_X1   g633(.A1(new_n834), .A2(new_n689), .ZN(new_n835));
  NAND3_X1  g634(.A1(new_n835), .A2(new_n602), .A3(new_n722), .ZN(new_n836));
  NAND2_X1  g635(.A1(new_n828), .A2(new_n836), .ZN(G1336gat));
  NAND3_X1  g636(.A1(new_n835), .A2(new_n603), .A3(new_n461), .ZN(new_n838));
  NOR2_X1   g637(.A1(new_n827), .A2(new_n703), .ZN(new_n839));
  OAI21_X1  g638(.A(new_n838), .B1(new_n839), .B2(new_n603), .ZN(new_n840));
  NAND2_X1  g639(.A1(new_n840), .A2(KEYINPUT52), .ZN(new_n841));
  INV_X1    g640(.A(KEYINPUT52), .ZN(new_n842));
  OAI211_X1 g641(.A(new_n838), .B(new_n842), .C1(new_n839), .C2(new_n603), .ZN(new_n843));
  NAND2_X1  g642(.A1(new_n841), .A2(new_n843), .ZN(G1337gat));
  AND2_X1   g643(.A1(new_n824), .A2(new_n826), .ZN(new_n845));
  AND3_X1   g644(.A1(new_n845), .A2(G99gat), .A3(new_n736), .ZN(new_n846));
  AOI21_X1  g645(.A(G99gat), .B1(new_n835), .B2(new_n309), .ZN(new_n847));
  NOR2_X1   g646(.A1(new_n846), .A2(new_n847), .ZN(G1338gat));
  INV_X1    g647(.A(G106gat), .ZN(new_n849));
  AOI21_X1  g648(.A(new_n849), .B1(new_n845), .B2(new_n486), .ZN(new_n850));
  NOR2_X1   g649(.A1(new_n380), .A2(G106gat), .ZN(new_n851));
  OAI211_X1 g650(.A(new_n688), .B(new_n851), .C1(new_n832), .C2(new_n833), .ZN(new_n852));
  XNOR2_X1  g651(.A(new_n852), .B(KEYINPUT115), .ZN(new_n853));
  OAI21_X1  g652(.A(KEYINPUT53), .B1(new_n850), .B2(new_n853), .ZN(new_n854));
  NOR2_X1   g653(.A1(KEYINPUT116), .A2(KEYINPUT53), .ZN(new_n855));
  AND2_X1   g654(.A1(KEYINPUT116), .A2(KEYINPUT53), .ZN(new_n856));
  OAI21_X1  g655(.A(new_n852), .B1(new_n855), .B2(new_n856), .ZN(new_n857));
  OAI21_X1  g656(.A(new_n854), .B1(new_n850), .B2(new_n857), .ZN(G1339gat));
  INV_X1    g657(.A(KEYINPUT54), .ZN(new_n859));
  AOI21_X1  g658(.A(new_n859), .B1(new_n685), .B2(new_n676), .ZN(new_n860));
  NAND2_X1  g659(.A1(new_n675), .A2(new_n860), .ZN(new_n861));
  OAI211_X1 g660(.A(new_n859), .B(new_n674), .C1(new_n665), .C2(new_n672), .ZN(new_n862));
  AND3_X1   g661(.A1(new_n862), .A2(KEYINPUT55), .A3(new_n681), .ZN(new_n863));
  AOI22_X1  g662(.A1(new_n861), .A2(new_n863), .B1(new_n675), .B2(new_n683), .ZN(new_n864));
  NAND2_X1  g663(.A1(new_n862), .A2(new_n681), .ZN(new_n865));
  AOI21_X1  g664(.A(new_n865), .B1(new_n675), .B2(new_n860), .ZN(new_n866));
  OR2_X1    g665(.A1(new_n866), .A2(KEYINPUT55), .ZN(new_n867));
  NAND4_X1  g666(.A1(new_n728), .A2(new_n729), .A3(new_n864), .A4(new_n867), .ZN(new_n868));
  AOI21_X1  g667(.A(new_n568), .B1(new_n567), .B2(new_n572), .ZN(new_n869));
  AND3_X1   g668(.A1(new_n572), .A2(new_n579), .A3(new_n578), .ZN(new_n870));
  OAI21_X1  g669(.A(new_n587), .B1(new_n869), .B2(new_n870), .ZN(new_n871));
  NAND2_X1  g670(.A1(new_n593), .A2(new_n871), .ZN(new_n872));
  INV_X1    g671(.A(new_n872), .ZN(new_n873));
  NAND2_X1  g672(.A1(new_n873), .A2(new_n688), .ZN(new_n874));
  AOI21_X1  g673(.A(new_n628), .B1(new_n868), .B2(new_n874), .ZN(new_n875));
  INV_X1    g674(.A(new_n627), .ZN(new_n876));
  NAND3_X1  g675(.A1(new_n876), .A2(new_n873), .A3(new_n625), .ZN(new_n877));
  NAND2_X1  g676(.A1(new_n867), .A2(new_n864), .ZN(new_n878));
  NOR2_X1   g677(.A1(new_n877), .A2(new_n878), .ZN(new_n879));
  OAI21_X1  g678(.A(new_n658), .B1(new_n875), .B2(new_n879), .ZN(new_n880));
  NAND3_X1  g679(.A1(new_n659), .A2(new_n689), .A3(new_n730), .ZN(new_n881));
  AOI211_X1 g680(.A(new_n711), .B(new_n486), .C1(new_n880), .C2(new_n881), .ZN(new_n882));
  NAND3_X1  g681(.A1(new_n882), .A2(new_n722), .A3(new_n703), .ZN(new_n883));
  XNOR2_X1  g682(.A(new_n883), .B(KEYINPUT117), .ZN(new_n884));
  OAI21_X1  g683(.A(G113gat), .B1(new_n884), .B2(new_n595), .ZN(new_n885));
  AOI21_X1  g684(.A(new_n696), .B1(new_n880), .B2(new_n881), .ZN(new_n886));
  AND3_X1   g685(.A1(new_n886), .A2(new_n751), .A3(new_n703), .ZN(new_n887));
  INV_X1    g686(.A(new_n730), .ZN(new_n888));
  NAND4_X1  g687(.A1(new_n887), .A2(new_n203), .A3(new_n205), .A4(new_n888), .ZN(new_n889));
  NAND2_X1  g688(.A1(new_n885), .A2(new_n889), .ZN(G1340gat));
  NOR3_X1   g689(.A1(new_n884), .A2(new_n209), .A3(new_n689), .ZN(new_n891));
  AOI21_X1  g690(.A(G120gat), .B1(new_n887), .B2(new_n688), .ZN(new_n892));
  NOR2_X1   g691(.A1(new_n891), .A2(new_n892), .ZN(G1341gat));
  OAI21_X1  g692(.A(G127gat), .B1(new_n884), .B2(new_n658), .ZN(new_n894));
  NAND3_X1  g693(.A1(new_n887), .A2(new_n214), .A3(new_n718), .ZN(new_n895));
  NAND2_X1  g694(.A1(new_n894), .A2(new_n895), .ZN(G1342gat));
  NAND3_X1  g695(.A1(new_n887), .A2(new_n212), .A3(new_n628), .ZN(new_n897));
  XOR2_X1   g696(.A(new_n897), .B(KEYINPUT56), .Z(new_n898));
  OAI21_X1  g697(.A(G134gat), .B1(new_n884), .B2(new_n717), .ZN(new_n899));
  NAND2_X1  g698(.A1(new_n898), .A2(new_n899), .ZN(G1343gat));
  NOR3_X1   g699(.A1(new_n736), .A2(new_n696), .A3(new_n461), .ZN(new_n901));
  AOI21_X1  g700(.A(new_n380), .B1(new_n880), .B2(new_n881), .ZN(new_n902));
  XOR2_X1   g701(.A(KEYINPUT118), .B(KEYINPUT57), .Z(new_n903));
  INV_X1    g702(.A(new_n903), .ZN(new_n904));
  OAI21_X1  g703(.A(KEYINPUT119), .B1(new_n902), .B2(new_n904), .ZN(new_n905));
  OR3_X1    g704(.A1(new_n866), .A2(KEYINPUT121), .A3(KEYINPUT55), .ZN(new_n906));
  OAI21_X1  g705(.A(KEYINPUT121), .B1(new_n866), .B2(KEYINPUT55), .ZN(new_n907));
  AND4_X1   g706(.A1(new_n594), .A2(new_n906), .A3(new_n864), .A4(new_n907), .ZN(new_n908));
  NAND3_X1  g707(.A1(new_n873), .A2(KEYINPUT120), .A3(new_n688), .ZN(new_n909));
  INV_X1    g708(.A(KEYINPUT120), .ZN(new_n910));
  OAI21_X1  g709(.A(new_n910), .B1(new_n689), .B2(new_n872), .ZN(new_n911));
  NAND2_X1  g710(.A1(new_n909), .A2(new_n911), .ZN(new_n912));
  OAI21_X1  g711(.A(new_n717), .B1(new_n908), .B2(new_n912), .ZN(new_n913));
  INV_X1    g712(.A(new_n879), .ZN(new_n914));
  AOI21_X1  g713(.A(new_n718), .B1(new_n913), .B2(new_n914), .ZN(new_n915));
  INV_X1    g714(.A(new_n881), .ZN(new_n916));
  OAI211_X1 g715(.A(KEYINPUT57), .B(new_n486), .C1(new_n915), .C2(new_n916), .ZN(new_n917));
  NAND2_X1  g716(.A1(new_n905), .A2(new_n917), .ZN(new_n918));
  NOR3_X1   g717(.A1(new_n902), .A2(KEYINPUT119), .A3(new_n904), .ZN(new_n919));
  OAI211_X1 g718(.A(new_n888), .B(new_n901), .C1(new_n918), .C2(new_n919), .ZN(new_n920));
  NAND2_X1  g719(.A1(new_n920), .A2(G141gat), .ZN(new_n921));
  NOR3_X1   g720(.A1(new_n736), .A2(new_n380), .A3(new_n461), .ZN(new_n922));
  AND2_X1   g721(.A1(new_n886), .A2(new_n922), .ZN(new_n923));
  NAND3_X1  g722(.A1(new_n923), .A2(new_n318), .A3(new_n594), .ZN(new_n924));
  NAND2_X1  g723(.A1(new_n921), .A2(new_n924), .ZN(new_n925));
  NAND2_X1  g724(.A1(new_n925), .A2(KEYINPUT58), .ZN(new_n926));
  OAI211_X1 g725(.A(new_n594), .B(new_n901), .C1(new_n918), .C2(new_n919), .ZN(new_n927));
  NAND2_X1  g726(.A1(new_n927), .A2(KEYINPUT122), .ZN(new_n928));
  NOR2_X1   g727(.A1(new_n902), .A2(new_n904), .ZN(new_n929));
  INV_X1    g728(.A(KEYINPUT119), .ZN(new_n930));
  NAND2_X1  g729(.A1(new_n929), .A2(new_n930), .ZN(new_n931));
  NAND3_X1  g730(.A1(new_n931), .A2(new_n917), .A3(new_n905), .ZN(new_n932));
  INV_X1    g731(.A(KEYINPUT122), .ZN(new_n933));
  NAND4_X1  g732(.A1(new_n932), .A2(new_n933), .A3(new_n594), .A4(new_n901), .ZN(new_n934));
  AND3_X1   g733(.A1(new_n928), .A2(G141gat), .A3(new_n934), .ZN(new_n935));
  INV_X1    g734(.A(KEYINPUT58), .ZN(new_n936));
  NAND2_X1  g735(.A1(new_n924), .A2(new_n936), .ZN(new_n937));
  OAI21_X1  g736(.A(new_n926), .B1(new_n935), .B2(new_n937), .ZN(G1344gat));
  NOR2_X1   g737(.A1(new_n319), .A2(KEYINPUT59), .ZN(new_n939));
  NAND2_X1  g738(.A1(new_n932), .A2(new_n901), .ZN(new_n940));
  OAI21_X1  g739(.A(new_n939), .B1(new_n940), .B2(new_n689), .ZN(new_n941));
  NAND2_X1  g740(.A1(new_n901), .A2(new_n688), .ZN(new_n942));
  AND3_X1   g741(.A1(new_n691), .A2(new_n595), .A3(new_n693), .ZN(new_n943));
  OAI21_X1  g742(.A(new_n486), .B1(new_n943), .B2(new_n915), .ZN(new_n944));
  INV_X1    g743(.A(KEYINPUT57), .ZN(new_n945));
  NAND2_X1  g744(.A1(new_n944), .A2(new_n945), .ZN(new_n946));
  NAND2_X1  g745(.A1(new_n902), .A2(new_n904), .ZN(new_n947));
  AOI21_X1  g746(.A(new_n942), .B1(new_n946), .B2(new_n947), .ZN(new_n948));
  OAI21_X1  g747(.A(KEYINPUT59), .B1(new_n948), .B2(new_n319), .ZN(new_n949));
  NAND2_X1  g748(.A1(new_n941), .A2(new_n949), .ZN(new_n950));
  NAND3_X1  g749(.A1(new_n923), .A2(new_n319), .A3(new_n688), .ZN(new_n951));
  NAND2_X1  g750(.A1(new_n950), .A2(new_n951), .ZN(G1345gat));
  OAI21_X1  g751(.A(G155gat), .B1(new_n940), .B2(new_n658), .ZN(new_n953));
  INV_X1    g752(.A(G155gat), .ZN(new_n954));
  NAND3_X1  g753(.A1(new_n923), .A2(new_n954), .A3(new_n718), .ZN(new_n955));
  NAND2_X1  g754(.A1(new_n953), .A2(new_n955), .ZN(G1346gat));
  INV_X1    g755(.A(G162gat), .ZN(new_n957));
  NOR3_X1   g756(.A1(new_n940), .A2(new_n957), .A3(new_n717), .ZN(new_n958));
  AOI21_X1  g757(.A(G162gat), .B1(new_n923), .B2(new_n628), .ZN(new_n959));
  NOR2_X1   g758(.A1(new_n958), .A2(new_n959), .ZN(G1347gat));
  AOI211_X1 g759(.A(new_n722), .B(new_n703), .C1(new_n880), .C2(new_n881), .ZN(new_n961));
  NAND2_X1  g760(.A1(new_n961), .A2(new_n751), .ZN(new_n962));
  INV_X1    g761(.A(new_n962), .ZN(new_n963));
  NAND3_X1  g762(.A1(new_n963), .A2(new_n227), .A3(new_n888), .ZN(new_n964));
  XNOR2_X1  g763(.A(new_n964), .B(KEYINPUT123), .ZN(new_n965));
  NOR2_X1   g764(.A1(new_n722), .A2(new_n703), .ZN(new_n966));
  NAND2_X1  g765(.A1(new_n882), .A2(new_n966), .ZN(new_n967));
  OAI21_X1  g766(.A(G169gat), .B1(new_n967), .B2(new_n595), .ZN(new_n968));
  NAND2_X1  g767(.A1(new_n965), .A2(new_n968), .ZN(G1348gat));
  OAI21_X1  g768(.A(G176gat), .B1(new_n967), .B2(new_n689), .ZN(new_n970));
  NAND2_X1  g769(.A1(new_n688), .A2(new_n228), .ZN(new_n971));
  OAI21_X1  g770(.A(new_n970), .B1(new_n962), .B2(new_n971), .ZN(G1349gat));
  OAI21_X1  g771(.A(G183gat), .B1(new_n967), .B2(new_n658), .ZN(new_n973));
  NAND3_X1  g772(.A1(new_n718), .A2(new_n245), .A3(new_n247), .ZN(new_n974));
  OAI21_X1  g773(.A(new_n973), .B1(new_n962), .B2(new_n974), .ZN(new_n975));
  XNOR2_X1  g774(.A(KEYINPUT124), .B(KEYINPUT60), .ZN(new_n976));
  XNOR2_X1  g775(.A(new_n975), .B(new_n976), .ZN(G1350gat));
  OAI21_X1  g776(.A(G190gat), .B1(new_n967), .B2(new_n717), .ZN(new_n978));
  XNOR2_X1  g777(.A(new_n978), .B(KEYINPUT61), .ZN(new_n979));
  NAND3_X1  g778(.A1(new_n963), .A2(new_n248), .A3(new_n628), .ZN(new_n980));
  NAND2_X1  g779(.A1(new_n979), .A2(new_n980), .ZN(G1351gat));
  NOR3_X1   g780(.A1(new_n736), .A2(new_n703), .A3(new_n722), .ZN(new_n982));
  INV_X1    g781(.A(new_n946), .ZN(new_n983));
  INV_X1    g782(.A(new_n947), .ZN(new_n984));
  OAI21_X1  g783(.A(new_n982), .B1(new_n983), .B2(new_n984), .ZN(new_n985));
  OAI21_X1  g784(.A(G197gat), .B1(new_n985), .B2(new_n595), .ZN(new_n986));
  NOR2_X1   g785(.A1(new_n736), .A2(new_n380), .ZN(new_n987));
  NAND2_X1  g786(.A1(new_n961), .A2(new_n987), .ZN(new_n988));
  NOR3_X1   g787(.A1(new_n988), .A2(G197gat), .A3(new_n730), .ZN(new_n989));
  XNOR2_X1  g788(.A(new_n989), .B(KEYINPUT125), .ZN(new_n990));
  NAND2_X1  g789(.A1(new_n986), .A2(new_n990), .ZN(G1352gat));
  NAND4_X1  g790(.A1(new_n961), .A2(new_n331), .A3(new_n688), .A4(new_n987), .ZN(new_n992));
  OR2_X1    g791(.A1(new_n992), .A2(KEYINPUT126), .ZN(new_n993));
  INV_X1    g792(.A(KEYINPUT62), .ZN(new_n994));
  NAND2_X1  g793(.A1(new_n992), .A2(KEYINPUT126), .ZN(new_n995));
  NAND3_X1  g794(.A1(new_n993), .A2(new_n994), .A3(new_n995), .ZN(new_n996));
  OAI21_X1  g795(.A(G204gat), .B1(new_n985), .B2(new_n689), .ZN(new_n997));
  INV_X1    g796(.A(KEYINPUT127), .ZN(new_n998));
  NAND2_X1  g797(.A1(new_n993), .A2(new_n995), .ZN(new_n999));
  AOI21_X1  g798(.A(new_n998), .B1(new_n999), .B2(KEYINPUT62), .ZN(new_n1000));
  AOI211_X1 g799(.A(KEYINPUT127), .B(new_n994), .C1(new_n993), .C2(new_n995), .ZN(new_n1001));
  OAI211_X1 g800(.A(new_n996), .B(new_n997), .C1(new_n1000), .C2(new_n1001), .ZN(G1353gat));
  OR3_X1    g801(.A1(new_n988), .A2(G211gat), .A3(new_n658), .ZN(new_n1003));
  OAI211_X1 g802(.A(new_n718), .B(new_n982), .C1(new_n983), .C2(new_n984), .ZN(new_n1004));
  AND3_X1   g803(.A1(new_n1004), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n1005));
  AOI21_X1  g804(.A(KEYINPUT63), .B1(new_n1004), .B2(G211gat), .ZN(new_n1006));
  OAI21_X1  g805(.A(new_n1003), .B1(new_n1005), .B2(new_n1006), .ZN(G1354gat));
  OAI21_X1  g806(.A(G218gat), .B1(new_n985), .B2(new_n717), .ZN(new_n1008));
  OR2_X1    g807(.A1(new_n717), .A2(G218gat), .ZN(new_n1009));
  OAI21_X1  g808(.A(new_n1008), .B1(new_n988), .B2(new_n1009), .ZN(G1355gat));
endmodule


