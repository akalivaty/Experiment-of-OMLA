//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 1 1 0 1 0 1 0 0 1 0 0 0 0 0 0 0 0 1 1 0 1 1 1 0 0 1 1 0 1 0 1 1 0 1 1 1 1 1 0 0 0 1 1 1 1 0 0 0 0 0 0 0 1 0 0 1 1 1 0 1 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:38:04 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n238, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n245, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1087,
    new_n1088, new_n1089, new_n1090, new_n1091, new_n1092, new_n1093,
    new_n1094, new_n1095, new_n1096, new_n1097, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1108, new_n1109, new_n1110, new_n1111, new_n1112,
    new_n1113, new_n1114, new_n1115, new_n1116, new_n1117, new_n1118,
    new_n1119, new_n1120, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1251, new_n1252,
    new_n1253, new_n1254, new_n1255, new_n1256, new_n1257, new_n1258,
    new_n1260, new_n1261, new_n1262, new_n1263, new_n1264, new_n1265,
    new_n1266, new_n1267, new_n1268, new_n1269, new_n1270, new_n1271,
    new_n1272, new_n1273, new_n1274, new_n1275, new_n1276, new_n1277,
    new_n1278, new_n1279, new_n1280, new_n1281, new_n1282, new_n1283,
    new_n1284, new_n1285, new_n1286, new_n1288, new_n1289, new_n1290,
    new_n1291, new_n1292, new_n1293, new_n1294, new_n1295, new_n1296,
    new_n1297, new_n1298, new_n1299, new_n1300, new_n1302, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1346,
    new_n1348, new_n1349, new_n1350, new_n1351, new_n1352, new_n1353,
    new_n1354, new_n1355;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0005(.A1(G1), .A2(G20), .ZN(new_n206));
  NOR2_X1   g0006(.A1(new_n206), .A2(G13), .ZN(new_n207));
  OAI211_X1 g0007(.A(new_n207), .B(G250), .C1(G257), .C2(G264), .ZN(new_n208));
  XNOR2_X1  g0008(.A(new_n208), .B(KEYINPUT0), .ZN(new_n209));
  INV_X1    g0009(.A(new_n201), .ZN(new_n210));
  NAND2_X1  g0010(.A1(new_n210), .A2(G50), .ZN(new_n211));
  INV_X1    g0011(.A(new_n211), .ZN(new_n212));
  NAND2_X1  g0012(.A1(G1), .A2(G13), .ZN(new_n213));
  INV_X1    g0013(.A(G20), .ZN(new_n214));
  NOR2_X1   g0014(.A1(new_n213), .A2(new_n214), .ZN(new_n215));
  NAND2_X1  g0015(.A1(new_n212), .A2(new_n215), .ZN(new_n216));
  AOI22_X1  g0016(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n217));
  INV_X1    g0017(.A(G68), .ZN(new_n218));
  INV_X1    g0018(.A(G238), .ZN(new_n219));
  INV_X1    g0019(.A(G87), .ZN(new_n220));
  INV_X1    g0020(.A(G250), .ZN(new_n221));
  OAI221_X1 g0021(.A(new_n217), .B1(new_n218), .B2(new_n219), .C1(new_n220), .C2(new_n221), .ZN(new_n222));
  AOI22_X1  g0022(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n223));
  AOI22_X1  g0023(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n224));
  NAND2_X1  g0024(.A1(new_n223), .A2(new_n224), .ZN(new_n225));
  OAI21_X1  g0025(.A(new_n206), .B1(new_n222), .B2(new_n225), .ZN(new_n226));
  OAI211_X1 g0026(.A(new_n209), .B(new_n216), .C1(KEYINPUT1), .C2(new_n226), .ZN(new_n227));
  AOI21_X1  g0027(.A(new_n227), .B1(KEYINPUT1), .B2(new_n226), .ZN(G361));
  XOR2_X1   g0028(.A(G238), .B(G244), .Z(new_n229));
  XNOR2_X1  g0029(.A(G226), .B(G232), .ZN(new_n230));
  XNOR2_X1  g0030(.A(new_n229), .B(new_n230), .ZN(new_n231));
  XNOR2_X1  g0031(.A(KEYINPUT64), .B(KEYINPUT2), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n231), .B(new_n232), .ZN(new_n233));
  XOR2_X1   g0033(.A(G264), .B(G270), .Z(new_n234));
  XNOR2_X1  g0034(.A(G250), .B(G257), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n233), .B(new_n236), .ZN(G358));
  XOR2_X1   g0037(.A(G87), .B(G97), .Z(new_n238));
  XOR2_X1   g0038(.A(G107), .B(G116), .Z(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  NAND2_X1  g0040(.A1(new_n202), .A2(G68), .ZN(new_n241));
  NAND2_X1  g0041(.A1(new_n218), .A2(G50), .ZN(new_n242));
  NAND2_X1  g0042(.A1(new_n241), .A2(new_n242), .ZN(new_n243));
  XNOR2_X1  g0043(.A(G58), .B(G77), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XOR2_X1   g0045(.A(new_n240), .B(new_n245), .Z(G351));
  INV_X1    g0046(.A(G169), .ZN(new_n247));
  INV_X1    g0047(.A(KEYINPUT3), .ZN(new_n248));
  INV_X1    g0048(.A(G33), .ZN(new_n249));
  NAND2_X1  g0049(.A1(new_n248), .A2(new_n249), .ZN(new_n250));
  NAND2_X1  g0050(.A1(KEYINPUT3), .A2(G33), .ZN(new_n251));
  NAND2_X1  g0051(.A1(new_n250), .A2(new_n251), .ZN(new_n252));
  INV_X1    g0052(.A(G232), .ZN(new_n253));
  NAND2_X1  g0053(.A1(new_n253), .A2(G1698), .ZN(new_n254));
  OAI211_X1 g0054(.A(new_n252), .B(new_n254), .C1(G226), .C2(G1698), .ZN(new_n255));
  INV_X1    g0055(.A(KEYINPUT73), .ZN(new_n256));
  NAND2_X1  g0056(.A1(G33), .A2(G97), .ZN(new_n257));
  AND3_X1   g0057(.A1(new_n255), .A2(new_n256), .A3(new_n257), .ZN(new_n258));
  AOI21_X1  g0058(.A(new_n256), .B1(new_n255), .B2(new_n257), .ZN(new_n259));
  NAND2_X1  g0059(.A1(G33), .A2(G41), .ZN(new_n260));
  NAND3_X1  g0060(.A1(new_n260), .A2(G1), .A3(G13), .ZN(new_n261));
  NOR3_X1   g0061(.A1(new_n258), .A2(new_n259), .A3(new_n261), .ZN(new_n262));
  INV_X1    g0062(.A(new_n262), .ZN(new_n263));
  INV_X1    g0063(.A(G1), .ZN(new_n264));
  OAI21_X1  g0064(.A(new_n264), .B1(G41), .B2(G45), .ZN(new_n265));
  AND3_X1   g0065(.A1(new_n261), .A2(KEYINPUT75), .A3(new_n265), .ZN(new_n266));
  AOI21_X1  g0066(.A(KEYINPUT75), .B1(new_n261), .B2(new_n265), .ZN(new_n267));
  NOR3_X1   g0067(.A1(new_n266), .A2(new_n267), .A3(new_n219), .ZN(new_n268));
  AND2_X1   g0068(.A1(G33), .A2(G41), .ZN(new_n269));
  OAI21_X1  g0069(.A(G274), .B1(new_n269), .B2(new_n213), .ZN(new_n270));
  INV_X1    g0070(.A(KEYINPUT65), .ZN(new_n271));
  NOR3_X1   g0071(.A1(new_n270), .A2(new_n271), .A3(new_n265), .ZN(new_n272));
  INV_X1    g0072(.A(G274), .ZN(new_n273));
  AND2_X1   g0073(.A1(G1), .A2(G13), .ZN(new_n274));
  AOI21_X1  g0074(.A(new_n273), .B1(new_n274), .B2(new_n260), .ZN(new_n275));
  INV_X1    g0075(.A(new_n265), .ZN(new_n276));
  AOI21_X1  g0076(.A(KEYINPUT65), .B1(new_n275), .B2(new_n276), .ZN(new_n277));
  OAI21_X1  g0077(.A(KEYINPUT74), .B1(new_n272), .B2(new_n277), .ZN(new_n278));
  OAI21_X1  g0078(.A(new_n271), .B1(new_n270), .B2(new_n265), .ZN(new_n279));
  INV_X1    g0079(.A(KEYINPUT74), .ZN(new_n280));
  NAND3_X1  g0080(.A1(new_n275), .A2(KEYINPUT65), .A3(new_n276), .ZN(new_n281));
  NAND3_X1  g0081(.A1(new_n279), .A2(new_n280), .A3(new_n281), .ZN(new_n282));
  AOI211_X1 g0082(.A(KEYINPUT76), .B(new_n268), .C1(new_n278), .C2(new_n282), .ZN(new_n283));
  INV_X1    g0083(.A(KEYINPUT76), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n278), .A2(new_n282), .ZN(new_n285));
  OR3_X1    g0085(.A1(new_n266), .A2(new_n267), .A3(new_n219), .ZN(new_n286));
  AOI21_X1  g0086(.A(new_n284), .B1(new_n285), .B2(new_n286), .ZN(new_n287));
  OAI21_X1  g0087(.A(new_n263), .B1(new_n283), .B2(new_n287), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n288), .A2(KEYINPUT13), .ZN(new_n289));
  AND3_X1   g0089(.A1(new_n279), .A2(new_n280), .A3(new_n281), .ZN(new_n290));
  AOI21_X1  g0090(.A(new_n280), .B1(new_n279), .B2(new_n281), .ZN(new_n291));
  OAI21_X1  g0091(.A(new_n286), .B1(new_n290), .B2(new_n291), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n292), .A2(KEYINPUT76), .ZN(new_n293));
  NAND3_X1  g0093(.A1(new_n285), .A2(new_n284), .A3(new_n286), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n293), .A2(new_n294), .ZN(new_n295));
  INV_X1    g0095(.A(KEYINPUT13), .ZN(new_n296));
  NAND3_X1  g0096(.A1(new_n295), .A2(new_n296), .A3(new_n263), .ZN(new_n297));
  AOI21_X1  g0097(.A(new_n247), .B1(new_n289), .B2(new_n297), .ZN(new_n298));
  INV_X1    g0098(.A(KEYINPUT14), .ZN(new_n299));
  AOI21_X1  g0099(.A(new_n296), .B1(new_n295), .B2(new_n263), .ZN(new_n300));
  AOI211_X1 g0100(.A(KEYINPUT13), .B(new_n262), .C1(new_n293), .C2(new_n294), .ZN(new_n301));
  NOR2_X1   g0101(.A1(new_n300), .A2(new_n301), .ZN(new_n302));
  AOI22_X1  g0102(.A1(new_n298), .A2(new_n299), .B1(new_n302), .B2(G179), .ZN(new_n303));
  INV_X1    g0103(.A(KEYINPUT79), .ZN(new_n304));
  NOR3_X1   g0104(.A1(new_n298), .A2(new_n304), .A3(new_n299), .ZN(new_n305));
  OAI21_X1  g0105(.A(G169), .B1(new_n300), .B2(new_n301), .ZN(new_n306));
  AOI21_X1  g0106(.A(KEYINPUT79), .B1(new_n306), .B2(KEYINPUT14), .ZN(new_n307));
  OAI21_X1  g0107(.A(new_n303), .B1(new_n305), .B2(new_n307), .ZN(new_n308));
  NOR2_X1   g0108(.A1(new_n249), .A2(G20), .ZN(new_n309));
  AOI22_X1  g0109(.A1(new_n309), .A2(G77), .B1(G20), .B2(new_n218), .ZN(new_n310));
  NOR2_X1   g0110(.A1(G20), .A2(G33), .ZN(new_n311));
  INV_X1    g0111(.A(new_n311), .ZN(new_n312));
  OAI21_X1  g0112(.A(new_n310), .B1(new_n202), .B2(new_n312), .ZN(new_n313));
  NAND3_X1  g0113(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n314), .A2(new_n213), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n313), .A2(new_n315), .ZN(new_n316));
  XNOR2_X1  g0116(.A(new_n316), .B(KEYINPUT11), .ZN(new_n317));
  NAND3_X1  g0117(.A1(new_n264), .A2(G13), .A3(G20), .ZN(new_n318));
  INV_X1    g0118(.A(KEYINPUT68), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n318), .A2(new_n319), .ZN(new_n320));
  NAND4_X1  g0120(.A1(new_n264), .A2(KEYINPUT68), .A3(G13), .A4(G20), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n320), .A2(new_n321), .ZN(new_n322));
  INV_X1    g0122(.A(new_n322), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n323), .A2(new_n218), .ZN(new_n324));
  XNOR2_X1  g0124(.A(new_n324), .B(KEYINPUT12), .ZN(new_n325));
  NOR2_X1   g0125(.A1(new_n323), .A2(new_n315), .ZN(new_n326));
  OAI211_X1 g0126(.A(new_n326), .B(G68), .C1(G1), .C2(new_n214), .ZN(new_n327));
  NAND3_X1  g0127(.A1(new_n317), .A2(new_n325), .A3(new_n327), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n328), .A2(KEYINPUT77), .ZN(new_n329));
  INV_X1    g0129(.A(KEYINPUT77), .ZN(new_n330));
  NAND4_X1  g0130(.A1(new_n317), .A2(new_n325), .A3(new_n330), .A4(new_n327), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n329), .A2(new_n331), .ZN(new_n332));
  INV_X1    g0132(.A(new_n332), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n308), .A2(new_n333), .ZN(new_n334));
  INV_X1    g0134(.A(new_n334), .ZN(new_n335));
  OAI21_X1  g0135(.A(G200), .B1(new_n300), .B2(new_n301), .ZN(new_n336));
  NAND3_X1  g0136(.A1(new_n289), .A2(G190), .A3(new_n297), .ZN(new_n337));
  NAND3_X1  g0137(.A1(new_n336), .A2(new_n337), .A3(new_n332), .ZN(new_n338));
  INV_X1    g0138(.A(KEYINPUT78), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n338), .A2(new_n339), .ZN(new_n340));
  NAND4_X1  g0140(.A1(new_n336), .A2(new_n337), .A3(KEYINPUT78), .A4(new_n332), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n340), .A2(new_n341), .ZN(new_n342));
  XNOR2_X1  g0142(.A(KEYINPUT8), .B(G58), .ZN(new_n343));
  NAND2_X1  g0143(.A1(new_n343), .A2(KEYINPUT66), .ZN(new_n344));
  INV_X1    g0144(.A(G58), .ZN(new_n345));
  OR3_X1    g0145(.A1(new_n345), .A2(KEYINPUT66), .A3(KEYINPUT8), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n344), .A2(new_n346), .ZN(new_n347));
  AOI21_X1  g0147(.A(new_n347), .B1(new_n264), .B2(G20), .ZN(new_n348));
  AOI22_X1  g0148(.A1(new_n348), .A2(new_n326), .B1(new_n323), .B2(new_n347), .ZN(new_n349));
  INV_X1    g0149(.A(KEYINPUT16), .ZN(new_n350));
  NOR2_X1   g0150(.A1(new_n345), .A2(new_n218), .ZN(new_n351));
  OAI21_X1  g0151(.A(G20), .B1(new_n351), .B2(new_n201), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n311), .A2(G159), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n352), .A2(new_n353), .ZN(new_n354));
  NAND3_X1  g0154(.A1(new_n250), .A2(new_n214), .A3(new_n251), .ZN(new_n355));
  INV_X1    g0155(.A(KEYINPUT7), .ZN(new_n356));
  INV_X1    g0156(.A(KEYINPUT80), .ZN(new_n357));
  NOR2_X1   g0157(.A1(new_n357), .A2(KEYINPUT7), .ZN(new_n358));
  NAND3_X1  g0158(.A1(new_n355), .A2(new_n356), .A3(new_n358), .ZN(new_n359));
  AND2_X1   g0159(.A1(new_n359), .A2(G68), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n355), .A2(new_n356), .ZN(new_n361));
  NAND4_X1  g0161(.A1(new_n250), .A2(KEYINPUT7), .A3(new_n214), .A4(new_n251), .ZN(new_n362));
  NAND3_X1  g0162(.A1(new_n361), .A2(new_n357), .A3(new_n362), .ZN(new_n363));
  AOI211_X1 g0163(.A(new_n350), .B(new_n354), .C1(new_n360), .C2(new_n363), .ZN(new_n364));
  AOI21_X1  g0164(.A(new_n218), .B1(new_n361), .B2(new_n362), .ZN(new_n365));
  OAI21_X1  g0165(.A(new_n350), .B1(new_n365), .B2(new_n354), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n366), .A2(new_n315), .ZN(new_n367));
  OAI21_X1  g0167(.A(new_n349), .B1(new_n364), .B2(new_n367), .ZN(new_n368));
  INV_X1    g0168(.A(G1698), .ZN(new_n369));
  AND2_X1   g0169(.A1(KEYINPUT3), .A2(G33), .ZN(new_n370));
  NOR2_X1   g0170(.A1(KEYINPUT3), .A2(G33), .ZN(new_n371));
  OAI211_X1 g0171(.A(G223), .B(new_n369), .C1(new_n370), .C2(new_n371), .ZN(new_n372));
  INV_X1    g0172(.A(KEYINPUT81), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n372), .A2(new_n373), .ZN(new_n374));
  NAND4_X1  g0174(.A1(new_n252), .A2(KEYINPUT81), .A3(G223), .A4(new_n369), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n374), .A2(new_n375), .ZN(new_n376));
  AOI21_X1  g0176(.A(new_n369), .B1(new_n250), .B2(new_n251), .ZN(new_n377));
  AOI22_X1  g0177(.A1(new_n377), .A2(G226), .B1(G33), .B2(G87), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n376), .A2(new_n378), .ZN(new_n379));
  INV_X1    g0179(.A(new_n261), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n379), .A2(new_n380), .ZN(new_n381));
  INV_X1    g0181(.A(G179), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n261), .A2(new_n265), .ZN(new_n383));
  OAI22_X1  g0183(.A1(new_n272), .A2(new_n277), .B1(new_n253), .B2(new_n383), .ZN(new_n384));
  INV_X1    g0184(.A(new_n384), .ZN(new_n385));
  NAND3_X1  g0185(.A1(new_n381), .A2(new_n382), .A3(new_n385), .ZN(new_n386));
  AOI21_X1  g0186(.A(new_n261), .B1(new_n376), .B2(new_n378), .ZN(new_n387));
  OAI21_X1  g0187(.A(new_n247), .B1(new_n387), .B2(new_n384), .ZN(new_n388));
  INV_X1    g0188(.A(KEYINPUT82), .ZN(new_n389));
  AND3_X1   g0189(.A1(new_n386), .A2(new_n388), .A3(new_n389), .ZN(new_n390));
  AOI21_X1  g0190(.A(new_n389), .B1(new_n386), .B2(new_n388), .ZN(new_n391));
  OAI21_X1  g0191(.A(new_n368), .B1(new_n390), .B2(new_n391), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n392), .A2(KEYINPUT18), .ZN(new_n393));
  INV_X1    g0193(.A(KEYINPUT17), .ZN(new_n394));
  AOI21_X1  g0194(.A(new_n354), .B1(new_n360), .B2(new_n363), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n395), .A2(KEYINPUT16), .ZN(new_n396));
  NAND3_X1  g0196(.A1(new_n396), .A2(new_n315), .A3(new_n366), .ZN(new_n397));
  NAND3_X1  g0197(.A1(new_n381), .A2(G190), .A3(new_n385), .ZN(new_n398));
  OAI21_X1  g0198(.A(G200), .B1(new_n387), .B2(new_n384), .ZN(new_n399));
  NAND4_X1  g0199(.A1(new_n397), .A2(new_n349), .A3(new_n398), .A4(new_n399), .ZN(new_n400));
  INV_X1    g0200(.A(KEYINPUT83), .ZN(new_n401));
  OAI21_X1  g0201(.A(new_n394), .B1(new_n400), .B2(new_n401), .ZN(new_n402));
  AOI21_X1  g0202(.A(G169), .B1(new_n381), .B2(new_n385), .ZN(new_n403));
  NOR3_X1   g0203(.A1(new_n387), .A2(G179), .A3(new_n384), .ZN(new_n404));
  OAI21_X1  g0204(.A(KEYINPUT82), .B1(new_n403), .B2(new_n404), .ZN(new_n405));
  NAND3_X1  g0205(.A1(new_n386), .A2(new_n388), .A3(new_n389), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n405), .A2(new_n406), .ZN(new_n407));
  INV_X1    g0207(.A(KEYINPUT18), .ZN(new_n408));
  NAND3_X1  g0208(.A1(new_n407), .A2(new_n408), .A3(new_n368), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n398), .A2(new_n399), .ZN(new_n410));
  NOR2_X1   g0210(.A1(new_n368), .A2(new_n410), .ZN(new_n411));
  NAND3_X1  g0211(.A1(new_n411), .A2(KEYINPUT83), .A3(KEYINPUT17), .ZN(new_n412));
  NAND4_X1  g0212(.A1(new_n393), .A2(new_n402), .A3(new_n409), .A4(new_n412), .ZN(new_n413));
  NAND2_X1  g0213(.A1(new_n279), .A2(new_n281), .ZN(new_n414));
  INV_X1    g0214(.A(new_n383), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n415), .A2(G226), .ZN(new_n416));
  AND2_X1   g0216(.A1(new_n414), .A2(new_n416), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n377), .A2(G223), .ZN(new_n418));
  NAND3_X1  g0218(.A1(new_n252), .A2(G222), .A3(new_n369), .ZN(new_n419));
  NOR2_X1   g0219(.A1(new_n370), .A2(new_n371), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n420), .A2(G77), .ZN(new_n421));
  NAND3_X1  g0221(.A1(new_n418), .A2(new_n419), .A3(new_n421), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n422), .A2(new_n380), .ZN(new_n423));
  NAND4_X1  g0223(.A1(new_n417), .A2(KEYINPUT72), .A3(G190), .A4(new_n423), .ZN(new_n424));
  NAND4_X1  g0224(.A1(new_n423), .A2(G190), .A3(new_n414), .A4(new_n416), .ZN(new_n425));
  INV_X1    g0225(.A(KEYINPUT72), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n425), .A2(new_n426), .ZN(new_n427));
  INV_X1    g0227(.A(G200), .ZN(new_n428));
  AOI21_X1  g0228(.A(new_n428), .B1(new_n417), .B2(new_n423), .ZN(new_n429));
  OAI21_X1  g0229(.A(new_n424), .B1(new_n427), .B2(new_n429), .ZN(new_n430));
  NAND3_X1  g0230(.A1(new_n344), .A2(new_n309), .A3(new_n346), .ZN(new_n431));
  INV_X1    g0231(.A(KEYINPUT67), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n311), .A2(G150), .ZN(new_n433));
  NAND3_X1  g0233(.A1(new_n431), .A2(new_n432), .A3(new_n433), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n203), .A2(G20), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n434), .A2(new_n435), .ZN(new_n436));
  AOI21_X1  g0236(.A(new_n432), .B1(new_n431), .B2(new_n433), .ZN(new_n437));
  OAI21_X1  g0237(.A(new_n315), .B1(new_n436), .B2(new_n437), .ZN(new_n438));
  INV_X1    g0238(.A(KEYINPUT9), .ZN(new_n439));
  AOI21_X1  g0239(.A(new_n202), .B1(new_n264), .B2(G20), .ZN(new_n440));
  AOI22_X1  g0240(.A1(new_n326), .A2(new_n440), .B1(new_n202), .B2(new_n323), .ZN(new_n441));
  AND3_X1   g0241(.A1(new_n438), .A2(new_n439), .A3(new_n441), .ZN(new_n442));
  AOI21_X1  g0242(.A(new_n439), .B1(new_n438), .B2(new_n441), .ZN(new_n443));
  OAI21_X1  g0243(.A(new_n430), .B1(new_n442), .B2(new_n443), .ZN(new_n444));
  INV_X1    g0244(.A(KEYINPUT71), .ZN(new_n445));
  AOI21_X1  g0245(.A(KEYINPUT10), .B1(new_n430), .B2(new_n445), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n444), .A2(new_n446), .ZN(new_n447));
  OAI221_X1 g0247(.A(new_n430), .B1(new_n445), .B2(KEYINPUT10), .C1(new_n442), .C2(new_n443), .ZN(new_n448));
  NAND2_X1  g0248(.A1(new_n447), .A2(new_n448), .ZN(new_n449));
  NAND2_X1  g0249(.A1(new_n438), .A2(new_n441), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n417), .A2(new_n423), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n451), .A2(new_n247), .ZN(new_n452));
  NAND3_X1  g0252(.A1(new_n417), .A2(new_n382), .A3(new_n423), .ZN(new_n453));
  NAND3_X1  g0253(.A1(new_n450), .A2(new_n452), .A3(new_n453), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n415), .A2(G244), .ZN(new_n455));
  AND2_X1   g0255(.A1(new_n414), .A2(new_n455), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n377), .A2(G238), .ZN(new_n457));
  NAND3_X1  g0257(.A1(new_n252), .A2(G232), .A3(new_n369), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n420), .A2(G107), .ZN(new_n459));
  NAND3_X1  g0259(.A1(new_n457), .A2(new_n458), .A3(new_n459), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n460), .A2(new_n380), .ZN(new_n461));
  NAND3_X1  g0261(.A1(new_n456), .A2(new_n382), .A3(new_n461), .ZN(new_n462));
  INV_X1    g0262(.A(KEYINPUT70), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  NAND4_X1  g0264(.A1(new_n456), .A2(KEYINPUT70), .A3(new_n382), .A4(new_n461), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n456), .A2(new_n461), .ZN(new_n467));
  XNOR2_X1  g0267(.A(KEYINPUT15), .B(G87), .ZN(new_n468));
  INV_X1    g0268(.A(new_n468), .ZN(new_n469));
  NAND3_X1  g0269(.A1(new_n469), .A2(KEYINPUT69), .A3(new_n309), .ZN(new_n470));
  NAND2_X1  g0270(.A1(G20), .A2(G77), .ZN(new_n471));
  OAI211_X1 g0271(.A(new_n470), .B(new_n471), .C1(new_n312), .C2(new_n343), .ZN(new_n472));
  AOI21_X1  g0272(.A(KEYINPUT69), .B1(new_n469), .B2(new_n309), .ZN(new_n473));
  OAI21_X1  g0273(.A(new_n315), .B1(new_n472), .B2(new_n473), .ZN(new_n474));
  INV_X1    g0274(.A(G77), .ZN(new_n475));
  AOI21_X1  g0275(.A(new_n475), .B1(new_n264), .B2(G20), .ZN(new_n476));
  AOI22_X1  g0276(.A1(new_n326), .A2(new_n476), .B1(new_n475), .B2(new_n323), .ZN(new_n477));
  AOI22_X1  g0277(.A1(new_n467), .A2(new_n247), .B1(new_n474), .B2(new_n477), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n466), .A2(new_n478), .ZN(new_n479));
  AND2_X1   g0279(.A1(new_n474), .A2(new_n477), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n467), .A2(G200), .ZN(new_n481));
  INV_X1    g0281(.A(G190), .ZN(new_n482));
  OAI211_X1 g0282(.A(new_n480), .B(new_n481), .C1(new_n482), .C2(new_n467), .ZN(new_n483));
  NAND3_X1  g0283(.A1(new_n454), .A2(new_n479), .A3(new_n483), .ZN(new_n484));
  NOR3_X1   g0284(.A1(new_n413), .A2(new_n449), .A3(new_n484), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n342), .A2(new_n485), .ZN(new_n486));
  NOR2_X1   g0286(.A1(new_n335), .A2(new_n486), .ZN(new_n487));
  INV_X1    g0287(.A(KEYINPUT84), .ZN(new_n488));
  NOR2_X1   g0288(.A1(new_n312), .A2(new_n475), .ZN(new_n489));
  INV_X1    g0289(.A(new_n489), .ZN(new_n490));
  XNOR2_X1  g0290(.A(G97), .B(G107), .ZN(new_n491));
  INV_X1    g0291(.A(KEYINPUT6), .ZN(new_n492));
  INV_X1    g0292(.A(G107), .ZN(new_n493));
  INV_X1    g0293(.A(G97), .ZN(new_n494));
  NOR2_X1   g0294(.A1(new_n492), .A2(new_n494), .ZN(new_n495));
  AOI22_X1  g0295(.A1(new_n491), .A2(new_n492), .B1(new_n493), .B2(new_n495), .ZN(new_n496));
  OAI211_X1 g0296(.A(new_n488), .B(new_n490), .C1(new_n496), .C2(new_n214), .ZN(new_n497));
  AND2_X1   g0297(.A1(G97), .A2(G107), .ZN(new_n498));
  NOR2_X1   g0298(.A1(G97), .A2(G107), .ZN(new_n499));
  OAI21_X1  g0299(.A(new_n492), .B1(new_n498), .B2(new_n499), .ZN(new_n500));
  NAND3_X1  g0300(.A1(new_n493), .A2(KEYINPUT6), .A3(G97), .ZN(new_n501));
  AOI21_X1  g0301(.A(new_n214), .B1(new_n500), .B2(new_n501), .ZN(new_n502));
  OAI21_X1  g0302(.A(KEYINPUT84), .B1(new_n502), .B2(new_n489), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n361), .A2(new_n362), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n504), .A2(G107), .ZN(new_n505));
  NAND3_X1  g0305(.A1(new_n497), .A2(new_n503), .A3(new_n505), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n506), .A2(new_n315), .ZN(new_n507));
  AOI21_X1  g0307(.A(G97), .B1(new_n320), .B2(new_n321), .ZN(new_n508));
  INV_X1    g0308(.A(new_n315), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n264), .A2(G33), .ZN(new_n510));
  NAND3_X1  g0310(.A1(new_n322), .A2(new_n509), .A3(new_n510), .ZN(new_n511));
  AOI21_X1  g0311(.A(new_n508), .B1(new_n511), .B2(G97), .ZN(new_n512));
  INV_X1    g0312(.A(new_n512), .ZN(new_n513));
  AOI21_X1  g0313(.A(KEYINPUT87), .B1(new_n507), .B2(new_n513), .ZN(new_n514));
  INV_X1    g0314(.A(KEYINPUT87), .ZN(new_n515));
  AOI211_X1 g0315(.A(new_n515), .B(new_n512), .C1(new_n506), .C2(new_n315), .ZN(new_n516));
  NOR2_X1   g0316(.A1(new_n514), .A2(new_n516), .ZN(new_n517));
  XNOR2_X1  g0317(.A(KEYINPUT5), .B(G41), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n264), .A2(G45), .ZN(new_n519));
  INV_X1    g0319(.A(new_n519), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n518), .A2(new_n520), .ZN(new_n521));
  NAND3_X1  g0321(.A1(new_n521), .A2(G257), .A3(new_n261), .ZN(new_n522));
  OR2_X1    g0322(.A1(KEYINPUT5), .A2(G41), .ZN(new_n523));
  NAND2_X1  g0323(.A1(KEYINPUT5), .A2(G41), .ZN(new_n524));
  AOI21_X1  g0324(.A(new_n519), .B1(new_n523), .B2(new_n524), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n525), .A2(new_n275), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n522), .A2(new_n526), .ZN(new_n527));
  OAI211_X1 g0327(.A(G244), .B(new_n369), .C1(new_n370), .C2(new_n371), .ZN(new_n528));
  XNOR2_X1  g0328(.A(KEYINPUT85), .B(KEYINPUT4), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  NAND4_X1  g0330(.A1(new_n252), .A2(KEYINPUT4), .A3(G244), .A4(new_n369), .ZN(new_n531));
  NAND2_X1  g0331(.A1(G33), .A2(G283), .ZN(new_n532));
  OAI211_X1 g0332(.A(G250), .B(G1698), .C1(new_n370), .C2(new_n371), .ZN(new_n533));
  NAND4_X1  g0333(.A1(new_n530), .A2(new_n531), .A3(new_n532), .A4(new_n533), .ZN(new_n534));
  AOI21_X1  g0334(.A(new_n527), .B1(new_n380), .B2(new_n534), .ZN(new_n535));
  INV_X1    g0335(.A(KEYINPUT88), .ZN(new_n536));
  NAND3_X1  g0336(.A1(new_n535), .A2(new_n536), .A3(new_n382), .ZN(new_n537));
  INV_X1    g0337(.A(KEYINPUT4), .ZN(new_n538));
  OAI211_X1 g0338(.A(new_n532), .B(new_n533), .C1(new_n528), .C2(new_n538), .ZN(new_n539));
  AND2_X1   g0339(.A1(new_n528), .A2(new_n529), .ZN(new_n540));
  OAI21_X1  g0340(.A(new_n380), .B1(new_n539), .B2(new_n540), .ZN(new_n541));
  AND2_X1   g0341(.A1(new_n522), .A2(new_n526), .ZN(new_n542));
  NAND3_X1  g0342(.A1(new_n541), .A2(new_n542), .A3(new_n382), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n543), .A2(KEYINPUT88), .ZN(new_n544));
  AOI21_X1  g0344(.A(G169), .B1(new_n541), .B2(new_n542), .ZN(new_n545));
  OAI21_X1  g0345(.A(new_n537), .B1(new_n544), .B2(new_n545), .ZN(new_n546));
  AOI21_X1  g0346(.A(new_n512), .B1(new_n506), .B2(new_n315), .ZN(new_n547));
  NAND2_X1  g0347(.A1(KEYINPUT86), .A2(G200), .ZN(new_n548));
  NOR2_X1   g0348(.A1(new_n535), .A2(new_n548), .ZN(new_n549));
  OAI21_X1  g0349(.A(new_n482), .B1(new_n428), .B2(KEYINPUT86), .ZN(new_n550));
  AOI21_X1  g0350(.A(new_n549), .B1(new_n535), .B2(new_n550), .ZN(new_n551));
  AOI22_X1  g0351(.A1(new_n517), .A2(new_n546), .B1(new_n547), .B2(new_n551), .ZN(new_n552));
  OAI211_X1 g0352(.A(new_n214), .B(G87), .C1(new_n370), .C2(new_n371), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n553), .A2(KEYINPUT22), .ZN(new_n554));
  INV_X1    g0354(.A(KEYINPUT22), .ZN(new_n555));
  NAND4_X1  g0355(.A1(new_n252), .A2(new_n555), .A3(new_n214), .A4(G87), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n554), .A2(new_n556), .ZN(new_n557));
  INV_X1    g0357(.A(KEYINPUT24), .ZN(new_n558));
  INV_X1    g0358(.A(KEYINPUT23), .ZN(new_n559));
  OAI21_X1  g0359(.A(new_n559), .B1(new_n214), .B2(G107), .ZN(new_n560));
  NAND3_X1  g0360(.A1(new_n493), .A2(KEYINPUT23), .A3(G20), .ZN(new_n561));
  AOI22_X1  g0361(.A1(new_n560), .A2(new_n561), .B1(new_n309), .B2(G116), .ZN(new_n562));
  AND3_X1   g0362(.A1(new_n557), .A2(new_n558), .A3(new_n562), .ZN(new_n563));
  AOI21_X1  g0363(.A(new_n558), .B1(new_n557), .B2(new_n562), .ZN(new_n564));
  OAI21_X1  g0364(.A(new_n315), .B1(new_n563), .B2(new_n564), .ZN(new_n565));
  INV_X1    g0365(.A(KEYINPUT25), .ZN(new_n566));
  OAI21_X1  g0366(.A(new_n566), .B1(new_n322), .B2(G107), .ZN(new_n567));
  NAND3_X1  g0367(.A1(new_n323), .A2(KEYINPUT25), .A3(new_n493), .ZN(new_n568));
  INV_X1    g0368(.A(new_n511), .ZN(new_n569));
  AOI22_X1  g0369(.A1(new_n567), .A2(new_n568), .B1(new_n569), .B2(G107), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n565), .A2(new_n570), .ZN(new_n571));
  OAI211_X1 g0371(.A(G257), .B(G1698), .C1(new_n370), .C2(new_n371), .ZN(new_n572));
  OAI211_X1 g0372(.A(G250), .B(new_n369), .C1(new_n370), .C2(new_n371), .ZN(new_n573));
  INV_X1    g0373(.A(G294), .ZN(new_n574));
  OAI211_X1 g0374(.A(new_n572), .B(new_n573), .C1(new_n249), .C2(new_n574), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n575), .A2(new_n380), .ZN(new_n576));
  NOR2_X1   g0376(.A1(new_n525), .A2(new_n380), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n577), .A2(G264), .ZN(new_n578));
  NAND3_X1  g0378(.A1(new_n576), .A2(new_n526), .A3(new_n578), .ZN(new_n579));
  NOR2_X1   g0379(.A1(new_n579), .A2(new_n482), .ZN(new_n580));
  AOI22_X1  g0380(.A1(new_n575), .A2(new_n380), .B1(new_n577), .B2(G264), .ZN(new_n581));
  AOI21_X1  g0381(.A(new_n428), .B1(new_n581), .B2(new_n526), .ZN(new_n582));
  NOR3_X1   g0382(.A1(new_n571), .A2(new_n580), .A3(new_n582), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n579), .A2(G169), .ZN(new_n584));
  NAND3_X1  g0384(.A1(new_n581), .A2(G179), .A3(new_n526), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n584), .A2(new_n585), .ZN(new_n586));
  INV_X1    g0386(.A(KEYINPUT91), .ZN(new_n587));
  AOI22_X1  g0387(.A1(new_n586), .A2(new_n587), .B1(new_n565), .B2(new_n570), .ZN(new_n588));
  NAND3_X1  g0388(.A1(new_n584), .A2(KEYINPUT91), .A3(new_n585), .ZN(new_n589));
  AOI21_X1  g0389(.A(new_n583), .B1(new_n588), .B2(new_n589), .ZN(new_n590));
  INV_X1    g0390(.A(KEYINPUT21), .ZN(new_n591));
  AOI22_X1  g0391(.A1(new_n577), .A2(G270), .B1(new_n275), .B2(new_n525), .ZN(new_n592));
  OAI211_X1 g0392(.A(G264), .B(G1698), .C1(new_n370), .C2(new_n371), .ZN(new_n593));
  OAI211_X1 g0393(.A(G257), .B(new_n369), .C1(new_n370), .C2(new_n371), .ZN(new_n594));
  INV_X1    g0394(.A(G303), .ZN(new_n595));
  OAI211_X1 g0395(.A(new_n593), .B(new_n594), .C1(new_n595), .C2(new_n252), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n596), .A2(new_n380), .ZN(new_n597));
  AOI21_X1  g0397(.A(new_n247), .B1(new_n592), .B2(new_n597), .ZN(new_n598));
  INV_X1    g0398(.A(new_n598), .ZN(new_n599));
  INV_X1    g0399(.A(G116), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n323), .A2(new_n600), .ZN(new_n601));
  OAI21_X1  g0401(.A(new_n601), .B1(new_n511), .B2(new_n600), .ZN(new_n602));
  AOI22_X1  g0402(.A1(new_n314), .A2(new_n213), .B1(G20), .B2(new_n600), .ZN(new_n603));
  OAI211_X1 g0403(.A(new_n532), .B(new_n214), .C1(G33), .C2(new_n494), .ZN(new_n604));
  AND3_X1   g0404(.A1(new_n603), .A2(KEYINPUT20), .A3(new_n604), .ZN(new_n605));
  AOI21_X1  g0405(.A(KEYINPUT20), .B1(new_n603), .B2(new_n604), .ZN(new_n606));
  NOR2_X1   g0406(.A1(new_n605), .A2(new_n606), .ZN(new_n607));
  NOR2_X1   g0407(.A1(new_n602), .A2(new_n607), .ZN(new_n608));
  OAI21_X1  g0408(.A(new_n591), .B1(new_n599), .B2(new_n608), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n592), .A2(new_n597), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n610), .A2(G200), .ZN(new_n611));
  OAI211_X1 g0411(.A(new_n611), .B(new_n608), .C1(new_n482), .C2(new_n610), .ZN(new_n612));
  NAND3_X1  g0412(.A1(new_n592), .A2(G179), .A3(new_n597), .ZN(new_n613));
  INV_X1    g0413(.A(new_n613), .ZN(new_n614));
  OAI221_X1 g0414(.A(new_n601), .B1(new_n605), .B2(new_n606), .C1(new_n511), .C2(new_n600), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  NAND3_X1  g0416(.A1(new_n615), .A2(new_n598), .A3(KEYINPUT21), .ZN(new_n617));
  NAND4_X1  g0417(.A1(new_n609), .A2(new_n612), .A3(new_n616), .A4(new_n617), .ZN(new_n618));
  NAND3_X1  g0418(.A1(new_n214), .A2(G33), .A3(G97), .ZN(new_n619));
  INV_X1    g0419(.A(KEYINPUT19), .ZN(new_n620));
  AND3_X1   g0420(.A1(new_n619), .A2(KEYINPUT89), .A3(new_n620), .ZN(new_n621));
  AOI21_X1  g0421(.A(KEYINPUT89), .B1(new_n619), .B2(new_n620), .ZN(new_n622));
  NOR2_X1   g0422(.A1(new_n621), .A2(new_n622), .ZN(new_n623));
  OAI21_X1  g0423(.A(new_n214), .B1(new_n257), .B2(new_n620), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n499), .A2(new_n220), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  OAI211_X1 g0426(.A(new_n214), .B(G68), .C1(new_n370), .C2(new_n371), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  OAI21_X1  g0428(.A(new_n315), .B1(new_n623), .B2(new_n628), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n323), .A2(new_n468), .ZN(new_n630));
  NAND4_X1  g0430(.A1(new_n322), .A2(new_n509), .A3(new_n469), .A4(new_n510), .ZN(new_n631));
  NAND3_X1  g0431(.A1(new_n629), .A2(new_n630), .A3(new_n631), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n632), .A2(KEYINPUT90), .ZN(new_n633));
  OAI211_X1 g0433(.A(G244), .B(G1698), .C1(new_n370), .C2(new_n371), .ZN(new_n634));
  OAI211_X1 g0434(.A(G238), .B(new_n369), .C1(new_n370), .C2(new_n371), .ZN(new_n635));
  OAI211_X1 g0435(.A(new_n634), .B(new_n635), .C1(new_n249), .C2(new_n600), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n636), .A2(new_n380), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n519), .A2(G250), .ZN(new_n638));
  OAI22_X1  g0438(.A1(new_n270), .A2(new_n519), .B1(new_n380), .B2(new_n638), .ZN(new_n639));
  INV_X1    g0439(.A(new_n639), .ZN(new_n640));
  NAND3_X1  g0440(.A1(new_n637), .A2(G179), .A3(new_n640), .ZN(new_n641));
  AOI21_X1  g0441(.A(new_n639), .B1(new_n636), .B2(new_n380), .ZN(new_n642));
  OAI21_X1  g0442(.A(new_n641), .B1(new_n247), .B2(new_n642), .ZN(new_n643));
  INV_X1    g0443(.A(KEYINPUT90), .ZN(new_n644));
  NAND4_X1  g0444(.A1(new_n629), .A2(new_n644), .A3(new_n630), .A4(new_n631), .ZN(new_n645));
  NAND3_X1  g0445(.A1(new_n633), .A2(new_n643), .A3(new_n645), .ZN(new_n646));
  NAND4_X1  g0446(.A1(new_n322), .A2(new_n509), .A3(G87), .A4(new_n510), .ZN(new_n647));
  AND3_X1   g0447(.A1(new_n629), .A2(new_n630), .A3(new_n647), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n642), .A2(G190), .ZN(new_n649));
  OAI211_X1 g0449(.A(new_n648), .B(new_n649), .C1(new_n428), .C2(new_n642), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n646), .A2(new_n650), .ZN(new_n651));
  NOR2_X1   g0451(.A1(new_n618), .A2(new_n651), .ZN(new_n652));
  AND4_X1   g0452(.A1(new_n487), .A2(new_n552), .A3(new_n590), .A4(new_n652), .ZN(G372));
  INV_X1    g0453(.A(new_n454), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n393), .A2(new_n409), .ZN(new_n655));
  INV_X1    g0455(.A(new_n655), .ZN(new_n656));
  INV_X1    g0456(.A(new_n479), .ZN(new_n657));
  AOI22_X1  g0457(.A1(new_n308), .A2(new_n333), .B1(new_n338), .B2(new_n657), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n402), .A2(new_n412), .ZN(new_n659));
  OAI21_X1  g0459(.A(new_n656), .B1(new_n658), .B2(new_n659), .ZN(new_n660));
  INV_X1    g0460(.A(KEYINPUT94), .ZN(new_n661));
  XNOR2_X1  g0461(.A(new_n449), .B(new_n661), .ZN(new_n662));
  AOI21_X1  g0462(.A(new_n654), .B1(new_n660), .B2(new_n662), .ZN(new_n663));
  INV_X1    g0463(.A(KEYINPUT93), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n643), .A2(new_n632), .ZN(new_n665));
  INV_X1    g0465(.A(new_n665), .ZN(new_n666));
  AND2_X1   g0466(.A1(new_n646), .A2(new_n650), .ZN(new_n667));
  XOR2_X1   g0467(.A(KEYINPUT92), .B(KEYINPUT26), .Z(new_n668));
  INV_X1    g0468(.A(new_n668), .ZN(new_n669));
  NAND4_X1  g0469(.A1(new_n667), .A2(new_n546), .A3(new_n517), .A4(new_n669), .ZN(new_n670));
  INV_X1    g0470(.A(new_n547), .ZN(new_n671));
  NAND4_X1  g0471(.A1(new_n546), .A2(new_n671), .A3(new_n650), .A4(new_n665), .ZN(new_n672));
  INV_X1    g0472(.A(KEYINPUT26), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  AOI211_X1 g0474(.A(new_n664), .B(new_n666), .C1(new_n670), .C2(new_n674), .ZN(new_n675));
  NAND3_X1  g0475(.A1(new_n609), .A2(new_n616), .A3(new_n617), .ZN(new_n676));
  INV_X1    g0476(.A(new_n676), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n571), .A2(new_n586), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n650), .A2(new_n665), .ZN(new_n680));
  NOR2_X1   g0480(.A1(new_n583), .A2(new_n680), .ZN(new_n681));
  NAND3_X1  g0481(.A1(new_n679), .A2(new_n552), .A3(new_n681), .ZN(new_n682));
  AOI21_X1  g0482(.A(new_n666), .B1(new_n670), .B2(new_n674), .ZN(new_n683));
  OAI21_X1  g0483(.A(new_n682), .B1(new_n683), .B2(KEYINPUT93), .ZN(new_n684));
  OAI21_X1  g0484(.A(new_n487), .B1(new_n675), .B2(new_n684), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n663), .A2(new_n685), .ZN(new_n686));
  XOR2_X1   g0486(.A(new_n686), .B(KEYINPUT95), .Z(G369));
  NAND3_X1  g0487(.A1(new_n264), .A2(new_n214), .A3(G13), .ZN(new_n688));
  OR2_X1    g0488(.A1(new_n688), .A2(KEYINPUT27), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n688), .A2(KEYINPUT27), .ZN(new_n690));
  NAND3_X1  g0490(.A1(new_n689), .A2(G213), .A3(new_n690), .ZN(new_n691));
  INV_X1    g0491(.A(G343), .ZN(new_n692));
  NOR2_X1   g0492(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  INV_X1    g0493(.A(new_n693), .ZN(new_n694));
  NOR2_X1   g0494(.A1(new_n608), .A2(new_n694), .ZN(new_n695));
  OR2_X1    g0495(.A1(new_n618), .A2(new_n695), .ZN(new_n696));
  NAND2_X1  g0496(.A1(new_n676), .A2(new_n695), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n696), .A2(new_n697), .ZN(new_n698));
  NAND2_X1  g0498(.A1(new_n698), .A2(G330), .ZN(new_n699));
  INV_X1    g0499(.A(new_n571), .ZN(new_n700));
  OAI21_X1  g0500(.A(new_n590), .B1(new_n700), .B2(new_n694), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n586), .A2(new_n587), .ZN(new_n702));
  NAND3_X1  g0502(.A1(new_n702), .A2(new_n571), .A3(new_n589), .ZN(new_n703));
  INV_X1    g0503(.A(new_n703), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n704), .A2(new_n693), .ZN(new_n705));
  AOI21_X1  g0505(.A(new_n699), .B1(new_n701), .B2(new_n705), .ZN(new_n706));
  INV_X1    g0506(.A(new_n706), .ZN(new_n707));
  NOR2_X1   g0507(.A1(new_n678), .A2(new_n693), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n676), .A2(new_n694), .ZN(new_n709));
  INV_X1    g0509(.A(new_n709), .ZN(new_n710));
  AOI21_X1  g0510(.A(new_n708), .B1(new_n590), .B2(new_n710), .ZN(new_n711));
  NAND2_X1  g0511(.A1(new_n707), .A2(new_n711), .ZN(G399));
  INV_X1    g0512(.A(new_n207), .ZN(new_n713));
  NOR2_X1   g0513(.A1(new_n713), .A2(G41), .ZN(new_n714));
  INV_X1    g0514(.A(new_n714), .ZN(new_n715));
  NOR2_X1   g0515(.A1(new_n625), .A2(G116), .ZN(new_n716));
  NAND3_X1  g0516(.A1(new_n715), .A2(G1), .A3(new_n716), .ZN(new_n717));
  OAI21_X1  g0517(.A(new_n717), .B1(new_n211), .B2(new_n715), .ZN(new_n718));
  XNOR2_X1  g0518(.A(new_n718), .B(KEYINPUT96), .ZN(new_n719));
  XNOR2_X1  g0519(.A(new_n719), .B(KEYINPUT28), .ZN(new_n720));
  OAI21_X1  g0520(.A(new_n694), .B1(new_n684), .B2(new_n675), .ZN(new_n721));
  INV_X1    g0521(.A(KEYINPUT29), .ZN(new_n722));
  AOI21_X1  g0522(.A(KEYINPUT98), .B1(new_n721), .B2(new_n722), .ZN(new_n723));
  INV_X1    g0523(.A(new_n723), .ZN(new_n724));
  NAND3_X1  g0524(.A1(new_n721), .A2(KEYINPUT98), .A3(new_n722), .ZN(new_n725));
  INV_X1    g0525(.A(KEYINPUT100), .ZN(new_n726));
  OAI21_X1  g0526(.A(new_n726), .B1(new_n704), .B2(new_n676), .ZN(new_n727));
  NAND3_X1  g0527(.A1(new_n677), .A2(new_n703), .A3(KEYINPUT100), .ZN(new_n728));
  NAND4_X1  g0528(.A1(new_n727), .A2(new_n552), .A3(new_n681), .A4(new_n728), .ZN(new_n729));
  INV_X1    g0529(.A(new_n514), .ZN(new_n730));
  INV_X1    g0530(.A(new_n516), .ZN(new_n731));
  NAND3_X1  g0531(.A1(new_n730), .A2(new_n731), .A3(new_n546), .ZN(new_n732));
  OAI21_X1  g0532(.A(new_n668), .B1(new_n732), .B2(new_n651), .ZN(new_n733));
  AND2_X1   g0533(.A1(new_n546), .A2(new_n671), .ZN(new_n734));
  INV_X1    g0534(.A(new_n680), .ZN(new_n735));
  NAND4_X1  g0535(.A1(new_n734), .A2(KEYINPUT99), .A3(new_n735), .A4(KEYINPUT26), .ZN(new_n736));
  INV_X1    g0536(.A(KEYINPUT99), .ZN(new_n737));
  OAI21_X1  g0537(.A(new_n737), .B1(new_n672), .B2(new_n673), .ZN(new_n738));
  NAND3_X1  g0538(.A1(new_n733), .A2(new_n736), .A3(new_n738), .ZN(new_n739));
  NAND3_X1  g0539(.A1(new_n729), .A2(new_n739), .A3(new_n665), .ZN(new_n740));
  AND2_X1   g0540(.A1(new_n740), .A2(new_n694), .ZN(new_n741));
  AOI22_X1  g0541(.A1(new_n724), .A2(new_n725), .B1(KEYINPUT29), .B2(new_n741), .ZN(new_n742));
  AND2_X1   g0542(.A1(new_n642), .A2(new_n581), .ZN(new_n743));
  NAND4_X1  g0543(.A1(new_n743), .A2(new_n614), .A3(KEYINPUT30), .A4(new_n535), .ZN(new_n744));
  INV_X1    g0544(.A(new_n535), .ZN(new_n745));
  NOR2_X1   g0545(.A1(new_n642), .A2(G179), .ZN(new_n746));
  NAND4_X1  g0546(.A1(new_n745), .A2(new_n579), .A3(new_n610), .A4(new_n746), .ZN(new_n747));
  INV_X1    g0547(.A(KEYINPUT30), .ZN(new_n748));
  NAND4_X1  g0548(.A1(new_n581), .A2(new_n642), .A3(new_n541), .A4(new_n542), .ZN(new_n749));
  OAI21_X1  g0549(.A(new_n748), .B1(new_n749), .B2(new_n613), .ZN(new_n750));
  NAND3_X1  g0550(.A1(new_n744), .A2(new_n747), .A3(new_n750), .ZN(new_n751));
  AOI21_X1  g0551(.A(KEYINPUT31), .B1(new_n751), .B2(new_n693), .ZN(new_n752));
  NAND2_X1  g0552(.A1(new_n747), .A2(new_n750), .ZN(new_n753));
  NAND2_X1  g0553(.A1(new_n753), .A2(KEYINPUT97), .ZN(new_n754));
  INV_X1    g0554(.A(KEYINPUT97), .ZN(new_n755));
  NAND3_X1  g0555(.A1(new_n747), .A2(new_n750), .A3(new_n755), .ZN(new_n756));
  NAND3_X1  g0556(.A1(new_n754), .A2(new_n744), .A3(new_n756), .ZN(new_n757));
  AND2_X1   g0557(.A1(new_n693), .A2(KEYINPUT31), .ZN(new_n758));
  AOI21_X1  g0558(.A(new_n752), .B1(new_n757), .B2(new_n758), .ZN(new_n759));
  NAND4_X1  g0559(.A1(new_n590), .A2(new_n552), .A3(new_n652), .A4(new_n694), .ZN(new_n760));
  NAND2_X1  g0560(.A1(new_n759), .A2(new_n760), .ZN(new_n761));
  NAND2_X1  g0561(.A1(new_n761), .A2(G330), .ZN(new_n762));
  INV_X1    g0562(.A(new_n762), .ZN(new_n763));
  NOR2_X1   g0563(.A1(new_n742), .A2(new_n763), .ZN(new_n764));
  OAI21_X1  g0564(.A(new_n720), .B1(new_n764), .B2(G1), .ZN(G364));
  AND2_X1   g0565(.A1(new_n214), .A2(G13), .ZN(new_n766));
  AOI21_X1  g0566(.A(new_n264), .B1(new_n766), .B2(G45), .ZN(new_n767));
  INV_X1    g0567(.A(new_n767), .ZN(new_n768));
  NOR2_X1   g0568(.A1(new_n768), .A2(new_n714), .ZN(new_n769));
  OR2_X1    g0569(.A1(new_n698), .A2(G330), .ZN(new_n770));
  AOI21_X1  g0570(.A(new_n769), .B1(new_n770), .B2(new_n699), .ZN(new_n771));
  INV_X1    g0571(.A(new_n769), .ZN(new_n772));
  NOR2_X1   g0572(.A1(G13), .A2(G33), .ZN(new_n773));
  INV_X1    g0573(.A(new_n773), .ZN(new_n774));
  NOR2_X1   g0574(.A1(new_n774), .A2(G20), .ZN(new_n775));
  AOI21_X1  g0575(.A(new_n213), .B1(G20), .B2(new_n247), .ZN(new_n776));
  NOR2_X1   g0576(.A1(new_n775), .A2(new_n776), .ZN(new_n777));
  XOR2_X1   g0577(.A(new_n777), .B(KEYINPUT102), .Z(new_n778));
  INV_X1    g0578(.A(G45), .ZN(new_n779));
  NOR2_X1   g0579(.A1(new_n245), .A2(new_n779), .ZN(new_n780));
  INV_X1    g0580(.A(KEYINPUT101), .ZN(new_n781));
  NOR2_X1   g0581(.A1(new_n713), .A2(new_n252), .ZN(new_n782));
  INV_X1    g0582(.A(new_n782), .ZN(new_n783));
  AOI21_X1  g0583(.A(new_n783), .B1(new_n779), .B2(new_n212), .ZN(new_n784));
  AOI21_X1  g0584(.A(new_n780), .B1(new_n781), .B2(new_n784), .ZN(new_n785));
  OAI21_X1  g0585(.A(new_n785), .B1(new_n781), .B2(new_n784), .ZN(new_n786));
  NOR2_X1   g0586(.A1(new_n713), .A2(new_n420), .ZN(new_n787));
  AOI22_X1  g0587(.A1(new_n787), .A2(G355), .B1(new_n600), .B2(new_n713), .ZN(new_n788));
  AOI21_X1  g0588(.A(new_n778), .B1(new_n786), .B2(new_n788), .ZN(new_n789));
  NOR2_X1   g0589(.A1(new_n214), .A2(G179), .ZN(new_n790));
  NAND3_X1  g0590(.A1(new_n790), .A2(new_n482), .A3(G200), .ZN(new_n791));
  NOR2_X1   g0591(.A1(new_n791), .A2(new_n493), .ZN(new_n792));
  INV_X1    g0592(.A(new_n792), .ZN(new_n793));
  NOR2_X1   g0593(.A1(G179), .A2(G200), .ZN(new_n794));
  AOI21_X1  g0594(.A(new_n214), .B1(new_n794), .B2(G190), .ZN(new_n795));
  NOR2_X1   g0595(.A1(new_n214), .A2(G190), .ZN(new_n796));
  NAND2_X1  g0596(.A1(new_n796), .A2(new_n794), .ZN(new_n797));
  INV_X1    g0597(.A(G159), .ZN(new_n798));
  NOR2_X1   g0598(.A1(new_n797), .A2(new_n798), .ZN(new_n799));
  INV_X1    g0599(.A(KEYINPUT32), .ZN(new_n800));
  OAI221_X1 g0600(.A(new_n793), .B1(new_n494), .B2(new_n795), .C1(new_n799), .C2(new_n800), .ZN(new_n801));
  NOR2_X1   g0601(.A1(new_n382), .A2(G200), .ZN(new_n802));
  NAND2_X1  g0602(.A1(new_n796), .A2(new_n802), .ZN(new_n803));
  NAND3_X1  g0603(.A1(new_n802), .A2(G20), .A3(G190), .ZN(new_n804));
  OAI221_X1 g0604(.A(new_n252), .B1(new_n803), .B2(new_n475), .C1(new_n345), .C2(new_n804), .ZN(new_n805));
  NAND2_X1  g0605(.A1(new_n799), .A2(new_n800), .ZN(new_n806));
  NAND3_X1  g0606(.A1(new_n790), .A2(G190), .A3(G200), .ZN(new_n807));
  OAI21_X1  g0607(.A(new_n806), .B1(new_n220), .B2(new_n807), .ZN(new_n808));
  NOR3_X1   g0608(.A1(new_n801), .A2(new_n805), .A3(new_n808), .ZN(new_n809));
  NAND3_X1  g0609(.A1(G20), .A2(G179), .A3(G200), .ZN(new_n810));
  XNOR2_X1  g0610(.A(new_n810), .B(KEYINPUT103), .ZN(new_n811));
  NOR2_X1   g0611(.A1(new_n811), .A2(new_n482), .ZN(new_n812));
  INV_X1    g0612(.A(new_n812), .ZN(new_n813));
  NOR2_X1   g0613(.A1(new_n811), .A2(G190), .ZN(new_n814));
  INV_X1    g0614(.A(new_n814), .ZN(new_n815));
  OAI221_X1 g0615(.A(new_n809), .B1(new_n202), .B2(new_n813), .C1(new_n218), .C2(new_n815), .ZN(new_n816));
  OR2_X1    g0616(.A1(new_n816), .A2(KEYINPUT104), .ZN(new_n817));
  INV_X1    g0617(.A(new_n797), .ZN(new_n818));
  OR2_X1    g0618(.A1(new_n818), .A2(KEYINPUT105), .ZN(new_n819));
  NAND2_X1  g0619(.A1(new_n818), .A2(KEYINPUT105), .ZN(new_n820));
  NAND2_X1  g0620(.A1(new_n819), .A2(new_n820), .ZN(new_n821));
  INV_X1    g0621(.A(new_n821), .ZN(new_n822));
  NAND2_X1  g0622(.A1(new_n822), .A2(G329), .ZN(new_n823));
  INV_X1    g0623(.A(G283), .ZN(new_n824));
  OAI22_X1  g0624(.A1(new_n791), .A2(new_n824), .B1(new_n807), .B2(new_n595), .ZN(new_n825));
  INV_X1    g0625(.A(new_n795), .ZN(new_n826));
  AOI21_X1  g0626(.A(new_n825), .B1(G294), .B2(new_n826), .ZN(new_n827));
  INV_X1    g0627(.A(G322), .ZN(new_n828));
  OAI21_X1  g0628(.A(new_n420), .B1(new_n804), .B2(new_n828), .ZN(new_n829));
  INV_X1    g0629(.A(new_n803), .ZN(new_n830));
  AOI21_X1  g0630(.A(new_n829), .B1(G311), .B2(new_n830), .ZN(new_n831));
  XNOR2_X1  g0631(.A(KEYINPUT33), .B(G317), .ZN(new_n832));
  AOI22_X1  g0632(.A1(G326), .A2(new_n812), .B1(new_n814), .B2(new_n832), .ZN(new_n833));
  NAND4_X1  g0633(.A1(new_n823), .A2(new_n827), .A3(new_n831), .A4(new_n833), .ZN(new_n834));
  NAND2_X1  g0634(.A1(new_n816), .A2(KEYINPUT104), .ZN(new_n835));
  NAND3_X1  g0635(.A1(new_n817), .A2(new_n834), .A3(new_n835), .ZN(new_n836));
  AOI21_X1  g0636(.A(new_n789), .B1(new_n836), .B2(new_n776), .ZN(new_n837));
  NAND3_X1  g0637(.A1(new_n696), .A2(new_n697), .A3(new_n775), .ZN(new_n838));
  AOI21_X1  g0638(.A(new_n772), .B1(new_n837), .B2(new_n838), .ZN(new_n839));
  NOR2_X1   g0639(.A1(new_n771), .A2(new_n839), .ZN(new_n840));
  XNOR2_X1  g0640(.A(new_n840), .B(KEYINPUT106), .ZN(new_n841));
  INV_X1    g0641(.A(new_n841), .ZN(G396));
  OR2_X1    g0642(.A1(new_n480), .A2(new_n694), .ZN(new_n843));
  OR2_X1    g0643(.A1(new_n479), .A2(new_n843), .ZN(new_n844));
  NAND3_X1  g0644(.A1(new_n479), .A2(new_n843), .A3(new_n483), .ZN(new_n845));
  NAND2_X1  g0645(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  INV_X1    g0646(.A(new_n846), .ZN(new_n847));
  NAND2_X1  g0647(.A1(new_n721), .A2(new_n847), .ZN(new_n848));
  OAI211_X1 g0648(.A(new_n694), .B(new_n846), .C1(new_n684), .C2(new_n675), .ZN(new_n849));
  NAND2_X1  g0649(.A1(new_n848), .A2(new_n849), .ZN(new_n850));
  OAI21_X1  g0650(.A(new_n772), .B1(new_n850), .B2(new_n762), .ZN(new_n851));
  AOI22_X1  g0651(.A1(new_n851), .A2(KEYINPUT109), .B1(new_n762), .B2(new_n850), .ZN(new_n852));
  OAI21_X1  g0652(.A(new_n852), .B1(KEYINPUT109), .B2(new_n851), .ZN(new_n853));
  NOR2_X1   g0653(.A1(new_n776), .A2(new_n773), .ZN(new_n854));
  XOR2_X1   g0654(.A(new_n854), .B(KEYINPUT107), .Z(new_n855));
  INV_X1    g0655(.A(new_n855), .ZN(new_n856));
  AOI21_X1  g0656(.A(new_n772), .B1(new_n856), .B2(new_n475), .ZN(new_n857));
  INV_X1    g0657(.A(new_n804), .ZN(new_n858));
  AOI22_X1  g0658(.A1(new_n858), .A2(G143), .B1(new_n830), .B2(G159), .ZN(new_n859));
  INV_X1    g0659(.A(G150), .ZN(new_n860));
  OAI21_X1  g0660(.A(new_n859), .B1(new_n815), .B2(new_n860), .ZN(new_n861));
  AOI21_X1  g0661(.A(new_n861), .B1(G137), .B2(new_n812), .ZN(new_n862));
  XOR2_X1   g0662(.A(new_n862), .B(KEYINPUT34), .Z(new_n863));
  NOR2_X1   g0663(.A1(new_n791), .A2(new_n218), .ZN(new_n864));
  AOI21_X1  g0664(.A(new_n864), .B1(G58), .B2(new_n826), .ZN(new_n865));
  OAI211_X1 g0665(.A(new_n865), .B(new_n252), .C1(new_n202), .C2(new_n807), .ZN(new_n866));
  AOI21_X1  g0666(.A(new_n866), .B1(G132), .B2(new_n822), .ZN(new_n867));
  OAI22_X1  g0667(.A1(new_n804), .A2(new_n574), .B1(new_n795), .B2(new_n494), .ZN(new_n868));
  XOR2_X1   g0668(.A(new_n868), .B(KEYINPUT108), .Z(new_n869));
  AOI21_X1  g0669(.A(new_n252), .B1(new_n830), .B2(G116), .ZN(new_n870));
  INV_X1    g0670(.A(new_n791), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n871), .A2(G87), .ZN(new_n872));
  OAI211_X1 g0672(.A(new_n870), .B(new_n872), .C1(new_n493), .C2(new_n807), .ZN(new_n873));
  OAI22_X1  g0673(.A1(new_n824), .A2(new_n815), .B1(new_n813), .B2(new_n595), .ZN(new_n874));
  AOI211_X1 g0674(.A(new_n873), .B(new_n874), .C1(G311), .C2(new_n822), .ZN(new_n875));
  AOI22_X1  g0675(.A1(new_n863), .A2(new_n867), .B1(new_n869), .B2(new_n875), .ZN(new_n876));
  INV_X1    g0676(.A(new_n776), .ZN(new_n877));
  OAI221_X1 g0677(.A(new_n857), .B1(new_n876), .B2(new_n877), .C1(new_n774), .C2(new_n846), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n853), .A2(new_n878), .ZN(G384));
  INV_X1    g0679(.A(new_n496), .ZN(new_n880));
  OR2_X1    g0680(.A1(new_n880), .A2(KEYINPUT35), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n880), .A2(KEYINPUT35), .ZN(new_n882));
  NAND4_X1  g0682(.A1(new_n881), .A2(new_n882), .A3(G116), .A4(new_n215), .ZN(new_n883));
  XOR2_X1   g0683(.A(new_n883), .B(KEYINPUT36), .Z(new_n884));
  OR3_X1    g0684(.A1(new_n211), .A2(new_n475), .A3(new_n351), .ZN(new_n885));
  AOI211_X1 g0685(.A(new_n264), .B(G13), .C1(new_n885), .C2(new_n241), .ZN(new_n886));
  NOR2_X1   g0686(.A1(new_n884), .A2(new_n886), .ZN(new_n887));
  NAND3_X1  g0687(.A1(new_n289), .A2(G179), .A3(new_n297), .ZN(new_n888));
  OAI21_X1  g0688(.A(new_n888), .B1(new_n306), .B2(KEYINPUT14), .ZN(new_n889));
  OAI21_X1  g0689(.A(new_n304), .B1(new_n298), .B2(new_n299), .ZN(new_n890));
  NAND3_X1  g0690(.A1(new_n306), .A2(KEYINPUT79), .A3(KEYINPUT14), .ZN(new_n891));
  AOI21_X1  g0691(.A(new_n889), .B1(new_n890), .B2(new_n891), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n892), .A2(new_n342), .ZN(new_n893));
  NAND3_X1  g0693(.A1(new_n329), .A2(new_n331), .A3(new_n693), .ZN(new_n894));
  INV_X1    g0694(.A(new_n894), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n893), .A2(new_n895), .ZN(new_n896));
  XNOR2_X1  g0696(.A(new_n894), .B(KEYINPUT110), .ZN(new_n897));
  OAI211_X1 g0697(.A(new_n338), .B(new_n897), .C1(new_n892), .C2(new_n332), .ZN(new_n898));
  NOR2_X1   g0698(.A1(new_n479), .A2(new_n693), .ZN(new_n899));
  INV_X1    g0699(.A(new_n899), .ZN(new_n900));
  AOI22_X1  g0700(.A1(new_n896), .A2(new_n898), .B1(new_n849), .B2(new_n900), .ZN(new_n901));
  INV_X1    g0701(.A(KEYINPUT38), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n392), .A2(KEYINPUT113), .ZN(new_n903));
  INV_X1    g0703(.A(KEYINPUT37), .ZN(new_n904));
  INV_X1    g0704(.A(new_n691), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n368), .A2(new_n905), .ZN(new_n906));
  AND3_X1   g0706(.A1(new_n400), .A2(new_n904), .A3(new_n906), .ZN(new_n907));
  INV_X1    g0707(.A(KEYINPUT113), .ZN(new_n908));
  NAND3_X1  g0708(.A1(new_n407), .A2(new_n908), .A3(new_n368), .ZN(new_n909));
  AND3_X1   g0709(.A1(new_n903), .A2(new_n907), .A3(new_n909), .ZN(new_n910));
  INV_X1    g0710(.A(KEYINPUT112), .ZN(new_n911));
  INV_X1    g0711(.A(KEYINPUT111), .ZN(new_n912));
  NAND3_X1  g0712(.A1(new_n363), .A2(G68), .A3(new_n359), .ZN(new_n913));
  INV_X1    g0713(.A(new_n354), .ZN(new_n914));
  AOI21_X1  g0714(.A(KEYINPUT16), .B1(new_n913), .B2(new_n914), .ZN(new_n915));
  OAI21_X1  g0715(.A(new_n912), .B1(new_n915), .B2(new_n509), .ZN(new_n916));
  OAI211_X1 g0716(.A(KEYINPUT111), .B(new_n315), .C1(new_n395), .C2(KEYINPUT16), .ZN(new_n917));
  NAND3_X1  g0717(.A1(new_n916), .A2(new_n396), .A3(new_n917), .ZN(new_n918));
  AOI22_X1  g0718(.A1(new_n918), .A2(new_n349), .B1(new_n405), .B2(new_n406), .ZN(new_n919));
  OAI21_X1  g0719(.A(new_n911), .B1(new_n919), .B2(new_n411), .ZN(new_n920));
  INV_X1    g0720(.A(new_n349), .ZN(new_n921));
  OAI21_X1  g0721(.A(new_n315), .B1(new_n395), .B2(KEYINPUT16), .ZN(new_n922));
  AOI21_X1  g0722(.A(new_n364), .B1(new_n922), .B2(new_n912), .ZN(new_n923));
  AOI21_X1  g0723(.A(new_n921), .B1(new_n923), .B2(new_n917), .ZN(new_n924));
  NOR2_X1   g0724(.A1(new_n390), .A2(new_n391), .ZN(new_n925));
  OAI211_X1 g0725(.A(KEYINPUT112), .B(new_n400), .C1(new_n924), .C2(new_n925), .ZN(new_n926));
  NAND2_X1  g0726(.A1(new_n918), .A2(new_n349), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n927), .A2(new_n905), .ZN(new_n928));
  NAND3_X1  g0728(.A1(new_n920), .A2(new_n926), .A3(new_n928), .ZN(new_n929));
  AOI21_X1  g0729(.A(new_n910), .B1(new_n929), .B2(KEYINPUT37), .ZN(new_n930));
  NOR2_X1   g0730(.A1(new_n924), .A2(new_n691), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n413), .A2(new_n931), .ZN(new_n932));
  INV_X1    g0732(.A(new_n932), .ZN(new_n933));
  OAI21_X1  g0733(.A(new_n902), .B1(new_n930), .B2(new_n933), .ZN(new_n934));
  AOI21_X1  g0734(.A(new_n411), .B1(new_n927), .B2(new_n407), .ZN(new_n935));
  AOI21_X1  g0735(.A(new_n931), .B1(new_n935), .B2(KEYINPUT112), .ZN(new_n936));
  AOI21_X1  g0736(.A(new_n904), .B1(new_n936), .B2(new_n920), .ZN(new_n937));
  OAI211_X1 g0737(.A(KEYINPUT38), .B(new_n932), .C1(new_n937), .C2(new_n910), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n934), .A2(new_n938), .ZN(new_n939));
  AOI22_X1  g0739(.A1(new_n901), .A2(new_n939), .B1(new_n655), .B2(new_n691), .ZN(new_n940));
  NAND3_X1  g0740(.A1(new_n934), .A2(new_n938), .A3(KEYINPUT39), .ZN(new_n941));
  NOR2_X1   g0741(.A1(new_n334), .A2(new_n693), .ZN(new_n942));
  NAND3_X1  g0742(.A1(new_n903), .A2(new_n907), .A3(new_n909), .ZN(new_n943));
  INV_X1    g0743(.A(new_n906), .ZN(new_n944));
  AOI211_X1 g0744(.A(new_n411), .B(new_n944), .C1(new_n368), .C2(new_n407), .ZN(new_n945));
  OAI21_X1  g0745(.A(new_n943), .B1(new_n945), .B2(new_n904), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n413), .A2(new_n944), .ZN(new_n947));
  AOI21_X1  g0747(.A(KEYINPUT38), .B1(new_n946), .B2(new_n947), .ZN(new_n948));
  NOR2_X1   g0748(.A1(new_n930), .A2(new_n933), .ZN(new_n949));
  AOI21_X1  g0749(.A(new_n948), .B1(new_n949), .B2(KEYINPUT38), .ZN(new_n950));
  OAI211_X1 g0750(.A(new_n941), .B(new_n942), .C1(new_n950), .C2(KEYINPUT39), .ZN(new_n951));
  AND2_X1   g0751(.A1(new_n940), .A2(new_n951), .ZN(new_n952));
  NAND3_X1  g0752(.A1(new_n740), .A2(KEYINPUT29), .A3(new_n694), .ZN(new_n953));
  AND2_X1   g0753(.A1(new_n342), .A2(new_n485), .ZN(new_n954));
  AND3_X1   g0754(.A1(new_n953), .A2(new_n954), .A3(new_n334), .ZN(new_n955));
  AND3_X1   g0755(.A1(new_n721), .A2(KEYINPUT98), .A3(new_n722), .ZN(new_n956));
  OAI21_X1  g0756(.A(new_n955), .B1(new_n956), .B2(new_n723), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n957), .A2(new_n663), .ZN(new_n958));
  XNOR2_X1  g0758(.A(new_n952), .B(new_n958), .ZN(new_n959));
  INV_X1    g0759(.A(KEYINPUT40), .ZN(new_n960));
  AND2_X1   g0760(.A1(new_n934), .A2(new_n938), .ZN(new_n961));
  AND3_X1   g0761(.A1(new_n751), .A2(KEYINPUT31), .A3(new_n693), .ZN(new_n962));
  NOR2_X1   g0762(.A1(new_n962), .A2(new_n752), .ZN(new_n963));
  NAND2_X1  g0763(.A1(new_n760), .A2(new_n963), .ZN(new_n964));
  NAND2_X1  g0764(.A1(new_n964), .A2(new_n846), .ZN(new_n965));
  INV_X1    g0765(.A(new_n965), .ZN(new_n966));
  AOI21_X1  g0766(.A(new_n894), .B1(new_n892), .B2(new_n342), .ZN(new_n967));
  NAND2_X1  g0767(.A1(new_n897), .A2(new_n338), .ZN(new_n968));
  AOI21_X1  g0768(.A(new_n968), .B1(new_n308), .B2(new_n333), .ZN(new_n969));
  OAI21_X1  g0769(.A(new_n966), .B1(new_n967), .B2(new_n969), .ZN(new_n970));
  OAI21_X1  g0770(.A(new_n960), .B1(new_n961), .B2(new_n970), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n896), .A2(new_n898), .ZN(new_n972));
  NAND2_X1  g0772(.A1(new_n946), .A2(new_n947), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n973), .A2(new_n902), .ZN(new_n974));
  NAND2_X1  g0774(.A1(new_n938), .A2(new_n974), .ZN(new_n975));
  NAND4_X1  g0775(.A1(new_n972), .A2(new_n975), .A3(KEYINPUT40), .A4(new_n966), .ZN(new_n976));
  NAND4_X1  g0776(.A1(new_n971), .A2(new_n487), .A3(new_n964), .A4(new_n976), .ZN(new_n977));
  NAND2_X1  g0777(.A1(new_n977), .A2(G330), .ZN(new_n978));
  AOI22_X1  g0778(.A1(new_n971), .A2(new_n976), .B1(new_n487), .B2(new_n964), .ZN(new_n979));
  NOR2_X1   g0779(.A1(new_n978), .A2(new_n979), .ZN(new_n980));
  OAI22_X1  g0780(.A1(new_n959), .A2(new_n980), .B1(new_n264), .B2(new_n766), .ZN(new_n981));
  AND2_X1   g0781(.A1(new_n959), .A2(new_n980), .ZN(new_n982));
  OAI21_X1  g0782(.A(new_n887), .B1(new_n981), .B2(new_n982), .ZN(G367));
  OAI21_X1  g0783(.A(new_n552), .B1(new_n547), .B2(new_n694), .ZN(new_n984));
  NAND2_X1  g0784(.A1(new_n734), .A2(new_n693), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n984), .A2(new_n985), .ZN(new_n986));
  NAND2_X1  g0786(.A1(new_n986), .A2(new_n711), .ZN(new_n987));
  XNOR2_X1  g0787(.A(new_n987), .B(KEYINPUT45), .ZN(new_n988));
  AOI21_X1  g0788(.A(new_n988), .B1(KEYINPUT116), .B2(new_n706), .ZN(new_n989));
  NOR2_X1   g0789(.A1(new_n986), .A2(new_n711), .ZN(new_n990));
  XNOR2_X1  g0790(.A(new_n990), .B(KEYINPUT44), .ZN(new_n991));
  NAND2_X1  g0791(.A1(new_n989), .A2(new_n991), .ZN(new_n992));
  NOR2_X1   g0792(.A1(new_n706), .A2(KEYINPUT116), .ZN(new_n993));
  NAND2_X1  g0793(.A1(new_n992), .A2(new_n993), .ZN(new_n994));
  OAI211_X1 g0794(.A(new_n989), .B(new_n991), .C1(KEYINPUT116), .C2(new_n706), .ZN(new_n995));
  NAND2_X1  g0795(.A1(new_n994), .A2(new_n995), .ZN(new_n996));
  NAND3_X1  g0796(.A1(new_n701), .A2(new_n705), .A3(new_n709), .ZN(new_n997));
  NAND2_X1  g0797(.A1(new_n590), .A2(new_n710), .ZN(new_n998));
  NAND2_X1  g0798(.A1(new_n997), .A2(new_n998), .ZN(new_n999));
  XNOR2_X1  g0799(.A(new_n999), .B(new_n699), .ZN(new_n1000));
  INV_X1    g0800(.A(new_n1000), .ZN(new_n1001));
  NAND3_X1  g0801(.A1(new_n996), .A2(new_n764), .A3(new_n1001), .ZN(new_n1002));
  NAND2_X1  g0802(.A1(new_n1002), .A2(new_n764), .ZN(new_n1003));
  INV_X1    g0803(.A(new_n1003), .ZN(new_n1004));
  XOR2_X1   g0804(.A(new_n714), .B(KEYINPUT41), .Z(new_n1005));
  OAI21_X1  g0805(.A(new_n767), .B1(new_n1004), .B2(new_n1005), .ZN(new_n1006));
  INV_X1    g0806(.A(new_n986), .ZN(new_n1007));
  OR3_X1    g0807(.A1(new_n1007), .A2(KEYINPUT42), .A3(new_n998), .ZN(new_n1008));
  OAI21_X1  g0808(.A(KEYINPUT42), .B1(new_n1007), .B2(new_n998), .ZN(new_n1009));
  AOI22_X1  g0809(.A1(new_n986), .A2(new_n704), .B1(new_n546), .B2(new_n517), .ZN(new_n1010));
  OAI211_X1 g0810(.A(new_n1008), .B(new_n1009), .C1(new_n1010), .C2(new_n693), .ZN(new_n1011));
  NOR2_X1   g0811(.A1(new_n648), .A2(new_n694), .ZN(new_n1012));
  NAND2_X1  g0812(.A1(new_n666), .A2(new_n1012), .ZN(new_n1013));
  OAI21_X1  g0813(.A(new_n1013), .B1(new_n680), .B2(new_n1012), .ZN(new_n1014));
  NAND2_X1  g0814(.A1(new_n1014), .A2(KEYINPUT43), .ZN(new_n1015));
  NAND2_X1  g0815(.A1(new_n1011), .A2(new_n1015), .ZN(new_n1016));
  NAND2_X1  g0816(.A1(new_n1016), .A2(KEYINPUT114), .ZN(new_n1017));
  INV_X1    g0817(.A(KEYINPUT114), .ZN(new_n1018));
  NAND3_X1  g0818(.A1(new_n1011), .A2(new_n1018), .A3(new_n1015), .ZN(new_n1019));
  NAND2_X1  g0819(.A1(new_n1017), .A2(new_n1019), .ZN(new_n1020));
  NOR2_X1   g0820(.A1(new_n1014), .A2(KEYINPUT43), .ZN(new_n1021));
  INV_X1    g0821(.A(new_n1021), .ZN(new_n1022));
  NAND2_X1  g0822(.A1(new_n1020), .A2(new_n1022), .ZN(new_n1023));
  NOR2_X1   g0823(.A1(new_n707), .A2(new_n1007), .ZN(new_n1024));
  NAND3_X1  g0824(.A1(new_n1017), .A2(new_n1021), .A3(new_n1019), .ZN(new_n1025));
  NAND3_X1  g0825(.A1(new_n1023), .A2(new_n1024), .A3(new_n1025), .ZN(new_n1026));
  NAND2_X1  g0826(.A1(new_n1026), .A2(KEYINPUT115), .ZN(new_n1027));
  INV_X1    g0827(.A(KEYINPUT115), .ZN(new_n1028));
  NAND4_X1  g0828(.A1(new_n1023), .A2(new_n1028), .A3(new_n1024), .A4(new_n1025), .ZN(new_n1029));
  NAND2_X1  g0829(.A1(new_n1023), .A2(new_n1025), .ZN(new_n1030));
  INV_X1    g0830(.A(new_n1024), .ZN(new_n1031));
  NAND2_X1  g0831(.A1(new_n1030), .A2(new_n1031), .ZN(new_n1032));
  AND3_X1   g0832(.A1(new_n1027), .A2(new_n1029), .A3(new_n1032), .ZN(new_n1033));
  OAI211_X1 g0833(.A(new_n1013), .B(new_n775), .C1(new_n680), .C2(new_n1012), .ZN(new_n1034));
  INV_X1    g0834(.A(new_n778), .ZN(new_n1035));
  OAI21_X1  g0835(.A(new_n1035), .B1(new_n207), .B2(new_n468), .ZN(new_n1036));
  NOR2_X1   g0836(.A1(new_n236), .A2(new_n783), .ZN(new_n1037));
  OAI21_X1  g0837(.A(new_n769), .B1(new_n1036), .B2(new_n1037), .ZN(new_n1038));
  NOR2_X1   g0838(.A1(new_n795), .A2(new_n218), .ZN(new_n1039));
  NOR2_X1   g0839(.A1(new_n791), .A2(new_n475), .ZN(new_n1040));
  INV_X1    g0840(.A(new_n807), .ZN(new_n1041));
  AOI211_X1 g0841(.A(new_n1039), .B(new_n1040), .C1(G58), .C2(new_n1041), .ZN(new_n1042));
  AOI22_X1  g0842(.A1(G143), .A2(new_n812), .B1(new_n814), .B2(G159), .ZN(new_n1043));
  AOI21_X1  g0843(.A(new_n420), .B1(new_n858), .B2(G150), .ZN(new_n1044));
  XNOR2_X1  g0844(.A(KEYINPUT117), .B(G137), .ZN(new_n1045));
  INV_X1    g0845(.A(new_n1045), .ZN(new_n1046));
  AOI22_X1  g0846(.A1(G50), .A2(new_n830), .B1(new_n818), .B2(new_n1046), .ZN(new_n1047));
  NAND4_X1  g0847(.A1(new_n1042), .A2(new_n1043), .A3(new_n1044), .A4(new_n1047), .ZN(new_n1048));
  NAND2_X1  g0848(.A1(new_n1041), .A2(G116), .ZN(new_n1049));
  XNOR2_X1  g0849(.A(new_n1049), .B(KEYINPUT46), .ZN(new_n1050));
  AOI21_X1  g0850(.A(new_n252), .B1(new_n818), .B2(G317), .ZN(new_n1051));
  AOI22_X1  g0851(.A1(new_n858), .A2(G303), .B1(new_n830), .B2(G283), .ZN(new_n1052));
  NOR2_X1   g0852(.A1(new_n791), .A2(new_n494), .ZN(new_n1053));
  AOI21_X1  g0853(.A(new_n1053), .B1(G107), .B2(new_n826), .ZN(new_n1054));
  NAND4_X1  g0854(.A1(new_n1050), .A2(new_n1051), .A3(new_n1052), .A4(new_n1054), .ZN(new_n1055));
  INV_X1    g0855(.A(G311), .ZN(new_n1056));
  OAI22_X1  g0856(.A1(new_n574), .A2(new_n815), .B1(new_n813), .B2(new_n1056), .ZN(new_n1057));
  OAI21_X1  g0857(.A(new_n1048), .B1(new_n1055), .B2(new_n1057), .ZN(new_n1058));
  XNOR2_X1  g0858(.A(new_n1058), .B(KEYINPUT47), .ZN(new_n1059));
  AOI21_X1  g0859(.A(new_n1038), .B1(new_n1059), .B2(new_n776), .ZN(new_n1060));
  AOI22_X1  g0860(.A1(new_n1006), .A2(new_n1033), .B1(new_n1034), .B2(new_n1060), .ZN(new_n1061));
  INV_X1    g0861(.A(new_n1061), .ZN(G387));
  NAND2_X1  g0862(.A1(new_n764), .A2(new_n1001), .ZN(new_n1063));
  OAI21_X1  g0863(.A(new_n1000), .B1(new_n742), .B2(new_n763), .ZN(new_n1064));
  NAND3_X1  g0864(.A1(new_n1063), .A2(new_n714), .A3(new_n1064), .ZN(new_n1065));
  NAND3_X1  g0865(.A1(new_n701), .A2(new_n705), .A3(new_n775), .ZN(new_n1066));
  INV_X1    g0866(.A(new_n787), .ZN(new_n1067));
  OAI22_X1  g0867(.A1(new_n1067), .A2(new_n716), .B1(G107), .B2(new_n207), .ZN(new_n1068));
  OR2_X1    g0868(.A1(new_n233), .A2(new_n779), .ZN(new_n1069));
  INV_X1    g0869(.A(new_n716), .ZN(new_n1070));
  AOI211_X1 g0870(.A(G45), .B(new_n1070), .C1(G68), .C2(G77), .ZN(new_n1071));
  NOR2_X1   g0871(.A1(new_n343), .A2(G50), .ZN(new_n1072));
  XNOR2_X1  g0872(.A(new_n1072), .B(KEYINPUT50), .ZN(new_n1073));
  AOI21_X1  g0873(.A(new_n783), .B1(new_n1071), .B2(new_n1073), .ZN(new_n1074));
  AOI21_X1  g0874(.A(new_n1068), .B1(new_n1069), .B2(new_n1074), .ZN(new_n1075));
  OAI21_X1  g0875(.A(new_n769), .B1(new_n1075), .B2(new_n778), .ZN(new_n1076));
  AOI21_X1  g0876(.A(new_n420), .B1(new_n830), .B2(G68), .ZN(new_n1077));
  XOR2_X1   g0877(.A(KEYINPUT118), .B(G150), .Z(new_n1078));
  OAI221_X1 g0878(.A(new_n1077), .B1(new_n202), .B2(new_n804), .C1(new_n797), .C2(new_n1078), .ZN(new_n1079));
  NOR2_X1   g0879(.A1(new_n807), .A2(new_n475), .ZN(new_n1080));
  NOR2_X1   g0880(.A1(new_n795), .A2(new_n468), .ZN(new_n1081));
  NOR4_X1   g0881(.A1(new_n1079), .A2(new_n1053), .A3(new_n1080), .A4(new_n1081), .ZN(new_n1082));
  NAND2_X1  g0882(.A1(new_n812), .A2(G159), .ZN(new_n1083));
  XOR2_X1   g0883(.A(new_n1083), .B(KEYINPUT119), .Z(new_n1084));
  OAI211_X1 g0884(.A(new_n1082), .B(new_n1084), .C1(new_n347), .C2(new_n815), .ZN(new_n1085));
  OAI22_X1  g0885(.A1(new_n807), .A2(new_n574), .B1(new_n795), .B2(new_n824), .ZN(new_n1086));
  AOI22_X1  g0886(.A1(new_n858), .A2(G317), .B1(new_n830), .B2(G303), .ZN(new_n1087));
  OAI221_X1 g0887(.A(new_n1087), .B1(new_n815), .B2(new_n1056), .C1(new_n828), .C2(new_n813), .ZN(new_n1088));
  INV_X1    g0888(.A(KEYINPUT48), .ZN(new_n1089));
  AOI21_X1  g0889(.A(new_n1086), .B1(new_n1088), .B2(new_n1089), .ZN(new_n1090));
  OAI21_X1  g0890(.A(new_n1090), .B1(new_n1089), .B2(new_n1088), .ZN(new_n1091));
  XOR2_X1   g0891(.A(new_n1091), .B(KEYINPUT49), .Z(new_n1092));
  AOI21_X1  g0892(.A(new_n252), .B1(new_n818), .B2(G326), .ZN(new_n1093));
  OAI21_X1  g0893(.A(new_n1093), .B1(new_n600), .B2(new_n791), .ZN(new_n1094));
  OAI21_X1  g0894(.A(new_n1085), .B1(new_n1092), .B2(new_n1094), .ZN(new_n1095));
  AOI21_X1  g0895(.A(new_n1076), .B1(new_n1095), .B2(new_n776), .ZN(new_n1096));
  AOI22_X1  g0896(.A1(new_n1001), .A2(new_n768), .B1(new_n1066), .B2(new_n1096), .ZN(new_n1097));
  NAND2_X1  g0897(.A1(new_n1065), .A2(new_n1097), .ZN(G393));
  NAND2_X1  g0898(.A1(new_n996), .A2(new_n768), .ZN(new_n1099));
  NAND2_X1  g0899(.A1(new_n1007), .A2(new_n775), .ZN(new_n1100));
  XNOR2_X1  g0900(.A(new_n1100), .B(KEYINPUT120), .ZN(new_n1101));
  INV_X1    g0901(.A(new_n1101), .ZN(new_n1102));
  AOI21_X1  g0902(.A(new_n778), .B1(G97), .B2(new_n713), .ZN(new_n1103));
  NAND2_X1  g0903(.A1(new_n240), .A2(new_n782), .ZN(new_n1104));
  AOI21_X1  g0904(.A(new_n772), .B1(new_n1103), .B2(new_n1104), .ZN(new_n1105));
  AOI22_X1  g0905(.A1(new_n812), .A2(G317), .B1(G311), .B2(new_n858), .ZN(new_n1106));
  XOR2_X1   g0906(.A(new_n1106), .B(KEYINPUT52), .Z(new_n1107));
  OAI221_X1 g0907(.A(new_n420), .B1(new_n797), .B2(new_n828), .C1(new_n574), .C2(new_n803), .ZN(new_n1108));
  OAI221_X1 g0908(.A(new_n793), .B1(new_n600), .B2(new_n795), .C1(new_n824), .C2(new_n807), .ZN(new_n1109));
  AOI211_X1 g0909(.A(new_n1108), .B(new_n1109), .C1(G303), .C2(new_n814), .ZN(new_n1110));
  AOI21_X1  g0910(.A(new_n420), .B1(new_n818), .B2(G143), .ZN(new_n1111));
  OAI21_X1  g0911(.A(new_n1111), .B1(new_n343), .B2(new_n803), .ZN(new_n1112));
  OAI221_X1 g0912(.A(new_n872), .B1(new_n218), .B2(new_n807), .C1(new_n475), .C2(new_n795), .ZN(new_n1113));
  AOI211_X1 g0913(.A(new_n1112), .B(new_n1113), .C1(G50), .C2(new_n814), .ZN(new_n1114));
  AOI22_X1  g0914(.A1(new_n812), .A2(G150), .B1(G159), .B2(new_n858), .ZN(new_n1115));
  XOR2_X1   g0915(.A(new_n1115), .B(KEYINPUT51), .Z(new_n1116));
  AOI22_X1  g0916(.A1(new_n1107), .A2(new_n1110), .B1(new_n1114), .B2(new_n1116), .ZN(new_n1117));
  OAI211_X1 g0917(.A(new_n1102), .B(new_n1105), .C1(new_n877), .C2(new_n1117), .ZN(new_n1118));
  NAND2_X1  g0918(.A1(new_n1002), .A2(new_n714), .ZN(new_n1119));
  AOI21_X1  g0919(.A(new_n996), .B1(new_n764), .B2(new_n1001), .ZN(new_n1120));
  OAI211_X1 g0920(.A(new_n1099), .B(new_n1118), .C1(new_n1119), .C2(new_n1120), .ZN(G390));
  OAI211_X1 g0921(.A(G330), .B(new_n966), .C1(new_n967), .C2(new_n969), .ZN(new_n1122));
  INV_X1    g0922(.A(new_n941), .ZN(new_n1123));
  AOI21_X1  g0923(.A(KEYINPUT39), .B1(new_n938), .B2(new_n974), .ZN(new_n1124));
  OAI22_X1  g0924(.A1(new_n1123), .A2(new_n1124), .B1(new_n901), .B2(new_n942), .ZN(new_n1125));
  NOR2_X1   g0925(.A1(new_n950), .A2(new_n942), .ZN(new_n1126));
  NAND2_X1  g0926(.A1(new_n740), .A2(new_n694), .ZN(new_n1127));
  OAI21_X1  g0927(.A(new_n900), .B1(new_n1127), .B2(new_n847), .ZN(new_n1128));
  NAND2_X1  g0928(.A1(new_n972), .A2(new_n1128), .ZN(new_n1129));
  NAND2_X1  g0929(.A1(new_n1126), .A2(new_n1129), .ZN(new_n1130));
  AOI21_X1  g0930(.A(new_n1122), .B1(new_n1125), .B2(new_n1130), .ZN(new_n1131));
  OAI211_X1 g0931(.A(new_n763), .B(new_n846), .C1(new_n967), .C2(new_n969), .ZN(new_n1132));
  OR2_X1    g0932(.A1(new_n901), .A2(new_n942), .ZN(new_n1133));
  OAI21_X1  g0933(.A(new_n941), .B1(new_n950), .B2(KEYINPUT39), .ZN(new_n1134));
  AOI22_X1  g0934(.A1(new_n1133), .A2(new_n1134), .B1(new_n1129), .B2(new_n1126), .ZN(new_n1135));
  AOI21_X1  g0935(.A(new_n1131), .B1(new_n1132), .B2(new_n1135), .ZN(new_n1136));
  NAND2_X1  g0936(.A1(new_n1136), .A2(new_n768), .ZN(new_n1137));
  NAND2_X1  g0937(.A1(new_n1134), .A2(new_n773), .ZN(new_n1138));
  NOR2_X1   g0938(.A1(new_n821), .A2(new_n574), .ZN(new_n1139));
  AOI21_X1  g0939(.A(new_n864), .B1(G87), .B2(new_n1041), .ZN(new_n1140));
  OAI21_X1  g0940(.A(new_n1140), .B1(new_n475), .B2(new_n795), .ZN(new_n1141));
  OAI221_X1 g0941(.A(new_n420), .B1(new_n803), .B2(new_n494), .C1(new_n600), .C2(new_n804), .ZN(new_n1142));
  NOR3_X1   g0942(.A1(new_n1139), .A2(new_n1141), .A3(new_n1142), .ZN(new_n1143));
  OAI221_X1 g0943(.A(new_n1143), .B1(new_n493), .B2(new_n815), .C1(new_n824), .C2(new_n813), .ZN(new_n1144));
  OR2_X1    g0944(.A1(new_n1078), .A2(new_n807), .ZN(new_n1145));
  AOI22_X1  g0945(.A1(new_n822), .A2(G125), .B1(KEYINPUT53), .B2(new_n1145), .ZN(new_n1146));
  OAI21_X1  g0946(.A(new_n1146), .B1(KEYINPUT53), .B2(new_n1145), .ZN(new_n1147));
  NAND2_X1  g0947(.A1(new_n812), .A2(G128), .ZN(new_n1148));
  XNOR2_X1  g0948(.A(KEYINPUT54), .B(G143), .ZN(new_n1149));
  OAI21_X1  g0949(.A(new_n252), .B1(new_n803), .B2(new_n1149), .ZN(new_n1150));
  AOI21_X1  g0950(.A(new_n1150), .B1(G132), .B2(new_n858), .ZN(new_n1151));
  NAND2_X1  g0951(.A1(new_n814), .A2(new_n1046), .ZN(new_n1152));
  AOI22_X1  g0952(.A1(new_n871), .A2(G50), .B1(new_n826), .B2(G159), .ZN(new_n1153));
  NAND4_X1  g0953(.A1(new_n1148), .A2(new_n1151), .A3(new_n1152), .A4(new_n1153), .ZN(new_n1154));
  OAI21_X1  g0954(.A(new_n1144), .B1(new_n1147), .B2(new_n1154), .ZN(new_n1155));
  NAND2_X1  g0955(.A1(new_n1155), .A2(new_n776), .ZN(new_n1156));
  AOI21_X1  g0956(.A(new_n772), .B1(new_n856), .B2(new_n347), .ZN(new_n1157));
  NAND3_X1  g0957(.A1(new_n1138), .A2(new_n1156), .A3(new_n1157), .ZN(new_n1158));
  INV_X1    g0958(.A(KEYINPUT122), .ZN(new_n1159));
  AOI21_X1  g0959(.A(new_n899), .B1(new_n741), .B2(new_n846), .ZN(new_n1160));
  AND2_X1   g0960(.A1(new_n1132), .A2(new_n1160), .ZN(new_n1161));
  NAND2_X1  g0961(.A1(new_n964), .A2(G330), .ZN(new_n1162));
  NAND2_X1  g0962(.A1(new_n1162), .A2(KEYINPUT121), .ZN(new_n1163));
  INV_X1    g0963(.A(KEYINPUT121), .ZN(new_n1164));
  NAND3_X1  g0964(.A1(new_n964), .A2(new_n1164), .A3(G330), .ZN(new_n1165));
  NAND3_X1  g0965(.A1(new_n1163), .A2(new_n846), .A3(new_n1165), .ZN(new_n1166));
  NAND3_X1  g0966(.A1(new_n1166), .A2(new_n896), .A3(new_n898), .ZN(new_n1167));
  NAND3_X1  g0967(.A1(new_n761), .A2(G330), .A3(new_n846), .ZN(new_n1168));
  NAND3_X1  g0968(.A1(new_n896), .A2(new_n898), .A3(new_n1168), .ZN(new_n1169));
  NAND2_X1  g0969(.A1(new_n1122), .A2(new_n1169), .ZN(new_n1170));
  NAND2_X1  g0970(.A1(new_n849), .A2(new_n900), .ZN(new_n1171));
  AOI22_X1  g0971(.A1(new_n1161), .A2(new_n1167), .B1(new_n1170), .B2(new_n1171), .ZN(new_n1172));
  NAND3_X1  g0972(.A1(new_n487), .A2(G330), .A3(new_n964), .ZN(new_n1173));
  NAND3_X1  g0973(.A1(new_n957), .A2(new_n663), .A3(new_n1173), .ZN(new_n1174));
  OAI21_X1  g0974(.A(new_n1159), .B1(new_n1172), .B2(new_n1174), .ZN(new_n1175));
  AND3_X1   g0975(.A1(new_n957), .A2(new_n663), .A3(new_n1173), .ZN(new_n1176));
  NAND2_X1  g0976(.A1(new_n1170), .A2(new_n1171), .ZN(new_n1177));
  NAND3_X1  g0977(.A1(new_n1167), .A2(new_n1132), .A3(new_n1160), .ZN(new_n1178));
  NAND2_X1  g0978(.A1(new_n1177), .A2(new_n1178), .ZN(new_n1179));
  NAND3_X1  g0979(.A1(new_n1176), .A2(new_n1179), .A3(KEYINPUT122), .ZN(new_n1180));
  NAND2_X1  g0980(.A1(new_n1175), .A2(new_n1180), .ZN(new_n1181));
  OAI21_X1  g0981(.A(new_n714), .B1(new_n1181), .B2(new_n1136), .ZN(new_n1182));
  NAND3_X1  g0982(.A1(new_n1125), .A2(new_n1132), .A3(new_n1130), .ZN(new_n1183));
  OAI21_X1  g0983(.A(new_n1183), .B1(new_n1135), .B2(new_n1122), .ZN(new_n1184));
  AOI21_X1  g0984(.A(new_n1184), .B1(new_n1175), .B2(new_n1180), .ZN(new_n1185));
  OAI211_X1 g0985(.A(new_n1137), .B(new_n1158), .C1(new_n1182), .C2(new_n1185), .ZN(G378));
  XNOR2_X1  g0986(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1187));
  INV_X1    g0987(.A(new_n1187), .ZN(new_n1188));
  NAND2_X1  g0988(.A1(new_n450), .A2(new_n905), .ZN(new_n1189));
  AOI21_X1  g0989(.A(new_n1189), .B1(new_n662), .B2(new_n454), .ZN(new_n1190));
  NOR2_X1   g0990(.A1(new_n449), .A2(new_n661), .ZN(new_n1191));
  AOI21_X1  g0991(.A(KEYINPUT94), .B1(new_n447), .B2(new_n448), .ZN(new_n1192));
  OAI211_X1 g0992(.A(new_n454), .B(new_n1189), .C1(new_n1191), .C2(new_n1192), .ZN(new_n1193));
  INV_X1    g0993(.A(new_n1193), .ZN(new_n1194));
  OAI21_X1  g0994(.A(new_n1188), .B1(new_n1190), .B2(new_n1194), .ZN(new_n1195));
  NOR2_X1   g0995(.A1(new_n1191), .A2(new_n1192), .ZN(new_n1196));
  OAI211_X1 g0996(.A(new_n450), .B(new_n905), .C1(new_n1196), .C2(new_n654), .ZN(new_n1197));
  NAND3_X1  g0997(.A1(new_n1197), .A2(new_n1193), .A3(new_n1187), .ZN(new_n1198));
  NAND2_X1  g0998(.A1(new_n1195), .A2(new_n1198), .ZN(new_n1199));
  INV_X1    g0999(.A(new_n1199), .ZN(new_n1200));
  AOI21_X1  g1000(.A(new_n965), .B1(new_n896), .B2(new_n898), .ZN(new_n1201));
  AOI21_X1  g1001(.A(KEYINPUT40), .B1(new_n1201), .B2(new_n939), .ZN(new_n1202));
  OAI211_X1 g1002(.A(KEYINPUT40), .B(new_n966), .C1(new_n967), .C2(new_n969), .ZN(new_n1203));
  OAI21_X1  g1003(.A(G330), .B1(new_n1203), .B2(new_n950), .ZN(new_n1204));
  OAI21_X1  g1004(.A(new_n1200), .B1(new_n1202), .B2(new_n1204), .ZN(new_n1205));
  NAND4_X1  g1005(.A1(new_n971), .A2(G330), .A3(new_n976), .A4(new_n1199), .ZN(new_n1206));
  NAND2_X1  g1006(.A1(new_n1205), .A2(new_n1206), .ZN(new_n1207));
  NAND2_X1  g1007(.A1(new_n940), .A2(new_n951), .ZN(new_n1208));
  NAND2_X1  g1008(.A1(new_n1207), .A2(new_n1208), .ZN(new_n1209));
  NAND3_X1  g1009(.A1(new_n952), .A2(new_n1205), .A3(new_n1206), .ZN(new_n1210));
  AOI21_X1  g1010(.A(new_n767), .B1(new_n1209), .B2(new_n1210), .ZN(new_n1211));
  NOR2_X1   g1011(.A1(new_n252), .A2(G41), .ZN(new_n1212));
  OAI221_X1 g1012(.A(new_n1212), .B1(new_n493), .B2(new_n804), .C1(new_n468), .C2(new_n803), .ZN(new_n1213));
  AOI21_X1  g1013(.A(new_n1213), .B1(new_n822), .B2(G283), .ZN(new_n1214));
  AOI211_X1 g1014(.A(new_n1039), .B(new_n1080), .C1(G58), .C2(new_n871), .ZN(new_n1215));
  AOI22_X1  g1015(.A1(G97), .A2(new_n814), .B1(new_n812), .B2(G116), .ZN(new_n1216));
  NAND3_X1  g1016(.A1(new_n1214), .A2(new_n1215), .A3(new_n1216), .ZN(new_n1217));
  INV_X1    g1017(.A(KEYINPUT58), .ZN(new_n1218));
  INV_X1    g1018(.A(new_n1212), .ZN(new_n1219));
  INV_X1    g1019(.A(G41), .ZN(new_n1220));
  AOI21_X1  g1020(.A(G50), .B1(new_n249), .B2(new_n1220), .ZN(new_n1221));
  AOI22_X1  g1021(.A1(new_n1217), .A2(new_n1218), .B1(new_n1219), .B2(new_n1221), .ZN(new_n1222));
  AOI211_X1 g1022(.A(G33), .B(G41), .C1(new_n818), .C2(G124), .ZN(new_n1223));
  NAND2_X1  g1023(.A1(new_n814), .A2(G132), .ZN(new_n1224));
  AOI22_X1  g1024(.A1(new_n858), .A2(G128), .B1(new_n830), .B2(G137), .ZN(new_n1225));
  OAI211_X1 g1025(.A(new_n1224), .B(new_n1225), .C1(new_n807), .C2(new_n1149), .ZN(new_n1226));
  AOI22_X1  g1026(.A1(new_n812), .A2(G125), .B1(G150), .B2(new_n826), .ZN(new_n1227));
  OR2_X1    g1027(.A1(new_n1227), .A2(KEYINPUT123), .ZN(new_n1228));
  NAND2_X1  g1028(.A1(new_n1227), .A2(KEYINPUT123), .ZN(new_n1229));
  AOI21_X1  g1029(.A(new_n1226), .B1(new_n1228), .B2(new_n1229), .ZN(new_n1230));
  INV_X1    g1030(.A(KEYINPUT59), .ZN(new_n1231));
  OAI221_X1 g1031(.A(new_n1223), .B1(new_n798), .B2(new_n791), .C1(new_n1230), .C2(new_n1231), .ZN(new_n1232));
  AND2_X1   g1032(.A1(new_n1230), .A2(new_n1231), .ZN(new_n1233));
  OAI221_X1 g1033(.A(new_n1222), .B1(new_n1218), .B2(new_n1217), .C1(new_n1232), .C2(new_n1233), .ZN(new_n1234));
  NAND2_X1  g1034(.A1(new_n1234), .A2(new_n776), .ZN(new_n1235));
  AOI21_X1  g1035(.A(new_n772), .B1(new_n202), .B2(new_n854), .ZN(new_n1236));
  OAI211_X1 g1036(.A(new_n1235), .B(new_n1236), .C1(new_n1199), .C2(new_n774), .ZN(new_n1237));
  INV_X1    g1037(.A(new_n1237), .ZN(new_n1238));
  OAI21_X1  g1038(.A(KEYINPUT124), .B1(new_n1211), .B2(new_n1238), .ZN(new_n1239));
  AND3_X1   g1039(.A1(new_n952), .A2(new_n1205), .A3(new_n1206), .ZN(new_n1240));
  AOI22_X1  g1040(.A1(new_n1205), .A2(new_n1206), .B1(new_n951), .B2(new_n940), .ZN(new_n1241));
  OAI21_X1  g1041(.A(new_n768), .B1(new_n1240), .B2(new_n1241), .ZN(new_n1242));
  INV_X1    g1042(.A(KEYINPUT124), .ZN(new_n1243));
  NAND3_X1  g1043(.A1(new_n1242), .A2(new_n1243), .A3(new_n1237), .ZN(new_n1244));
  NAND2_X1  g1044(.A1(new_n1239), .A2(new_n1244), .ZN(new_n1245));
  NOR3_X1   g1045(.A1(new_n1172), .A2(new_n1159), .A3(new_n1174), .ZN(new_n1246));
  AOI21_X1  g1046(.A(KEYINPUT122), .B1(new_n1176), .B2(new_n1179), .ZN(new_n1247));
  NOR2_X1   g1047(.A1(new_n1246), .A2(new_n1247), .ZN(new_n1248));
  OAI21_X1  g1048(.A(new_n1176), .B1(new_n1248), .B2(new_n1184), .ZN(new_n1249));
  NAND2_X1  g1049(.A1(new_n1209), .A2(new_n1210), .ZN(new_n1250));
  AOI21_X1  g1050(.A(KEYINPUT57), .B1(new_n1249), .B2(new_n1250), .ZN(new_n1251));
  AOI21_X1  g1051(.A(new_n1174), .B1(new_n1181), .B2(new_n1136), .ZN(new_n1252));
  OAI21_X1  g1052(.A(KEYINPUT57), .B1(new_n1240), .B2(new_n1241), .ZN(new_n1253));
  OAI21_X1  g1053(.A(new_n714), .B1(new_n1252), .B2(new_n1253), .ZN(new_n1254));
  OAI21_X1  g1054(.A(new_n1245), .B1(new_n1251), .B2(new_n1254), .ZN(new_n1255));
  INV_X1    g1055(.A(KEYINPUT125), .ZN(new_n1256));
  AND2_X1   g1056(.A1(new_n1255), .A2(new_n1256), .ZN(new_n1257));
  NOR2_X1   g1057(.A1(new_n1255), .A2(new_n1256), .ZN(new_n1258));
  NOR2_X1   g1058(.A1(new_n1257), .A2(new_n1258), .ZN(G375));
  NAND2_X1  g1059(.A1(new_n1172), .A2(new_n1174), .ZN(new_n1260));
  NAND3_X1  g1060(.A1(new_n1175), .A2(new_n1180), .A3(new_n1260), .ZN(new_n1261));
  INV_X1    g1061(.A(new_n1261), .ZN(new_n1262));
  INV_X1    g1062(.A(new_n1005), .ZN(new_n1263));
  NAND2_X1  g1063(.A1(new_n1262), .A2(new_n1263), .ZN(new_n1264));
  NAND2_X1  g1064(.A1(new_n822), .A2(G303), .ZN(new_n1265));
  AOI211_X1 g1065(.A(new_n1081), .B(new_n1040), .C1(G97), .C2(new_n1041), .ZN(new_n1266));
  OAI21_X1  g1066(.A(new_n420), .B1(new_n804), .B2(new_n824), .ZN(new_n1267));
  AOI21_X1  g1067(.A(new_n1267), .B1(G107), .B2(new_n830), .ZN(new_n1268));
  AOI22_X1  g1068(.A1(G116), .A2(new_n814), .B1(new_n812), .B2(G294), .ZN(new_n1269));
  NAND4_X1  g1069(.A1(new_n1265), .A2(new_n1266), .A3(new_n1268), .A4(new_n1269), .ZN(new_n1270));
  NAND2_X1  g1070(.A1(new_n812), .A2(G132), .ZN(new_n1271));
  OAI221_X1 g1071(.A(new_n1271), .B1(new_n804), .B2(new_n1045), .C1(new_n815), .C2(new_n1149), .ZN(new_n1272));
  INV_X1    g1072(.A(KEYINPUT126), .ZN(new_n1273));
  NAND2_X1  g1073(.A1(new_n1272), .A2(new_n1273), .ZN(new_n1274));
  NAND2_X1  g1074(.A1(new_n822), .A2(G128), .ZN(new_n1275));
  OAI21_X1  g1075(.A(new_n252), .B1(new_n803), .B2(new_n860), .ZN(new_n1276));
  OAI22_X1  g1076(.A1(new_n807), .A2(new_n798), .B1(new_n795), .B2(new_n202), .ZN(new_n1277));
  AOI211_X1 g1077(.A(new_n1276), .B(new_n1277), .C1(G58), .C2(new_n871), .ZN(new_n1278));
  NAND3_X1  g1078(.A1(new_n1274), .A2(new_n1275), .A3(new_n1278), .ZN(new_n1279));
  NOR2_X1   g1079(.A1(new_n1272), .A2(new_n1273), .ZN(new_n1280));
  OAI21_X1  g1080(.A(new_n1270), .B1(new_n1279), .B2(new_n1280), .ZN(new_n1281));
  NAND2_X1  g1081(.A1(new_n1281), .A2(new_n776), .ZN(new_n1282));
  AOI21_X1  g1082(.A(new_n772), .B1(new_n856), .B2(new_n218), .ZN(new_n1283));
  OAI211_X1 g1083(.A(new_n1282), .B(new_n1283), .C1(new_n972), .C2(new_n774), .ZN(new_n1284));
  OAI21_X1  g1084(.A(new_n1284), .B1(new_n1172), .B2(new_n767), .ZN(new_n1285));
  INV_X1    g1085(.A(new_n1285), .ZN(new_n1286));
  NAND2_X1  g1086(.A1(new_n1264), .A2(new_n1286), .ZN(G381));
  INV_X1    g1087(.A(G390), .ZN(new_n1288));
  NAND2_X1  g1088(.A1(new_n1137), .A2(new_n1158), .ZN(new_n1289));
  INV_X1    g1089(.A(new_n1182), .ZN(new_n1290));
  INV_X1    g1090(.A(new_n1185), .ZN(new_n1291));
  AOI21_X1  g1091(.A(new_n1289), .B1(new_n1290), .B2(new_n1291), .ZN(new_n1292));
  NAND3_X1  g1092(.A1(new_n1061), .A2(new_n1288), .A3(new_n1292), .ZN(new_n1293));
  NOR2_X1   g1093(.A1(G393), .A2(G396), .ZN(new_n1294));
  INV_X1    g1094(.A(new_n1294), .ZN(new_n1295));
  INV_X1    g1095(.A(KEYINPUT127), .ZN(new_n1296));
  NOR3_X1   g1096(.A1(new_n1295), .A2(new_n1296), .A3(G384), .ZN(new_n1297));
  INV_X1    g1097(.A(G384), .ZN(new_n1298));
  AOI21_X1  g1098(.A(KEYINPUT127), .B1(new_n1294), .B2(new_n1298), .ZN(new_n1299));
  NOR4_X1   g1099(.A1(new_n1293), .A2(G381), .A3(new_n1297), .A4(new_n1299), .ZN(new_n1300));
  OAI21_X1  g1100(.A(new_n1300), .B1(new_n1257), .B2(new_n1258), .ZN(G407));
  OAI21_X1  g1101(.A(new_n1292), .B1(new_n1257), .B2(new_n1258), .ZN(new_n1302));
  OAI211_X1 g1102(.A(G407), .B(G213), .C1(G343), .C2(new_n1302), .ZN(G409));
  INV_X1    g1103(.A(KEYINPUT61), .ZN(new_n1304));
  NAND2_X1  g1104(.A1(new_n692), .A2(G213), .ZN(new_n1305));
  INV_X1    g1105(.A(new_n1305), .ZN(new_n1306));
  OAI211_X1 g1106(.A(new_n1245), .B(G378), .C1(new_n1251), .C2(new_n1254), .ZN(new_n1307));
  OAI211_X1 g1107(.A(new_n1263), .B(new_n1250), .C1(new_n1185), .C2(new_n1174), .ZN(new_n1308));
  NOR2_X1   g1108(.A1(new_n1211), .A2(new_n1238), .ZN(new_n1309));
  NAND2_X1  g1109(.A1(new_n1308), .A2(new_n1309), .ZN(new_n1310));
  NAND2_X1  g1110(.A1(new_n1310), .A2(new_n1292), .ZN(new_n1311));
  AOI21_X1  g1111(.A(new_n1306), .B1(new_n1307), .B2(new_n1311), .ZN(new_n1312));
  NAND2_X1  g1112(.A1(new_n1306), .A2(G2897), .ZN(new_n1313));
  INV_X1    g1113(.A(new_n1313), .ZN(new_n1314));
  NOR2_X1   g1114(.A1(new_n1176), .A2(new_n1179), .ZN(new_n1315));
  OAI21_X1  g1115(.A(new_n714), .B1(new_n1315), .B2(KEYINPUT60), .ZN(new_n1316));
  INV_X1    g1116(.A(new_n1316), .ZN(new_n1317));
  INV_X1    g1117(.A(KEYINPUT60), .ZN(new_n1318));
  OAI21_X1  g1118(.A(new_n1317), .B1(new_n1262), .B2(new_n1318), .ZN(new_n1319));
  AOI21_X1  g1119(.A(G384), .B1(new_n1319), .B2(new_n1286), .ZN(new_n1320));
  AOI21_X1  g1120(.A(new_n1316), .B1(KEYINPUT60), .B2(new_n1261), .ZN(new_n1321));
  NOR3_X1   g1121(.A1(new_n1321), .A2(new_n1298), .A3(new_n1285), .ZN(new_n1322));
  OAI21_X1  g1122(.A(new_n1314), .B1(new_n1320), .B2(new_n1322), .ZN(new_n1323));
  NAND3_X1  g1123(.A1(new_n1319), .A2(G384), .A3(new_n1286), .ZN(new_n1324));
  OAI21_X1  g1124(.A(new_n1298), .B1(new_n1321), .B2(new_n1285), .ZN(new_n1325));
  NAND3_X1  g1125(.A1(new_n1324), .A2(new_n1325), .A3(new_n1313), .ZN(new_n1326));
  NAND2_X1  g1126(.A1(new_n1323), .A2(new_n1326), .ZN(new_n1327));
  OAI21_X1  g1127(.A(new_n1304), .B1(new_n1312), .B2(new_n1327), .ZN(new_n1328));
  INV_X1    g1128(.A(new_n1328), .ZN(new_n1329));
  NOR2_X1   g1129(.A1(new_n1320), .A2(new_n1322), .ZN(new_n1330));
  NAND2_X1  g1130(.A1(new_n1312), .A2(new_n1330), .ZN(new_n1331));
  INV_X1    g1131(.A(KEYINPUT63), .ZN(new_n1332));
  NAND2_X1  g1132(.A1(new_n1331), .A2(new_n1332), .ZN(new_n1333));
  AOI21_X1  g1133(.A(new_n841), .B1(new_n1065), .B2(new_n1097), .ZN(new_n1334));
  OAI21_X1  g1134(.A(new_n1288), .B1(new_n1294), .B2(new_n1334), .ZN(new_n1335));
  NOR2_X1   g1135(.A1(new_n1294), .A2(new_n1334), .ZN(new_n1336));
  NAND2_X1  g1136(.A1(new_n1336), .A2(G390), .ZN(new_n1337));
  AND3_X1   g1137(.A1(new_n1061), .A2(new_n1335), .A3(new_n1337), .ZN(new_n1338));
  AOI21_X1  g1138(.A(new_n1061), .B1(new_n1337), .B2(new_n1335), .ZN(new_n1339));
  NOR2_X1   g1139(.A1(new_n1338), .A2(new_n1339), .ZN(new_n1340));
  NAND3_X1  g1140(.A1(new_n1312), .A2(KEYINPUT63), .A3(new_n1330), .ZN(new_n1341));
  NAND4_X1  g1141(.A1(new_n1329), .A2(new_n1333), .A3(new_n1340), .A4(new_n1341), .ZN(new_n1342));
  INV_X1    g1142(.A(KEYINPUT62), .ZN(new_n1343));
  AND3_X1   g1143(.A1(new_n1312), .A2(new_n1343), .A3(new_n1330), .ZN(new_n1344));
  AOI21_X1  g1144(.A(new_n1343), .B1(new_n1312), .B2(new_n1330), .ZN(new_n1345));
  NOR3_X1   g1145(.A1(new_n1344), .A2(new_n1328), .A3(new_n1345), .ZN(new_n1346));
  OAI21_X1  g1146(.A(new_n1342), .B1(new_n1346), .B2(new_n1340), .ZN(G405));
  NAND2_X1  g1147(.A1(new_n1255), .A2(G378), .ZN(new_n1348));
  NAND2_X1  g1148(.A1(new_n1302), .A2(new_n1348), .ZN(new_n1349));
  OAI22_X1  g1149(.A1(new_n1338), .A2(new_n1339), .B1(new_n1320), .B2(new_n1322), .ZN(new_n1350));
  NAND2_X1  g1150(.A1(new_n1335), .A2(new_n1337), .ZN(new_n1351));
  NAND2_X1  g1151(.A1(new_n1351), .A2(G387), .ZN(new_n1352));
  NAND3_X1  g1152(.A1(new_n1061), .A2(new_n1335), .A3(new_n1337), .ZN(new_n1353));
  NAND3_X1  g1153(.A1(new_n1352), .A2(new_n1330), .A3(new_n1353), .ZN(new_n1354));
  NAND2_X1  g1154(.A1(new_n1350), .A2(new_n1354), .ZN(new_n1355));
  XNOR2_X1  g1155(.A(new_n1349), .B(new_n1355), .ZN(G402));
endmodule


