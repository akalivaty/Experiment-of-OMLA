//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 1 1 1 0 1 0 0 1 1 1 1 0 1 1 0 0 1 1 1 0 1 0 1 0 0 0 0 0 0 1 1 1 1 1 0 0 0 0 0 1 1 0 0 0 0 0 0 1 0 0 1 0 0 1 0 0 0 0 1 0 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:35:42 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n245, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1233, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1246, new_n1247,
    new_n1248, new_n1249, new_n1250, new_n1251, new_n1252, new_n1253,
    new_n1254, new_n1255, new_n1257, new_n1258, new_n1259, new_n1260,
    new_n1261, new_n1262, new_n1263, new_n1264, new_n1265, new_n1267,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1323,
    new_n1324, new_n1325, new_n1326, new_n1327, new_n1328, new_n1329,
    new_n1330, new_n1331, new_n1332, new_n1333, new_n1334, new_n1335,
    new_n1336, new_n1337, new_n1338;
  XNOR2_X1  g0000(.A(KEYINPUT64), .B(G50), .ZN(new_n201));
  INV_X1    g0001(.A(G58), .ZN(new_n202));
  INV_X1    g0002(.A(G68), .ZN(new_n203));
  NAND2_X1  g0003(.A1(new_n202), .A2(new_n203), .ZN(new_n204));
  NOR3_X1   g0004(.A1(new_n201), .A2(G77), .A3(new_n204), .ZN(G353));
  OAI21_X1  g0005(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0006(.A1(new_n204), .A2(G50), .ZN(new_n207));
  INV_X1    g0007(.A(G20), .ZN(new_n208));
  NAND2_X1  g0008(.A1(G1), .A2(G13), .ZN(new_n209));
  NOR3_X1   g0009(.A1(new_n207), .A2(new_n208), .A3(new_n209), .ZN(new_n210));
  NAND2_X1  g0010(.A1(G1), .A2(G20), .ZN(new_n211));
  INV_X1    g0011(.A(KEYINPUT1), .ZN(new_n212));
  XOR2_X1   g0012(.A(KEYINPUT65), .B(G238), .Z(new_n213));
  AOI22_X1  g0013(.A1(new_n213), .A2(G68), .B1(G77), .B2(G244), .ZN(new_n214));
  INV_X1    g0014(.A(G232), .ZN(new_n215));
  OAI21_X1  g0015(.A(new_n214), .B1(new_n202), .B2(new_n215), .ZN(new_n216));
  AOI21_X1  g0016(.A(new_n216), .B1(G107), .B2(G264), .ZN(new_n217));
  NAND2_X1  g0017(.A1(G116), .A2(G270), .ZN(new_n218));
  NAND2_X1  g0018(.A1(G97), .A2(G257), .ZN(new_n219));
  NAND2_X1  g0019(.A1(G50), .A2(G226), .ZN(new_n220));
  NAND4_X1  g0020(.A1(new_n217), .A2(new_n218), .A3(new_n219), .A4(new_n220), .ZN(new_n221));
  AND2_X1   g0021(.A1(G87), .A2(G250), .ZN(new_n222));
  OAI221_X1 g0022(.A(new_n211), .B1(KEYINPUT66), .B2(new_n212), .C1(new_n221), .C2(new_n222), .ZN(new_n223));
  NAND2_X1  g0023(.A1(new_n212), .A2(KEYINPUT66), .ZN(new_n224));
  XNOR2_X1  g0024(.A(new_n223), .B(new_n224), .ZN(new_n225));
  NOR2_X1   g0025(.A1(new_n211), .A2(G13), .ZN(new_n226));
  OAI211_X1 g0026(.A(new_n226), .B(G250), .C1(G257), .C2(G264), .ZN(new_n227));
  NAND2_X1  g0027(.A1(new_n227), .A2(KEYINPUT0), .ZN(new_n228));
  OR2_X1    g0028(.A1(new_n227), .A2(KEYINPUT0), .ZN(new_n229));
  AOI211_X1 g0029(.A(new_n210), .B(new_n225), .C1(new_n228), .C2(new_n229), .ZN(G361));
  XNOR2_X1  g0030(.A(G238), .B(G244), .ZN(new_n231));
  XNOR2_X1  g0031(.A(new_n231), .B(new_n215), .ZN(new_n232));
  XOR2_X1   g0032(.A(KEYINPUT2), .B(G226), .Z(new_n233));
  XNOR2_X1  g0033(.A(new_n232), .B(new_n233), .ZN(new_n234));
  XNOR2_X1  g0034(.A(G250), .B(G257), .ZN(new_n235));
  XNOR2_X1  g0035(.A(G264), .B(G270), .ZN(new_n236));
  XOR2_X1   g0036(.A(new_n235), .B(new_n236), .Z(new_n237));
  XNOR2_X1  g0037(.A(new_n234), .B(new_n237), .ZN(G358));
  XOR2_X1   g0038(.A(G68), .B(G77), .Z(new_n239));
  XNOR2_X1  g0039(.A(new_n239), .B(KEYINPUT67), .ZN(new_n240));
  XNOR2_X1  g0040(.A(G50), .B(G58), .ZN(new_n241));
  XOR2_X1   g0041(.A(new_n240), .B(new_n241), .Z(new_n242));
  XNOR2_X1  g0042(.A(G87), .B(G97), .ZN(new_n243));
  XNOR2_X1  g0043(.A(G107), .B(G116), .ZN(new_n244));
  XOR2_X1   g0044(.A(new_n243), .B(new_n244), .Z(new_n245));
  XOR2_X1   g0045(.A(new_n242), .B(new_n245), .Z(G351));
  NAND2_X1  g0046(.A1(G33), .A2(G41), .ZN(new_n247));
  NAND3_X1  g0047(.A1(new_n247), .A2(G1), .A3(G13), .ZN(new_n248));
  INV_X1    g0048(.A(G1), .ZN(new_n249));
  OAI21_X1  g0049(.A(new_n249), .B1(G41), .B2(G45), .ZN(new_n250));
  NAND2_X1  g0050(.A1(new_n248), .A2(new_n250), .ZN(new_n251));
  INV_X1    g0051(.A(G226), .ZN(new_n252));
  NOR2_X1   g0052(.A1(new_n251), .A2(new_n252), .ZN(new_n253));
  INV_X1    g0053(.A(G274), .ZN(new_n254));
  NOR2_X1   g0054(.A1(new_n250), .A2(new_n254), .ZN(new_n255));
  OAI21_X1  g0055(.A(KEYINPUT68), .B1(new_n253), .B2(new_n255), .ZN(new_n256));
  INV_X1    g0056(.A(KEYINPUT3), .ZN(new_n257));
  INV_X1    g0057(.A(G33), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n257), .A2(new_n258), .ZN(new_n259));
  NAND2_X1  g0059(.A1(KEYINPUT3), .A2(G33), .ZN(new_n260));
  NAND2_X1  g0060(.A1(new_n259), .A2(new_n260), .ZN(new_n261));
  NOR2_X1   g0061(.A1(G222), .A2(G1698), .ZN(new_n262));
  INV_X1    g0062(.A(G1698), .ZN(new_n263));
  NOR2_X1   g0063(.A1(new_n263), .A2(G223), .ZN(new_n264));
  OAI21_X1  g0064(.A(new_n261), .B1(new_n262), .B2(new_n264), .ZN(new_n265));
  AND2_X1   g0065(.A1(G33), .A2(G41), .ZN(new_n266));
  OAI21_X1  g0066(.A(KEYINPUT69), .B1(new_n266), .B2(new_n209), .ZN(new_n267));
  INV_X1    g0067(.A(KEYINPUT69), .ZN(new_n268));
  NAND4_X1  g0068(.A1(new_n247), .A2(new_n268), .A3(G1), .A4(G13), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n267), .A2(new_n269), .ZN(new_n270));
  OAI211_X1 g0070(.A(new_n265), .B(new_n270), .C1(G77), .C2(new_n261), .ZN(new_n271));
  INV_X1    g0071(.A(new_n255), .ZN(new_n272));
  INV_X1    g0072(.A(KEYINPUT68), .ZN(new_n273));
  OAI211_X1 g0073(.A(new_n272), .B(new_n273), .C1(new_n252), .C2(new_n251), .ZN(new_n274));
  NAND3_X1  g0074(.A1(new_n256), .A2(new_n271), .A3(new_n274), .ZN(new_n275));
  OR2_X1    g0075(.A1(new_n275), .A2(G179), .ZN(new_n276));
  OAI21_X1  g0076(.A(G20), .B1(new_n201), .B2(new_n204), .ZN(new_n277));
  INV_X1    g0077(.A(G150), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n208), .A2(new_n258), .ZN(new_n279));
  NAND2_X1  g0079(.A1(new_n208), .A2(G33), .ZN(new_n280));
  XNOR2_X1  g0080(.A(KEYINPUT8), .B(G58), .ZN(new_n281));
  OAI221_X1 g0081(.A(new_n277), .B1(new_n278), .B2(new_n279), .C1(new_n280), .C2(new_n281), .ZN(new_n282));
  NAND3_X1  g0082(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n283), .A2(new_n209), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n282), .A2(new_n284), .ZN(new_n285));
  NAND2_X1  g0085(.A1(new_n249), .A2(G20), .ZN(new_n286));
  INV_X1    g0086(.A(new_n286), .ZN(new_n287));
  NOR2_X1   g0087(.A1(new_n287), .A2(new_n284), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n288), .A2(G50), .ZN(new_n289));
  NAND3_X1  g0089(.A1(new_n249), .A2(G13), .A3(G20), .ZN(new_n290));
  INV_X1    g0090(.A(new_n290), .ZN(new_n291));
  INV_X1    g0091(.A(G50), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n291), .A2(new_n292), .ZN(new_n293));
  NAND3_X1  g0093(.A1(new_n285), .A2(new_n289), .A3(new_n293), .ZN(new_n294));
  INV_X1    g0094(.A(G169), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n275), .A2(new_n295), .ZN(new_n296));
  NAND3_X1  g0096(.A1(new_n276), .A2(new_n294), .A3(new_n296), .ZN(new_n297));
  INV_X1    g0097(.A(KEYINPUT9), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n294), .A2(new_n298), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n275), .A2(G200), .ZN(new_n300));
  NAND4_X1  g0100(.A1(new_n285), .A2(KEYINPUT9), .A3(new_n289), .A4(new_n293), .ZN(new_n301));
  INV_X1    g0101(.A(G190), .ZN(new_n302));
  OR2_X1    g0102(.A1(new_n275), .A2(new_n302), .ZN(new_n303));
  NAND4_X1  g0103(.A1(new_n299), .A2(new_n300), .A3(new_n301), .A4(new_n303), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n304), .A2(KEYINPUT10), .ZN(new_n305));
  INV_X1    g0105(.A(new_n305), .ZN(new_n306));
  NOR2_X1   g0106(.A1(new_n304), .A2(KEYINPUT10), .ZN(new_n307));
  OAI21_X1  g0107(.A(new_n297), .B1(new_n306), .B2(new_n307), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n281), .A2(new_n290), .ZN(new_n309));
  OAI21_X1  g0109(.A(new_n309), .B1(new_n288), .B2(new_n281), .ZN(new_n310));
  INV_X1    g0110(.A(new_n310), .ZN(new_n311));
  XNOR2_X1  g0111(.A(G58), .B(G68), .ZN(new_n312));
  INV_X1    g0112(.A(new_n279), .ZN(new_n313));
  AOI22_X1  g0113(.A1(G20), .A2(new_n312), .B1(new_n313), .B2(G159), .ZN(new_n314));
  NAND4_X1  g0114(.A1(new_n259), .A2(KEYINPUT7), .A3(new_n208), .A4(new_n260), .ZN(new_n315));
  INV_X1    g0115(.A(KEYINPUT74), .ZN(new_n316));
  NOR2_X1   g0116(.A1(new_n315), .A2(new_n316), .ZN(new_n317));
  AND2_X1   g0117(.A1(KEYINPUT3), .A2(G33), .ZN(new_n318));
  NOR2_X1   g0118(.A1(KEYINPUT3), .A2(G33), .ZN(new_n319));
  NOR3_X1   g0119(.A1(new_n318), .A2(new_n319), .A3(G20), .ZN(new_n320));
  XNOR2_X1  g0120(.A(KEYINPUT73), .B(KEYINPUT7), .ZN(new_n321));
  OAI21_X1  g0121(.A(KEYINPUT74), .B1(new_n320), .B2(new_n321), .ZN(new_n322));
  AOI21_X1  g0122(.A(new_n317), .B1(new_n322), .B2(new_n315), .ZN(new_n323));
  OAI21_X1  g0123(.A(new_n314), .B1(new_n323), .B2(new_n203), .ZN(new_n324));
  INV_X1    g0124(.A(KEYINPUT16), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n324), .A2(new_n325), .ZN(new_n326));
  INV_X1    g0126(.A(KEYINPUT7), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n327), .A2(KEYINPUT73), .ZN(new_n328));
  INV_X1    g0128(.A(KEYINPUT73), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n329), .A2(KEYINPUT7), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n328), .A2(new_n330), .ZN(new_n331));
  NOR2_X1   g0131(.A1(new_n318), .A2(new_n319), .ZN(new_n332));
  NAND3_X1  g0132(.A1(new_n331), .A2(new_n332), .A3(new_n208), .ZN(new_n333));
  NAND3_X1  g0133(.A1(new_n259), .A2(new_n208), .A3(new_n260), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n334), .A2(KEYINPUT7), .ZN(new_n335));
  NAND3_X1  g0135(.A1(new_n333), .A2(new_n335), .A3(G68), .ZN(new_n336));
  NAND3_X1  g0136(.A1(new_n336), .A2(KEYINPUT16), .A3(new_n314), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n337), .A2(new_n284), .ZN(new_n338));
  INV_X1    g0138(.A(new_n338), .ZN(new_n339));
  AOI21_X1  g0139(.A(new_n311), .B1(new_n326), .B2(new_n339), .ZN(new_n340));
  OR2_X1    g0140(.A1(G223), .A2(G1698), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n252), .A2(G1698), .ZN(new_n342));
  OAI211_X1 g0142(.A(new_n341), .B(new_n342), .C1(new_n318), .C2(new_n319), .ZN(new_n343));
  NAND2_X1  g0143(.A1(G33), .A2(G87), .ZN(new_n344));
  AOI22_X1  g0144(.A1(new_n343), .A2(new_n344), .B1(new_n267), .B2(new_n269), .ZN(new_n345));
  AND3_X1   g0145(.A1(new_n248), .A2(G232), .A3(new_n250), .ZN(new_n346));
  NOR3_X1   g0146(.A1(new_n345), .A2(new_n255), .A3(new_n346), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n347), .A2(G190), .ZN(new_n348));
  INV_X1    g0148(.A(G200), .ZN(new_n349));
  OR2_X1    g0149(.A1(new_n347), .A2(new_n349), .ZN(new_n350));
  NAND4_X1  g0150(.A1(new_n340), .A2(KEYINPUT17), .A3(new_n348), .A4(new_n350), .ZN(new_n351));
  INV_X1    g0151(.A(KEYINPUT75), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n343), .A2(new_n344), .ZN(new_n353));
  AOI21_X1  g0153(.A(new_n255), .B1(new_n353), .B2(new_n270), .ZN(new_n354));
  INV_X1    g0154(.A(new_n346), .ZN(new_n355));
  AOI21_X1  g0155(.A(new_n295), .B1(new_n354), .B2(new_n355), .ZN(new_n356));
  INV_X1    g0156(.A(G179), .ZN(new_n357));
  NOR4_X1   g0157(.A1(new_n345), .A2(new_n357), .A3(new_n346), .A4(new_n255), .ZN(new_n358));
  OAI21_X1  g0158(.A(new_n352), .B1(new_n356), .B2(new_n358), .ZN(new_n359));
  NAND3_X1  g0159(.A1(new_n354), .A2(G179), .A3(new_n355), .ZN(new_n360));
  OAI211_X1 g0160(.A(new_n360), .B(KEYINPUT75), .C1(new_n295), .C2(new_n347), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n359), .A2(new_n361), .ZN(new_n362));
  OAI21_X1  g0162(.A(KEYINPUT18), .B1(new_n340), .B2(new_n362), .ZN(new_n363));
  INV_X1    g0163(.A(new_n314), .ZN(new_n364));
  NAND3_X1  g0164(.A1(new_n320), .A2(KEYINPUT74), .A3(KEYINPUT7), .ZN(new_n365));
  AOI21_X1  g0165(.A(new_n316), .B1(new_n334), .B2(new_n331), .ZN(new_n366));
  INV_X1    g0166(.A(new_n315), .ZN(new_n367));
  OAI21_X1  g0167(.A(new_n365), .B1(new_n366), .B2(new_n367), .ZN(new_n368));
  AOI21_X1  g0168(.A(new_n364), .B1(new_n368), .B2(G68), .ZN(new_n369));
  OAI211_X1 g0169(.A(new_n284), .B(new_n337), .C1(new_n369), .C2(KEYINPUT16), .ZN(new_n370));
  NAND4_X1  g0170(.A1(new_n370), .A2(new_n348), .A3(new_n310), .A4(new_n350), .ZN(new_n371));
  INV_X1    g0171(.A(KEYINPUT17), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n371), .A2(new_n372), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n368), .A2(G68), .ZN(new_n374));
  AOI21_X1  g0174(.A(KEYINPUT16), .B1(new_n374), .B2(new_n314), .ZN(new_n375));
  OAI21_X1  g0175(.A(new_n310), .B1(new_n375), .B2(new_n338), .ZN(new_n376));
  INV_X1    g0176(.A(KEYINPUT18), .ZN(new_n377));
  NAND4_X1  g0177(.A1(new_n376), .A2(new_n377), .A3(new_n359), .A4(new_n361), .ZN(new_n378));
  NAND4_X1  g0178(.A1(new_n351), .A2(new_n363), .A3(new_n373), .A4(new_n378), .ZN(new_n379));
  NOR2_X1   g0179(.A1(new_n308), .A2(new_n379), .ZN(new_n380));
  NAND3_X1  g0180(.A1(new_n213), .A2(G1698), .A3(new_n261), .ZN(new_n381));
  OAI211_X1 g0181(.A(G232), .B(new_n263), .C1(new_n318), .C2(new_n319), .ZN(new_n382));
  INV_X1    g0182(.A(KEYINPUT70), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n382), .A2(new_n383), .ZN(new_n384));
  NAND4_X1  g0184(.A1(new_n261), .A2(KEYINPUT70), .A3(G232), .A4(new_n263), .ZN(new_n385));
  NAND2_X1  g0185(.A1(new_n332), .A2(G107), .ZN(new_n386));
  NAND4_X1  g0186(.A1(new_n381), .A2(new_n384), .A3(new_n385), .A4(new_n386), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n387), .A2(new_n270), .ZN(new_n388));
  INV_X1    g0188(.A(new_n251), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n389), .A2(G244), .ZN(new_n390));
  NAND3_X1  g0190(.A1(new_n388), .A2(new_n272), .A3(new_n390), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n391), .A2(G200), .ZN(new_n392));
  AOI21_X1  g0192(.A(new_n255), .B1(new_n387), .B2(new_n270), .ZN(new_n393));
  NAND3_X1  g0193(.A1(new_n393), .A2(G190), .A3(new_n390), .ZN(new_n394));
  NAND2_X1  g0194(.A1(G20), .A2(G77), .ZN(new_n395));
  XNOR2_X1  g0195(.A(KEYINPUT15), .B(G87), .ZN(new_n396));
  OAI221_X1 g0196(.A(new_n395), .B1(new_n281), .B2(new_n279), .C1(new_n280), .C2(new_n396), .ZN(new_n397));
  INV_X1    g0197(.A(G77), .ZN(new_n398));
  AOI22_X1  g0198(.A1(new_n397), .A2(new_n284), .B1(new_n398), .B2(new_n291), .ZN(new_n399));
  AND2_X1   g0199(.A1(new_n283), .A2(new_n209), .ZN(new_n400));
  INV_X1    g0200(.A(KEYINPUT71), .ZN(new_n401));
  NAND3_X1  g0201(.A1(new_n400), .A2(new_n401), .A3(new_n290), .ZN(new_n402));
  OAI21_X1  g0202(.A(KEYINPUT71), .B1(new_n291), .B2(new_n284), .ZN(new_n403));
  AOI21_X1  g0203(.A(new_n287), .B1(new_n402), .B2(new_n403), .ZN(new_n404));
  INV_X1    g0204(.A(KEYINPUT72), .ZN(new_n405));
  AND3_X1   g0205(.A1(new_n404), .A2(new_n405), .A3(G77), .ZN(new_n406));
  AOI21_X1  g0206(.A(new_n405), .B1(new_n404), .B2(G77), .ZN(new_n407));
  NOR2_X1   g0207(.A1(new_n406), .A2(new_n407), .ZN(new_n408));
  NAND4_X1  g0208(.A1(new_n392), .A2(new_n394), .A3(new_n399), .A4(new_n408), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n252), .A2(new_n263), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n215), .A2(G1698), .ZN(new_n411));
  OAI211_X1 g0211(.A(new_n410), .B(new_n411), .C1(new_n318), .C2(new_n319), .ZN(new_n412));
  NAND2_X1  g0212(.A1(G33), .A2(G97), .ZN(new_n413));
  NAND2_X1  g0213(.A1(new_n412), .A2(new_n413), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n414), .A2(new_n270), .ZN(new_n415));
  AND3_X1   g0215(.A1(new_n248), .A2(G238), .A3(new_n250), .ZN(new_n416));
  INV_X1    g0216(.A(new_n416), .ZN(new_n417));
  NAND3_X1  g0217(.A1(new_n415), .A2(new_n272), .A3(new_n417), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n418), .A2(KEYINPUT13), .ZN(new_n419));
  AOI21_X1  g0219(.A(new_n255), .B1(new_n414), .B2(new_n270), .ZN(new_n420));
  INV_X1    g0220(.A(KEYINPUT13), .ZN(new_n421));
  NAND3_X1  g0221(.A1(new_n420), .A2(new_n421), .A3(new_n417), .ZN(new_n422));
  NAND3_X1  g0222(.A1(new_n419), .A2(G190), .A3(new_n422), .ZN(new_n423));
  AOI21_X1  g0223(.A(new_n421), .B1(new_n420), .B2(new_n417), .ZN(new_n424));
  AOI22_X1  g0224(.A1(new_n412), .A2(new_n413), .B1(new_n267), .B2(new_n269), .ZN(new_n425));
  NOR4_X1   g0225(.A1(new_n425), .A2(KEYINPUT13), .A3(new_n416), .A4(new_n255), .ZN(new_n426));
  OAI21_X1  g0226(.A(G200), .B1(new_n424), .B2(new_n426), .ZN(new_n427));
  NAND3_X1  g0227(.A1(new_n208), .A2(G33), .A3(G77), .ZN(new_n428));
  OAI221_X1 g0228(.A(new_n428), .B1(new_n208), .B2(G68), .C1(new_n279), .C2(new_n292), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n429), .A2(new_n284), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n430), .A2(KEYINPUT11), .ZN(new_n431));
  INV_X1    g0231(.A(KEYINPUT11), .ZN(new_n432));
  NAND3_X1  g0232(.A1(new_n429), .A2(new_n432), .A3(new_n284), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n431), .A2(new_n433), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n404), .A2(G68), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n291), .A2(new_n203), .ZN(new_n436));
  XNOR2_X1  g0236(.A(new_n436), .B(KEYINPUT12), .ZN(new_n437));
  AND3_X1   g0237(.A1(new_n434), .A2(new_n435), .A3(new_n437), .ZN(new_n438));
  AND3_X1   g0238(.A1(new_n423), .A2(new_n427), .A3(new_n438), .ZN(new_n439));
  OAI21_X1  g0239(.A(G169), .B1(new_n424), .B2(new_n426), .ZN(new_n440));
  NAND2_X1  g0240(.A1(new_n440), .A2(KEYINPUT14), .ZN(new_n441));
  NAND3_X1  g0241(.A1(new_n419), .A2(G179), .A3(new_n422), .ZN(new_n442));
  INV_X1    g0242(.A(KEYINPUT14), .ZN(new_n443));
  OAI211_X1 g0243(.A(new_n443), .B(G169), .C1(new_n424), .C2(new_n426), .ZN(new_n444));
  NAND3_X1  g0244(.A1(new_n441), .A2(new_n442), .A3(new_n444), .ZN(new_n445));
  INV_X1    g0245(.A(new_n438), .ZN(new_n446));
  AOI21_X1  g0246(.A(new_n439), .B1(new_n445), .B2(new_n446), .ZN(new_n447));
  NAND2_X1  g0247(.A1(new_n391), .A2(new_n295), .ZN(new_n448));
  NAND2_X1  g0248(.A1(new_n404), .A2(G77), .ZN(new_n449));
  NAND2_X1  g0249(.A1(new_n449), .A2(KEYINPUT72), .ZN(new_n450));
  NAND3_X1  g0250(.A1(new_n404), .A2(new_n405), .A3(G77), .ZN(new_n451));
  NAND3_X1  g0251(.A1(new_n450), .A2(new_n399), .A3(new_n451), .ZN(new_n452));
  NAND3_X1  g0252(.A1(new_n393), .A2(new_n357), .A3(new_n390), .ZN(new_n453));
  NAND3_X1  g0253(.A1(new_n448), .A2(new_n452), .A3(new_n453), .ZN(new_n454));
  AND4_X1   g0254(.A1(new_n380), .A2(new_n409), .A3(new_n447), .A4(new_n454), .ZN(new_n455));
  OAI211_X1 g0255(.A(G264), .B(G1698), .C1(new_n318), .C2(new_n319), .ZN(new_n456));
  OAI211_X1 g0256(.A(G257), .B(new_n263), .C1(new_n318), .C2(new_n319), .ZN(new_n457));
  NAND3_X1  g0257(.A1(new_n259), .A2(G303), .A3(new_n260), .ZN(new_n458));
  NAND3_X1  g0258(.A1(new_n456), .A2(new_n457), .A3(new_n458), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n459), .A2(KEYINPUT83), .ZN(new_n460));
  INV_X1    g0260(.A(KEYINPUT83), .ZN(new_n461));
  NAND4_X1  g0261(.A1(new_n456), .A2(new_n457), .A3(new_n461), .A4(new_n458), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n460), .A2(new_n462), .ZN(new_n463));
  AOI21_X1  g0263(.A(KEYINPUT84), .B1(new_n463), .B2(new_n270), .ZN(new_n464));
  INV_X1    g0264(.A(KEYINPUT84), .ZN(new_n465));
  INV_X1    g0265(.A(new_n270), .ZN(new_n466));
  AOI211_X1 g0266(.A(new_n465), .B(new_n466), .C1(new_n460), .C2(new_n462), .ZN(new_n467));
  INV_X1    g0267(.A(G41), .ZN(new_n468));
  OAI211_X1 g0268(.A(new_n249), .B(G45), .C1(new_n468), .C2(KEYINPUT5), .ZN(new_n469));
  INV_X1    g0269(.A(KEYINPUT5), .ZN(new_n470));
  NOR2_X1   g0270(.A1(new_n470), .A2(G41), .ZN(new_n471));
  OR2_X1    g0271(.A1(new_n469), .A2(new_n471), .ZN(new_n472));
  AND2_X1   g0272(.A1(new_n472), .A2(new_n248), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n473), .A2(G270), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n469), .A2(KEYINPUT78), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n470), .A2(G41), .ZN(new_n476));
  INV_X1    g0276(.A(KEYINPUT78), .ZN(new_n477));
  NAND4_X1  g0277(.A1(new_n476), .A2(new_n477), .A3(new_n249), .A4(G45), .ZN(new_n478));
  NOR2_X1   g0278(.A1(new_n471), .A2(new_n254), .ZN(new_n479));
  NAND4_X1  g0279(.A1(new_n475), .A2(new_n478), .A3(new_n479), .A4(new_n248), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n474), .A2(new_n480), .ZN(new_n481));
  NOR3_X1   g0281(.A1(new_n464), .A2(new_n467), .A3(new_n481), .ZN(new_n482));
  NAND2_X1  g0282(.A1(G33), .A2(G283), .ZN(new_n483));
  INV_X1    g0283(.A(G97), .ZN(new_n484));
  OAI211_X1 g0284(.A(new_n483), .B(new_n208), .C1(G33), .C2(new_n484), .ZN(new_n485));
  OAI211_X1 g0285(.A(new_n485), .B(new_n284), .C1(new_n208), .C2(G116), .ZN(new_n486));
  INV_X1    g0286(.A(KEYINPUT20), .ZN(new_n487));
  XNOR2_X1  g0287(.A(new_n486), .B(new_n487), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n402), .A2(new_n403), .ZN(new_n489));
  NOR2_X1   g0289(.A1(new_n258), .A2(G1), .ZN(new_n490));
  XNOR2_X1  g0290(.A(new_n490), .B(KEYINPUT77), .ZN(new_n491));
  NAND3_X1  g0291(.A1(new_n489), .A2(G116), .A3(new_n491), .ZN(new_n492));
  OAI211_X1 g0292(.A(new_n488), .B(new_n492), .C1(G116), .C2(new_n290), .ZN(new_n493));
  NAND3_X1  g0293(.A1(new_n482), .A2(G179), .A3(new_n493), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n463), .A2(new_n270), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n495), .A2(new_n465), .ZN(new_n496));
  AND2_X1   g0296(.A1(new_n474), .A2(new_n480), .ZN(new_n497));
  NAND3_X1  g0297(.A1(new_n463), .A2(KEYINPUT84), .A3(new_n270), .ZN(new_n498));
  NAND4_X1  g0298(.A1(new_n496), .A2(G190), .A3(new_n497), .A4(new_n498), .ZN(new_n499));
  INV_X1    g0299(.A(new_n493), .ZN(new_n500));
  OAI211_X1 g0300(.A(new_n499), .B(new_n500), .C1(new_n482), .C2(new_n349), .ZN(new_n501));
  INV_X1    g0301(.A(KEYINPUT21), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n493), .A2(G169), .ZN(new_n503));
  OAI21_X1  g0303(.A(new_n502), .B1(new_n482), .B2(new_n503), .ZN(new_n504));
  NAND3_X1  g0304(.A1(new_n496), .A2(new_n497), .A3(new_n498), .ZN(new_n505));
  NAND4_X1  g0305(.A1(new_n505), .A2(KEYINPUT21), .A3(G169), .A4(new_n493), .ZN(new_n506));
  AND4_X1   g0306(.A1(new_n494), .A2(new_n501), .A3(new_n504), .A4(new_n506), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n291), .A2(new_n484), .ZN(new_n508));
  NOR2_X1   g0308(.A1(new_n291), .A2(new_n284), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n491), .A2(new_n509), .ZN(new_n510));
  OAI21_X1  g0310(.A(new_n508), .B1(new_n510), .B2(new_n484), .ZN(new_n511));
  NOR2_X1   g0311(.A1(new_n279), .A2(new_n398), .ZN(new_n512));
  OR2_X1    g0312(.A1(new_n512), .A2(KEYINPUT76), .ZN(new_n513));
  XNOR2_X1  g0313(.A(G97), .B(G107), .ZN(new_n514));
  INV_X1    g0314(.A(KEYINPUT6), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  NOR3_X1   g0316(.A1(new_n515), .A2(new_n484), .A3(G107), .ZN(new_n517));
  INV_X1    g0317(.A(new_n517), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n516), .A2(new_n518), .ZN(new_n519));
  AOI22_X1  g0319(.A1(new_n519), .A2(G20), .B1(KEYINPUT76), .B2(new_n512), .ZN(new_n520));
  INV_X1    g0320(.A(G107), .ZN(new_n521));
  OAI211_X1 g0321(.A(new_n513), .B(new_n520), .C1(new_n323), .C2(new_n521), .ZN(new_n522));
  AOI21_X1  g0322(.A(new_n511), .B1(new_n522), .B2(new_n284), .ZN(new_n523));
  INV_X1    g0323(.A(G244), .ZN(new_n524));
  NOR2_X1   g0324(.A1(new_n524), .A2(G1698), .ZN(new_n525));
  OAI21_X1  g0325(.A(new_n525), .B1(new_n318), .B2(new_n319), .ZN(new_n526));
  INV_X1    g0326(.A(KEYINPUT4), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  NAND3_X1  g0328(.A1(new_n261), .A2(G250), .A3(G1698), .ZN(new_n529));
  NAND3_X1  g0329(.A1(new_n261), .A2(KEYINPUT4), .A3(new_n525), .ZN(new_n530));
  NAND4_X1  g0330(.A1(new_n528), .A2(new_n529), .A3(new_n530), .A4(new_n483), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n531), .A2(new_n270), .ZN(new_n532));
  OAI211_X1 g0332(.A(G257), .B(new_n248), .C1(new_n469), .C2(new_n471), .ZN(new_n533));
  AND2_X1   g0333(.A1(new_n480), .A2(new_n533), .ZN(new_n534));
  AND2_X1   g0334(.A1(new_n532), .A2(new_n534), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n535), .A2(G190), .ZN(new_n536));
  INV_X1    g0336(.A(KEYINPUT79), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n532), .A2(new_n534), .ZN(new_n538));
  AOI21_X1  g0338(.A(new_n537), .B1(new_n538), .B2(G200), .ZN(new_n539));
  AOI211_X1 g0339(.A(KEYINPUT79), .B(new_n349), .C1(new_n532), .C2(new_n534), .ZN(new_n540));
  OAI211_X1 g0340(.A(new_n523), .B(new_n536), .C1(new_n539), .C2(new_n540), .ZN(new_n541));
  AND2_X1   g0341(.A1(KEYINPUT85), .A2(KEYINPUT22), .ZN(new_n542));
  NOR2_X1   g0342(.A1(KEYINPUT85), .A2(KEYINPUT22), .ZN(new_n543));
  NOR2_X1   g0343(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  NAND4_X1  g0344(.A1(new_n261), .A2(new_n544), .A3(new_n208), .A4(G87), .ZN(new_n545));
  OAI211_X1 g0345(.A(new_n208), .B(G87), .C1(new_n318), .C2(new_n319), .ZN(new_n546));
  XNOR2_X1  g0346(.A(KEYINPUT85), .B(KEYINPUT22), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n546), .A2(new_n547), .ZN(new_n548));
  OAI21_X1  g0348(.A(KEYINPUT23), .B1(new_n208), .B2(G107), .ZN(new_n549));
  INV_X1    g0349(.A(KEYINPUT23), .ZN(new_n550));
  NAND3_X1  g0350(.A1(new_n550), .A2(new_n521), .A3(G20), .ZN(new_n551));
  NAND3_X1  g0351(.A1(new_n208), .A2(G33), .A3(G116), .ZN(new_n552));
  AND3_X1   g0352(.A1(new_n549), .A2(new_n551), .A3(new_n552), .ZN(new_n553));
  NAND3_X1  g0353(.A1(new_n545), .A2(new_n548), .A3(new_n553), .ZN(new_n554));
  INV_X1    g0354(.A(KEYINPUT24), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  NAND4_X1  g0356(.A1(new_n545), .A2(new_n548), .A3(KEYINPUT24), .A4(new_n553), .ZN(new_n557));
  NAND3_X1  g0357(.A1(new_n556), .A2(new_n284), .A3(new_n557), .ZN(new_n558));
  NOR2_X1   g0358(.A1(new_n290), .A2(G107), .ZN(new_n559));
  XNOR2_X1  g0359(.A(new_n559), .B(KEYINPUT25), .ZN(new_n560));
  AND2_X1   g0360(.A1(new_n558), .A2(new_n560), .ZN(new_n561));
  NAND3_X1  g0361(.A1(new_n261), .A2(G257), .A3(G1698), .ZN(new_n562));
  NAND3_X1  g0362(.A1(new_n261), .A2(G250), .A3(new_n263), .ZN(new_n563));
  INV_X1    g0363(.A(G294), .ZN(new_n564));
  OAI211_X1 g0364(.A(new_n562), .B(new_n563), .C1(new_n258), .C2(new_n564), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n565), .A2(new_n270), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n473), .A2(G264), .ZN(new_n567));
  NAND4_X1  g0367(.A1(new_n566), .A2(new_n567), .A3(G190), .A4(new_n480), .ZN(new_n568));
  INV_X1    g0368(.A(new_n510), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n569), .A2(G107), .ZN(new_n570));
  NAND3_X1  g0370(.A1(new_n566), .A2(new_n567), .A3(new_n480), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n571), .A2(G200), .ZN(new_n572));
  NAND4_X1  g0372(.A1(new_n561), .A2(new_n568), .A3(new_n570), .A4(new_n572), .ZN(new_n573));
  NAND3_X1  g0373(.A1(new_n532), .A2(new_n357), .A3(new_n534), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n538), .A2(new_n295), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n512), .A2(KEYINPUT76), .ZN(new_n576));
  AOI21_X1  g0376(.A(new_n517), .B1(new_n515), .B2(new_n514), .ZN(new_n577));
  OAI21_X1  g0377(.A(new_n576), .B1(new_n577), .B2(new_n208), .ZN(new_n578));
  AOI21_X1  g0378(.A(new_n578), .B1(G107), .B2(new_n368), .ZN(new_n579));
  AOI21_X1  g0379(.A(new_n400), .B1(new_n579), .B2(new_n513), .ZN(new_n580));
  OAI211_X1 g0380(.A(new_n574), .B(new_n575), .C1(new_n580), .C2(new_n511), .ZN(new_n581));
  NAND3_X1  g0381(.A1(new_n558), .A2(new_n570), .A3(new_n560), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n571), .A2(new_n295), .ZN(new_n583));
  NAND4_X1  g0383(.A1(new_n566), .A2(new_n567), .A3(new_n357), .A4(new_n480), .ZN(new_n584));
  NAND3_X1  g0384(.A1(new_n582), .A2(new_n583), .A3(new_n584), .ZN(new_n585));
  NAND4_X1  g0385(.A1(new_n541), .A2(new_n573), .A3(new_n581), .A4(new_n585), .ZN(new_n586));
  INV_X1    g0386(.A(KEYINPUT19), .ZN(new_n587));
  OAI21_X1  g0387(.A(new_n208), .B1(new_n413), .B2(new_n587), .ZN(new_n588));
  INV_X1    g0388(.A(G87), .ZN(new_n589));
  AND4_X1   g0389(.A1(KEYINPUT81), .A2(new_n589), .A3(new_n484), .A4(new_n521), .ZN(new_n590));
  NOR2_X1   g0390(.A1(G97), .A2(G107), .ZN(new_n591));
  AOI21_X1  g0391(.A(KEYINPUT81), .B1(new_n591), .B2(new_n589), .ZN(new_n592));
  OAI21_X1  g0392(.A(new_n588), .B1(new_n590), .B2(new_n592), .ZN(new_n593));
  INV_X1    g0393(.A(KEYINPUT82), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  AOI21_X1  g0395(.A(G20), .B1(new_n259), .B2(new_n260), .ZN(new_n596));
  NAND3_X1  g0396(.A1(new_n208), .A2(G33), .A3(G97), .ZN(new_n597));
  AOI22_X1  g0397(.A1(new_n596), .A2(G68), .B1(new_n597), .B2(new_n587), .ZN(new_n598));
  OAI211_X1 g0398(.A(KEYINPUT82), .B(new_n588), .C1(new_n590), .C2(new_n592), .ZN(new_n599));
  NAND3_X1  g0399(.A1(new_n595), .A2(new_n598), .A3(new_n599), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n600), .A2(new_n284), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n396), .A2(new_n291), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n569), .A2(G87), .ZN(new_n603));
  AND3_X1   g0403(.A1(new_n601), .A2(new_n602), .A3(new_n603), .ZN(new_n604));
  INV_X1    g0404(.A(KEYINPUT80), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n249), .A2(G45), .ZN(new_n606));
  OAI21_X1  g0406(.A(new_n605), .B1(new_n606), .B2(new_n254), .ZN(new_n607));
  NAND4_X1  g0407(.A1(new_n249), .A2(KEYINPUT80), .A3(G45), .A4(G274), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  NAND3_X1  g0409(.A1(new_n248), .A2(G250), .A3(new_n606), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n609), .A2(new_n610), .ZN(new_n611));
  INV_X1    g0411(.A(new_n611), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n524), .A2(G1698), .ZN(new_n613));
  OAI221_X1 g0413(.A(new_n613), .B1(G238), .B2(G1698), .C1(new_n318), .C2(new_n319), .ZN(new_n614));
  NAND2_X1  g0414(.A1(G33), .A2(G116), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n616), .A2(new_n270), .ZN(new_n617));
  NAND3_X1  g0417(.A1(new_n612), .A2(new_n617), .A3(G190), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n612), .A2(new_n617), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n619), .A2(G200), .ZN(new_n620));
  NAND3_X1  g0420(.A1(new_n604), .A2(new_n618), .A3(new_n620), .ZN(new_n621));
  INV_X1    g0421(.A(new_n396), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n569), .A2(new_n622), .ZN(new_n623));
  NAND3_X1  g0423(.A1(new_n601), .A2(new_n602), .A3(new_n623), .ZN(new_n624));
  INV_X1    g0424(.A(new_n619), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n625), .A2(new_n357), .ZN(new_n626));
  OAI211_X1 g0426(.A(new_n624), .B(new_n626), .C1(G169), .C2(new_n625), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n621), .A2(new_n627), .ZN(new_n628));
  NOR2_X1   g0428(.A1(new_n586), .A2(new_n628), .ZN(new_n629));
  AND3_X1   g0429(.A1(new_n455), .A2(new_n507), .A3(new_n629), .ZN(G372));
  AND3_X1   g0430(.A1(new_n609), .A2(KEYINPUT86), .A3(new_n610), .ZN(new_n631));
  AOI21_X1  g0431(.A(KEYINPUT86), .B1(new_n609), .B2(new_n610), .ZN(new_n632));
  OAI21_X1  g0432(.A(new_n617), .B1(new_n631), .B2(new_n632), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n633), .A2(G200), .ZN(new_n634));
  AOI22_X1  g0434(.A1(new_n600), .A2(new_n284), .B1(new_n291), .B2(new_n396), .ZN(new_n635));
  NAND4_X1  g0435(.A1(new_n634), .A2(new_n635), .A3(new_n603), .A4(new_n618), .ZN(new_n636));
  AND4_X1   g0436(.A1(new_n581), .A2(new_n541), .A3(new_n573), .A4(new_n636), .ZN(new_n637));
  NAND4_X1  g0437(.A1(new_n504), .A2(new_n506), .A3(new_n494), .A4(new_n585), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n633), .A2(new_n295), .ZN(new_n640));
  NAND3_X1  g0440(.A1(new_n624), .A2(new_n626), .A3(new_n640), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n575), .A2(new_n574), .ZN(new_n642));
  NOR2_X1   g0442(.A1(new_n642), .A2(new_n523), .ZN(new_n643));
  INV_X1    g0443(.A(KEYINPUT26), .ZN(new_n644));
  NAND4_X1  g0444(.A1(new_n643), .A2(new_n644), .A3(new_n641), .A4(new_n636), .ZN(new_n645));
  OAI21_X1  g0445(.A(KEYINPUT26), .B1(new_n628), .B2(new_n581), .ZN(new_n646));
  NAND4_X1  g0446(.A1(new_n639), .A2(new_n641), .A3(new_n645), .A4(new_n646), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n455), .A2(new_n647), .ZN(new_n648));
  XOR2_X1   g0448(.A(new_n648), .B(KEYINPUT87), .Z(new_n649));
  INV_X1    g0449(.A(new_n297), .ZN(new_n650));
  OAI21_X1  g0450(.A(new_n360), .B1(new_n295), .B2(new_n347), .ZN(new_n651));
  AOI21_X1  g0451(.A(new_n338), .B1(new_n324), .B2(new_n325), .ZN(new_n652));
  OAI21_X1  g0452(.A(new_n651), .B1(new_n652), .B2(new_n311), .ZN(new_n653));
  NOR2_X1   g0453(.A1(new_n653), .A2(new_n377), .ZN(new_n654));
  AOI21_X1  g0454(.A(KEYINPUT18), .B1(new_n376), .B2(new_n651), .ZN(new_n655));
  OR2_X1    g0455(.A1(new_n654), .A2(new_n655), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n445), .A2(new_n446), .ZN(new_n657));
  OAI21_X1  g0457(.A(new_n657), .B1(new_n439), .B2(new_n454), .ZN(new_n658));
  XOR2_X1   g0458(.A(new_n658), .B(KEYINPUT88), .Z(new_n659));
  AND2_X1   g0459(.A1(new_n351), .A2(new_n373), .ZN(new_n660));
  INV_X1    g0460(.A(new_n660), .ZN(new_n661));
  OAI21_X1  g0461(.A(new_n656), .B1(new_n659), .B2(new_n661), .ZN(new_n662));
  AND2_X1   g0462(.A1(new_n299), .A2(new_n301), .ZN(new_n663));
  INV_X1    g0463(.A(KEYINPUT10), .ZN(new_n664));
  NAND4_X1  g0464(.A1(new_n663), .A2(new_n664), .A3(new_n300), .A4(new_n303), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n665), .A2(new_n305), .ZN(new_n666));
  AOI21_X1  g0466(.A(new_n650), .B1(new_n662), .B2(new_n666), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n649), .A2(new_n667), .ZN(G369));
  NAND3_X1  g0468(.A1(new_n504), .A2(new_n506), .A3(new_n494), .ZN(new_n669));
  INV_X1    g0469(.A(G13), .ZN(new_n670));
  NOR2_X1   g0470(.A1(new_n670), .A2(G20), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n671), .A2(new_n249), .ZN(new_n672));
  OR2_X1    g0472(.A1(new_n672), .A2(KEYINPUT27), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n672), .A2(KEYINPUT27), .ZN(new_n674));
  NAND3_X1  g0474(.A1(new_n673), .A2(G213), .A3(new_n674), .ZN(new_n675));
  INV_X1    g0475(.A(G343), .ZN(new_n676));
  NOR2_X1   g0476(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n493), .A2(new_n677), .ZN(new_n678));
  MUX2_X1   g0478(.A(new_n669), .B(new_n507), .S(new_n678), .Z(new_n679));
  NAND2_X1  g0479(.A1(new_n582), .A2(new_n677), .ZN(new_n680));
  AND2_X1   g0480(.A1(new_n573), .A2(new_n680), .ZN(new_n681));
  MUX2_X1   g0481(.A(new_n677), .B(new_n681), .S(new_n585), .Z(new_n682));
  NAND3_X1  g0482(.A1(new_n679), .A2(G330), .A3(new_n682), .ZN(new_n683));
  INV_X1    g0483(.A(new_n677), .ZN(new_n684));
  AND2_X1   g0484(.A1(new_n669), .A2(new_n684), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n682), .A2(new_n685), .ZN(new_n686));
  INV_X1    g0486(.A(KEYINPUT89), .ZN(new_n687));
  OR2_X1    g0487(.A1(new_n585), .A2(new_n677), .ZN(new_n688));
  NAND3_X1  g0488(.A1(new_n686), .A2(new_n687), .A3(new_n688), .ZN(new_n689));
  INV_X1    g0489(.A(new_n689), .ZN(new_n690));
  AOI21_X1  g0490(.A(new_n687), .B1(new_n686), .B2(new_n688), .ZN(new_n691));
  OAI21_X1  g0491(.A(new_n683), .B1(new_n690), .B2(new_n691), .ZN(G399));
  INV_X1    g0492(.A(new_n226), .ZN(new_n693));
  NOR2_X1   g0493(.A1(new_n693), .A2(G41), .ZN(new_n694));
  INV_X1    g0494(.A(new_n694), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n695), .A2(G1), .ZN(new_n696));
  NOR2_X1   g0496(.A1(new_n590), .A2(new_n592), .ZN(new_n697));
  INV_X1    g0497(.A(G116), .ZN(new_n698));
  NAND2_X1  g0498(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  OAI22_X1  g0499(.A1(new_n696), .A2(new_n699), .B1(new_n207), .B2(new_n695), .ZN(new_n700));
  XOR2_X1   g0500(.A(KEYINPUT90), .B(KEYINPUT28), .Z(new_n701));
  XNOR2_X1  g0501(.A(new_n700), .B(new_n701), .ZN(new_n702));
  INV_X1    g0502(.A(new_n641), .ZN(new_n703));
  AOI21_X1  g0503(.A(new_n703), .B1(new_n637), .B2(new_n638), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n641), .A2(new_n636), .ZN(new_n705));
  OAI21_X1  g0505(.A(KEYINPUT26), .B1(new_n705), .B2(new_n581), .ZN(new_n706));
  NAND4_X1  g0506(.A1(new_n643), .A2(new_n621), .A3(new_n627), .A4(new_n644), .ZN(new_n707));
  AND2_X1   g0507(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  AOI21_X1  g0508(.A(new_n677), .B1(new_n704), .B2(new_n708), .ZN(new_n709));
  NAND2_X1  g0509(.A1(new_n709), .A2(KEYINPUT29), .ZN(new_n710));
  AND2_X1   g0510(.A1(new_n647), .A2(new_n684), .ZN(new_n711));
  OAI21_X1  g0511(.A(new_n710), .B1(new_n711), .B2(KEYINPUT29), .ZN(new_n712));
  INV_X1    g0512(.A(KEYINPUT30), .ZN(new_n713));
  NAND4_X1  g0513(.A1(new_n496), .A2(G179), .A3(new_n497), .A4(new_n498), .ZN(new_n714));
  NAND4_X1  g0514(.A1(new_n535), .A2(new_n625), .A3(new_n566), .A4(new_n567), .ZN(new_n715));
  OAI21_X1  g0515(.A(new_n713), .B1(new_n714), .B2(new_n715), .ZN(new_n716));
  NAND2_X1  g0516(.A1(new_n566), .A2(new_n567), .ZN(new_n717));
  NOR3_X1   g0517(.A1(new_n717), .A2(new_n538), .A3(new_n619), .ZN(new_n718));
  NAND4_X1  g0518(.A1(new_n482), .A2(new_n718), .A3(KEYINPUT30), .A4(G179), .ZN(new_n719));
  NAND4_X1  g0519(.A1(new_n505), .A2(new_n357), .A3(new_n571), .A4(new_n633), .ZN(new_n720));
  OAI211_X1 g0520(.A(new_n716), .B(new_n719), .C1(new_n720), .C2(new_n535), .ZN(new_n721));
  NAND2_X1  g0521(.A1(new_n721), .A2(new_n677), .ZN(new_n722));
  INV_X1    g0522(.A(KEYINPUT31), .ZN(new_n723));
  NAND2_X1  g0523(.A1(new_n722), .A2(new_n723), .ZN(new_n724));
  NAND3_X1  g0524(.A1(new_n507), .A2(new_n629), .A3(new_n684), .ZN(new_n725));
  NAND3_X1  g0525(.A1(new_n721), .A2(KEYINPUT31), .A3(new_n677), .ZN(new_n726));
  NAND3_X1  g0526(.A1(new_n724), .A2(new_n725), .A3(new_n726), .ZN(new_n727));
  NAND2_X1  g0527(.A1(new_n727), .A2(G330), .ZN(new_n728));
  NAND2_X1  g0528(.A1(new_n712), .A2(new_n728), .ZN(new_n729));
  INV_X1    g0529(.A(new_n729), .ZN(new_n730));
  OAI21_X1  g0530(.A(new_n702), .B1(new_n730), .B2(G1), .ZN(G364));
  OR2_X1    g0531(.A1(new_n679), .A2(G330), .ZN(new_n732));
  NAND2_X1  g0532(.A1(new_n679), .A2(G330), .ZN(new_n733));
  NAND2_X1  g0533(.A1(new_n671), .A2(G45), .ZN(new_n734));
  NAND3_X1  g0534(.A1(new_n695), .A2(G1), .A3(new_n734), .ZN(new_n735));
  NAND3_X1  g0535(.A1(new_n732), .A2(new_n733), .A3(new_n735), .ZN(new_n736));
  NOR2_X1   g0536(.A1(new_n208), .A2(new_n357), .ZN(new_n737));
  NAND3_X1  g0537(.A1(new_n737), .A2(new_n302), .A3(G200), .ZN(new_n738));
  OR2_X1    g0538(.A1(KEYINPUT33), .A2(G317), .ZN(new_n739));
  NAND2_X1  g0539(.A1(KEYINPUT33), .A2(G317), .ZN(new_n740));
  AOI21_X1  g0540(.A(new_n738), .B1(new_n739), .B2(new_n740), .ZN(new_n741));
  NOR2_X1   g0541(.A1(new_n349), .A2(G179), .ZN(new_n742));
  NOR2_X1   g0542(.A1(new_n208), .A2(G190), .ZN(new_n743));
  NAND2_X1  g0543(.A1(new_n742), .A2(new_n743), .ZN(new_n744));
  INV_X1    g0544(.A(new_n744), .ZN(new_n745));
  NAND2_X1  g0545(.A1(new_n745), .A2(G283), .ZN(new_n746));
  INV_X1    g0546(.A(new_n737), .ZN(new_n747));
  NOR3_X1   g0547(.A1(new_n747), .A2(G190), .A3(G200), .ZN(new_n748));
  INV_X1    g0548(.A(new_n748), .ZN(new_n749));
  INV_X1    g0549(.A(G311), .ZN(new_n750));
  OAI211_X1 g0550(.A(new_n332), .B(new_n746), .C1(new_n749), .C2(new_n750), .ZN(new_n751));
  NOR3_X1   g0551(.A1(new_n747), .A2(new_n302), .A3(G200), .ZN(new_n752));
  AOI211_X1 g0552(.A(new_n741), .B(new_n751), .C1(G322), .C2(new_n752), .ZN(new_n753));
  NAND3_X1  g0553(.A1(new_n742), .A2(G20), .A3(G190), .ZN(new_n754));
  INV_X1    g0554(.A(new_n754), .ZN(new_n755));
  NAND2_X1  g0555(.A1(new_n755), .A2(G303), .ZN(new_n756));
  NAND3_X1  g0556(.A1(new_n737), .A2(G190), .A3(G200), .ZN(new_n757));
  AND2_X1   g0557(.A1(new_n757), .A2(KEYINPUT93), .ZN(new_n758));
  NOR2_X1   g0558(.A1(new_n757), .A2(KEYINPUT93), .ZN(new_n759));
  NOR2_X1   g0559(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  INV_X1    g0560(.A(new_n760), .ZN(new_n761));
  XNOR2_X1  g0561(.A(KEYINPUT96), .B(G326), .ZN(new_n762));
  NAND2_X1  g0562(.A1(new_n761), .A2(new_n762), .ZN(new_n763));
  NOR2_X1   g0563(.A1(G179), .A2(G200), .ZN(new_n764));
  NAND2_X1  g0564(.A1(new_n743), .A2(new_n764), .ZN(new_n765));
  INV_X1    g0565(.A(new_n765), .ZN(new_n766));
  AOI21_X1  g0566(.A(new_n208), .B1(new_n764), .B2(G190), .ZN(new_n767));
  INV_X1    g0567(.A(new_n767), .ZN(new_n768));
  AOI22_X1  g0568(.A1(G329), .A2(new_n766), .B1(new_n768), .B2(G294), .ZN(new_n769));
  NAND4_X1  g0569(.A1(new_n753), .A2(new_n756), .A3(new_n763), .A4(new_n769), .ZN(new_n770));
  INV_X1    g0570(.A(new_n752), .ZN(new_n771));
  OAI22_X1  g0571(.A1(new_n749), .A2(new_n398), .B1(new_n771), .B2(new_n202), .ZN(new_n772));
  AOI21_X1  g0572(.A(new_n772), .B1(G50), .B2(new_n761), .ZN(new_n773));
  XOR2_X1   g0573(.A(new_n773), .B(KEYINPUT94), .Z(new_n774));
  INV_X1    g0574(.A(new_n738), .ZN(new_n775));
  NAND2_X1  g0575(.A1(new_n775), .A2(G68), .ZN(new_n776));
  NOR2_X1   g0576(.A1(new_n754), .A2(new_n589), .ZN(new_n777));
  AOI211_X1 g0577(.A(new_n332), .B(new_n777), .C1(G107), .C2(new_n745), .ZN(new_n778));
  XNOR2_X1  g0578(.A(new_n778), .B(KEYINPUT95), .ZN(new_n779));
  NOR2_X1   g0579(.A1(new_n767), .A2(new_n484), .ZN(new_n780));
  NAND2_X1  g0580(.A1(new_n766), .A2(G159), .ZN(new_n781));
  AOI21_X1  g0581(.A(new_n780), .B1(new_n781), .B2(KEYINPUT32), .ZN(new_n782));
  NAND4_X1  g0582(.A1(new_n774), .A2(new_n776), .A3(new_n779), .A4(new_n782), .ZN(new_n783));
  NOR2_X1   g0583(.A1(new_n781), .A2(KEYINPUT32), .ZN(new_n784));
  OAI21_X1  g0584(.A(new_n770), .B1(new_n783), .B2(new_n784), .ZN(new_n785));
  AOI21_X1  g0585(.A(new_n209), .B1(G20), .B2(new_n295), .ZN(new_n786));
  NOR2_X1   g0586(.A1(G13), .A2(G33), .ZN(new_n787));
  INV_X1    g0587(.A(new_n787), .ZN(new_n788));
  NOR2_X1   g0588(.A1(new_n788), .A2(G20), .ZN(new_n789));
  NOR2_X1   g0589(.A1(new_n789), .A2(new_n786), .ZN(new_n790));
  NOR2_X1   g0590(.A1(new_n693), .A2(new_n261), .ZN(new_n791));
  OAI21_X1  g0591(.A(new_n791), .B1(G45), .B2(new_n207), .ZN(new_n792));
  XNOR2_X1  g0592(.A(new_n792), .B(KEYINPUT92), .ZN(new_n793));
  INV_X1    g0593(.A(new_n242), .ZN(new_n794));
  INV_X1    g0594(.A(G45), .ZN(new_n795));
  OAI21_X1  g0595(.A(new_n793), .B1(new_n794), .B2(new_n795), .ZN(new_n796));
  NAND2_X1  g0596(.A1(new_n261), .A2(new_n226), .ZN(new_n797));
  XNOR2_X1  g0597(.A(new_n797), .B(KEYINPUT91), .ZN(new_n798));
  AOI22_X1  g0598(.A1(new_n798), .A2(G355), .B1(new_n698), .B2(new_n693), .ZN(new_n799));
  NAND2_X1  g0599(.A1(new_n796), .A2(new_n799), .ZN(new_n800));
  AOI22_X1  g0600(.A1(new_n785), .A2(new_n786), .B1(new_n790), .B2(new_n800), .ZN(new_n801));
  INV_X1    g0601(.A(new_n735), .ZN(new_n802));
  INV_X1    g0602(.A(new_n789), .ZN(new_n803));
  OAI211_X1 g0603(.A(new_n801), .B(new_n802), .C1(new_n679), .C2(new_n803), .ZN(new_n804));
  NAND2_X1  g0604(.A1(new_n736), .A2(new_n804), .ZN(G396));
  NAND2_X1  g0605(.A1(new_n452), .A2(new_n677), .ZN(new_n806));
  AOI22_X1  g0606(.A1(new_n408), .A2(new_n399), .B1(new_n391), .B2(new_n295), .ZN(new_n807));
  AOI22_X1  g0607(.A1(new_n409), .A2(new_n806), .B1(new_n807), .B2(new_n453), .ZN(new_n808));
  NOR2_X1   g0608(.A1(new_n454), .A2(new_n677), .ZN(new_n809));
  OAI21_X1  g0609(.A(KEYINPUT99), .B1(new_n808), .B2(new_n809), .ZN(new_n810));
  INV_X1    g0610(.A(new_n454), .ZN(new_n811));
  NAND2_X1  g0611(.A1(new_n811), .A2(new_n684), .ZN(new_n812));
  INV_X1    g0612(.A(KEYINPUT99), .ZN(new_n813));
  AOI21_X1  g0613(.A(new_n349), .B1(new_n393), .B2(new_n390), .ZN(new_n814));
  NOR2_X1   g0614(.A1(new_n452), .A2(new_n814), .ZN(new_n815));
  AOI22_X1  g0615(.A1(new_n815), .A2(new_n394), .B1(new_n452), .B2(new_n677), .ZN(new_n816));
  OAI211_X1 g0616(.A(new_n812), .B(new_n813), .C1(new_n816), .C2(new_n811), .ZN(new_n817));
  NAND2_X1  g0617(.A1(new_n810), .A2(new_n817), .ZN(new_n818));
  XNOR2_X1  g0618(.A(new_n711), .B(new_n818), .ZN(new_n819));
  XNOR2_X1  g0619(.A(new_n819), .B(new_n728), .ZN(new_n820));
  NAND2_X1  g0620(.A1(new_n820), .A2(new_n735), .ZN(new_n821));
  NAND2_X1  g0621(.A1(new_n818), .A2(new_n787), .ZN(new_n822));
  AOI22_X1  g0622(.A1(new_n752), .A2(G143), .B1(new_n775), .B2(G150), .ZN(new_n823));
  INV_X1    g0623(.A(G159), .ZN(new_n824));
  INV_X1    g0624(.A(G137), .ZN(new_n825));
  OAI221_X1 g0625(.A(new_n823), .B1(new_n824), .B2(new_n749), .C1(new_n760), .C2(new_n825), .ZN(new_n826));
  XOR2_X1   g0626(.A(new_n826), .B(KEYINPUT34), .Z(new_n827));
  NOR2_X1   g0627(.A1(new_n767), .A2(new_n202), .ZN(new_n828));
  AOI22_X1  g0628(.A1(new_n755), .A2(G50), .B1(new_n745), .B2(G68), .ZN(new_n829));
  INV_X1    g0629(.A(G132), .ZN(new_n830));
  OAI21_X1  g0630(.A(new_n829), .B1(new_n830), .B2(new_n765), .ZN(new_n831));
  NOR4_X1   g0631(.A1(new_n827), .A2(new_n332), .A3(new_n828), .A4(new_n831), .ZN(new_n832));
  INV_X1    g0632(.A(KEYINPUT98), .ZN(new_n833));
  XNOR2_X1  g0633(.A(KEYINPUT97), .B(G283), .ZN(new_n834));
  AOI22_X1  g0634(.A1(new_n748), .A2(G116), .B1(new_n775), .B2(new_n834), .ZN(new_n835));
  AOI22_X1  g0635(.A1(new_n761), .A2(G303), .B1(new_n833), .B2(new_n835), .ZN(new_n836));
  AOI211_X1 g0636(.A(new_n261), .B(new_n780), .C1(new_n752), .C2(G294), .ZN(new_n837));
  OAI211_X1 g0637(.A(new_n836), .B(new_n837), .C1(new_n833), .C2(new_n835), .ZN(new_n838));
  NOR2_X1   g0638(.A1(new_n754), .A2(new_n521), .ZN(new_n839));
  NOR2_X1   g0639(.A1(new_n765), .A2(new_n750), .ZN(new_n840));
  NOR2_X1   g0640(.A1(new_n744), .A2(new_n589), .ZN(new_n841));
  NOR4_X1   g0641(.A1(new_n838), .A2(new_n839), .A3(new_n840), .A4(new_n841), .ZN(new_n842));
  OAI21_X1  g0642(.A(new_n786), .B1(new_n832), .B2(new_n842), .ZN(new_n843));
  NOR2_X1   g0643(.A1(new_n786), .A2(new_n787), .ZN(new_n844));
  NAND2_X1  g0644(.A1(new_n844), .A2(new_n398), .ZN(new_n845));
  NAND4_X1  g0645(.A1(new_n822), .A2(new_n802), .A3(new_n843), .A4(new_n845), .ZN(new_n846));
  NAND2_X1  g0646(.A1(new_n821), .A2(new_n846), .ZN(G384));
  INV_X1    g0647(.A(KEYINPUT104), .ZN(new_n848));
  NAND3_X1  g0648(.A1(new_n721), .A2(new_n848), .A3(new_n677), .ZN(new_n849));
  NAND2_X1  g0649(.A1(new_n849), .A2(new_n723), .ZN(new_n850));
  AOI21_X1  g0650(.A(new_n848), .B1(new_n721), .B2(new_n677), .ZN(new_n851));
  OAI211_X1 g0651(.A(new_n726), .B(new_n725), .C1(new_n850), .C2(new_n851), .ZN(new_n852));
  NAND3_X1  g0652(.A1(new_n455), .A2(G330), .A3(new_n852), .ZN(new_n853));
  INV_X1    g0653(.A(KEYINPUT38), .ZN(new_n854));
  NAND3_X1  g0654(.A1(new_n376), .A2(new_n359), .A3(new_n361), .ZN(new_n855));
  INV_X1    g0655(.A(new_n675), .ZN(new_n856));
  NAND2_X1  g0656(.A1(new_n376), .A2(new_n856), .ZN(new_n857));
  INV_X1    g0657(.A(KEYINPUT37), .ZN(new_n858));
  NAND4_X1  g0658(.A1(new_n855), .A2(new_n857), .A3(new_n858), .A4(new_n371), .ZN(new_n859));
  INV_X1    g0659(.A(new_n859), .ZN(new_n860));
  NAND2_X1  g0660(.A1(new_n653), .A2(new_n371), .ZN(new_n861));
  INV_X1    g0661(.A(KEYINPUT102), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n861), .A2(new_n862), .ZN(new_n863));
  NAND3_X1  g0663(.A1(new_n653), .A2(new_n371), .A3(KEYINPUT102), .ZN(new_n864));
  NAND3_X1  g0664(.A1(new_n863), .A2(new_n857), .A3(new_n864), .ZN(new_n865));
  AOI21_X1  g0665(.A(new_n860), .B1(new_n865), .B2(KEYINPUT37), .ZN(new_n866));
  AOI21_X1  g0666(.A(new_n857), .B1(new_n656), .B2(new_n660), .ZN(new_n867));
  OAI21_X1  g0667(.A(new_n854), .B1(new_n866), .B2(new_n867), .ZN(new_n868));
  AOI21_X1  g0668(.A(KEYINPUT16), .B1(new_n336), .B2(new_n314), .ZN(new_n869));
  OAI21_X1  g0669(.A(new_n310), .B1(new_n338), .B2(new_n869), .ZN(new_n870));
  NAND3_X1  g0670(.A1(new_n379), .A2(new_n856), .A3(new_n870), .ZN(new_n871));
  OAI21_X1  g0671(.A(new_n870), .B1(new_n651), .B2(new_n856), .ZN(new_n872));
  AND2_X1   g0672(.A1(new_n371), .A2(new_n872), .ZN(new_n873));
  OAI21_X1  g0673(.A(new_n859), .B1(new_n858), .B2(new_n873), .ZN(new_n874));
  NAND3_X1  g0674(.A1(new_n871), .A2(KEYINPUT38), .A3(new_n874), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n868), .A2(new_n875), .ZN(new_n876));
  NOR2_X1   g0676(.A1(new_n657), .A2(new_n684), .ZN(new_n877));
  INV_X1    g0677(.A(new_n877), .ZN(new_n878));
  INV_X1    g0678(.A(new_n439), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n446), .A2(new_n677), .ZN(new_n880));
  AND4_X1   g0680(.A1(KEYINPUT101), .A2(new_n657), .A3(new_n879), .A4(new_n880), .ZN(new_n881));
  AOI21_X1  g0681(.A(KEYINPUT101), .B1(new_n447), .B2(new_n880), .ZN(new_n882));
  OAI21_X1  g0682(.A(new_n878), .B1(new_n881), .B2(new_n882), .ZN(new_n883));
  AND2_X1   g0683(.A1(new_n810), .A2(new_n817), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  AND2_X1   g0685(.A1(new_n725), .A2(new_n726), .ZN(new_n886));
  INV_X1    g0686(.A(new_n851), .ZN(new_n887));
  NAND3_X1  g0687(.A1(new_n887), .A2(new_n723), .A3(new_n849), .ZN(new_n888));
  AOI21_X1  g0688(.A(new_n885), .B1(new_n886), .B2(new_n888), .ZN(new_n889));
  INV_X1    g0689(.A(KEYINPUT105), .ZN(new_n890));
  OAI21_X1  g0690(.A(new_n876), .B1(new_n889), .B2(new_n890), .ZN(new_n891));
  NAND3_X1  g0691(.A1(new_n657), .A2(new_n879), .A3(new_n880), .ZN(new_n892));
  INV_X1    g0692(.A(KEYINPUT101), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n892), .A2(new_n893), .ZN(new_n894));
  NAND3_X1  g0694(.A1(new_n447), .A2(KEYINPUT101), .A3(new_n880), .ZN(new_n895));
  AOI21_X1  g0695(.A(new_n877), .B1(new_n894), .B2(new_n895), .ZN(new_n896));
  NOR2_X1   g0696(.A1(new_n896), .A2(new_n818), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n852), .A2(new_n897), .ZN(new_n898));
  AND3_X1   g0698(.A1(new_n871), .A2(KEYINPUT38), .A3(new_n874), .ZN(new_n899));
  AOI21_X1  g0699(.A(KEYINPUT38), .B1(new_n871), .B2(new_n874), .ZN(new_n900));
  NOR3_X1   g0700(.A1(new_n899), .A2(new_n900), .A3(KEYINPUT40), .ZN(new_n901));
  NOR2_X1   g0701(.A1(new_n898), .A2(new_n901), .ZN(new_n902));
  NAND2_X1  g0702(.A1(KEYINPUT105), .A2(KEYINPUT40), .ZN(new_n903));
  AOI22_X1  g0703(.A1(new_n891), .A2(KEYINPUT40), .B1(new_n902), .B2(new_n903), .ZN(new_n904));
  INV_X1    g0704(.A(G330), .ZN(new_n905));
  OAI21_X1  g0705(.A(new_n853), .B1(new_n904), .B2(new_n905), .ZN(new_n906));
  AOI21_X1  g0706(.A(new_n890), .B1(new_n852), .B2(new_n897), .ZN(new_n907));
  OAI211_X1 g0707(.A(new_n373), .B(new_n351), .C1(new_n654), .C2(new_n655), .ZN(new_n908));
  INV_X1    g0708(.A(new_n857), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  AOI21_X1  g0710(.A(KEYINPUT102), .B1(new_n653), .B2(new_n371), .ZN(new_n911));
  NOR2_X1   g0711(.A1(new_n911), .A2(new_n909), .ZN(new_n912));
  AOI21_X1  g0712(.A(new_n858), .B1(new_n912), .B2(new_n864), .ZN(new_n913));
  OAI21_X1  g0713(.A(new_n910), .B1(new_n913), .B2(new_n860), .ZN(new_n914));
  AOI21_X1  g0714(.A(new_n899), .B1(new_n854), .B2(new_n914), .ZN(new_n915));
  OAI21_X1  g0715(.A(KEYINPUT40), .B1(new_n907), .B2(new_n915), .ZN(new_n916));
  OR3_X1    g0716(.A1(new_n899), .A2(new_n900), .A3(KEYINPUT40), .ZN(new_n917));
  NAND3_X1  g0717(.A1(new_n917), .A2(new_n889), .A3(new_n903), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n916), .A2(new_n918), .ZN(new_n919));
  NAND3_X1  g0719(.A1(new_n919), .A2(new_n455), .A3(new_n852), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n906), .A2(new_n920), .ZN(new_n921));
  OAI211_X1 g0721(.A(new_n455), .B(new_n710), .C1(new_n711), .C2(KEYINPUT29), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n667), .A2(new_n922), .ZN(new_n923));
  XNOR2_X1  g0723(.A(new_n921), .B(new_n923), .ZN(new_n924));
  NAND3_X1  g0724(.A1(new_n647), .A2(new_n684), .A3(new_n884), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n925), .A2(new_n812), .ZN(new_n926));
  INV_X1    g0726(.A(new_n900), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n927), .A2(new_n875), .ZN(new_n928));
  NAND3_X1  g0728(.A1(new_n926), .A2(new_n928), .A3(new_n883), .ZN(new_n929));
  NOR2_X1   g0729(.A1(new_n656), .A2(new_n856), .ZN(new_n930));
  INV_X1    g0730(.A(new_n930), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n929), .A2(new_n931), .ZN(new_n932));
  AOI21_X1  g0732(.A(KEYINPUT39), .B1(new_n868), .B2(new_n875), .ZN(new_n933));
  INV_X1    g0733(.A(KEYINPUT39), .ZN(new_n934));
  NOR3_X1   g0734(.A1(new_n899), .A2(new_n900), .A3(new_n934), .ZN(new_n935));
  NOR2_X1   g0735(.A1(new_n657), .A2(new_n677), .ZN(new_n936));
  INV_X1    g0736(.A(new_n936), .ZN(new_n937));
  NOR3_X1   g0737(.A1(new_n933), .A2(new_n935), .A3(new_n937), .ZN(new_n938));
  OAI21_X1  g0738(.A(KEYINPUT103), .B1(new_n932), .B2(new_n938), .ZN(new_n939));
  AOI21_X1  g0739(.A(new_n896), .B1(new_n925), .B2(new_n812), .ZN(new_n940));
  AOI21_X1  g0740(.A(new_n930), .B1(new_n940), .B2(new_n928), .ZN(new_n941));
  NAND3_X1  g0741(.A1(new_n927), .A2(KEYINPUT39), .A3(new_n875), .ZN(new_n942));
  OAI211_X1 g0742(.A(new_n936), .B(new_n942), .C1(new_n915), .C2(KEYINPUT39), .ZN(new_n943));
  INV_X1    g0743(.A(KEYINPUT103), .ZN(new_n944));
  NAND3_X1  g0744(.A1(new_n941), .A2(new_n943), .A3(new_n944), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n939), .A2(new_n945), .ZN(new_n946));
  XNOR2_X1  g0746(.A(new_n924), .B(new_n946), .ZN(new_n947));
  OAI21_X1  g0747(.A(new_n947), .B1(new_n249), .B2(new_n671), .ZN(new_n948));
  AOI211_X1 g0748(.A(new_n398), .B(new_n207), .C1(G58), .C2(G68), .ZN(new_n949));
  NOR2_X1   g0749(.A1(new_n201), .A2(new_n203), .ZN(new_n950));
  OAI211_X1 g0750(.A(G1), .B(new_n670), .C1(new_n949), .C2(new_n950), .ZN(new_n951));
  AOI21_X1  g0751(.A(new_n698), .B1(new_n519), .B2(KEYINPUT35), .ZN(new_n952));
  NOR2_X1   g0752(.A1(new_n209), .A2(new_n208), .ZN(new_n953));
  OAI211_X1 g0753(.A(new_n952), .B(new_n953), .C1(KEYINPUT35), .C2(new_n519), .ZN(new_n954));
  XOR2_X1   g0754(.A(KEYINPUT100), .B(KEYINPUT36), .Z(new_n955));
  XNOR2_X1  g0755(.A(new_n954), .B(new_n955), .ZN(new_n956));
  NAND3_X1  g0756(.A1(new_n948), .A2(new_n951), .A3(new_n956), .ZN(G367));
  OAI211_X1 g0757(.A(new_n541), .B(new_n581), .C1(new_n523), .C2(new_n684), .ZN(new_n958));
  OAI21_X1  g0758(.A(new_n958), .B1(new_n581), .B2(new_n684), .ZN(new_n959));
  XOR2_X1   g0759(.A(new_n959), .B(KEYINPUT106), .Z(new_n960));
  OR3_X1    g0760(.A1(new_n683), .A2(new_n960), .A3(KEYINPUT107), .ZN(new_n961));
  OAI21_X1  g0761(.A(KEYINPUT107), .B1(new_n683), .B2(new_n960), .ZN(new_n962));
  NAND2_X1  g0762(.A1(new_n961), .A2(new_n962), .ZN(new_n963));
  NOR2_X1   g0763(.A1(new_n604), .A2(new_n684), .ZN(new_n964));
  NAND2_X1  g0764(.A1(new_n703), .A2(new_n964), .ZN(new_n965));
  OAI21_X1  g0765(.A(new_n965), .B1(new_n705), .B2(new_n964), .ZN(new_n966));
  NOR2_X1   g0766(.A1(new_n966), .A2(KEYINPUT43), .ZN(new_n967));
  XOR2_X1   g0767(.A(new_n963), .B(new_n967), .Z(new_n968));
  NOR2_X1   g0768(.A1(new_n960), .A2(new_n686), .ZN(new_n969));
  XNOR2_X1  g0769(.A(new_n969), .B(KEYINPUT42), .ZN(new_n970));
  OAI21_X1  g0770(.A(new_n581), .B1(new_n960), .B2(new_n585), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n971), .A2(new_n684), .ZN(new_n972));
  AOI22_X1  g0772(.A1(new_n970), .A2(new_n972), .B1(KEYINPUT43), .B2(new_n966), .ZN(new_n973));
  XNOR2_X1  g0773(.A(new_n968), .B(new_n973), .ZN(new_n974));
  XNOR2_X1  g0774(.A(KEYINPUT108), .B(KEYINPUT41), .ZN(new_n975));
  XOR2_X1   g0775(.A(new_n694), .B(new_n975), .Z(new_n976));
  INV_X1    g0776(.A(new_n976), .ZN(new_n977));
  INV_X1    g0777(.A(new_n691), .ZN(new_n978));
  NAND3_X1  g0778(.A1(new_n978), .A2(new_n689), .A3(new_n960), .ZN(new_n979));
  XOR2_X1   g0779(.A(new_n979), .B(KEYINPUT44), .Z(new_n980));
  AOI21_X1  g0780(.A(new_n960), .B1(new_n978), .B2(new_n689), .ZN(new_n981));
  XNOR2_X1  g0781(.A(new_n981), .B(KEYINPUT45), .ZN(new_n982));
  NAND3_X1  g0782(.A1(new_n980), .A2(new_n683), .A3(new_n982), .ZN(new_n983));
  AOI21_X1  g0783(.A(new_n685), .B1(new_n679), .B2(G330), .ZN(new_n984));
  INV_X1    g0784(.A(new_n682), .ZN(new_n985));
  XNOR2_X1  g0785(.A(new_n984), .B(new_n985), .ZN(new_n986));
  NOR2_X1   g0786(.A1(new_n986), .A2(new_n729), .ZN(new_n987));
  NAND2_X1  g0787(.A1(new_n983), .A2(new_n987), .ZN(new_n988));
  AOI21_X1  g0788(.A(new_n977), .B1(new_n988), .B2(new_n730), .ZN(new_n989));
  NAND2_X1  g0789(.A1(new_n734), .A2(G1), .ZN(new_n990));
  OAI21_X1  g0790(.A(new_n974), .B1(new_n989), .B2(new_n990), .ZN(new_n991));
  INV_X1    g0791(.A(new_n791), .ZN(new_n992));
  OAI221_X1 g0792(.A(new_n790), .B1(new_n226), .B2(new_n396), .C1(new_n237), .C2(new_n992), .ZN(new_n993));
  NOR2_X1   g0793(.A1(new_n754), .A2(new_n698), .ZN(new_n994));
  AOI22_X1  g0794(.A1(new_n761), .A2(G311), .B1(KEYINPUT46), .B2(new_n994), .ZN(new_n995));
  INV_X1    g0795(.A(new_n834), .ZN(new_n996));
  OAI221_X1 g0796(.A(new_n995), .B1(KEYINPUT46), .B2(new_n994), .C1(new_n749), .C2(new_n996), .ZN(new_n997));
  AOI21_X1  g0797(.A(new_n997), .B1(G303), .B2(new_n752), .ZN(new_n998));
  INV_X1    g0798(.A(G317), .ZN(new_n999));
  OAI21_X1  g0799(.A(new_n998), .B1(new_n999), .B2(new_n765), .ZN(new_n1000));
  NOR2_X1   g0800(.A1(new_n744), .A2(new_n484), .ZN(new_n1001));
  NOR2_X1   g0801(.A1(new_n738), .A2(new_n564), .ZN(new_n1002));
  NOR3_X1   g0802(.A1(new_n1000), .A2(new_n1001), .A3(new_n1002), .ZN(new_n1003));
  OAI211_X1 g0803(.A(new_n1003), .B(new_n332), .C1(new_n521), .C2(new_n767), .ZN(new_n1004));
  NOR2_X1   g0804(.A1(new_n767), .A2(new_n203), .ZN(new_n1005));
  NOR2_X1   g0805(.A1(new_n744), .A2(new_n398), .ZN(new_n1006));
  NOR2_X1   g0806(.A1(new_n1006), .A2(new_n332), .ZN(new_n1007));
  NOR2_X1   g0807(.A1(new_n1007), .A2(KEYINPUT109), .ZN(new_n1008));
  AOI22_X1  g0808(.A1(new_n761), .A2(G143), .B1(G150), .B2(new_n752), .ZN(new_n1009));
  OAI21_X1  g0809(.A(new_n1009), .B1(new_n825), .B2(new_n765), .ZN(new_n1010));
  AOI211_X1 g0810(.A(new_n1008), .B(new_n1010), .C1(G159), .C2(new_n775), .ZN(new_n1011));
  AOI22_X1  g0811(.A1(new_n1007), .A2(KEYINPUT109), .B1(G58), .B2(new_n755), .ZN(new_n1012));
  INV_X1    g0812(.A(new_n201), .ZN(new_n1013));
  OAI211_X1 g0813(.A(new_n1011), .B(new_n1012), .C1(new_n1013), .C2(new_n749), .ZN(new_n1014));
  OAI21_X1  g0814(.A(new_n1004), .B1(new_n1005), .B2(new_n1014), .ZN(new_n1015));
  XOR2_X1   g0815(.A(new_n1015), .B(KEYINPUT47), .Z(new_n1016));
  INV_X1    g0816(.A(new_n786), .ZN(new_n1017));
  OAI211_X1 g0817(.A(new_n802), .B(new_n993), .C1(new_n1016), .C2(new_n1017), .ZN(new_n1018));
  XNOR2_X1  g0818(.A(new_n1018), .B(KEYINPUT110), .ZN(new_n1019));
  OAI21_X1  g0819(.A(new_n1019), .B1(new_n803), .B2(new_n966), .ZN(new_n1020));
  NAND2_X1  g0820(.A1(new_n991), .A2(new_n1020), .ZN(G387));
  AOI211_X1 g0821(.A(G45), .B(new_n699), .C1(G68), .C2(G77), .ZN(new_n1022));
  XNOR2_X1  g0822(.A(new_n1022), .B(KEYINPUT111), .ZN(new_n1023));
  INV_X1    g0823(.A(new_n281), .ZN(new_n1024));
  NAND2_X1  g0824(.A1(new_n1024), .A2(new_n292), .ZN(new_n1025));
  XNOR2_X1  g0825(.A(new_n1025), .B(KEYINPUT50), .ZN(new_n1026));
  OAI221_X1 g0826(.A(new_n791), .B1(new_n795), .B2(new_n234), .C1(new_n1023), .C2(new_n1026), .ZN(new_n1027));
  NAND2_X1  g0827(.A1(new_n798), .A2(new_n699), .ZN(new_n1028));
  OAI211_X1 g0828(.A(new_n1027), .B(new_n1028), .C1(G107), .C2(new_n226), .ZN(new_n1029));
  AOI22_X1  g0829(.A1(new_n985), .A2(new_n789), .B1(new_n790), .B2(new_n1029), .ZN(new_n1030));
  NOR2_X1   g0830(.A1(new_n760), .A2(new_n824), .ZN(new_n1031));
  NOR2_X1   g0831(.A1(new_n767), .A2(new_n396), .ZN(new_n1032));
  AOI21_X1  g0832(.A(new_n1032), .B1(new_n1024), .B2(new_n775), .ZN(new_n1033));
  NAND2_X1  g0833(.A1(new_n766), .A2(G150), .ZN(new_n1034));
  AOI21_X1  g0834(.A(new_n332), .B1(new_n755), .B2(G77), .ZN(new_n1035));
  NAND2_X1  g0835(.A1(new_n752), .A2(G50), .ZN(new_n1036));
  NAND4_X1  g0836(.A1(new_n1033), .A2(new_n1034), .A3(new_n1035), .A4(new_n1036), .ZN(new_n1037));
  NOR2_X1   g0837(.A1(new_n749), .A2(new_n203), .ZN(new_n1038));
  NOR4_X1   g0838(.A1(new_n1031), .A2(new_n1037), .A3(new_n1001), .A4(new_n1038), .ZN(new_n1039));
  NOR2_X1   g0839(.A1(new_n754), .A2(new_n564), .ZN(new_n1040));
  INV_X1    g0840(.A(G322), .ZN(new_n1041));
  OAI22_X1  g0841(.A1(new_n760), .A2(new_n1041), .B1(new_n750), .B2(new_n738), .ZN(new_n1042));
  XNOR2_X1  g0842(.A(new_n1042), .B(KEYINPUT112), .ZN(new_n1043));
  AOI22_X1  g0843(.A1(G303), .A2(new_n748), .B1(new_n752), .B2(G317), .ZN(new_n1044));
  NAND2_X1  g0844(.A1(new_n1043), .A2(new_n1044), .ZN(new_n1045));
  INV_X1    g0845(.A(KEYINPUT48), .ZN(new_n1046));
  NOR2_X1   g0846(.A1(new_n1045), .A2(new_n1046), .ZN(new_n1047));
  AOI211_X1 g0847(.A(new_n1040), .B(new_n1047), .C1(new_n768), .C2(new_n834), .ZN(new_n1048));
  OR2_X1    g0848(.A1(new_n1048), .A2(KEYINPUT113), .ZN(new_n1049));
  NAND2_X1  g0849(.A1(new_n1048), .A2(KEYINPUT113), .ZN(new_n1050));
  AOI22_X1  g0850(.A1(new_n1049), .A2(new_n1050), .B1(new_n1046), .B2(new_n1045), .ZN(new_n1051));
  XOR2_X1   g0851(.A(new_n1051), .B(KEYINPUT49), .Z(new_n1052));
  NOR2_X1   g0852(.A1(new_n744), .A2(new_n698), .ZN(new_n1053));
  AOI211_X1 g0853(.A(new_n261), .B(new_n1053), .C1(new_n762), .C2(new_n766), .ZN(new_n1054));
  AOI21_X1  g0854(.A(new_n1039), .B1(new_n1052), .B2(new_n1054), .ZN(new_n1055));
  OAI211_X1 g0855(.A(new_n802), .B(new_n1030), .C1(new_n1055), .C2(new_n1017), .ZN(new_n1056));
  INV_X1    g0856(.A(new_n987), .ZN(new_n1057));
  AOI21_X1  g0857(.A(new_n695), .B1(new_n986), .B2(new_n729), .ZN(new_n1058));
  NAND2_X1  g0858(.A1(new_n1057), .A2(new_n1058), .ZN(new_n1059));
  INV_X1    g0859(.A(new_n990), .ZN(new_n1060));
  OAI211_X1 g0860(.A(new_n1056), .B(new_n1059), .C1(new_n1060), .C2(new_n986), .ZN(G393));
  OAI22_X1  g0861(.A1(new_n760), .A2(new_n999), .B1(new_n750), .B2(new_n771), .ZN(new_n1062));
  XNOR2_X1  g0862(.A(new_n1062), .B(KEYINPUT52), .ZN(new_n1063));
  NAND2_X1  g0863(.A1(new_n775), .A2(G303), .ZN(new_n1064));
  AOI22_X1  g0864(.A1(new_n748), .A2(G294), .B1(G116), .B2(new_n768), .ZN(new_n1065));
  OAI22_X1  g0865(.A1(new_n996), .A2(new_n754), .B1(new_n744), .B2(new_n521), .ZN(new_n1066));
  AOI211_X1 g0866(.A(new_n261), .B(new_n1066), .C1(G322), .C2(new_n766), .ZN(new_n1067));
  NAND4_X1  g0867(.A1(new_n1063), .A2(new_n1064), .A3(new_n1065), .A4(new_n1067), .ZN(new_n1068));
  AOI211_X1 g0868(.A(new_n332), .B(new_n841), .C1(G143), .C2(new_n766), .ZN(new_n1069));
  OAI21_X1  g0869(.A(new_n1069), .B1(new_n203), .B2(new_n754), .ZN(new_n1070));
  XOR2_X1   g0870(.A(new_n1070), .B(KEYINPUT116), .Z(new_n1071));
  AOI22_X1  g0871(.A1(new_n775), .A2(new_n201), .B1(new_n768), .B2(G77), .ZN(new_n1072));
  OAI22_X1  g0872(.A1(new_n760), .A2(new_n278), .B1(new_n824), .B2(new_n771), .ZN(new_n1073));
  XNOR2_X1  g0873(.A(new_n1073), .B(KEYINPUT51), .ZN(new_n1074));
  NAND3_X1  g0874(.A1(new_n1071), .A2(new_n1072), .A3(new_n1074), .ZN(new_n1075));
  NOR2_X1   g0875(.A1(new_n749), .A2(new_n281), .ZN(new_n1076));
  OAI21_X1  g0876(.A(new_n1068), .B1(new_n1075), .B2(new_n1076), .ZN(new_n1077));
  AND2_X1   g0877(.A1(new_n1077), .A2(new_n786), .ZN(new_n1078));
  OAI221_X1 g0878(.A(new_n790), .B1(new_n484), .B2(new_n226), .C1(new_n245), .C2(new_n992), .ZN(new_n1079));
  NAND2_X1  g0879(.A1(new_n1079), .A2(new_n802), .ZN(new_n1080));
  XOR2_X1   g0880(.A(new_n1080), .B(KEYINPUT115), .Z(new_n1081));
  AOI211_X1 g0881(.A(new_n1078), .B(new_n1081), .C1(new_n960), .C2(new_n789), .ZN(new_n1082));
  INV_X1    g0882(.A(new_n983), .ZN(new_n1083));
  AOI21_X1  g0883(.A(new_n683), .B1(new_n980), .B2(new_n982), .ZN(new_n1084));
  OAI21_X1  g0884(.A(new_n1057), .B1(new_n1083), .B2(new_n1084), .ZN(new_n1085));
  AOI21_X1  g0885(.A(new_n695), .B1(new_n983), .B2(new_n987), .ZN(new_n1086));
  AOI21_X1  g0886(.A(new_n1082), .B1(new_n1085), .B2(new_n1086), .ZN(new_n1087));
  INV_X1    g0887(.A(KEYINPUT114), .ZN(new_n1088));
  OAI21_X1  g0888(.A(new_n1088), .B1(new_n1083), .B2(new_n1084), .ZN(new_n1089));
  INV_X1    g0889(.A(new_n1084), .ZN(new_n1090));
  NAND3_X1  g0890(.A1(new_n1090), .A2(KEYINPUT114), .A3(new_n983), .ZN(new_n1091));
  NAND3_X1  g0891(.A1(new_n1089), .A2(new_n1091), .A3(new_n990), .ZN(new_n1092));
  NAND2_X1  g0892(.A1(new_n1087), .A2(new_n1092), .ZN(G390));
  OAI22_X1  g0893(.A1(new_n936), .A2(new_n940), .B1(new_n933), .B2(new_n935), .ZN(new_n1094));
  NAND4_X1  g0894(.A1(new_n727), .A2(G330), .A3(new_n884), .A4(new_n883), .ZN(new_n1095));
  INV_X1    g0895(.A(new_n1095), .ZN(new_n1096));
  INV_X1    g0896(.A(new_n864), .ZN(new_n1097));
  NOR3_X1   g0897(.A1(new_n1097), .A2(new_n911), .A3(new_n909), .ZN(new_n1098));
  OAI21_X1  g0898(.A(new_n859), .B1(new_n1098), .B2(new_n858), .ZN(new_n1099));
  AOI21_X1  g0899(.A(KEYINPUT38), .B1(new_n1099), .B2(new_n910), .ZN(new_n1100));
  OAI21_X1  g0900(.A(new_n937), .B1(new_n1100), .B2(new_n899), .ZN(new_n1101));
  NAND3_X1  g0901(.A1(new_n639), .A2(new_n708), .A3(new_n641), .ZN(new_n1102));
  NAND3_X1  g0902(.A1(new_n1102), .A2(new_n884), .A3(new_n684), .ZN(new_n1103));
  AOI21_X1  g0903(.A(new_n896), .B1(new_n1103), .B2(new_n812), .ZN(new_n1104));
  INV_X1    g0904(.A(KEYINPUT117), .ZN(new_n1105));
  NOR3_X1   g0905(.A1(new_n1101), .A2(new_n1104), .A3(new_n1105), .ZN(new_n1106));
  NAND2_X1  g0906(.A1(new_n1103), .A2(new_n812), .ZN(new_n1107));
  NAND2_X1  g0907(.A1(new_n1107), .A2(new_n883), .ZN(new_n1108));
  AOI21_X1  g0908(.A(new_n936), .B1(new_n868), .B2(new_n875), .ZN(new_n1109));
  AOI21_X1  g0909(.A(KEYINPUT117), .B1(new_n1108), .B2(new_n1109), .ZN(new_n1110));
  OAI211_X1 g0910(.A(new_n1094), .B(new_n1096), .C1(new_n1106), .C2(new_n1110), .ZN(new_n1111));
  OAI21_X1  g0911(.A(new_n1105), .B1(new_n1101), .B2(new_n1104), .ZN(new_n1112));
  NAND3_X1  g0912(.A1(new_n1108), .A2(KEYINPUT117), .A3(new_n1109), .ZN(new_n1113));
  OR2_X1    g0913(.A1(new_n940), .A2(new_n936), .ZN(new_n1114));
  OAI21_X1  g0914(.A(new_n942), .B1(new_n915), .B2(KEYINPUT39), .ZN(new_n1115));
  AOI22_X1  g0915(.A1(new_n1112), .A2(new_n1113), .B1(new_n1114), .B2(new_n1115), .ZN(new_n1116));
  NAND3_X1  g0916(.A1(new_n852), .A2(G330), .A3(new_n897), .ZN(new_n1117));
  INV_X1    g0917(.A(new_n1117), .ZN(new_n1118));
  OAI21_X1  g0918(.A(new_n1111), .B1(new_n1116), .B2(new_n1118), .ZN(new_n1119));
  NAND3_X1  g0919(.A1(new_n727), .A2(G330), .A3(new_n884), .ZN(new_n1120));
  NAND2_X1  g0920(.A1(new_n1120), .A2(new_n896), .ZN(new_n1121));
  NAND2_X1  g0921(.A1(new_n1121), .A2(new_n1117), .ZN(new_n1122));
  AOI21_X1  g0922(.A(new_n809), .B1(new_n709), .B2(new_n884), .ZN(new_n1123));
  AND2_X1   g0923(.A1(new_n1095), .A2(new_n1123), .ZN(new_n1124));
  NAND3_X1  g0924(.A1(new_n852), .A2(G330), .A3(new_n884), .ZN(new_n1125));
  NAND2_X1  g0925(.A1(new_n1125), .A2(new_n896), .ZN(new_n1126));
  AOI22_X1  g0926(.A1(new_n926), .A2(new_n1122), .B1(new_n1124), .B2(new_n1126), .ZN(new_n1127));
  NAND3_X1  g0927(.A1(new_n667), .A2(new_n922), .A3(new_n853), .ZN(new_n1128));
  NOR3_X1   g0928(.A1(new_n1127), .A2(KEYINPUT118), .A3(new_n1128), .ZN(new_n1129));
  INV_X1    g0929(.A(KEYINPUT118), .ZN(new_n1130));
  NAND2_X1  g0930(.A1(new_n1122), .A2(new_n926), .ZN(new_n1131));
  NAND2_X1  g0931(.A1(new_n1124), .A2(new_n1126), .ZN(new_n1132));
  NAND2_X1  g0932(.A1(new_n1131), .A2(new_n1132), .ZN(new_n1133));
  AND3_X1   g0933(.A1(new_n667), .A2(new_n922), .A3(new_n853), .ZN(new_n1134));
  AOI21_X1  g0934(.A(new_n1130), .B1(new_n1133), .B2(new_n1134), .ZN(new_n1135));
  OAI21_X1  g0935(.A(new_n1119), .B1(new_n1129), .B2(new_n1135), .ZN(new_n1136));
  OAI21_X1  g0936(.A(KEYINPUT118), .B1(new_n1127), .B2(new_n1128), .ZN(new_n1137));
  OAI21_X1  g0937(.A(new_n1094), .B1(new_n1106), .B2(new_n1110), .ZN(new_n1138));
  NAND2_X1  g0938(.A1(new_n1138), .A2(new_n1117), .ZN(new_n1139));
  AND2_X1   g0939(.A1(new_n1124), .A2(new_n1126), .ZN(new_n1140));
  AOI22_X1  g0940(.A1(new_n1121), .A2(new_n1117), .B1(new_n812), .B2(new_n925), .ZN(new_n1141));
  OAI211_X1 g0941(.A(new_n1134), .B(new_n1130), .C1(new_n1140), .C2(new_n1141), .ZN(new_n1142));
  NAND4_X1  g0942(.A1(new_n1137), .A2(new_n1139), .A3(new_n1142), .A4(new_n1111), .ZN(new_n1143));
  NAND3_X1  g0943(.A1(new_n1136), .A2(new_n694), .A3(new_n1143), .ZN(new_n1144));
  NAND2_X1  g0944(.A1(new_n1119), .A2(new_n990), .ZN(new_n1145));
  NAND2_X1  g0945(.A1(new_n1115), .A2(new_n787), .ZN(new_n1146));
  NAND2_X1  g0946(.A1(new_n761), .A2(G283), .ZN(new_n1147));
  NAND2_X1  g0947(.A1(new_n748), .A2(G97), .ZN(new_n1148));
  AOI21_X1  g0948(.A(new_n261), .B1(new_n745), .B2(G68), .ZN(new_n1149));
  OAI22_X1  g0949(.A1(new_n738), .A2(new_n521), .B1(new_n765), .B2(new_n564), .ZN(new_n1150));
  AOI21_X1  g0950(.A(new_n1150), .B1(G116), .B2(new_n752), .ZN(new_n1151));
  NAND4_X1  g0951(.A1(new_n1147), .A2(new_n1148), .A3(new_n1149), .A4(new_n1151), .ZN(new_n1152));
  AOI211_X1 g0952(.A(new_n777), .B(new_n1152), .C1(G77), .C2(new_n768), .ZN(new_n1153));
  AOI22_X1  g0953(.A1(new_n761), .A2(G128), .B1(new_n201), .B2(new_n745), .ZN(new_n1154));
  OAI211_X1 g0954(.A(new_n1154), .B(new_n261), .C1(new_n825), .C2(new_n738), .ZN(new_n1155));
  NOR2_X1   g0955(.A1(new_n771), .A2(new_n830), .ZN(new_n1156));
  AOI22_X1  g0956(.A1(G125), .A2(new_n766), .B1(new_n768), .B2(G159), .ZN(new_n1157));
  XOR2_X1   g0957(.A(KEYINPUT54), .B(G143), .Z(new_n1158));
  INV_X1    g0958(.A(new_n1158), .ZN(new_n1159));
  OAI21_X1  g0959(.A(new_n1157), .B1(new_n749), .B2(new_n1159), .ZN(new_n1160));
  NOR2_X1   g0960(.A1(new_n754), .A2(new_n278), .ZN(new_n1161));
  XOR2_X1   g0961(.A(KEYINPUT119), .B(KEYINPUT53), .Z(new_n1162));
  XNOR2_X1  g0962(.A(new_n1161), .B(new_n1162), .ZN(new_n1163));
  NOR4_X1   g0963(.A1(new_n1155), .A2(new_n1156), .A3(new_n1160), .A4(new_n1163), .ZN(new_n1164));
  OAI21_X1  g0964(.A(new_n786), .B1(new_n1153), .B2(new_n1164), .ZN(new_n1165));
  NAND2_X1  g0965(.A1(new_n844), .A2(new_n281), .ZN(new_n1166));
  NAND4_X1  g0966(.A1(new_n1146), .A2(new_n802), .A3(new_n1165), .A4(new_n1166), .ZN(new_n1167));
  NAND3_X1  g0967(.A1(new_n1144), .A2(new_n1145), .A3(new_n1167), .ZN(G378));
  NAND2_X1  g0968(.A1(new_n1136), .A2(new_n1134), .ZN(new_n1169));
  AND3_X1   g0969(.A1(new_n941), .A2(new_n943), .A3(new_n944), .ZN(new_n1170));
  AOI21_X1  g0970(.A(new_n944), .B1(new_n941), .B2(new_n943), .ZN(new_n1171));
  NOR2_X1   g0971(.A1(new_n1170), .A2(new_n1171), .ZN(new_n1172));
  NAND2_X1  g0972(.A1(new_n294), .A2(new_n856), .ZN(new_n1173));
  INV_X1    g0973(.A(new_n1173), .ZN(new_n1174));
  AOI21_X1  g0974(.A(KEYINPUT121), .B1(new_n666), .B2(new_n297), .ZN(new_n1175));
  INV_X1    g0975(.A(KEYINPUT121), .ZN(new_n1176));
  AOI211_X1 g0976(.A(new_n1176), .B(new_n650), .C1(new_n665), .C2(new_n305), .ZN(new_n1177));
  OAI21_X1  g0977(.A(new_n1174), .B1(new_n1175), .B2(new_n1177), .ZN(new_n1178));
  NAND2_X1  g0978(.A1(new_n308), .A2(new_n1176), .ZN(new_n1179));
  NAND3_X1  g0979(.A1(new_n666), .A2(KEYINPUT121), .A3(new_n297), .ZN(new_n1180));
  NAND3_X1  g0980(.A1(new_n1179), .A2(new_n1173), .A3(new_n1180), .ZN(new_n1181));
  XOR2_X1   g0981(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1182));
  AND3_X1   g0982(.A1(new_n1178), .A2(new_n1181), .A3(new_n1182), .ZN(new_n1183));
  AOI21_X1  g0983(.A(new_n1182), .B1(new_n1178), .B2(new_n1181), .ZN(new_n1184));
  NOR2_X1   g0984(.A1(new_n1183), .A2(new_n1184), .ZN(new_n1185));
  INV_X1    g0985(.A(new_n1185), .ZN(new_n1186));
  AOI21_X1  g0986(.A(new_n1186), .B1(new_n919), .B2(G330), .ZN(new_n1187));
  AOI211_X1 g0987(.A(new_n905), .B(new_n1185), .C1(new_n916), .C2(new_n918), .ZN(new_n1188));
  OAI21_X1  g0988(.A(new_n1172), .B1(new_n1187), .B2(new_n1188), .ZN(new_n1189));
  OAI21_X1  g0989(.A(new_n1185), .B1(new_n904), .B2(new_n905), .ZN(new_n1190));
  NAND3_X1  g0990(.A1(new_n919), .A2(G330), .A3(new_n1186), .ZN(new_n1191));
  NAND3_X1  g0991(.A1(new_n1190), .A2(new_n946), .A3(new_n1191), .ZN(new_n1192));
  AND2_X1   g0992(.A1(new_n1189), .A2(new_n1192), .ZN(new_n1193));
  NAND3_X1  g0993(.A1(new_n1169), .A2(new_n1193), .A3(KEYINPUT57), .ZN(new_n1194));
  INV_X1    g0994(.A(KEYINPUT57), .ZN(new_n1195));
  NAND2_X1  g0995(.A1(new_n1137), .A2(new_n1142), .ZN(new_n1196));
  AOI21_X1  g0996(.A(new_n1128), .B1(new_n1196), .B2(new_n1119), .ZN(new_n1197));
  NAND2_X1  g0997(.A1(new_n1189), .A2(new_n1192), .ZN(new_n1198));
  OAI21_X1  g0998(.A(new_n1195), .B1(new_n1197), .B2(new_n1198), .ZN(new_n1199));
  NAND3_X1  g0999(.A1(new_n1194), .A2(new_n1199), .A3(new_n694), .ZN(new_n1200));
  AOI22_X1  g1000(.A1(new_n775), .A2(G97), .B1(new_n766), .B2(G283), .ZN(new_n1201));
  NAND2_X1  g1001(.A1(new_n745), .A2(G58), .ZN(new_n1202));
  NAND4_X1  g1002(.A1(new_n1201), .A2(new_n468), .A3(new_n332), .A4(new_n1202), .ZN(new_n1203));
  NOR2_X1   g1003(.A1(new_n1203), .A2(new_n1005), .ZN(new_n1204));
  OAI21_X1  g1004(.A(new_n1204), .B1(new_n396), .B2(new_n749), .ZN(new_n1205));
  AOI21_X1  g1005(.A(new_n1205), .B1(G77), .B2(new_n755), .ZN(new_n1206));
  OAI221_X1 g1006(.A(new_n1206), .B1(new_n521), .B2(new_n771), .C1(new_n698), .C2(new_n760), .ZN(new_n1207));
  INV_X1    g1007(.A(KEYINPUT58), .ZN(new_n1208));
  NAND2_X1  g1008(.A1(new_n1207), .A2(new_n1208), .ZN(new_n1209));
  OAI21_X1  g1009(.A(new_n292), .B1(new_n318), .B2(G41), .ZN(new_n1210));
  OR3_X1    g1010(.A1(new_n1159), .A2(KEYINPUT120), .A3(new_n754), .ZN(new_n1211));
  OAI21_X1  g1011(.A(KEYINPUT120), .B1(new_n1159), .B2(new_n754), .ZN(new_n1212));
  NAND2_X1  g1012(.A1(new_n752), .A2(G128), .ZN(new_n1213));
  NAND3_X1  g1013(.A1(new_n1211), .A2(new_n1212), .A3(new_n1213), .ZN(new_n1214));
  NAND2_X1  g1014(.A1(new_n761), .A2(G125), .ZN(new_n1215));
  OAI221_X1 g1015(.A(new_n1215), .B1(new_n830), .B2(new_n738), .C1(new_n278), .C2(new_n767), .ZN(new_n1216));
  AOI211_X1 g1016(.A(new_n1214), .B(new_n1216), .C1(G137), .C2(new_n748), .ZN(new_n1217));
  INV_X1    g1017(.A(KEYINPUT59), .ZN(new_n1218));
  AOI21_X1  g1018(.A(G33), .B1(new_n1217), .B2(new_n1218), .ZN(new_n1219));
  AOI21_X1  g1019(.A(G41), .B1(new_n766), .B2(G124), .ZN(new_n1220));
  OAI211_X1 g1020(.A(new_n1219), .B(new_n1220), .C1(new_n824), .C2(new_n744), .ZN(new_n1221));
  NOR2_X1   g1021(.A1(new_n1217), .A2(new_n1218), .ZN(new_n1222));
  OAI211_X1 g1022(.A(new_n1209), .B(new_n1210), .C1(new_n1221), .C2(new_n1222), .ZN(new_n1223));
  NOR2_X1   g1023(.A1(new_n1207), .A2(new_n1208), .ZN(new_n1224));
  NOR2_X1   g1024(.A1(new_n1223), .A2(new_n1224), .ZN(new_n1225));
  NOR2_X1   g1025(.A1(new_n1225), .A2(new_n1017), .ZN(new_n1226));
  NOR2_X1   g1026(.A1(new_n1185), .A2(new_n788), .ZN(new_n1227));
  AOI211_X1 g1027(.A(new_n1226), .B(new_n1227), .C1(new_n1013), .C2(new_n844), .ZN(new_n1228));
  NAND2_X1  g1028(.A1(new_n1228), .A2(new_n802), .ZN(new_n1229));
  OAI21_X1  g1029(.A(new_n1229), .B1(new_n1198), .B2(new_n1060), .ZN(new_n1230));
  INV_X1    g1030(.A(new_n1230), .ZN(new_n1231));
  NAND2_X1  g1031(.A1(new_n1200), .A2(new_n1231), .ZN(G375));
  NAND2_X1  g1032(.A1(new_n844), .A2(new_n203), .ZN(new_n1233));
  OAI21_X1  g1033(.A(new_n1233), .B1(new_n883), .B2(new_n788), .ZN(new_n1234));
  OAI21_X1  g1034(.A(new_n1202), .B1(new_n824), .B2(new_n754), .ZN(new_n1235));
  AOI211_X1 g1035(.A(new_n332), .B(new_n1235), .C1(G128), .C2(new_n766), .ZN(new_n1236));
  OAI22_X1  g1036(.A1(new_n749), .A2(new_n278), .B1(new_n771), .B2(new_n825), .ZN(new_n1237));
  AOI21_X1  g1037(.A(new_n1237), .B1(new_n775), .B2(new_n1158), .ZN(new_n1238));
  NAND2_X1  g1038(.A1(new_n768), .A2(G50), .ZN(new_n1239));
  NAND2_X1  g1039(.A1(new_n761), .A2(G132), .ZN(new_n1240));
  NAND4_X1  g1040(.A1(new_n1236), .A2(new_n1238), .A3(new_n1239), .A4(new_n1240), .ZN(new_n1241));
  OAI22_X1  g1041(.A1(new_n749), .A2(new_n521), .B1(new_n738), .B2(new_n698), .ZN(new_n1242));
  AOI21_X1  g1042(.A(new_n1242), .B1(G294), .B2(new_n761), .ZN(new_n1243));
  XOR2_X1   g1043(.A(new_n1243), .B(KEYINPUT123), .Z(new_n1244));
  NAND2_X1  g1044(.A1(new_n766), .A2(G303), .ZN(new_n1245));
  AOI211_X1 g1045(.A(new_n1032), .B(new_n1006), .C1(G283), .C2(new_n752), .ZN(new_n1246));
  NAND4_X1  g1046(.A1(new_n1244), .A2(new_n332), .A3(new_n1245), .A4(new_n1246), .ZN(new_n1247));
  NOR2_X1   g1047(.A1(new_n754), .A2(new_n484), .ZN(new_n1248));
  OAI21_X1  g1048(.A(new_n1241), .B1(new_n1247), .B2(new_n1248), .ZN(new_n1249));
  AOI211_X1 g1049(.A(new_n735), .B(new_n1234), .C1(new_n786), .C2(new_n1249), .ZN(new_n1250));
  AOI21_X1  g1050(.A(new_n1250), .B1(new_n1133), .B2(new_n990), .ZN(new_n1251));
  NAND3_X1  g1051(.A1(new_n1131), .A2(new_n1128), .A3(new_n1132), .ZN(new_n1252));
  NAND3_X1  g1052(.A1(new_n1137), .A2(new_n1142), .A3(new_n1252), .ZN(new_n1253));
  XOR2_X1   g1053(.A(new_n976), .B(KEYINPUT122), .Z(new_n1254));
  INV_X1    g1054(.A(new_n1254), .ZN(new_n1255));
  OAI21_X1  g1055(.A(new_n1251), .B1(new_n1253), .B2(new_n1255), .ZN(G381));
  AOI22_X1  g1056(.A1(new_n1142), .A2(new_n1137), .B1(new_n1139), .B2(new_n1111), .ZN(new_n1257));
  OAI211_X1 g1057(.A(new_n1192), .B(new_n1189), .C1(new_n1257), .C2(new_n1128), .ZN(new_n1258));
  AOI21_X1  g1058(.A(new_n695), .B1(new_n1258), .B2(new_n1195), .ZN(new_n1259));
  AOI21_X1  g1059(.A(new_n1230), .B1(new_n1259), .B2(new_n1194), .ZN(new_n1260));
  XNOR2_X1  g1060(.A(new_n1260), .B(KEYINPUT124), .ZN(new_n1261));
  INV_X1    g1061(.A(G384), .ZN(new_n1262));
  INV_X1    g1062(.A(G378), .ZN(new_n1263));
  NAND4_X1  g1063(.A1(new_n991), .A2(new_n1020), .A3(new_n1087), .A4(new_n1092), .ZN(new_n1264));
  NOR4_X1   g1064(.A1(new_n1264), .A2(G396), .A3(G393), .A4(G381), .ZN(new_n1265));
  NAND4_X1  g1065(.A1(new_n1261), .A2(new_n1262), .A3(new_n1263), .A4(new_n1265), .ZN(G407));
  NAND3_X1  g1066(.A1(new_n1261), .A2(new_n676), .A3(new_n1263), .ZN(new_n1267));
  NAND3_X1  g1067(.A1(G407), .A2(G213), .A3(new_n1267), .ZN(G409));
  NAND2_X1  g1068(.A1(G387), .A2(G390), .ZN(new_n1269));
  NAND2_X1  g1069(.A1(new_n1269), .A2(new_n1264), .ZN(new_n1270));
  XNOR2_X1  g1070(.A(G393), .B(G396), .ZN(new_n1271));
  INV_X1    g1071(.A(new_n1271), .ZN(new_n1272));
  NAND2_X1  g1072(.A1(new_n1270), .A2(new_n1272), .ZN(new_n1273));
  NAND3_X1  g1073(.A1(new_n1269), .A2(new_n1264), .A3(new_n1271), .ZN(new_n1274));
  NAND2_X1  g1074(.A1(new_n1273), .A2(new_n1274), .ZN(new_n1275));
  INV_X1    g1075(.A(G213), .ZN(new_n1276));
  NOR2_X1   g1076(.A1(new_n1276), .A2(G343), .ZN(new_n1277));
  NAND2_X1  g1077(.A1(new_n1277), .A2(G2897), .ZN(new_n1278));
  INV_X1    g1078(.A(new_n1278), .ZN(new_n1279));
  NAND2_X1  g1079(.A1(new_n1253), .A2(KEYINPUT60), .ZN(new_n1280));
  INV_X1    g1080(.A(KEYINPUT60), .ZN(new_n1281));
  NAND2_X1  g1081(.A1(new_n1252), .A2(new_n1281), .ZN(new_n1282));
  NAND2_X1  g1082(.A1(new_n1282), .A2(new_n694), .ZN(new_n1283));
  INV_X1    g1083(.A(new_n1283), .ZN(new_n1284));
  NAND2_X1  g1084(.A1(new_n1280), .A2(new_n1284), .ZN(new_n1285));
  INV_X1    g1085(.A(KEYINPUT125), .ZN(new_n1286));
  NAND2_X1  g1086(.A1(new_n1285), .A2(new_n1286), .ZN(new_n1287));
  NAND3_X1  g1087(.A1(new_n1280), .A2(KEYINPUT125), .A3(new_n1284), .ZN(new_n1288));
  NAND2_X1  g1088(.A1(new_n1287), .A2(new_n1288), .ZN(new_n1289));
  AOI21_X1  g1089(.A(G384), .B1(new_n1289), .B2(new_n1251), .ZN(new_n1290));
  AOI211_X1 g1090(.A(new_n1286), .B(new_n1283), .C1(KEYINPUT60), .C2(new_n1253), .ZN(new_n1291));
  AOI21_X1  g1091(.A(KEYINPUT125), .B1(new_n1280), .B2(new_n1284), .ZN(new_n1292));
  OAI211_X1 g1092(.A(G384), .B(new_n1251), .C1(new_n1291), .C2(new_n1292), .ZN(new_n1293));
  INV_X1    g1093(.A(new_n1293), .ZN(new_n1294));
  OAI21_X1  g1094(.A(new_n1279), .B1(new_n1290), .B2(new_n1294), .ZN(new_n1295));
  OAI21_X1  g1095(.A(new_n1251), .B1(new_n1291), .B2(new_n1292), .ZN(new_n1296));
  NAND2_X1  g1096(.A1(new_n1296), .A2(new_n1262), .ZN(new_n1297));
  NAND3_X1  g1097(.A1(new_n1297), .A2(new_n1293), .A3(new_n1278), .ZN(new_n1298));
  NAND3_X1  g1098(.A1(new_n1169), .A2(new_n1193), .A3(new_n1254), .ZN(new_n1299));
  AOI21_X1  g1099(.A(G378), .B1(new_n1231), .B2(new_n1299), .ZN(new_n1300));
  AOI21_X1  g1100(.A(new_n1300), .B1(new_n1260), .B2(G378), .ZN(new_n1301));
  OAI211_X1 g1101(.A(new_n1295), .B(new_n1298), .C1(new_n1301), .C2(new_n1277), .ZN(new_n1302));
  NOR2_X1   g1102(.A1(new_n1290), .A2(new_n1294), .ZN(new_n1303));
  INV_X1    g1103(.A(new_n1277), .ZN(new_n1304));
  NAND3_X1  g1104(.A1(new_n1200), .A2(G378), .A3(new_n1231), .ZN(new_n1305));
  NAND2_X1  g1105(.A1(new_n1231), .A2(new_n1299), .ZN(new_n1306));
  NAND2_X1  g1106(.A1(new_n1306), .A2(new_n1263), .ZN(new_n1307));
  NAND2_X1  g1107(.A1(new_n1305), .A2(new_n1307), .ZN(new_n1308));
  NAND3_X1  g1108(.A1(new_n1303), .A2(new_n1304), .A3(new_n1308), .ZN(new_n1309));
  AOI21_X1  g1109(.A(KEYINPUT62), .B1(new_n1302), .B2(new_n1309), .ZN(new_n1310));
  NAND2_X1  g1110(.A1(new_n1309), .A2(KEYINPUT62), .ZN(new_n1311));
  INV_X1    g1111(.A(KEYINPUT61), .ZN(new_n1312));
  NAND2_X1  g1112(.A1(new_n1311), .A2(new_n1312), .ZN(new_n1313));
  OAI21_X1  g1113(.A(new_n1275), .B1(new_n1310), .B2(new_n1313), .ZN(new_n1314));
  NAND2_X1  g1114(.A1(new_n1295), .A2(new_n1298), .ZN(new_n1315));
  AOI21_X1  g1115(.A(new_n1277), .B1(new_n1305), .B2(new_n1307), .ZN(new_n1316));
  OAI21_X1  g1116(.A(new_n1309), .B1(new_n1315), .B2(new_n1316), .ZN(new_n1317));
  NAND2_X1  g1117(.A1(new_n1317), .A2(KEYINPUT63), .ZN(new_n1318));
  AOI21_X1  g1118(.A(KEYINPUT63), .B1(new_n1316), .B2(new_n1303), .ZN(new_n1319));
  NOR3_X1   g1119(.A1(new_n1319), .A2(new_n1275), .A3(KEYINPUT61), .ZN(new_n1320));
  NAND2_X1  g1120(.A1(new_n1318), .A2(new_n1320), .ZN(new_n1321));
  NAND2_X1  g1121(.A1(new_n1314), .A2(new_n1321), .ZN(G405));
  INV_X1    g1122(.A(KEYINPUT127), .ZN(new_n1323));
  NAND2_X1  g1123(.A1(G375), .A2(new_n1263), .ZN(new_n1324));
  NAND2_X1  g1124(.A1(new_n1324), .A2(new_n1305), .ZN(new_n1325));
  INV_X1    g1125(.A(new_n1325), .ZN(new_n1326));
  INV_X1    g1126(.A(KEYINPUT126), .ZN(new_n1327));
  OAI21_X1  g1127(.A(new_n1327), .B1(new_n1290), .B2(new_n1294), .ZN(new_n1328));
  NAND2_X1  g1128(.A1(new_n1303), .A2(KEYINPUT126), .ZN(new_n1329));
  AOI21_X1  g1129(.A(new_n1326), .B1(new_n1328), .B2(new_n1329), .ZN(new_n1330));
  AOI21_X1  g1130(.A(new_n1325), .B1(KEYINPUT126), .B2(new_n1303), .ZN(new_n1331));
  OAI211_X1 g1131(.A(new_n1275), .B(new_n1323), .C1(new_n1330), .C2(new_n1331), .ZN(new_n1332));
  NAND2_X1  g1132(.A1(new_n1329), .A2(new_n1328), .ZN(new_n1333));
  NAND2_X1  g1133(.A1(new_n1333), .A2(new_n1325), .ZN(new_n1334));
  NAND2_X1  g1134(.A1(new_n1275), .A2(new_n1323), .ZN(new_n1335));
  NAND3_X1  g1135(.A1(new_n1273), .A2(KEYINPUT127), .A3(new_n1274), .ZN(new_n1336));
  NAND2_X1  g1136(.A1(new_n1326), .A2(new_n1329), .ZN(new_n1337));
  NAND4_X1  g1137(.A1(new_n1334), .A2(new_n1335), .A3(new_n1336), .A4(new_n1337), .ZN(new_n1338));
  NAND2_X1  g1138(.A1(new_n1332), .A2(new_n1338), .ZN(G402));
endmodule


