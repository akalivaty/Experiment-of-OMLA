//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 0 1 1 1 1 0 0 1 0 1 1 0 1 1 1 1 1 0 1 1 1 0 1 1 1 1 0 0 0 1 1 0 0 1 1 1 0 1 1 0 0 0 0 1 0 0 0 0 1 1 1 1 0 0 1 0 0 0 0 0 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:39:33 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1234, new_n1236,
    new_n1237, new_n1238, new_n1239, new_n1240, new_n1241, new_n1242,
    new_n1243, new_n1244, new_n1246, new_n1247, new_n1248, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1308, new_n1309, new_n1310, new_n1311,
    new_n1312, new_n1313, new_n1314, new_n1315, new_n1316, new_n1317,
    new_n1318;
  INV_X1    g0000(.A(G50), .ZN(new_n201));
  INV_X1    g0001(.A(G58), .ZN(new_n202));
  INV_X1    g0002(.A(G68), .ZN(new_n203));
  NAND3_X1  g0003(.A1(new_n201), .A2(new_n202), .A3(new_n203), .ZN(new_n204));
  NOR2_X1   g0004(.A1(new_n204), .A2(G77), .ZN(G353));
  OAI21_X1  g0005(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0006(.A(G1), .ZN(new_n207));
  INV_X1    g0007(.A(G20), .ZN(new_n208));
  NOR2_X1   g0008(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  INV_X1    g0009(.A(new_n209), .ZN(new_n210));
  NOR2_X1   g0010(.A1(new_n210), .A2(G13), .ZN(new_n211));
  OAI211_X1 g0011(.A(new_n211), .B(G250), .C1(G257), .C2(G264), .ZN(new_n212));
  XNOR2_X1  g0012(.A(KEYINPUT64), .B(KEYINPUT0), .ZN(new_n213));
  XNOR2_X1  g0013(.A(new_n212), .B(new_n213), .ZN(new_n214));
  NAND2_X1  g0014(.A1(G1), .A2(G13), .ZN(new_n215));
  NOR2_X1   g0015(.A1(new_n215), .A2(new_n208), .ZN(new_n216));
  OAI21_X1  g0016(.A(G50), .B1(G58), .B2(G68), .ZN(new_n217));
  INV_X1    g0017(.A(new_n217), .ZN(new_n218));
  AOI21_X1  g0018(.A(new_n214), .B1(new_n216), .B2(new_n218), .ZN(new_n219));
  AOI22_X1  g0019(.A1(G107), .A2(G264), .B1(G116), .B2(G270), .ZN(new_n220));
  INV_X1    g0020(.A(G77), .ZN(new_n221));
  INV_X1    g0021(.A(G244), .ZN(new_n222));
  INV_X1    g0022(.A(G87), .ZN(new_n223));
  INV_X1    g0023(.A(G250), .ZN(new_n224));
  OAI221_X1 g0024(.A(new_n220), .B1(new_n221), .B2(new_n222), .C1(new_n223), .C2(new_n224), .ZN(new_n225));
  AOI22_X1  g0025(.A1(G50), .A2(G226), .B1(G97), .B2(G257), .ZN(new_n226));
  INV_X1    g0026(.A(G232), .ZN(new_n227));
  INV_X1    g0027(.A(G238), .ZN(new_n228));
  OAI221_X1 g0028(.A(new_n226), .B1(new_n202), .B2(new_n227), .C1(new_n203), .C2(new_n228), .ZN(new_n229));
  OAI21_X1  g0029(.A(new_n210), .B1(new_n225), .B2(new_n229), .ZN(new_n230));
  OR2_X1    g0030(.A1(new_n230), .A2(KEYINPUT1), .ZN(new_n231));
  NAND2_X1  g0031(.A1(new_n230), .A2(KEYINPUT1), .ZN(new_n232));
  AND3_X1   g0032(.A1(new_n219), .A2(new_n231), .A3(new_n232), .ZN(G361));
  XNOR2_X1  g0033(.A(G238), .B(G244), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n234), .B(KEYINPUT2), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n235), .B(G226), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n236), .B(new_n227), .ZN(new_n237));
  XNOR2_X1  g0037(.A(G250), .B(G257), .ZN(new_n238));
  XNOR2_X1  g0038(.A(G264), .B(G270), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n237), .B(new_n240), .ZN(G358));
  XOR2_X1   g0041(.A(G68), .B(G77), .Z(new_n242));
  XNOR2_X1  g0042(.A(G50), .B(G58), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XOR2_X1   g0044(.A(G87), .B(G97), .Z(new_n245));
  XNOR2_X1  g0045(.A(G107), .B(G116), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n245), .B(new_n246), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n244), .B(new_n247), .ZN(G351));
  INV_X1    g0048(.A(KEYINPUT73), .ZN(new_n249));
  AND2_X1   g0049(.A1(KEYINPUT3), .A2(G33), .ZN(new_n250));
  NOR2_X1   g0050(.A1(KEYINPUT3), .A2(G33), .ZN(new_n251));
  NOR2_X1   g0051(.A1(new_n250), .A2(new_n251), .ZN(new_n252));
  AOI21_X1  g0052(.A(KEYINPUT7), .B1(new_n252), .B2(new_n208), .ZN(new_n253));
  OR2_X1    g0053(.A1(KEYINPUT3), .A2(G33), .ZN(new_n254));
  NAND2_X1  g0054(.A1(KEYINPUT3), .A2(G33), .ZN(new_n255));
  NAND4_X1  g0055(.A1(new_n254), .A2(KEYINPUT7), .A3(new_n208), .A4(new_n255), .ZN(new_n256));
  INV_X1    g0056(.A(new_n256), .ZN(new_n257));
  OAI21_X1  g0057(.A(G68), .B1(new_n253), .B2(new_n257), .ZN(new_n258));
  AND2_X1   g0058(.A1(G58), .A2(G68), .ZN(new_n259));
  NOR2_X1   g0059(.A1(G58), .A2(G68), .ZN(new_n260));
  OAI21_X1  g0060(.A(G20), .B1(new_n259), .B2(new_n260), .ZN(new_n261));
  NOR2_X1   g0061(.A1(G20), .A2(G33), .ZN(new_n262));
  AND3_X1   g0062(.A1(new_n262), .A2(KEYINPUT71), .A3(G159), .ZN(new_n263));
  AOI21_X1  g0063(.A(KEYINPUT71), .B1(new_n262), .B2(G159), .ZN(new_n264));
  OAI21_X1  g0064(.A(new_n261), .B1(new_n263), .B2(new_n264), .ZN(new_n265));
  INV_X1    g0065(.A(new_n265), .ZN(new_n266));
  AOI21_X1  g0066(.A(KEYINPUT16), .B1(new_n258), .B2(new_n266), .ZN(new_n267));
  NAND3_X1  g0067(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n268));
  NAND2_X1  g0068(.A1(new_n268), .A2(new_n215), .ZN(new_n269));
  NAND3_X1  g0069(.A1(new_n254), .A2(new_n208), .A3(new_n255), .ZN(new_n270));
  INV_X1    g0070(.A(KEYINPUT7), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n270), .A2(new_n271), .ZN(new_n272));
  AOI21_X1  g0072(.A(new_n203), .B1(new_n272), .B2(new_n256), .ZN(new_n273));
  OAI211_X1 g0073(.A(KEYINPUT16), .B(new_n261), .C1(new_n263), .C2(new_n264), .ZN(new_n274));
  OAI21_X1  g0074(.A(new_n269), .B1(new_n273), .B2(new_n274), .ZN(new_n275));
  NOR2_X1   g0075(.A1(new_n267), .A2(new_n275), .ZN(new_n276));
  INV_X1    g0076(.A(KEYINPUT66), .ZN(new_n277));
  OAI21_X1  g0077(.A(new_n277), .B1(new_n208), .B2(G1), .ZN(new_n278));
  NAND3_X1  g0078(.A1(new_n207), .A2(KEYINPUT66), .A3(G20), .ZN(new_n279));
  NAND2_X1  g0079(.A1(new_n278), .A2(new_n279), .ZN(new_n280));
  AND2_X1   g0080(.A1(new_n268), .A2(new_n215), .ZN(new_n281));
  NAND3_X1  g0081(.A1(new_n207), .A2(G13), .A3(G20), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n202), .A2(KEYINPUT8), .ZN(new_n283));
  INV_X1    g0083(.A(KEYINPUT8), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n284), .A2(G58), .ZN(new_n285));
  NAND2_X1  g0085(.A1(new_n283), .A2(new_n285), .ZN(new_n286));
  NAND4_X1  g0086(.A1(new_n280), .A2(new_n281), .A3(new_n282), .A4(new_n286), .ZN(new_n287));
  XNOR2_X1  g0087(.A(KEYINPUT8), .B(G58), .ZN(new_n288));
  INV_X1    g0088(.A(new_n282), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n288), .A2(new_n289), .ZN(new_n290));
  NAND2_X1  g0090(.A1(new_n287), .A2(new_n290), .ZN(new_n291));
  INV_X1    g0091(.A(KEYINPUT72), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n291), .A2(new_n292), .ZN(new_n293));
  NAND3_X1  g0093(.A1(new_n287), .A2(KEYINPUT72), .A3(new_n290), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n293), .A2(new_n294), .ZN(new_n295));
  OAI21_X1  g0095(.A(new_n249), .B1(new_n276), .B2(new_n295), .ZN(new_n296));
  INV_X1    g0096(.A(new_n274), .ZN(new_n297));
  AOI21_X1  g0097(.A(new_n281), .B1(new_n258), .B2(new_n297), .ZN(new_n298));
  INV_X1    g0098(.A(KEYINPUT16), .ZN(new_n299));
  OAI21_X1  g0099(.A(new_n299), .B1(new_n273), .B2(new_n265), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n298), .A2(new_n300), .ZN(new_n301));
  AND3_X1   g0101(.A1(new_n287), .A2(KEYINPUT72), .A3(new_n290), .ZN(new_n302));
  AOI21_X1  g0102(.A(KEYINPUT72), .B1(new_n287), .B2(new_n290), .ZN(new_n303));
  NOR2_X1   g0103(.A1(new_n302), .A2(new_n303), .ZN(new_n304));
  NAND3_X1  g0104(.A1(new_n301), .A2(KEYINPUT73), .A3(new_n304), .ZN(new_n305));
  OR2_X1    g0105(.A1(G223), .A2(G1698), .ZN(new_n306));
  INV_X1    g0106(.A(G226), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n307), .A2(G1698), .ZN(new_n308));
  OAI211_X1 g0108(.A(new_n306), .B(new_n308), .C1(new_n250), .C2(new_n251), .ZN(new_n309));
  NAND2_X1  g0109(.A1(G33), .A2(G87), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n309), .A2(new_n310), .ZN(new_n311));
  AOI21_X1  g0111(.A(new_n215), .B1(G33), .B2(G41), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n311), .A2(new_n312), .ZN(new_n313));
  INV_X1    g0113(.A(G41), .ZN(new_n314));
  INV_X1    g0114(.A(G45), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n314), .A2(new_n315), .ZN(new_n316));
  AND2_X1   g0116(.A1(G1), .A2(G13), .ZN(new_n317));
  NAND2_X1  g0117(.A1(G33), .A2(G41), .ZN(new_n318));
  AOI22_X1  g0118(.A1(new_n207), .A2(new_n316), .B1(new_n317), .B2(new_n318), .ZN(new_n319));
  OR2_X1    g0119(.A1(KEYINPUT65), .A2(G41), .ZN(new_n320));
  NAND2_X1  g0120(.A1(KEYINPUT65), .A2(G41), .ZN(new_n321));
  NAND3_X1  g0121(.A1(new_n320), .A2(new_n315), .A3(new_n321), .ZN(new_n322));
  INV_X1    g0122(.A(G274), .ZN(new_n323));
  NOR2_X1   g0123(.A1(new_n323), .A2(G1), .ZN(new_n324));
  AOI22_X1  g0124(.A1(new_n319), .A2(G232), .B1(new_n322), .B2(new_n324), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n313), .A2(new_n325), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n326), .A2(G169), .ZN(new_n327));
  INV_X1    g0127(.A(G179), .ZN(new_n328));
  OAI21_X1  g0128(.A(new_n327), .B1(new_n328), .B2(new_n326), .ZN(new_n329));
  NAND3_X1  g0129(.A1(new_n296), .A2(new_n305), .A3(new_n329), .ZN(new_n330));
  INV_X1    g0130(.A(KEYINPUT18), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n330), .A2(new_n331), .ZN(new_n332));
  NAND4_X1  g0132(.A1(new_n296), .A2(KEYINPUT18), .A3(new_n305), .A4(new_n329), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n332), .A2(new_n333), .ZN(new_n334));
  INV_X1    g0134(.A(KEYINPUT17), .ZN(new_n335));
  INV_X1    g0135(.A(G190), .ZN(new_n336));
  NAND3_X1  g0136(.A1(new_n313), .A2(new_n336), .A3(new_n325), .ZN(new_n337));
  INV_X1    g0137(.A(G200), .ZN(new_n338));
  NAND3_X1  g0138(.A1(new_n318), .A2(G1), .A3(G13), .ZN(new_n339));
  AOI21_X1  g0139(.A(new_n339), .B1(new_n309), .B2(new_n310), .ZN(new_n340));
  OAI21_X1  g0140(.A(new_n207), .B1(G41), .B2(G45), .ZN(new_n341));
  NAND3_X1  g0141(.A1(new_n339), .A2(G232), .A3(new_n341), .ZN(new_n342));
  AND2_X1   g0142(.A1(KEYINPUT65), .A2(G41), .ZN(new_n343));
  NOR2_X1   g0143(.A1(KEYINPUT65), .A2(G41), .ZN(new_n344));
  NOR3_X1   g0144(.A1(new_n343), .A2(new_n344), .A3(G45), .ZN(new_n345));
  INV_X1    g0145(.A(new_n324), .ZN(new_n346));
  OAI21_X1  g0146(.A(new_n342), .B1(new_n345), .B2(new_n346), .ZN(new_n347));
  OAI21_X1  g0147(.A(new_n338), .B1(new_n340), .B2(new_n347), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n337), .A2(new_n348), .ZN(new_n349));
  OAI211_X1 g0149(.A(new_n349), .B(new_n304), .C1(new_n267), .C2(new_n275), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n350), .A2(KEYINPUT74), .ZN(new_n351));
  INV_X1    g0151(.A(KEYINPUT74), .ZN(new_n352));
  NAND4_X1  g0152(.A1(new_n301), .A2(new_n352), .A3(new_n304), .A4(new_n349), .ZN(new_n353));
  AOI21_X1  g0153(.A(new_n335), .B1(new_n351), .B2(new_n353), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n350), .A2(new_n335), .ZN(new_n355));
  INV_X1    g0155(.A(new_n355), .ZN(new_n356));
  NOR2_X1   g0156(.A1(new_n354), .A2(new_n356), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n334), .A2(new_n357), .ZN(new_n358));
  NOR2_X1   g0158(.A1(new_n289), .A2(new_n269), .ZN(new_n359));
  AOI21_X1  g0159(.A(new_n201), .B1(new_n278), .B2(new_n279), .ZN(new_n360));
  INV_X1    g0160(.A(KEYINPUT67), .ZN(new_n361));
  OAI21_X1  g0161(.A(new_n359), .B1(new_n360), .B2(new_n361), .ZN(new_n362));
  AND2_X1   g0162(.A1(new_n360), .A2(new_n361), .ZN(new_n363));
  OR2_X1    g0163(.A1(new_n362), .A2(new_n363), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n204), .A2(G20), .ZN(new_n365));
  INV_X1    g0165(.A(G150), .ZN(new_n366));
  INV_X1    g0166(.A(G33), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n208), .A2(new_n367), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n208), .A2(G33), .ZN(new_n369));
  OAI221_X1 g0169(.A(new_n365), .B1(new_n366), .B2(new_n368), .C1(new_n369), .C2(new_n288), .ZN(new_n370));
  AOI22_X1  g0170(.A1(new_n370), .A2(new_n269), .B1(new_n201), .B2(new_n289), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n364), .A2(new_n371), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n372), .A2(KEYINPUT9), .ZN(new_n373));
  INV_X1    g0173(.A(KEYINPUT9), .ZN(new_n374));
  NAND3_X1  g0174(.A1(new_n364), .A2(new_n371), .A3(new_n374), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n254), .A2(new_n255), .ZN(new_n376));
  INV_X1    g0176(.A(G1698), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n377), .A2(G222), .ZN(new_n378));
  NAND2_X1  g0178(.A1(G223), .A2(G1698), .ZN(new_n379));
  NAND3_X1  g0179(.A1(new_n376), .A2(new_n378), .A3(new_n379), .ZN(new_n380));
  OAI211_X1 g0180(.A(new_n380), .B(new_n312), .C1(G77), .C2(new_n376), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n322), .A2(new_n324), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n319), .A2(G226), .ZN(new_n383));
  NAND3_X1  g0183(.A1(new_n381), .A2(new_n382), .A3(new_n383), .ZN(new_n384));
  INV_X1    g0184(.A(new_n384), .ZN(new_n385));
  AOI22_X1  g0185(.A1(new_n373), .A2(new_n375), .B1(G190), .B2(new_n385), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n384), .A2(G200), .ZN(new_n387));
  INV_X1    g0187(.A(KEYINPUT68), .ZN(new_n388));
  OAI211_X1 g0188(.A(new_n386), .B(new_n387), .C1(new_n388), .C2(KEYINPUT10), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n385), .A2(G190), .ZN(new_n390));
  INV_X1    g0190(.A(new_n375), .ZN(new_n391));
  AOI21_X1  g0191(.A(new_n374), .B1(new_n364), .B2(new_n371), .ZN(new_n392));
  OAI211_X1 g0192(.A(new_n390), .B(new_n387), .C1(new_n391), .C2(new_n392), .ZN(new_n393));
  OAI211_X1 g0193(.A(new_n390), .B(new_n388), .C1(new_n391), .C2(new_n392), .ZN(new_n394));
  INV_X1    g0194(.A(KEYINPUT10), .ZN(new_n395));
  NAND3_X1  g0195(.A1(new_n393), .A2(new_n394), .A3(new_n395), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n389), .A2(new_n396), .ZN(new_n397));
  INV_X1    g0197(.A(G169), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n384), .A2(new_n398), .ZN(new_n399));
  OAI21_X1  g0199(.A(new_n399), .B1(G179), .B2(new_n384), .ZN(new_n400));
  INV_X1    g0200(.A(new_n372), .ZN(new_n401));
  OR2_X1    g0201(.A1(new_n400), .A2(new_n401), .ZN(new_n402));
  INV_X1    g0202(.A(new_n402), .ZN(new_n403));
  NOR3_X1   g0203(.A1(new_n358), .A2(new_n397), .A3(new_n403), .ZN(new_n404));
  OAI22_X1  g0204(.A1(new_n369), .A2(new_n221), .B1(new_n208), .B2(G68), .ZN(new_n405));
  NOR2_X1   g0205(.A1(new_n368), .A2(new_n201), .ZN(new_n406));
  OAI21_X1  g0206(.A(new_n269), .B1(new_n405), .B2(new_n406), .ZN(new_n407));
  XNOR2_X1  g0207(.A(new_n407), .B(KEYINPUT11), .ZN(new_n408));
  INV_X1    g0208(.A(KEYINPUT70), .ZN(new_n409));
  OR2_X1    g0209(.A1(new_n408), .A2(new_n409), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n408), .A2(new_n409), .ZN(new_n411));
  NOR2_X1   g0211(.A1(new_n282), .A2(G68), .ZN(new_n412));
  XNOR2_X1  g0212(.A(new_n412), .B(KEYINPUT12), .ZN(new_n413));
  AND2_X1   g0213(.A1(new_n359), .A2(new_n280), .ZN(new_n414));
  AOI21_X1  g0214(.A(new_n413), .B1(G68), .B2(new_n414), .ZN(new_n415));
  NAND3_X1  g0215(.A1(new_n410), .A2(new_n411), .A3(new_n415), .ZN(new_n416));
  INV_X1    g0216(.A(KEYINPUT14), .ZN(new_n417));
  NAND4_X1  g0217(.A1(new_n376), .A2(KEYINPUT69), .A3(G232), .A4(G1698), .ZN(new_n418));
  INV_X1    g0218(.A(G97), .ZN(new_n419));
  NOR2_X1   g0219(.A1(new_n367), .A2(new_n419), .ZN(new_n420));
  NOR2_X1   g0220(.A1(new_n307), .A2(G1698), .ZN(new_n421));
  AOI21_X1  g0221(.A(new_n420), .B1(new_n376), .B2(new_n421), .ZN(new_n422));
  INV_X1    g0222(.A(KEYINPUT69), .ZN(new_n423));
  NAND2_X1  g0223(.A1(G232), .A2(G1698), .ZN(new_n424));
  OAI21_X1  g0224(.A(new_n423), .B1(new_n252), .B2(new_n424), .ZN(new_n425));
  NAND3_X1  g0225(.A1(new_n418), .A2(new_n422), .A3(new_n425), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n426), .A2(new_n312), .ZN(new_n427));
  NAND3_X1  g0227(.A1(new_n339), .A2(G238), .A3(new_n341), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n382), .A2(new_n428), .ZN(new_n429));
  INV_X1    g0229(.A(new_n429), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n427), .A2(new_n430), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n431), .A2(KEYINPUT13), .ZN(new_n432));
  INV_X1    g0232(.A(KEYINPUT13), .ZN(new_n433));
  NAND3_X1  g0233(.A1(new_n427), .A2(new_n433), .A3(new_n430), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n432), .A2(new_n434), .ZN(new_n435));
  AOI21_X1  g0235(.A(new_n417), .B1(new_n435), .B2(G169), .ZN(new_n436));
  AOI21_X1  g0236(.A(new_n433), .B1(new_n427), .B2(new_n430), .ZN(new_n437));
  AOI211_X1 g0237(.A(KEYINPUT13), .B(new_n429), .C1(new_n426), .C2(new_n312), .ZN(new_n438));
  OAI211_X1 g0238(.A(new_n417), .B(G169), .C1(new_n437), .C2(new_n438), .ZN(new_n439));
  NAND3_X1  g0239(.A1(new_n432), .A2(G179), .A3(new_n434), .ZN(new_n440));
  NAND2_X1  g0240(.A1(new_n439), .A2(new_n440), .ZN(new_n441));
  OAI21_X1  g0241(.A(new_n416), .B1(new_n436), .B2(new_n441), .ZN(new_n442));
  INV_X1    g0242(.A(new_n416), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n435), .A2(G200), .ZN(new_n444));
  OAI211_X1 g0244(.A(new_n443), .B(new_n444), .C1(new_n336), .C2(new_n435), .ZN(new_n445));
  NAND2_X1  g0245(.A1(G238), .A2(G1698), .ZN(new_n446));
  OAI211_X1 g0246(.A(new_n376), .B(new_n446), .C1(new_n227), .C2(G1698), .ZN(new_n447));
  OAI211_X1 g0247(.A(new_n447), .B(new_n312), .C1(G107), .C2(new_n376), .ZN(new_n448));
  NAND2_X1  g0248(.A1(new_n319), .A2(G244), .ZN(new_n449));
  NAND3_X1  g0249(.A1(new_n448), .A2(new_n382), .A3(new_n449), .ZN(new_n450));
  OR2_X1    g0250(.A1(new_n450), .A2(G179), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n450), .A2(new_n398), .ZN(new_n452));
  NAND2_X1  g0252(.A1(G20), .A2(G77), .ZN(new_n453));
  XNOR2_X1  g0253(.A(KEYINPUT15), .B(G87), .ZN(new_n454));
  OAI221_X1 g0254(.A(new_n453), .B1(new_n288), .B2(new_n368), .C1(new_n369), .C2(new_n454), .ZN(new_n455));
  AOI22_X1  g0255(.A1(new_n455), .A2(new_n269), .B1(new_n221), .B2(new_n289), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n414), .A2(G77), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n456), .A2(new_n457), .ZN(new_n458));
  NAND3_X1  g0258(.A1(new_n451), .A2(new_n452), .A3(new_n458), .ZN(new_n459));
  INV_X1    g0259(.A(new_n458), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n450), .A2(G200), .ZN(new_n461));
  OAI211_X1 g0261(.A(new_n460), .B(new_n461), .C1(new_n336), .C2(new_n450), .ZN(new_n462));
  NAND4_X1  g0262(.A1(new_n442), .A2(new_n445), .A3(new_n459), .A4(new_n462), .ZN(new_n463));
  INV_X1    g0263(.A(new_n463), .ZN(new_n464));
  AOI21_X1  g0264(.A(KEYINPUT75), .B1(new_n404), .B2(new_n464), .ZN(new_n465));
  AND3_X1   g0265(.A1(new_n389), .A2(new_n396), .A3(new_n402), .ZN(new_n466));
  NAND3_X1  g0266(.A1(new_n466), .A2(new_n357), .A3(new_n334), .ZN(new_n467));
  INV_X1    g0267(.A(KEYINPUT75), .ZN(new_n468));
  NOR3_X1   g0268(.A1(new_n467), .A2(new_n468), .A3(new_n463), .ZN(new_n469));
  OR2_X1    g0269(.A1(new_n465), .A2(new_n469), .ZN(new_n470));
  INV_X1    g0270(.A(KEYINPUT4), .ZN(new_n471));
  NOR2_X1   g0271(.A1(new_n471), .A2(G1698), .ZN(new_n472));
  OAI211_X1 g0272(.A(new_n472), .B(G244), .C1(new_n251), .C2(new_n250), .ZN(new_n473));
  NAND2_X1  g0273(.A1(G33), .A2(G283), .ZN(new_n474));
  AOI21_X1  g0274(.A(new_n222), .B1(new_n254), .B2(new_n255), .ZN(new_n475));
  OAI211_X1 g0275(.A(new_n473), .B(new_n474), .C1(new_n475), .C2(KEYINPUT4), .ZN(new_n476));
  OAI21_X1  g0276(.A(G250), .B1(new_n250), .B2(new_n251), .ZN(new_n477));
  AOI21_X1  g0277(.A(new_n377), .B1(new_n477), .B2(KEYINPUT4), .ZN(new_n478));
  OAI21_X1  g0278(.A(new_n312), .B1(new_n476), .B2(new_n478), .ZN(new_n479));
  INV_X1    g0279(.A(KEYINPUT5), .ZN(new_n480));
  OAI211_X1 g0280(.A(new_n207), .B(G45), .C1(new_n480), .C2(G41), .ZN(new_n481));
  INV_X1    g0281(.A(new_n481), .ZN(new_n482));
  OAI21_X1  g0282(.A(new_n480), .B1(new_n343), .B2(new_n344), .ZN(new_n483));
  AOI21_X1  g0283(.A(new_n312), .B1(new_n482), .B2(new_n483), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n320), .A2(new_n321), .ZN(new_n485));
  AOI21_X1  g0285(.A(new_n481), .B1(new_n485), .B2(new_n480), .ZN(new_n486));
  NOR2_X1   g0286(.A1(new_n312), .A2(new_n323), .ZN(new_n487));
  AOI22_X1  g0287(.A1(new_n484), .A2(G257), .B1(new_n486), .B2(new_n487), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n479), .A2(new_n488), .ZN(new_n489));
  NOR2_X1   g0289(.A1(new_n489), .A2(G179), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n289), .A2(new_n419), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n207), .A2(G33), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n359), .A2(new_n492), .ZN(new_n493));
  OAI21_X1  g0293(.A(new_n491), .B1(new_n493), .B2(new_n419), .ZN(new_n494));
  INV_X1    g0294(.A(KEYINPUT6), .ZN(new_n495));
  AND2_X1   g0295(.A1(G97), .A2(G107), .ZN(new_n496));
  NOR2_X1   g0296(.A1(G97), .A2(G107), .ZN(new_n497));
  OAI21_X1  g0297(.A(new_n495), .B1(new_n496), .B2(new_n497), .ZN(new_n498));
  INV_X1    g0298(.A(KEYINPUT76), .ZN(new_n499));
  NAND2_X1  g0299(.A1(KEYINPUT6), .A2(G97), .ZN(new_n500));
  OAI21_X1  g0300(.A(new_n499), .B1(new_n500), .B2(G107), .ZN(new_n501));
  INV_X1    g0301(.A(G107), .ZN(new_n502));
  NAND4_X1  g0302(.A1(new_n502), .A2(KEYINPUT76), .A3(KEYINPUT6), .A4(G97), .ZN(new_n503));
  NAND3_X1  g0303(.A1(new_n498), .A2(new_n501), .A3(new_n503), .ZN(new_n504));
  AOI22_X1  g0304(.A1(new_n504), .A2(G20), .B1(G77), .B2(new_n262), .ZN(new_n505));
  OAI21_X1  g0305(.A(G107), .B1(new_n253), .B2(new_n257), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  AOI21_X1  g0307(.A(new_n494), .B1(new_n507), .B2(new_n269), .ZN(new_n508));
  AOI21_X1  g0308(.A(G169), .B1(new_n479), .B2(new_n488), .ZN(new_n509));
  NOR3_X1   g0309(.A1(new_n490), .A2(new_n508), .A3(new_n509), .ZN(new_n510));
  NAND3_X1  g0310(.A1(new_n479), .A2(new_n488), .A3(G190), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n508), .A2(new_n511), .ZN(new_n512));
  INV_X1    g0312(.A(KEYINPUT77), .ZN(new_n513));
  AOI21_X1  g0313(.A(new_n513), .B1(new_n489), .B2(G200), .ZN(new_n514));
  NOR2_X1   g0314(.A1(new_n512), .A2(new_n514), .ZN(new_n515));
  NAND3_X1  g0315(.A1(new_n489), .A2(new_n513), .A3(G200), .ZN(new_n516));
  AOI21_X1  g0316(.A(new_n510), .B1(new_n515), .B2(new_n516), .ZN(new_n517));
  NAND4_X1  g0317(.A1(new_n207), .A2(new_n502), .A3(G13), .A4(G20), .ZN(new_n518));
  INV_X1    g0318(.A(KEYINPUT25), .ZN(new_n519));
  OAI21_X1  g0319(.A(KEYINPUT81), .B1(new_n518), .B2(new_n519), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n518), .A2(new_n519), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  NAND3_X1  g0322(.A1(new_n518), .A2(KEYINPUT81), .A3(new_n519), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  OAI21_X1  g0324(.A(new_n524), .B1(new_n502), .B2(new_n493), .ZN(new_n525));
  INV_X1    g0325(.A(new_n525), .ZN(new_n526));
  INV_X1    g0326(.A(KEYINPUT23), .ZN(new_n527));
  OAI21_X1  g0327(.A(new_n527), .B1(new_n208), .B2(G107), .ZN(new_n528));
  NAND3_X1  g0328(.A1(new_n502), .A2(KEYINPUT23), .A3(G20), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  NAND3_X1  g0330(.A1(new_n208), .A2(G33), .A3(G116), .ZN(new_n531));
  INV_X1    g0331(.A(KEYINPUT80), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n532), .A2(KEYINPUT24), .ZN(new_n533));
  NAND3_X1  g0333(.A1(new_n530), .A2(new_n531), .A3(new_n533), .ZN(new_n534));
  OAI211_X1 g0334(.A(new_n208), .B(G87), .C1(new_n250), .C2(new_n251), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n535), .A2(KEYINPUT22), .ZN(new_n536));
  INV_X1    g0336(.A(KEYINPUT22), .ZN(new_n537));
  NAND4_X1  g0337(.A1(new_n376), .A2(new_n537), .A3(new_n208), .A4(G87), .ZN(new_n538));
  AOI21_X1  g0338(.A(new_n534), .B1(new_n536), .B2(new_n538), .ZN(new_n539));
  NOR2_X1   g0339(.A1(new_n532), .A2(KEYINPUT24), .ZN(new_n540));
  INV_X1    g0340(.A(new_n540), .ZN(new_n541));
  OAI21_X1  g0341(.A(new_n269), .B1(new_n539), .B2(new_n541), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n536), .A2(new_n538), .ZN(new_n543));
  INV_X1    g0343(.A(new_n534), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n543), .A2(new_n544), .ZN(new_n545));
  NOR2_X1   g0345(.A1(new_n545), .A2(new_n540), .ZN(new_n546));
  OAI21_X1  g0346(.A(new_n526), .B1(new_n542), .B2(new_n546), .ZN(new_n547));
  OAI211_X1 g0347(.A(G257), .B(G1698), .C1(new_n250), .C2(new_n251), .ZN(new_n548));
  NAND2_X1  g0348(.A1(G33), .A2(G294), .ZN(new_n549));
  OAI211_X1 g0349(.A(new_n548), .B(new_n549), .C1(new_n477), .C2(G1698), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n550), .A2(new_n312), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n486), .A2(new_n487), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n484), .A2(G264), .ZN(new_n553));
  NAND3_X1  g0353(.A1(new_n551), .A2(new_n552), .A3(new_n553), .ZN(new_n554));
  INV_X1    g0354(.A(KEYINPUT82), .ZN(new_n555));
  AND3_X1   g0355(.A1(new_n554), .A2(new_n555), .A3(new_n338), .ZN(new_n556));
  NOR2_X1   g0356(.A1(new_n547), .A2(new_n556), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n554), .A2(new_n338), .ZN(new_n558));
  OAI211_X1 g0358(.A(new_n558), .B(KEYINPUT82), .C1(G190), .C2(new_n554), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n554), .A2(new_n398), .ZN(new_n560));
  AOI22_X1  g0360(.A1(new_n550), .A2(new_n312), .B1(new_n484), .B2(G264), .ZN(new_n561));
  NAND3_X1  g0361(.A1(new_n561), .A2(new_n328), .A3(new_n552), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n560), .A2(new_n562), .ZN(new_n563));
  INV_X1    g0363(.A(new_n563), .ZN(new_n564));
  AOI22_X1  g0364(.A1(new_n557), .A2(new_n559), .B1(new_n547), .B2(new_n564), .ZN(new_n565));
  NAND2_X1  g0365(.A1(G244), .A2(G1698), .ZN(new_n566));
  OAI21_X1  g0366(.A(new_n566), .B1(new_n228), .B2(G1698), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n376), .A2(new_n567), .ZN(new_n568));
  NAND2_X1  g0368(.A1(G33), .A2(G116), .ZN(new_n569));
  AOI21_X1  g0369(.A(new_n339), .B1(new_n568), .B2(new_n569), .ZN(new_n570));
  OAI21_X1  g0370(.A(new_n224), .B1(new_n315), .B2(G1), .ZN(new_n571));
  NAND3_X1  g0371(.A1(new_n207), .A2(new_n323), .A3(G45), .ZN(new_n572));
  NAND3_X1  g0372(.A1(new_n339), .A2(new_n571), .A3(new_n572), .ZN(new_n573));
  INV_X1    g0373(.A(new_n573), .ZN(new_n574));
  OAI21_X1  g0374(.A(G200), .B1(new_n570), .B2(new_n574), .ZN(new_n575));
  XOR2_X1   g0375(.A(KEYINPUT15), .B(G87), .Z(new_n576));
  NOR2_X1   g0376(.A1(new_n576), .A2(new_n282), .ZN(new_n577));
  NAND3_X1  g0377(.A1(new_n223), .A2(new_n419), .A3(new_n502), .ZN(new_n578));
  OAI211_X1 g0378(.A(KEYINPUT19), .B(new_n578), .C1(new_n420), .C2(G20), .ZN(new_n579));
  OAI211_X1 g0379(.A(new_n208), .B(G68), .C1(new_n250), .C2(new_n251), .ZN(new_n580));
  INV_X1    g0380(.A(KEYINPUT19), .ZN(new_n581));
  OAI21_X1  g0381(.A(new_n581), .B1(new_n369), .B2(new_n419), .ZN(new_n582));
  NAND3_X1  g0382(.A1(new_n579), .A2(new_n580), .A3(new_n582), .ZN(new_n583));
  AOI21_X1  g0383(.A(new_n577), .B1(new_n583), .B2(new_n269), .ZN(new_n584));
  NAND3_X1  g0384(.A1(new_n359), .A2(G87), .A3(new_n492), .ZN(new_n585));
  NAND3_X1  g0385(.A1(new_n575), .A2(new_n584), .A3(new_n585), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n586), .A2(KEYINPUT79), .ZN(new_n587));
  INV_X1    g0387(.A(KEYINPUT79), .ZN(new_n588));
  NAND4_X1  g0388(.A1(new_n575), .A2(new_n584), .A3(new_n588), .A4(new_n585), .ZN(new_n589));
  AOI22_X1  g0389(.A1(new_n376), .A2(new_n567), .B1(G33), .B2(G116), .ZN(new_n590));
  OAI211_X1 g0390(.A(G190), .B(new_n573), .C1(new_n590), .C2(new_n339), .ZN(new_n591));
  NAND3_X1  g0391(.A1(new_n587), .A2(new_n589), .A3(new_n591), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n583), .A2(new_n269), .ZN(new_n593));
  INV_X1    g0393(.A(new_n577), .ZN(new_n594));
  INV_X1    g0394(.A(KEYINPUT78), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n576), .A2(new_n595), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n454), .A2(KEYINPUT78), .ZN(new_n597));
  NAND4_X1  g0397(.A1(new_n596), .A2(new_n359), .A3(new_n492), .A4(new_n597), .ZN(new_n598));
  NAND3_X1  g0398(.A1(new_n593), .A2(new_n594), .A3(new_n598), .ZN(new_n599));
  OAI211_X1 g0399(.A(new_n328), .B(new_n573), .C1(new_n590), .C2(new_n339), .ZN(new_n600));
  OAI21_X1  g0400(.A(new_n573), .B1(new_n590), .B2(new_n339), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n601), .A2(new_n398), .ZN(new_n602));
  NAND3_X1  g0402(.A1(new_n599), .A2(new_n600), .A3(new_n602), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n592), .A2(new_n603), .ZN(new_n604));
  NAND3_X1  g0404(.A1(new_n359), .A2(G116), .A3(new_n492), .ZN(new_n605));
  INV_X1    g0405(.A(G116), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n289), .A2(new_n606), .ZN(new_n607));
  AOI22_X1  g0407(.A1(new_n268), .A2(new_n215), .B1(G20), .B2(new_n606), .ZN(new_n608));
  OAI211_X1 g0408(.A(new_n474), .B(new_n208), .C1(G33), .C2(new_n419), .ZN(new_n609));
  AND3_X1   g0409(.A1(new_n608), .A2(KEYINPUT20), .A3(new_n609), .ZN(new_n610));
  AOI21_X1  g0410(.A(KEYINPUT20), .B1(new_n608), .B2(new_n609), .ZN(new_n611));
  OAI211_X1 g0411(.A(new_n605), .B(new_n607), .C1(new_n610), .C2(new_n611), .ZN(new_n612));
  AOI21_X1  g0412(.A(KEYINPUT5), .B1(new_n320), .B2(new_n321), .ZN(new_n613));
  OAI211_X1 g0413(.A(G270), .B(new_n339), .C1(new_n613), .C2(new_n481), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n377), .A2(G257), .ZN(new_n615));
  NAND2_X1  g0415(.A1(G264), .A2(G1698), .ZN(new_n616));
  OAI211_X1 g0416(.A(new_n615), .B(new_n616), .C1(new_n250), .C2(new_n251), .ZN(new_n617));
  OAI211_X1 g0417(.A(new_n617), .B(new_n312), .C1(G303), .C2(new_n376), .ZN(new_n618));
  NAND3_X1  g0418(.A1(new_n552), .A2(new_n614), .A3(new_n618), .ZN(new_n619));
  NAND3_X1  g0419(.A1(new_n612), .A2(G169), .A3(new_n619), .ZN(new_n620));
  INV_X1    g0420(.A(KEYINPUT21), .ZN(new_n621));
  NAND4_X1  g0421(.A1(new_n552), .A2(new_n614), .A3(new_n618), .A4(G179), .ZN(new_n622));
  INV_X1    g0422(.A(new_n622), .ZN(new_n623));
  AOI22_X1  g0423(.A1(new_n620), .A2(new_n621), .B1(new_n623), .B2(new_n612), .ZN(new_n624));
  NAND4_X1  g0424(.A1(new_n612), .A2(new_n619), .A3(KEYINPUT21), .A4(G169), .ZN(new_n625));
  INV_X1    g0425(.A(new_n612), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n619), .A2(G200), .ZN(new_n627));
  OAI211_X1 g0427(.A(new_n626), .B(new_n627), .C1(new_n336), .C2(new_n619), .ZN(new_n628));
  NAND3_X1  g0428(.A1(new_n624), .A2(new_n625), .A3(new_n628), .ZN(new_n629));
  NOR2_X1   g0429(.A1(new_n604), .A2(new_n629), .ZN(new_n630));
  AND4_X1   g0430(.A1(new_n470), .A2(new_n517), .A3(new_n565), .A4(new_n630), .ZN(G372));
  INV_X1    g0431(.A(new_n517), .ZN(new_n632));
  NAND4_X1  g0432(.A1(new_n575), .A2(new_n584), .A3(new_n585), .A4(new_n591), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n603), .A2(new_n633), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n634), .A2(KEYINPUT83), .ZN(new_n635));
  INV_X1    g0435(.A(KEYINPUT83), .ZN(new_n636));
  NAND3_X1  g0436(.A1(new_n603), .A2(new_n636), .A3(new_n633), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n635), .A2(new_n637), .ZN(new_n638));
  AOI21_X1  g0438(.A(new_n281), .B1(new_n545), .B2(new_n540), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n539), .A2(new_n541), .ZN(new_n640));
  AOI21_X1  g0440(.A(new_n525), .B1(new_n639), .B2(new_n640), .ZN(new_n641));
  OAI211_X1 g0441(.A(new_n624), .B(new_n625), .C1(new_n641), .C2(new_n563), .ZN(new_n642));
  INV_X1    g0442(.A(new_n556), .ZN(new_n643));
  NAND3_X1  g0443(.A1(new_n559), .A2(new_n643), .A3(new_n641), .ZN(new_n644));
  NAND3_X1  g0444(.A1(new_n638), .A2(new_n642), .A3(new_n644), .ZN(new_n645));
  OAI21_X1  g0445(.A(new_n603), .B1(new_n632), .B2(new_n645), .ZN(new_n646));
  NAND3_X1  g0446(.A1(new_n510), .A2(new_n603), .A3(new_n592), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n647), .A2(KEYINPUT26), .ZN(new_n648));
  INV_X1    g0448(.A(KEYINPUT26), .ZN(new_n649));
  NAND3_X1  g0449(.A1(new_n638), .A2(new_n649), .A3(new_n510), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n648), .A2(new_n650), .ZN(new_n651));
  OAI21_X1  g0451(.A(new_n470), .B1(new_n646), .B2(new_n651), .ZN(new_n652));
  XNOR2_X1  g0452(.A(new_n652), .B(KEYINPUT84), .ZN(new_n653));
  AND4_X1   g0453(.A1(new_n445), .A2(new_n458), .A3(new_n452), .A4(new_n451), .ZN(new_n654));
  INV_X1    g0454(.A(new_n442), .ZN(new_n655));
  OAI21_X1  g0455(.A(new_n357), .B1(new_n654), .B2(new_n655), .ZN(new_n656));
  OAI21_X1  g0456(.A(new_n329), .B1(new_n276), .B2(new_n295), .ZN(new_n657));
  XNOR2_X1  g0457(.A(new_n657), .B(new_n331), .ZN(new_n658));
  AOI21_X1  g0458(.A(new_n397), .B1(new_n656), .B2(new_n658), .ZN(new_n659));
  NOR2_X1   g0459(.A1(new_n659), .A2(new_n403), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n653), .A2(new_n660), .ZN(G369));
  NAND3_X1  g0461(.A1(new_n207), .A2(new_n208), .A3(G13), .ZN(new_n662));
  OR2_X1    g0462(.A1(new_n662), .A2(KEYINPUT27), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n662), .A2(KEYINPUT27), .ZN(new_n664));
  NAND3_X1  g0464(.A1(new_n663), .A2(G213), .A3(new_n664), .ZN(new_n665));
  XOR2_X1   g0465(.A(KEYINPUT85), .B(G343), .Z(new_n666));
  NOR2_X1   g0466(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  INV_X1    g0467(.A(new_n667), .ZN(new_n668));
  OAI21_X1  g0468(.A(new_n565), .B1(new_n641), .B2(new_n668), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n564), .A2(new_n547), .ZN(new_n670));
  OAI21_X1  g0470(.A(new_n669), .B1(new_n670), .B2(new_n668), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n624), .A2(new_n625), .ZN(new_n672));
  NOR2_X1   g0472(.A1(new_n626), .A2(new_n668), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  OAI21_X1  g0474(.A(new_n674), .B1(new_n629), .B2(new_n673), .ZN(new_n675));
  AND2_X1   g0475(.A1(new_n675), .A2(G330), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n671), .A2(new_n676), .ZN(new_n677));
  AND4_X1   g0477(.A1(new_n670), .A2(new_n644), .A3(new_n672), .A4(new_n668), .ZN(new_n678));
  NOR2_X1   g0478(.A1(new_n670), .A2(new_n667), .ZN(new_n679));
  NOR2_X1   g0479(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n677), .A2(new_n680), .ZN(G399));
  INV_X1    g0481(.A(new_n211), .ZN(new_n682));
  NOR2_X1   g0482(.A1(new_n682), .A2(new_n485), .ZN(new_n683));
  INV_X1    g0483(.A(new_n683), .ZN(new_n684));
  NOR2_X1   g0484(.A1(new_n578), .A2(G116), .ZN(new_n685));
  NAND3_X1  g0485(.A1(new_n684), .A2(G1), .A3(new_n685), .ZN(new_n686));
  INV_X1    g0486(.A(KEYINPUT86), .ZN(new_n687));
  AOI22_X1  g0487(.A1(new_n686), .A2(new_n687), .B1(new_n218), .B2(new_n683), .ZN(new_n688));
  OAI21_X1  g0488(.A(new_n688), .B1(new_n687), .B2(new_n686), .ZN(new_n689));
  XNOR2_X1  g0489(.A(new_n689), .B(KEYINPUT28), .ZN(new_n690));
  INV_X1    g0490(.A(KEYINPUT30), .ZN(new_n691));
  INV_X1    g0491(.A(KEYINPUT87), .ZN(new_n692));
  XNOR2_X1  g0492(.A(new_n622), .B(new_n692), .ZN(new_n693));
  INV_X1    g0493(.A(new_n601), .ZN(new_n694));
  NAND4_X1  g0494(.A1(new_n479), .A2(new_n561), .A3(new_n694), .A4(new_n488), .ZN(new_n695));
  OAI21_X1  g0495(.A(new_n691), .B1(new_n693), .B2(new_n695), .ZN(new_n696));
  XNOR2_X1  g0496(.A(new_n622), .B(KEYINPUT87), .ZN(new_n697));
  INV_X1    g0497(.A(new_n695), .ZN(new_n698));
  NAND3_X1  g0498(.A1(new_n697), .A2(new_n698), .A3(KEYINPUT30), .ZN(new_n699));
  NOR2_X1   g0499(.A1(new_n694), .A2(G179), .ZN(new_n700));
  NAND4_X1  g0500(.A1(new_n700), .A2(new_n489), .A3(new_n554), .A4(new_n619), .ZN(new_n701));
  NAND3_X1  g0501(.A1(new_n696), .A2(new_n699), .A3(new_n701), .ZN(new_n702));
  NAND2_X1  g0502(.A1(new_n702), .A2(new_n667), .ZN(new_n703));
  INV_X1    g0503(.A(KEYINPUT31), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n703), .A2(new_n704), .ZN(new_n705));
  NAND4_X1  g0505(.A1(new_n630), .A2(new_n517), .A3(new_n565), .A4(new_n668), .ZN(new_n706));
  NAND3_X1  g0506(.A1(new_n702), .A2(KEYINPUT31), .A3(new_n667), .ZN(new_n707));
  NAND3_X1  g0507(.A1(new_n705), .A2(new_n706), .A3(new_n707), .ZN(new_n708));
  AND3_X1   g0508(.A1(new_n708), .A2(KEYINPUT88), .A3(G330), .ZN(new_n709));
  AOI21_X1  g0509(.A(KEYINPUT88), .B1(new_n708), .B2(G330), .ZN(new_n710));
  NOR2_X1   g0510(.A1(new_n709), .A2(new_n710), .ZN(new_n711));
  INV_X1    g0511(.A(new_n603), .ZN(new_n712));
  AND3_X1   g0512(.A1(new_n638), .A2(new_n644), .A3(new_n642), .ZN(new_n713));
  AOI21_X1  g0513(.A(new_n712), .B1(new_n713), .B2(new_n517), .ZN(new_n714));
  INV_X1    g0514(.A(new_n637), .ZN(new_n715));
  AOI21_X1  g0515(.A(new_n636), .B1(new_n603), .B2(new_n633), .ZN(new_n716));
  OAI211_X1 g0516(.A(new_n510), .B(KEYINPUT26), .C1(new_n715), .C2(new_n716), .ZN(new_n717));
  INV_X1    g0517(.A(KEYINPUT89), .ZN(new_n718));
  NAND2_X1  g0518(.A1(new_n717), .A2(new_n718), .ZN(new_n719));
  NAND4_X1  g0519(.A1(new_n638), .A2(KEYINPUT89), .A3(KEYINPUT26), .A4(new_n510), .ZN(new_n720));
  NAND2_X1  g0520(.A1(new_n647), .A2(new_n649), .ZN(new_n721));
  NAND3_X1  g0521(.A1(new_n719), .A2(new_n720), .A3(new_n721), .ZN(new_n722));
  AOI21_X1  g0522(.A(new_n667), .B1(new_n714), .B2(new_n722), .ZN(new_n723));
  NAND2_X1  g0523(.A1(new_n723), .A2(KEYINPUT29), .ZN(new_n724));
  OAI21_X1  g0524(.A(new_n668), .B1(new_n646), .B2(new_n651), .ZN(new_n725));
  INV_X1    g0525(.A(KEYINPUT29), .ZN(new_n726));
  NAND2_X1  g0526(.A1(new_n725), .A2(new_n726), .ZN(new_n727));
  NAND2_X1  g0527(.A1(new_n724), .A2(new_n727), .ZN(new_n728));
  NAND2_X1  g0528(.A1(new_n711), .A2(new_n728), .ZN(new_n729));
  INV_X1    g0529(.A(new_n729), .ZN(new_n730));
  OAI21_X1  g0530(.A(new_n690), .B1(new_n730), .B2(G1), .ZN(G364));
  AND2_X1   g0531(.A1(new_n208), .A2(G13), .ZN(new_n732));
  AOI21_X1  g0532(.A(new_n207), .B1(new_n732), .B2(G45), .ZN(new_n733));
  INV_X1    g0533(.A(new_n733), .ZN(new_n734));
  NOR2_X1   g0534(.A1(new_n683), .A2(new_n734), .ZN(new_n735));
  INV_X1    g0535(.A(new_n735), .ZN(new_n736));
  AOI21_X1  g0536(.A(new_n215), .B1(G20), .B2(new_n398), .ZN(new_n737));
  INV_X1    g0537(.A(new_n737), .ZN(new_n738));
  NOR2_X1   g0538(.A1(new_n208), .A2(G190), .ZN(new_n739));
  NAND3_X1  g0539(.A1(new_n739), .A2(new_n328), .A3(new_n338), .ZN(new_n740));
  INV_X1    g0540(.A(KEYINPUT94), .ZN(new_n741));
  OR2_X1    g0541(.A1(new_n740), .A2(new_n741), .ZN(new_n742));
  NAND2_X1  g0542(.A1(new_n740), .A2(new_n741), .ZN(new_n743));
  NAND2_X1  g0543(.A1(new_n742), .A2(new_n743), .ZN(new_n744));
  INV_X1    g0544(.A(G159), .ZN(new_n745));
  NOR2_X1   g0545(.A1(new_n744), .A2(new_n745), .ZN(new_n746));
  XNOR2_X1  g0546(.A(new_n746), .B(KEYINPUT32), .ZN(new_n747));
  NOR2_X1   g0547(.A1(new_n208), .A2(new_n336), .ZN(new_n748));
  NOR2_X1   g0548(.A1(new_n338), .A2(G179), .ZN(new_n749));
  NAND2_X1  g0549(.A1(new_n748), .A2(new_n749), .ZN(new_n750));
  INV_X1    g0550(.A(new_n750), .ZN(new_n751));
  NOR2_X1   g0551(.A1(new_n328), .A2(G200), .ZN(new_n752));
  NAND2_X1  g0552(.A1(new_n739), .A2(new_n752), .ZN(new_n753));
  INV_X1    g0553(.A(new_n753), .ZN(new_n754));
  AOI22_X1  g0554(.A1(G87), .A2(new_n751), .B1(new_n754), .B2(G77), .ZN(new_n755));
  NAND2_X1  g0555(.A1(new_n748), .A2(new_n752), .ZN(new_n756));
  OAI21_X1  g0556(.A(new_n755), .B1(new_n202), .B2(new_n756), .ZN(new_n757));
  NOR3_X1   g0557(.A1(new_n336), .A2(G179), .A3(G200), .ZN(new_n758));
  NOR2_X1   g0558(.A1(new_n758), .A2(new_n208), .ZN(new_n759));
  NOR2_X1   g0559(.A1(new_n759), .A2(new_n419), .ZN(new_n760));
  NAND2_X1  g0560(.A1(new_n739), .A2(new_n749), .ZN(new_n761));
  NAND3_X1  g0561(.A1(G20), .A2(G179), .A3(G200), .ZN(new_n762));
  NOR2_X1   g0562(.A1(new_n762), .A2(G190), .ZN(new_n763));
  INV_X1    g0563(.A(new_n763), .ZN(new_n764));
  OAI221_X1 g0564(.A(new_n376), .B1(new_n761), .B2(new_n502), .C1(new_n764), .C2(new_n203), .ZN(new_n765));
  NOR3_X1   g0565(.A1(new_n757), .A2(new_n760), .A3(new_n765), .ZN(new_n766));
  NOR2_X1   g0566(.A1(new_n762), .A2(new_n336), .ZN(new_n767));
  INV_X1    g0567(.A(KEYINPUT93), .ZN(new_n768));
  NOR2_X1   g0568(.A1(new_n767), .A2(new_n768), .ZN(new_n769));
  NOR3_X1   g0569(.A1(new_n762), .A2(KEYINPUT93), .A3(new_n336), .ZN(new_n770));
  NOR2_X1   g0570(.A1(new_n769), .A2(new_n770), .ZN(new_n771));
  OAI211_X1 g0571(.A(new_n747), .B(new_n766), .C1(new_n201), .C2(new_n771), .ZN(new_n772));
  INV_X1    g0572(.A(G303), .ZN(new_n773));
  OAI21_X1  g0573(.A(new_n252), .B1(new_n750), .B2(new_n773), .ZN(new_n774));
  OR2_X1    g0574(.A1(KEYINPUT33), .A2(G317), .ZN(new_n775));
  NAND2_X1  g0575(.A1(KEYINPUT33), .A2(G317), .ZN(new_n776));
  AOI21_X1  g0576(.A(new_n764), .B1(new_n775), .B2(new_n776), .ZN(new_n777));
  INV_X1    g0577(.A(new_n759), .ZN(new_n778));
  AOI211_X1 g0578(.A(new_n774), .B(new_n777), .C1(G294), .C2(new_n778), .ZN(new_n779));
  INV_X1    g0579(.A(new_n771), .ZN(new_n780));
  NAND2_X1  g0580(.A1(new_n780), .A2(G326), .ZN(new_n781));
  INV_X1    g0581(.A(new_n744), .ZN(new_n782));
  NAND2_X1  g0582(.A1(new_n782), .A2(G329), .ZN(new_n783));
  INV_X1    g0583(.A(G283), .ZN(new_n784));
  INV_X1    g0584(.A(G311), .ZN(new_n785));
  OAI22_X1  g0585(.A1(new_n784), .A2(new_n761), .B1(new_n753), .B2(new_n785), .ZN(new_n786));
  INV_X1    g0586(.A(new_n756), .ZN(new_n787));
  AOI21_X1  g0587(.A(new_n786), .B1(G322), .B2(new_n787), .ZN(new_n788));
  NAND4_X1  g0588(.A1(new_n779), .A2(new_n781), .A3(new_n783), .A4(new_n788), .ZN(new_n789));
  AOI21_X1  g0589(.A(new_n738), .B1(new_n772), .B2(new_n789), .ZN(new_n790));
  NOR2_X1   g0590(.A1(G13), .A2(G33), .ZN(new_n791));
  XNOR2_X1  g0591(.A(new_n791), .B(KEYINPUT92), .ZN(new_n792));
  NOR2_X1   g0592(.A1(new_n792), .A2(G20), .ZN(new_n793));
  NOR2_X1   g0593(.A1(new_n793), .A2(new_n737), .ZN(new_n794));
  NAND2_X1  g0594(.A1(new_n211), .A2(new_n376), .ZN(new_n795));
  INV_X1    g0595(.A(KEYINPUT90), .ZN(new_n796));
  AOI21_X1  g0596(.A(new_n795), .B1(new_n796), .B2(G355), .ZN(new_n797));
  OAI21_X1  g0597(.A(new_n797), .B1(new_n796), .B2(G355), .ZN(new_n798));
  OAI21_X1  g0598(.A(new_n798), .B1(G116), .B2(new_n211), .ZN(new_n799));
  OR2_X1    g0599(.A1(new_n799), .A2(KEYINPUT91), .ZN(new_n800));
  NOR2_X1   g0600(.A1(new_n682), .A2(new_n376), .ZN(new_n801));
  INV_X1    g0601(.A(new_n801), .ZN(new_n802));
  AOI21_X1  g0602(.A(new_n802), .B1(new_n315), .B2(new_n218), .ZN(new_n803));
  OAI21_X1  g0603(.A(new_n803), .B1(new_n244), .B2(new_n315), .ZN(new_n804));
  NAND2_X1  g0604(.A1(new_n799), .A2(KEYINPUT91), .ZN(new_n805));
  NAND3_X1  g0605(.A1(new_n800), .A2(new_n804), .A3(new_n805), .ZN(new_n806));
  AOI211_X1 g0606(.A(new_n736), .B(new_n790), .C1(new_n794), .C2(new_n806), .ZN(new_n807));
  INV_X1    g0607(.A(new_n793), .ZN(new_n808));
  OAI21_X1  g0608(.A(new_n807), .B1(new_n675), .B2(new_n808), .ZN(new_n809));
  XNOR2_X1  g0609(.A(new_n809), .B(KEYINPUT95), .ZN(new_n810));
  NOR2_X1   g0610(.A1(new_n676), .A2(new_n735), .ZN(new_n811));
  OAI21_X1  g0611(.A(new_n811), .B1(G330), .B2(new_n675), .ZN(new_n812));
  NAND2_X1  g0612(.A1(new_n810), .A2(new_n812), .ZN(G396));
  OAI21_X1  g0613(.A(new_n462), .B1(new_n460), .B2(new_n668), .ZN(new_n814));
  NAND2_X1  g0614(.A1(new_n814), .A2(new_n459), .ZN(new_n815));
  OR2_X1    g0615(.A1(new_n459), .A2(new_n667), .ZN(new_n816));
  NAND2_X1  g0616(.A1(new_n815), .A2(new_n816), .ZN(new_n817));
  NAND2_X1  g0617(.A1(new_n725), .A2(new_n817), .ZN(new_n818));
  INV_X1    g0618(.A(new_n817), .ZN(new_n819));
  OAI211_X1 g0619(.A(new_n819), .B(new_n668), .C1(new_n646), .C2(new_n651), .ZN(new_n820));
  NAND2_X1  g0620(.A1(new_n818), .A2(new_n820), .ZN(new_n821));
  AOI21_X1  g0621(.A(new_n735), .B1(new_n711), .B2(new_n821), .ZN(new_n822));
  OAI21_X1  g0622(.A(new_n822), .B1(new_n711), .B2(new_n821), .ZN(new_n823));
  INV_X1    g0623(.A(new_n761), .ZN(new_n824));
  AOI21_X1  g0624(.A(new_n252), .B1(new_n824), .B2(G68), .ZN(new_n825));
  OAI221_X1 g0625(.A(new_n825), .B1(new_n201), .B2(new_n750), .C1(new_n202), .C2(new_n759), .ZN(new_n826));
  AOI22_X1  g0626(.A1(G143), .A2(new_n787), .B1(new_n754), .B2(G159), .ZN(new_n827));
  INV_X1    g0627(.A(G137), .ZN(new_n828));
  OAI221_X1 g0628(.A(new_n827), .B1(new_n366), .B2(new_n764), .C1(new_n771), .C2(new_n828), .ZN(new_n829));
  XOR2_X1   g0629(.A(new_n829), .B(KEYINPUT34), .Z(new_n830));
  AOI211_X1 g0630(.A(new_n826), .B(new_n830), .C1(G132), .C2(new_n782), .ZN(new_n831));
  INV_X1    g0631(.A(G294), .ZN(new_n832));
  OAI21_X1  g0632(.A(new_n252), .B1(new_n756), .B2(new_n832), .ZN(new_n833));
  AOI211_X1 g0633(.A(new_n833), .B(new_n760), .C1(G283), .C2(new_n763), .ZN(new_n834));
  OAI22_X1  g0634(.A1(new_n223), .A2(new_n761), .B1(new_n753), .B2(new_n606), .ZN(new_n835));
  AOI21_X1  g0635(.A(new_n835), .B1(G107), .B2(new_n751), .ZN(new_n836));
  OAI211_X1 g0636(.A(new_n834), .B(new_n836), .C1(new_n785), .C2(new_n744), .ZN(new_n837));
  AOI21_X1  g0637(.A(new_n837), .B1(G303), .B2(new_n780), .ZN(new_n838));
  OAI21_X1  g0638(.A(new_n737), .B1(new_n831), .B2(new_n838), .ZN(new_n839));
  NOR2_X1   g0639(.A1(new_n737), .A2(new_n791), .ZN(new_n840));
  AOI21_X1  g0640(.A(new_n736), .B1(new_n221), .B2(new_n840), .ZN(new_n841));
  OAI211_X1 g0641(.A(new_n839), .B(new_n841), .C1(new_n792), .C2(new_n819), .ZN(new_n842));
  NAND2_X1  g0642(.A1(new_n823), .A2(new_n842), .ZN(G384));
  NAND2_X1  g0643(.A1(new_n416), .A2(new_n667), .ZN(new_n844));
  NAND3_X1  g0644(.A1(new_n442), .A2(new_n445), .A3(new_n844), .ZN(new_n845));
  OAI211_X1 g0645(.A(new_n416), .B(new_n667), .C1(new_n436), .C2(new_n441), .ZN(new_n846));
  AOI21_X1  g0646(.A(new_n817), .B1(new_n845), .B2(new_n846), .ZN(new_n847));
  NOR2_X1   g0647(.A1(KEYINPUT97), .A2(KEYINPUT31), .ZN(new_n848));
  NAND2_X1  g0648(.A1(new_n703), .A2(new_n848), .ZN(new_n849));
  OAI211_X1 g0649(.A(new_n702), .B(new_n667), .C1(KEYINPUT97), .C2(KEYINPUT31), .ZN(new_n850));
  NAND3_X1  g0650(.A1(new_n849), .A2(new_n706), .A3(new_n850), .ZN(new_n851));
  NAND2_X1  g0651(.A1(new_n847), .A2(new_n851), .ZN(new_n852));
  INV_X1    g0652(.A(KEYINPUT40), .ZN(new_n853));
  NOR2_X1   g0653(.A1(new_n852), .A2(new_n853), .ZN(new_n854));
  NAND3_X1  g0654(.A1(new_n301), .A2(new_n287), .A3(new_n290), .ZN(new_n855));
  INV_X1    g0655(.A(new_n665), .ZN(new_n856));
  NAND2_X1  g0656(.A1(new_n855), .A2(new_n856), .ZN(new_n857));
  INV_X1    g0657(.A(new_n857), .ZN(new_n858));
  NAND2_X1  g0658(.A1(new_n358), .A2(new_n858), .ZN(new_n859));
  AOI21_X1  g0659(.A(new_n295), .B1(new_n300), .B2(new_n298), .ZN(new_n860));
  AOI21_X1  g0660(.A(new_n352), .B1(new_n860), .B2(new_n349), .ZN(new_n861));
  INV_X1    g0661(.A(new_n353), .ZN(new_n862));
  NOR3_X1   g0662(.A1(new_n861), .A2(new_n862), .A3(KEYINPUT37), .ZN(new_n863));
  OAI211_X1 g0663(.A(new_n296), .B(new_n305), .C1(new_n329), .C2(new_n856), .ZN(new_n864));
  OAI21_X1  g0664(.A(new_n855), .B1(new_n329), .B2(new_n856), .ZN(new_n865));
  NAND3_X1  g0665(.A1(new_n865), .A2(new_n351), .A3(new_n353), .ZN(new_n866));
  AOI22_X1  g0666(.A1(new_n863), .A2(new_n864), .B1(new_n866), .B2(KEYINPUT37), .ZN(new_n867));
  INV_X1    g0667(.A(new_n867), .ZN(new_n868));
  NAND3_X1  g0668(.A1(new_n859), .A2(KEYINPUT38), .A3(new_n868), .ZN(new_n869));
  NAND3_X1  g0669(.A1(new_n296), .A2(new_n305), .A3(new_n856), .ZN(new_n870));
  NAND3_X1  g0670(.A1(new_n870), .A2(new_n350), .A3(new_n657), .ZN(new_n871));
  AOI22_X1  g0671(.A1(new_n864), .A2(new_n863), .B1(new_n871), .B2(KEYINPUT37), .ZN(new_n872));
  OAI21_X1  g0672(.A(KEYINPUT17), .B1(new_n861), .B2(new_n862), .ZN(new_n873));
  INV_X1    g0673(.A(KEYINPUT96), .ZN(new_n874));
  NAND3_X1  g0674(.A1(new_n873), .A2(new_n874), .A3(new_n355), .ZN(new_n875));
  OAI21_X1  g0675(.A(KEYINPUT96), .B1(new_n354), .B2(new_n356), .ZN(new_n876));
  NAND3_X1  g0676(.A1(new_n875), .A2(new_n658), .A3(new_n876), .ZN(new_n877));
  INV_X1    g0677(.A(new_n870), .ZN(new_n878));
  AOI21_X1  g0678(.A(new_n872), .B1(new_n877), .B2(new_n878), .ZN(new_n879));
  OAI21_X1  g0679(.A(new_n869), .B1(new_n879), .B2(KEYINPUT38), .ZN(new_n880));
  AND2_X1   g0680(.A1(new_n854), .A2(new_n880), .ZN(new_n881));
  INV_X1    g0681(.A(KEYINPUT98), .ZN(new_n882));
  INV_X1    g0682(.A(KEYINPUT38), .ZN(new_n883));
  AOI21_X1  g0683(.A(new_n857), .B1(new_n334), .B2(new_n357), .ZN(new_n884));
  OAI21_X1  g0684(.A(new_n883), .B1(new_n884), .B2(new_n867), .ZN(new_n885));
  AOI21_X1  g0685(.A(new_n852), .B1(new_n869), .B2(new_n885), .ZN(new_n886));
  OAI21_X1  g0686(.A(new_n882), .B1(new_n886), .B2(KEYINPUT40), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n869), .A2(new_n885), .ZN(new_n888));
  AND2_X1   g0688(.A1(new_n847), .A2(new_n851), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  NAND3_X1  g0690(.A1(new_n890), .A2(KEYINPUT98), .A3(new_n853), .ZN(new_n891));
  AOI21_X1  g0691(.A(new_n881), .B1(new_n887), .B2(new_n891), .ZN(new_n892));
  INV_X1    g0692(.A(new_n892), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n470), .A2(new_n851), .ZN(new_n894));
  OAI21_X1  g0694(.A(G330), .B1(new_n893), .B2(new_n894), .ZN(new_n895));
  AOI21_X1  g0695(.A(new_n895), .B1(new_n894), .B2(new_n893), .ZN(new_n896));
  NOR2_X1   g0696(.A1(new_n658), .A2(new_n856), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n820), .A2(new_n816), .ZN(new_n898));
  INV_X1    g0698(.A(new_n898), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n845), .A2(new_n846), .ZN(new_n900));
  INV_X1    g0700(.A(new_n900), .ZN(new_n901));
  NOR2_X1   g0701(.A1(new_n899), .A2(new_n901), .ZN(new_n902));
  AOI21_X1  g0702(.A(new_n897), .B1(new_n902), .B2(new_n888), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n888), .A2(KEYINPUT39), .ZN(new_n904));
  INV_X1    g0704(.A(KEYINPUT39), .ZN(new_n905));
  OAI211_X1 g0705(.A(new_n869), .B(new_n905), .C1(new_n879), .C2(KEYINPUT38), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n904), .A2(new_n906), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n655), .A2(new_n668), .ZN(new_n908));
  INV_X1    g0708(.A(new_n908), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n907), .A2(new_n909), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n903), .A2(new_n910), .ZN(new_n911));
  OAI211_X1 g0711(.A(new_n724), .B(new_n727), .C1(new_n465), .C2(new_n469), .ZN(new_n912));
  AND2_X1   g0712(.A1(new_n912), .A2(new_n660), .ZN(new_n913));
  XNOR2_X1  g0713(.A(new_n911), .B(new_n913), .ZN(new_n914));
  OAI22_X1  g0714(.A1(new_n896), .A2(new_n914), .B1(new_n207), .B2(new_n732), .ZN(new_n915));
  AOI21_X1  g0715(.A(new_n915), .B1(new_n914), .B2(new_n896), .ZN(new_n916));
  OR2_X1    g0716(.A1(new_n504), .A2(KEYINPUT35), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n504), .A2(KEYINPUT35), .ZN(new_n918));
  NAND4_X1  g0718(.A1(new_n917), .A2(G116), .A3(new_n216), .A4(new_n918), .ZN(new_n919));
  XOR2_X1   g0719(.A(new_n919), .B(KEYINPUT36), .Z(new_n920));
  OAI211_X1 g0720(.A(new_n218), .B(G77), .C1(new_n202), .C2(new_n203), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n201), .A2(G68), .ZN(new_n922));
  AOI211_X1 g0722(.A(new_n207), .B(G13), .C1(new_n921), .C2(new_n922), .ZN(new_n923));
  NOR3_X1   g0723(.A1(new_n916), .A2(new_n920), .A3(new_n923), .ZN(new_n924));
  XOR2_X1   g0724(.A(new_n924), .B(KEYINPUT99), .Z(G367));
  AOI21_X1  g0725(.A(new_n668), .B1(new_n584), .B2(new_n585), .ZN(new_n926));
  XNOR2_X1  g0726(.A(new_n926), .B(KEYINPUT100), .ZN(new_n927));
  AND2_X1   g0727(.A1(new_n927), .A2(new_n712), .ZN(new_n928));
  OR2_X1    g0728(.A1(new_n928), .A2(KEYINPUT101), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n928), .A2(KEYINPUT101), .ZN(new_n930));
  INV_X1    g0730(.A(new_n638), .ZN(new_n931));
  OAI211_X1 g0731(.A(new_n929), .B(new_n930), .C1(new_n931), .C2(new_n927), .ZN(new_n932));
  OR2_X1    g0732(.A1(new_n932), .A2(new_n808), .ZN(new_n933));
  OAI21_X1  g0733(.A(new_n794), .B1(new_n211), .B2(new_n454), .ZN(new_n934));
  AND2_X1   g0734(.A1(new_n801), .A2(new_n240), .ZN(new_n935));
  OAI21_X1  g0735(.A(new_n735), .B1(new_n934), .B2(new_n935), .ZN(new_n936));
  XNOR2_X1  g0736(.A(new_n936), .B(KEYINPUT104), .ZN(new_n937));
  OAI221_X1 g0737(.A(new_n376), .B1(new_n756), .B2(new_n366), .C1(new_n745), .C2(new_n764), .ZN(new_n938));
  AOI21_X1  g0738(.A(new_n938), .B1(G68), .B2(new_n778), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n782), .A2(G137), .ZN(new_n940));
  NAND2_X1  g0740(.A1(new_n780), .A2(G143), .ZN(new_n941));
  OAI22_X1  g0741(.A1(new_n750), .A2(new_n202), .B1(new_n753), .B2(new_n201), .ZN(new_n942));
  AOI21_X1  g0742(.A(new_n942), .B1(G77), .B2(new_n824), .ZN(new_n943));
  NAND4_X1  g0743(.A1(new_n939), .A2(new_n940), .A3(new_n941), .A4(new_n943), .ZN(new_n944));
  OAI22_X1  g0744(.A1(new_n756), .A2(new_n773), .B1(new_n761), .B2(new_n419), .ZN(new_n945));
  AOI211_X1 g0745(.A(new_n376), .B(new_n945), .C1(G283), .C2(new_n754), .ZN(new_n946));
  XOR2_X1   g0746(.A(KEYINPUT106), .B(G317), .Z(new_n947));
  NAND2_X1  g0747(.A1(new_n782), .A2(new_n947), .ZN(new_n948));
  INV_X1    g0748(.A(KEYINPUT46), .ZN(new_n949));
  OAI21_X1  g0749(.A(new_n949), .B1(new_n750), .B2(new_n606), .ZN(new_n950));
  OR2_X1    g0750(.A1(new_n950), .A2(KEYINPUT105), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n950), .A2(KEYINPUT105), .ZN(new_n952));
  NAND4_X1  g0752(.A1(new_n946), .A2(new_n948), .A3(new_n951), .A4(new_n952), .ZN(new_n953));
  NOR3_X1   g0753(.A1(new_n750), .A2(new_n949), .A3(new_n606), .ZN(new_n954));
  AOI21_X1  g0754(.A(new_n954), .B1(G294), .B2(new_n763), .ZN(new_n955));
  OAI221_X1 g0755(.A(new_n955), .B1(new_n502), .B2(new_n759), .C1(new_n771), .C2(new_n785), .ZN(new_n956));
  OAI21_X1  g0756(.A(new_n944), .B1(new_n953), .B2(new_n956), .ZN(new_n957));
  INV_X1    g0757(.A(KEYINPUT47), .ZN(new_n958));
  OR2_X1    g0758(.A1(new_n957), .A2(new_n958), .ZN(new_n959));
  AOI21_X1  g0759(.A(new_n738), .B1(new_n957), .B2(new_n958), .ZN(new_n960));
  AOI21_X1  g0760(.A(new_n937), .B1(new_n959), .B2(new_n960), .ZN(new_n961));
  NAND2_X1  g0761(.A1(new_n933), .A2(new_n961), .ZN(new_n962));
  INV_X1    g0762(.A(KEYINPUT103), .ZN(new_n963));
  NAND2_X1  g0763(.A1(new_n672), .A2(new_n668), .ZN(new_n964));
  INV_X1    g0764(.A(new_n964), .ZN(new_n965));
  NAND2_X1  g0765(.A1(new_n965), .A2(new_n565), .ZN(new_n966));
  OAI21_X1  g0766(.A(new_n966), .B1(new_n671), .B2(new_n965), .ZN(new_n967));
  XNOR2_X1  g0767(.A(new_n967), .B(new_n676), .ZN(new_n968));
  NAND3_X1  g0768(.A1(new_n968), .A2(new_n711), .A3(new_n728), .ZN(new_n969));
  INV_X1    g0769(.A(new_n969), .ZN(new_n970));
  INV_X1    g0770(.A(new_n677), .ZN(new_n971));
  OR2_X1    g0771(.A1(new_n508), .A2(new_n668), .ZN(new_n972));
  NAND2_X1  g0772(.A1(new_n517), .A2(new_n972), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n510), .A2(new_n667), .ZN(new_n974));
  NAND2_X1  g0774(.A1(new_n973), .A2(new_n974), .ZN(new_n975));
  AND3_X1   g0775(.A1(new_n680), .A2(KEYINPUT45), .A3(new_n975), .ZN(new_n976));
  AOI21_X1  g0776(.A(KEYINPUT45), .B1(new_n680), .B2(new_n975), .ZN(new_n977));
  NOR2_X1   g0777(.A1(new_n976), .A2(new_n977), .ZN(new_n978));
  INV_X1    g0778(.A(new_n975), .ZN(new_n979));
  OAI21_X1  g0779(.A(new_n966), .B1(new_n670), .B2(new_n667), .ZN(new_n980));
  INV_X1    g0780(.A(KEYINPUT44), .ZN(new_n981));
  NAND3_X1  g0781(.A1(new_n979), .A2(new_n980), .A3(new_n981), .ZN(new_n982));
  OAI21_X1  g0782(.A(KEYINPUT44), .B1(new_n680), .B2(new_n975), .ZN(new_n983));
  NAND2_X1  g0783(.A1(new_n982), .A2(new_n983), .ZN(new_n984));
  OAI21_X1  g0784(.A(new_n971), .B1(new_n978), .B2(new_n984), .ZN(new_n985));
  INV_X1    g0785(.A(KEYINPUT45), .ZN(new_n986));
  OAI21_X1  g0786(.A(new_n986), .B1(new_n979), .B2(new_n980), .ZN(new_n987));
  NAND3_X1  g0787(.A1(new_n680), .A2(KEYINPUT45), .A3(new_n975), .ZN(new_n988));
  NAND2_X1  g0788(.A1(new_n987), .A2(new_n988), .ZN(new_n989));
  NAND4_X1  g0789(.A1(new_n989), .A2(new_n677), .A3(new_n983), .A4(new_n982), .ZN(new_n990));
  AND2_X1   g0790(.A1(new_n985), .A2(new_n990), .ZN(new_n991));
  AOI21_X1  g0791(.A(new_n963), .B1(new_n970), .B2(new_n991), .ZN(new_n992));
  NAND2_X1  g0792(.A1(new_n985), .A2(new_n990), .ZN(new_n993));
  NOR3_X1   g0793(.A1(new_n969), .A2(new_n993), .A3(KEYINPUT103), .ZN(new_n994));
  OAI21_X1  g0794(.A(new_n730), .B1(new_n992), .B2(new_n994), .ZN(new_n995));
  XNOR2_X1  g0795(.A(KEYINPUT102), .B(KEYINPUT41), .ZN(new_n996));
  XNOR2_X1  g0796(.A(new_n683), .B(new_n996), .ZN(new_n997));
  INV_X1    g0797(.A(new_n997), .ZN(new_n998));
  AOI21_X1  g0798(.A(new_n734), .B1(new_n995), .B2(new_n998), .ZN(new_n999));
  OR2_X1    g0799(.A1(new_n973), .A2(new_n670), .ZN(new_n1000));
  INV_X1    g0800(.A(new_n510), .ZN(new_n1001));
  AOI21_X1  g0801(.A(new_n667), .B1(new_n1000), .B2(new_n1001), .ZN(new_n1002));
  NAND2_X1  g0802(.A1(new_n975), .A2(new_n678), .ZN(new_n1003));
  AOI21_X1  g0803(.A(new_n1002), .B1(KEYINPUT42), .B2(new_n1003), .ZN(new_n1004));
  OR2_X1    g0804(.A1(new_n1003), .A2(KEYINPUT42), .ZN(new_n1005));
  AOI22_X1  g0805(.A1(new_n1004), .A2(new_n1005), .B1(KEYINPUT43), .B2(new_n932), .ZN(new_n1006));
  OR2_X1    g0806(.A1(new_n932), .A2(KEYINPUT43), .ZN(new_n1007));
  XNOR2_X1  g0807(.A(new_n1006), .B(new_n1007), .ZN(new_n1008));
  NOR2_X1   g0808(.A1(new_n677), .A2(new_n979), .ZN(new_n1009));
  INV_X1    g0809(.A(new_n1009), .ZN(new_n1010));
  XNOR2_X1  g0810(.A(new_n1008), .B(new_n1010), .ZN(new_n1011));
  OAI21_X1  g0811(.A(new_n962), .B1(new_n999), .B2(new_n1011), .ZN(G387));
  INV_X1    g0812(.A(KEYINPUT109), .ZN(new_n1013));
  OAI21_X1  g0813(.A(new_n1013), .B1(new_n730), .B2(new_n968), .ZN(new_n1014));
  INV_X1    g0814(.A(new_n968), .ZN(new_n1015));
  NAND3_X1  g0815(.A1(new_n1015), .A2(new_n729), .A3(KEYINPUT109), .ZN(new_n1016));
  NAND4_X1  g0816(.A1(new_n1014), .A2(new_n683), .A3(new_n969), .A4(new_n1016), .ZN(new_n1017));
  NOR2_X1   g0817(.A1(new_n671), .A2(new_n808), .ZN(new_n1018));
  NAND2_X1  g0818(.A1(new_n237), .A2(G45), .ZN(new_n1019));
  XNOR2_X1  g0819(.A(new_n1019), .B(KEYINPUT107), .ZN(new_n1020));
  XNOR2_X1  g0820(.A(KEYINPUT108), .B(KEYINPUT50), .ZN(new_n1021));
  INV_X1    g0821(.A(new_n1021), .ZN(new_n1022));
  OAI21_X1  g0822(.A(new_n1022), .B1(G50), .B2(new_n288), .ZN(new_n1023));
  NAND3_X1  g0823(.A1(new_n286), .A2(new_n1021), .A3(new_n201), .ZN(new_n1024));
  AOI21_X1  g0824(.A(G45), .B1(G68), .B2(G77), .ZN(new_n1025));
  AND4_X1   g0825(.A1(new_n685), .A2(new_n1023), .A3(new_n1024), .A4(new_n1025), .ZN(new_n1026));
  NOR3_X1   g0826(.A1(new_n1020), .A2(new_n802), .A3(new_n1026), .ZN(new_n1027));
  OAI22_X1  g0827(.A1(new_n795), .A2(new_n685), .B1(G107), .B2(new_n211), .ZN(new_n1028));
  OAI21_X1  g0828(.A(new_n794), .B1(new_n1027), .B2(new_n1028), .ZN(new_n1029));
  NAND2_X1  g0829(.A1(new_n1029), .A2(new_n735), .ZN(new_n1030));
  OAI22_X1  g0830(.A1(new_n756), .A2(new_n201), .B1(new_n753), .B2(new_n203), .ZN(new_n1031));
  OAI221_X1 g0831(.A(new_n376), .B1(new_n761), .B2(new_n419), .C1(new_n764), .C2(new_n288), .ZN(new_n1032));
  AOI211_X1 g0832(.A(new_n1031), .B(new_n1032), .C1(G77), .C2(new_n751), .ZN(new_n1033));
  NAND2_X1  g0833(.A1(new_n780), .A2(G159), .ZN(new_n1034));
  NAND2_X1  g0834(.A1(new_n782), .A2(G150), .ZN(new_n1035));
  NAND2_X1  g0835(.A1(new_n596), .A2(new_n597), .ZN(new_n1036));
  INV_X1    g0836(.A(new_n1036), .ZN(new_n1037));
  NAND2_X1  g0837(.A1(new_n1037), .A2(new_n778), .ZN(new_n1038));
  NAND4_X1  g0838(.A1(new_n1033), .A2(new_n1034), .A3(new_n1035), .A4(new_n1038), .ZN(new_n1039));
  NAND2_X1  g0839(.A1(new_n782), .A2(G326), .ZN(new_n1040));
  AOI21_X1  g0840(.A(new_n376), .B1(new_n824), .B2(G116), .ZN(new_n1041));
  OAI22_X1  g0841(.A1(new_n759), .A2(new_n784), .B1(new_n750), .B2(new_n832), .ZN(new_n1042));
  AOI22_X1  g0842(.A1(new_n787), .A2(new_n947), .B1(new_n754), .B2(G303), .ZN(new_n1043));
  INV_X1    g0843(.A(G322), .ZN(new_n1044));
  OAI221_X1 g0844(.A(new_n1043), .B1(new_n785), .B2(new_n764), .C1(new_n771), .C2(new_n1044), .ZN(new_n1045));
  INV_X1    g0845(.A(KEYINPUT48), .ZN(new_n1046));
  AOI21_X1  g0846(.A(new_n1042), .B1(new_n1045), .B2(new_n1046), .ZN(new_n1047));
  OAI21_X1  g0847(.A(new_n1047), .B1(new_n1046), .B2(new_n1045), .ZN(new_n1048));
  INV_X1    g0848(.A(KEYINPUT49), .ZN(new_n1049));
  OAI211_X1 g0849(.A(new_n1040), .B(new_n1041), .C1(new_n1048), .C2(new_n1049), .ZN(new_n1050));
  AND2_X1   g0850(.A1(new_n1048), .A2(new_n1049), .ZN(new_n1051));
  OAI21_X1  g0851(.A(new_n1039), .B1(new_n1050), .B2(new_n1051), .ZN(new_n1052));
  AOI211_X1 g0852(.A(new_n1018), .B(new_n1030), .C1(new_n737), .C2(new_n1052), .ZN(new_n1053));
  AOI21_X1  g0853(.A(new_n1053), .B1(new_n734), .B2(new_n968), .ZN(new_n1054));
  NAND2_X1  g0854(.A1(new_n1017), .A2(new_n1054), .ZN(G393));
  NAND3_X1  g0855(.A1(new_n970), .A2(new_n991), .A3(new_n963), .ZN(new_n1056));
  OAI21_X1  g0856(.A(KEYINPUT103), .B1(new_n969), .B2(new_n993), .ZN(new_n1057));
  NAND2_X1  g0857(.A1(new_n1056), .A2(new_n1057), .ZN(new_n1058));
  INV_X1    g0858(.A(KEYINPUT110), .ZN(new_n1059));
  NAND2_X1  g0859(.A1(new_n990), .A2(new_n1059), .ZN(new_n1060));
  XOR2_X1   g0860(.A(new_n1060), .B(new_n985), .Z(new_n1061));
  OAI211_X1 g0861(.A(new_n683), .B(new_n1058), .C1(new_n1061), .C2(new_n970), .ZN(new_n1062));
  NAND2_X1  g0862(.A1(new_n979), .A2(new_n793), .ZN(new_n1063));
  NOR2_X1   g0863(.A1(new_n802), .A2(new_n247), .ZN(new_n1064));
  OAI21_X1  g0864(.A(new_n794), .B1(new_n419), .B2(new_n211), .ZN(new_n1065));
  OAI22_X1  g0865(.A1(new_n771), .A2(new_n366), .B1(new_n745), .B2(new_n756), .ZN(new_n1066));
  XOR2_X1   g0866(.A(new_n1066), .B(KEYINPUT111), .Z(new_n1067));
  XNOR2_X1  g0867(.A(new_n1067), .B(KEYINPUT51), .ZN(new_n1068));
  NAND2_X1  g0868(.A1(new_n778), .A2(G77), .ZN(new_n1069));
  OAI21_X1  g0869(.A(new_n1069), .B1(new_n764), .B2(new_n201), .ZN(new_n1070));
  AOI21_X1  g0870(.A(new_n252), .B1(new_n824), .B2(G87), .ZN(new_n1071));
  OAI221_X1 g0871(.A(new_n1071), .B1(new_n203), .B2(new_n750), .C1(new_n288), .C2(new_n753), .ZN(new_n1072));
  AOI211_X1 g0872(.A(new_n1070), .B(new_n1072), .C1(G143), .C2(new_n782), .ZN(new_n1073));
  AOI22_X1  g0873(.A1(new_n780), .A2(G317), .B1(G311), .B2(new_n787), .ZN(new_n1074));
  XOR2_X1   g0874(.A(new_n1074), .B(KEYINPUT52), .Z(new_n1075));
  OAI22_X1  g0875(.A1(new_n759), .A2(new_n606), .B1(new_n764), .B2(new_n773), .ZN(new_n1076));
  AOI21_X1  g0876(.A(new_n376), .B1(new_n824), .B2(G107), .ZN(new_n1077));
  OAI221_X1 g0877(.A(new_n1077), .B1(new_n784), .B2(new_n750), .C1(new_n832), .C2(new_n753), .ZN(new_n1078));
  AOI211_X1 g0878(.A(new_n1076), .B(new_n1078), .C1(G322), .C2(new_n782), .ZN(new_n1079));
  AOI22_X1  g0879(.A1(new_n1068), .A2(new_n1073), .B1(new_n1075), .B2(new_n1079), .ZN(new_n1080));
  OAI221_X1 g0880(.A(new_n735), .B1(new_n1064), .B2(new_n1065), .C1(new_n1080), .C2(new_n738), .ZN(new_n1081));
  XNOR2_X1  g0881(.A(new_n1081), .B(KEYINPUT112), .ZN(new_n1082));
  AOI22_X1  g0882(.A1(new_n1061), .A2(new_n734), .B1(new_n1063), .B2(new_n1082), .ZN(new_n1083));
  NAND2_X1  g0883(.A1(new_n1062), .A2(new_n1083), .ZN(G390));
  INV_X1    g0884(.A(KEYINPUT113), .ZN(new_n1085));
  NAND2_X1  g0885(.A1(new_n880), .A2(new_n908), .ZN(new_n1086));
  INV_X1    g0886(.A(new_n722), .ZN(new_n1087));
  OAI211_X1 g0887(.A(new_n668), .B(new_n815), .C1(new_n1087), .C2(new_n646), .ZN(new_n1088));
  AOI21_X1  g0888(.A(new_n901), .B1(new_n1088), .B2(new_n816), .ZN(new_n1089));
  OAI21_X1  g0889(.A(new_n1085), .B1(new_n1086), .B2(new_n1089), .ZN(new_n1090));
  INV_X1    g0890(.A(new_n815), .ZN(new_n1091));
  AOI211_X1 g0891(.A(new_n667), .B(new_n1091), .C1(new_n714), .C2(new_n722), .ZN(new_n1092));
  INV_X1    g0892(.A(new_n816), .ZN(new_n1093));
  OAI21_X1  g0893(.A(new_n900), .B1(new_n1092), .B2(new_n1093), .ZN(new_n1094));
  NAND4_X1  g0894(.A1(new_n1094), .A2(KEYINPUT113), .A3(new_n908), .A4(new_n880), .ZN(new_n1095));
  NAND2_X1  g0895(.A1(new_n1090), .A2(new_n1095), .ZN(new_n1096));
  OAI211_X1 g0896(.A(new_n904), .B(new_n906), .C1(new_n902), .C2(new_n909), .ZN(new_n1097));
  OAI211_X1 g0897(.A(new_n819), .B(new_n900), .C1(new_n709), .C2(new_n710), .ZN(new_n1098));
  NAND3_X1  g0898(.A1(new_n1096), .A2(new_n1097), .A3(new_n1098), .ZN(new_n1099));
  AND2_X1   g0899(.A1(new_n1096), .A2(new_n1097), .ZN(new_n1100));
  NAND2_X1  g0900(.A1(new_n851), .A2(G330), .ZN(new_n1101));
  NOR3_X1   g0901(.A1(new_n1101), .A2(new_n901), .A3(new_n817), .ZN(new_n1102));
  INV_X1    g0902(.A(new_n1102), .ZN(new_n1103));
  OAI21_X1  g0903(.A(new_n1099), .B1(new_n1100), .B2(new_n1103), .ZN(new_n1104));
  INV_X1    g0904(.A(new_n1101), .ZN(new_n1105));
  OAI21_X1  g0905(.A(new_n1105), .B1(new_n465), .B2(new_n469), .ZN(new_n1106));
  NAND3_X1  g0906(.A1(new_n912), .A2(new_n660), .A3(new_n1106), .ZN(new_n1107));
  NAND2_X1  g0907(.A1(new_n708), .A2(G330), .ZN(new_n1108));
  INV_X1    g0908(.A(KEYINPUT88), .ZN(new_n1109));
  NAND2_X1  g0909(.A1(new_n1108), .A2(new_n1109), .ZN(new_n1110));
  NAND3_X1  g0910(.A1(new_n708), .A2(KEYINPUT88), .A3(G330), .ZN(new_n1111));
  AOI21_X1  g0911(.A(new_n817), .B1(new_n1110), .B2(new_n1111), .ZN(new_n1112));
  OAI21_X1  g0912(.A(new_n1103), .B1(new_n1112), .B2(new_n900), .ZN(new_n1113));
  NAND2_X1  g0913(.A1(new_n1113), .A2(new_n898), .ZN(new_n1114));
  AOI21_X1  g0914(.A(new_n1093), .B1(new_n723), .B2(new_n815), .ZN(new_n1115));
  OAI21_X1  g0915(.A(new_n901), .B1(new_n1101), .B2(new_n817), .ZN(new_n1116));
  NAND3_X1  g0916(.A1(new_n1098), .A2(new_n1115), .A3(new_n1116), .ZN(new_n1117));
  AOI21_X1  g0917(.A(new_n1107), .B1(new_n1114), .B2(new_n1117), .ZN(new_n1118));
  INV_X1    g0918(.A(new_n1118), .ZN(new_n1119));
  AOI21_X1  g0919(.A(new_n684), .B1(new_n1104), .B2(new_n1119), .ZN(new_n1120));
  OAI211_X1 g0920(.A(new_n1099), .B(new_n1118), .C1(new_n1100), .C2(new_n1103), .ZN(new_n1121));
  NAND2_X1  g0921(.A1(new_n1120), .A2(new_n1121), .ZN(new_n1122));
  AOI21_X1  g0922(.A(new_n736), .B1(new_n288), .B2(new_n840), .ZN(new_n1123));
  XOR2_X1   g0923(.A(new_n1123), .B(KEYINPUT114), .Z(new_n1124));
  NAND2_X1  g0924(.A1(new_n782), .A2(G125), .ZN(new_n1125));
  NOR2_X1   g0925(.A1(new_n761), .A2(new_n201), .ZN(new_n1126));
  INV_X1    g0926(.A(G132), .ZN(new_n1127));
  OAI21_X1  g0927(.A(new_n376), .B1(new_n756), .B2(new_n1127), .ZN(new_n1128));
  AOI211_X1 g0928(.A(new_n1126), .B(new_n1128), .C1(G159), .C2(new_n778), .ZN(new_n1129));
  NAND2_X1  g0929(.A1(new_n780), .A2(G128), .ZN(new_n1130));
  NOR2_X1   g0930(.A1(new_n750), .A2(new_n366), .ZN(new_n1131));
  XNOR2_X1  g0931(.A(new_n1131), .B(KEYINPUT53), .ZN(new_n1132));
  NAND4_X1  g0932(.A1(new_n1125), .A2(new_n1129), .A3(new_n1130), .A4(new_n1132), .ZN(new_n1133));
  XNOR2_X1  g0933(.A(KEYINPUT54), .B(G143), .ZN(new_n1134));
  OAI22_X1  g0934(.A1(new_n764), .A2(new_n828), .B1(new_n753), .B2(new_n1134), .ZN(new_n1135));
  XNOR2_X1  g0935(.A(new_n1135), .B(KEYINPUT115), .ZN(new_n1136));
  NAND2_X1  g0936(.A1(new_n782), .A2(G294), .ZN(new_n1137));
  AOI21_X1  g0937(.A(new_n376), .B1(new_n751), .B2(G87), .ZN(new_n1138));
  AOI22_X1  g0938(.A1(new_n787), .A2(G116), .B1(new_n824), .B2(G68), .ZN(new_n1139));
  NAND4_X1  g0939(.A1(new_n1137), .A2(new_n1069), .A3(new_n1138), .A4(new_n1139), .ZN(new_n1140));
  OAI22_X1  g0940(.A1(new_n764), .A2(new_n502), .B1(new_n753), .B2(new_n419), .ZN(new_n1141));
  AOI22_X1  g0941(.A1(new_n780), .A2(G283), .B1(KEYINPUT116), .B2(new_n1141), .ZN(new_n1142));
  OAI21_X1  g0942(.A(new_n1142), .B1(KEYINPUT116), .B2(new_n1141), .ZN(new_n1143));
  OAI22_X1  g0943(.A1(new_n1133), .A2(new_n1136), .B1(new_n1140), .B2(new_n1143), .ZN(new_n1144));
  AOI21_X1  g0944(.A(new_n1124), .B1(new_n1144), .B2(new_n737), .ZN(new_n1145));
  OAI21_X1  g0945(.A(new_n1145), .B1(new_n907), .B2(new_n792), .ZN(new_n1146));
  XNOR2_X1  g0946(.A(new_n1146), .B(KEYINPUT117), .ZN(new_n1147));
  AND3_X1   g0947(.A1(new_n1096), .A2(new_n1097), .A3(new_n1098), .ZN(new_n1148));
  AOI21_X1  g0948(.A(new_n1103), .B1(new_n1096), .B2(new_n1097), .ZN(new_n1149));
  NOR2_X1   g0949(.A1(new_n1148), .A2(new_n1149), .ZN(new_n1150));
  NAND2_X1  g0950(.A1(new_n1150), .A2(new_n734), .ZN(new_n1151));
  NAND3_X1  g0951(.A1(new_n1122), .A2(new_n1147), .A3(new_n1151), .ZN(G378));
  INV_X1    g0952(.A(KEYINPUT57), .ZN(new_n1153));
  OAI21_X1  g0953(.A(new_n819), .B1(new_n709), .B2(new_n710), .ZN(new_n1154));
  AOI21_X1  g0954(.A(new_n1102), .B1(new_n1154), .B2(new_n901), .ZN(new_n1155));
  OAI21_X1  g0955(.A(new_n1117), .B1(new_n1155), .B2(new_n899), .ZN(new_n1156));
  AOI21_X1  g0956(.A(new_n1107), .B1(new_n1150), .B2(new_n1156), .ZN(new_n1157));
  NAND2_X1  g0957(.A1(new_n887), .A2(new_n891), .ZN(new_n1158));
  INV_X1    g0958(.A(new_n881), .ZN(new_n1159));
  NAND2_X1  g0959(.A1(new_n372), .A2(new_n856), .ZN(new_n1160));
  XNOR2_X1  g0960(.A(new_n1160), .B(KEYINPUT55), .ZN(new_n1161));
  XNOR2_X1  g0961(.A(new_n466), .B(new_n1161), .ZN(new_n1162));
  XNOR2_X1  g0962(.A(KEYINPUT119), .B(KEYINPUT56), .ZN(new_n1163));
  XNOR2_X1  g0963(.A(new_n1162), .B(new_n1163), .ZN(new_n1164));
  INV_X1    g0964(.A(new_n1164), .ZN(new_n1165));
  AND4_X1   g0965(.A1(G330), .A2(new_n1158), .A3(new_n1159), .A4(new_n1165), .ZN(new_n1166));
  AOI21_X1  g0966(.A(new_n1165), .B1(new_n892), .B2(G330), .ZN(new_n1167));
  OAI21_X1  g0967(.A(new_n911), .B1(new_n1166), .B2(new_n1167), .ZN(new_n1168));
  NAND3_X1  g0968(.A1(new_n1158), .A2(G330), .A3(new_n1159), .ZN(new_n1169));
  NAND2_X1  g0969(.A1(new_n1169), .A2(new_n1164), .ZN(new_n1170));
  INV_X1    g0970(.A(new_n911), .ZN(new_n1171));
  NAND3_X1  g0971(.A1(new_n892), .A2(G330), .A3(new_n1165), .ZN(new_n1172));
  NAND3_X1  g0972(.A1(new_n1170), .A2(new_n1171), .A3(new_n1172), .ZN(new_n1173));
  NAND2_X1  g0973(.A1(new_n1168), .A2(new_n1173), .ZN(new_n1174));
  OAI21_X1  g0974(.A(new_n1153), .B1(new_n1157), .B2(new_n1174), .ZN(new_n1175));
  INV_X1    g0975(.A(new_n1107), .ZN(new_n1176));
  NAND2_X1  g0976(.A1(new_n1121), .A2(new_n1176), .ZN(new_n1177));
  NAND4_X1  g0977(.A1(new_n1177), .A2(KEYINPUT57), .A3(new_n1173), .A4(new_n1168), .ZN(new_n1178));
  NAND3_X1  g0978(.A1(new_n1175), .A2(new_n683), .A3(new_n1178), .ZN(new_n1179));
  NAND3_X1  g0979(.A1(new_n1168), .A2(new_n1173), .A3(new_n734), .ZN(new_n1180));
  AOI21_X1  g0980(.A(new_n736), .B1(new_n201), .B2(new_n840), .ZN(new_n1181));
  OAI22_X1  g0981(.A1(new_n756), .A2(new_n502), .B1(new_n761), .B2(new_n202), .ZN(new_n1182));
  INV_X1    g0982(.A(new_n485), .ZN(new_n1183));
  OAI211_X1 g0983(.A(new_n1183), .B(new_n252), .C1(new_n750), .C2(new_n221), .ZN(new_n1184));
  AOI211_X1 g0984(.A(new_n1182), .B(new_n1184), .C1(G97), .C2(new_n763), .ZN(new_n1185));
  OAI221_X1 g0985(.A(new_n1185), .B1(new_n784), .B2(new_n744), .C1(new_n1036), .C2(new_n753), .ZN(new_n1186));
  OAI22_X1  g0986(.A1(new_n771), .A2(new_n606), .B1(new_n203), .B2(new_n759), .ZN(new_n1187));
  XOR2_X1   g0987(.A(new_n1187), .B(KEYINPUT118), .Z(new_n1188));
  NOR2_X1   g0988(.A1(new_n1186), .A2(new_n1188), .ZN(new_n1189));
  OR2_X1    g0989(.A1(new_n1189), .A2(KEYINPUT58), .ZN(new_n1190));
  OAI221_X1 g0990(.A(new_n201), .B1(G33), .B2(G41), .C1(new_n376), .C2(new_n485), .ZN(new_n1191));
  NAND2_X1  g0991(.A1(new_n780), .A2(G125), .ZN(new_n1192));
  INV_X1    g0992(.A(G128), .ZN(new_n1193));
  OAI22_X1  g0993(.A1(new_n1193), .A2(new_n756), .B1(new_n750), .B2(new_n1134), .ZN(new_n1194));
  AOI21_X1  g0994(.A(new_n1194), .B1(G137), .B2(new_n754), .ZN(new_n1195));
  AOI22_X1  g0995(.A1(new_n778), .A2(G150), .B1(new_n763), .B2(G132), .ZN(new_n1196));
  NAND3_X1  g0996(.A1(new_n1192), .A2(new_n1195), .A3(new_n1196), .ZN(new_n1197));
  OR2_X1    g0997(.A1(new_n1197), .A2(KEYINPUT59), .ZN(new_n1198));
  NAND2_X1  g0998(.A1(new_n1197), .A2(KEYINPUT59), .ZN(new_n1199));
  NAND2_X1  g0999(.A1(new_n782), .A2(G124), .ZN(new_n1200));
  AOI211_X1 g1000(.A(G33), .B(G41), .C1(new_n824), .C2(G159), .ZN(new_n1201));
  NAND4_X1  g1001(.A1(new_n1198), .A2(new_n1199), .A3(new_n1200), .A4(new_n1201), .ZN(new_n1202));
  NAND3_X1  g1002(.A1(new_n1190), .A2(new_n1191), .A3(new_n1202), .ZN(new_n1203));
  AOI21_X1  g1003(.A(new_n1203), .B1(KEYINPUT58), .B2(new_n1189), .ZN(new_n1204));
  OAI221_X1 g1004(.A(new_n1181), .B1(new_n738), .B2(new_n1204), .C1(new_n1164), .C2(new_n792), .ZN(new_n1205));
  NAND2_X1  g1005(.A1(new_n1180), .A2(new_n1205), .ZN(new_n1206));
  INV_X1    g1006(.A(new_n1206), .ZN(new_n1207));
  NAND2_X1  g1007(.A1(new_n1179), .A2(new_n1207), .ZN(G375));
  INV_X1    g1008(.A(KEYINPUT120), .ZN(new_n1209));
  AND2_X1   g1009(.A1(new_n1116), .A2(new_n1115), .ZN(new_n1210));
  AOI22_X1  g1010(.A1(new_n1113), .A2(new_n898), .B1(new_n1098), .B2(new_n1210), .ZN(new_n1211));
  OAI21_X1  g1011(.A(new_n1209), .B1(new_n1211), .B2(new_n733), .ZN(new_n1212));
  NAND3_X1  g1012(.A1(new_n1156), .A2(KEYINPUT120), .A3(new_n734), .ZN(new_n1213));
  OAI22_X1  g1013(.A1(new_n764), .A2(new_n1134), .B1(new_n756), .B2(new_n828), .ZN(new_n1214));
  OAI22_X1  g1014(.A1(new_n750), .A2(new_n745), .B1(new_n753), .B2(new_n366), .ZN(new_n1215));
  AOI211_X1 g1015(.A(new_n252), .B(new_n1215), .C1(G58), .C2(new_n824), .ZN(new_n1216));
  OAI221_X1 g1016(.A(new_n1216), .B1(new_n201), .B2(new_n759), .C1(new_n1193), .C2(new_n744), .ZN(new_n1217));
  XOR2_X1   g1017(.A(new_n1217), .B(KEYINPUT121), .Z(new_n1218));
  AOI211_X1 g1018(.A(new_n1214), .B(new_n1218), .C1(G132), .C2(new_n780), .ZN(new_n1219));
  OAI21_X1  g1019(.A(new_n1038), .B1(new_n773), .B2(new_n744), .ZN(new_n1220));
  NOR2_X1   g1020(.A1(new_n771), .A2(new_n832), .ZN(new_n1221));
  AOI22_X1  g1021(.A1(G97), .A2(new_n751), .B1(new_n787), .B2(G283), .ZN(new_n1222));
  OAI21_X1  g1022(.A(new_n1222), .B1(new_n502), .B2(new_n753), .ZN(new_n1223));
  OAI221_X1 g1023(.A(new_n252), .B1(new_n761), .B2(new_n221), .C1(new_n764), .C2(new_n606), .ZN(new_n1224));
  NOR4_X1   g1024(.A1(new_n1220), .A2(new_n1221), .A3(new_n1223), .A4(new_n1224), .ZN(new_n1225));
  OAI21_X1  g1025(.A(new_n737), .B1(new_n1219), .B2(new_n1225), .ZN(new_n1226));
  AOI21_X1  g1026(.A(new_n736), .B1(new_n203), .B2(new_n840), .ZN(new_n1227));
  NAND2_X1  g1027(.A1(new_n1226), .A2(new_n1227), .ZN(new_n1228));
  AOI21_X1  g1028(.A(new_n1228), .B1(new_n791), .B2(new_n901), .ZN(new_n1229));
  INV_X1    g1029(.A(new_n1229), .ZN(new_n1230));
  NAND3_X1  g1030(.A1(new_n1212), .A2(new_n1213), .A3(new_n1230), .ZN(new_n1231));
  INV_X1    g1031(.A(new_n1231), .ZN(new_n1232));
  OAI211_X1 g1032(.A(new_n1107), .B(new_n1117), .C1(new_n1155), .C2(new_n899), .ZN(new_n1233));
  NAND3_X1  g1033(.A1(new_n1119), .A2(new_n998), .A3(new_n1233), .ZN(new_n1234));
  NAND2_X1  g1034(.A1(new_n1232), .A2(new_n1234), .ZN(G381));
  NOR2_X1   g1035(.A1(G375), .A2(G378), .ZN(new_n1236));
  INV_X1    g1036(.A(new_n962), .ZN(new_n1237));
  AOI21_X1  g1037(.A(new_n729), .B1(new_n1056), .B2(new_n1057), .ZN(new_n1238));
  OAI21_X1  g1038(.A(new_n733), .B1(new_n1238), .B2(new_n997), .ZN(new_n1239));
  XNOR2_X1  g1039(.A(new_n1008), .B(new_n1009), .ZN(new_n1240));
  AOI21_X1  g1040(.A(new_n1237), .B1(new_n1239), .B2(new_n1240), .ZN(new_n1241));
  INV_X1    g1041(.A(G396), .ZN(new_n1242));
  NAND3_X1  g1042(.A1(new_n1017), .A2(new_n1242), .A3(new_n1054), .ZN(new_n1243));
  NOR4_X1   g1043(.A1(G381), .A2(G390), .A3(new_n1243), .A4(G384), .ZN(new_n1244));
  NAND3_X1  g1044(.A1(new_n1236), .A2(new_n1241), .A3(new_n1244), .ZN(G407));
  NAND2_X1  g1045(.A1(new_n666), .A2(G213), .ZN(new_n1246));
  INV_X1    g1046(.A(new_n1246), .ZN(new_n1247));
  NAND2_X1  g1047(.A1(new_n1236), .A2(new_n1247), .ZN(new_n1248));
  NAND3_X1  g1048(.A1(G407), .A2(G213), .A3(new_n1248), .ZN(G409));
  INV_X1    g1049(.A(KEYINPUT61), .ZN(new_n1250));
  INV_X1    g1050(.A(KEYINPUT125), .ZN(new_n1251));
  INV_X1    g1051(.A(G390), .ZN(new_n1252));
  NAND2_X1  g1052(.A1(G387), .A2(new_n1252), .ZN(new_n1253));
  NAND2_X1  g1053(.A1(new_n1241), .A2(G390), .ZN(new_n1254));
  XNOR2_X1  g1054(.A(G393), .B(new_n1242), .ZN(new_n1255));
  AND4_X1   g1055(.A1(new_n1251), .A2(new_n1253), .A3(new_n1254), .A4(new_n1255), .ZN(new_n1256));
  OAI21_X1  g1056(.A(KEYINPUT125), .B1(new_n1241), .B2(G390), .ZN(new_n1257));
  AOI22_X1  g1057(.A1(new_n1257), .A2(new_n1255), .B1(new_n1253), .B2(new_n1254), .ZN(new_n1258));
  NOR2_X1   g1058(.A1(new_n1256), .A2(new_n1258), .ZN(new_n1259));
  NAND3_X1  g1059(.A1(new_n1179), .A2(G378), .A3(new_n1207), .ZN(new_n1260));
  NAND2_X1  g1060(.A1(new_n1151), .A2(new_n1147), .ZN(new_n1261));
  AOI21_X1  g1061(.A(new_n1261), .B1(new_n1121), .B2(new_n1120), .ZN(new_n1262));
  NOR3_X1   g1062(.A1(new_n1157), .A2(new_n1174), .A3(new_n997), .ZN(new_n1263));
  OAI21_X1  g1063(.A(new_n1262), .B1(new_n1206), .B2(new_n1263), .ZN(new_n1264));
  AOI21_X1  g1064(.A(new_n1247), .B1(new_n1260), .B2(new_n1264), .ZN(new_n1265));
  NAND2_X1  g1065(.A1(new_n1247), .A2(G2897), .ZN(new_n1266));
  INV_X1    g1066(.A(new_n1266), .ZN(new_n1267));
  INV_X1    g1067(.A(KEYINPUT122), .ZN(new_n1268));
  NAND2_X1  g1068(.A1(new_n1233), .A2(new_n1268), .ZN(new_n1269));
  NAND2_X1  g1069(.A1(new_n1269), .A2(KEYINPUT60), .ZN(new_n1270));
  INV_X1    g1070(.A(KEYINPUT60), .ZN(new_n1271));
  NAND3_X1  g1071(.A1(new_n1233), .A2(new_n1268), .A3(new_n1271), .ZN(new_n1272));
  AOI21_X1  g1072(.A(new_n684), .B1(new_n1156), .B2(new_n1176), .ZN(new_n1273));
  NAND3_X1  g1073(.A1(new_n1270), .A2(new_n1272), .A3(new_n1273), .ZN(new_n1274));
  NAND3_X1  g1074(.A1(new_n1232), .A2(new_n1274), .A3(G384), .ZN(new_n1275));
  AOI21_X1  g1075(.A(G384), .B1(new_n1232), .B2(new_n1274), .ZN(new_n1276));
  INV_X1    g1076(.A(KEYINPUT123), .ZN(new_n1277));
  OAI21_X1  g1077(.A(new_n1275), .B1(new_n1276), .B2(new_n1277), .ZN(new_n1278));
  AND2_X1   g1078(.A1(new_n1272), .A2(new_n1273), .ZN(new_n1279));
  AOI21_X1  g1079(.A(new_n1231), .B1(new_n1279), .B2(new_n1270), .ZN(new_n1280));
  NOR3_X1   g1080(.A1(new_n1280), .A2(KEYINPUT123), .A3(G384), .ZN(new_n1281));
  OAI21_X1  g1081(.A(new_n1267), .B1(new_n1278), .B2(new_n1281), .ZN(new_n1282));
  OAI21_X1  g1082(.A(KEYINPUT123), .B1(new_n1280), .B2(G384), .ZN(new_n1283));
  NAND2_X1  g1083(.A1(new_n1232), .A2(new_n1274), .ZN(new_n1284));
  INV_X1    g1084(.A(G384), .ZN(new_n1285));
  NAND3_X1  g1085(.A1(new_n1284), .A2(new_n1277), .A3(new_n1285), .ZN(new_n1286));
  NAND4_X1  g1086(.A1(new_n1283), .A2(new_n1286), .A3(new_n1275), .A4(new_n1266), .ZN(new_n1287));
  NAND2_X1  g1087(.A1(new_n1282), .A2(new_n1287), .ZN(new_n1288));
  OAI211_X1 g1088(.A(new_n1250), .B(new_n1259), .C1(new_n1265), .C2(new_n1288), .ZN(new_n1289));
  INV_X1    g1089(.A(new_n1289), .ZN(new_n1290));
  NAND3_X1  g1090(.A1(new_n1283), .A2(new_n1286), .A3(new_n1275), .ZN(new_n1291));
  AOI211_X1 g1091(.A(new_n1247), .B(new_n1291), .C1(new_n1260), .C2(new_n1264), .ZN(new_n1292));
  OAI21_X1  g1092(.A(KEYINPUT63), .B1(new_n1292), .B2(KEYINPUT124), .ZN(new_n1293));
  INV_X1    g1093(.A(new_n1291), .ZN(new_n1294));
  NAND2_X1  g1094(.A1(new_n1265), .A2(new_n1294), .ZN(new_n1295));
  INV_X1    g1095(.A(KEYINPUT124), .ZN(new_n1296));
  INV_X1    g1096(.A(KEYINPUT63), .ZN(new_n1297));
  NAND3_X1  g1097(.A1(new_n1295), .A2(new_n1296), .A3(new_n1297), .ZN(new_n1298));
  NAND3_X1  g1098(.A1(new_n1290), .A2(new_n1293), .A3(new_n1298), .ZN(new_n1299));
  XNOR2_X1  g1099(.A(KEYINPUT126), .B(KEYINPUT62), .ZN(new_n1300));
  AND3_X1   g1100(.A1(new_n1265), .A2(new_n1294), .A3(new_n1300), .ZN(new_n1301));
  OAI21_X1  g1101(.A(new_n1250), .B1(new_n1265), .B2(new_n1288), .ZN(new_n1302));
  INV_X1    g1102(.A(KEYINPUT126), .ZN(new_n1303));
  NAND2_X1  g1103(.A1(new_n1303), .A2(KEYINPUT62), .ZN(new_n1304));
  AOI21_X1  g1104(.A(new_n1304), .B1(new_n1265), .B2(new_n1294), .ZN(new_n1305));
  NOR3_X1   g1105(.A1(new_n1301), .A2(new_n1302), .A3(new_n1305), .ZN(new_n1306));
  OAI21_X1  g1106(.A(new_n1299), .B1(new_n1306), .B2(new_n1259), .ZN(G405));
  NAND2_X1  g1107(.A1(G375), .A2(new_n1262), .ZN(new_n1308));
  AOI21_X1  g1108(.A(KEYINPUT127), .B1(new_n1308), .B2(new_n1260), .ZN(new_n1309));
  NOR2_X1   g1109(.A1(new_n1309), .A2(new_n1294), .ZN(new_n1310));
  NAND2_X1  g1110(.A1(new_n1257), .A2(new_n1255), .ZN(new_n1311));
  NAND2_X1  g1111(.A1(new_n1253), .A2(new_n1254), .ZN(new_n1312));
  XNOR2_X1  g1112(.A(new_n1311), .B(new_n1312), .ZN(new_n1313));
  NAND4_X1  g1113(.A1(new_n1313), .A2(KEYINPUT127), .A3(new_n1260), .A4(new_n1308), .ZN(new_n1314));
  NAND3_X1  g1114(.A1(new_n1308), .A2(KEYINPUT127), .A3(new_n1260), .ZN(new_n1315));
  NAND2_X1  g1115(.A1(new_n1315), .A2(new_n1259), .ZN(new_n1316));
  AND3_X1   g1116(.A1(new_n1310), .A2(new_n1314), .A3(new_n1316), .ZN(new_n1317));
  AOI21_X1  g1117(.A(new_n1310), .B1(new_n1316), .B2(new_n1314), .ZN(new_n1318));
  NOR2_X1   g1118(.A1(new_n1317), .A2(new_n1318), .ZN(G402));
endmodule


