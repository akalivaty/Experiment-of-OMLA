

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n522, n523, n524, n525,
         n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536,
         n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547,
         n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558,
         n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569,
         n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580,
         n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591,
         n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602,
         n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, n613,
         n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624,
         n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635,
         n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, n646,
         n647, n648, n649, n650, n651, n652, n653, n654, n655, n656, n657,
         n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668,
         n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679,
         n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690,
         n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701,
         n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712,
         n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723,
         n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, n734,
         n735, n736, n737, n738, n739, n740, n741, n742, n743, n744, n745,
         n746, n747, n748, n749, n750, n751, n752, n753, n754, n755, n756,
         n757, n758, n759, n760, n761, n762, n763, n764, n765, n766, n767,
         n768, n769, n770, n771, n772, n773, n774, n775, n776, n777, n778,
         n779, n780, n781, n782, n783, n784, n785, n786, n787, n788, n789,
         n790, n791, n792, n793, n794, n795, n796, n797, n798, n799, n800,
         n801, n802, n803, n804, n805, n806, n807, n808, n809, n810, n811,
         n812, n813, n814, n815, n816, n817, n818, n819, n820, n821, n822,
         n823, n824, n825, n826, n827, n828, n829, n830, n831, n832, n833,
         n834, n835, n836, n837, n838, n839, n840, n841, n842, n843, n844,
         n845, n846, n847, n848, n849, n850, n851, n852, n853, n854, n855,
         n856, n857, n858, n859, n860, n861, n862, n863, n864, n865, n866,
         n867, n868, n869, n870, n871, n872, n873, n874, n875, n876, n877,
         n878, n879, n880, n881, n882, n883, n884, n885, n886, n887, n888,
         n889, n890, n891, n892, n893, n894, n895, n896, n897, n898, n899,
         n900, n901, n902, n903, n904, n905, n906, n907, n908, n909, n910,
         n911, n912, n913, n914, n915, n916, n917, n918, n919, n920, n921,
         n922, n923, n924, n925, n926, n927, n928, n929, n930, n931, n932,
         n933, n934, n935, n936, n937, n938, n939, n940, n941, n942, n943,
         n944, n945, n946, n947, n948, n949, n950, n951, n952, n953, n954,
         n955, n956, n957, n958, n959, n960, n961, n962, n963, n964, n965,
         n966, n967, n968, n969, n970, n971, n972, n973, n974, n975, n976,
         n977, n978, n979, n980, n981, n982, n983, n984, n985, n986, n987,
         n988, n989, n990, n991, n992, n993, n994, n995, n996, n997, n998,
         n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008,
         n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018,
         n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028,
         n1029, n1030;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  AND2_X1 U557 ( .A1(n822), .A2(n821), .ZN(n823) );
  NOR2_X1 U558 ( .A1(n726), .A2(n725), .ZN(n727) );
  INV_X1 U559 ( .A(n776), .ZN(n698) );
  XNOR2_X1 U560 ( .A(n745), .B(n744), .ZN(n751) );
  NOR2_X1 U561 ( .A1(n818), .A2(n817), .ZN(n522) );
  INV_X1 U562 ( .A(KEYINPUT27), .ZN(n715) );
  XNOR2_X1 U563 ( .A(n719), .B(KEYINPUT96), .ZN(n723) );
  INV_X1 U564 ( .A(KEYINPUT102), .ZN(n744) );
  INV_X1 U565 ( .A(n819), .ZN(n820) );
  NOR2_X1 U566 ( .A1(n522), .A2(n820), .ZN(n821) );
  OR2_X1 U567 ( .A1(n697), .A2(n696), .ZN(n776) );
  NOR2_X1 U568 ( .A1(G2104), .A2(n547), .ZN(n896) );
  NOR2_X1 U569 ( .A1(G651), .A2(G543), .ZN(n651) );
  NOR2_X1 U570 ( .A1(G651), .A2(n638), .ZN(n659) );
  XOR2_X1 U571 ( .A(KEYINPUT0), .B(G543), .Z(n638) );
  INV_X1 U572 ( .A(G651), .ZN(n523) );
  NOR2_X1 U573 ( .A1(n638), .A2(n523), .ZN(n655) );
  NAND2_X1 U574 ( .A1(G78), .A2(n655), .ZN(n527) );
  NOR2_X1 U575 ( .A1(G543), .A2(n523), .ZN(n524) );
  XOR2_X1 U576 ( .A(KEYINPUT66), .B(n524), .Z(n525) );
  XNOR2_X1 U577 ( .A(KEYINPUT1), .B(n525), .ZN(n652) );
  NAND2_X1 U578 ( .A1(G65), .A2(n652), .ZN(n526) );
  NAND2_X1 U579 ( .A1(n527), .A2(n526), .ZN(n531) );
  NAND2_X1 U580 ( .A1(G91), .A2(n651), .ZN(n529) );
  NAND2_X1 U581 ( .A1(G53), .A2(n659), .ZN(n528) );
  NAND2_X1 U582 ( .A1(n529), .A2(n528), .ZN(n530) );
  NOR2_X1 U583 ( .A1(n531), .A2(n530), .ZN(n532) );
  XOR2_X1 U584 ( .A(KEYINPUT68), .B(n532), .Z(G299) );
  NAND2_X1 U585 ( .A1(n659), .A2(G51), .ZN(n534) );
  NAND2_X1 U586 ( .A1(G63), .A2(n652), .ZN(n533) );
  NAND2_X1 U587 ( .A1(n534), .A2(n533), .ZN(n535) );
  XNOR2_X1 U588 ( .A(KEYINPUT6), .B(n535), .ZN(n542) );
  NAND2_X1 U589 ( .A1(n651), .A2(G89), .ZN(n536) );
  XNOR2_X1 U590 ( .A(n536), .B(KEYINPUT4), .ZN(n538) );
  NAND2_X1 U591 ( .A1(G76), .A2(n655), .ZN(n537) );
  NAND2_X1 U592 ( .A1(n538), .A2(n537), .ZN(n539) );
  XOR2_X1 U593 ( .A(KEYINPUT74), .B(n539), .Z(n540) );
  XNOR2_X1 U594 ( .A(KEYINPUT5), .B(n540), .ZN(n541) );
  NOR2_X1 U595 ( .A1(n542), .A2(n541), .ZN(n543) );
  XOR2_X1 U596 ( .A(KEYINPUT7), .B(n543), .Z(G168) );
  XOR2_X1 U597 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NOR2_X1 U598 ( .A1(G2105), .A2(G2104), .ZN(n544) );
  XOR2_X2 U599 ( .A(KEYINPUT17), .B(n544), .Z(n900) );
  NAND2_X1 U600 ( .A1(G138), .A2(n900), .ZN(n546) );
  INV_X1 U601 ( .A(G2105), .ZN(n547) );
  AND2_X1 U602 ( .A1(n547), .A2(G2104), .ZN(n619) );
  NAND2_X1 U603 ( .A1(G102), .A2(n619), .ZN(n545) );
  NAND2_X1 U604 ( .A1(n546), .A2(n545), .ZN(n551) );
  NAND2_X1 U605 ( .A1(G126), .A2(n896), .ZN(n549) );
  AND2_X1 U606 ( .A1(G2105), .A2(G2104), .ZN(n897) );
  NAND2_X1 U607 ( .A1(G114), .A2(n897), .ZN(n548) );
  NAND2_X1 U608 ( .A1(n549), .A2(n548), .ZN(n550) );
  NOR2_X1 U609 ( .A1(n551), .A2(n550), .ZN(G164) );
  XOR2_X1 U610 ( .A(G2443), .B(G2446), .Z(n553) );
  XNOR2_X1 U611 ( .A(G2427), .B(G2451), .ZN(n552) );
  XNOR2_X1 U612 ( .A(n553), .B(n552), .ZN(n559) );
  XOR2_X1 U613 ( .A(G2430), .B(G2454), .Z(n555) );
  XNOR2_X1 U614 ( .A(G1348), .B(G1341), .ZN(n554) );
  XNOR2_X1 U615 ( .A(n555), .B(n554), .ZN(n557) );
  XOR2_X1 U616 ( .A(G2435), .B(G2438), .Z(n556) );
  XNOR2_X1 U617 ( .A(n557), .B(n556), .ZN(n558) );
  XOR2_X1 U618 ( .A(n559), .B(n558), .Z(n560) );
  AND2_X1 U619 ( .A1(G14), .A2(n560), .ZN(G401) );
  XNOR2_X1 U620 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NAND2_X1 U621 ( .A1(n659), .A2(G52), .ZN(n562) );
  NAND2_X1 U622 ( .A1(G64), .A2(n652), .ZN(n561) );
  NAND2_X1 U623 ( .A1(n562), .A2(n561), .ZN(n567) );
  NAND2_X1 U624 ( .A1(G77), .A2(n655), .ZN(n564) );
  NAND2_X1 U625 ( .A1(G90), .A2(n651), .ZN(n563) );
  NAND2_X1 U626 ( .A1(n564), .A2(n563), .ZN(n565) );
  XOR2_X1 U627 ( .A(KEYINPUT9), .B(n565), .Z(n566) );
  NOR2_X1 U628 ( .A1(n567), .A2(n566), .ZN(n568) );
  XOR2_X1 U629 ( .A(KEYINPUT67), .B(n568), .Z(G171) );
  AND2_X1 U630 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U631 ( .A(G132), .ZN(G219) );
  INV_X1 U632 ( .A(G82), .ZN(G220) );
  INV_X1 U633 ( .A(G120), .ZN(G236) );
  NAND2_X1 U634 ( .A1(G75), .A2(n655), .ZN(n570) );
  NAND2_X1 U635 ( .A1(G88), .A2(n651), .ZN(n569) );
  NAND2_X1 U636 ( .A1(n570), .A2(n569), .ZN(n571) );
  XNOR2_X1 U637 ( .A(KEYINPUT83), .B(n571), .ZN(n576) );
  NAND2_X1 U638 ( .A1(n659), .A2(G50), .ZN(n573) );
  NAND2_X1 U639 ( .A1(G62), .A2(n652), .ZN(n572) );
  NAND2_X1 U640 ( .A1(n573), .A2(n572), .ZN(n574) );
  XOR2_X1 U641 ( .A(KEYINPUT82), .B(n574), .Z(n575) );
  NAND2_X1 U642 ( .A1(n576), .A2(n575), .ZN(G303) );
  NAND2_X1 U643 ( .A1(n896), .A2(G125), .ZN(n579) );
  NAND2_X1 U644 ( .A1(n619), .A2(G101), .ZN(n577) );
  XOR2_X1 U645 ( .A(n577), .B(KEYINPUT23), .Z(n578) );
  NAND2_X1 U646 ( .A1(n579), .A2(n578), .ZN(n580) );
  XNOR2_X1 U647 ( .A(n580), .B(KEYINPUT64), .ZN(n697) );
  NAND2_X1 U648 ( .A1(G137), .A2(n900), .ZN(n582) );
  NAND2_X1 U649 ( .A1(G113), .A2(n897), .ZN(n581) );
  NAND2_X1 U650 ( .A1(n582), .A2(n581), .ZN(n695) );
  NOR2_X1 U651 ( .A1(n697), .A2(n695), .ZN(G160) );
  NAND2_X1 U652 ( .A1(G7), .A2(G661), .ZN(n583) );
  XNOR2_X1 U653 ( .A(n583), .B(KEYINPUT70), .ZN(n584) );
  XOR2_X1 U654 ( .A(KEYINPUT10), .B(n584), .Z(n848) );
  NAND2_X1 U655 ( .A1(n848), .A2(G567), .ZN(n585) );
  XOR2_X1 U656 ( .A(KEYINPUT11), .B(n585), .Z(G234) );
  NAND2_X1 U657 ( .A1(G56), .A2(n652), .ZN(n586) );
  XOR2_X1 U658 ( .A(KEYINPUT14), .B(n586), .Z(n594) );
  NAND2_X1 U659 ( .A1(G68), .A2(n655), .ZN(n590) );
  XOR2_X1 U660 ( .A(KEYINPUT12), .B(KEYINPUT71), .Z(n588) );
  NAND2_X1 U661 ( .A1(G81), .A2(n651), .ZN(n587) );
  XNOR2_X1 U662 ( .A(n588), .B(n587), .ZN(n589) );
  NAND2_X1 U663 ( .A1(n590), .A2(n589), .ZN(n591) );
  XNOR2_X1 U664 ( .A(n591), .B(KEYINPUT13), .ZN(n592) );
  XOR2_X1 U665 ( .A(KEYINPUT72), .B(n592), .Z(n593) );
  NOR2_X1 U666 ( .A1(n594), .A2(n593), .ZN(n596) );
  NAND2_X1 U667 ( .A1(n659), .A2(G43), .ZN(n595) );
  NAND2_X1 U668 ( .A1(n596), .A2(n595), .ZN(n973) );
  INV_X1 U669 ( .A(G860), .ZN(n610) );
  OR2_X1 U670 ( .A1(n973), .A2(n610), .ZN(G153) );
  XNOR2_X1 U671 ( .A(G171), .B(KEYINPUT73), .ZN(G301) );
  NAND2_X1 U672 ( .A1(G868), .A2(G301), .ZN(n605) );
  NAND2_X1 U673 ( .A1(G79), .A2(n655), .ZN(n598) );
  NAND2_X1 U674 ( .A1(G66), .A2(n652), .ZN(n597) );
  NAND2_X1 U675 ( .A1(n598), .A2(n597), .ZN(n602) );
  NAND2_X1 U676 ( .A1(G92), .A2(n651), .ZN(n600) );
  NAND2_X1 U677 ( .A1(G54), .A2(n659), .ZN(n599) );
  NAND2_X1 U678 ( .A1(n600), .A2(n599), .ZN(n601) );
  NOR2_X1 U679 ( .A1(n602), .A2(n601), .ZN(n603) );
  XOR2_X1 U680 ( .A(KEYINPUT15), .B(n603), .Z(n972) );
  OR2_X1 U681 ( .A1(n972), .A2(G868), .ZN(n604) );
  NAND2_X1 U682 ( .A1(n605), .A2(n604), .ZN(G284) );
  INV_X1 U683 ( .A(G868), .ZN(n674) );
  XOR2_X1 U684 ( .A(KEYINPUT75), .B(n674), .Z(n606) );
  NOR2_X1 U685 ( .A1(G286), .A2(n606), .ZN(n608) );
  NOR2_X1 U686 ( .A1(G299), .A2(G868), .ZN(n607) );
  NOR2_X1 U687 ( .A1(n608), .A2(n607), .ZN(n609) );
  XNOR2_X1 U688 ( .A(KEYINPUT76), .B(n609), .ZN(G297) );
  NAND2_X1 U689 ( .A1(n610), .A2(G559), .ZN(n611) );
  NAND2_X1 U690 ( .A1(n611), .A2(n972), .ZN(n612) );
  XNOR2_X1 U691 ( .A(n612), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U692 ( .A1(G559), .A2(n674), .ZN(n613) );
  NAND2_X1 U693 ( .A1(n972), .A2(n613), .ZN(n614) );
  XNOR2_X1 U694 ( .A(n614), .B(KEYINPUT77), .ZN(n616) );
  NOR2_X1 U695 ( .A1(n973), .A2(G868), .ZN(n615) );
  NOR2_X1 U696 ( .A1(n616), .A2(n615), .ZN(G282) );
  NAND2_X1 U697 ( .A1(G123), .A2(n896), .ZN(n617) );
  XNOR2_X1 U698 ( .A(n617), .B(KEYINPUT18), .ZN(n618) );
  XNOR2_X1 U699 ( .A(n618), .B(KEYINPUT78), .ZN(n621) );
  NAND2_X1 U700 ( .A1(G99), .A2(n619), .ZN(n620) );
  NAND2_X1 U701 ( .A1(n621), .A2(n620), .ZN(n625) );
  NAND2_X1 U702 ( .A1(G135), .A2(n900), .ZN(n623) );
  NAND2_X1 U703 ( .A1(G111), .A2(n897), .ZN(n622) );
  NAND2_X1 U704 ( .A1(n623), .A2(n622), .ZN(n624) );
  NOR2_X1 U705 ( .A1(n625), .A2(n624), .ZN(n922) );
  XNOR2_X1 U706 ( .A(n922), .B(G2096), .ZN(n626) );
  INV_X1 U707 ( .A(G2100), .ZN(n852) );
  NAND2_X1 U708 ( .A1(n626), .A2(n852), .ZN(G156) );
  NAND2_X1 U709 ( .A1(n659), .A2(G55), .ZN(n628) );
  NAND2_X1 U710 ( .A1(G67), .A2(n652), .ZN(n627) );
  NAND2_X1 U711 ( .A1(n628), .A2(n627), .ZN(n633) );
  NAND2_X1 U712 ( .A1(G80), .A2(n655), .ZN(n630) );
  NAND2_X1 U713 ( .A1(G93), .A2(n651), .ZN(n629) );
  NAND2_X1 U714 ( .A1(n630), .A2(n629), .ZN(n631) );
  XOR2_X1 U715 ( .A(KEYINPUT81), .B(n631), .Z(n632) );
  OR2_X1 U716 ( .A1(n633), .A2(n632), .ZN(n673) );
  NAND2_X1 U717 ( .A1(G559), .A2(n972), .ZN(n634) );
  XNOR2_X1 U718 ( .A(n634), .B(KEYINPUT79), .ZN(n670) );
  XOR2_X1 U719 ( .A(n670), .B(KEYINPUT80), .Z(n635) );
  XNOR2_X1 U720 ( .A(n973), .B(n635), .ZN(n636) );
  NOR2_X1 U721 ( .A1(G860), .A2(n636), .ZN(n637) );
  XOR2_X1 U722 ( .A(n673), .B(n637), .Z(G145) );
  NAND2_X1 U723 ( .A1(G87), .A2(n638), .ZN(n640) );
  NAND2_X1 U724 ( .A1(G74), .A2(G651), .ZN(n639) );
  NAND2_X1 U725 ( .A1(n640), .A2(n639), .ZN(n641) );
  NOR2_X1 U726 ( .A1(n652), .A2(n641), .ZN(n643) );
  NAND2_X1 U727 ( .A1(n659), .A2(G49), .ZN(n642) );
  NAND2_X1 U728 ( .A1(n643), .A2(n642), .ZN(G288) );
  NAND2_X1 U729 ( .A1(n659), .A2(G47), .ZN(n645) );
  NAND2_X1 U730 ( .A1(G60), .A2(n652), .ZN(n644) );
  NAND2_X1 U731 ( .A1(n645), .A2(n644), .ZN(n648) );
  NAND2_X1 U732 ( .A1(G72), .A2(n655), .ZN(n646) );
  XNOR2_X1 U733 ( .A(KEYINPUT65), .B(n646), .ZN(n647) );
  NOR2_X1 U734 ( .A1(n648), .A2(n647), .ZN(n650) );
  NAND2_X1 U735 ( .A1(n651), .A2(G85), .ZN(n649) );
  NAND2_X1 U736 ( .A1(n650), .A2(n649), .ZN(G290) );
  NAND2_X1 U737 ( .A1(n651), .A2(G86), .ZN(n654) );
  NAND2_X1 U738 ( .A1(G61), .A2(n652), .ZN(n653) );
  NAND2_X1 U739 ( .A1(n654), .A2(n653), .ZN(n658) );
  NAND2_X1 U740 ( .A1(n655), .A2(G73), .ZN(n656) );
  XOR2_X1 U741 ( .A(KEYINPUT2), .B(n656), .Z(n657) );
  NOR2_X1 U742 ( .A1(n658), .A2(n657), .ZN(n661) );
  NAND2_X1 U743 ( .A1(n659), .A2(G48), .ZN(n660) );
  NAND2_X1 U744 ( .A1(n661), .A2(n660), .ZN(G305) );
  XOR2_X1 U745 ( .A(KEYINPUT85), .B(KEYINPUT84), .Z(n663) );
  XOR2_X1 U746 ( .A(n673), .B(KEYINPUT19), .Z(n662) );
  XNOR2_X1 U747 ( .A(n663), .B(n662), .ZN(n664) );
  XNOR2_X1 U748 ( .A(n664), .B(G288), .ZN(n667) );
  XOR2_X1 U749 ( .A(G299), .B(G303), .Z(n665) );
  XNOR2_X1 U750 ( .A(n665), .B(n973), .ZN(n666) );
  XNOR2_X1 U751 ( .A(n667), .B(n666), .ZN(n668) );
  XNOR2_X1 U752 ( .A(n668), .B(G290), .ZN(n669) );
  XNOR2_X1 U753 ( .A(n669), .B(G305), .ZN(n910) );
  XNOR2_X1 U754 ( .A(n910), .B(n670), .ZN(n671) );
  NAND2_X1 U755 ( .A1(n671), .A2(G868), .ZN(n672) );
  XNOR2_X1 U756 ( .A(n672), .B(KEYINPUT86), .ZN(n676) );
  NAND2_X1 U757 ( .A1(n674), .A2(n673), .ZN(n675) );
  NAND2_X1 U758 ( .A1(n676), .A2(n675), .ZN(G295) );
  NAND2_X1 U759 ( .A1(G2084), .A2(G2078), .ZN(n677) );
  XOR2_X1 U760 ( .A(KEYINPUT20), .B(n677), .Z(n678) );
  NAND2_X1 U761 ( .A1(G2090), .A2(n678), .ZN(n679) );
  XNOR2_X1 U762 ( .A(KEYINPUT21), .B(n679), .ZN(n680) );
  NAND2_X1 U763 ( .A1(n680), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U764 ( .A(KEYINPUT69), .B(G57), .ZN(G237) );
  NOR2_X1 U765 ( .A1(G237), .A2(G236), .ZN(n681) );
  NAND2_X1 U766 ( .A1(G69), .A2(n681), .ZN(n682) );
  XNOR2_X1 U767 ( .A(KEYINPUT87), .B(n682), .ZN(n683) );
  NAND2_X1 U768 ( .A1(n683), .A2(G108), .ZN(n684) );
  XNOR2_X1 U769 ( .A(KEYINPUT88), .B(n684), .ZN(n919) );
  NAND2_X1 U770 ( .A1(n919), .A2(G567), .ZN(n685) );
  XNOR2_X1 U771 ( .A(n685), .B(KEYINPUT89), .ZN(n690) );
  NOR2_X1 U772 ( .A1(G220), .A2(G219), .ZN(n686) );
  XNOR2_X1 U773 ( .A(KEYINPUT22), .B(n686), .ZN(n687) );
  NAND2_X1 U774 ( .A1(n687), .A2(G96), .ZN(n688) );
  OR2_X1 U775 ( .A1(G218), .A2(n688), .ZN(n920) );
  AND2_X1 U776 ( .A1(G2106), .A2(n920), .ZN(n689) );
  NOR2_X1 U777 ( .A1(n690), .A2(n689), .ZN(G319) );
  NAND2_X1 U778 ( .A1(G483), .A2(G661), .ZN(n692) );
  INV_X1 U779 ( .A(G319), .ZN(n691) );
  NOR2_X1 U780 ( .A1(n692), .A2(n691), .ZN(n693) );
  XNOR2_X1 U781 ( .A(n693), .B(KEYINPUT90), .ZN(n851) );
  NAND2_X1 U782 ( .A1(G36), .A2(n851), .ZN(G176) );
  NOR2_X1 U783 ( .A1(G164), .A2(G1384), .ZN(n777) );
  INV_X1 U784 ( .A(G40), .ZN(n694) );
  OR2_X1 U785 ( .A1(n695), .A2(n694), .ZN(n696) );
  NAND2_X2 U786 ( .A1(n777), .A2(n698), .ZN(n752) );
  NOR2_X1 U787 ( .A1(n752), .A2(G2084), .ZN(n699) );
  XNOR2_X1 U788 ( .A(n699), .B(KEYINPUT94), .ZN(n733) );
  NAND2_X1 U789 ( .A1(n733), .A2(G8), .ZN(n749) );
  NAND2_X1 U790 ( .A1(G8), .A2(n752), .ZN(n817) );
  NOR2_X1 U791 ( .A1(G1966), .A2(n817), .ZN(n746) );
  XOR2_X1 U792 ( .A(KEYINPUT95), .B(n752), .Z(n714) );
  INV_X1 U793 ( .A(n714), .ZN(n728) );
  NAND2_X1 U794 ( .A1(G2067), .A2(n728), .ZN(n700) );
  XNOR2_X1 U795 ( .A(KEYINPUT98), .B(n700), .ZN(n703) );
  NAND2_X1 U796 ( .A1(G1348), .A2(n752), .ZN(n701) );
  XOR2_X1 U797 ( .A(KEYINPUT97), .B(n701), .Z(n702) );
  NAND2_X1 U798 ( .A1(n703), .A2(n702), .ZN(n709) );
  INV_X1 U799 ( .A(G1996), .ZN(n952) );
  NOR2_X1 U800 ( .A1(n752), .A2(n952), .ZN(n704) );
  XOR2_X1 U801 ( .A(KEYINPUT26), .B(n704), .Z(n706) );
  NAND2_X1 U802 ( .A1(n752), .A2(G1341), .ZN(n705) );
  NAND2_X1 U803 ( .A1(n706), .A2(n705), .ZN(n707) );
  NOR2_X1 U804 ( .A1(n973), .A2(n707), .ZN(n711) );
  NAND2_X1 U805 ( .A1(n972), .A2(n711), .ZN(n708) );
  NAND2_X1 U806 ( .A1(n709), .A2(n708), .ZN(n710) );
  XOR2_X1 U807 ( .A(n710), .B(KEYINPUT99), .Z(n713) );
  OR2_X1 U808 ( .A1(n972), .A2(n711), .ZN(n712) );
  AND2_X1 U809 ( .A1(n713), .A2(n712), .ZN(n721) );
  NAND2_X1 U810 ( .A1(n714), .A2(G1956), .ZN(n718) );
  NAND2_X1 U811 ( .A1(n728), .A2(G2072), .ZN(n716) );
  XNOR2_X1 U812 ( .A(n716), .B(n715), .ZN(n717) );
  NAND2_X1 U813 ( .A1(n718), .A2(n717), .ZN(n719) );
  NOR2_X1 U814 ( .A1(n723), .A2(G299), .ZN(n720) );
  NOR2_X1 U815 ( .A1(n721), .A2(n720), .ZN(n722) );
  XNOR2_X1 U816 ( .A(n722), .B(KEYINPUT100), .ZN(n726) );
  NAND2_X1 U817 ( .A1(G299), .A2(n723), .ZN(n724) );
  XOR2_X1 U818 ( .A(KEYINPUT28), .B(n724), .Z(n725) );
  XNOR2_X1 U819 ( .A(n727), .B(KEYINPUT29), .ZN(n732) );
  INV_X1 U820 ( .A(G1961), .ZN(n1018) );
  NAND2_X1 U821 ( .A1(n1018), .A2(n752), .ZN(n730) );
  XNOR2_X1 U822 ( .A(G2078), .B(KEYINPUT25), .ZN(n960) );
  NAND2_X1 U823 ( .A1(n728), .A2(n960), .ZN(n729) );
  NAND2_X1 U824 ( .A1(n730), .A2(n729), .ZN(n738) );
  NAND2_X1 U825 ( .A1(G171), .A2(n738), .ZN(n731) );
  NAND2_X1 U826 ( .A1(n732), .A2(n731), .ZN(n743) );
  NOR2_X1 U827 ( .A1(n746), .A2(n733), .ZN(n734) );
  NAND2_X1 U828 ( .A1(n734), .A2(G8), .ZN(n735) );
  XOR2_X1 U829 ( .A(KEYINPUT30), .B(n735), .Z(n736) );
  XNOR2_X1 U830 ( .A(KEYINPUT101), .B(n736), .ZN(n737) );
  NOR2_X1 U831 ( .A1(G168), .A2(n737), .ZN(n740) );
  NOR2_X1 U832 ( .A1(G171), .A2(n738), .ZN(n739) );
  NOR2_X1 U833 ( .A1(n740), .A2(n739), .ZN(n741) );
  XOR2_X1 U834 ( .A(KEYINPUT31), .B(n741), .Z(n742) );
  NAND2_X1 U835 ( .A1(n743), .A2(n742), .ZN(n745) );
  NOR2_X1 U836 ( .A1(n746), .A2(n751), .ZN(n747) );
  XOR2_X1 U837 ( .A(KEYINPUT103), .B(n747), .Z(n748) );
  NAND2_X1 U838 ( .A1(n749), .A2(n748), .ZN(n761) );
  INV_X1 U839 ( .A(G286), .ZN(n750) );
  OR2_X1 U840 ( .A1(n751), .A2(n750), .ZN(n757) );
  NOR2_X1 U841 ( .A1(G1971), .A2(n817), .ZN(n754) );
  NOR2_X1 U842 ( .A1(G2090), .A2(n752), .ZN(n753) );
  NOR2_X1 U843 ( .A1(n754), .A2(n753), .ZN(n755) );
  NAND2_X1 U844 ( .A1(n755), .A2(G303), .ZN(n756) );
  NAND2_X1 U845 ( .A1(n757), .A2(n756), .ZN(n758) );
  NAND2_X1 U846 ( .A1(n758), .A2(G8), .ZN(n759) );
  XNOR2_X1 U847 ( .A(n759), .B(KEYINPUT32), .ZN(n760) );
  NAND2_X1 U848 ( .A1(n761), .A2(n760), .ZN(n816) );
  NOR2_X1 U849 ( .A1(G1971), .A2(G303), .ZN(n763) );
  NOR2_X1 U850 ( .A1(G288), .A2(G1976), .ZN(n762) );
  XNOR2_X1 U851 ( .A(n762), .B(KEYINPUT104), .ZN(n976) );
  NOR2_X1 U852 ( .A1(n763), .A2(n976), .ZN(n765) );
  INV_X1 U853 ( .A(KEYINPUT33), .ZN(n764) );
  AND2_X1 U854 ( .A1(n765), .A2(n764), .ZN(n766) );
  NAND2_X1 U855 ( .A1(n816), .A2(n766), .ZN(n770) );
  INV_X1 U856 ( .A(n817), .ZN(n767) );
  NAND2_X1 U857 ( .A1(G1976), .A2(G288), .ZN(n977) );
  AND2_X1 U858 ( .A1(n767), .A2(n977), .ZN(n768) );
  OR2_X1 U859 ( .A1(KEYINPUT33), .A2(n768), .ZN(n769) );
  AND2_X1 U860 ( .A1(n770), .A2(n769), .ZN(n809) );
  NAND2_X1 U861 ( .A1(KEYINPUT33), .A2(n976), .ZN(n771) );
  XOR2_X1 U862 ( .A(KEYINPUT105), .B(n771), .Z(n772) );
  NOR2_X1 U863 ( .A1(n817), .A2(n772), .ZN(n773) );
  XNOR2_X1 U864 ( .A(n773), .B(KEYINPUT106), .ZN(n775) );
  XOR2_X1 U865 ( .A(G1981), .B(G305), .Z(n991) );
  INV_X1 U866 ( .A(n991), .ZN(n774) );
  NOR2_X1 U867 ( .A1(n775), .A2(n774), .ZN(n805) );
  NOR2_X1 U868 ( .A1(n777), .A2(n776), .ZN(n841) );
  XNOR2_X1 U869 ( .A(KEYINPUT34), .B(KEYINPUT92), .ZN(n781) );
  NAND2_X1 U870 ( .A1(G140), .A2(n900), .ZN(n779) );
  NAND2_X1 U871 ( .A1(G104), .A2(n619), .ZN(n778) );
  NAND2_X1 U872 ( .A1(n779), .A2(n778), .ZN(n780) );
  XNOR2_X1 U873 ( .A(n781), .B(n780), .ZN(n787) );
  XNOR2_X1 U874 ( .A(KEYINPUT35), .B(KEYINPUT93), .ZN(n785) );
  NAND2_X1 U875 ( .A1(G128), .A2(n896), .ZN(n783) );
  NAND2_X1 U876 ( .A1(G116), .A2(n897), .ZN(n782) );
  NAND2_X1 U877 ( .A1(n783), .A2(n782), .ZN(n784) );
  XNOR2_X1 U878 ( .A(n785), .B(n784), .ZN(n786) );
  NOR2_X1 U879 ( .A1(n787), .A2(n786), .ZN(n788) );
  XOR2_X1 U880 ( .A(n788), .B(KEYINPUT36), .Z(n885) );
  XOR2_X1 U881 ( .A(KEYINPUT37), .B(G2067), .Z(n838) );
  AND2_X1 U882 ( .A1(n885), .A2(n838), .ZN(n927) );
  NAND2_X1 U883 ( .A1(n841), .A2(n927), .ZN(n836) );
  NAND2_X1 U884 ( .A1(G131), .A2(n900), .ZN(n790) );
  NAND2_X1 U885 ( .A1(G95), .A2(n619), .ZN(n789) );
  NAND2_X1 U886 ( .A1(n790), .A2(n789), .ZN(n794) );
  NAND2_X1 U887 ( .A1(G119), .A2(n896), .ZN(n792) );
  NAND2_X1 U888 ( .A1(G107), .A2(n897), .ZN(n791) );
  NAND2_X1 U889 ( .A1(n792), .A2(n791), .ZN(n793) );
  NOR2_X1 U890 ( .A1(n794), .A2(n793), .ZN(n888) );
  INV_X1 U891 ( .A(G1991), .ZN(n829) );
  NOR2_X1 U892 ( .A1(n888), .A2(n829), .ZN(n803) );
  NAND2_X1 U893 ( .A1(G141), .A2(n900), .ZN(n796) );
  NAND2_X1 U894 ( .A1(G129), .A2(n896), .ZN(n795) );
  NAND2_X1 U895 ( .A1(n796), .A2(n795), .ZN(n799) );
  NAND2_X1 U896 ( .A1(n619), .A2(G105), .ZN(n797) );
  XOR2_X1 U897 ( .A(KEYINPUT38), .B(n797), .Z(n798) );
  NOR2_X1 U898 ( .A1(n799), .A2(n798), .ZN(n801) );
  NAND2_X1 U899 ( .A1(n897), .A2(G117), .ZN(n800) );
  NAND2_X1 U900 ( .A1(n801), .A2(n800), .ZN(n893) );
  AND2_X1 U901 ( .A1(G1996), .A2(n893), .ZN(n802) );
  NOR2_X1 U902 ( .A1(n803), .A2(n802), .ZN(n925) );
  INV_X1 U903 ( .A(n925), .ZN(n804) );
  NAND2_X1 U904 ( .A1(n804), .A2(n841), .ZN(n828) );
  AND2_X1 U905 ( .A1(n836), .A2(n828), .ZN(n819) );
  AND2_X1 U906 ( .A1(n805), .A2(n819), .ZN(n807) );
  XOR2_X1 U907 ( .A(G1986), .B(KEYINPUT91), .Z(n806) );
  XNOR2_X1 U908 ( .A(G290), .B(n806), .ZN(n985) );
  NAND2_X1 U909 ( .A1(n985), .A2(n841), .ZN(n824) );
  AND2_X1 U910 ( .A1(n807), .A2(n824), .ZN(n808) );
  NAND2_X1 U911 ( .A1(n809), .A2(n808), .ZN(n826) );
  NOR2_X1 U912 ( .A1(G2090), .A2(G303), .ZN(n810) );
  NAND2_X1 U913 ( .A1(G8), .A2(n810), .ZN(n814) );
  NOR2_X1 U914 ( .A1(G1981), .A2(G305), .ZN(n811) );
  XOR2_X1 U915 ( .A(n811), .B(KEYINPUT24), .Z(n812) );
  NOR2_X1 U916 ( .A1(n817), .A2(n812), .ZN(n818) );
  INV_X1 U917 ( .A(n818), .ZN(n813) );
  AND2_X1 U918 ( .A1(n814), .A2(n813), .ZN(n815) );
  NAND2_X1 U919 ( .A1(n816), .A2(n815), .ZN(n822) );
  NAND2_X1 U920 ( .A1(n824), .A2(n823), .ZN(n825) );
  AND2_X1 U921 ( .A1(n826), .A2(n825), .ZN(n844) );
  NOR2_X1 U922 ( .A1(G1996), .A2(n893), .ZN(n827) );
  XOR2_X1 U923 ( .A(KEYINPUT107), .B(n827), .Z(n936) );
  INV_X1 U924 ( .A(n828), .ZN(n832) );
  AND2_X1 U925 ( .A1(n829), .A2(n888), .ZN(n921) );
  NOR2_X1 U926 ( .A1(G1986), .A2(G290), .ZN(n830) );
  NOR2_X1 U927 ( .A1(n921), .A2(n830), .ZN(n831) );
  NOR2_X1 U928 ( .A1(n832), .A2(n831), .ZN(n833) );
  XNOR2_X1 U929 ( .A(n833), .B(KEYINPUT108), .ZN(n834) );
  NOR2_X1 U930 ( .A1(n936), .A2(n834), .ZN(n835) );
  XNOR2_X1 U931 ( .A(n835), .B(KEYINPUT39), .ZN(n837) );
  NAND2_X1 U932 ( .A1(n837), .A2(n836), .ZN(n840) );
  NOR2_X1 U933 ( .A1(n838), .A2(n885), .ZN(n839) );
  XNOR2_X1 U934 ( .A(n839), .B(KEYINPUT109), .ZN(n940) );
  NAND2_X1 U935 ( .A1(n840), .A2(n940), .ZN(n842) );
  NAND2_X1 U936 ( .A1(n842), .A2(n841), .ZN(n843) );
  NAND2_X1 U937 ( .A1(n844), .A2(n843), .ZN(n847) );
  XOR2_X1 U938 ( .A(KEYINPUT111), .B(KEYINPUT40), .Z(n845) );
  XNOR2_X1 U939 ( .A(KEYINPUT110), .B(n845), .ZN(n846) );
  XNOR2_X1 U940 ( .A(n847), .B(n846), .ZN(G329) );
  NAND2_X1 U941 ( .A1(G2106), .A2(n848), .ZN(G217) );
  INV_X1 U942 ( .A(n848), .ZN(G223) );
  AND2_X1 U943 ( .A1(G15), .A2(G2), .ZN(n849) );
  NAND2_X1 U944 ( .A1(G661), .A2(n849), .ZN(G259) );
  NAND2_X1 U945 ( .A1(G3), .A2(G1), .ZN(n850) );
  NAND2_X1 U946 ( .A1(n851), .A2(n850), .ZN(G188) );
  XNOR2_X1 U947 ( .A(n852), .B(G2096), .ZN(n854) );
  XNOR2_X1 U948 ( .A(KEYINPUT42), .B(G2678), .ZN(n853) );
  XNOR2_X1 U949 ( .A(n854), .B(n853), .ZN(n858) );
  XOR2_X1 U950 ( .A(KEYINPUT43), .B(G2090), .Z(n856) );
  XNOR2_X1 U951 ( .A(G2067), .B(G2072), .ZN(n855) );
  XNOR2_X1 U952 ( .A(n856), .B(n855), .ZN(n857) );
  XOR2_X1 U953 ( .A(n858), .B(n857), .Z(n860) );
  XNOR2_X1 U954 ( .A(G2084), .B(G2078), .ZN(n859) );
  XNOR2_X1 U955 ( .A(n860), .B(n859), .ZN(G227) );
  XOR2_X1 U956 ( .A(G1976), .B(G1971), .Z(n862) );
  XNOR2_X1 U957 ( .A(G1986), .B(G1956), .ZN(n861) );
  XNOR2_X1 U958 ( .A(n862), .B(n861), .ZN(n863) );
  XOR2_X1 U959 ( .A(n863), .B(G2474), .Z(n865) );
  XOR2_X1 U960 ( .A(n952), .B(G1991), .Z(n864) );
  XNOR2_X1 U961 ( .A(n865), .B(n864), .ZN(n869) );
  XOR2_X1 U962 ( .A(KEYINPUT41), .B(G1981), .Z(n867) );
  XOR2_X1 U963 ( .A(G1966), .B(n1018), .Z(n866) );
  XNOR2_X1 U964 ( .A(n867), .B(n866), .ZN(n868) );
  XNOR2_X1 U965 ( .A(n869), .B(n868), .ZN(G229) );
  NAND2_X1 U966 ( .A1(G124), .A2(n896), .ZN(n870) );
  XNOR2_X1 U967 ( .A(n870), .B(KEYINPUT44), .ZN(n872) );
  NAND2_X1 U968 ( .A1(n619), .A2(G100), .ZN(n871) );
  NAND2_X1 U969 ( .A1(n872), .A2(n871), .ZN(n876) );
  NAND2_X1 U970 ( .A1(G136), .A2(n900), .ZN(n874) );
  NAND2_X1 U971 ( .A1(G112), .A2(n897), .ZN(n873) );
  NAND2_X1 U972 ( .A1(n874), .A2(n873), .ZN(n875) );
  NOR2_X1 U973 ( .A1(n876), .A2(n875), .ZN(G162) );
  NAND2_X1 U974 ( .A1(G139), .A2(n900), .ZN(n878) );
  NAND2_X1 U975 ( .A1(G103), .A2(n619), .ZN(n877) );
  NAND2_X1 U976 ( .A1(n878), .A2(n877), .ZN(n879) );
  XNOR2_X1 U977 ( .A(KEYINPUT112), .B(n879), .ZN(n884) );
  NAND2_X1 U978 ( .A1(G127), .A2(n896), .ZN(n881) );
  NAND2_X1 U979 ( .A1(G115), .A2(n897), .ZN(n880) );
  NAND2_X1 U980 ( .A1(n881), .A2(n880), .ZN(n882) );
  XOR2_X1 U981 ( .A(KEYINPUT47), .B(n882), .Z(n883) );
  NOR2_X1 U982 ( .A1(n884), .A2(n883), .ZN(n931) );
  XOR2_X1 U983 ( .A(G162), .B(n931), .Z(n887) );
  XNOR2_X1 U984 ( .A(n885), .B(n922), .ZN(n886) );
  XNOR2_X1 U985 ( .A(n887), .B(n886), .ZN(n892) );
  XOR2_X1 U986 ( .A(KEYINPUT48), .B(KEYINPUT113), .Z(n890) );
  XNOR2_X1 U987 ( .A(n888), .B(KEYINPUT46), .ZN(n889) );
  XNOR2_X1 U988 ( .A(n890), .B(n889), .ZN(n891) );
  XOR2_X1 U989 ( .A(n892), .B(n891), .Z(n895) );
  XOR2_X1 U990 ( .A(G164), .B(n893), .Z(n894) );
  XNOR2_X1 U991 ( .A(n895), .B(n894), .ZN(n908) );
  NAND2_X1 U992 ( .A1(G130), .A2(n896), .ZN(n899) );
  NAND2_X1 U993 ( .A1(G118), .A2(n897), .ZN(n898) );
  NAND2_X1 U994 ( .A1(n899), .A2(n898), .ZN(n905) );
  NAND2_X1 U995 ( .A1(G142), .A2(n900), .ZN(n902) );
  NAND2_X1 U996 ( .A1(G106), .A2(n619), .ZN(n901) );
  NAND2_X1 U997 ( .A1(n902), .A2(n901), .ZN(n903) );
  XOR2_X1 U998 ( .A(KEYINPUT45), .B(n903), .Z(n904) );
  NOR2_X1 U999 ( .A1(n905), .A2(n904), .ZN(n906) );
  XOR2_X1 U1000 ( .A(G160), .B(n906), .Z(n907) );
  XNOR2_X1 U1001 ( .A(n908), .B(n907), .ZN(n909) );
  NOR2_X1 U1002 ( .A1(G37), .A2(n909), .ZN(G395) );
  XNOR2_X1 U1003 ( .A(n972), .B(G286), .ZN(n911) );
  XNOR2_X1 U1004 ( .A(n911), .B(n910), .ZN(n912) );
  XNOR2_X1 U1005 ( .A(n912), .B(G171), .ZN(n913) );
  NOR2_X1 U1006 ( .A1(G37), .A2(n913), .ZN(G397) );
  NOR2_X1 U1007 ( .A1(G227), .A2(G229), .ZN(n914) );
  XNOR2_X1 U1008 ( .A(KEYINPUT49), .B(n914), .ZN(n915) );
  NOR2_X1 U1009 ( .A1(G401), .A2(n915), .ZN(n916) );
  AND2_X1 U1010 ( .A1(G319), .A2(n916), .ZN(n918) );
  NOR2_X1 U1011 ( .A1(G395), .A2(G397), .ZN(n917) );
  NAND2_X1 U1012 ( .A1(n918), .A2(n917), .ZN(G225) );
  XOR2_X1 U1013 ( .A(KEYINPUT114), .B(G225), .Z(G308) );
  INV_X1 U1015 ( .A(G108), .ZN(G238) );
  INV_X1 U1016 ( .A(G96), .ZN(G221) );
  NOR2_X1 U1017 ( .A1(n920), .A2(n919), .ZN(G325) );
  INV_X1 U1018 ( .A(G325), .ZN(G261) );
  INV_X1 U1019 ( .A(G303), .ZN(G166) );
  INV_X1 U1020 ( .A(G69), .ZN(G235) );
  XNOR2_X1 U1021 ( .A(G160), .B(G2084), .ZN(n929) );
  NOR2_X1 U1022 ( .A1(n922), .A2(n921), .ZN(n923) );
  XOR2_X1 U1023 ( .A(KEYINPUT115), .B(n923), .Z(n924) );
  NAND2_X1 U1024 ( .A1(n925), .A2(n924), .ZN(n926) );
  NOR2_X1 U1025 ( .A1(n927), .A2(n926), .ZN(n928) );
  NAND2_X1 U1026 ( .A1(n929), .A2(n928), .ZN(n930) );
  XNOR2_X1 U1027 ( .A(n930), .B(KEYINPUT116), .ZN(n943) );
  XOR2_X1 U1028 ( .A(G2072), .B(n931), .Z(n933) );
  XOR2_X1 U1029 ( .A(G164), .B(G2078), .Z(n932) );
  NOR2_X1 U1030 ( .A1(n933), .A2(n932), .ZN(n934) );
  XOR2_X1 U1031 ( .A(KEYINPUT50), .B(n934), .Z(n939) );
  XOR2_X1 U1032 ( .A(G2090), .B(G162), .Z(n935) );
  NOR2_X1 U1033 ( .A1(n936), .A2(n935), .ZN(n937) );
  XNOR2_X1 U1034 ( .A(KEYINPUT51), .B(n937), .ZN(n938) );
  NOR2_X1 U1035 ( .A1(n939), .A2(n938), .ZN(n941) );
  NAND2_X1 U1036 ( .A1(n941), .A2(n940), .ZN(n942) );
  NOR2_X1 U1037 ( .A1(n943), .A2(n942), .ZN(n944) );
  XNOR2_X1 U1038 ( .A(KEYINPUT52), .B(n944), .ZN(n945) );
  INV_X1 U1039 ( .A(KEYINPUT55), .ZN(n967) );
  NAND2_X1 U1040 ( .A1(n945), .A2(n967), .ZN(n946) );
  NAND2_X1 U1041 ( .A1(n946), .A2(G29), .ZN(n1029) );
  XOR2_X1 U1042 ( .A(G29), .B(KEYINPUT120), .Z(n970) );
  XNOR2_X1 U1043 ( .A(KEYINPUT54), .B(KEYINPUT119), .ZN(n947) );
  XNOR2_X1 U1044 ( .A(n947), .B(G34), .ZN(n948) );
  XNOR2_X1 U1045 ( .A(G2084), .B(n948), .ZN(n951) );
  XNOR2_X1 U1046 ( .A(G2090), .B(KEYINPUT117), .ZN(n949) );
  XNOR2_X1 U1047 ( .A(n949), .B(G35), .ZN(n950) );
  NAND2_X1 U1048 ( .A1(n951), .A2(n950), .ZN(n966) );
  XOR2_X1 U1049 ( .A(n952), .B(G32), .Z(n954) );
  XNOR2_X1 U1050 ( .A(G33), .B(G2072), .ZN(n953) );
  NOR2_X1 U1051 ( .A1(n954), .A2(n953), .ZN(n959) );
  XOR2_X1 U1052 ( .A(G25), .B(G1991), .Z(n955) );
  NAND2_X1 U1053 ( .A1(n955), .A2(G28), .ZN(n957) );
  XNOR2_X1 U1054 ( .A(G26), .B(G2067), .ZN(n956) );
  NOR2_X1 U1055 ( .A1(n957), .A2(n956), .ZN(n958) );
  NAND2_X1 U1056 ( .A1(n959), .A2(n958), .ZN(n962) );
  XOR2_X1 U1057 ( .A(G27), .B(n960), .Z(n961) );
  NOR2_X1 U1058 ( .A1(n962), .A2(n961), .ZN(n963) );
  XNOR2_X1 U1059 ( .A(KEYINPUT53), .B(n963), .ZN(n964) );
  XNOR2_X1 U1060 ( .A(KEYINPUT118), .B(n964), .ZN(n965) );
  NOR2_X1 U1061 ( .A1(n966), .A2(n965), .ZN(n968) );
  XOR2_X1 U1062 ( .A(n968), .B(n967), .Z(n969) );
  NAND2_X1 U1063 ( .A1(n970), .A2(n969), .ZN(n971) );
  NAND2_X1 U1064 ( .A1(G11), .A2(n971), .ZN(n1027) );
  XNOR2_X1 U1065 ( .A(G16), .B(KEYINPUT56), .ZN(n997) );
  XOR2_X1 U1066 ( .A(G1348), .B(n972), .Z(n975) );
  XNOR2_X1 U1067 ( .A(n973), .B(G1341), .ZN(n974) );
  NOR2_X1 U1068 ( .A1(n975), .A2(n974), .ZN(n988) );
  XNOR2_X1 U1069 ( .A(KEYINPUT121), .B(n976), .ZN(n983) );
  XOR2_X1 U1070 ( .A(G299), .B(G1956), .Z(n978) );
  NAND2_X1 U1071 ( .A1(n978), .A2(n977), .ZN(n981) );
  XNOR2_X1 U1072 ( .A(G1971), .B(G303), .ZN(n979) );
  XNOR2_X1 U1073 ( .A(KEYINPUT122), .B(n979), .ZN(n980) );
  NOR2_X1 U1074 ( .A1(n981), .A2(n980), .ZN(n982) );
  NAND2_X1 U1075 ( .A1(n983), .A2(n982), .ZN(n984) );
  NOR2_X1 U1076 ( .A1(n985), .A2(n984), .ZN(n986) );
  XOR2_X1 U1077 ( .A(KEYINPUT123), .B(n986), .Z(n987) );
  NAND2_X1 U1078 ( .A1(n988), .A2(n987), .ZN(n990) );
  XNOR2_X1 U1079 ( .A(G171), .B(n1018), .ZN(n989) );
  NOR2_X1 U1080 ( .A1(n990), .A2(n989), .ZN(n995) );
  XNOR2_X1 U1081 ( .A(G1966), .B(G168), .ZN(n992) );
  NAND2_X1 U1082 ( .A1(n992), .A2(n991), .ZN(n993) );
  XNOR2_X1 U1083 ( .A(n993), .B(KEYINPUT57), .ZN(n994) );
  NAND2_X1 U1084 ( .A1(n995), .A2(n994), .ZN(n996) );
  NAND2_X1 U1085 ( .A1(n997), .A2(n996), .ZN(n1025) );
  XOR2_X1 U1086 ( .A(G16), .B(KEYINPUT124), .Z(n1023) );
  XNOR2_X1 U1087 ( .A(KEYINPUT125), .B(G1966), .ZN(n998) );
  XNOR2_X1 U1088 ( .A(n998), .B(G21), .ZN(n1017) );
  XOR2_X1 U1089 ( .A(G1348), .B(KEYINPUT59), .Z(n999) );
  XNOR2_X1 U1090 ( .A(G4), .B(n999), .ZN(n1001) );
  XNOR2_X1 U1091 ( .A(G20), .B(G1956), .ZN(n1000) );
  NOR2_X1 U1092 ( .A1(n1001), .A2(n1000), .ZN(n1005) );
  XNOR2_X1 U1093 ( .A(G1341), .B(G19), .ZN(n1003) );
  XNOR2_X1 U1094 ( .A(G1981), .B(G6), .ZN(n1002) );
  NOR2_X1 U1095 ( .A1(n1003), .A2(n1002), .ZN(n1004) );
  NAND2_X1 U1096 ( .A1(n1005), .A2(n1004), .ZN(n1006) );
  XNOR2_X1 U1097 ( .A(n1006), .B(KEYINPUT60), .ZN(n1015) );
  XNOR2_X1 U1098 ( .A(G1971), .B(G22), .ZN(n1008) );
  XNOR2_X1 U1099 ( .A(G1976), .B(G23), .ZN(n1007) );
  NOR2_X1 U1100 ( .A1(n1008), .A2(n1007), .ZN(n1009) );
  XOR2_X1 U1101 ( .A(KEYINPUT126), .B(n1009), .Z(n1011) );
  XNOR2_X1 U1102 ( .A(G1986), .B(G24), .ZN(n1010) );
  NOR2_X1 U1103 ( .A1(n1011), .A2(n1010), .ZN(n1012) );
  XNOR2_X1 U1104 ( .A(KEYINPUT58), .B(n1012), .ZN(n1013) );
  XNOR2_X1 U1105 ( .A(KEYINPUT127), .B(n1013), .ZN(n1014) );
  NOR2_X1 U1106 ( .A1(n1015), .A2(n1014), .ZN(n1016) );
  NAND2_X1 U1107 ( .A1(n1017), .A2(n1016), .ZN(n1020) );
  XOR2_X1 U1108 ( .A(G5), .B(n1018), .Z(n1019) );
  NOR2_X1 U1109 ( .A1(n1020), .A2(n1019), .ZN(n1021) );
  XNOR2_X1 U1110 ( .A(n1021), .B(KEYINPUT61), .ZN(n1022) );
  NAND2_X1 U1111 ( .A1(n1023), .A2(n1022), .ZN(n1024) );
  NAND2_X1 U1112 ( .A1(n1025), .A2(n1024), .ZN(n1026) );
  NOR2_X1 U1113 ( .A1(n1027), .A2(n1026), .ZN(n1028) );
  NAND2_X1 U1114 ( .A1(n1029), .A2(n1028), .ZN(n1030) );
  XNOR2_X1 U1115 ( .A(KEYINPUT62), .B(n1030), .ZN(G150) );
  INV_X1 U1116 ( .A(G150), .ZN(G311) );
endmodule

