

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363,
         n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374,
         n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385,
         n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n396,
         n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407,
         n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418,
         n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429,
         n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440,
         n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451,
         n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462,
         n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473,
         n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484,
         n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495,
         n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506,
         n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517,
         n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528,
         n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539,
         n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550,
         n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561,
         n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572,
         n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583,
         n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594,
         n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605,
         n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616,
         n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627,
         n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, n638,
         n639, n640, n641, n642, n643, n644, n645, n646, n647, n648, n649,
         n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, n660,
         n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, n671,
         n672, n673, n674, n675, n676, n677, n678, n679, n680, n681, n682,
         n683, n684, n685, n686, n687, n688, n689, n690, n691, n692, n693,
         n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, n704,
         n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n715,
         n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726,
         n727, n728, n729, n730, n731, n732, n733, n734, n735, n736, n737,
         n738, n739, n740, n741, n742, n743, n744, n745, n746, n747, n748,
         n749, n750, n751, n752, n753, n754, n755, n756, n757, n758, n759,
         n760, n761, n762;

  BUF_X1 U374 ( .A(n724), .Z(n353) );
  NOR2_X1 U375 ( .A1(n651), .A2(n652), .ZN(n555) );
  NAND2_X1 U376 ( .A1(n383), .A2(n382), .ZN(n581) );
  XNOR2_X1 U377 ( .A(n752), .B(G146), .ZN(n540) );
  XNOR2_X2 U378 ( .A(n375), .B(n516), .ZN(n752) );
  XNOR2_X2 U379 ( .A(n444), .B(n486), .ZN(n375) );
  XNOR2_X1 U380 ( .A(G110), .B(G128), .ZN(n396) );
  AND2_X2 U381 ( .A1(n381), .A2(n379), .ZN(n378) );
  XNOR2_X2 U382 ( .A(n416), .B(KEYINPUT32), .ZN(n762) );
  NOR2_X2 U383 ( .A1(n591), .A2(n590), .ZN(n410) );
  XNOR2_X2 U384 ( .A(n447), .B(n363), .ZN(n567) );
  NAND2_X2 U385 ( .A1(n378), .A2(n376), .ZN(n447) );
  XNOR2_X2 U386 ( .A(n511), .B(n510), .ZN(n553) );
  NOR2_X2 U387 ( .A1(G902), .A2(n689), .ZN(n511) );
  NAND2_X1 U388 ( .A1(n546), .A2(n645), .ZN(n393) );
  OR2_X2 U389 ( .A1(n682), .A2(G902), .ZN(n543) );
  NOR2_X1 U390 ( .A1(n449), .A2(n419), .ZN(n418) );
  NAND2_X1 U391 ( .A1(n399), .A2(n397), .ZN(n753) );
  NAND2_X1 U392 ( .A1(n377), .A2(n549), .ZN(n376) );
  NOR2_X1 U393 ( .A1(n596), .A2(n632), .ZN(n417) );
  INV_X1 U394 ( .A(n554), .ZN(n354) );
  NOR2_X1 U395 ( .A1(n652), .A2(n581), .ZN(n557) );
  AND2_X2 U396 ( .A1(n553), .A2(n552), .ZN(n602) );
  XNOR2_X1 U397 ( .A(n623), .B(n572), .ZN(n632) );
  XOR2_X1 U398 ( .A(n544), .B(n647), .Z(n603) );
  XNOR2_X1 U399 ( .A(n455), .B(n527), .ZN(n737) );
  XNOR2_X1 U400 ( .A(n467), .B(n466), .ZN(n535) );
  XNOR2_X1 U401 ( .A(n465), .B(G119), .ZN(n467) );
  INV_X4 U402 ( .A(G953), .ZN(n754) );
  XNOR2_X1 U403 ( .A(G146), .B(G125), .ZN(n497) );
  XNOR2_X1 U404 ( .A(G101), .B(G116), .ZN(n466) );
  XNOR2_X1 U405 ( .A(KEYINPUT64), .B(KEYINPUT4), .ZN(n444) );
  INV_X1 U406 ( .A(KEYINPUT3), .ZN(n465) );
  INV_X1 U407 ( .A(n723), .ZN(n730) );
  NAND2_X1 U408 ( .A1(n673), .A2(n672), .ZN(n723) );
  NAND2_X1 U409 ( .A1(n631), .A2(n745), .ZN(n672) );
  XNOR2_X1 U410 ( .A(n581), .B(KEYINPUT1), .ZN(n651) );
  AND2_X1 U411 ( .A1(n442), .A2(n570), .ZN(n441) );
  XNOR2_X1 U412 ( .A(n373), .B(KEYINPUT83), .ZN(n372) );
  XNOR2_X1 U413 ( .A(G137), .B(G134), .ZN(n516) );
  XNOR2_X1 U414 ( .A(n473), .B(n472), .ZN(n571) );
  XNOR2_X1 U415 ( .A(n471), .B(KEYINPUT90), .ZN(n472) );
  XNOR2_X1 U416 ( .A(n430), .B(n429), .ZN(n631) );
  INV_X1 U417 ( .A(KEYINPUT79), .ZN(n429) );
  NOR2_X1 U418 ( .A1(n753), .A2(n431), .ZN(n430) );
  XNOR2_X1 U419 ( .A(n515), .B(n446), .ZN(n405) );
  INV_X1 U420 ( .A(KEYINPUT22), .ZN(n446) );
  XNOR2_X1 U421 ( .A(n564), .B(KEYINPUT85), .ZN(n569) );
  XNOR2_X1 U422 ( .A(n368), .B(n428), .ZN(n404) );
  INV_X1 U423 ( .A(KEYINPUT48), .ZN(n428) );
  NAND2_X1 U424 ( .A1(n374), .A2(n439), .ZN(n373) );
  AND2_X1 U425 ( .A1(n560), .A2(n440), .ZN(n439) );
  XNOR2_X1 U426 ( .A(n550), .B(KEYINPUT84), .ZN(n374) );
  INV_X1 U427 ( .A(G902), .ZN(n386) );
  NAND2_X1 U428 ( .A1(n722), .A2(G902), .ZN(n387) );
  NAND2_X1 U429 ( .A1(n721), .A2(KEYINPUT80), .ZN(n401) );
  INV_X1 U430 ( .A(n761), .ZN(n426) );
  INV_X1 U431 ( .A(n404), .ZN(n398) );
  XNOR2_X1 U432 ( .A(KEYINPUT12), .B(KEYINPUT11), .ZN(n499) );
  XOR2_X1 U433 ( .A(KEYINPUT99), .B(KEYINPUT100), .Z(n500) );
  XNOR2_X1 U434 ( .A(G143), .B(G122), .ZN(n501) );
  INV_X1 U435 ( .A(n753), .ZN(n630) );
  NOR2_X1 U436 ( .A1(n578), .A2(n590), .ZN(n606) );
  NOR2_X1 U437 ( .A1(n737), .A2(G902), .ZN(n394) );
  XNOR2_X1 U438 ( .A(KEYINPUT70), .B(KEYINPUT5), .ZN(n532) );
  XNOR2_X1 U439 ( .A(G131), .B(G113), .ZN(n533) );
  INV_X1 U440 ( .A(KEYINPUT71), .ZN(n503) );
  NOR2_X1 U441 ( .A1(G953), .A2(G237), .ZN(n504) );
  XOR2_X1 U442 ( .A(G122), .B(G107), .Z(n488) );
  XNOR2_X1 U443 ( .A(n396), .B(n395), .ZN(n456) );
  XNOR2_X1 U444 ( .A(G119), .B(G137), .ZN(n395) );
  XNOR2_X1 U445 ( .A(n497), .B(KEYINPUT10), .ZN(n523) );
  XOR2_X1 U446 ( .A(G116), .B(KEYINPUT102), .Z(n487) );
  XNOR2_X1 U447 ( .A(n740), .B(n406), .ZN(n674) );
  XNOR2_X1 U448 ( .A(n407), .B(n470), .ZN(n406) );
  XNOR2_X1 U449 ( .A(n375), .B(n408), .ZN(n407) );
  NAND2_X1 U450 ( .A1(n434), .A2(n432), .ZN(n584) );
  AND2_X1 U451 ( .A1(n435), .A2(n437), .ZN(n434) );
  NAND2_X1 U452 ( .A1(n433), .A2(n436), .ZN(n432) );
  XNOR2_X1 U453 ( .A(n509), .B(n687), .ZN(n510) );
  XNOR2_X1 U454 ( .A(n557), .B(KEYINPUT96), .ZN(n592) );
  BUF_X1 U455 ( .A(n647), .Z(n411) );
  INV_X1 U456 ( .A(KEYINPUT65), .ZN(n670) );
  XNOR2_X1 U457 ( .A(n540), .B(n522), .ZN(n724) );
  NAND2_X1 U458 ( .A1(n730), .A2(G210), .ZN(n425) );
  INV_X1 U459 ( .A(KEYINPUT47), .ZN(n412) );
  NOR2_X1 U460 ( .A1(n569), .A2(n565), .ZN(n443) );
  NAND2_X1 U461 ( .A1(G234), .A2(G237), .ZN(n477) );
  AND2_X1 U462 ( .A1(n635), .A2(n587), .ZN(n438) );
  OR2_X1 U463 ( .A1(G237), .A2(G902), .ZN(n474) );
  XNOR2_X1 U464 ( .A(KEYINPUT17), .B(KEYINPUT18), .ZN(n408) );
  NOR2_X1 U465 ( .A1(n630), .A2(KEYINPUT2), .ZN(n452) );
  AND2_X1 U466 ( .A1(n438), .A2(KEYINPUT41), .ZN(n436) );
  OR2_X1 U467 ( .A1(n438), .A2(KEYINPUT41), .ZN(n437) );
  OR2_X1 U468 ( .A1(n724), .A2(n385), .ZN(n382) );
  AND2_X1 U469 ( .A1(n384), .A2(n387), .ZN(n383) );
  NAND2_X1 U470 ( .A1(G469), .A2(n386), .ZN(n385) );
  AND2_X1 U471 ( .A1(n402), .A2(n400), .ZN(n399) );
  NAND2_X1 U472 ( .A1(n398), .A2(KEYINPUT80), .ZN(n397) );
  AND2_X1 U473 ( .A1(n401), .A2(n426), .ZN(n400) );
  XNOR2_X1 U474 ( .A(n508), .B(n507), .ZN(n689) );
  XNOR2_X1 U475 ( .A(n750), .B(n461), .ZN(n508) );
  NAND2_X1 U476 ( .A1(n459), .A2(KEYINPUT2), .ZN(n457) );
  XOR2_X1 U477 ( .A(G131), .B(G140), .Z(n519) );
  XOR2_X1 U478 ( .A(G110), .B(G107), .Z(n518) );
  XNOR2_X1 U479 ( .A(G101), .B(G104), .ZN(n517) );
  INV_X1 U480 ( .A(n584), .ZN(n666) );
  AND2_X1 U481 ( .A1(n380), .A2(n361), .ZN(n379) );
  NAND2_X1 U482 ( .A1(n354), .A2(n549), .ZN(n380) );
  BUF_X1 U483 ( .A(n546), .Z(n574) );
  XNOR2_X1 U484 ( .A(n540), .B(n539), .ZN(n682) );
  XNOR2_X1 U485 ( .A(n409), .B(n468), .ZN(n740) );
  XNOR2_X1 U486 ( .A(n535), .B(n356), .ZN(n409) );
  XNOR2_X1 U487 ( .A(n526), .B(n456), .ZN(n455) );
  XNOR2_X1 U488 ( .A(n414), .B(n491), .ZN(n731) );
  XNOR2_X1 U489 ( .A(n357), .B(n494), .ZN(n414) );
  XOR2_X1 U490 ( .A(KEYINPUT9), .B(KEYINPUT7), .Z(n490) );
  NOR2_X1 U491 ( .A1(n584), .A2(n610), .ZN(n586) );
  NOR2_X1 U492 ( .A1(n621), .A2(n623), .ZN(n607) );
  NAND2_X1 U493 ( .A1(n405), .A2(n464), .ZN(n416) );
  XNOR2_X1 U494 ( .A(n556), .B(n415), .ZN(n716) );
  XNOR2_X1 U495 ( .A(KEYINPUT98), .B(KEYINPUT31), .ZN(n415) );
  XNOR2_X1 U496 ( .A(n602), .B(n413), .ZN(n710) );
  INV_X1 U497 ( .A(KEYINPUT107), .ZN(n413) );
  XNOR2_X1 U498 ( .A(n392), .B(KEYINPUT109), .ZN(n597) );
  AND2_X1 U499 ( .A1(n592), .A2(n391), .ZN(n370) );
  XNOR2_X1 U500 ( .A(n725), .B(n420), .ZN(n729) );
  XNOR2_X1 U501 ( .A(n353), .B(n728), .ZN(n420) );
  INV_X1 U502 ( .A(KEYINPUT56), .ZN(n422) );
  XOR2_X1 U503 ( .A(G140), .B(KEYINPUT24), .Z(n355) );
  XNOR2_X1 U504 ( .A(G110), .B(KEYINPUT16), .ZN(n356) );
  XOR2_X1 U505 ( .A(n486), .B(n487), .Z(n357) );
  XOR2_X1 U506 ( .A(KEYINPUT94), .B(KEYINPUT23), .Z(n358) );
  AND2_X1 U507 ( .A1(n745), .A2(n630), .ZN(n359) );
  BUF_X1 U508 ( .A(n571), .Z(n623) );
  OR2_X1 U509 ( .A1(n359), .A2(n628), .ZN(n360) );
  AND2_X1 U510 ( .A1(n551), .A2(n553), .ZN(n361) );
  AND2_X1 U511 ( .A1(n554), .A2(n448), .ZN(n362) );
  XNOR2_X1 U512 ( .A(KEYINPUT72), .B(KEYINPUT35), .ZN(n363) );
  XOR2_X1 U513 ( .A(KEYINPUT82), .B(KEYINPUT39), .Z(n364) );
  INV_X1 U514 ( .A(KEYINPUT41), .ZN(n454) );
  XNOR2_X1 U515 ( .A(n676), .B(n675), .ZN(n365) );
  INV_X1 U516 ( .A(n669), .ZN(n459) );
  XNOR2_X1 U517 ( .A(G902), .B(KEYINPUT15), .ZN(n669) );
  INV_X1 U518 ( .A(KEYINPUT2), .ZN(n431) );
  XOR2_X1 U519 ( .A(KEYINPUT53), .B(KEYINPUT122), .Z(n366) );
  XNOR2_X1 U520 ( .A(n678), .B(KEYINPUT89), .ZN(n739) );
  XNOR2_X2 U521 ( .A(n367), .B(KEYINPUT45), .ZN(n629) );
  NAND2_X1 U522 ( .A1(n441), .A2(n372), .ZN(n367) );
  INV_X1 U523 ( .A(n620), .ZN(n445) );
  XNOR2_X1 U524 ( .A(n671), .B(n670), .ZN(n673) );
  NAND2_X1 U525 ( .A1(n369), .A2(n457), .ZN(n671) );
  NAND2_X1 U526 ( .A1(n618), .A2(n619), .ZN(n368) );
  NOR2_X1 U527 ( .A1(n753), .A2(n669), .ZN(n458) );
  XNOR2_X1 U528 ( .A(n425), .B(n365), .ZN(n424) );
  NAND2_X1 U529 ( .A1(n458), .A2(n629), .ZN(n369) );
  NAND2_X1 U530 ( .A1(n370), .A2(n410), .ZN(n392) );
  XNOR2_X1 U531 ( .A(n601), .B(n600), .ZN(n617) );
  BUF_X2 U532 ( .A(n629), .Z(n745) );
  NAND2_X1 U533 ( .A1(n371), .A2(n668), .ZN(n390) );
  NAND2_X1 U534 ( .A1(n418), .A2(n360), .ZN(n371) );
  NAND2_X2 U535 ( .A1(n597), .A2(n361), .ZN(n709) );
  INV_X1 U536 ( .A(n642), .ZN(n377) );
  NAND2_X1 U537 ( .A1(n642), .A2(n362), .ZN(n381) );
  XNOR2_X2 U538 ( .A(n548), .B(KEYINPUT33), .ZN(n642) );
  NAND2_X1 U539 ( .A1(n724), .A2(n722), .ZN(n384) );
  XNOR2_X1 U540 ( .A(n388), .B(n366), .ZN(G75) );
  NAND2_X1 U541 ( .A1(n389), .A2(n754), .ZN(n388) );
  XNOR2_X1 U542 ( .A(n390), .B(KEYINPUT121), .ZN(n389) );
  NAND2_X1 U543 ( .A1(n592), .A2(n410), .ZN(n596) );
  INV_X1 U544 ( .A(n623), .ZN(n391) );
  XNOR2_X2 U545 ( .A(n393), .B(KEYINPUT68), .ZN(n652) );
  XNOR2_X1 U546 ( .A(n394), .B(n531), .ZN(n546) );
  NAND2_X1 U547 ( .A1(n404), .A2(n403), .ZN(n402) );
  AND2_X1 U548 ( .A1(n427), .A2(n625), .ZN(n403) );
  AND2_X1 U549 ( .A1(n405), .A2(n445), .ZN(n563) );
  NAND2_X1 U550 ( .A1(n674), .A2(n669), .ZN(n473) );
  NOR2_X1 U551 ( .A1(n667), .A2(n460), .ZN(n668) );
  AND2_X1 U552 ( .A1(n451), .A2(n450), .ZN(n449) );
  NAND2_X1 U553 ( .A1(n554), .A2(n514), .ZN(n515) );
  XNOR2_X1 U554 ( .A(n711), .B(n412), .ZN(n614) );
  NOR2_X1 U555 ( .A1(n610), .A2(n611), .ZN(n711) );
  NOR2_X1 U556 ( .A1(n571), .A2(n633), .ZN(n476) );
  NAND2_X1 U557 ( .A1(n603), .A2(n710), .ZN(n604) );
  XNOR2_X1 U558 ( .A(n417), .B(n364), .ZN(n626) );
  INV_X1 U559 ( .A(n672), .ZN(n419) );
  NAND2_X1 U560 ( .A1(n421), .A2(n453), .ZN(n595) );
  XNOR2_X1 U561 ( .A(n421), .B(G131), .ZN(G33) );
  XNOR2_X2 U562 ( .A(n593), .B(KEYINPUT40), .ZN(n421) );
  XNOR2_X1 U563 ( .A(n423), .B(n422), .ZN(G51) );
  NAND2_X1 U564 ( .A1(n424), .A2(n692), .ZN(n423) );
  INV_X1 U565 ( .A(n721), .ZN(n427) );
  INV_X1 U566 ( .A(n632), .ZN(n433) );
  NAND2_X1 U567 ( .A1(n632), .A2(n454), .ZN(n435) );
  NOR2_X1 U568 ( .A1(n632), .A2(n633), .ZN(n638) );
  INV_X1 U569 ( .A(n696), .ZN(n440) );
  XNOR2_X1 U570 ( .A(n443), .B(n566), .ZN(n442) );
  XNOR2_X2 U571 ( .A(G143), .B(G128), .ZN(n486) );
  NAND2_X1 U572 ( .A1(n567), .A2(KEYINPUT44), .ZN(n550) );
  INV_X1 U573 ( .A(n549), .ZN(n448) );
  INV_X1 U574 ( .A(KEYINPUT78), .ZN(n450) );
  NAND2_X1 U575 ( .A1(n745), .A2(n452), .ZN(n451) );
  XNOR2_X1 U576 ( .A(n586), .B(n585), .ZN(n453) );
  XNOR2_X1 U577 ( .A(n453), .B(G137), .ZN(G39) );
  XNOR2_X1 U578 ( .A(n358), .B(n355), .ZN(n524) );
  NOR2_X2 U579 ( .A1(n611), .A2(n483), .ZN(n485) );
  AND2_X1 U580 ( .A1(n642), .A2(n666), .ZN(n460) );
  XOR2_X1 U581 ( .A(n500), .B(n499), .Z(n461) );
  AND2_X1 U582 ( .A1(G227), .A2(n754), .ZN(n462) );
  OR2_X1 U583 ( .A1(n644), .A2(n445), .ZN(n463) );
  NOR2_X1 U584 ( .A1(n561), .A2(n463), .ZN(n464) );
  INV_X1 U585 ( .A(KEYINPUT75), .ZN(n600) );
  INV_X1 U586 ( .A(KEYINPUT66), .ZN(n566) );
  INV_X1 U587 ( .A(KEYINPUT80), .ZN(n625) );
  XNOR2_X1 U588 ( .A(n519), .B(n462), .ZN(n520) );
  INV_X1 U589 ( .A(KEYINPUT42), .ZN(n585) );
  XNOR2_X1 U590 ( .A(G113), .B(G104), .ZN(n502) );
  XOR2_X1 U591 ( .A(n502), .B(n488), .Z(n468) );
  NAND2_X1 U592 ( .A1(G224), .A2(n754), .ZN(n469) );
  XNOR2_X1 U593 ( .A(n497), .B(n469), .ZN(n470) );
  NAND2_X1 U594 ( .A1(n474), .A2(G210), .ZN(n471) );
  NAND2_X1 U595 ( .A1(n474), .A2(G214), .ZN(n475) );
  XNOR2_X1 U596 ( .A(n475), .B(KEYINPUT91), .ZN(n633) );
  XNOR2_X1 U597 ( .A(n476), .B(KEYINPUT19), .ZN(n611) );
  XOR2_X1 U598 ( .A(KEYINPUT14), .B(KEYINPUT92), .Z(n478) );
  XOR2_X1 U599 ( .A(n478), .B(n477), .Z(n480) );
  NAND2_X1 U600 ( .A1(n480), .A2(G952), .ZN(n479) );
  XOR2_X1 U601 ( .A(KEYINPUT93), .B(n479), .Z(n664) );
  NOR2_X1 U602 ( .A1(n664), .A2(G953), .ZN(n577) );
  AND2_X1 U603 ( .A1(n480), .A2(G953), .ZN(n481) );
  NAND2_X1 U604 ( .A1(G902), .A2(n481), .ZN(n575) );
  NOR2_X1 U605 ( .A1(G898), .A2(n575), .ZN(n482) );
  NOR2_X1 U606 ( .A1(n577), .A2(n482), .ZN(n483) );
  XOR2_X1 U607 ( .A(KEYINPUT67), .B(KEYINPUT0), .Z(n484) );
  XNOR2_X2 U608 ( .A(n485), .B(n484), .ZN(n554) );
  XNOR2_X1 U609 ( .A(G134), .B(n488), .ZN(n489) );
  XNOR2_X1 U610 ( .A(n490), .B(n489), .ZN(n491) );
  NAND2_X1 U611 ( .A1(n754), .A2(G234), .ZN(n493) );
  XNOR2_X1 U612 ( .A(KEYINPUT77), .B(KEYINPUT8), .ZN(n492) );
  XNOR2_X1 U613 ( .A(n493), .B(n492), .ZN(n525) );
  NAND2_X1 U614 ( .A1(G217), .A2(n525), .ZN(n494) );
  NOR2_X1 U615 ( .A1(G902), .A2(n731), .ZN(n496) );
  XNOR2_X1 U616 ( .A(KEYINPUT103), .B(G478), .ZN(n495) );
  XNOR2_X1 U617 ( .A(n496), .B(n495), .ZN(n551) );
  INV_X1 U618 ( .A(n519), .ZN(n498) );
  XNOR2_X1 U619 ( .A(n523), .B(n498), .ZN(n750) );
  XNOR2_X1 U620 ( .A(n502), .B(n501), .ZN(n506) );
  XNOR2_X1 U621 ( .A(n504), .B(n503), .ZN(n536) );
  NAND2_X1 U622 ( .A1(n536), .A2(G214), .ZN(n505) );
  XNOR2_X1 U623 ( .A(n506), .B(n505), .ZN(n507) );
  XNOR2_X1 U624 ( .A(KEYINPUT101), .B(KEYINPUT13), .ZN(n509) );
  INV_X1 U625 ( .A(G475), .ZN(n687) );
  NOR2_X1 U626 ( .A1(n551), .A2(n553), .ZN(n635) );
  NAND2_X1 U627 ( .A1(G234), .A2(n669), .ZN(n512) );
  XNOR2_X1 U628 ( .A(KEYINPUT20), .B(n512), .ZN(n528) );
  NAND2_X1 U629 ( .A1(n528), .A2(G221), .ZN(n513) );
  XOR2_X1 U630 ( .A(KEYINPUT21), .B(n513), .Z(n645) );
  AND2_X1 U631 ( .A1(n635), .A2(n645), .ZN(n514) );
  XNOR2_X1 U632 ( .A(n518), .B(n517), .ZN(n521) );
  XNOR2_X1 U633 ( .A(n521), .B(n520), .ZN(n522) );
  INV_X1 U634 ( .A(G469), .ZN(n722) );
  INV_X1 U635 ( .A(n651), .ZN(n620) );
  XNOR2_X1 U636 ( .A(n524), .B(n523), .ZN(n527) );
  NAND2_X1 U637 ( .A1(G221), .A2(n525), .ZN(n526) );
  XOR2_X1 U638 ( .A(KEYINPUT25), .B(KEYINPUT95), .Z(n530) );
  NAND2_X1 U639 ( .A1(n528), .A2(G217), .ZN(n529) );
  XNOR2_X1 U640 ( .A(n530), .B(n529), .ZN(n531) );
  XOR2_X1 U641 ( .A(n574), .B(KEYINPUT105), .Z(n644) );
  NAND2_X1 U642 ( .A1(n563), .A2(n644), .ZN(n545) );
  XNOR2_X1 U643 ( .A(KEYINPUT104), .B(KEYINPUT6), .ZN(n544) );
  XNOR2_X1 U644 ( .A(n533), .B(n532), .ZN(n534) );
  XNOR2_X1 U645 ( .A(n535), .B(n534), .ZN(n538) );
  AND2_X1 U646 ( .A1(n536), .A2(G210), .ZN(n537) );
  XNOR2_X1 U647 ( .A(n538), .B(n537), .ZN(n539) );
  XNOR2_X1 U648 ( .A(G472), .B(KEYINPUT97), .ZN(n541) );
  XNOR2_X1 U649 ( .A(n541), .B(KEYINPUT69), .ZN(n542) );
  XNOR2_X2 U650 ( .A(n543), .B(n542), .ZN(n647) );
  NOR2_X1 U651 ( .A1(n545), .A2(n603), .ZN(n696) );
  XOR2_X1 U652 ( .A(KEYINPUT34), .B(KEYINPUT73), .Z(n549) );
  XNOR2_X1 U653 ( .A(n555), .B(KEYINPUT106), .ZN(n547) );
  NAND2_X1 U654 ( .A1(n547), .A2(n603), .ZN(n548) );
  INV_X1 U655 ( .A(n551), .ZN(n552) );
  NOR2_X1 U656 ( .A1(n553), .A2(n552), .ZN(n706) );
  NOR2_X1 U657 ( .A1(n602), .A2(n706), .ZN(n612) );
  INV_X1 U658 ( .A(n612), .ZN(n637) );
  NAND2_X1 U659 ( .A1(n555), .A2(n411), .ZN(n656) );
  NOR2_X1 U660 ( .A1(n354), .A2(n656), .ZN(n556) );
  NOR2_X1 U661 ( .A1(n354), .A2(n411), .ZN(n558) );
  NAND2_X1 U662 ( .A1(n558), .A2(n592), .ZN(n700) );
  NAND2_X1 U663 ( .A1(n716), .A2(n700), .ZN(n559) );
  NAND2_X1 U664 ( .A1(n637), .A2(n559), .ZN(n560) );
  XNOR2_X1 U665 ( .A(n603), .B(KEYINPUT74), .ZN(n561) );
  NOR2_X1 U666 ( .A1(n574), .A2(n411), .ZN(n562) );
  NAND2_X1 U667 ( .A1(n563), .A2(n562), .ZN(n705) );
  NAND2_X1 U668 ( .A1(n762), .A2(n705), .ZN(n564) );
  INV_X1 U669 ( .A(KEYINPUT44), .ZN(n565) );
  NOR2_X1 U670 ( .A1(KEYINPUT44), .A2(n567), .ZN(n568) );
  NAND2_X1 U671 ( .A1(n569), .A2(n568), .ZN(n570) );
  INV_X1 U672 ( .A(KEYINPUT38), .ZN(n572) );
  INV_X1 U673 ( .A(n645), .ZN(n573) );
  OR2_X1 U674 ( .A1(n574), .A2(n573), .ZN(n578) );
  NOR2_X1 U675 ( .A1(n575), .A2(G900), .ZN(n576) );
  NOR2_X1 U676 ( .A1(n577), .A2(n576), .ZN(n590) );
  NAND2_X1 U677 ( .A1(n606), .A2(n411), .ZN(n580) );
  INV_X1 U678 ( .A(KEYINPUT28), .ZN(n579) );
  XNOR2_X1 U679 ( .A(n580), .B(n579), .ZN(n583) );
  INV_X1 U680 ( .A(n581), .ZN(n582) );
  NAND2_X1 U681 ( .A1(n583), .A2(n582), .ZN(n610) );
  INV_X1 U682 ( .A(n633), .ZN(n587) );
  NAND2_X1 U683 ( .A1(n647), .A2(n587), .ZN(n589) );
  XNOR2_X1 U684 ( .A(KEYINPUT108), .B(KEYINPUT30), .ZN(n588) );
  XNOR2_X1 U685 ( .A(n589), .B(n588), .ZN(n591) );
  NAND2_X1 U686 ( .A1(n626), .A2(n602), .ZN(n593) );
  XNOR2_X1 U687 ( .A(KEYINPUT81), .B(KEYINPUT46), .ZN(n594) );
  XNOR2_X1 U688 ( .A(n595), .B(n594), .ZN(n619) );
  XNOR2_X1 U689 ( .A(n709), .B(KEYINPUT76), .ZN(n599) );
  NAND2_X1 U690 ( .A1(n612), .A2(KEYINPUT47), .ZN(n598) );
  NAND2_X1 U691 ( .A1(n599), .A2(n598), .ZN(n601) );
  XOR2_X1 U692 ( .A(KEYINPUT110), .B(KEYINPUT36), .Z(n608) );
  NOR2_X1 U693 ( .A1(n633), .A2(n604), .ZN(n605) );
  NAND2_X1 U694 ( .A1(n606), .A2(n605), .ZN(n621) );
  XOR2_X1 U695 ( .A(n608), .B(n607), .Z(n609) );
  NAND2_X1 U696 ( .A1(n609), .A2(n620), .ZN(n719) );
  NAND2_X1 U697 ( .A1(n711), .A2(n612), .ZN(n613) );
  NAND2_X1 U698 ( .A1(n614), .A2(n613), .ZN(n615) );
  NAND2_X1 U699 ( .A1(n719), .A2(n615), .ZN(n616) );
  NOR2_X1 U700 ( .A1(n617), .A2(n616), .ZN(n618) );
  NOR2_X1 U701 ( .A1(n621), .A2(n620), .ZN(n622) );
  XNOR2_X1 U702 ( .A(n622), .B(KEYINPUT43), .ZN(n624) );
  NOR2_X1 U703 ( .A1(n624), .A2(n391), .ZN(n721) );
  NAND2_X1 U704 ( .A1(n626), .A2(n706), .ZN(n627) );
  XNOR2_X1 U705 ( .A(n627), .B(KEYINPUT111), .ZN(n761) );
  NAND2_X1 U706 ( .A1(n431), .A2(KEYINPUT78), .ZN(n628) );
  NAND2_X1 U707 ( .A1(n633), .A2(n632), .ZN(n634) );
  NAND2_X1 U708 ( .A1(n635), .A2(n634), .ZN(n636) );
  XNOR2_X1 U709 ( .A(KEYINPUT118), .B(n636), .ZN(n641) );
  NAND2_X1 U710 ( .A1(n638), .A2(n637), .ZN(n639) );
  XOR2_X1 U711 ( .A(KEYINPUT119), .B(n639), .Z(n640) );
  NAND2_X1 U712 ( .A1(n641), .A2(n640), .ZN(n643) );
  NAND2_X1 U713 ( .A1(n643), .A2(n642), .ZN(n661) );
  NOR2_X1 U714 ( .A1(n645), .A2(n644), .ZN(n646) );
  XNOR2_X1 U715 ( .A(n646), .B(KEYINPUT49), .ZN(n649) );
  INV_X1 U716 ( .A(n411), .ZN(n648) );
  NAND2_X1 U717 ( .A1(n649), .A2(n648), .ZN(n650) );
  XNOR2_X1 U718 ( .A(n650), .B(KEYINPUT117), .ZN(n655) );
  NAND2_X1 U719 ( .A1(n652), .A2(n445), .ZN(n653) );
  XNOR2_X1 U720 ( .A(n653), .B(KEYINPUT50), .ZN(n654) );
  NAND2_X1 U721 ( .A1(n655), .A2(n654), .ZN(n657) );
  NAND2_X1 U722 ( .A1(n657), .A2(n656), .ZN(n658) );
  XOR2_X1 U723 ( .A(KEYINPUT51), .B(n658), .Z(n659) );
  NAND2_X1 U724 ( .A1(n666), .A2(n659), .ZN(n660) );
  NAND2_X1 U725 ( .A1(n661), .A2(n660), .ZN(n662) );
  XNOR2_X1 U726 ( .A(n662), .B(KEYINPUT52), .ZN(n663) );
  XOR2_X1 U727 ( .A(KEYINPUT120), .B(n663), .Z(n665) );
  NOR2_X1 U728 ( .A1(n665), .A2(n664), .ZN(n667) );
  XOR2_X1 U729 ( .A(KEYINPUT86), .B(KEYINPUT55), .Z(n676) );
  XNOR2_X1 U730 ( .A(n674), .B(KEYINPUT54), .ZN(n675) );
  INV_X1 U731 ( .A(G952), .ZN(n677) );
  NAND2_X1 U732 ( .A1(n677), .A2(G953), .ZN(n678) );
  INV_X1 U733 ( .A(G472), .ZN(n679) );
  NOR2_X1 U734 ( .A1(n723), .A2(n679), .ZN(n684) );
  XOR2_X1 U735 ( .A(KEYINPUT87), .B(KEYINPUT112), .Z(n680) );
  XNOR2_X1 U736 ( .A(n680), .B(KEYINPUT62), .ZN(n681) );
  XNOR2_X1 U737 ( .A(n682), .B(n681), .ZN(n683) );
  XNOR2_X1 U738 ( .A(n684), .B(n683), .ZN(n685) );
  INV_X1 U739 ( .A(n739), .ZN(n692) );
  NAND2_X1 U740 ( .A1(n685), .A2(n692), .ZN(n686) );
  XNOR2_X1 U741 ( .A(n686), .B(KEYINPUT63), .ZN(G57) );
  NOR2_X1 U742 ( .A1(n723), .A2(n687), .ZN(n691) );
  XOR2_X1 U743 ( .A(KEYINPUT88), .B(KEYINPUT59), .Z(n688) );
  XNOR2_X1 U744 ( .A(n689), .B(n688), .ZN(n690) );
  XNOR2_X1 U745 ( .A(n691), .B(n690), .ZN(n693) );
  NAND2_X1 U746 ( .A1(n693), .A2(n692), .ZN(n695) );
  INV_X1 U747 ( .A(KEYINPUT60), .ZN(n694) );
  XNOR2_X1 U748 ( .A(n695), .B(n694), .ZN(G60) );
  XOR2_X1 U749 ( .A(G101), .B(n696), .Z(G3) );
  INV_X1 U750 ( .A(n710), .ZN(n713) );
  NOR2_X1 U751 ( .A1(n700), .A2(n713), .ZN(n697) );
  XOR2_X1 U752 ( .A(G104), .B(n697), .Z(G6) );
  XOR2_X1 U753 ( .A(KEYINPUT115), .B(KEYINPUT27), .Z(n699) );
  XNOR2_X1 U754 ( .A(KEYINPUT113), .B(KEYINPUT114), .ZN(n698) );
  XNOR2_X1 U755 ( .A(n699), .B(n698), .ZN(n704) );
  INV_X1 U756 ( .A(n706), .ZN(n715) );
  NOR2_X1 U757 ( .A1(n700), .A2(n715), .ZN(n702) );
  XNOR2_X1 U758 ( .A(G107), .B(KEYINPUT26), .ZN(n701) );
  XNOR2_X1 U759 ( .A(n702), .B(n701), .ZN(n703) );
  XOR2_X1 U760 ( .A(n704), .B(n703), .Z(G9) );
  XNOR2_X1 U761 ( .A(G110), .B(n705), .ZN(G12) );
  XOR2_X1 U762 ( .A(G128), .B(KEYINPUT29), .Z(n708) );
  NAND2_X1 U763 ( .A1(n711), .A2(n706), .ZN(n707) );
  XNOR2_X1 U764 ( .A(n708), .B(n707), .ZN(G30) );
  XNOR2_X1 U765 ( .A(n709), .B(G143), .ZN(G45) );
  NAND2_X1 U766 ( .A1(n711), .A2(n710), .ZN(n712) );
  XNOR2_X1 U767 ( .A(n712), .B(G146), .ZN(G48) );
  NOR2_X1 U768 ( .A1(n716), .A2(n713), .ZN(n714) );
  XOR2_X1 U769 ( .A(G113), .B(n714), .Z(G15) );
  NOR2_X1 U770 ( .A1(n716), .A2(n715), .ZN(n717) );
  XOR2_X1 U771 ( .A(G116), .B(n717), .Z(G18) );
  XOR2_X1 U772 ( .A(KEYINPUT37), .B(KEYINPUT116), .Z(n718) );
  XNOR2_X1 U773 ( .A(n719), .B(n718), .ZN(n720) );
  XNOR2_X1 U774 ( .A(G125), .B(n720), .ZN(G27) );
  XOR2_X1 U775 ( .A(G140), .B(n721), .Z(G42) );
  NOR2_X1 U776 ( .A1(n723), .A2(n722), .ZN(n725) );
  XOR2_X1 U777 ( .A(KEYINPUT58), .B(KEYINPUT57), .Z(n727) );
  XNOR2_X1 U778 ( .A(KEYINPUT124), .B(KEYINPUT123), .ZN(n726) );
  XNOR2_X1 U779 ( .A(n727), .B(n726), .ZN(n728) );
  NOR2_X1 U780 ( .A1(n739), .A2(n729), .ZN(G54) );
  BUF_X2 U781 ( .A(n730), .Z(n735) );
  NAND2_X1 U782 ( .A1(n735), .A2(G478), .ZN(n733) );
  XOR2_X1 U783 ( .A(n731), .B(KEYINPUT125), .Z(n732) );
  XNOR2_X1 U784 ( .A(n733), .B(n732), .ZN(n734) );
  NOR2_X1 U785 ( .A1(n739), .A2(n734), .ZN(G63) );
  NAND2_X1 U786 ( .A1(n735), .A2(G217), .ZN(n736) );
  XNOR2_X1 U787 ( .A(n737), .B(n736), .ZN(n738) );
  NOR2_X1 U788 ( .A1(n739), .A2(n738), .ZN(G66) );
  OR2_X1 U789 ( .A1(G898), .A2(n754), .ZN(n741) );
  NAND2_X1 U790 ( .A1(n741), .A2(n740), .ZN(n742) );
  XNOR2_X1 U791 ( .A(n742), .B(KEYINPUT126), .ZN(n749) );
  NAND2_X1 U792 ( .A1(G953), .A2(G224), .ZN(n743) );
  XNOR2_X1 U793 ( .A(KEYINPUT61), .B(n743), .ZN(n744) );
  NAND2_X1 U794 ( .A1(n744), .A2(G898), .ZN(n747) );
  NAND2_X1 U795 ( .A1(n745), .A2(n754), .ZN(n746) );
  NAND2_X1 U796 ( .A1(n747), .A2(n746), .ZN(n748) );
  XOR2_X1 U797 ( .A(n749), .B(n748), .Z(G69) );
  XNOR2_X1 U798 ( .A(n750), .B(KEYINPUT127), .ZN(n751) );
  XNOR2_X1 U799 ( .A(n752), .B(n751), .ZN(n756) );
  XNOR2_X1 U800 ( .A(n753), .B(n756), .ZN(n755) );
  NAND2_X1 U801 ( .A1(n755), .A2(n754), .ZN(n760) );
  XNOR2_X1 U802 ( .A(n756), .B(G227), .ZN(n757) );
  NAND2_X1 U803 ( .A1(n757), .A2(G900), .ZN(n758) );
  NAND2_X1 U804 ( .A1(G953), .A2(n758), .ZN(n759) );
  NAND2_X1 U805 ( .A1(n760), .A2(n759), .ZN(G72) );
  XOR2_X1 U806 ( .A(G134), .B(n761), .Z(G36) );
  XOR2_X1 U807 ( .A(n567), .B(G122), .Z(G24) );
  XNOR2_X1 U808 ( .A(G119), .B(n762), .ZN(G21) );
endmodule

