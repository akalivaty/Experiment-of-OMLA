//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 0 1 1 0 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 1 0 1 1 1 1 1 1 1 0 0 0 1 1 1 0 0 1 0 1 1 0 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:25:44 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n617, new_n618, new_n619, new_n620, new_n621, new_n622,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n631, new_n632, new_n633, new_n634, new_n635, new_n636, new_n637,
    new_n638, new_n639, new_n640, new_n641, new_n642, new_n644, new_n645,
    new_n646, new_n647, new_n648, new_n649, new_n650, new_n651, new_n652,
    new_n653, new_n654, new_n655, new_n656, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n708, new_n709, new_n710, new_n712, new_n713, new_n714,
    new_n715, new_n716, new_n717, new_n718, new_n720, new_n721, new_n722,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n744, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n774, new_n775,
    new_n776, new_n777, new_n778, new_n779, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n890, new_n891,
    new_n892, new_n894, new_n895, new_n896, new_n897, new_n898, new_n899,
    new_n900, new_n901, new_n902, new_n903, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n917, new_n918, new_n919, new_n920, new_n921, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n946, new_n947, new_n948, new_n949, new_n950, new_n951, new_n952,
    new_n953, new_n954, new_n955, new_n956;
  INV_X1    g000(.A(KEYINPUT69), .ZN(new_n187));
  OR2_X1    g001(.A1(KEYINPUT65), .A2(G116), .ZN(new_n188));
  NAND2_X1  g002(.A1(KEYINPUT65), .A2(G116), .ZN(new_n189));
  NAND3_X1  g003(.A1(new_n188), .A2(G119), .A3(new_n189), .ZN(new_n190));
  INV_X1    g004(.A(G116), .ZN(new_n191));
  OAI21_X1  g005(.A(new_n190), .B1(new_n191), .B2(G119), .ZN(new_n192));
  XNOR2_X1  g006(.A(KEYINPUT2), .B(G113), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n192), .A2(new_n193), .ZN(new_n194));
  INV_X1    g008(.A(new_n193), .ZN(new_n195));
  OAI211_X1 g009(.A(new_n195), .B(new_n190), .C1(new_n191), .C2(G119), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n194), .A2(new_n196), .ZN(new_n197));
  INV_X1    g011(.A(KEYINPUT30), .ZN(new_n198));
  INV_X1    g012(.A(KEYINPUT66), .ZN(new_n199));
  INV_X1    g013(.A(KEYINPUT64), .ZN(new_n200));
  INV_X1    g014(.A(G143), .ZN(new_n201));
  OAI21_X1  g015(.A(new_n200), .B1(new_n201), .B2(G146), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n201), .A2(G146), .ZN(new_n203));
  INV_X1    g017(.A(G146), .ZN(new_n204));
  NAND3_X1  g018(.A1(new_n204), .A2(KEYINPUT64), .A3(G143), .ZN(new_n205));
  NAND3_X1  g019(.A1(new_n202), .A2(new_n203), .A3(new_n205), .ZN(new_n206));
  AND2_X1   g020(.A1(KEYINPUT0), .A2(G128), .ZN(new_n207));
  NOR2_X1   g021(.A1(KEYINPUT0), .A2(G128), .ZN(new_n208));
  NOR2_X1   g022(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  AND2_X1   g023(.A1(new_n206), .A2(new_n209), .ZN(new_n210));
  XNOR2_X1  g024(.A(G143), .B(G146), .ZN(new_n211));
  AND2_X1   g025(.A1(new_n211), .A2(new_n207), .ZN(new_n212));
  OAI21_X1  g026(.A(new_n199), .B1(new_n210), .B2(new_n212), .ZN(new_n213));
  INV_X1    g027(.A(KEYINPUT11), .ZN(new_n214));
  INV_X1    g028(.A(G134), .ZN(new_n215));
  OAI21_X1  g029(.A(new_n214), .B1(new_n215), .B2(G137), .ZN(new_n216));
  INV_X1    g030(.A(G137), .ZN(new_n217));
  NAND3_X1  g031(.A1(new_n217), .A2(KEYINPUT11), .A3(G134), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n215), .A2(G137), .ZN(new_n219));
  NAND3_X1  g033(.A1(new_n216), .A2(new_n218), .A3(new_n219), .ZN(new_n220));
  OR2_X1    g034(.A1(new_n220), .A2(G131), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n220), .A2(G131), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  AOI22_X1  g037(.A1(new_n206), .A2(new_n209), .B1(new_n211), .B2(new_n207), .ZN(new_n224));
  NAND2_X1  g038(.A1(new_n224), .A2(KEYINPUT66), .ZN(new_n225));
  NAND3_X1  g039(.A1(new_n213), .A2(new_n223), .A3(new_n225), .ZN(new_n226));
  NOR2_X1   g040(.A1(new_n201), .A2(G146), .ZN(new_n227));
  INV_X1    g041(.A(KEYINPUT1), .ZN(new_n228));
  OAI21_X1  g042(.A(G128), .B1(new_n227), .B2(new_n228), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n206), .A2(new_n229), .ZN(new_n230));
  NAND3_X1  g044(.A1(new_n211), .A2(new_n228), .A3(G128), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n230), .A2(new_n231), .ZN(new_n232));
  INV_X1    g046(.A(new_n219), .ZN(new_n233));
  NOR2_X1   g047(.A1(new_n215), .A2(G137), .ZN(new_n234));
  OAI21_X1  g048(.A(G131), .B1(new_n233), .B2(new_n234), .ZN(new_n235));
  NAND3_X1  g049(.A1(new_n232), .A2(new_n221), .A3(new_n235), .ZN(new_n236));
  AOI21_X1  g050(.A(new_n198), .B1(new_n226), .B2(new_n236), .ZN(new_n237));
  INV_X1    g051(.A(new_n222), .ZN(new_n238));
  NOR2_X1   g052(.A1(new_n220), .A2(G131), .ZN(new_n239));
  OAI21_X1  g053(.A(new_n224), .B1(new_n238), .B2(new_n239), .ZN(new_n240));
  AND3_X1   g054(.A1(new_n236), .A2(new_n240), .A3(new_n198), .ZN(new_n241));
  OAI21_X1  g055(.A(new_n197), .B1(new_n237), .B2(new_n241), .ZN(new_n242));
  NAND4_X1  g056(.A1(new_n226), .A2(new_n194), .A3(new_n196), .A4(new_n236), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n242), .A2(new_n243), .ZN(new_n244));
  INV_X1    g058(.A(new_n244), .ZN(new_n245));
  AND2_X1   g059(.A1(KEYINPUT68), .A2(G953), .ZN(new_n246));
  NOR2_X1   g060(.A1(KEYINPUT68), .A2(G953), .ZN(new_n247));
  NOR2_X1   g061(.A1(new_n246), .A2(new_n247), .ZN(new_n248));
  XNOR2_X1  g062(.A(KEYINPUT67), .B(G237), .ZN(new_n249));
  NAND3_X1  g063(.A1(new_n248), .A2(new_n249), .A3(G210), .ZN(new_n250));
  XNOR2_X1  g064(.A(new_n250), .B(KEYINPUT27), .ZN(new_n251));
  XNOR2_X1  g065(.A(KEYINPUT26), .B(G101), .ZN(new_n252));
  XNOR2_X1  g066(.A(new_n251), .B(new_n252), .ZN(new_n253));
  OAI21_X1  g067(.A(new_n187), .B1(new_n245), .B2(new_n253), .ZN(new_n254));
  INV_X1    g068(.A(KEYINPUT29), .ZN(new_n255));
  INV_X1    g069(.A(new_n253), .ZN(new_n256));
  NAND3_X1  g070(.A1(new_n244), .A2(KEYINPUT69), .A3(new_n256), .ZN(new_n257));
  INV_X1    g071(.A(KEYINPUT28), .ZN(new_n258));
  AND2_X1   g072(.A1(new_n243), .A2(new_n258), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n236), .A2(new_n240), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n260), .A2(new_n197), .ZN(new_n261));
  AOI21_X1  g075(.A(new_n258), .B1(new_n243), .B2(new_n261), .ZN(new_n262));
  OR3_X1    g076(.A1(new_n259), .A2(new_n262), .A3(new_n256), .ZN(new_n263));
  NAND4_X1  g077(.A1(new_n254), .A2(new_n255), .A3(new_n257), .A4(new_n263), .ZN(new_n264));
  INV_X1    g078(.A(G902), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n226), .A2(new_n236), .ZN(new_n266));
  NAND2_X1  g080(.A1(new_n266), .A2(new_n197), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n267), .A2(new_n243), .ZN(new_n268));
  AOI21_X1  g082(.A(new_n259), .B1(new_n268), .B2(KEYINPUT28), .ZN(new_n269));
  NOR2_X1   g083(.A1(new_n256), .A2(new_n255), .ZN(new_n270));
  NAND2_X1  g084(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n271), .A2(KEYINPUT70), .ZN(new_n272));
  INV_X1    g086(.A(KEYINPUT70), .ZN(new_n273));
  NAND3_X1  g087(.A1(new_n269), .A2(new_n273), .A3(new_n270), .ZN(new_n274));
  NAND4_X1  g088(.A1(new_n264), .A2(new_n265), .A3(new_n272), .A4(new_n274), .ZN(new_n275));
  NAND3_X1  g089(.A1(new_n242), .A2(new_n243), .A3(new_n253), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n276), .A2(KEYINPUT31), .ZN(new_n277));
  INV_X1    g091(.A(KEYINPUT31), .ZN(new_n278));
  NAND4_X1  g092(.A1(new_n242), .A2(new_n278), .A3(new_n243), .A4(new_n253), .ZN(new_n279));
  OAI21_X1  g093(.A(new_n256), .B1(new_n259), .B2(new_n262), .ZN(new_n280));
  NAND3_X1  g094(.A1(new_n277), .A2(new_n279), .A3(new_n280), .ZN(new_n281));
  INV_X1    g095(.A(G472), .ZN(new_n282));
  NAND3_X1  g096(.A1(new_n281), .A2(new_n282), .A3(new_n265), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n283), .A2(KEYINPUT32), .ZN(new_n284));
  INV_X1    g098(.A(KEYINPUT32), .ZN(new_n285));
  NAND4_X1  g099(.A1(new_n281), .A2(new_n285), .A3(new_n282), .A4(new_n265), .ZN(new_n286));
  AOI22_X1  g100(.A1(new_n275), .A2(G472), .B1(new_n284), .B2(new_n286), .ZN(new_n287));
  INV_X1    g101(.A(G128), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n288), .A2(G119), .ZN(new_n289));
  INV_X1    g103(.A(G119), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n290), .A2(G128), .ZN(new_n291));
  INV_X1    g105(.A(KEYINPUT72), .ZN(new_n292));
  AND3_X1   g106(.A1(new_n289), .A2(new_n291), .A3(new_n292), .ZN(new_n293));
  AOI21_X1  g107(.A(new_n292), .B1(new_n289), .B2(new_n291), .ZN(new_n294));
  XNOR2_X1  g108(.A(KEYINPUT24), .B(G110), .ZN(new_n295));
  NOR3_X1   g109(.A1(new_n293), .A2(new_n294), .A3(new_n295), .ZN(new_n296));
  INV_X1    g110(.A(KEYINPUT23), .ZN(new_n297));
  OAI21_X1  g111(.A(new_n297), .B1(new_n290), .B2(G128), .ZN(new_n298));
  NAND3_X1  g112(.A1(new_n288), .A2(KEYINPUT23), .A3(G119), .ZN(new_n299));
  NAND3_X1  g113(.A1(new_n298), .A2(new_n291), .A3(new_n299), .ZN(new_n300));
  AOI21_X1  g114(.A(new_n296), .B1(G110), .B2(new_n300), .ZN(new_n301));
  XNOR2_X1  g115(.A(KEYINPUT74), .B(G125), .ZN(new_n302));
  NOR2_X1   g116(.A1(KEYINPUT16), .A2(G140), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n302), .A2(new_n303), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n304), .A2(KEYINPUT75), .ZN(new_n305));
  INV_X1    g119(.A(KEYINPUT75), .ZN(new_n306));
  NAND3_X1  g120(.A1(new_n302), .A2(new_n306), .A3(new_n303), .ZN(new_n307));
  AND2_X1   g121(.A1(new_n305), .A2(new_n307), .ZN(new_n308));
  INV_X1    g122(.A(KEYINPUT73), .ZN(new_n309));
  INV_X1    g123(.A(G125), .ZN(new_n310));
  OAI21_X1  g124(.A(new_n309), .B1(new_n310), .B2(G140), .ZN(new_n311));
  INV_X1    g125(.A(G140), .ZN(new_n312));
  NAND3_X1  g126(.A1(new_n312), .A2(KEYINPUT73), .A3(G125), .ZN(new_n313));
  NAND2_X1  g127(.A1(new_n311), .A2(new_n313), .ZN(new_n314));
  OAI211_X1 g128(.A(new_n314), .B(KEYINPUT16), .C1(new_n312), .C2(new_n302), .ZN(new_n315));
  AOI21_X1  g129(.A(G146), .B1(new_n308), .B2(new_n315), .ZN(new_n316));
  NAND4_X1  g130(.A1(new_n315), .A2(new_n305), .A3(G146), .A4(new_n307), .ZN(new_n317));
  INV_X1    g131(.A(new_n317), .ZN(new_n318));
  OAI21_X1  g132(.A(new_n301), .B1(new_n316), .B2(new_n318), .ZN(new_n319));
  INV_X1    g133(.A(G110), .ZN(new_n320));
  NAND4_X1  g134(.A1(new_n298), .A2(new_n299), .A3(new_n320), .A4(new_n291), .ZN(new_n321));
  OR2_X1    g135(.A1(new_n321), .A2(KEYINPUT76), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n321), .A2(KEYINPUT76), .ZN(new_n323));
  OAI21_X1  g137(.A(new_n295), .B1(new_n293), .B2(new_n294), .ZN(new_n324));
  NAND3_X1  g138(.A1(new_n322), .A2(new_n323), .A3(new_n324), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n325), .A2(KEYINPUT77), .ZN(new_n326));
  INV_X1    g140(.A(KEYINPUT77), .ZN(new_n327));
  NAND4_X1  g141(.A1(new_n322), .A2(new_n327), .A3(new_n324), .A4(new_n323), .ZN(new_n328));
  XNOR2_X1  g142(.A(G125), .B(G140), .ZN(new_n329));
  XNOR2_X1  g143(.A(new_n329), .B(KEYINPUT78), .ZN(new_n330));
  OR2_X1    g144(.A1(new_n330), .A2(G146), .ZN(new_n331));
  NAND4_X1  g145(.A1(new_n326), .A2(new_n317), .A3(new_n328), .A4(new_n331), .ZN(new_n332));
  NAND3_X1  g146(.A1(new_n248), .A2(G221), .A3(G234), .ZN(new_n333));
  XOR2_X1   g147(.A(KEYINPUT22), .B(G137), .Z(new_n334));
  XNOR2_X1  g148(.A(new_n333), .B(new_n334), .ZN(new_n335));
  AND3_X1   g149(.A1(new_n319), .A2(new_n332), .A3(new_n335), .ZN(new_n336));
  AOI21_X1  g150(.A(new_n335), .B1(new_n319), .B2(new_n332), .ZN(new_n337));
  OAI21_X1  g151(.A(new_n265), .B1(new_n336), .B2(new_n337), .ZN(new_n338));
  INV_X1    g152(.A(G217), .ZN(new_n339));
  AOI21_X1  g153(.A(new_n339), .B1(G234), .B2(new_n265), .ZN(new_n340));
  OR2_X1    g154(.A1(new_n338), .A2(new_n340), .ZN(new_n341));
  XNOR2_X1  g155(.A(new_n341), .B(KEYINPUT80), .ZN(new_n342));
  INV_X1    g156(.A(KEYINPUT79), .ZN(new_n343));
  INV_X1    g157(.A(KEYINPUT25), .ZN(new_n344));
  NOR2_X1   g158(.A1(new_n343), .A2(new_n344), .ZN(new_n345));
  NOR2_X1   g159(.A1(KEYINPUT79), .A2(KEYINPUT25), .ZN(new_n346));
  INV_X1    g160(.A(new_n346), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n338), .A2(new_n347), .ZN(new_n348));
  OAI211_X1 g162(.A(new_n265), .B(new_n346), .C1(new_n336), .C2(new_n337), .ZN(new_n349));
  AOI21_X1  g163(.A(new_n345), .B1(new_n348), .B2(new_n349), .ZN(new_n350));
  XOR2_X1   g164(.A(new_n340), .B(KEYINPUT71), .Z(new_n351));
  OR2_X1    g165(.A1(new_n350), .A2(new_n351), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n342), .A2(new_n352), .ZN(new_n353));
  NOR2_X1   g167(.A1(new_n287), .A2(new_n353), .ZN(new_n354));
  OAI21_X1  g168(.A(G214), .B1(G237), .B2(G902), .ZN(new_n355));
  INV_X1    g169(.A(new_n355), .ZN(new_n356));
  XNOR2_X1  g170(.A(G110), .B(G122), .ZN(new_n357));
  XNOR2_X1  g171(.A(new_n357), .B(KEYINPUT82), .ZN(new_n358));
  XNOR2_X1  g172(.A(new_n358), .B(KEYINPUT8), .ZN(new_n359));
  INV_X1    g173(.A(G113), .ZN(new_n360));
  NOR3_X1   g174(.A1(new_n191), .A2(KEYINPUT5), .A3(G119), .ZN(new_n361));
  AOI21_X1  g175(.A(new_n360), .B1(new_n361), .B2(KEYINPUT81), .ZN(new_n362));
  INV_X1    g176(.A(KEYINPUT5), .ZN(new_n363));
  OAI221_X1 g177(.A(new_n362), .B1(KEYINPUT81), .B2(new_n361), .C1(new_n192), .C2(new_n363), .ZN(new_n364));
  INV_X1    g178(.A(G104), .ZN(new_n365));
  OAI21_X1  g179(.A(KEYINPUT3), .B1(new_n365), .B2(G107), .ZN(new_n366));
  INV_X1    g180(.A(KEYINPUT3), .ZN(new_n367));
  INV_X1    g181(.A(G107), .ZN(new_n368));
  NAND3_X1  g182(.A1(new_n367), .A2(new_n368), .A3(G104), .ZN(new_n369));
  INV_X1    g183(.A(G101), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n365), .A2(G107), .ZN(new_n371));
  NAND4_X1  g185(.A1(new_n366), .A2(new_n369), .A3(new_n370), .A4(new_n371), .ZN(new_n372));
  NOR2_X1   g186(.A1(new_n365), .A2(G107), .ZN(new_n373));
  NOR2_X1   g187(.A1(new_n368), .A2(G104), .ZN(new_n374));
  OAI21_X1  g188(.A(G101), .B1(new_n373), .B2(new_n374), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n372), .A2(new_n375), .ZN(new_n376));
  INV_X1    g190(.A(new_n376), .ZN(new_n377));
  NAND3_X1  g191(.A1(new_n364), .A2(new_n196), .A3(new_n377), .ZN(new_n378));
  INV_X1    g192(.A(new_n378), .ZN(new_n379));
  AOI21_X1  g193(.A(new_n377), .B1(new_n364), .B2(new_n196), .ZN(new_n380));
  OAI21_X1  g194(.A(new_n359), .B1(new_n379), .B2(new_n380), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n381), .A2(KEYINPUT83), .ZN(new_n382));
  INV_X1    g196(.A(new_n302), .ZN(new_n383));
  NAND2_X1  g197(.A1(new_n232), .A2(new_n383), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n224), .A2(new_n302), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n384), .A2(new_n385), .ZN(new_n386));
  INV_X1    g200(.A(G224), .ZN(new_n387));
  NOR2_X1   g201(.A1(new_n387), .A2(G953), .ZN(new_n388));
  INV_X1    g202(.A(KEYINPUT7), .ZN(new_n389));
  NOR2_X1   g203(.A1(new_n388), .A2(new_n389), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n386), .A2(new_n390), .ZN(new_n391));
  XNOR2_X1  g205(.A(new_n391), .B(KEYINPUT84), .ZN(new_n392));
  NAND3_X1  g206(.A1(new_n366), .A2(new_n369), .A3(new_n371), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n393), .A2(G101), .ZN(new_n394));
  OR2_X1    g208(.A1(new_n394), .A2(KEYINPUT4), .ZN(new_n395));
  NAND3_X1  g209(.A1(new_n394), .A2(KEYINPUT4), .A3(new_n372), .ZN(new_n396));
  NAND3_X1  g210(.A1(new_n197), .A2(new_n395), .A3(new_n396), .ZN(new_n397));
  NAND3_X1  g211(.A1(new_n378), .A2(new_n358), .A3(new_n397), .ZN(new_n398));
  OR2_X1    g212(.A1(new_n386), .A2(new_n390), .ZN(new_n399));
  AND2_X1   g213(.A1(new_n398), .A2(new_n399), .ZN(new_n400));
  INV_X1    g214(.A(KEYINPUT83), .ZN(new_n401));
  OAI211_X1 g215(.A(new_n401), .B(new_n359), .C1(new_n379), .C2(new_n380), .ZN(new_n402));
  NAND4_X1  g216(.A1(new_n382), .A2(new_n392), .A3(new_n400), .A4(new_n402), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n378), .A2(new_n397), .ZN(new_n404));
  INV_X1    g218(.A(new_n358), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n404), .A2(new_n405), .ZN(new_n406));
  NAND3_X1  g220(.A1(new_n406), .A2(KEYINPUT6), .A3(new_n398), .ZN(new_n407));
  INV_X1    g221(.A(KEYINPUT6), .ZN(new_n408));
  NAND3_X1  g222(.A1(new_n404), .A2(new_n408), .A3(new_n405), .ZN(new_n409));
  XOR2_X1   g223(.A(new_n386), .B(new_n388), .Z(new_n410));
  NAND3_X1  g224(.A1(new_n407), .A2(new_n409), .A3(new_n410), .ZN(new_n411));
  NAND3_X1  g225(.A1(new_n403), .A2(new_n265), .A3(new_n411), .ZN(new_n412));
  OAI21_X1  g226(.A(G210), .B1(G237), .B2(G902), .ZN(new_n413));
  XOR2_X1   g227(.A(new_n413), .B(KEYINPUT85), .Z(new_n414));
  NAND2_X1  g228(.A1(new_n412), .A2(new_n414), .ZN(new_n415));
  INV_X1    g229(.A(new_n414), .ZN(new_n416));
  NAND4_X1  g230(.A1(new_n403), .A2(new_n411), .A3(new_n265), .A4(new_n416), .ZN(new_n417));
  AOI21_X1  g231(.A(new_n356), .B1(new_n415), .B2(new_n417), .ZN(new_n418));
  INV_X1    g232(.A(new_n418), .ZN(new_n419));
  NAND2_X1  g233(.A1(new_n248), .A2(G227), .ZN(new_n420));
  XNOR2_X1  g234(.A(G110), .B(G140), .ZN(new_n421));
  XNOR2_X1  g235(.A(new_n420), .B(new_n421), .ZN(new_n422));
  INV_X1    g236(.A(new_n422), .ZN(new_n423));
  INV_X1    g237(.A(KEYINPUT10), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n204), .A2(G143), .ZN(new_n425));
  AOI21_X1  g239(.A(new_n288), .B1(new_n425), .B2(KEYINPUT1), .ZN(new_n426));
  NOR2_X1   g240(.A1(new_n426), .A2(new_n211), .ZN(new_n427));
  AND4_X1   g241(.A1(new_n228), .A2(new_n425), .A3(new_n203), .A4(G128), .ZN(new_n428));
  OAI211_X1 g242(.A(new_n372), .B(new_n375), .C1(new_n427), .C2(new_n428), .ZN(new_n429));
  AOI21_X1  g243(.A(new_n424), .B1(new_n230), .B2(new_n231), .ZN(new_n430));
  AOI22_X1  g244(.A1(new_n424), .A2(new_n429), .B1(new_n430), .B2(new_n377), .ZN(new_n431));
  NAND4_X1  g245(.A1(new_n213), .A2(new_n395), .A3(new_n225), .A4(new_n396), .ZN(new_n432));
  INV_X1    g246(.A(new_n223), .ZN(new_n433));
  AND3_X1   g247(.A1(new_n431), .A2(new_n432), .A3(new_n433), .ZN(new_n434));
  AOI21_X1  g248(.A(new_n433), .B1(new_n431), .B2(new_n432), .ZN(new_n435));
  OAI21_X1  g249(.A(new_n423), .B1(new_n434), .B2(new_n435), .ZN(new_n436));
  NAND3_X1  g250(.A1(new_n431), .A2(new_n432), .A3(new_n433), .ZN(new_n437));
  OAI21_X1  g251(.A(new_n429), .B1(new_n232), .B2(new_n377), .ZN(new_n438));
  AND3_X1   g252(.A1(new_n438), .A2(KEYINPUT12), .A3(new_n223), .ZN(new_n439));
  AOI21_X1  g253(.A(KEYINPUT12), .B1(new_n438), .B2(new_n223), .ZN(new_n440));
  OAI211_X1 g254(.A(new_n437), .B(new_n422), .C1(new_n439), .C2(new_n440), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n436), .A2(new_n441), .ZN(new_n442));
  INV_X1    g256(.A(G469), .ZN(new_n443));
  NAND3_X1  g257(.A1(new_n442), .A2(new_n443), .A3(new_n265), .ZN(new_n444));
  OAI21_X1  g258(.A(new_n437), .B1(new_n439), .B2(new_n440), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n445), .A2(new_n423), .ZN(new_n446));
  INV_X1    g260(.A(new_n435), .ZN(new_n447));
  NAND3_X1  g261(.A1(new_n447), .A2(new_n437), .A3(new_n422), .ZN(new_n448));
  AOI21_X1  g262(.A(G902), .B1(new_n446), .B2(new_n448), .ZN(new_n449));
  OAI21_X1  g263(.A(new_n444), .B1(new_n449), .B2(new_n443), .ZN(new_n450));
  XNOR2_X1  g264(.A(KEYINPUT9), .B(G234), .ZN(new_n451));
  OAI21_X1  g265(.A(G221), .B1(new_n451), .B2(G902), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n450), .A2(new_n452), .ZN(new_n453));
  NOR2_X1   g267(.A1(new_n419), .A2(new_n453), .ZN(new_n454));
  XNOR2_X1  g268(.A(G113), .B(G122), .ZN(new_n455));
  XNOR2_X1  g269(.A(new_n455), .B(new_n365), .ZN(new_n456));
  NAND3_X1  g270(.A1(new_n248), .A2(new_n249), .A3(G214), .ZN(new_n457));
  NOR2_X1   g271(.A1(new_n457), .A2(new_n201), .ZN(new_n458));
  INV_X1    g272(.A(new_n458), .ZN(new_n459));
  AND3_X1   g273(.A1(new_n457), .A2(KEYINPUT86), .A3(new_n201), .ZN(new_n460));
  AOI21_X1  g274(.A(KEYINPUT86), .B1(new_n457), .B2(new_n201), .ZN(new_n461));
  OAI21_X1  g275(.A(new_n459), .B1(new_n460), .B2(new_n461), .ZN(new_n462));
  NAND3_X1  g276(.A1(new_n462), .A2(KEYINPUT18), .A3(G131), .ZN(new_n463));
  AOI22_X1  g277(.A1(new_n383), .A2(G140), .B1(new_n311), .B2(new_n313), .ZN(new_n464));
  OAI21_X1  g278(.A(new_n331), .B1(new_n204), .B2(new_n464), .ZN(new_n465));
  AND2_X1   g279(.A1(KEYINPUT18), .A2(G131), .ZN(new_n466));
  OAI211_X1 g280(.A(new_n463), .B(new_n465), .C1(new_n462), .C2(new_n466), .ZN(new_n467));
  INV_X1    g281(.A(KEYINPUT68), .ZN(new_n468));
  INV_X1    g282(.A(G953), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  NAND2_X1  g284(.A1(KEYINPUT68), .A2(G953), .ZN(new_n471));
  AND2_X1   g285(.A1(KEYINPUT67), .A2(G237), .ZN(new_n472));
  NOR2_X1   g286(.A1(KEYINPUT67), .A2(G237), .ZN(new_n473));
  OAI211_X1 g287(.A(new_n470), .B(new_n471), .C1(new_n472), .C2(new_n473), .ZN(new_n474));
  INV_X1    g288(.A(G214), .ZN(new_n475));
  OAI21_X1  g289(.A(new_n201), .B1(new_n474), .B2(new_n475), .ZN(new_n476));
  INV_X1    g290(.A(KEYINPUT86), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  NAND3_X1  g292(.A1(new_n457), .A2(KEYINPUT86), .A3(new_n201), .ZN(new_n479));
  AOI211_X1 g293(.A(G131), .B(new_n458), .C1(new_n478), .C2(new_n479), .ZN(new_n480));
  AOI21_X1  g294(.A(new_n458), .B1(new_n478), .B2(new_n479), .ZN(new_n481));
  INV_X1    g295(.A(G131), .ZN(new_n482));
  OAI21_X1  g296(.A(KEYINPUT87), .B1(new_n481), .B2(new_n482), .ZN(new_n483));
  INV_X1    g297(.A(KEYINPUT87), .ZN(new_n484));
  NAND3_X1  g298(.A1(new_n462), .A2(new_n484), .A3(G131), .ZN(new_n485));
  AOI211_X1 g299(.A(KEYINPUT17), .B(new_n480), .C1(new_n483), .C2(new_n485), .ZN(new_n486));
  NAND3_X1  g300(.A1(new_n483), .A2(KEYINPUT17), .A3(new_n485), .ZN(new_n487));
  NOR2_X1   g301(.A1(new_n316), .A2(new_n318), .ZN(new_n488));
  NAND2_X1  g302(.A1(new_n487), .A2(new_n488), .ZN(new_n489));
  OAI211_X1 g303(.A(new_n456), .B(new_n467), .C1(new_n486), .C2(new_n489), .ZN(new_n490));
  NAND2_X1  g304(.A1(new_n490), .A2(KEYINPUT89), .ZN(new_n491));
  INV_X1    g305(.A(new_n480), .ZN(new_n492));
  NOR3_X1   g306(.A1(new_n481), .A2(KEYINPUT87), .A3(new_n482), .ZN(new_n493));
  AOI21_X1  g307(.A(new_n484), .B1(new_n462), .B2(G131), .ZN(new_n494));
  OAI21_X1  g308(.A(new_n492), .B1(new_n493), .B2(new_n494), .ZN(new_n495));
  OAI211_X1 g309(.A(new_n488), .B(new_n487), .C1(new_n495), .C2(KEYINPUT17), .ZN(new_n496));
  INV_X1    g310(.A(KEYINPUT89), .ZN(new_n497));
  NAND4_X1  g311(.A1(new_n496), .A2(new_n497), .A3(new_n456), .A4(new_n467), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n491), .A2(new_n498), .ZN(new_n499));
  INV_X1    g313(.A(KEYINPUT19), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n330), .A2(new_n500), .ZN(new_n501));
  NAND2_X1  g315(.A1(new_n464), .A2(KEYINPUT19), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  AOI21_X1  g317(.A(new_n318), .B1(new_n503), .B2(new_n204), .ZN(new_n504));
  INV_X1    g318(.A(KEYINPUT88), .ZN(new_n505));
  OR2_X1    g319(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  NAND2_X1  g320(.A1(new_n504), .A2(new_n505), .ZN(new_n507));
  NAND3_X1  g321(.A1(new_n495), .A2(new_n506), .A3(new_n507), .ZN(new_n508));
  AOI21_X1  g322(.A(new_n456), .B1(new_n508), .B2(new_n467), .ZN(new_n509));
  INV_X1    g323(.A(new_n509), .ZN(new_n510));
  NAND2_X1  g324(.A1(new_n499), .A2(new_n510), .ZN(new_n511));
  NOR2_X1   g325(.A1(G475), .A2(G902), .ZN(new_n512));
  INV_X1    g326(.A(new_n512), .ZN(new_n513));
  NOR2_X1   g327(.A1(new_n513), .A2(KEYINPUT20), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n511), .A2(new_n514), .ZN(new_n515));
  INV_X1    g329(.A(new_n515), .ZN(new_n516));
  INV_X1    g330(.A(KEYINPUT90), .ZN(new_n517));
  NAND2_X1  g331(.A1(new_n511), .A2(new_n517), .ZN(new_n518));
  NAND3_X1  g332(.A1(new_n499), .A2(KEYINPUT90), .A3(new_n510), .ZN(new_n519));
  NAND3_X1  g333(.A1(new_n518), .A2(new_n512), .A3(new_n519), .ZN(new_n520));
  AOI21_X1  g334(.A(new_n516), .B1(new_n520), .B2(KEYINPUT20), .ZN(new_n521));
  INV_X1    g335(.A(new_n499), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n496), .A2(new_n467), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n523), .A2(KEYINPUT92), .ZN(new_n524));
  INV_X1    g338(.A(KEYINPUT92), .ZN(new_n525));
  NAND3_X1  g339(.A1(new_n496), .A2(new_n525), .A3(new_n467), .ZN(new_n526));
  AOI21_X1  g340(.A(new_n456), .B1(new_n524), .B2(new_n526), .ZN(new_n527));
  OAI21_X1  g341(.A(new_n265), .B1(new_n522), .B2(new_n527), .ZN(new_n528));
  XNOR2_X1  g342(.A(KEYINPUT91), .B(G475), .ZN(new_n529));
  NAND2_X1  g343(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  INV_X1    g344(.A(new_n530), .ZN(new_n531));
  NOR2_X1   g345(.A1(new_n521), .A2(new_n531), .ZN(new_n532));
  NAND3_X1  g346(.A1(new_n188), .A2(G122), .A3(new_n189), .ZN(new_n533));
  INV_X1    g347(.A(KEYINPUT94), .ZN(new_n534));
  OR2_X1    g348(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n533), .A2(new_n534), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  NOR2_X1   g351(.A1(new_n191), .A2(G122), .ZN(new_n538));
  XOR2_X1   g352(.A(new_n538), .B(KEYINPUT93), .Z(new_n539));
  NAND2_X1  g353(.A1(new_n537), .A2(new_n539), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n540), .A2(G107), .ZN(new_n541));
  NAND3_X1  g355(.A1(new_n537), .A2(new_n368), .A3(new_n539), .ZN(new_n542));
  NAND2_X1  g356(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  OAI21_X1  g357(.A(KEYINPUT95), .B1(new_n201), .B2(G128), .ZN(new_n544));
  INV_X1    g358(.A(KEYINPUT95), .ZN(new_n545));
  NAND3_X1  g359(.A1(new_n545), .A2(new_n288), .A3(G143), .ZN(new_n546));
  AOI21_X1  g360(.A(KEYINPUT13), .B1(new_n544), .B2(new_n546), .ZN(new_n547));
  NOR2_X1   g361(.A1(new_n547), .A2(new_n215), .ZN(new_n548));
  AOI22_X1  g362(.A1(new_n544), .A2(new_n546), .B1(G128), .B2(new_n201), .ZN(new_n549));
  XNOR2_X1  g363(.A(new_n548), .B(new_n549), .ZN(new_n550));
  NAND2_X1  g364(.A1(new_n543), .A2(new_n550), .ZN(new_n551));
  XNOR2_X1  g365(.A(new_n549), .B(new_n215), .ZN(new_n552));
  AND2_X1   g366(.A1(new_n542), .A2(new_n552), .ZN(new_n553));
  INV_X1    g367(.A(KEYINPUT14), .ZN(new_n554));
  NAND3_X1  g368(.A1(new_n535), .A2(new_n554), .A3(new_n536), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n555), .A2(new_n539), .ZN(new_n556));
  AOI21_X1  g370(.A(new_n554), .B1(new_n535), .B2(new_n536), .ZN(new_n557));
  OAI21_X1  g371(.A(G107), .B1(new_n556), .B2(new_n557), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n553), .A2(new_n558), .ZN(new_n559));
  NOR3_X1   g373(.A1(new_n451), .A2(new_n339), .A3(G953), .ZN(new_n560));
  NAND3_X1  g374(.A1(new_n551), .A2(new_n559), .A3(new_n560), .ZN(new_n561));
  INV_X1    g375(.A(KEYINPUT96), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  NAND4_X1  g377(.A1(new_n551), .A2(new_n559), .A3(KEYINPUT96), .A4(new_n560), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n551), .A2(new_n559), .ZN(new_n565));
  INV_X1    g379(.A(new_n560), .ZN(new_n566));
  AOI22_X1  g380(.A1(new_n563), .A2(new_n564), .B1(new_n565), .B2(new_n566), .ZN(new_n567));
  INV_X1    g381(.A(G478), .ZN(new_n568));
  NOR2_X1   g382(.A1(new_n568), .A2(KEYINPUT15), .ZN(new_n569));
  OR3_X1    g383(.A1(new_n567), .A2(G902), .A3(new_n569), .ZN(new_n570));
  OAI21_X1  g384(.A(new_n569), .B1(new_n567), .B2(G902), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n570), .A2(new_n571), .ZN(new_n572));
  INV_X1    g386(.A(new_n572), .ZN(new_n573));
  AND2_X1   g387(.A1(new_n469), .A2(G952), .ZN(new_n574));
  NAND2_X1  g388(.A1(G234), .A2(G237), .ZN(new_n575));
  AND2_X1   g389(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  INV_X1    g390(.A(new_n248), .ZN(new_n577));
  AND3_X1   g391(.A1(new_n577), .A2(G902), .A3(new_n575), .ZN(new_n578));
  XNOR2_X1  g392(.A(KEYINPUT21), .B(G898), .ZN(new_n579));
  AOI21_X1  g393(.A(new_n576), .B1(new_n578), .B2(new_n579), .ZN(new_n580));
  INV_X1    g394(.A(new_n580), .ZN(new_n581));
  NAND2_X1  g395(.A1(new_n573), .A2(new_n581), .ZN(new_n582));
  INV_X1    g396(.A(new_n582), .ZN(new_n583));
  AOI21_X1  g397(.A(KEYINPUT97), .B1(new_n532), .B2(new_n583), .ZN(new_n584));
  AOI21_X1  g398(.A(KEYINPUT90), .B1(new_n499), .B2(new_n510), .ZN(new_n585));
  AOI211_X1 g399(.A(new_n517), .B(new_n509), .C1(new_n491), .C2(new_n498), .ZN(new_n586));
  NOR3_X1   g400(.A1(new_n585), .A2(new_n586), .A3(new_n513), .ZN(new_n587));
  INV_X1    g401(.A(KEYINPUT20), .ZN(new_n588));
  OAI21_X1  g402(.A(new_n515), .B1(new_n587), .B2(new_n588), .ZN(new_n589));
  AND4_X1   g403(.A1(KEYINPUT97), .A2(new_n589), .A3(new_n530), .A4(new_n583), .ZN(new_n590));
  OAI211_X1 g404(.A(new_n354), .B(new_n454), .C1(new_n584), .C2(new_n590), .ZN(new_n591));
  XOR2_X1   g405(.A(KEYINPUT98), .B(G101), .Z(new_n592));
  XNOR2_X1  g406(.A(new_n591), .B(new_n592), .ZN(G3));
  NAND2_X1  g407(.A1(new_n565), .A2(new_n566), .ZN(new_n594));
  XNOR2_X1  g408(.A(new_n594), .B(KEYINPUT99), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n595), .A2(new_n561), .ZN(new_n596));
  NAND2_X1  g410(.A1(new_n596), .A2(KEYINPUT33), .ZN(new_n597));
  INV_X1    g411(.A(new_n567), .ZN(new_n598));
  OAI21_X1  g412(.A(new_n597), .B1(KEYINPUT33), .B2(new_n598), .ZN(new_n599));
  NOR2_X1   g413(.A1(new_n568), .A2(G902), .ZN(new_n600));
  NAND2_X1  g414(.A1(new_n598), .A2(new_n265), .ZN(new_n601));
  AOI22_X1  g415(.A1(new_n599), .A2(new_n600), .B1(new_n568), .B2(new_n601), .ZN(new_n602));
  AOI21_X1  g416(.A(new_n602), .B1(new_n589), .B2(new_n530), .ZN(new_n603));
  INV_X1    g417(.A(new_n353), .ZN(new_n604));
  INV_X1    g418(.A(new_n453), .ZN(new_n605));
  NAND2_X1  g419(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  NAND2_X1  g420(.A1(new_n281), .A2(new_n265), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n607), .A2(G472), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n608), .A2(new_n283), .ZN(new_n609));
  NOR2_X1   g423(.A1(new_n606), .A2(new_n609), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n418), .A2(new_n581), .ZN(new_n611));
  INV_X1    g425(.A(new_n611), .ZN(new_n612));
  NAND3_X1  g426(.A1(new_n603), .A2(new_n610), .A3(new_n612), .ZN(new_n613));
  XNOR2_X1  g427(.A(new_n613), .B(KEYINPUT100), .ZN(new_n614));
  XNOR2_X1  g428(.A(new_n614), .B(KEYINPUT34), .ZN(new_n615));
  XNOR2_X1  g429(.A(new_n615), .B(new_n365), .ZN(G6));
  NOR2_X1   g430(.A1(new_n585), .A2(new_n586), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n617), .A2(new_n514), .ZN(new_n618));
  OAI21_X1  g432(.A(new_n618), .B1(new_n588), .B2(new_n587), .ZN(new_n619));
  AOI21_X1  g433(.A(new_n573), .B1(new_n528), .B2(new_n529), .ZN(new_n620));
  NAND3_X1  g434(.A1(new_n619), .A2(new_n581), .A3(new_n620), .ZN(new_n621));
  INV_X1    g435(.A(KEYINPUT101), .ZN(new_n622));
  AOI21_X1  g436(.A(new_n419), .B1(new_n621), .B2(new_n622), .ZN(new_n623));
  INV_X1    g437(.A(KEYINPUT102), .ZN(new_n624));
  NAND4_X1  g438(.A1(new_n619), .A2(KEYINPUT101), .A3(new_n581), .A4(new_n620), .ZN(new_n625));
  AND3_X1   g439(.A1(new_n623), .A2(new_n624), .A3(new_n625), .ZN(new_n626));
  AOI21_X1  g440(.A(new_n624), .B1(new_n623), .B2(new_n625), .ZN(new_n627));
  OAI21_X1  g441(.A(new_n610), .B1(new_n626), .B2(new_n627), .ZN(new_n628));
  XOR2_X1   g442(.A(KEYINPUT35), .B(G107), .Z(new_n629));
  XNOR2_X1  g443(.A(new_n628), .B(new_n629), .ZN(G9));
  NAND2_X1  g444(.A1(new_n319), .A2(new_n332), .ZN(new_n631));
  NOR2_X1   g445(.A1(new_n335), .A2(KEYINPUT36), .ZN(new_n632));
  XNOR2_X1  g446(.A(new_n631), .B(new_n632), .ZN(new_n633));
  OAI211_X1 g447(.A(new_n633), .B(new_n265), .C1(new_n339), .C2(G234), .ZN(new_n634));
  OAI21_X1  g448(.A(new_n634), .B1(new_n350), .B2(new_n351), .ZN(new_n635));
  INV_X1    g449(.A(KEYINPUT103), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n635), .A2(new_n636), .ZN(new_n637));
  OAI211_X1 g451(.A(KEYINPUT103), .B(new_n634), .C1(new_n350), .C2(new_n351), .ZN(new_n638));
  AND2_X1   g452(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  AND3_X1   g453(.A1(new_n639), .A2(new_n283), .A3(new_n608), .ZN(new_n640));
  OAI211_X1 g454(.A(new_n454), .B(new_n640), .C1(new_n584), .C2(new_n590), .ZN(new_n641));
  XOR2_X1   g455(.A(KEYINPUT37), .B(G110), .Z(new_n642));
  XNOR2_X1  g456(.A(new_n641), .B(new_n642), .ZN(G12));
  AOI22_X1  g457(.A1(new_n520), .A2(KEYINPUT20), .B1(new_n617), .B2(new_n514), .ZN(new_n644));
  NAND2_X1  g458(.A1(new_n530), .A2(new_n572), .ZN(new_n645));
  INV_X1    g459(.A(KEYINPUT104), .ZN(new_n646));
  INV_X1    g460(.A(new_n578), .ZN(new_n647));
  OAI21_X1  g461(.A(new_n646), .B1(new_n647), .B2(G900), .ZN(new_n648));
  INV_X1    g462(.A(new_n576), .ZN(new_n649));
  INV_X1    g463(.A(G900), .ZN(new_n650));
  NAND3_X1  g464(.A1(new_n578), .A2(KEYINPUT104), .A3(new_n650), .ZN(new_n651));
  AND3_X1   g465(.A1(new_n648), .A2(new_n649), .A3(new_n651), .ZN(new_n652));
  NOR3_X1   g466(.A1(new_n644), .A2(new_n645), .A3(new_n652), .ZN(new_n653));
  NAND3_X1  g467(.A1(new_n637), .A2(new_n418), .A3(new_n638), .ZN(new_n654));
  NOR3_X1   g468(.A1(new_n654), .A2(new_n287), .A3(new_n453), .ZN(new_n655));
  NAND2_X1  g469(.A1(new_n653), .A2(new_n655), .ZN(new_n656));
  XNOR2_X1  g470(.A(new_n656), .B(G128), .ZN(G30));
  XOR2_X1   g471(.A(new_n652), .B(KEYINPUT39), .Z(new_n658));
  NAND2_X1  g472(.A1(new_n605), .A2(new_n658), .ZN(new_n659));
  XOR2_X1   g473(.A(KEYINPUT107), .B(KEYINPUT40), .Z(new_n660));
  XNOR2_X1  g474(.A(new_n659), .B(new_n660), .ZN(new_n661));
  NAND2_X1  g475(.A1(new_n415), .A2(new_n417), .ZN(new_n662));
  XOR2_X1   g476(.A(new_n662), .B(KEYINPUT38), .Z(new_n663));
  INV_X1    g477(.A(new_n663), .ZN(new_n664));
  NAND2_X1  g478(.A1(new_n661), .A2(new_n664), .ZN(new_n665));
  NAND2_X1  g479(.A1(new_n284), .A2(new_n286), .ZN(new_n666));
  AOI21_X1  g480(.A(new_n253), .B1(new_n267), .B2(new_n243), .ZN(new_n667));
  INV_X1    g481(.A(KEYINPUT105), .ZN(new_n668));
  OR2_X1    g482(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  NAND2_X1  g483(.A1(new_n667), .A2(new_n668), .ZN(new_n670));
  AND3_X1   g484(.A1(new_n669), .A2(new_n276), .A3(new_n670), .ZN(new_n671));
  OAI21_X1  g485(.A(G472), .B1(new_n671), .B2(G902), .ZN(new_n672));
  NAND2_X1  g486(.A1(new_n666), .A2(new_n672), .ZN(new_n673));
  NAND2_X1  g487(.A1(new_n673), .A2(KEYINPUT106), .ZN(new_n674));
  INV_X1    g488(.A(KEYINPUT106), .ZN(new_n675));
  NAND3_X1  g489(.A1(new_n666), .A2(new_n675), .A3(new_n672), .ZN(new_n676));
  AND2_X1   g490(.A1(new_n674), .A2(new_n676), .ZN(new_n677));
  NOR4_X1   g491(.A1(new_n665), .A2(new_n677), .A3(new_n356), .A4(new_n635), .ZN(new_n678));
  NOR2_X1   g492(.A1(new_n532), .A2(new_n573), .ZN(new_n679));
  NAND2_X1  g493(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  XNOR2_X1  g494(.A(new_n680), .B(G143), .ZN(G45));
  AOI21_X1  g495(.A(new_n588), .B1(new_n617), .B2(new_n512), .ZN(new_n682));
  OAI21_X1  g496(.A(new_n530), .B1(new_n682), .B2(new_n516), .ZN(new_n683));
  INV_X1    g497(.A(new_n602), .ZN(new_n684));
  INV_X1    g498(.A(new_n652), .ZN(new_n685));
  NAND4_X1  g499(.A1(new_n683), .A2(new_n655), .A3(new_n684), .A4(new_n685), .ZN(new_n686));
  XNOR2_X1  g500(.A(new_n686), .B(G146), .ZN(G48));
  NAND3_X1  g501(.A1(new_n683), .A2(new_n684), .A3(new_n612), .ZN(new_n688));
  NAND2_X1  g502(.A1(new_n442), .A2(new_n265), .ZN(new_n689));
  NAND2_X1  g503(.A1(new_n689), .A2(G469), .ZN(new_n690));
  NAND2_X1  g504(.A1(new_n690), .A2(new_n444), .ZN(new_n691));
  INV_X1    g505(.A(new_n691), .ZN(new_n692));
  AND2_X1   g506(.A1(new_n692), .A2(new_n452), .ZN(new_n693));
  NAND2_X1  g507(.A1(new_n354), .A2(new_n693), .ZN(new_n694));
  OAI21_X1  g508(.A(KEYINPUT108), .B1(new_n688), .B2(new_n694), .ZN(new_n695));
  INV_X1    g509(.A(new_n694), .ZN(new_n696));
  INV_X1    g510(.A(KEYINPUT108), .ZN(new_n697));
  NAND4_X1  g511(.A1(new_n696), .A2(new_n603), .A3(new_n697), .A4(new_n612), .ZN(new_n698));
  NAND2_X1  g512(.A1(new_n695), .A2(new_n698), .ZN(new_n699));
  XNOR2_X1  g513(.A(KEYINPUT41), .B(G113), .ZN(new_n700));
  XNOR2_X1  g514(.A(new_n699), .B(new_n700), .ZN(G15));
  NAND2_X1  g515(.A1(new_n621), .A2(new_n622), .ZN(new_n702));
  NAND3_X1  g516(.A1(new_n702), .A2(new_n418), .A3(new_n625), .ZN(new_n703));
  NAND2_X1  g517(.A1(new_n703), .A2(KEYINPUT102), .ZN(new_n704));
  NAND3_X1  g518(.A1(new_n623), .A2(new_n624), .A3(new_n625), .ZN(new_n705));
  AOI21_X1  g519(.A(new_n694), .B1(new_n704), .B2(new_n705), .ZN(new_n706));
  XNOR2_X1  g520(.A(new_n706), .B(new_n191), .ZN(G18));
  INV_X1    g521(.A(new_n693), .ZN(new_n708));
  NOR3_X1   g522(.A1(new_n654), .A2(new_n287), .A3(new_n708), .ZN(new_n709));
  OAI21_X1  g523(.A(new_n709), .B1(new_n584), .B2(new_n590), .ZN(new_n710));
  XNOR2_X1  g524(.A(new_n710), .B(G119), .ZN(G21));
  OAI21_X1  g525(.A(new_n277), .B1(new_n253), .B2(new_n269), .ZN(new_n712));
  AND2_X1   g526(.A1(new_n712), .A2(KEYINPUT109), .ZN(new_n713));
  OAI21_X1  g527(.A(new_n279), .B1(new_n712), .B2(KEYINPUT109), .ZN(new_n714));
  OAI211_X1 g528(.A(new_n282), .B(new_n265), .C1(new_n713), .C2(new_n714), .ZN(new_n715));
  AND3_X1   g529(.A1(new_n715), .A2(new_n604), .A3(new_n608), .ZN(new_n716));
  NOR2_X1   g530(.A1(new_n708), .A2(new_n580), .ZN(new_n717));
  NAND4_X1  g531(.A1(new_n679), .A2(new_n418), .A3(new_n716), .A4(new_n717), .ZN(new_n718));
  XNOR2_X1  g532(.A(new_n718), .B(G122), .ZN(G24));
  NOR2_X1   g533(.A1(new_n708), .A2(new_n419), .ZN(new_n720));
  AND3_X1   g534(.A1(new_n715), .A2(new_n608), .A3(new_n635), .ZN(new_n721));
  NAND4_X1  g535(.A1(new_n603), .A2(new_n685), .A3(new_n720), .A4(new_n721), .ZN(new_n722));
  XNOR2_X1  g536(.A(new_n722), .B(G125), .ZN(G27));
  INV_X1    g537(.A(KEYINPUT42), .ZN(new_n724));
  OR2_X1    g538(.A1(new_n724), .A2(KEYINPUT112), .ZN(new_n725));
  NAND2_X1  g539(.A1(new_n724), .A2(KEYINPUT112), .ZN(new_n726));
  NAND3_X1  g540(.A1(new_n683), .A2(new_n684), .A3(new_n685), .ZN(new_n727));
  INV_X1    g541(.A(KEYINPUT110), .ZN(new_n728));
  NAND2_X1  g542(.A1(new_n450), .A2(new_n728), .ZN(new_n729));
  OAI211_X1 g543(.A(new_n444), .B(KEYINPUT110), .C1(new_n443), .C2(new_n449), .ZN(new_n730));
  NAND2_X1  g544(.A1(new_n729), .A2(new_n730), .ZN(new_n731));
  NAND4_X1  g545(.A1(new_n415), .A2(new_n452), .A3(new_n355), .A4(new_n417), .ZN(new_n732));
  INV_X1    g546(.A(KEYINPUT111), .ZN(new_n733));
  OR3_X1    g547(.A1(new_n731), .A2(new_n732), .A3(new_n733), .ZN(new_n734));
  OAI21_X1  g548(.A(new_n733), .B1(new_n731), .B2(new_n732), .ZN(new_n735));
  NAND2_X1  g549(.A1(new_n734), .A2(new_n735), .ZN(new_n736));
  NAND2_X1  g550(.A1(new_n736), .A2(new_n354), .ZN(new_n737));
  OAI211_X1 g551(.A(new_n725), .B(new_n726), .C1(new_n727), .C2(new_n737), .ZN(new_n738));
  AOI211_X1 g552(.A(new_n652), .B(new_n602), .C1(new_n589), .C2(new_n530), .ZN(new_n739));
  AND2_X1   g553(.A1(new_n736), .A2(new_n354), .ZN(new_n740));
  NAND4_X1  g554(.A1(new_n739), .A2(KEYINPUT112), .A3(new_n724), .A4(new_n740), .ZN(new_n741));
  NAND2_X1  g555(.A1(new_n738), .A2(new_n741), .ZN(new_n742));
  XNOR2_X1  g556(.A(new_n742), .B(new_n482), .ZN(G33));
  NAND2_X1  g557(.A1(new_n740), .A2(new_n653), .ZN(new_n744));
  XNOR2_X1  g558(.A(new_n744), .B(G134), .ZN(G36));
  NAND3_X1  g559(.A1(new_n415), .A2(new_n355), .A3(new_n417), .ZN(new_n746));
  INV_X1    g560(.A(new_n746), .ZN(new_n747));
  OR3_X1    g561(.A1(new_n521), .A2(KEYINPUT113), .A3(new_n531), .ZN(new_n748));
  NAND2_X1  g562(.A1(new_n683), .A2(KEYINPUT113), .ZN(new_n749));
  AOI21_X1  g563(.A(new_n602), .B1(new_n748), .B2(new_n749), .ZN(new_n750));
  NAND2_X1  g564(.A1(new_n750), .A2(KEYINPUT43), .ZN(new_n751));
  INV_X1    g565(.A(KEYINPUT43), .ZN(new_n752));
  OAI21_X1  g566(.A(new_n752), .B1(new_n683), .B2(new_n602), .ZN(new_n753));
  NAND2_X1  g567(.A1(new_n751), .A2(new_n753), .ZN(new_n754));
  NAND2_X1  g568(.A1(new_n609), .A2(new_n635), .ZN(new_n755));
  XNOR2_X1  g569(.A(new_n755), .B(KEYINPUT114), .ZN(new_n756));
  NAND2_X1  g570(.A1(new_n754), .A2(new_n756), .ZN(new_n757));
  INV_X1    g571(.A(KEYINPUT44), .ZN(new_n758));
  OAI21_X1  g572(.A(new_n747), .B1(new_n757), .B2(new_n758), .ZN(new_n759));
  INV_X1    g573(.A(KEYINPUT115), .ZN(new_n760));
  NAND2_X1  g574(.A1(new_n759), .A2(new_n760), .ZN(new_n761));
  NAND2_X1  g575(.A1(new_n446), .A2(new_n448), .ZN(new_n762));
  XNOR2_X1  g576(.A(new_n762), .B(KEYINPUT45), .ZN(new_n763));
  OAI21_X1  g577(.A(G469), .B1(new_n763), .B2(G902), .ZN(new_n764));
  OR2_X1    g578(.A1(new_n764), .A2(KEYINPUT46), .ZN(new_n765));
  NAND2_X1  g579(.A1(new_n764), .A2(KEYINPUT46), .ZN(new_n766));
  NAND3_X1  g580(.A1(new_n765), .A2(new_n444), .A3(new_n766), .ZN(new_n767));
  NAND3_X1  g581(.A1(new_n767), .A2(new_n452), .A3(new_n658), .ZN(new_n768));
  AOI21_X1  g582(.A(new_n768), .B1(new_n757), .B2(new_n758), .ZN(new_n769));
  NAND2_X1  g583(.A1(new_n761), .A2(new_n769), .ZN(new_n770));
  NOR2_X1   g584(.A1(new_n759), .A2(new_n760), .ZN(new_n771));
  NOR2_X1   g585(.A1(new_n770), .A2(new_n771), .ZN(new_n772));
  XNOR2_X1  g586(.A(new_n772), .B(new_n217), .ZN(G39));
  NAND2_X1  g587(.A1(new_n767), .A2(new_n452), .ZN(new_n774));
  XNOR2_X1  g588(.A(new_n774), .B(KEYINPUT47), .ZN(new_n775));
  NAND2_X1  g589(.A1(new_n275), .A2(G472), .ZN(new_n776));
  NAND2_X1  g590(.A1(new_n776), .A2(new_n666), .ZN(new_n777));
  NOR4_X1   g591(.A1(new_n775), .A2(new_n777), .A3(new_n604), .A4(new_n746), .ZN(new_n778));
  NAND2_X1  g592(.A1(new_n778), .A2(new_n739), .ZN(new_n779));
  XNOR2_X1  g593(.A(new_n779), .B(G140), .ZN(G42));
  INV_X1    g594(.A(KEYINPUT120), .ZN(new_n781));
  INV_X1    g595(.A(KEYINPUT51), .ZN(new_n782));
  AND2_X1   g596(.A1(new_n677), .A2(new_n604), .ZN(new_n783));
  NOR2_X1   g597(.A1(new_n732), .A2(new_n691), .ZN(new_n784));
  NAND3_X1  g598(.A1(new_n783), .A2(new_n576), .A3(new_n784), .ZN(new_n785));
  NOR3_X1   g599(.A1(new_n785), .A2(new_n683), .A3(new_n684), .ZN(new_n786));
  AND3_X1   g600(.A1(new_n754), .A2(new_n576), .A3(new_n716), .ZN(new_n787));
  OR2_X1    g601(.A1(new_n691), .A2(new_n452), .ZN(new_n788));
  AOI21_X1  g602(.A(new_n746), .B1(new_n775), .B2(new_n788), .ZN(new_n789));
  AOI21_X1  g603(.A(new_n786), .B1(new_n787), .B2(new_n789), .ZN(new_n790));
  NOR3_X1   g604(.A1(new_n664), .A2(new_n708), .A3(new_n355), .ZN(new_n791));
  AOI21_X1  g605(.A(KEYINPUT50), .B1(new_n787), .B2(new_n791), .ZN(new_n792));
  AOI21_X1  g606(.A(new_n649), .B1(new_n751), .B2(new_n753), .ZN(new_n793));
  AND4_X1   g607(.A1(KEYINPUT50), .A2(new_n793), .A3(new_n716), .A4(new_n791), .ZN(new_n794));
  OAI21_X1  g608(.A(new_n790), .B1(new_n792), .B2(new_n794), .ZN(new_n795));
  INV_X1    g609(.A(new_n721), .ZN(new_n796));
  AOI21_X1  g610(.A(KEYINPUT121), .B1(new_n793), .B2(new_n784), .ZN(new_n797));
  INV_X1    g611(.A(new_n797), .ZN(new_n798));
  NAND3_X1  g612(.A1(new_n793), .A2(KEYINPUT121), .A3(new_n784), .ZN(new_n799));
  AOI21_X1  g613(.A(new_n796), .B1(new_n798), .B2(new_n799), .ZN(new_n800));
  OAI211_X1 g614(.A(new_n781), .B(new_n782), .C1(new_n795), .C2(new_n800), .ZN(new_n801));
  NAND2_X1  g615(.A1(new_n787), .A2(new_n720), .ZN(new_n802));
  NAND2_X1  g616(.A1(new_n683), .A2(new_n684), .ZN(new_n803));
  OAI211_X1 g617(.A(new_n802), .B(new_n574), .C1(new_n803), .C2(new_n785), .ZN(new_n804));
  INV_X1    g618(.A(new_n799), .ZN(new_n805));
  OAI21_X1  g619(.A(new_n354), .B1(new_n805), .B2(new_n797), .ZN(new_n806));
  NAND2_X1  g620(.A1(new_n806), .A2(KEYINPUT48), .ZN(new_n807));
  INV_X1    g621(.A(KEYINPUT48), .ZN(new_n808));
  OAI211_X1 g622(.A(new_n808), .B(new_n354), .C1(new_n805), .C2(new_n797), .ZN(new_n809));
  AOI21_X1  g623(.A(new_n804), .B1(new_n807), .B2(new_n809), .ZN(new_n810));
  AND2_X1   g624(.A1(new_n801), .A2(new_n810), .ZN(new_n811));
  INV_X1    g625(.A(KEYINPUT53), .ZN(new_n812));
  NAND2_X1  g626(.A1(new_n685), .A2(new_n452), .ZN(new_n813));
  OR3_X1    g627(.A1(new_n731), .A2(new_n635), .A3(new_n813), .ZN(new_n814));
  AOI21_X1  g628(.A(new_n814), .B1(new_n674), .B2(new_n676), .ZN(new_n815));
  NAND4_X1  g629(.A1(new_n815), .A2(new_n683), .A3(new_n572), .A4(new_n418), .ZN(new_n816));
  NAND4_X1  g630(.A1(new_n722), .A2(new_n656), .A3(new_n686), .A4(new_n816), .ZN(new_n817));
  INV_X1    g631(.A(KEYINPUT52), .ZN(new_n818));
  NAND2_X1  g632(.A1(new_n817), .A2(new_n818), .ZN(new_n819));
  NOR2_X1   g633(.A1(new_n644), .A2(new_n645), .ZN(new_n820));
  OAI211_X1 g634(.A(new_n685), .B(new_n655), .C1(new_n603), .C2(new_n820), .ZN(new_n821));
  NAND4_X1  g635(.A1(new_n821), .A2(new_n722), .A3(KEYINPUT52), .A4(new_n816), .ZN(new_n822));
  NAND2_X1  g636(.A1(new_n819), .A2(new_n822), .ZN(new_n823));
  OAI21_X1  g637(.A(new_n803), .B1(new_n683), .B2(new_n573), .ZN(new_n824));
  NOR3_X1   g638(.A1(new_n606), .A2(new_n609), .A3(new_n611), .ZN(new_n825));
  NAND2_X1  g639(.A1(new_n824), .A2(new_n825), .ZN(new_n826));
  AND3_X1   g640(.A1(new_n591), .A2(new_n641), .A3(new_n826), .ZN(new_n827));
  NAND3_X1  g641(.A1(new_n570), .A2(new_n571), .A3(new_n685), .ZN(new_n828));
  NOR3_X1   g642(.A1(new_n828), .A2(new_n746), .A3(new_n453), .ZN(new_n829));
  AND3_X1   g643(.A1(new_n639), .A2(new_n530), .A3(new_n829), .ZN(new_n830));
  INV_X1    g644(.A(KEYINPUT116), .ZN(new_n831));
  NAND4_X1  g645(.A1(new_n830), .A2(new_n619), .A3(new_n831), .A4(new_n777), .ZN(new_n832));
  NAND4_X1  g646(.A1(new_n639), .A2(new_n777), .A3(new_n829), .A4(new_n530), .ZN(new_n833));
  OAI21_X1  g647(.A(KEYINPUT116), .B1(new_n833), .B2(new_n644), .ZN(new_n834));
  AOI22_X1  g648(.A1(new_n832), .A2(new_n834), .B1(new_n653), .B2(new_n740), .ZN(new_n835));
  NAND3_X1  g649(.A1(new_n739), .A2(new_n721), .A3(new_n736), .ZN(new_n836));
  AND4_X1   g650(.A1(new_n741), .A2(new_n835), .A3(new_n738), .A4(new_n836), .ZN(new_n837));
  NAND3_X1  g651(.A1(new_n823), .A2(new_n827), .A3(new_n837), .ZN(new_n838));
  AND3_X1   g652(.A1(new_n699), .A2(new_n710), .A3(new_n718), .ZN(new_n839));
  OAI21_X1  g653(.A(new_n696), .B1(new_n626), .B2(new_n627), .ZN(new_n840));
  NAND2_X1  g654(.A1(new_n839), .A2(new_n840), .ZN(new_n841));
  OAI21_X1  g655(.A(new_n812), .B1(new_n838), .B2(new_n841), .ZN(new_n842));
  INV_X1    g656(.A(KEYINPUT117), .ZN(new_n843));
  NAND2_X1  g657(.A1(new_n842), .A2(new_n843), .ZN(new_n844));
  NAND3_X1  g658(.A1(new_n699), .A2(new_n710), .A3(new_n718), .ZN(new_n845));
  NOR2_X1   g659(.A1(new_n706), .A2(new_n845), .ZN(new_n846));
  NAND3_X1  g660(.A1(new_n591), .A2(new_n641), .A3(new_n826), .ZN(new_n847));
  NAND4_X1  g661(.A1(new_n835), .A2(new_n738), .A3(new_n741), .A4(new_n836), .ZN(new_n848));
  NOR2_X1   g662(.A1(new_n847), .A2(new_n848), .ZN(new_n849));
  NAND4_X1  g663(.A1(new_n846), .A2(KEYINPUT53), .A3(new_n823), .A4(new_n849), .ZN(new_n850));
  INV_X1    g664(.A(KEYINPUT118), .ZN(new_n851));
  NAND2_X1  g665(.A1(new_n850), .A2(new_n851), .ZN(new_n852));
  AND3_X1   g666(.A1(new_n823), .A2(new_n827), .A3(new_n837), .ZN(new_n853));
  NAND4_X1  g667(.A1(new_n853), .A2(KEYINPUT118), .A3(KEYINPUT53), .A4(new_n846), .ZN(new_n854));
  OAI211_X1 g668(.A(KEYINPUT117), .B(new_n812), .C1(new_n838), .C2(new_n841), .ZN(new_n855));
  NAND4_X1  g669(.A1(new_n844), .A2(new_n852), .A3(new_n854), .A4(new_n855), .ZN(new_n856));
  NAND2_X1  g670(.A1(new_n856), .A2(KEYINPUT54), .ZN(new_n857));
  INV_X1    g671(.A(KEYINPUT54), .ZN(new_n858));
  NAND3_X1  g672(.A1(new_n842), .A2(new_n858), .A3(new_n850), .ZN(new_n859));
  INV_X1    g673(.A(KEYINPUT119), .ZN(new_n860));
  NAND2_X1  g674(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  NAND4_X1  g675(.A1(new_n842), .A2(new_n850), .A3(KEYINPUT119), .A4(new_n858), .ZN(new_n862));
  NAND2_X1  g676(.A1(new_n861), .A2(new_n862), .ZN(new_n863));
  OAI21_X1  g677(.A(new_n781), .B1(new_n795), .B2(new_n800), .ZN(new_n864));
  NAND2_X1  g678(.A1(new_n864), .A2(KEYINPUT51), .ZN(new_n865));
  NAND4_X1  g679(.A1(new_n811), .A2(new_n857), .A3(new_n863), .A4(new_n865), .ZN(new_n866));
  OAI21_X1  g680(.A(new_n866), .B1(G952), .B2(G953), .ZN(new_n867));
  XOR2_X1   g681(.A(new_n691), .B(KEYINPUT49), .Z(new_n868));
  AND4_X1   g682(.A1(new_n452), .A2(new_n663), .A3(new_n355), .A4(new_n868), .ZN(new_n869));
  NAND3_X1  g683(.A1(new_n750), .A2(new_n783), .A3(new_n869), .ZN(new_n870));
  NAND2_X1  g684(.A1(new_n867), .A2(new_n870), .ZN(G75));
  NOR2_X1   g685(.A1(new_n248), .A2(G952), .ZN(new_n872));
  INV_X1    g686(.A(new_n872), .ZN(new_n873));
  AOI21_X1  g687(.A(new_n265), .B1(new_n842), .B2(new_n850), .ZN(new_n874));
  AOI21_X1  g688(.A(KEYINPUT56), .B1(new_n874), .B2(new_n414), .ZN(new_n875));
  NAND2_X1  g689(.A1(new_n407), .A2(new_n409), .ZN(new_n876));
  XNOR2_X1  g690(.A(new_n876), .B(new_n410), .ZN(new_n877));
  XNOR2_X1  g691(.A(new_n877), .B(KEYINPUT55), .ZN(new_n878));
  OAI21_X1  g692(.A(new_n873), .B1(new_n875), .B2(new_n878), .ZN(new_n879));
  AOI21_X1  g693(.A(new_n879), .B1(new_n875), .B2(new_n878), .ZN(G51));
  NAND2_X1  g694(.A1(new_n842), .A2(new_n850), .ZN(new_n881));
  NAND2_X1  g695(.A1(new_n881), .A2(KEYINPUT54), .ZN(new_n882));
  NAND2_X1  g696(.A1(new_n882), .A2(new_n859), .ZN(new_n883));
  NAND2_X1  g697(.A1(G469), .A2(G902), .ZN(new_n884));
  XOR2_X1   g698(.A(new_n884), .B(KEYINPUT57), .Z(new_n885));
  NAND2_X1  g699(.A1(new_n883), .A2(new_n885), .ZN(new_n886));
  NAND2_X1  g700(.A1(new_n886), .A2(new_n442), .ZN(new_n887));
  NAND3_X1  g701(.A1(new_n874), .A2(G469), .A3(new_n763), .ZN(new_n888));
  AOI21_X1  g702(.A(new_n872), .B1(new_n887), .B2(new_n888), .ZN(G54));
  NAND3_X1  g703(.A1(new_n874), .A2(KEYINPUT58), .A3(G475), .ZN(new_n890));
  INV_X1    g704(.A(new_n617), .ZN(new_n891));
  OAI21_X1  g705(.A(new_n873), .B1(new_n890), .B2(new_n891), .ZN(new_n892));
  AOI21_X1  g706(.A(new_n892), .B1(new_n891), .B2(new_n890), .ZN(G60));
  NAND2_X1  g707(.A1(G478), .A2(G902), .ZN(new_n894));
  XOR2_X1   g708(.A(new_n894), .B(KEYINPUT59), .Z(new_n895));
  INV_X1    g709(.A(new_n895), .ZN(new_n896));
  AND2_X1   g710(.A1(new_n599), .A2(new_n896), .ZN(new_n897));
  AOI21_X1  g711(.A(new_n872), .B1(new_n883), .B2(new_n897), .ZN(new_n898));
  AOI21_X1  g712(.A(new_n895), .B1(new_n857), .B2(new_n863), .ZN(new_n899));
  OAI21_X1  g713(.A(new_n898), .B1(new_n899), .B2(new_n599), .ZN(new_n900));
  NAND2_X1  g714(.A1(new_n900), .A2(KEYINPUT122), .ZN(new_n901));
  INV_X1    g715(.A(KEYINPUT122), .ZN(new_n902));
  OAI211_X1 g716(.A(new_n898), .B(new_n902), .C1(new_n899), .C2(new_n599), .ZN(new_n903));
  NAND2_X1  g717(.A1(new_n901), .A2(new_n903), .ZN(G63));
  INV_X1    g718(.A(KEYINPUT61), .ZN(new_n905));
  NOR2_X1   g719(.A1(new_n905), .A2(KEYINPUT124), .ZN(new_n906));
  XNOR2_X1  g720(.A(KEYINPUT123), .B(KEYINPUT60), .ZN(new_n907));
  NOR2_X1   g721(.A1(new_n339), .A2(new_n265), .ZN(new_n908));
  XNOR2_X1  g722(.A(new_n907), .B(new_n908), .ZN(new_n909));
  NAND2_X1  g723(.A1(new_n881), .A2(new_n909), .ZN(new_n910));
  NOR2_X1   g724(.A1(new_n336), .A2(new_n337), .ZN(new_n911));
  AOI21_X1  g725(.A(new_n872), .B1(new_n910), .B2(new_n911), .ZN(new_n912));
  NAND3_X1  g726(.A1(new_n881), .A2(new_n633), .A3(new_n909), .ZN(new_n913));
  AOI21_X1  g727(.A(new_n906), .B1(new_n912), .B2(new_n913), .ZN(new_n914));
  NAND2_X1  g728(.A1(new_n905), .A2(KEYINPUT124), .ZN(new_n915));
  XOR2_X1   g729(.A(new_n914), .B(new_n915), .Z(G66));
  OAI21_X1  g730(.A(G953), .B1(new_n579), .B2(new_n387), .ZN(new_n917));
  NOR2_X1   g731(.A1(new_n841), .A2(new_n847), .ZN(new_n918));
  OAI21_X1  g732(.A(new_n917), .B1(new_n918), .B2(new_n577), .ZN(new_n919));
  XOR2_X1   g733(.A(new_n919), .B(KEYINPUT125), .Z(new_n920));
  OAI21_X1  g734(.A(new_n876), .B1(G898), .B2(new_n248), .ZN(new_n921));
  XNOR2_X1  g735(.A(new_n920), .B(new_n921), .ZN(G69));
  NOR2_X1   g736(.A1(new_n237), .A2(new_n241), .ZN(new_n923));
  XNOR2_X1  g737(.A(new_n503), .B(KEYINPUT126), .ZN(new_n924));
  XNOR2_X1  g738(.A(new_n923), .B(new_n924), .ZN(new_n925));
  XOR2_X1   g739(.A(new_n925), .B(G227), .Z(new_n926));
  NOR3_X1   g740(.A1(new_n926), .A2(new_n650), .A3(new_n248), .ZN(new_n927));
  INV_X1    g741(.A(new_n354), .ZN(new_n928));
  NOR3_X1   g742(.A1(new_n928), .A2(new_n659), .A3(new_n746), .ZN(new_n929));
  NAND2_X1  g743(.A1(new_n824), .A2(new_n929), .ZN(new_n930));
  NAND2_X1  g744(.A1(new_n779), .A2(new_n930), .ZN(new_n931));
  NAND2_X1  g745(.A1(new_n821), .A2(new_n722), .ZN(new_n932));
  INV_X1    g746(.A(new_n932), .ZN(new_n933));
  NAND4_X1  g747(.A1(new_n933), .A2(KEYINPUT127), .A3(new_n680), .A4(KEYINPUT62), .ZN(new_n934));
  NAND2_X1  g748(.A1(new_n933), .A2(new_n680), .ZN(new_n935));
  XOR2_X1   g749(.A(KEYINPUT127), .B(KEYINPUT62), .Z(new_n936));
  NAND2_X1  g750(.A1(new_n935), .A2(new_n936), .ZN(new_n937));
  AOI21_X1  g751(.A(new_n931), .B1(new_n934), .B2(new_n937), .ZN(new_n938));
  OAI211_X1 g752(.A(new_n925), .B(new_n938), .C1(new_n770), .C2(new_n771), .ZN(new_n939));
  NOR2_X1   g753(.A1(new_n768), .A2(new_n928), .ZN(new_n940));
  NAND3_X1  g754(.A1(new_n679), .A2(new_n940), .A3(new_n418), .ZN(new_n941));
  NAND3_X1  g755(.A1(new_n779), .A2(new_n744), .A3(new_n941), .ZN(new_n942));
  NOR4_X1   g756(.A1(new_n772), .A2(new_n742), .A3(new_n932), .A4(new_n942), .ZN(new_n943));
  OAI21_X1  g757(.A(new_n939), .B1(new_n943), .B2(new_n925), .ZN(new_n944));
  AOI21_X1  g758(.A(new_n927), .B1(new_n944), .B2(new_n248), .ZN(G72));
  NAND2_X1  g759(.A1(G472), .A2(G902), .ZN(new_n946));
  XOR2_X1   g760(.A(new_n946), .B(KEYINPUT63), .Z(new_n947));
  NAND3_X1  g761(.A1(new_n254), .A2(new_n257), .A3(new_n276), .ZN(new_n948));
  NAND3_X1  g762(.A1(new_n856), .A2(new_n947), .A3(new_n948), .ZN(new_n949));
  NOR2_X1   g763(.A1(new_n245), .A2(new_n256), .ZN(new_n950));
  NOR2_X1   g764(.A1(new_n244), .A2(new_n253), .ZN(new_n951));
  NOR2_X1   g765(.A1(new_n950), .A2(new_n951), .ZN(new_n952));
  OAI211_X1 g766(.A(new_n949), .B(new_n873), .C1(new_n947), .C2(new_n952), .ZN(new_n953));
  NAND2_X1  g767(.A1(new_n943), .A2(new_n951), .ZN(new_n954));
  OAI211_X1 g768(.A(new_n938), .B(new_n950), .C1(new_n770), .C2(new_n771), .ZN(new_n955));
  NAND2_X1  g769(.A1(new_n954), .A2(new_n955), .ZN(new_n956));
  AOI21_X1  g770(.A(new_n953), .B1(new_n956), .B2(new_n918), .ZN(G57));
endmodule


