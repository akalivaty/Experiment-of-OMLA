//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 0 1 0 1 0 1 1 0 0 1 0 0 1 1 1 0 1 0 1 1 0 0 1 0 0 1 1 1 1 1 1 0 0 1 0 1 0 1 0 0 0 0 0 1 1 1 0 0 0 1 0 0 0 0 0 1 0 0 1 1 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:38:41 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n228, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n237, new_n238, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n245, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1087,
    new_n1088, new_n1089, new_n1090, new_n1091, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1108, new_n1109, new_n1110, new_n1111, new_n1112,
    new_n1113, new_n1114, new_n1115, new_n1116, new_n1117, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1186, new_n1187, new_n1188, new_n1189, new_n1190, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1251, new_n1252, new_n1253,
    new_n1254, new_n1255, new_n1256, new_n1257, new_n1258, new_n1259,
    new_n1260, new_n1261, new_n1262, new_n1263, new_n1264, new_n1265,
    new_n1266, new_n1267, new_n1268, new_n1269, new_n1270, new_n1271,
    new_n1272, new_n1273, new_n1274, new_n1275, new_n1277, new_n1278,
    new_n1279, new_n1280, new_n1282, new_n1283, new_n1284, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1346,
    new_n1347, new_n1348, new_n1349, new_n1351, new_n1352, new_n1353,
    new_n1354, new_n1355;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0005(.A1(G1), .A2(G20), .ZN(new_n206));
  AOI22_X1  g0006(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n207));
  XOR2_X1   g0007(.A(new_n207), .B(KEYINPUT64), .Z(new_n208));
  AOI22_X1  g0008(.A1(G87), .A2(G250), .B1(G116), .B2(G270), .ZN(new_n209));
  AOI22_X1  g0009(.A1(G50), .A2(G226), .B1(G68), .B2(G238), .ZN(new_n210));
  AOI22_X1  g0010(.A1(G77), .A2(G244), .B1(G97), .B2(G257), .ZN(new_n211));
  NAND3_X1  g0011(.A1(new_n209), .A2(new_n210), .A3(new_n211), .ZN(new_n212));
  OAI21_X1  g0012(.A(new_n206), .B1(new_n208), .B2(new_n212), .ZN(new_n213));
  NAND2_X1  g0013(.A1(new_n213), .A2(KEYINPUT1), .ZN(new_n214));
  XOR2_X1   g0014(.A(new_n214), .B(KEYINPUT65), .Z(new_n215));
  INV_X1    g0015(.A(new_n201), .ZN(new_n216));
  NAND2_X1  g0016(.A1(new_n216), .A2(G50), .ZN(new_n217));
  INV_X1    g0017(.A(new_n217), .ZN(new_n218));
  NAND2_X1  g0018(.A1(G1), .A2(G13), .ZN(new_n219));
  INV_X1    g0019(.A(G20), .ZN(new_n220));
  NOR2_X1   g0020(.A1(new_n219), .A2(new_n220), .ZN(new_n221));
  NAND2_X1  g0021(.A1(new_n218), .A2(new_n221), .ZN(new_n222));
  NOR2_X1   g0022(.A1(new_n206), .A2(G13), .ZN(new_n223));
  OAI211_X1 g0023(.A(new_n223), .B(G250), .C1(G257), .C2(G264), .ZN(new_n224));
  XNOR2_X1  g0024(.A(new_n224), .B(KEYINPUT0), .ZN(new_n225));
  OAI211_X1 g0025(.A(new_n222), .B(new_n225), .C1(new_n213), .C2(KEYINPUT1), .ZN(new_n226));
  NOR2_X1   g0026(.A1(new_n215), .A2(new_n226), .ZN(G361));
  XNOR2_X1  g0027(.A(G238), .B(G244), .ZN(new_n228));
  INV_X1    g0028(.A(G232), .ZN(new_n229));
  XNOR2_X1  g0029(.A(new_n228), .B(new_n229), .ZN(new_n230));
  XOR2_X1   g0030(.A(KEYINPUT2), .B(G226), .Z(new_n231));
  XNOR2_X1  g0031(.A(new_n230), .B(new_n231), .ZN(new_n232));
  XOR2_X1   g0032(.A(G264), .B(G270), .Z(new_n233));
  XNOR2_X1  g0033(.A(G250), .B(G257), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n233), .B(new_n234), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n232), .B(new_n235), .ZN(G358));
  XOR2_X1   g0036(.A(G87), .B(G97), .Z(new_n237));
  XNOR2_X1  g0037(.A(G107), .B(G116), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  NAND2_X1  g0039(.A1(new_n202), .A2(G68), .ZN(new_n240));
  INV_X1    g0040(.A(G68), .ZN(new_n241));
  NAND2_X1  g0041(.A1(new_n241), .A2(G50), .ZN(new_n242));
  NAND2_X1  g0042(.A1(new_n240), .A2(new_n242), .ZN(new_n243));
  XNOR2_X1  g0043(.A(G58), .B(G77), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n239), .B(new_n245), .ZN(G351));
  XNOR2_X1  g0046(.A(KEYINPUT66), .B(G45), .ZN(new_n247));
  INV_X1    g0047(.A(G41), .ZN(new_n248));
  NAND2_X1  g0048(.A1(new_n247), .A2(new_n248), .ZN(new_n249));
  INV_X1    g0049(.A(G1), .ZN(new_n250));
  NAND3_X1  g0050(.A1(new_n249), .A2(new_n250), .A3(G274), .ZN(new_n251));
  NOR2_X1   g0051(.A1(G226), .A2(G1698), .ZN(new_n252));
  AOI21_X1  g0052(.A(new_n252), .B1(new_n229), .B2(G1698), .ZN(new_n253));
  XNOR2_X1  g0053(.A(KEYINPUT3), .B(G33), .ZN(new_n254));
  AOI22_X1  g0054(.A1(new_n253), .A2(new_n254), .B1(G33), .B2(G97), .ZN(new_n255));
  AOI21_X1  g0055(.A(new_n219), .B1(G33), .B2(G41), .ZN(new_n256));
  INV_X1    g0056(.A(new_n256), .ZN(new_n257));
  INV_X1    g0057(.A(G238), .ZN(new_n258));
  XNOR2_X1  g0058(.A(KEYINPUT67), .B(G1), .ZN(new_n259));
  NOR2_X1   g0059(.A1(G41), .A2(G45), .ZN(new_n260));
  OAI21_X1  g0060(.A(new_n257), .B1(new_n259), .B2(new_n260), .ZN(new_n261));
  OAI221_X1 g0061(.A(new_n251), .B1(new_n255), .B2(new_n257), .C1(new_n258), .C2(new_n261), .ZN(new_n262));
  NAND2_X1  g0062(.A1(new_n262), .A2(KEYINPUT13), .ZN(new_n263));
  INV_X1    g0063(.A(new_n263), .ZN(new_n264));
  NOR2_X1   g0064(.A1(new_n262), .A2(KEYINPUT13), .ZN(new_n265));
  OAI21_X1  g0065(.A(G169), .B1(new_n264), .B2(new_n265), .ZN(new_n266));
  NAND2_X1  g0066(.A1(new_n266), .A2(KEYINPUT14), .ZN(new_n267));
  INV_X1    g0067(.A(new_n265), .ZN(new_n268));
  NAND2_X1  g0068(.A1(new_n268), .A2(new_n263), .ZN(new_n269));
  INV_X1    g0069(.A(KEYINPUT14), .ZN(new_n270));
  NAND3_X1  g0070(.A1(new_n269), .A2(new_n270), .A3(G169), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n264), .A2(KEYINPUT72), .ZN(new_n272));
  INV_X1    g0072(.A(KEYINPUT72), .ZN(new_n273));
  NAND2_X1  g0073(.A1(new_n263), .A2(new_n273), .ZN(new_n274));
  NAND3_X1  g0074(.A1(new_n272), .A2(new_n274), .A3(new_n268), .ZN(new_n275));
  INV_X1    g0075(.A(G179), .ZN(new_n276));
  OAI211_X1 g0076(.A(new_n267), .B(new_n271), .C1(new_n275), .C2(new_n276), .ZN(new_n277));
  NOR2_X1   g0077(.A1(G20), .A2(G33), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n278), .A2(G50), .ZN(new_n279));
  INV_X1    g0079(.A(G77), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n220), .A2(G33), .ZN(new_n281));
  OAI221_X1 g0081(.A(new_n279), .B1(new_n220), .B2(G68), .C1(new_n280), .C2(new_n281), .ZN(new_n282));
  NAND3_X1  g0082(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n283), .A2(new_n219), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n282), .A2(new_n284), .ZN(new_n285));
  XOR2_X1   g0085(.A(new_n285), .B(KEYINPUT11), .Z(new_n286));
  INV_X1    g0086(.A(KEYINPUT73), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n286), .A2(new_n287), .ZN(new_n288));
  XNOR2_X1  g0088(.A(new_n285), .B(KEYINPUT11), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n289), .A2(KEYINPUT73), .ZN(new_n290));
  OR2_X1    g0090(.A1(KEYINPUT67), .A2(G1), .ZN(new_n291));
  NAND2_X1  g0091(.A1(KEYINPUT67), .A2(G1), .ZN(new_n292));
  NAND4_X1  g0092(.A1(new_n291), .A2(G13), .A3(G20), .A4(new_n292), .ZN(new_n293));
  OR3_X1    g0093(.A1(new_n293), .A2(KEYINPUT12), .A3(G68), .ZN(new_n294));
  OAI21_X1  g0094(.A(KEYINPUT12), .B1(new_n293), .B2(G68), .ZN(new_n295));
  AND2_X1   g0095(.A1(new_n291), .A2(new_n292), .ZN(new_n296));
  AOI21_X1  g0096(.A(new_n284), .B1(new_n296), .B2(G20), .ZN(new_n297));
  AOI22_X1  g0097(.A1(new_n294), .A2(new_n295), .B1(G68), .B2(new_n297), .ZN(new_n298));
  NAND3_X1  g0098(.A1(new_n288), .A2(new_n290), .A3(new_n298), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n277), .A2(new_n299), .ZN(new_n300));
  INV_X1    g0100(.A(new_n300), .ZN(new_n301));
  AOI21_X1  g0101(.A(new_n299), .B1(new_n269), .B2(G200), .ZN(new_n302));
  NAND4_X1  g0102(.A1(new_n272), .A2(G190), .A3(new_n274), .A4(new_n268), .ZN(new_n303));
  AND2_X1   g0103(.A1(new_n302), .A2(new_n303), .ZN(new_n304));
  NOR2_X1   g0104(.A1(new_n301), .A2(new_n304), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n297), .A2(G50), .ZN(new_n306));
  OAI21_X1  g0106(.A(new_n306), .B1(G50), .B2(new_n293), .ZN(new_n307));
  INV_X1    g0107(.A(new_n284), .ZN(new_n308));
  NOR2_X1   g0108(.A1(KEYINPUT8), .A2(G58), .ZN(new_n309));
  INV_X1    g0109(.A(G58), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n310), .A2(KEYINPUT68), .ZN(new_n311));
  INV_X1    g0111(.A(KEYINPUT68), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n312), .A2(G58), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n311), .A2(new_n313), .ZN(new_n314));
  AOI21_X1  g0114(.A(new_n309), .B1(new_n314), .B2(KEYINPUT8), .ZN(new_n315));
  INV_X1    g0115(.A(G33), .ZN(new_n316));
  NOR2_X1   g0116(.A1(new_n316), .A2(G20), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n315), .A2(new_n317), .ZN(new_n318));
  AOI22_X1  g0118(.A1(new_n203), .A2(G20), .B1(G150), .B2(new_n278), .ZN(new_n319));
  AOI21_X1  g0119(.A(new_n308), .B1(new_n318), .B2(new_n319), .ZN(new_n320));
  NOR2_X1   g0120(.A1(new_n307), .A2(new_n320), .ZN(new_n321));
  INV_X1    g0121(.A(G169), .ZN(new_n322));
  INV_X1    g0122(.A(G1698), .ZN(new_n323));
  NAND3_X1  g0123(.A1(new_n254), .A2(G222), .A3(new_n323), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n254), .A2(G1698), .ZN(new_n325));
  INV_X1    g0125(.A(G223), .ZN(new_n326));
  OAI221_X1 g0126(.A(new_n324), .B1(new_n280), .B2(new_n254), .C1(new_n325), .C2(new_n326), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n327), .A2(new_n256), .ZN(new_n328));
  INV_X1    g0128(.A(G274), .ZN(new_n329));
  AOI211_X1 g0129(.A(G1), .B(new_n329), .C1(new_n247), .C2(new_n248), .ZN(new_n330));
  NOR2_X1   g0130(.A1(new_n259), .A2(new_n260), .ZN(new_n331));
  NOR2_X1   g0131(.A1(new_n331), .A2(new_n256), .ZN(new_n332));
  AOI21_X1  g0132(.A(new_n330), .B1(new_n332), .B2(G226), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n328), .A2(new_n333), .ZN(new_n334));
  AOI21_X1  g0134(.A(new_n321), .B1(new_n322), .B2(new_n334), .ZN(new_n335));
  OAI21_X1  g0135(.A(new_n335), .B1(G179), .B2(new_n334), .ZN(new_n336));
  XNOR2_X1  g0136(.A(new_n336), .B(KEYINPUT69), .ZN(new_n337));
  OR2_X1    g0137(.A1(new_n321), .A2(KEYINPUT9), .ZN(new_n338));
  AOI22_X1  g0138(.A1(new_n321), .A2(KEYINPUT9), .B1(new_n334), .B2(G200), .ZN(new_n339));
  NAND3_X1  g0139(.A1(new_n328), .A2(G190), .A3(new_n333), .ZN(new_n340));
  NAND3_X1  g0140(.A1(new_n338), .A2(new_n339), .A3(new_n340), .ZN(new_n341));
  XNOR2_X1  g0141(.A(new_n341), .B(KEYINPUT10), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n297), .A2(G77), .ZN(new_n343));
  XOR2_X1   g0143(.A(new_n343), .B(KEYINPUT70), .Z(new_n344));
  NOR2_X1   g0144(.A1(new_n293), .A2(G77), .ZN(new_n345));
  XOR2_X1   g0145(.A(KEYINPUT8), .B(G58), .Z(new_n346));
  AOI22_X1  g0146(.A1(new_n346), .A2(new_n278), .B1(G20), .B2(G77), .ZN(new_n347));
  XNOR2_X1  g0147(.A(KEYINPUT15), .B(G87), .ZN(new_n348));
  OAI21_X1  g0148(.A(new_n347), .B1(new_n281), .B2(new_n348), .ZN(new_n349));
  AOI21_X1  g0149(.A(new_n345), .B1(new_n349), .B2(new_n284), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n344), .A2(new_n350), .ZN(new_n351));
  OR2_X1    g0151(.A1(new_n351), .A2(KEYINPUT71), .ZN(new_n352));
  NAND3_X1  g0152(.A1(new_n254), .A2(G232), .A3(new_n323), .ZN(new_n353));
  INV_X1    g0153(.A(G107), .ZN(new_n354));
  OAI221_X1 g0154(.A(new_n353), .B1(new_n354), .B2(new_n254), .C1(new_n325), .C2(new_n258), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n355), .A2(new_n256), .ZN(new_n356));
  AOI21_X1  g0156(.A(new_n330), .B1(new_n332), .B2(G244), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n356), .A2(new_n357), .ZN(new_n358));
  INV_X1    g0158(.A(new_n358), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n359), .A2(G190), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n351), .A2(KEYINPUT71), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n358), .A2(G200), .ZN(new_n362));
  NAND4_X1  g0162(.A1(new_n352), .A2(new_n360), .A3(new_n361), .A4(new_n362), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n359), .A2(new_n276), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n358), .A2(new_n322), .ZN(new_n365));
  NAND3_X1  g0165(.A1(new_n351), .A2(new_n364), .A3(new_n365), .ZN(new_n366));
  AND4_X1   g0166(.A1(new_n337), .A2(new_n342), .A3(new_n363), .A4(new_n366), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n326), .A2(new_n323), .ZN(new_n368));
  INV_X1    g0168(.A(G226), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n369), .A2(G1698), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n368), .A2(new_n370), .ZN(new_n371));
  INV_X1    g0171(.A(KEYINPUT3), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n372), .A2(G33), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n316), .A2(KEYINPUT3), .ZN(new_n374));
  INV_X1    g0174(.A(KEYINPUT74), .ZN(new_n375));
  NAND3_X1  g0175(.A1(new_n373), .A2(new_n374), .A3(new_n375), .ZN(new_n376));
  NAND3_X1  g0176(.A1(new_n372), .A2(KEYINPUT74), .A3(G33), .ZN(new_n377));
  AOI21_X1  g0177(.A(new_n371), .B1(new_n376), .B2(new_n377), .ZN(new_n378));
  NAND2_X1  g0178(.A1(G33), .A2(G87), .ZN(new_n379));
  INV_X1    g0179(.A(new_n379), .ZN(new_n380));
  OAI21_X1  g0180(.A(KEYINPUT76), .B1(new_n378), .B2(new_n380), .ZN(new_n381));
  INV_X1    g0181(.A(KEYINPUT76), .ZN(new_n382));
  AND3_X1   g0182(.A1(new_n372), .A2(KEYINPUT74), .A3(G33), .ZN(new_n383));
  AOI21_X1  g0183(.A(new_n383), .B1(new_n254), .B2(new_n375), .ZN(new_n384));
  OAI211_X1 g0184(.A(new_n382), .B(new_n379), .C1(new_n384), .C2(new_n371), .ZN(new_n385));
  NAND3_X1  g0185(.A1(new_n381), .A2(new_n385), .A3(new_n256), .ZN(new_n386));
  OAI21_X1  g0186(.A(new_n251), .B1(new_n261), .B2(new_n229), .ZN(new_n387));
  INV_X1    g0187(.A(new_n387), .ZN(new_n388));
  NAND3_X1  g0188(.A1(new_n386), .A2(G179), .A3(new_n388), .ZN(new_n389));
  OAI21_X1  g0189(.A(new_n379), .B1(new_n384), .B2(new_n371), .ZN(new_n390));
  AOI21_X1  g0190(.A(new_n257), .B1(new_n390), .B2(KEYINPUT76), .ZN(new_n391));
  AOI21_X1  g0191(.A(new_n387), .B1(new_n391), .B2(new_n385), .ZN(new_n392));
  OAI21_X1  g0192(.A(new_n389), .B1(new_n392), .B2(new_n322), .ZN(new_n393));
  XNOR2_X1  g0193(.A(KEYINPUT68), .B(G58), .ZN(new_n394));
  OAI21_X1  g0194(.A(new_n216), .B1(new_n394), .B2(new_n241), .ZN(new_n395));
  AOI22_X1  g0195(.A1(new_n395), .A2(G20), .B1(G159), .B2(new_n278), .ZN(new_n396));
  NAND2_X1  g0196(.A1(KEYINPUT75), .A2(KEYINPUT7), .ZN(new_n397));
  INV_X1    g0197(.A(KEYINPUT75), .ZN(new_n398));
  INV_X1    g0198(.A(KEYINPUT7), .ZN(new_n399));
  AOI21_X1  g0199(.A(G20), .B1(new_n398), .B2(new_n399), .ZN(new_n400));
  AOI21_X1  g0200(.A(new_n397), .B1(new_n384), .B2(new_n400), .ZN(new_n401));
  NAND4_X1  g0201(.A1(new_n376), .A2(new_n377), .A3(new_n400), .A4(new_n397), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n402), .A2(G68), .ZN(new_n403));
  OAI211_X1 g0203(.A(KEYINPUT16), .B(new_n396), .C1(new_n401), .C2(new_n403), .ZN(new_n404));
  INV_X1    g0204(.A(KEYINPUT16), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n278), .A2(G159), .ZN(new_n406));
  AOI21_X1  g0206(.A(new_n201), .B1(new_n314), .B2(G68), .ZN(new_n407));
  OAI21_X1  g0207(.A(new_n406), .B1(new_n407), .B2(new_n220), .ZN(new_n408));
  OAI21_X1  g0208(.A(new_n399), .B1(new_n254), .B2(G20), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n373), .A2(new_n374), .ZN(new_n410));
  NAND3_X1  g0210(.A1(new_n410), .A2(KEYINPUT7), .A3(new_n220), .ZN(new_n411));
  AOI21_X1  g0211(.A(new_n241), .B1(new_n409), .B2(new_n411), .ZN(new_n412));
  OAI21_X1  g0212(.A(new_n405), .B1(new_n408), .B2(new_n412), .ZN(new_n413));
  NAND3_X1  g0213(.A1(new_n404), .A2(new_n413), .A3(new_n284), .ZN(new_n414));
  INV_X1    g0214(.A(new_n315), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n415), .A2(new_n293), .ZN(new_n416));
  OAI21_X1  g0216(.A(new_n416), .B1(new_n297), .B2(new_n415), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n414), .A2(new_n417), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n393), .A2(new_n418), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n419), .A2(KEYINPUT18), .ZN(new_n420));
  INV_X1    g0220(.A(G200), .ZN(new_n421));
  AOI21_X1  g0221(.A(new_n421), .B1(new_n386), .B2(new_n388), .ZN(new_n422));
  AOI21_X1  g0222(.A(new_n422), .B1(G190), .B2(new_n392), .ZN(new_n423));
  AND2_X1   g0223(.A1(new_n414), .A2(new_n417), .ZN(new_n424));
  NAND3_X1  g0224(.A1(new_n423), .A2(KEYINPUT17), .A3(new_n424), .ZN(new_n425));
  INV_X1    g0225(.A(KEYINPUT18), .ZN(new_n426));
  NAND3_X1  g0226(.A1(new_n393), .A2(new_n426), .A3(new_n418), .ZN(new_n427));
  INV_X1    g0227(.A(KEYINPUT17), .ZN(new_n428));
  NAND3_X1  g0228(.A1(new_n386), .A2(G190), .A3(new_n388), .ZN(new_n429));
  OAI21_X1  g0229(.A(new_n429), .B1(new_n392), .B2(new_n421), .ZN(new_n430));
  OAI21_X1  g0230(.A(new_n428), .B1(new_n430), .B2(new_n418), .ZN(new_n431));
  NAND4_X1  g0231(.A1(new_n420), .A2(new_n425), .A3(new_n427), .A4(new_n431), .ZN(new_n432));
  INV_X1    g0232(.A(new_n432), .ZN(new_n433));
  NAND3_X1  g0233(.A1(new_n305), .A2(new_n367), .A3(new_n433), .ZN(new_n434));
  INV_X1    g0234(.A(new_n434), .ZN(new_n435));
  INV_X1    g0235(.A(KEYINPUT79), .ZN(new_n436));
  INV_X1    g0236(.A(KEYINPUT77), .ZN(new_n437));
  OAI21_X1  g0237(.A(G45), .B1(new_n248), .B2(KEYINPUT5), .ZN(new_n438));
  OAI21_X1  g0238(.A(new_n437), .B1(new_n259), .B2(new_n438), .ZN(new_n439));
  INV_X1    g0239(.A(KEYINPUT5), .ZN(new_n440));
  OAI21_X1  g0240(.A(G274), .B1(new_n440), .B2(G41), .ZN(new_n441));
  NOR2_X1   g0241(.A1(new_n256), .A2(new_n441), .ZN(new_n442));
  INV_X1    g0242(.A(G45), .ZN(new_n443));
  AOI21_X1  g0243(.A(new_n443), .B1(new_n440), .B2(G41), .ZN(new_n444));
  NAND4_X1  g0244(.A1(new_n444), .A2(KEYINPUT77), .A3(new_n291), .A4(new_n292), .ZN(new_n445));
  NAND3_X1  g0245(.A1(new_n439), .A2(new_n442), .A3(new_n445), .ZN(new_n446));
  INV_X1    g0246(.A(KEYINPUT78), .ZN(new_n447));
  NAND2_X1  g0247(.A1(new_n440), .A2(G41), .ZN(new_n448));
  NAND4_X1  g0248(.A1(new_n291), .A2(new_n448), .A3(G45), .A4(new_n292), .ZN(new_n449));
  NOR2_X1   g0249(.A1(new_n440), .A2(G41), .ZN(new_n450));
  OAI211_X1 g0250(.A(new_n257), .B(G257), .C1(new_n449), .C2(new_n450), .ZN(new_n451));
  AND3_X1   g0251(.A1(new_n446), .A2(new_n447), .A3(new_n451), .ZN(new_n452));
  AOI21_X1  g0252(.A(new_n447), .B1(new_n446), .B2(new_n451), .ZN(new_n453));
  OAI21_X1  g0253(.A(new_n436), .B1(new_n452), .B2(new_n453), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n446), .A2(new_n451), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n455), .A2(KEYINPUT78), .ZN(new_n456));
  NAND3_X1  g0256(.A1(new_n446), .A2(new_n447), .A3(new_n451), .ZN(new_n457));
  NAND3_X1  g0257(.A1(new_n456), .A2(KEYINPUT79), .A3(new_n457), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n454), .A2(new_n458), .ZN(new_n459));
  INV_X1    g0259(.A(G244), .ZN(new_n460));
  AOI21_X1  g0260(.A(new_n460), .B1(new_n376), .B2(new_n377), .ZN(new_n461));
  AOI21_X1  g0261(.A(KEYINPUT4), .B1(new_n461), .B2(new_n323), .ZN(new_n462));
  NAND4_X1  g0262(.A1(new_n254), .A2(KEYINPUT4), .A3(G244), .A4(new_n323), .ZN(new_n463));
  NAND2_X1  g0263(.A1(G33), .A2(G283), .ZN(new_n464));
  NAND3_X1  g0264(.A1(new_n254), .A2(G250), .A3(G1698), .ZN(new_n465));
  NAND3_X1  g0265(.A1(new_n463), .A2(new_n464), .A3(new_n465), .ZN(new_n466));
  OAI21_X1  g0266(.A(new_n256), .B1(new_n462), .B2(new_n466), .ZN(new_n467));
  AOI21_X1  g0267(.A(new_n421), .B1(new_n459), .B2(new_n467), .ZN(new_n468));
  NAND4_X1  g0268(.A1(new_n467), .A2(new_n456), .A3(G190), .A4(new_n457), .ZN(new_n469));
  NAND3_X1  g0269(.A1(new_n291), .A2(G33), .A3(new_n292), .ZN(new_n470));
  NAND3_X1  g0270(.A1(new_n293), .A2(new_n308), .A3(new_n470), .ZN(new_n471));
  INV_X1    g0271(.A(new_n471), .ZN(new_n472));
  NAND2_X1  g0272(.A1(new_n472), .A2(G97), .ZN(new_n473));
  INV_X1    g0273(.A(G97), .ZN(new_n474));
  NAND4_X1  g0274(.A1(new_n296), .A2(G13), .A3(G20), .A4(new_n474), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n473), .A2(new_n475), .ZN(new_n476));
  INV_X1    g0276(.A(KEYINPUT6), .ZN(new_n477));
  NOR2_X1   g0277(.A1(new_n474), .A2(new_n354), .ZN(new_n478));
  NOR2_X1   g0278(.A1(G97), .A2(G107), .ZN(new_n479));
  OAI21_X1  g0279(.A(new_n477), .B1(new_n478), .B2(new_n479), .ZN(new_n480));
  NAND3_X1  g0280(.A1(new_n354), .A2(KEYINPUT6), .A3(G97), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n480), .A2(new_n481), .ZN(new_n482));
  AOI22_X1  g0282(.A1(new_n482), .A2(G20), .B1(G77), .B2(new_n278), .ZN(new_n483));
  AND2_X1   g0283(.A1(new_n409), .A2(new_n411), .ZN(new_n484));
  OAI21_X1  g0284(.A(new_n483), .B1(new_n484), .B2(new_n354), .ZN(new_n485));
  AOI21_X1  g0285(.A(new_n476), .B1(new_n485), .B2(new_n284), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n469), .A2(new_n486), .ZN(new_n487));
  OAI21_X1  g0287(.A(KEYINPUT80), .B1(new_n468), .B2(new_n487), .ZN(new_n488));
  INV_X1    g0288(.A(new_n487), .ZN(new_n489));
  INV_X1    g0289(.A(KEYINPUT80), .ZN(new_n490));
  INV_X1    g0290(.A(new_n467), .ZN(new_n491));
  AOI21_X1  g0291(.A(new_n491), .B1(new_n454), .B2(new_n458), .ZN(new_n492));
  OAI211_X1 g0292(.A(new_n489), .B(new_n490), .C1(new_n421), .C2(new_n492), .ZN(new_n493));
  NAND3_X1  g0293(.A1(new_n459), .A2(new_n276), .A3(new_n467), .ZN(new_n494));
  NAND3_X1  g0294(.A1(new_n467), .A2(new_n456), .A3(new_n457), .ZN(new_n495));
  AOI21_X1  g0295(.A(new_n486), .B1(new_n322), .B2(new_n495), .ZN(new_n496));
  AOI22_X1  g0296(.A1(new_n488), .A2(new_n493), .B1(new_n494), .B2(new_n496), .ZN(new_n497));
  NOR2_X1   g0297(.A1(new_n293), .A2(G107), .ZN(new_n498));
  OR2_X1    g0298(.A1(new_n498), .A2(KEYINPUT25), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n498), .A2(KEYINPUT25), .ZN(new_n500));
  AOI22_X1  g0300(.A1(new_n499), .A2(new_n500), .B1(G107), .B2(new_n472), .ZN(new_n501));
  OAI211_X1 g0301(.A(new_n257), .B(G264), .C1(new_n449), .C2(new_n450), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n376), .A2(new_n377), .ZN(new_n503));
  NOR2_X1   g0303(.A1(G250), .A2(G1698), .ZN(new_n504));
  INV_X1    g0304(.A(G257), .ZN(new_n505));
  AOI21_X1  g0305(.A(new_n504), .B1(new_n505), .B2(G1698), .ZN(new_n506));
  AOI22_X1  g0306(.A1(new_n503), .A2(new_n506), .B1(G33), .B2(G294), .ZN(new_n507));
  OAI211_X1 g0307(.A(new_n446), .B(new_n502), .C1(new_n507), .C2(new_n257), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n508), .A2(new_n421), .ZN(new_n509));
  INV_X1    g0309(.A(new_n506), .ZN(new_n510));
  INV_X1    g0310(.A(G294), .ZN(new_n511));
  OAI22_X1  g0311(.A1(new_n384), .A2(new_n510), .B1(new_n316), .B2(new_n511), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n512), .A2(new_n256), .ZN(new_n513));
  INV_X1    g0313(.A(G190), .ZN(new_n514));
  NAND4_X1  g0314(.A1(new_n513), .A2(new_n514), .A3(new_n446), .A4(new_n502), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n509), .A2(new_n515), .ZN(new_n516));
  XNOR2_X1  g0316(.A(KEYINPUT85), .B(KEYINPUT22), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n220), .A2(G87), .ZN(new_n518));
  NOR3_X1   g0318(.A1(new_n410), .A2(new_n517), .A3(new_n518), .ZN(new_n519));
  NAND3_X1  g0319(.A1(new_n503), .A2(new_n220), .A3(G87), .ZN(new_n520));
  AOI21_X1  g0320(.A(new_n519), .B1(new_n520), .B2(KEYINPUT22), .ZN(new_n521));
  OAI21_X1  g0321(.A(KEYINPUT23), .B1(new_n220), .B2(G107), .ZN(new_n522));
  INV_X1    g0322(.A(KEYINPUT23), .ZN(new_n523));
  NAND3_X1  g0323(.A1(new_n523), .A2(new_n354), .A3(G20), .ZN(new_n524));
  NAND2_X1  g0324(.A1(G33), .A2(G116), .ZN(new_n525));
  OAI211_X1 g0325(.A(new_n522), .B(new_n524), .C1(G20), .C2(new_n525), .ZN(new_n526));
  INV_X1    g0326(.A(KEYINPUT86), .ZN(new_n527));
  XNOR2_X1  g0327(.A(new_n526), .B(new_n527), .ZN(new_n528));
  OAI21_X1  g0328(.A(KEYINPUT24), .B1(new_n521), .B2(new_n528), .ZN(new_n529));
  XNOR2_X1  g0329(.A(new_n526), .B(KEYINPUT86), .ZN(new_n530));
  INV_X1    g0330(.A(KEYINPUT24), .ZN(new_n531));
  INV_X1    g0331(.A(KEYINPUT22), .ZN(new_n532));
  AOI21_X1  g0332(.A(G20), .B1(new_n376), .B2(new_n377), .ZN(new_n533));
  AOI21_X1  g0333(.A(new_n532), .B1(new_n533), .B2(G87), .ZN(new_n534));
  OAI211_X1 g0334(.A(new_n530), .B(new_n531), .C1(new_n534), .C2(new_n519), .ZN(new_n535));
  AND2_X1   g0335(.A1(new_n529), .A2(new_n535), .ZN(new_n536));
  OAI211_X1 g0336(.A(new_n501), .B(new_n516), .C1(new_n536), .C2(new_n308), .ZN(new_n537));
  AND2_X1   g0337(.A1(new_n513), .A2(new_n502), .ZN(new_n538));
  NAND3_X1  g0338(.A1(new_n538), .A2(new_n276), .A3(new_n446), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n508), .A2(new_n322), .ZN(new_n540));
  AOI21_X1  g0340(.A(new_n308), .B1(new_n529), .B2(new_n535), .ZN(new_n541));
  INV_X1    g0341(.A(new_n501), .ZN(new_n542));
  OAI211_X1 g0342(.A(new_n539), .B(new_n540), .C1(new_n541), .C2(new_n542), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n537), .A2(new_n543), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n544), .A2(KEYINPUT87), .ZN(new_n545));
  INV_X1    g0345(.A(KEYINPUT87), .ZN(new_n546));
  NAND3_X1  g0346(.A1(new_n537), .A2(new_n543), .A3(new_n546), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n545), .A2(new_n547), .ZN(new_n548));
  NAND3_X1  g0348(.A1(new_n296), .A2(G45), .A3(new_n329), .ZN(new_n549));
  INV_X1    g0349(.A(G250), .ZN(new_n550));
  OAI21_X1  g0350(.A(new_n550), .B1(new_n259), .B2(new_n443), .ZN(new_n551));
  NAND3_X1  g0351(.A1(new_n549), .A2(new_n257), .A3(new_n551), .ZN(new_n552));
  INV_X1    g0352(.A(new_n552), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n323), .A2(G238), .ZN(new_n554));
  OAI21_X1  g0354(.A(KEYINPUT81), .B1(new_n384), .B2(new_n554), .ZN(new_n555));
  INV_X1    g0355(.A(KEYINPUT81), .ZN(new_n556));
  NAND4_X1  g0356(.A1(new_n503), .A2(new_n556), .A3(G238), .A4(new_n323), .ZN(new_n557));
  NAND3_X1  g0357(.A1(new_n503), .A2(G244), .A3(G1698), .ZN(new_n558));
  NAND4_X1  g0358(.A1(new_n555), .A2(new_n557), .A3(new_n525), .A4(new_n558), .ZN(new_n559));
  AOI21_X1  g0359(.A(new_n553), .B1(new_n559), .B2(new_n256), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n560), .A2(new_n276), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n559), .A2(new_n256), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n562), .A2(new_n552), .ZN(new_n563));
  XNOR2_X1  g0363(.A(new_n348), .B(KEYINPUT82), .ZN(new_n564));
  INV_X1    g0364(.A(new_n564), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n565), .A2(new_n472), .ZN(new_n566));
  NAND3_X1  g0366(.A1(new_n503), .A2(new_n220), .A3(G68), .ZN(new_n567));
  AOI21_X1  g0367(.A(KEYINPUT19), .B1(new_n317), .B2(G97), .ZN(new_n568));
  NAND3_X1  g0368(.A1(KEYINPUT19), .A2(G33), .A3(G97), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n569), .A2(new_n220), .ZN(new_n570));
  INV_X1    g0370(.A(G87), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n479), .A2(new_n571), .ZN(new_n572));
  AOI21_X1  g0372(.A(new_n568), .B1(new_n570), .B2(new_n572), .ZN(new_n573));
  AOI21_X1  g0373(.A(new_n308), .B1(new_n567), .B2(new_n573), .ZN(new_n574));
  INV_X1    g0374(.A(new_n293), .ZN(new_n575));
  AND2_X1   g0375(.A1(new_n575), .A2(new_n348), .ZN(new_n576));
  NOR2_X1   g0376(.A1(new_n574), .A2(new_n576), .ZN(new_n577));
  AOI22_X1  g0377(.A1(new_n563), .A2(new_n322), .B1(new_n566), .B2(new_n577), .ZN(new_n578));
  NOR2_X1   g0378(.A1(new_n471), .A2(new_n571), .ZN(new_n579));
  OR3_X1    g0379(.A1(new_n574), .A2(new_n576), .A3(new_n579), .ZN(new_n580));
  AOI21_X1  g0380(.A(new_n580), .B1(G190), .B2(new_n560), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n563), .A2(G200), .ZN(new_n582));
  AOI22_X1  g0382(.A1(new_n561), .A2(new_n578), .B1(new_n581), .B2(new_n582), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n505), .A2(new_n323), .ZN(new_n584));
  INV_X1    g0384(.A(G264), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n585), .A2(G1698), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n584), .A2(new_n586), .ZN(new_n587));
  AOI21_X1  g0387(.A(new_n587), .B1(new_n376), .B2(new_n377), .ZN(new_n588));
  INV_X1    g0388(.A(G303), .ZN(new_n589));
  NOR2_X1   g0389(.A1(new_n254), .A2(new_n589), .ZN(new_n590));
  OAI21_X1  g0390(.A(new_n256), .B1(new_n588), .B2(new_n590), .ZN(new_n591));
  OAI211_X1 g0391(.A(new_n257), .B(G270), .C1(new_n449), .C2(new_n450), .ZN(new_n592));
  NAND3_X1  g0392(.A1(new_n591), .A2(new_n446), .A3(new_n592), .ZN(new_n593));
  INV_X1    g0393(.A(G116), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n575), .A2(new_n594), .ZN(new_n595));
  NAND4_X1  g0395(.A1(new_n293), .A2(new_n308), .A3(new_n470), .A4(G116), .ZN(new_n596));
  AOI22_X1  g0396(.A1(new_n283), .A2(new_n219), .B1(G20), .B2(new_n594), .ZN(new_n597));
  OAI211_X1 g0397(.A(new_n464), .B(new_n220), .C1(G33), .C2(new_n474), .ZN(new_n598));
  AND3_X1   g0398(.A1(new_n597), .A2(KEYINPUT20), .A3(new_n598), .ZN(new_n599));
  AOI21_X1  g0399(.A(KEYINPUT20), .B1(new_n597), .B2(new_n598), .ZN(new_n600));
  OAI211_X1 g0400(.A(new_n595), .B(new_n596), .C1(new_n599), .C2(new_n600), .ZN(new_n601));
  NAND3_X1  g0401(.A1(new_n593), .A2(G169), .A3(new_n601), .ZN(new_n602));
  INV_X1    g0402(.A(KEYINPUT21), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  NAND4_X1  g0404(.A1(new_n593), .A2(KEYINPUT21), .A3(G169), .A4(new_n601), .ZN(new_n605));
  AND2_X1   g0405(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  AND3_X1   g0406(.A1(new_n591), .A2(new_n446), .A3(new_n592), .ZN(new_n607));
  NAND4_X1  g0407(.A1(new_n607), .A2(KEYINPUT83), .A3(G179), .A4(new_n601), .ZN(new_n608));
  INV_X1    g0408(.A(KEYINPUT83), .ZN(new_n609));
  NAND4_X1  g0409(.A1(new_n591), .A2(G179), .A3(new_n446), .A4(new_n592), .ZN(new_n610));
  INV_X1    g0410(.A(new_n601), .ZN(new_n611));
  OAI21_X1  g0411(.A(new_n609), .B1(new_n610), .B2(new_n611), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n608), .A2(new_n612), .ZN(new_n613));
  AOI21_X1  g0413(.A(new_n601), .B1(new_n593), .B2(G200), .ZN(new_n614));
  OAI21_X1  g0414(.A(new_n614), .B1(new_n514), .B2(new_n593), .ZN(new_n615));
  NAND3_X1  g0415(.A1(new_n606), .A2(new_n613), .A3(new_n615), .ZN(new_n616));
  INV_X1    g0416(.A(KEYINPUT84), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  NAND4_X1  g0418(.A1(new_n606), .A2(KEYINPUT84), .A3(new_n613), .A4(new_n615), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  AND4_X1   g0420(.A1(new_n497), .A2(new_n548), .A3(new_n583), .A4(new_n620), .ZN(new_n621));
  AND2_X1   g0421(.A1(new_n435), .A2(new_n621), .ZN(G372));
  INV_X1    g0422(.A(new_n337), .ZN(new_n623));
  AND3_X1   g0423(.A1(new_n393), .A2(new_n426), .A3(new_n418), .ZN(new_n624));
  AOI21_X1  g0424(.A(new_n426), .B1(new_n393), .B2(new_n418), .ZN(new_n625));
  NOR2_X1   g0425(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n302), .A2(new_n303), .ZN(new_n627));
  INV_X1    g0427(.A(new_n366), .ZN(new_n628));
  AOI21_X1  g0428(.A(new_n301), .B1(new_n627), .B2(new_n628), .ZN(new_n629));
  AND2_X1   g0429(.A1(new_n425), .A2(new_n431), .ZN(new_n630));
  INV_X1    g0430(.A(new_n630), .ZN(new_n631));
  OAI21_X1  g0431(.A(new_n626), .B1(new_n629), .B2(new_n631), .ZN(new_n632));
  AOI21_X1  g0432(.A(new_n623), .B1(new_n632), .B2(new_n342), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n488), .A2(new_n493), .ZN(new_n634));
  INV_X1    g0434(.A(new_n516), .ZN(new_n635));
  NOR3_X1   g0435(.A1(new_n635), .A2(new_n541), .A3(new_n542), .ZN(new_n636));
  AND3_X1   g0436(.A1(new_n613), .A2(new_n604), .A3(new_n605), .ZN(new_n637));
  AOI21_X1  g0437(.A(new_n636), .B1(new_n637), .B2(new_n543), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n494), .A2(new_n496), .ZN(new_n639));
  NAND4_X1  g0439(.A1(new_n634), .A2(new_n638), .A3(new_n639), .A4(new_n583), .ZN(new_n640));
  INV_X1    g0440(.A(new_n640), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n578), .A2(new_n561), .ZN(new_n642));
  INV_X1    g0442(.A(new_n642), .ZN(new_n643));
  NOR3_X1   g0443(.A1(new_n574), .A2(new_n576), .A3(new_n579), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n560), .A2(G190), .ZN(new_n645));
  NAND3_X1  g0445(.A1(new_n582), .A2(new_n644), .A3(new_n645), .ZN(new_n646));
  NAND4_X1  g0446(.A1(new_n642), .A2(new_n646), .A3(new_n494), .A4(new_n496), .ZN(new_n647));
  AOI21_X1  g0447(.A(new_n643), .B1(new_n647), .B2(KEYINPUT26), .ZN(new_n648));
  AOI211_X1 g0448(.A(G179), .B(new_n491), .C1(new_n454), .C2(new_n458), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n495), .A2(new_n322), .ZN(new_n650));
  INV_X1    g0450(.A(new_n486), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  OAI21_X1  g0452(.A(KEYINPUT88), .B1(new_n649), .B2(new_n652), .ZN(new_n653));
  INV_X1    g0453(.A(KEYINPUT26), .ZN(new_n654));
  INV_X1    g0454(.A(KEYINPUT88), .ZN(new_n655));
  NAND3_X1  g0455(.A1(new_n494), .A2(new_n655), .A3(new_n496), .ZN(new_n656));
  NAND4_X1  g0456(.A1(new_n583), .A2(new_n653), .A3(new_n654), .A4(new_n656), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n648), .A2(new_n657), .ZN(new_n658));
  OAI21_X1  g0458(.A(new_n435), .B1(new_n641), .B2(new_n658), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n633), .A2(new_n659), .ZN(G369));
  INV_X1    g0460(.A(G13), .ZN(new_n661));
  NOR2_X1   g0461(.A1(new_n661), .A2(G20), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n296), .A2(new_n662), .ZN(new_n663));
  OR2_X1    g0463(.A1(new_n663), .A2(KEYINPUT27), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n663), .A2(KEYINPUT27), .ZN(new_n665));
  NAND3_X1  g0465(.A1(new_n664), .A2(G213), .A3(new_n665), .ZN(new_n666));
  INV_X1    g0466(.A(G343), .ZN(new_n667));
  NOR2_X1   g0467(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  OAI21_X1  g0468(.A(new_n668), .B1(new_n541), .B2(new_n542), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n548), .A2(new_n669), .ZN(new_n670));
  INV_X1    g0470(.A(KEYINPUT90), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  NAND3_X1  g0472(.A1(new_n548), .A2(KEYINPUT90), .A3(new_n669), .ZN(new_n673));
  AND2_X1   g0473(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  INV_X1    g0474(.A(new_n668), .ZN(new_n675));
  OR2_X1    g0475(.A1(new_n543), .A2(new_n675), .ZN(new_n676));
  INV_X1    g0476(.A(new_n676), .ZN(new_n677));
  NOR2_X1   g0477(.A1(new_n674), .A2(new_n677), .ZN(new_n678));
  OAI21_X1  g0478(.A(new_n620), .B1(new_n611), .B2(new_n675), .ZN(new_n679));
  INV_X1    g0479(.A(new_n637), .ZN(new_n680));
  NAND3_X1  g0480(.A1(new_n680), .A2(new_n601), .A3(new_n668), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n679), .A2(new_n681), .ZN(new_n682));
  XNOR2_X1  g0482(.A(KEYINPUT89), .B(G330), .ZN(new_n683));
  INV_X1    g0483(.A(new_n683), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n682), .A2(new_n684), .ZN(new_n685));
  NOR2_X1   g0485(.A1(new_n678), .A2(new_n685), .ZN(new_n686));
  NOR2_X1   g0486(.A1(new_n637), .A2(new_n668), .ZN(new_n687));
  NAND3_X1  g0487(.A1(new_n672), .A2(new_n673), .A3(new_n687), .ZN(new_n688));
  OR2_X1    g0488(.A1(new_n543), .A2(new_n668), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  OR2_X1    g0490(.A1(new_n686), .A2(new_n690), .ZN(G399));
  INV_X1    g0491(.A(new_n223), .ZN(new_n692));
  NOR2_X1   g0492(.A1(new_n692), .A2(G41), .ZN(new_n693));
  INV_X1    g0493(.A(new_n693), .ZN(new_n694));
  NOR2_X1   g0494(.A1(new_n572), .A2(G116), .ZN(new_n695));
  NAND3_X1  g0495(.A1(new_n694), .A2(G1), .A3(new_n695), .ZN(new_n696));
  OAI21_X1  g0496(.A(new_n696), .B1(new_n217), .B2(new_n694), .ZN(new_n697));
  XNOR2_X1  g0497(.A(new_n697), .B(KEYINPUT28), .ZN(new_n698));
  INV_X1    g0498(.A(KEYINPUT94), .ZN(new_n699));
  AND2_X1   g0499(.A1(new_n648), .A2(new_n657), .ZN(new_n700));
  AOI21_X1  g0500(.A(new_n668), .B1(new_n700), .B2(new_n640), .ZN(new_n701));
  OAI21_X1  g0501(.A(new_n699), .B1(new_n701), .B2(KEYINPUT29), .ZN(new_n702));
  NAND3_X1  g0502(.A1(new_n583), .A2(new_n653), .A3(new_n656), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n703), .A2(KEYINPUT26), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n645), .A2(new_n644), .ZN(new_n705));
  NOR2_X1   g0505(.A1(new_n560), .A2(new_n421), .ZN(new_n706));
  NAND2_X1  g0506(.A1(new_n577), .A2(new_n566), .ZN(new_n707));
  OAI21_X1  g0507(.A(new_n707), .B1(new_n560), .B2(G169), .ZN(new_n708));
  AND2_X1   g0508(.A1(new_n560), .A2(new_n276), .ZN(new_n709));
  OAI22_X1  g0509(.A1(new_n705), .A2(new_n706), .B1(new_n708), .B2(new_n709), .ZN(new_n710));
  NOR2_X1   g0510(.A1(new_n710), .A2(new_n639), .ZN(new_n711));
  AOI21_X1  g0511(.A(new_n643), .B1(new_n711), .B2(new_n654), .ZN(new_n712));
  NAND3_X1  g0512(.A1(new_n640), .A2(new_n704), .A3(new_n712), .ZN(new_n713));
  NAND3_X1  g0513(.A1(new_n713), .A2(KEYINPUT29), .A3(new_n675), .ZN(new_n714));
  OAI21_X1  g0514(.A(new_n675), .B1(new_n641), .B2(new_n658), .ZN(new_n715));
  INV_X1    g0515(.A(KEYINPUT29), .ZN(new_n716));
  NAND3_X1  g0516(.A1(new_n715), .A2(KEYINPUT94), .A3(new_n716), .ZN(new_n717));
  NAND3_X1  g0517(.A1(new_n702), .A2(new_n714), .A3(new_n717), .ZN(new_n718));
  AOI22_X1  g0518(.A1(new_n545), .A2(new_n547), .B1(new_n618), .B2(new_n619), .ZN(new_n719));
  NAND4_X1  g0519(.A1(new_n719), .A2(new_n497), .A3(new_n583), .A4(new_n675), .ZN(new_n720));
  NAND2_X1  g0520(.A1(new_n560), .A2(new_n538), .ZN(new_n721));
  NAND2_X1  g0521(.A1(new_n721), .A2(KEYINPUT92), .ZN(new_n722));
  NOR2_X1   g0522(.A1(new_n495), .A2(new_n610), .ZN(new_n723));
  INV_X1    g0523(.A(KEYINPUT92), .ZN(new_n724));
  NAND3_X1  g0524(.A1(new_n560), .A2(new_n724), .A3(new_n538), .ZN(new_n725));
  NAND4_X1  g0525(.A1(new_n722), .A2(new_n723), .A3(KEYINPUT30), .A4(new_n725), .ZN(new_n726));
  INV_X1    g0526(.A(KEYINPUT93), .ZN(new_n727));
  NAND2_X1  g0527(.A1(new_n726), .A2(new_n727), .ZN(new_n728));
  NAND3_X1  g0528(.A1(new_n722), .A2(new_n723), .A3(new_n725), .ZN(new_n729));
  INV_X1    g0529(.A(KEYINPUT30), .ZN(new_n730));
  NAND2_X1  g0530(.A1(new_n729), .A2(new_n730), .ZN(new_n731));
  AOI21_X1  g0531(.A(new_n724), .B1(new_n560), .B2(new_n538), .ZN(new_n732));
  NOR2_X1   g0532(.A1(new_n452), .A2(new_n453), .ZN(new_n733));
  NAND4_X1  g0533(.A1(new_n733), .A2(G179), .A3(new_n467), .A4(new_n607), .ZN(new_n734));
  NOR2_X1   g0534(.A1(new_n732), .A2(new_n734), .ZN(new_n735));
  NAND4_X1  g0535(.A1(new_n735), .A2(KEYINPUT93), .A3(KEYINPUT30), .A4(new_n725), .ZN(new_n736));
  NAND4_X1  g0536(.A1(new_n563), .A2(new_n276), .A3(new_n508), .A4(new_n593), .ZN(new_n737));
  OR2_X1    g0537(.A1(new_n737), .A2(new_n492), .ZN(new_n738));
  NAND4_X1  g0538(.A1(new_n728), .A2(new_n731), .A3(new_n736), .A4(new_n738), .ZN(new_n739));
  NAND2_X1  g0539(.A1(new_n739), .A2(new_n668), .ZN(new_n740));
  INV_X1    g0540(.A(KEYINPUT31), .ZN(new_n741));
  NAND2_X1  g0541(.A1(new_n740), .A2(new_n741), .ZN(new_n742));
  XOR2_X1   g0542(.A(KEYINPUT91), .B(KEYINPUT31), .Z(new_n743));
  INV_X1    g0543(.A(new_n743), .ZN(new_n744));
  NAND3_X1  g0544(.A1(new_n739), .A2(new_n668), .A3(new_n744), .ZN(new_n745));
  NAND3_X1  g0545(.A1(new_n720), .A2(new_n742), .A3(new_n745), .ZN(new_n746));
  NAND2_X1  g0546(.A1(new_n746), .A2(new_n684), .ZN(new_n747));
  NAND2_X1  g0547(.A1(new_n718), .A2(new_n747), .ZN(new_n748));
  INV_X1    g0548(.A(new_n748), .ZN(new_n749));
  OAI21_X1  g0549(.A(new_n698), .B1(new_n749), .B2(G1), .ZN(G364));
  AOI21_X1  g0550(.A(new_n250), .B1(new_n662), .B2(G45), .ZN(new_n751));
  INV_X1    g0551(.A(new_n751), .ZN(new_n752));
  OAI21_X1  g0552(.A(new_n685), .B1(new_n693), .B2(new_n752), .ZN(new_n753));
  INV_X1    g0553(.A(new_n682), .ZN(new_n754));
  AOI21_X1  g0554(.A(new_n753), .B1(new_n683), .B2(new_n754), .ZN(new_n755));
  AOI21_X1  g0555(.A(new_n219), .B1(G20), .B2(new_n322), .ZN(new_n756));
  INV_X1    g0556(.A(new_n756), .ZN(new_n757));
  NOR2_X1   g0557(.A1(new_n220), .A2(G190), .ZN(new_n758));
  INV_X1    g0558(.A(KEYINPUT99), .ZN(new_n759));
  XNOR2_X1  g0559(.A(new_n758), .B(new_n759), .ZN(new_n760));
  NOR3_X1   g0560(.A1(new_n760), .A2(G179), .A3(new_n421), .ZN(new_n761));
  OR2_X1    g0561(.A1(new_n761), .A2(KEYINPUT100), .ZN(new_n762));
  NAND2_X1  g0562(.A1(new_n761), .A2(KEYINPUT100), .ZN(new_n763));
  NAND2_X1  g0563(.A1(new_n762), .A2(new_n763), .ZN(new_n764));
  INV_X1    g0564(.A(new_n764), .ZN(new_n765));
  NAND2_X1  g0565(.A1(new_n765), .A2(G107), .ZN(new_n766));
  NOR3_X1   g0566(.A1(new_n760), .A2(G179), .A3(G200), .ZN(new_n767));
  NAND2_X1  g0567(.A1(new_n767), .A2(G159), .ZN(new_n768));
  XOR2_X1   g0568(.A(new_n768), .B(KEYINPUT32), .Z(new_n769));
  NOR2_X1   g0569(.A1(G179), .A2(G200), .ZN(new_n770));
  AOI21_X1  g0570(.A(new_n220), .B1(new_n770), .B2(G190), .ZN(new_n771));
  NOR2_X1   g0571(.A1(new_n771), .A2(new_n474), .ZN(new_n772));
  NAND3_X1  g0572(.A1(G20), .A2(G179), .A3(G200), .ZN(new_n773));
  NOR2_X1   g0573(.A1(new_n773), .A2(new_n514), .ZN(new_n774));
  INV_X1    g0574(.A(new_n774), .ZN(new_n775));
  NOR2_X1   g0575(.A1(new_n775), .A2(new_n202), .ZN(new_n776));
  NOR2_X1   g0576(.A1(new_n773), .A2(G190), .ZN(new_n777));
  AOI211_X1 g0577(.A(new_n772), .B(new_n776), .C1(G68), .C2(new_n777), .ZN(new_n778));
  NOR2_X1   g0578(.A1(new_n276), .A2(G200), .ZN(new_n779));
  NAND2_X1  g0579(.A1(new_n758), .A2(new_n779), .ZN(new_n780));
  NOR2_X1   g0580(.A1(new_n220), .A2(new_n514), .ZN(new_n781));
  NAND3_X1  g0581(.A1(new_n781), .A2(new_n276), .A3(G200), .ZN(new_n782));
  OAI221_X1 g0582(.A(new_n254), .B1(new_n780), .B2(new_n280), .C1(new_n782), .C2(new_n571), .ZN(new_n783));
  NAND2_X1  g0583(.A1(new_n781), .A2(new_n779), .ZN(new_n784));
  NAND2_X1  g0584(.A1(new_n784), .A2(KEYINPUT98), .ZN(new_n785));
  INV_X1    g0585(.A(new_n785), .ZN(new_n786));
  NOR2_X1   g0586(.A1(new_n784), .A2(KEYINPUT98), .ZN(new_n787));
  NOR2_X1   g0587(.A1(new_n786), .A2(new_n787), .ZN(new_n788));
  INV_X1    g0588(.A(new_n788), .ZN(new_n789));
  AOI21_X1  g0589(.A(new_n783), .B1(new_n789), .B2(new_n314), .ZN(new_n790));
  NAND4_X1  g0590(.A1(new_n766), .A2(new_n769), .A3(new_n778), .A4(new_n790), .ZN(new_n791));
  NAND2_X1  g0591(.A1(new_n765), .A2(G283), .ZN(new_n792));
  INV_X1    g0592(.A(new_n777), .ZN(new_n793));
  XOR2_X1   g0593(.A(KEYINPUT33), .B(G317), .Z(new_n794));
  INV_X1    g0594(.A(G326), .ZN(new_n795));
  OAI22_X1  g0595(.A1(new_n793), .A2(new_n794), .B1(new_n775), .B2(new_n795), .ZN(new_n796));
  INV_X1    g0596(.A(new_n771), .ZN(new_n797));
  AOI21_X1  g0597(.A(new_n796), .B1(G294), .B2(new_n797), .ZN(new_n798));
  NAND2_X1  g0598(.A1(new_n767), .A2(G329), .ZN(new_n799));
  INV_X1    g0599(.A(G311), .ZN(new_n800));
  OAI221_X1 g0600(.A(new_n410), .B1(new_n780), .B2(new_n800), .C1(new_n782), .C2(new_n589), .ZN(new_n801));
  AOI21_X1  g0601(.A(new_n801), .B1(new_n789), .B2(G322), .ZN(new_n802));
  NAND4_X1  g0602(.A1(new_n792), .A2(new_n798), .A3(new_n799), .A4(new_n802), .ZN(new_n803));
  AOI21_X1  g0603(.A(new_n757), .B1(new_n791), .B2(new_n803), .ZN(new_n804));
  NAND3_X1  g0604(.A1(new_n661), .A2(new_n316), .A3(KEYINPUT96), .ZN(new_n805));
  INV_X1    g0605(.A(KEYINPUT96), .ZN(new_n806));
  OAI21_X1  g0606(.A(new_n806), .B1(G13), .B2(G33), .ZN(new_n807));
  NAND2_X1  g0607(.A1(new_n805), .A2(new_n807), .ZN(new_n808));
  NAND2_X1  g0608(.A1(new_n808), .A2(new_n220), .ZN(new_n809));
  XOR2_X1   g0609(.A(new_n809), .B(KEYINPUT97), .Z(new_n810));
  INV_X1    g0610(.A(new_n810), .ZN(new_n811));
  NOR2_X1   g0611(.A1(new_n811), .A2(new_n756), .ZN(new_n812));
  NOR2_X1   g0612(.A1(new_n503), .A2(new_n692), .ZN(new_n813));
  INV_X1    g0613(.A(new_n813), .ZN(new_n814));
  NOR2_X1   g0614(.A1(new_n245), .A2(new_n443), .ZN(new_n815));
  AOI211_X1 g0615(.A(new_n814), .B(new_n815), .C1(new_n218), .C2(new_n247), .ZN(new_n816));
  NOR2_X1   g0616(.A1(new_n692), .A2(new_n410), .ZN(new_n817));
  AOI22_X1  g0617(.A1(new_n817), .A2(G355), .B1(new_n594), .B2(new_n692), .ZN(new_n818));
  XOR2_X1   g0618(.A(new_n818), .B(KEYINPUT95), .Z(new_n819));
  OAI21_X1  g0619(.A(new_n812), .B1(new_n816), .B2(new_n819), .ZN(new_n820));
  NOR2_X1   g0620(.A1(new_n693), .A2(new_n752), .ZN(new_n821));
  NAND2_X1  g0621(.A1(new_n820), .A2(new_n821), .ZN(new_n822));
  AOI211_X1 g0622(.A(new_n804), .B(new_n822), .C1(new_n754), .C2(new_n811), .ZN(new_n823));
  NOR2_X1   g0623(.A1(new_n755), .A2(new_n823), .ZN(new_n824));
  INV_X1    g0624(.A(new_n824), .ZN(G396));
  NOR2_X1   g0625(.A1(new_n366), .A2(new_n668), .ZN(new_n826));
  NAND2_X1  g0626(.A1(new_n351), .A2(new_n668), .ZN(new_n827));
  XNOR2_X1  g0627(.A(new_n827), .B(KEYINPUT103), .ZN(new_n828));
  NAND2_X1  g0628(.A1(new_n828), .A2(new_n363), .ZN(new_n829));
  AOI21_X1  g0629(.A(new_n826), .B1(new_n829), .B2(new_n366), .ZN(new_n830));
  INV_X1    g0630(.A(new_n830), .ZN(new_n831));
  NAND2_X1  g0631(.A1(new_n715), .A2(new_n831), .ZN(new_n832));
  OAI211_X1 g0632(.A(new_n675), .B(new_n830), .C1(new_n641), .C2(new_n658), .ZN(new_n833));
  NAND2_X1  g0633(.A1(new_n832), .A2(new_n833), .ZN(new_n834));
  AOI21_X1  g0634(.A(new_n821), .B1(new_n834), .B2(new_n747), .ZN(new_n835));
  OAI21_X1  g0635(.A(new_n835), .B1(new_n747), .B2(new_n834), .ZN(new_n836));
  INV_X1    g0636(.A(new_n808), .ZN(new_n837));
  NAND2_X1  g0637(.A1(new_n837), .A2(new_n757), .ZN(new_n838));
  OAI21_X1  g0638(.A(new_n821), .B1(G77), .B2(new_n838), .ZN(new_n839));
  NAND2_X1  g0639(.A1(new_n765), .A2(G87), .ZN(new_n840));
  NOR2_X1   g0640(.A1(new_n775), .A2(new_n589), .ZN(new_n841));
  AOI211_X1 g0641(.A(new_n772), .B(new_n841), .C1(G283), .C2(new_n777), .ZN(new_n842));
  NAND2_X1  g0642(.A1(new_n789), .A2(G294), .ZN(new_n843));
  OAI221_X1 g0643(.A(new_n410), .B1(new_n780), .B2(new_n594), .C1(new_n782), .C2(new_n354), .ZN(new_n844));
  AOI21_X1  g0644(.A(new_n844), .B1(new_n767), .B2(G311), .ZN(new_n845));
  NAND4_X1  g0645(.A1(new_n840), .A2(new_n842), .A3(new_n843), .A4(new_n845), .ZN(new_n846));
  NAND2_X1  g0646(.A1(new_n765), .A2(G68), .ZN(new_n847));
  INV_X1    g0647(.A(new_n780), .ZN(new_n848));
  AOI22_X1  g0648(.A1(new_n848), .A2(G159), .B1(G137), .B2(new_n774), .ZN(new_n849));
  INV_X1    g0649(.A(G150), .ZN(new_n850));
  INV_X1    g0650(.A(G143), .ZN(new_n851));
  OAI221_X1 g0651(.A(new_n849), .B1(new_n850), .B2(new_n793), .C1(new_n788), .C2(new_n851), .ZN(new_n852));
  XOR2_X1   g0652(.A(KEYINPUT101), .B(KEYINPUT34), .Z(new_n853));
  XNOR2_X1  g0653(.A(new_n853), .B(KEYINPUT102), .ZN(new_n854));
  INV_X1    g0654(.A(new_n854), .ZN(new_n855));
  NAND2_X1  g0655(.A1(new_n852), .A2(new_n855), .ZN(new_n856));
  OAI221_X1 g0656(.A(new_n503), .B1(new_n394), .B2(new_n771), .C1(new_n202), .C2(new_n782), .ZN(new_n857));
  AOI21_X1  g0657(.A(new_n857), .B1(G132), .B2(new_n767), .ZN(new_n858));
  NAND3_X1  g0658(.A1(new_n847), .A2(new_n856), .A3(new_n858), .ZN(new_n859));
  NOR2_X1   g0659(.A1(new_n852), .A2(new_n855), .ZN(new_n860));
  OAI21_X1  g0660(.A(new_n846), .B1(new_n859), .B2(new_n860), .ZN(new_n861));
  AOI21_X1  g0661(.A(new_n839), .B1(new_n861), .B2(new_n756), .ZN(new_n862));
  OAI21_X1  g0662(.A(new_n862), .B1(new_n830), .B2(new_n837), .ZN(new_n863));
  AND2_X1   g0663(.A1(new_n836), .A2(new_n863), .ZN(new_n864));
  INV_X1    g0664(.A(new_n864), .ZN(G384));
  OR2_X1    g0665(.A1(new_n482), .A2(KEYINPUT35), .ZN(new_n866));
  NAND2_X1  g0666(.A1(new_n482), .A2(KEYINPUT35), .ZN(new_n867));
  NAND4_X1  g0667(.A1(new_n866), .A2(G116), .A3(new_n221), .A4(new_n867), .ZN(new_n868));
  XOR2_X1   g0668(.A(new_n868), .B(KEYINPUT36), .Z(new_n869));
  OAI211_X1 g0669(.A(new_n218), .B(G77), .C1(new_n241), .C2(new_n394), .ZN(new_n870));
  AOI211_X1 g0670(.A(G13), .B(new_n296), .C1(new_n870), .C2(new_n240), .ZN(new_n871));
  NOR2_X1   g0671(.A1(new_n869), .A2(new_n871), .ZN(new_n872));
  OAI211_X1 g0672(.A(new_n299), .B(new_n668), .C1(new_n304), .C2(new_n277), .ZN(new_n873));
  NAND2_X1  g0673(.A1(new_n299), .A2(new_n668), .ZN(new_n874));
  NAND3_X1  g0674(.A1(new_n300), .A2(new_n627), .A3(new_n874), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n873), .A2(new_n875), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n876), .A2(new_n830), .ZN(new_n877));
  AOI21_X1  g0677(.A(new_n744), .B1(new_n739), .B2(new_n668), .ZN(new_n878));
  AOI21_X1  g0678(.A(new_n878), .B1(new_n621), .B2(new_n675), .ZN(new_n879));
  OAI21_X1  g0679(.A(KEYINPUT109), .B1(new_n740), .B2(new_n741), .ZN(new_n880));
  INV_X1    g0680(.A(KEYINPUT109), .ZN(new_n881));
  NAND4_X1  g0681(.A1(new_n739), .A2(new_n881), .A3(KEYINPUT31), .A4(new_n668), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n880), .A2(new_n882), .ZN(new_n883));
  AOI21_X1  g0683(.A(new_n877), .B1(new_n879), .B2(new_n883), .ZN(new_n884));
  INV_X1    g0684(.A(KEYINPUT107), .ZN(new_n885));
  INV_X1    g0685(.A(new_n422), .ZN(new_n886));
  NAND4_X1  g0686(.A1(new_n886), .A2(new_n414), .A3(new_n417), .A4(new_n429), .ZN(new_n887));
  INV_X1    g0687(.A(new_n417), .ZN(new_n888));
  OAI21_X1  g0688(.A(new_n396), .B1(new_n401), .B2(new_n403), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n889), .A2(KEYINPUT105), .ZN(new_n890));
  INV_X1    g0690(.A(KEYINPUT105), .ZN(new_n891));
  OAI211_X1 g0691(.A(new_n891), .B(new_n396), .C1(new_n401), .C2(new_n403), .ZN(new_n892));
  NAND3_X1  g0692(.A1(new_n890), .A2(new_n405), .A3(new_n892), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n404), .A2(new_n284), .ZN(new_n894));
  INV_X1    g0694(.A(new_n894), .ZN(new_n895));
  AOI21_X1  g0695(.A(new_n888), .B1(new_n893), .B2(new_n895), .ZN(new_n896));
  AOI21_X1  g0696(.A(new_n322), .B1(new_n386), .B2(new_n388), .ZN(new_n897));
  AOI21_X1  g0697(.A(new_n897), .B1(G179), .B2(new_n392), .ZN(new_n898));
  OAI21_X1  g0698(.A(new_n887), .B1(new_n896), .B2(new_n898), .ZN(new_n899));
  NOR2_X1   g0699(.A1(new_n896), .A2(new_n666), .ZN(new_n900));
  OAI21_X1  g0700(.A(KEYINPUT37), .B1(new_n899), .B2(new_n900), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n419), .A2(KEYINPUT106), .ZN(new_n902));
  AOI21_X1  g0702(.A(KEYINPUT37), .B1(new_n423), .B2(new_n424), .ZN(new_n903));
  INV_X1    g0703(.A(new_n666), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n418), .A2(new_n904), .ZN(new_n905));
  INV_X1    g0705(.A(KEYINPUT106), .ZN(new_n906));
  NAND3_X1  g0706(.A1(new_n393), .A2(new_n906), .A3(new_n418), .ZN(new_n907));
  NAND4_X1  g0707(.A1(new_n902), .A2(new_n903), .A3(new_n905), .A4(new_n907), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n901), .A2(new_n908), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n432), .A2(new_n900), .ZN(new_n910));
  AND3_X1   g0710(.A1(new_n909), .A2(KEYINPUT38), .A3(new_n910), .ZN(new_n911));
  AOI21_X1  g0711(.A(KEYINPUT38), .B1(new_n909), .B2(new_n910), .ZN(new_n912));
  OAI21_X1  g0712(.A(new_n885), .B1(new_n911), .B2(new_n912), .ZN(new_n913));
  INV_X1    g0713(.A(KEYINPUT38), .ZN(new_n914));
  INV_X1    g0714(.A(KEYINPUT37), .ZN(new_n915));
  AND3_X1   g0715(.A1(new_n887), .A2(new_n905), .A3(new_n915), .ZN(new_n916));
  INV_X1    g0716(.A(new_n907), .ZN(new_n917));
  AOI21_X1  g0717(.A(new_n906), .B1(new_n393), .B2(new_n418), .ZN(new_n918));
  NOR2_X1   g0718(.A1(new_n917), .A2(new_n918), .ZN(new_n919));
  AOI21_X1  g0719(.A(KEYINPUT16), .B1(new_n889), .B2(KEYINPUT105), .ZN(new_n920));
  AOI21_X1  g0720(.A(new_n894), .B1(new_n920), .B2(new_n892), .ZN(new_n921));
  OAI21_X1  g0721(.A(new_n904), .B1(new_n921), .B2(new_n888), .ZN(new_n922));
  OAI21_X1  g0722(.A(new_n393), .B1(new_n921), .B2(new_n888), .ZN(new_n923));
  NAND3_X1  g0723(.A1(new_n922), .A2(new_n923), .A3(new_n887), .ZN(new_n924));
  AOI22_X1  g0724(.A1(new_n916), .A2(new_n919), .B1(new_n924), .B2(KEYINPUT37), .ZN(new_n925));
  AOI21_X1  g0725(.A(new_n922), .B1(new_n630), .B2(new_n626), .ZN(new_n926));
  OAI21_X1  g0726(.A(new_n914), .B1(new_n925), .B2(new_n926), .ZN(new_n927));
  NAND3_X1  g0727(.A1(new_n909), .A2(KEYINPUT38), .A3(new_n910), .ZN(new_n928));
  NAND3_X1  g0728(.A1(new_n927), .A2(KEYINPUT107), .A3(new_n928), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n913), .A2(new_n929), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n884), .A2(new_n930), .ZN(new_n931));
  INV_X1    g0731(.A(KEYINPUT40), .ZN(new_n932));
  INV_X1    g0732(.A(KEYINPUT108), .ZN(new_n933));
  NAND3_X1  g0733(.A1(new_n419), .A2(new_n887), .A3(new_n905), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n934), .A2(KEYINPUT37), .ZN(new_n935));
  INV_X1    g0735(.A(new_n905), .ZN(new_n936));
  AOI22_X1  g0736(.A1(new_n908), .A2(new_n935), .B1(new_n432), .B2(new_n936), .ZN(new_n937));
  OAI21_X1  g0737(.A(new_n933), .B1(new_n937), .B2(KEYINPUT38), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n908), .A2(new_n935), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n432), .A2(new_n936), .ZN(new_n940));
  NAND2_X1  g0740(.A1(new_n939), .A2(new_n940), .ZN(new_n941));
  NAND3_X1  g0741(.A1(new_n941), .A2(KEYINPUT108), .A3(new_n914), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n938), .A2(new_n942), .ZN(new_n943));
  AOI21_X1  g0743(.A(new_n932), .B1(new_n943), .B2(new_n928), .ZN(new_n944));
  AOI22_X1  g0744(.A1(new_n931), .A2(new_n932), .B1(new_n884), .B2(new_n944), .ZN(new_n945));
  INV_X1    g0745(.A(new_n945), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n879), .A2(new_n883), .ZN(new_n947));
  INV_X1    g0747(.A(new_n947), .ZN(new_n948));
  OAI21_X1  g0748(.A(new_n946), .B1(new_n434), .B2(new_n948), .ZN(new_n949));
  NAND3_X1  g0749(.A1(new_n945), .A2(new_n435), .A3(new_n947), .ZN(new_n950));
  NAND3_X1  g0750(.A1(new_n949), .A2(new_n684), .A3(new_n950), .ZN(new_n951));
  NOR2_X1   g0751(.A1(new_n626), .A2(new_n904), .ZN(new_n952));
  AOI22_X1  g0752(.A1(new_n901), .A2(new_n908), .B1(new_n432), .B2(new_n900), .ZN(new_n953));
  AOI21_X1  g0753(.A(KEYINPUT39), .B1(new_n953), .B2(KEYINPUT38), .ZN(new_n954));
  AOI21_X1  g0754(.A(KEYINPUT108), .B1(new_n941), .B2(new_n914), .ZN(new_n955));
  AOI211_X1 g0755(.A(new_n933), .B(KEYINPUT38), .C1(new_n939), .C2(new_n940), .ZN(new_n956));
  OAI21_X1  g0756(.A(new_n954), .B1(new_n955), .B2(new_n956), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n927), .A2(new_n928), .ZN(new_n958));
  NAND2_X1  g0758(.A1(new_n958), .A2(KEYINPUT39), .ZN(new_n959));
  NAND2_X1  g0759(.A1(new_n957), .A2(new_n959), .ZN(new_n960));
  NOR2_X1   g0760(.A1(new_n300), .A2(new_n668), .ZN(new_n961));
  AOI21_X1  g0761(.A(new_n952), .B1(new_n960), .B2(new_n961), .ZN(new_n962));
  INV_X1    g0762(.A(new_n876), .ZN(new_n963));
  INV_X1    g0763(.A(KEYINPUT104), .ZN(new_n964));
  XNOR2_X1  g0764(.A(new_n826), .B(new_n964), .ZN(new_n965));
  INV_X1    g0765(.A(new_n965), .ZN(new_n966));
  AOI21_X1  g0766(.A(new_n963), .B1(new_n833), .B2(new_n966), .ZN(new_n967));
  NAND2_X1  g0767(.A1(new_n967), .A2(new_n930), .ZN(new_n968));
  NAND2_X1  g0768(.A1(new_n962), .A2(new_n968), .ZN(new_n969));
  NAND4_X1  g0769(.A1(new_n702), .A2(new_n435), .A3(new_n714), .A4(new_n717), .ZN(new_n970));
  NAND2_X1  g0770(.A1(new_n970), .A2(new_n633), .ZN(new_n971));
  XNOR2_X1  g0771(.A(new_n969), .B(new_n971), .ZN(new_n972));
  NAND2_X1  g0772(.A1(new_n951), .A2(new_n972), .ZN(new_n973));
  OAI21_X1  g0773(.A(new_n973), .B1(new_n296), .B2(new_n662), .ZN(new_n974));
  NOR2_X1   g0774(.A1(new_n951), .A2(new_n972), .ZN(new_n975));
  OAI21_X1  g0775(.A(new_n872), .B1(new_n974), .B2(new_n975), .ZN(G367));
  OAI21_X1  g0776(.A(new_n497), .B1(new_n486), .B2(new_n675), .ZN(new_n977));
  NAND3_X1  g0777(.A1(new_n494), .A2(new_n496), .A3(new_n668), .ZN(new_n978));
  AND2_X1   g0778(.A1(new_n977), .A2(new_n978), .ZN(new_n979));
  OR2_X1    g0779(.A1(new_n688), .A2(new_n979), .ZN(new_n980));
  OR2_X1    g0780(.A1(new_n980), .A2(KEYINPUT42), .ZN(new_n981));
  OR2_X1    g0781(.A1(new_n977), .A2(new_n543), .ZN(new_n982));
  AOI21_X1  g0782(.A(new_n668), .B1(new_n982), .B2(new_n639), .ZN(new_n983));
  AOI21_X1  g0783(.A(new_n983), .B1(new_n980), .B2(KEYINPUT42), .ZN(new_n984));
  NAND2_X1  g0784(.A1(new_n981), .A2(new_n984), .ZN(new_n985));
  NOR2_X1   g0785(.A1(new_n675), .A2(new_n644), .ZN(new_n986));
  NAND2_X1  g0786(.A1(new_n643), .A2(new_n986), .ZN(new_n987));
  OR2_X1    g0787(.A1(new_n987), .A2(KEYINPUT110), .ZN(new_n988));
  NOR2_X1   g0788(.A1(new_n710), .A2(new_n986), .ZN(new_n989));
  NAND2_X1  g0789(.A1(new_n987), .A2(KEYINPUT110), .ZN(new_n990));
  OAI21_X1  g0790(.A(new_n988), .B1(new_n989), .B2(new_n990), .ZN(new_n991));
  XNOR2_X1  g0791(.A(new_n991), .B(KEYINPUT111), .ZN(new_n992));
  INV_X1    g0792(.A(KEYINPUT43), .ZN(new_n993));
  NAND2_X1  g0793(.A1(new_n992), .A2(new_n993), .ZN(new_n994));
  OR2_X1    g0794(.A1(new_n992), .A2(new_n993), .ZN(new_n995));
  NAND3_X1  g0795(.A1(new_n985), .A2(new_n994), .A3(new_n995), .ZN(new_n996));
  NAND4_X1  g0796(.A1(new_n981), .A2(new_n984), .A3(new_n993), .A4(new_n992), .ZN(new_n997));
  NAND2_X1  g0797(.A1(new_n996), .A2(new_n997), .ZN(new_n998));
  INV_X1    g0798(.A(new_n686), .ZN(new_n999));
  NOR2_X1   g0799(.A1(new_n999), .A2(new_n979), .ZN(new_n1000));
  XNOR2_X1  g0800(.A(new_n998), .B(new_n1000), .ZN(new_n1001));
  XOR2_X1   g0801(.A(new_n693), .B(KEYINPUT41), .Z(new_n1002));
  NAND2_X1  g0802(.A1(new_n690), .A2(new_n979), .ZN(new_n1003));
  NAND2_X1  g0803(.A1(new_n1003), .A2(KEYINPUT112), .ZN(new_n1004));
  INV_X1    g0804(.A(KEYINPUT112), .ZN(new_n1005));
  NAND3_X1  g0805(.A1(new_n690), .A2(new_n1005), .A3(new_n979), .ZN(new_n1006));
  NAND2_X1  g0806(.A1(new_n1004), .A2(new_n1006), .ZN(new_n1007));
  INV_X1    g0807(.A(KEYINPUT44), .ZN(new_n1008));
  NAND2_X1  g0808(.A1(new_n1007), .A2(new_n1008), .ZN(new_n1009));
  NOR2_X1   g0809(.A1(new_n690), .A2(new_n979), .ZN(new_n1010));
  XNOR2_X1  g0810(.A(new_n1010), .B(KEYINPUT45), .ZN(new_n1011));
  NAND3_X1  g0811(.A1(new_n1004), .A2(KEYINPUT44), .A3(new_n1006), .ZN(new_n1012));
  NAND3_X1  g0812(.A1(new_n1009), .A2(new_n1011), .A3(new_n1012), .ZN(new_n1013));
  OR2_X1    g0813(.A1(new_n999), .A2(KEYINPUT113), .ZN(new_n1014));
  INV_X1    g0814(.A(new_n1014), .ZN(new_n1015));
  NAND2_X1  g0815(.A1(new_n1013), .A2(new_n1015), .ZN(new_n1016));
  NAND4_X1  g0816(.A1(new_n1014), .A2(new_n1009), .A3(new_n1011), .A4(new_n1012), .ZN(new_n1017));
  INV_X1    g0817(.A(new_n678), .ZN(new_n1018));
  OAI21_X1  g0818(.A(new_n688), .B1(new_n1018), .B2(new_n687), .ZN(new_n1019));
  NAND3_X1  g0819(.A1(new_n1019), .A2(new_n684), .A3(new_n682), .ZN(new_n1020));
  OAI211_X1 g0820(.A(new_n685), .B(new_n688), .C1(new_n1018), .C2(new_n687), .ZN(new_n1021));
  AOI21_X1  g0821(.A(new_n748), .B1(new_n1020), .B2(new_n1021), .ZN(new_n1022));
  NAND3_X1  g0822(.A1(new_n1016), .A2(new_n1017), .A3(new_n1022), .ZN(new_n1023));
  AOI21_X1  g0823(.A(new_n1002), .B1(new_n1023), .B2(new_n749), .ZN(new_n1024));
  OAI21_X1  g0824(.A(new_n1001), .B1(new_n1024), .B2(new_n752), .ZN(new_n1025));
  NAND2_X1  g0825(.A1(new_n992), .A2(new_n811), .ZN(new_n1026));
  INV_X1    g0826(.A(new_n812), .ZN(new_n1027));
  OAI22_X1  g0827(.A1(new_n814), .A2(new_n235), .B1(new_n223), .B2(new_n348), .ZN(new_n1028));
  OAI21_X1  g0828(.A(new_n821), .B1(new_n1027), .B2(new_n1028), .ZN(new_n1029));
  OAI21_X1  g0829(.A(KEYINPUT115), .B1(new_n782), .B2(new_n594), .ZN(new_n1030));
  AOI22_X1  g0830(.A1(new_n767), .A2(G317), .B1(KEYINPUT46), .B2(new_n1030), .ZN(new_n1031));
  OAI21_X1  g0831(.A(new_n1031), .B1(KEYINPUT46), .B2(new_n1030), .ZN(new_n1032));
  AOI22_X1  g0832(.A1(new_n797), .A2(G107), .B1(G294), .B2(new_n777), .ZN(new_n1033));
  XNOR2_X1  g0833(.A(KEYINPUT114), .B(G311), .ZN(new_n1034));
  OAI21_X1  g0834(.A(new_n1033), .B1(new_n775), .B2(new_n1034), .ZN(new_n1035));
  INV_X1    g0835(.A(G283), .ZN(new_n1036));
  OAI221_X1 g0836(.A(new_n384), .B1(new_n1036), .B2(new_n780), .C1(new_n788), .C2(new_n589), .ZN(new_n1037));
  OR3_X1    g0837(.A1(new_n1032), .A2(new_n1035), .A3(new_n1037), .ZN(new_n1038));
  NOR2_X1   g0838(.A1(new_n764), .A2(new_n474), .ZN(new_n1039));
  NOR2_X1   g0839(.A1(new_n764), .A2(new_n280), .ZN(new_n1040));
  NOR2_X1   g0840(.A1(new_n771), .A2(new_n241), .ZN(new_n1041));
  NOR2_X1   g0841(.A1(new_n775), .A2(new_n851), .ZN(new_n1042));
  AOI211_X1 g0842(.A(new_n1041), .B(new_n1042), .C1(G159), .C2(new_n777), .ZN(new_n1043));
  OAI221_X1 g0843(.A(new_n254), .B1(new_n780), .B2(new_n202), .C1(new_n782), .C2(new_n394), .ZN(new_n1044));
  AOI21_X1  g0844(.A(new_n1044), .B1(new_n789), .B2(G150), .ZN(new_n1045));
  INV_X1    g0845(.A(G137), .ZN(new_n1046));
  INV_X1    g0846(.A(new_n767), .ZN(new_n1047));
  OAI211_X1 g0847(.A(new_n1043), .B(new_n1045), .C1(new_n1046), .C2(new_n1047), .ZN(new_n1048));
  OAI22_X1  g0848(.A1(new_n1038), .A2(new_n1039), .B1(new_n1040), .B2(new_n1048), .ZN(new_n1049));
  XNOR2_X1  g0849(.A(new_n1049), .B(KEYINPUT47), .ZN(new_n1050));
  AOI21_X1  g0850(.A(new_n1029), .B1(new_n1050), .B2(new_n756), .ZN(new_n1051));
  NAND2_X1  g0851(.A1(new_n1026), .A2(new_n1051), .ZN(new_n1052));
  XOR2_X1   g0852(.A(new_n1052), .B(KEYINPUT116), .Z(new_n1053));
  NAND2_X1  g0853(.A1(new_n1025), .A2(new_n1053), .ZN(G387));
  NAND2_X1  g0854(.A1(new_n1020), .A2(new_n1021), .ZN(new_n1055));
  NAND2_X1  g0855(.A1(new_n1055), .A2(new_n752), .ZN(new_n1056));
  OR2_X1    g0856(.A1(new_n232), .A2(new_n247), .ZN(new_n1057));
  INV_X1    g0857(.A(new_n695), .ZN(new_n1058));
  AOI22_X1  g0858(.A1(new_n1057), .A2(new_n813), .B1(new_n1058), .B2(new_n817), .ZN(new_n1059));
  NAND2_X1  g0859(.A1(new_n346), .A2(new_n202), .ZN(new_n1060));
  XNOR2_X1  g0860(.A(new_n1060), .B(KEYINPUT50), .ZN(new_n1061));
  OAI21_X1  g0861(.A(new_n443), .B1(new_n241), .B2(new_n280), .ZN(new_n1062));
  NOR3_X1   g0862(.A1(new_n1061), .A2(new_n1058), .A3(new_n1062), .ZN(new_n1063));
  OAI22_X1  g0863(.A1(new_n1059), .A2(new_n1063), .B1(G107), .B2(new_n223), .ZN(new_n1064));
  AOI211_X1 g0864(.A(new_n693), .B(new_n752), .C1(new_n1064), .C2(new_n812), .ZN(new_n1065));
  AOI22_X1  g0865(.A1(new_n789), .A2(G50), .B1(new_n315), .B2(new_n777), .ZN(new_n1066));
  OAI22_X1  g0866(.A1(new_n782), .A2(new_n280), .B1(new_n780), .B2(new_n241), .ZN(new_n1067));
  AOI211_X1 g0867(.A(new_n384), .B(new_n1067), .C1(G159), .C2(new_n774), .ZN(new_n1068));
  XOR2_X1   g0868(.A(KEYINPUT117), .B(G150), .Z(new_n1069));
  NAND2_X1  g0869(.A1(new_n767), .A2(new_n1069), .ZN(new_n1070));
  NAND2_X1  g0870(.A1(new_n565), .A2(new_n797), .ZN(new_n1071));
  NAND4_X1  g0871(.A1(new_n1066), .A2(new_n1068), .A3(new_n1070), .A4(new_n1071), .ZN(new_n1072));
  NOR2_X1   g0872(.A1(new_n1039), .A2(new_n1072), .ZN(new_n1073));
  OAI21_X1  g0873(.A(new_n384), .B1(new_n1047), .B2(new_n795), .ZN(new_n1074));
  AOI22_X1  g0874(.A1(new_n848), .A2(G303), .B1(G322), .B2(new_n774), .ZN(new_n1075));
  INV_X1    g0875(.A(G317), .ZN(new_n1076));
  OAI221_X1 g0876(.A(new_n1075), .B1(new_n793), .B2(new_n1034), .C1(new_n788), .C2(new_n1076), .ZN(new_n1077));
  INV_X1    g0877(.A(KEYINPUT48), .ZN(new_n1078));
  OR2_X1    g0878(.A1(new_n1077), .A2(new_n1078), .ZN(new_n1079));
  NAND2_X1  g0879(.A1(new_n1077), .A2(new_n1078), .ZN(new_n1080));
  INV_X1    g0880(.A(new_n782), .ZN(new_n1081));
  AOI22_X1  g0881(.A1(new_n1081), .A2(G294), .B1(new_n797), .B2(G283), .ZN(new_n1082));
  NAND3_X1  g0882(.A1(new_n1079), .A2(new_n1080), .A3(new_n1082), .ZN(new_n1083));
  INV_X1    g0883(.A(KEYINPUT49), .ZN(new_n1084));
  NOR2_X1   g0884(.A1(new_n1083), .A2(new_n1084), .ZN(new_n1085));
  AOI211_X1 g0885(.A(new_n1074), .B(new_n1085), .C1(G116), .C2(new_n765), .ZN(new_n1086));
  NAND2_X1  g0886(.A1(new_n1083), .A2(new_n1084), .ZN(new_n1087));
  AOI21_X1  g0887(.A(new_n1073), .B1(new_n1086), .B2(new_n1087), .ZN(new_n1088));
  OAI221_X1 g0888(.A(new_n1065), .B1(new_n757), .B2(new_n1088), .C1(new_n1018), .C2(new_n810), .ZN(new_n1089));
  OR2_X1    g0889(.A1(new_n1022), .A2(new_n694), .ZN(new_n1090));
  NOR2_X1   g0890(.A1(new_n1055), .A2(new_n749), .ZN(new_n1091));
  OAI211_X1 g0891(.A(new_n1056), .B(new_n1089), .C1(new_n1090), .C2(new_n1091), .ZN(G393));
  OR2_X1    g0892(.A1(new_n1013), .A2(new_n686), .ZN(new_n1093));
  NAND2_X1  g0893(.A1(new_n1013), .A2(new_n686), .ZN(new_n1094));
  NAND3_X1  g0894(.A1(new_n1093), .A2(new_n752), .A3(new_n1094), .ZN(new_n1095));
  NAND2_X1  g0895(.A1(new_n979), .A2(new_n811), .ZN(new_n1096));
  XNOR2_X1  g0896(.A(new_n1096), .B(KEYINPUT118), .ZN(new_n1097));
  AOI22_X1  g0897(.A1(new_n789), .A2(G159), .B1(G150), .B2(new_n774), .ZN(new_n1098));
  XOR2_X1   g0898(.A(new_n1098), .B(KEYINPUT51), .Z(new_n1099));
  NOR2_X1   g0899(.A1(new_n771), .A2(new_n280), .ZN(new_n1100));
  AOI21_X1  g0900(.A(new_n1100), .B1(new_n777), .B2(G50), .ZN(new_n1101));
  AOI22_X1  g0901(.A1(new_n1081), .A2(G68), .B1(new_n848), .B2(new_n346), .ZN(new_n1102));
  NAND3_X1  g0902(.A1(new_n1101), .A2(new_n1102), .A3(new_n503), .ZN(new_n1103));
  AOI21_X1  g0903(.A(new_n1103), .B1(G143), .B2(new_n767), .ZN(new_n1104));
  NAND3_X1  g0904(.A1(new_n1099), .A2(new_n840), .A3(new_n1104), .ZN(new_n1105));
  OAI22_X1  g0905(.A1(new_n788), .A2(new_n800), .B1(new_n1076), .B2(new_n775), .ZN(new_n1106));
  XNOR2_X1  g0906(.A(new_n1106), .B(KEYINPUT52), .ZN(new_n1107));
  OAI22_X1  g0907(.A1(new_n793), .A2(new_n589), .B1(new_n771), .B2(new_n594), .ZN(new_n1108));
  OAI221_X1 g0908(.A(new_n410), .B1(new_n780), .B2(new_n511), .C1(new_n782), .C2(new_n1036), .ZN(new_n1109));
  AOI211_X1 g0909(.A(new_n1108), .B(new_n1109), .C1(G322), .C2(new_n767), .ZN(new_n1110));
  NAND3_X1  g0910(.A1(new_n766), .A2(new_n1107), .A3(new_n1110), .ZN(new_n1111));
  AOI21_X1  g0911(.A(new_n757), .B1(new_n1105), .B2(new_n1111), .ZN(new_n1112));
  OAI22_X1  g0912(.A1(new_n814), .A2(new_n239), .B1(new_n474), .B2(new_n223), .ZN(new_n1113));
  OAI21_X1  g0913(.A(new_n821), .B1(new_n1027), .B2(new_n1113), .ZN(new_n1114));
  OR3_X1    g0914(.A1(new_n1097), .A2(new_n1112), .A3(new_n1114), .ZN(new_n1115));
  NAND2_X1  g0915(.A1(new_n1023), .A2(new_n693), .ZN(new_n1116));
  AOI21_X1  g0916(.A(new_n1022), .B1(new_n1093), .B2(new_n1094), .ZN(new_n1117));
  OAI211_X1 g0917(.A(new_n1095), .B(new_n1115), .C1(new_n1116), .C2(new_n1117), .ZN(G390));
  INV_X1    g0918(.A(G330), .ZN(new_n1119));
  AOI21_X1  g0919(.A(new_n1119), .B1(new_n879), .B2(new_n883), .ZN(new_n1120));
  NAND2_X1  g0920(.A1(new_n1120), .A2(new_n435), .ZN(new_n1121));
  NAND3_X1  g0921(.A1(new_n1121), .A2(new_n970), .A3(new_n633), .ZN(new_n1122));
  NAND3_X1  g0922(.A1(new_n947), .A2(G330), .A3(new_n830), .ZN(new_n1123));
  NAND2_X1  g0923(.A1(new_n1123), .A2(new_n963), .ZN(new_n1124));
  NAND2_X1  g0924(.A1(new_n829), .A2(new_n366), .ZN(new_n1125));
  NAND3_X1  g0925(.A1(new_n713), .A2(new_n675), .A3(new_n1125), .ZN(new_n1126));
  INV_X1    g0926(.A(new_n826), .ZN(new_n1127));
  NAND2_X1  g0927(.A1(new_n1126), .A2(new_n1127), .ZN(new_n1128));
  NAND2_X1  g0928(.A1(new_n1128), .A2(KEYINPUT119), .ZN(new_n1129));
  INV_X1    g0929(.A(KEYINPUT119), .ZN(new_n1130));
  NAND3_X1  g0930(.A1(new_n1126), .A2(new_n1130), .A3(new_n1127), .ZN(new_n1131));
  NAND2_X1  g0931(.A1(new_n1129), .A2(new_n1131), .ZN(new_n1132));
  NAND4_X1  g0932(.A1(new_n746), .A2(new_n684), .A3(new_n830), .A4(new_n876), .ZN(new_n1133));
  NAND3_X1  g0933(.A1(new_n1124), .A2(new_n1132), .A3(new_n1133), .ZN(new_n1134));
  AOI21_X1  g0934(.A(new_n965), .B1(new_n701), .B2(new_n830), .ZN(new_n1135));
  INV_X1    g0935(.A(new_n1135), .ZN(new_n1136));
  AND2_X1   g0936(.A1(new_n746), .A2(new_n684), .ZN(new_n1137));
  AOI21_X1  g0937(.A(new_n876), .B1(new_n1137), .B2(new_n830), .ZN(new_n1138));
  AOI211_X1 g0938(.A(new_n1119), .B(new_n877), .C1(new_n883), .C2(new_n879), .ZN(new_n1139));
  OAI21_X1  g0939(.A(new_n1136), .B1(new_n1138), .B2(new_n1139), .ZN(new_n1140));
  AOI21_X1  g0940(.A(new_n1122), .B1(new_n1134), .B2(new_n1140), .ZN(new_n1141));
  AOI22_X1  g0941(.A1(new_n943), .A2(new_n954), .B1(new_n958), .B2(KEYINPUT39), .ZN(new_n1142));
  OAI21_X1  g0942(.A(new_n1142), .B1(new_n967), .B2(new_n961), .ZN(new_n1143));
  AND3_X1   g0943(.A1(new_n1126), .A2(new_n1130), .A3(new_n1127), .ZN(new_n1144));
  AOI21_X1  g0944(.A(new_n1130), .B1(new_n1126), .B2(new_n1127), .ZN(new_n1145));
  NOR3_X1   g0945(.A1(new_n1144), .A2(new_n1145), .A3(new_n963), .ZN(new_n1146));
  AOI21_X1  g0946(.A(new_n961), .B1(new_n943), .B2(new_n928), .ZN(new_n1147));
  INV_X1    g0947(.A(new_n1147), .ZN(new_n1148));
  OAI211_X1 g0948(.A(new_n1143), .B(new_n1133), .C1(new_n1146), .C2(new_n1148), .ZN(new_n1149));
  NAND3_X1  g0949(.A1(new_n1129), .A2(new_n876), .A3(new_n1131), .ZN(new_n1150));
  INV_X1    g0950(.A(new_n961), .ZN(new_n1151));
  OAI21_X1  g0951(.A(new_n1151), .B1(new_n1135), .B2(new_n963), .ZN(new_n1152));
  AOI22_X1  g0952(.A1(new_n1150), .A2(new_n1147), .B1(new_n1152), .B2(new_n1142), .ZN(new_n1153));
  NAND4_X1  g0953(.A1(new_n947), .A2(G330), .A3(new_n830), .A4(new_n876), .ZN(new_n1154));
  OAI211_X1 g0954(.A(new_n1141), .B(new_n1149), .C1(new_n1153), .C2(new_n1154), .ZN(new_n1155));
  OAI21_X1  g0955(.A(new_n1149), .B1(new_n1153), .B2(new_n1154), .ZN(new_n1156));
  AND3_X1   g0956(.A1(new_n1121), .A2(new_n970), .A3(new_n633), .ZN(new_n1157));
  AOI21_X1  g0957(.A(new_n876), .B1(new_n1120), .B2(new_n830), .ZN(new_n1158));
  OAI21_X1  g0958(.A(new_n1133), .B1(new_n1144), .B2(new_n1145), .ZN(new_n1159));
  NOR2_X1   g0959(.A1(new_n1158), .A2(new_n1159), .ZN(new_n1160));
  OAI21_X1  g0960(.A(new_n963), .B1(new_n747), .B2(new_n831), .ZN(new_n1161));
  AOI21_X1  g0961(.A(new_n1135), .B1(new_n1154), .B2(new_n1161), .ZN(new_n1162));
  OAI21_X1  g0962(.A(new_n1157), .B1(new_n1160), .B2(new_n1162), .ZN(new_n1163));
  AOI21_X1  g0963(.A(new_n694), .B1(new_n1156), .B2(new_n1163), .ZN(new_n1164));
  NAND2_X1  g0964(.A1(new_n1155), .A2(new_n1164), .ZN(new_n1165));
  OAI211_X1 g0965(.A(new_n1149), .B(new_n752), .C1(new_n1153), .C2(new_n1154), .ZN(new_n1166));
  OAI21_X1  g0966(.A(new_n821), .B1(new_n315), .B2(new_n838), .ZN(new_n1167));
  OAI22_X1  g0967(.A1(new_n793), .A2(new_n354), .B1(new_n775), .B2(new_n1036), .ZN(new_n1168));
  AOI211_X1 g0968(.A(new_n1100), .B(new_n1168), .C1(G97), .C2(new_n848), .ZN(new_n1169));
  AOI21_X1  g0969(.A(new_n254), .B1(new_n1081), .B2(G87), .ZN(new_n1170));
  AOI22_X1  g0970(.A1(new_n767), .A2(G294), .B1(new_n1170), .B2(KEYINPUT120), .ZN(new_n1171));
  NOR2_X1   g0971(.A1(new_n1170), .A2(KEYINPUT120), .ZN(new_n1172));
  AOI21_X1  g0972(.A(new_n1172), .B1(G116), .B2(new_n789), .ZN(new_n1173));
  NAND4_X1  g0973(.A1(new_n847), .A2(new_n1169), .A3(new_n1171), .A4(new_n1173), .ZN(new_n1174));
  NOR2_X1   g0974(.A1(new_n764), .A2(new_n202), .ZN(new_n1175));
  NAND2_X1  g0975(.A1(new_n1081), .A2(new_n1069), .ZN(new_n1176));
  XNOR2_X1  g0976(.A(new_n1176), .B(KEYINPUT53), .ZN(new_n1177));
  AOI21_X1  g0977(.A(new_n1177), .B1(G125), .B2(new_n767), .ZN(new_n1178));
  XNOR2_X1  g0978(.A(KEYINPUT54), .B(G143), .ZN(new_n1179));
  OAI21_X1  g0979(.A(new_n254), .B1(new_n780), .B2(new_n1179), .ZN(new_n1180));
  INV_X1    g0980(.A(G128), .ZN(new_n1181));
  OAI22_X1  g0981(.A1(new_n793), .A2(new_n1046), .B1(new_n775), .B2(new_n1181), .ZN(new_n1182));
  AOI211_X1 g0982(.A(new_n1180), .B(new_n1182), .C1(G159), .C2(new_n797), .ZN(new_n1183));
  NAND2_X1  g0983(.A1(new_n789), .A2(G132), .ZN(new_n1184));
  NAND3_X1  g0984(.A1(new_n1178), .A2(new_n1183), .A3(new_n1184), .ZN(new_n1185));
  OAI21_X1  g0985(.A(new_n1174), .B1(new_n1175), .B2(new_n1185), .ZN(new_n1186));
  AOI21_X1  g0986(.A(new_n1167), .B1(new_n1186), .B2(new_n756), .ZN(new_n1187));
  OAI21_X1  g0987(.A(new_n1187), .B1(new_n960), .B2(new_n837), .ZN(new_n1188));
  NAND2_X1  g0988(.A1(new_n1166), .A2(new_n1188), .ZN(new_n1189));
  INV_X1    g0989(.A(new_n1189), .ZN(new_n1190));
  NAND2_X1  g0990(.A1(new_n1165), .A2(new_n1190), .ZN(G378));
  OAI21_X1  g0991(.A(new_n1157), .B1(new_n1156), .B2(new_n1163), .ZN(new_n1192));
  INV_X1    g0992(.A(KEYINPUT57), .ZN(new_n1193));
  NAND2_X1  g0993(.A1(new_n931), .A2(new_n932), .ZN(new_n1194));
  NAND2_X1  g0994(.A1(new_n884), .A2(new_n944), .ZN(new_n1195));
  NAND3_X1  g0995(.A1(new_n1194), .A2(G330), .A3(new_n1195), .ZN(new_n1196));
  NAND2_X1  g0996(.A1(new_n342), .A2(new_n336), .ZN(new_n1197));
  OAI21_X1  g0997(.A(new_n904), .B1(new_n320), .B2(new_n307), .ZN(new_n1198));
  XNOR2_X1  g0998(.A(new_n1197), .B(new_n1198), .ZN(new_n1199));
  XNOR2_X1  g0999(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1200));
  XNOR2_X1  g1000(.A(new_n1199), .B(new_n1200), .ZN(new_n1201));
  AOI21_X1  g1001(.A(new_n1201), .B1(new_n962), .B2(new_n968), .ZN(new_n1202));
  INV_X1    g1002(.A(KEYINPUT39), .ZN(new_n1203));
  NAND2_X1  g1003(.A1(new_n928), .A2(new_n1203), .ZN(new_n1204));
  AOI21_X1  g1004(.A(new_n1204), .B1(new_n938), .B2(new_n942), .ZN(new_n1205));
  AOI21_X1  g1005(.A(new_n1203), .B1(new_n927), .B2(new_n928), .ZN(new_n1206));
  OAI21_X1  g1006(.A(new_n961), .B1(new_n1205), .B2(new_n1206), .ZN(new_n1207));
  INV_X1    g1007(.A(new_n952), .ZN(new_n1208));
  AND4_X1   g1008(.A1(new_n968), .A2(new_n1207), .A3(new_n1208), .A4(new_n1201), .ZN(new_n1209));
  OAI21_X1  g1009(.A(new_n1196), .B1(new_n1202), .B2(new_n1209), .ZN(new_n1210));
  INV_X1    g1010(.A(new_n1201), .ZN(new_n1211));
  OAI21_X1  g1011(.A(new_n1208), .B1(new_n1142), .B2(new_n1151), .ZN(new_n1212));
  AND2_X1   g1012(.A1(new_n967), .A2(new_n930), .ZN(new_n1213));
  OAI21_X1  g1013(.A(new_n1211), .B1(new_n1212), .B2(new_n1213), .ZN(new_n1214));
  NAND4_X1  g1014(.A1(new_n1207), .A2(new_n968), .A3(new_n1201), .A4(new_n1208), .ZN(new_n1215));
  NAND4_X1  g1015(.A1(new_n1214), .A2(G330), .A3(new_n945), .A4(new_n1215), .ZN(new_n1216));
  AOI21_X1  g1016(.A(new_n1193), .B1(new_n1210), .B2(new_n1216), .ZN(new_n1217));
  NAND2_X1  g1017(.A1(new_n1192), .A2(new_n1217), .ZN(new_n1218));
  NAND2_X1  g1018(.A1(new_n1218), .A2(new_n693), .ZN(new_n1219));
  NAND2_X1  g1019(.A1(new_n1210), .A2(new_n1216), .ZN(new_n1220));
  AOI21_X1  g1020(.A(KEYINPUT57), .B1(new_n1192), .B2(new_n1220), .ZN(new_n1221));
  OR2_X1    g1021(.A1(new_n1219), .A2(new_n1221), .ZN(new_n1222));
  OAI21_X1  g1022(.A(new_n821), .B1(G50), .B2(new_n838), .ZN(new_n1223));
  NAND2_X1  g1023(.A1(new_n765), .A2(new_n314), .ZN(new_n1224));
  OAI22_X1  g1024(.A1(new_n793), .A2(new_n474), .B1(new_n775), .B2(new_n594), .ZN(new_n1225));
  AOI211_X1 g1025(.A(new_n1041), .B(new_n1225), .C1(G77), .C2(new_n1081), .ZN(new_n1226));
  NAND2_X1  g1026(.A1(new_n384), .A2(new_n248), .ZN(new_n1227));
  AOI21_X1  g1027(.A(new_n1227), .B1(new_n565), .B2(new_n848), .ZN(new_n1228));
  AOI22_X1  g1028(.A1(new_n789), .A2(G107), .B1(new_n767), .B2(G283), .ZN(new_n1229));
  NAND4_X1  g1029(.A1(new_n1224), .A2(new_n1226), .A3(new_n1228), .A4(new_n1229), .ZN(new_n1230));
  INV_X1    g1030(.A(KEYINPUT58), .ZN(new_n1231));
  AOI21_X1  g1031(.A(G50), .B1(new_n316), .B2(new_n248), .ZN(new_n1232));
  AOI22_X1  g1032(.A1(new_n1230), .A2(new_n1231), .B1(new_n1227), .B2(new_n1232), .ZN(new_n1233));
  OAI22_X1  g1033(.A1(new_n782), .A2(new_n1179), .B1(new_n780), .B2(new_n1046), .ZN(new_n1234));
  AOI21_X1  g1034(.A(new_n1234), .B1(G132), .B2(new_n777), .ZN(new_n1235));
  AOI22_X1  g1035(.A1(new_n797), .A2(G150), .B1(G125), .B2(new_n774), .ZN(new_n1236));
  OAI211_X1 g1036(.A(new_n1235), .B(new_n1236), .C1(new_n1181), .C2(new_n788), .ZN(new_n1237));
  XOR2_X1   g1037(.A(new_n1237), .B(KEYINPUT59), .Z(new_n1238));
  INV_X1    g1038(.A(new_n1238), .ZN(new_n1239));
  NOR2_X1   g1039(.A1(new_n1239), .A2(KEYINPUT121), .ZN(new_n1240));
  NAND2_X1  g1040(.A1(new_n765), .A2(G159), .ZN(new_n1241));
  AOI211_X1 g1041(.A(G33), .B(G41), .C1(new_n767), .C2(G124), .ZN(new_n1242));
  INV_X1    g1042(.A(KEYINPUT121), .ZN(new_n1243));
  OAI211_X1 g1043(.A(new_n1241), .B(new_n1242), .C1(new_n1238), .C2(new_n1243), .ZN(new_n1244));
  OAI221_X1 g1044(.A(new_n1233), .B1(new_n1231), .B2(new_n1230), .C1(new_n1240), .C2(new_n1244), .ZN(new_n1245));
  AOI21_X1  g1045(.A(new_n1223), .B1(new_n1245), .B2(new_n756), .ZN(new_n1246));
  OAI21_X1  g1046(.A(new_n1246), .B1(new_n1201), .B2(new_n837), .ZN(new_n1247));
  XNOR2_X1  g1047(.A(new_n1247), .B(KEYINPUT122), .ZN(new_n1248));
  AOI21_X1  g1048(.A(new_n1248), .B1(new_n1220), .B2(new_n752), .ZN(new_n1249));
  NAND2_X1  g1049(.A1(new_n1222), .A2(new_n1249), .ZN(G375));
  NAND2_X1  g1050(.A1(new_n963), .A2(new_n808), .ZN(new_n1251));
  OAI21_X1  g1051(.A(new_n821), .B1(G68), .B2(new_n838), .ZN(new_n1252));
  NAND2_X1  g1052(.A1(new_n774), .A2(G132), .ZN(new_n1253));
  OAI21_X1  g1053(.A(new_n1253), .B1(new_n793), .B2(new_n1179), .ZN(new_n1254));
  AOI21_X1  g1054(.A(new_n1254), .B1(G50), .B2(new_n797), .ZN(new_n1255));
  NAND2_X1  g1055(.A1(new_n789), .A2(G137), .ZN(new_n1256));
  AOI21_X1  g1056(.A(new_n384), .B1(G150), .B2(new_n848), .ZN(new_n1257));
  NAND4_X1  g1057(.A1(new_n1224), .A2(new_n1255), .A3(new_n1256), .A4(new_n1257), .ZN(new_n1258));
  AOI22_X1  g1058(.A1(new_n767), .A2(G128), .B1(G159), .B2(new_n1081), .ZN(new_n1259));
  XNOR2_X1  g1059(.A(new_n1259), .B(KEYINPUT123), .ZN(new_n1260));
  OAI21_X1  g1060(.A(new_n410), .B1(new_n780), .B2(new_n354), .ZN(new_n1261));
  OAI22_X1  g1061(.A1(new_n793), .A2(new_n594), .B1(new_n775), .B2(new_n511), .ZN(new_n1262));
  AOI211_X1 g1062(.A(new_n1261), .B(new_n1262), .C1(G97), .C2(new_n1081), .ZN(new_n1263));
  NAND2_X1  g1063(.A1(new_n767), .A2(G303), .ZN(new_n1264));
  NAND2_X1  g1064(.A1(new_n789), .A2(G283), .ZN(new_n1265));
  NAND4_X1  g1065(.A1(new_n1263), .A2(new_n1071), .A3(new_n1264), .A4(new_n1265), .ZN(new_n1266));
  OAI22_X1  g1066(.A1(new_n1258), .A2(new_n1260), .B1(new_n1266), .B2(new_n1040), .ZN(new_n1267));
  AOI21_X1  g1067(.A(new_n1252), .B1(new_n1267), .B2(new_n756), .ZN(new_n1268));
  NAND2_X1  g1068(.A1(new_n1251), .A2(new_n1268), .ZN(new_n1269));
  NOR2_X1   g1069(.A1(new_n1160), .A2(new_n1162), .ZN(new_n1270));
  OAI21_X1  g1070(.A(new_n1269), .B1(new_n1270), .B2(new_n751), .ZN(new_n1271));
  INV_X1    g1071(.A(new_n1271), .ZN(new_n1272));
  NAND3_X1  g1072(.A1(new_n1134), .A2(new_n1140), .A3(new_n1122), .ZN(new_n1273));
  INV_X1    g1073(.A(new_n1002), .ZN(new_n1274));
  NAND3_X1  g1074(.A1(new_n1273), .A2(new_n1163), .A3(new_n1274), .ZN(new_n1275));
  NAND2_X1  g1075(.A1(new_n1272), .A2(new_n1275), .ZN(G381));
  INV_X1    g1076(.A(G390), .ZN(new_n1277));
  NOR4_X1   g1077(.A1(G393), .A2(G381), .A3(G396), .A4(G384), .ZN(new_n1278));
  AOI21_X1  g1078(.A(new_n1189), .B1(new_n1155), .B2(new_n1164), .ZN(new_n1279));
  NAND3_X1  g1079(.A1(new_n1277), .A2(new_n1278), .A3(new_n1279), .ZN(new_n1280));
  OR3_X1    g1080(.A1(new_n1280), .A2(G387), .A3(G375), .ZN(G407));
  NAND2_X1  g1081(.A1(new_n667), .A2(G213), .ZN(new_n1282));
  INV_X1    g1082(.A(new_n1282), .ZN(new_n1283));
  NAND2_X1  g1083(.A1(new_n1279), .A2(new_n1283), .ZN(new_n1284));
  OAI211_X1 g1084(.A(G407), .B(G213), .C1(G375), .C2(new_n1284), .ZN(G409));
  OAI211_X1 g1085(.A(G378), .B(new_n1249), .C1(new_n1219), .C2(new_n1221), .ZN(new_n1286));
  NAND3_X1  g1086(.A1(new_n1192), .A2(new_n1274), .A3(new_n1220), .ZN(new_n1287));
  NAND2_X1  g1087(.A1(new_n1287), .A2(new_n1247), .ZN(new_n1288));
  AND3_X1   g1088(.A1(new_n1210), .A2(new_n1216), .A3(KEYINPUT124), .ZN(new_n1289));
  AOI21_X1  g1089(.A(KEYINPUT124), .B1(new_n1210), .B2(new_n1216), .ZN(new_n1290));
  NOR3_X1   g1090(.A1(new_n1289), .A2(new_n1290), .A3(new_n751), .ZN(new_n1291));
  OAI21_X1  g1091(.A(new_n1279), .B1(new_n1288), .B2(new_n1291), .ZN(new_n1292));
  NAND2_X1  g1092(.A1(new_n1286), .A2(new_n1292), .ZN(new_n1293));
  NAND4_X1  g1093(.A1(new_n1134), .A2(new_n1140), .A3(KEYINPUT60), .A4(new_n1122), .ZN(new_n1294));
  AND2_X1   g1094(.A1(new_n1294), .A2(new_n693), .ZN(new_n1295));
  INV_X1    g1095(.A(KEYINPUT60), .ZN(new_n1296));
  OAI21_X1  g1096(.A(new_n1273), .B1(new_n1141), .B2(new_n1296), .ZN(new_n1297));
  NAND2_X1  g1097(.A1(new_n1295), .A2(new_n1297), .ZN(new_n1298));
  AOI21_X1  g1098(.A(G384), .B1(new_n1298), .B2(new_n1272), .ZN(new_n1299));
  AOI211_X1 g1099(.A(new_n864), .B(new_n1271), .C1(new_n1295), .C2(new_n1297), .ZN(new_n1300));
  NOR2_X1   g1100(.A1(new_n1299), .A2(new_n1300), .ZN(new_n1301));
  NAND3_X1  g1101(.A1(new_n1293), .A2(new_n1282), .A3(new_n1301), .ZN(new_n1302));
  INV_X1    g1102(.A(KEYINPUT125), .ZN(new_n1303));
  NAND2_X1  g1103(.A1(new_n1302), .A2(new_n1303), .ZN(new_n1304));
  AOI21_X1  g1104(.A(new_n1283), .B1(new_n1286), .B2(new_n1292), .ZN(new_n1305));
  NAND3_X1  g1105(.A1(new_n1305), .A2(KEYINPUT125), .A3(new_n1301), .ZN(new_n1306));
  AOI21_X1  g1106(.A(KEYINPUT62), .B1(new_n1304), .B2(new_n1306), .ZN(new_n1307));
  NAND2_X1  g1107(.A1(new_n1293), .A2(new_n1282), .ZN(new_n1308));
  NAND2_X1  g1108(.A1(new_n1283), .A2(G2897), .ZN(new_n1309));
  INV_X1    g1109(.A(new_n1309), .ZN(new_n1310));
  NOR3_X1   g1110(.A1(new_n1299), .A2(new_n1300), .A3(new_n1310), .ZN(new_n1311));
  NAND2_X1  g1111(.A1(new_n1294), .A2(new_n693), .ZN(new_n1312));
  NAND2_X1  g1112(.A1(new_n1163), .A2(KEYINPUT60), .ZN(new_n1313));
  AOI21_X1  g1113(.A(new_n1312), .B1(new_n1273), .B2(new_n1313), .ZN(new_n1314));
  OAI21_X1  g1114(.A(new_n864), .B1(new_n1314), .B2(new_n1271), .ZN(new_n1315));
  NAND3_X1  g1115(.A1(new_n1298), .A2(G384), .A3(new_n1272), .ZN(new_n1316));
  AOI21_X1  g1116(.A(new_n1309), .B1(new_n1315), .B2(new_n1316), .ZN(new_n1317));
  NOR2_X1   g1117(.A1(new_n1311), .A2(new_n1317), .ZN(new_n1318));
  AOI21_X1  g1118(.A(KEYINPUT61), .B1(new_n1308), .B2(new_n1318), .ZN(new_n1319));
  NAND2_X1  g1119(.A1(new_n1302), .A2(KEYINPUT62), .ZN(new_n1320));
  NAND2_X1  g1120(.A1(new_n1319), .A2(new_n1320), .ZN(new_n1321));
  OAI21_X1  g1121(.A(KEYINPUT126), .B1(new_n1307), .B2(new_n1321), .ZN(new_n1322));
  XNOR2_X1  g1122(.A(G393), .B(new_n824), .ZN(new_n1323));
  INV_X1    g1123(.A(new_n1323), .ZN(new_n1324));
  NAND3_X1  g1124(.A1(new_n1025), .A2(G390), .A3(new_n1053), .ZN(new_n1325));
  INV_X1    g1125(.A(new_n1325), .ZN(new_n1326));
  AOI21_X1  g1126(.A(G390), .B1(new_n1025), .B2(new_n1053), .ZN(new_n1327));
  OAI21_X1  g1127(.A(new_n1324), .B1(new_n1326), .B2(new_n1327), .ZN(new_n1328));
  NAND2_X1  g1128(.A1(G387), .A2(new_n1277), .ZN(new_n1329));
  NAND3_X1  g1129(.A1(new_n1329), .A2(new_n1323), .A3(new_n1325), .ZN(new_n1330));
  NAND2_X1  g1130(.A1(new_n1328), .A2(new_n1330), .ZN(new_n1331));
  INV_X1    g1131(.A(KEYINPUT62), .ZN(new_n1332));
  AND4_X1   g1132(.A1(KEYINPUT125), .A2(new_n1293), .A3(new_n1282), .A4(new_n1301), .ZN(new_n1333));
  AOI21_X1  g1133(.A(KEYINPUT125), .B1(new_n1305), .B2(new_n1301), .ZN(new_n1334));
  OAI21_X1  g1134(.A(new_n1332), .B1(new_n1333), .B2(new_n1334), .ZN(new_n1335));
  INV_X1    g1135(.A(KEYINPUT126), .ZN(new_n1336));
  INV_X1    g1136(.A(KEYINPUT61), .ZN(new_n1337));
  OAI21_X1  g1137(.A(new_n1310), .B1(new_n1299), .B2(new_n1300), .ZN(new_n1338));
  NAND3_X1  g1138(.A1(new_n1315), .A2(new_n1316), .A3(new_n1309), .ZN(new_n1339));
  NAND2_X1  g1139(.A1(new_n1338), .A2(new_n1339), .ZN(new_n1340));
  OAI21_X1  g1140(.A(new_n1337), .B1(new_n1305), .B2(new_n1340), .ZN(new_n1341));
  AOI21_X1  g1141(.A(new_n1332), .B1(new_n1305), .B2(new_n1301), .ZN(new_n1342));
  NOR2_X1   g1142(.A1(new_n1341), .A2(new_n1342), .ZN(new_n1343));
  NAND3_X1  g1143(.A1(new_n1335), .A2(new_n1336), .A3(new_n1343), .ZN(new_n1344));
  NAND3_X1  g1144(.A1(new_n1322), .A2(new_n1331), .A3(new_n1344), .ZN(new_n1345));
  INV_X1    g1145(.A(new_n1302), .ZN(new_n1346));
  AOI21_X1  g1146(.A(new_n1331), .B1(KEYINPUT63), .B2(new_n1346), .ZN(new_n1347));
  OR3_X1    g1147(.A1(new_n1333), .A2(new_n1334), .A3(KEYINPUT63), .ZN(new_n1348));
  NAND3_X1  g1148(.A1(new_n1347), .A2(new_n1348), .A3(new_n1319), .ZN(new_n1349));
  NAND2_X1  g1149(.A1(new_n1345), .A2(new_n1349), .ZN(G405));
  AOI21_X1  g1150(.A(G378), .B1(new_n1222), .B2(new_n1249), .ZN(new_n1351));
  INV_X1    g1151(.A(new_n1286), .ZN(new_n1352));
  NOR2_X1   g1152(.A1(new_n1351), .A2(new_n1352), .ZN(new_n1353));
  NOR3_X1   g1153(.A1(new_n1299), .A2(new_n1300), .A3(KEYINPUT127), .ZN(new_n1354));
  XNOR2_X1  g1154(.A(new_n1353), .B(new_n1354), .ZN(new_n1355));
  XOR2_X1   g1155(.A(new_n1355), .B(new_n1331), .Z(G402));
endmodule


