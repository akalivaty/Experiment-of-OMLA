//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 0 0 1 1 0 0 1 1 0 1 0 1 1 1 0 0 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 0 0 0 1 1 0 0 0 0 0 0 0 1 1 1 1 1 0 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:42:11 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n236, new_n237,
    new_n238, new_n239, new_n240, new_n241, new_n242, new_n244, new_n245,
    new_n246, new_n247, new_n248, new_n249, new_n250, new_n252, new_n253,
    new_n254, new_n255, new_n256, new_n257, new_n258, new_n259, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n609, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n699,
    new_n700, new_n701, new_n702, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n812, new_n813,
    new_n814, new_n815, new_n816, new_n817, new_n818, new_n819, new_n820,
    new_n821, new_n822, new_n823, new_n824, new_n825, new_n826, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n898,
    new_n899, new_n900, new_n901, new_n902, new_n903, new_n904, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n980, new_n981, new_n982, new_n983,
    new_n984, new_n985, new_n986, new_n987, new_n988, new_n989, new_n990,
    new_n991, new_n992, new_n993, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1019, new_n1020, new_n1021, new_n1022,
    new_n1023, new_n1024, new_n1025, new_n1026, new_n1027, new_n1028,
    new_n1029, new_n1030, new_n1031, new_n1032, new_n1033, new_n1034,
    new_n1035, new_n1036, new_n1037, new_n1038, new_n1039, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1045, new_n1047,
    new_n1048, new_n1049, new_n1050, new_n1051, new_n1052, new_n1053,
    new_n1054, new_n1055, new_n1056, new_n1057, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1106, new_n1107, new_n1108,
    new_n1109, new_n1110, new_n1111, new_n1112, new_n1113, new_n1114,
    new_n1115, new_n1116, new_n1117, new_n1118, new_n1119, new_n1120,
    new_n1121, new_n1122, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1177, new_n1178, new_n1179, new_n1180, new_n1181,
    new_n1182, new_n1183, new_n1184, new_n1185, new_n1186, new_n1187,
    new_n1188, new_n1189, new_n1190, new_n1191, new_n1192, new_n1193,
    new_n1194, new_n1195, new_n1196, new_n1197, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1212, new_n1213,
    new_n1215, new_n1216, new_n1217, new_n1218, new_n1219, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1273, new_n1274, new_n1275,
    new_n1276, new_n1277, new_n1278, new_n1279, new_n1280, new_n1281;
  INV_X1    g0000(.A(G58), .ZN(new_n201));
  INV_X1    g0001(.A(G68), .ZN(new_n202));
  NAND3_X1  g0002(.A1(new_n201), .A2(new_n202), .A3(KEYINPUT64), .ZN(new_n203));
  INV_X1    g0003(.A(KEYINPUT64), .ZN(new_n204));
  OAI21_X1  g0004(.A(new_n204), .B1(G58), .B2(G68), .ZN(new_n205));
  NAND2_X1  g0005(.A1(new_n203), .A2(new_n205), .ZN(new_n206));
  INV_X1    g0006(.A(G50), .ZN(new_n207));
  NAND2_X1  g0007(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  INV_X1    g0008(.A(KEYINPUT65), .ZN(new_n209));
  XNOR2_X1  g0009(.A(new_n208), .B(new_n209), .ZN(new_n210));
  INV_X1    g0010(.A(G77), .ZN(new_n211));
  NAND2_X1  g0011(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  XOR2_X1   g0012(.A(new_n212), .B(KEYINPUT66), .Z(G353));
  OAI21_X1  g0013(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND3_X1  g0014(.A1(new_n203), .A2(new_n205), .A3(G50), .ZN(new_n215));
  XOR2_X1   g0015(.A(new_n215), .B(KEYINPUT68), .Z(new_n216));
  XOR2_X1   g0016(.A(new_n216), .B(KEYINPUT69), .Z(new_n217));
  INV_X1    g0017(.A(new_n217), .ZN(new_n218));
  NAND2_X1  g0018(.A1(G1), .A2(G13), .ZN(new_n219));
  INV_X1    g0019(.A(G20), .ZN(new_n220));
  NAND2_X1  g0020(.A1(new_n220), .A2(KEYINPUT67), .ZN(new_n221));
  INV_X1    g0021(.A(KEYINPUT67), .ZN(new_n222));
  NAND2_X1  g0022(.A1(new_n222), .A2(G20), .ZN(new_n223));
  NAND2_X1  g0023(.A1(new_n221), .A2(new_n223), .ZN(new_n224));
  NOR3_X1   g0024(.A1(new_n218), .A2(new_n219), .A3(new_n224), .ZN(new_n225));
  NAND2_X1  g0025(.A1(G1), .A2(G20), .ZN(new_n226));
  NOR2_X1   g0026(.A1(new_n226), .A2(G13), .ZN(new_n227));
  OAI211_X1 g0027(.A(new_n227), .B(G250), .C1(G257), .C2(G264), .ZN(new_n228));
  XOR2_X1   g0028(.A(new_n228), .B(KEYINPUT0), .Z(new_n229));
  AOI22_X1  g0029(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n230));
  XOR2_X1   g0030(.A(new_n230), .B(KEYINPUT70), .Z(new_n231));
  INV_X1    g0031(.A(G232), .ZN(new_n232));
  INV_X1    g0032(.A(G107), .ZN(new_n233));
  INV_X1    g0033(.A(G264), .ZN(new_n234));
  OAI22_X1  g0034(.A1(new_n201), .A2(new_n232), .B1(new_n233), .B2(new_n234), .ZN(new_n235));
  AOI21_X1  g0035(.A(new_n235), .B1(G68), .B2(G238), .ZN(new_n236));
  AOI22_X1  g0036(.A1(G77), .A2(G244), .B1(G116), .B2(G270), .ZN(new_n237));
  NAND3_X1  g0037(.A1(new_n231), .A2(new_n236), .A3(new_n237), .ZN(new_n238));
  INV_X1    g0038(.A(G226), .ZN(new_n239));
  NOR2_X1   g0039(.A1(new_n207), .A2(new_n239), .ZN(new_n240));
  OAI21_X1  g0040(.A(new_n226), .B1(new_n238), .B2(new_n240), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n241), .B(KEYINPUT1), .ZN(new_n242));
  NOR3_X1   g0042(.A1(new_n225), .A2(new_n229), .A3(new_n242), .ZN(G361));
  XNOR2_X1  g0043(.A(G238), .B(G244), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n244), .B(new_n232), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n245), .B(KEYINPUT2), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n246), .B(new_n239), .ZN(new_n247));
  XNOR2_X1  g0047(.A(G250), .B(G257), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n248), .B(new_n234), .ZN(new_n249));
  XNOR2_X1  g0049(.A(new_n249), .B(G270), .ZN(new_n250));
  XNOR2_X1  g0050(.A(new_n247), .B(new_n250), .ZN(G358));
  XNOR2_X1  g0051(.A(G50), .B(G68), .ZN(new_n252));
  XNOR2_X1  g0052(.A(new_n252), .B(KEYINPUT71), .ZN(new_n253));
  XNOR2_X1  g0053(.A(new_n253), .B(G58), .ZN(new_n254));
  XNOR2_X1  g0054(.A(new_n254), .B(new_n211), .ZN(new_n255));
  XNOR2_X1  g0055(.A(G107), .B(G116), .ZN(new_n256));
  XNOR2_X1  g0056(.A(new_n256), .B(KEYINPUT72), .ZN(new_n257));
  XOR2_X1   g0057(.A(G87), .B(G97), .Z(new_n258));
  XOR2_X1   g0058(.A(new_n257), .B(new_n258), .Z(new_n259));
  XNOR2_X1  g0059(.A(new_n255), .B(new_n259), .ZN(G351));
  AND2_X1   g0060(.A1(KEYINPUT3), .A2(G33), .ZN(new_n261));
  NOR2_X1   g0061(.A1(KEYINPUT3), .A2(G33), .ZN(new_n262));
  NOR2_X1   g0062(.A1(new_n261), .A2(new_n262), .ZN(new_n263));
  NOR2_X1   g0063(.A1(new_n263), .A2(G1698), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n264), .A2(G226), .ZN(new_n265));
  INV_X1    g0065(.A(G1698), .ZN(new_n266));
  NOR2_X1   g0066(.A1(new_n263), .A2(new_n266), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n267), .A2(G232), .ZN(new_n268));
  NAND2_X1  g0068(.A1(G33), .A2(G97), .ZN(new_n269));
  NAND3_X1  g0069(.A1(new_n265), .A2(new_n268), .A3(new_n269), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n270), .A2(KEYINPUT76), .ZN(new_n271));
  AOI21_X1  g0071(.A(new_n219), .B1(G33), .B2(G41), .ZN(new_n272));
  INV_X1    g0072(.A(KEYINPUT76), .ZN(new_n273));
  NAND4_X1  g0073(.A1(new_n265), .A2(new_n268), .A3(new_n273), .A4(new_n269), .ZN(new_n274));
  NAND3_X1  g0074(.A1(new_n271), .A2(new_n272), .A3(new_n274), .ZN(new_n275));
  INV_X1    g0075(.A(G1), .ZN(new_n276));
  OAI21_X1  g0076(.A(new_n276), .B1(G41), .B2(G45), .ZN(new_n277));
  INV_X1    g0077(.A(G274), .ZN(new_n278));
  NOR2_X1   g0078(.A1(new_n277), .A2(new_n278), .ZN(new_n279));
  NAND2_X1  g0079(.A1(new_n277), .A2(KEYINPUT73), .ZN(new_n280));
  INV_X1    g0080(.A(KEYINPUT73), .ZN(new_n281));
  OAI211_X1 g0081(.A(new_n281), .B(new_n276), .C1(G41), .C2(G45), .ZN(new_n282));
  AOI21_X1  g0082(.A(new_n272), .B1(new_n280), .B2(new_n282), .ZN(new_n283));
  AOI21_X1  g0083(.A(new_n279), .B1(new_n283), .B2(G238), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n275), .A2(new_n284), .ZN(new_n285));
  INV_X1    g0085(.A(KEYINPUT13), .ZN(new_n286));
  XNOR2_X1  g0086(.A(new_n285), .B(new_n286), .ZN(new_n287));
  INV_X1    g0087(.A(G169), .ZN(new_n288));
  OAI21_X1  g0088(.A(KEYINPUT14), .B1(new_n287), .B2(new_n288), .ZN(new_n289));
  XNOR2_X1  g0089(.A(new_n285), .B(KEYINPUT13), .ZN(new_n290));
  INV_X1    g0090(.A(KEYINPUT14), .ZN(new_n291));
  NAND3_X1  g0091(.A1(new_n290), .A2(new_n291), .A3(G169), .ZN(new_n292));
  INV_X1    g0092(.A(G179), .ZN(new_n293));
  OAI211_X1 g0093(.A(new_n289), .B(new_n292), .C1(new_n293), .C2(new_n290), .ZN(new_n294));
  NOR2_X1   g0094(.A1(G20), .A2(G33), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n295), .A2(G50), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n224), .A2(G33), .ZN(new_n297));
  OAI221_X1 g0097(.A(new_n296), .B1(new_n220), .B2(G68), .C1(new_n297), .C2(new_n211), .ZN(new_n298));
  NAND3_X1  g0098(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n299), .A2(new_n219), .ZN(new_n300));
  NAND3_X1  g0100(.A1(new_n298), .A2(KEYINPUT11), .A3(new_n300), .ZN(new_n301));
  INV_X1    g0101(.A(new_n300), .ZN(new_n302));
  OAI21_X1  g0102(.A(new_n302), .B1(G1), .B2(new_n220), .ZN(new_n303));
  OAI21_X1  g0103(.A(new_n301), .B1(new_n202), .B2(new_n303), .ZN(new_n304));
  INV_X1    g0104(.A(G13), .ZN(new_n305));
  NOR3_X1   g0105(.A1(new_n305), .A2(new_n220), .A3(G1), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n306), .A2(new_n202), .ZN(new_n307));
  XOR2_X1   g0107(.A(new_n307), .B(KEYINPUT12), .Z(new_n308));
  AOI21_X1  g0108(.A(KEYINPUT11), .B1(new_n298), .B2(new_n300), .ZN(new_n309));
  NOR3_X1   g0109(.A1(new_n304), .A2(new_n308), .A3(new_n309), .ZN(new_n310));
  INV_X1    g0110(.A(new_n310), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n294), .A2(new_n311), .ZN(new_n312));
  INV_X1    g0112(.A(KEYINPUT3), .ZN(new_n313));
  INV_X1    g0113(.A(G33), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n313), .A2(new_n314), .ZN(new_n315));
  NAND2_X1  g0115(.A1(KEYINPUT3), .A2(G33), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n315), .A2(new_n316), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n317), .A2(new_n266), .ZN(new_n318));
  OAI21_X1  g0118(.A(KEYINPUT74), .B1(new_n318), .B2(new_n232), .ZN(new_n319));
  INV_X1    g0119(.A(KEYINPUT74), .ZN(new_n320));
  NAND3_X1  g0120(.A1(new_n264), .A2(new_n320), .A3(G232), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n263), .A2(G107), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n267), .A2(G238), .ZN(new_n323));
  NAND4_X1  g0123(.A1(new_n319), .A2(new_n321), .A3(new_n322), .A4(new_n323), .ZN(new_n324));
  AOI21_X1  g0124(.A(new_n279), .B1(new_n324), .B2(new_n272), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n283), .A2(G244), .ZN(new_n326));
  AOI21_X1  g0126(.A(G169), .B1(new_n325), .B2(new_n326), .ZN(new_n327));
  XOR2_X1   g0127(.A(KEYINPUT8), .B(G58), .Z(new_n328));
  NAND2_X1  g0128(.A1(new_n328), .A2(new_n295), .ZN(new_n329));
  XNOR2_X1  g0129(.A(KEYINPUT15), .B(G87), .ZN(new_n330));
  OAI221_X1 g0130(.A(new_n329), .B1(new_n211), .B2(new_n224), .C1(new_n297), .C2(new_n330), .ZN(new_n331));
  AOI22_X1  g0131(.A1(new_n331), .A2(new_n300), .B1(new_n211), .B2(new_n306), .ZN(new_n332));
  INV_X1    g0132(.A(new_n303), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n333), .A2(G77), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n332), .A2(new_n334), .ZN(new_n335));
  INV_X1    g0135(.A(new_n335), .ZN(new_n336));
  OAI21_X1  g0136(.A(KEYINPUT75), .B1(new_n327), .B2(new_n336), .ZN(new_n337));
  INV_X1    g0137(.A(new_n326), .ZN(new_n338));
  AOI211_X1 g0138(.A(new_n279), .B(new_n338), .C1(new_n324), .C2(new_n272), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n339), .A2(new_n293), .ZN(new_n340));
  INV_X1    g0140(.A(KEYINPUT75), .ZN(new_n341));
  OAI211_X1 g0141(.A(new_n335), .B(new_n341), .C1(new_n339), .C2(G169), .ZN(new_n342));
  NAND3_X1  g0142(.A1(new_n337), .A2(new_n340), .A3(new_n342), .ZN(new_n343));
  INV_X1    g0143(.A(new_n343), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n339), .A2(G190), .ZN(new_n345));
  INV_X1    g0145(.A(G200), .ZN(new_n346));
  OAI211_X1 g0146(.A(new_n345), .B(new_n336), .C1(new_n346), .C2(new_n339), .ZN(new_n347));
  INV_X1    g0147(.A(new_n347), .ZN(new_n348));
  NOR2_X1   g0148(.A1(new_n344), .A2(new_n348), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n287), .A2(G190), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n290), .A2(G200), .ZN(new_n351));
  NAND3_X1  g0151(.A1(new_n350), .A2(new_n351), .A3(new_n310), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n295), .A2(G150), .ZN(new_n353));
  INV_X1    g0153(.A(new_n328), .ZN(new_n354));
  OAI221_X1 g0154(.A(new_n353), .B1(new_n354), .B2(new_n297), .C1(new_n210), .C2(new_n220), .ZN(new_n355));
  AOI22_X1  g0155(.A1(new_n355), .A2(new_n300), .B1(new_n207), .B2(new_n306), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n333), .A2(G50), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n356), .A2(new_n357), .ZN(new_n358));
  AOI22_X1  g0158(.A1(new_n264), .A2(G222), .B1(G77), .B2(new_n263), .ZN(new_n359));
  INV_X1    g0159(.A(G223), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n317), .A2(G1698), .ZN(new_n361));
  OAI21_X1  g0161(.A(new_n359), .B1(new_n360), .B2(new_n361), .ZN(new_n362));
  AOI21_X1  g0162(.A(new_n279), .B1(new_n362), .B2(new_n272), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n283), .A2(G226), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n363), .A2(new_n364), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n365), .A2(new_n288), .ZN(new_n366));
  OAI211_X1 g0166(.A(new_n358), .B(new_n366), .C1(G179), .C2(new_n365), .ZN(new_n367));
  NAND4_X1  g0167(.A1(new_n312), .A2(new_n349), .A3(new_n352), .A4(new_n367), .ZN(new_n368));
  INV_X1    g0168(.A(new_n358), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n369), .A2(KEYINPUT9), .ZN(new_n370));
  NAND3_X1  g0170(.A1(new_n363), .A2(G190), .A3(new_n364), .ZN(new_n371));
  INV_X1    g0171(.A(KEYINPUT9), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n358), .A2(new_n372), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n365), .A2(G200), .ZN(new_n374));
  NAND4_X1  g0174(.A1(new_n370), .A2(new_n371), .A3(new_n373), .A4(new_n374), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n375), .A2(KEYINPUT10), .ZN(new_n376));
  AOI22_X1  g0176(.A1(new_n369), .A2(KEYINPUT9), .B1(G200), .B2(new_n365), .ZN(new_n377));
  INV_X1    g0177(.A(KEYINPUT10), .ZN(new_n378));
  NAND4_X1  g0178(.A1(new_n377), .A2(new_n378), .A3(new_n371), .A4(new_n373), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n376), .A2(new_n379), .ZN(new_n380));
  NOR3_X1   g0180(.A1(new_n261), .A2(new_n262), .A3(KEYINPUT77), .ZN(new_n381));
  INV_X1    g0181(.A(KEYINPUT77), .ZN(new_n382));
  AOI21_X1  g0182(.A(new_n382), .B1(new_n315), .B2(new_n316), .ZN(new_n383));
  OAI21_X1  g0183(.A(new_n224), .B1(new_n381), .B2(new_n383), .ZN(new_n384));
  INV_X1    g0184(.A(KEYINPUT7), .ZN(new_n385));
  NAND3_X1  g0185(.A1(new_n384), .A2(KEYINPUT78), .A3(new_n385), .ZN(new_n386));
  INV_X1    g0186(.A(KEYINPUT78), .ZN(new_n387));
  XNOR2_X1  g0187(.A(KEYINPUT67), .B(G20), .ZN(new_n388));
  OAI21_X1  g0188(.A(KEYINPUT77), .B1(new_n261), .B2(new_n262), .ZN(new_n389));
  NAND3_X1  g0189(.A1(new_n315), .A2(new_n382), .A3(new_n316), .ZN(new_n390));
  AOI21_X1  g0190(.A(new_n388), .B1(new_n389), .B2(new_n390), .ZN(new_n391));
  OAI21_X1  g0191(.A(new_n387), .B1(new_n391), .B2(KEYINPUT7), .ZN(new_n392));
  NAND3_X1  g0192(.A1(new_n263), .A2(KEYINPUT7), .A3(new_n220), .ZN(new_n393));
  NAND3_X1  g0193(.A1(new_n386), .A2(new_n392), .A3(new_n393), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n394), .A2(G68), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n295), .A2(G159), .ZN(new_n396));
  XNOR2_X1  g0196(.A(new_n396), .B(KEYINPUT79), .ZN(new_n397));
  NOR2_X1   g0197(.A1(new_n201), .A2(new_n202), .ZN(new_n398));
  OAI21_X1  g0198(.A(G20), .B1(new_n206), .B2(new_n398), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n397), .A2(new_n399), .ZN(new_n400));
  INV_X1    g0200(.A(new_n400), .ZN(new_n401));
  NAND3_X1  g0201(.A1(new_n395), .A2(KEYINPUT16), .A3(new_n401), .ZN(new_n402));
  INV_X1    g0202(.A(KEYINPUT16), .ZN(new_n403));
  NOR3_X1   g0203(.A1(new_n317), .A2(new_n388), .A3(new_n385), .ZN(new_n404));
  AOI21_X1  g0204(.A(KEYINPUT7), .B1(new_n263), .B2(new_n220), .ZN(new_n405));
  NOR2_X1   g0205(.A1(new_n404), .A2(new_n405), .ZN(new_n406));
  NOR2_X1   g0206(.A1(new_n406), .A2(new_n202), .ZN(new_n407));
  OAI21_X1  g0207(.A(new_n403), .B1(new_n407), .B2(new_n400), .ZN(new_n408));
  NAND3_X1  g0208(.A1(new_n402), .A2(new_n408), .A3(new_n300), .ZN(new_n409));
  NOR2_X1   g0209(.A1(new_n328), .A2(new_n306), .ZN(new_n410));
  AOI21_X1  g0210(.A(new_n410), .B1(new_n328), .B2(new_n303), .ZN(new_n411));
  INV_X1    g0211(.A(new_n411), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n409), .A2(new_n412), .ZN(new_n413));
  NAND3_X1  g0213(.A1(new_n317), .A2(G223), .A3(new_n266), .ZN(new_n414));
  NAND2_X1  g0214(.A1(G33), .A2(G87), .ZN(new_n415));
  OAI211_X1 g0215(.A(new_n414), .B(new_n415), .C1(new_n361), .C2(new_n239), .ZN(new_n416));
  AOI21_X1  g0216(.A(new_n279), .B1(new_n416), .B2(new_n272), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n283), .A2(G232), .ZN(new_n418));
  AOI21_X1  g0218(.A(new_n288), .B1(new_n417), .B2(new_n418), .ZN(new_n419));
  AND2_X1   g0219(.A1(new_n417), .A2(new_n418), .ZN(new_n420));
  AOI21_X1  g0220(.A(new_n419), .B1(G179), .B2(new_n420), .ZN(new_n421));
  INV_X1    g0221(.A(new_n421), .ZN(new_n422));
  AOI21_X1  g0222(.A(KEYINPUT18), .B1(new_n413), .B2(new_n422), .ZN(new_n423));
  INV_X1    g0223(.A(KEYINPUT18), .ZN(new_n424));
  AOI211_X1 g0224(.A(new_n424), .B(new_n421), .C1(new_n409), .C2(new_n412), .ZN(new_n425));
  NOR2_X1   g0225(.A1(new_n423), .A2(new_n425), .ZN(new_n426));
  INV_X1    g0226(.A(KEYINPUT80), .ZN(new_n427));
  INV_X1    g0227(.A(KEYINPUT17), .ZN(new_n428));
  AOI21_X1  g0228(.A(new_n400), .B1(new_n394), .B2(G68), .ZN(new_n429));
  AOI21_X1  g0229(.A(new_n302), .B1(new_n429), .B2(KEYINPUT16), .ZN(new_n430));
  AOI21_X1  g0230(.A(new_n411), .B1(new_n430), .B2(new_n408), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n417), .A2(new_n418), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n432), .A2(new_n346), .ZN(new_n433));
  OAI21_X1  g0233(.A(new_n433), .B1(G190), .B2(new_n432), .ZN(new_n434));
  AOI21_X1  g0234(.A(new_n428), .B1(new_n431), .B2(new_n434), .ZN(new_n435));
  NAND4_X1  g0235(.A1(new_n409), .A2(new_n428), .A3(new_n412), .A4(new_n434), .ZN(new_n436));
  INV_X1    g0236(.A(new_n436), .ZN(new_n437));
  OAI21_X1  g0237(.A(new_n427), .B1(new_n435), .B2(new_n437), .ZN(new_n438));
  NAND3_X1  g0238(.A1(new_n409), .A2(new_n412), .A3(new_n434), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n439), .A2(KEYINPUT17), .ZN(new_n440));
  NAND3_X1  g0240(.A1(new_n440), .A2(KEYINPUT80), .A3(new_n436), .ZN(new_n441));
  AOI21_X1  g0241(.A(new_n426), .B1(new_n438), .B2(new_n441), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n380), .A2(new_n442), .ZN(new_n443));
  NOR2_X1   g0243(.A1(new_n368), .A2(new_n443), .ZN(new_n444));
  INV_X1    g0244(.A(new_n306), .ZN(new_n445));
  NOR2_X1   g0245(.A1(new_n445), .A2(G97), .ZN(new_n446));
  OAI211_X1 g0246(.A(new_n445), .B(new_n302), .C1(G1), .C2(new_n314), .ZN(new_n447));
  INV_X1    g0247(.A(G97), .ZN(new_n448));
  NOR2_X1   g0248(.A1(new_n447), .A2(new_n448), .ZN(new_n449));
  NAND3_X1  g0249(.A1(new_n233), .A2(KEYINPUT6), .A3(G97), .ZN(new_n450));
  XOR2_X1   g0250(.A(G97), .B(G107), .Z(new_n451));
  OAI21_X1  g0251(.A(new_n450), .B1(new_n451), .B2(KEYINPUT6), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n295), .A2(G77), .ZN(new_n453));
  AOI22_X1  g0253(.A1(new_n452), .A2(new_n388), .B1(KEYINPUT81), .B2(new_n453), .ZN(new_n454));
  OR2_X1    g0254(.A1(new_n453), .A2(KEYINPUT81), .ZN(new_n455));
  OAI211_X1 g0255(.A(new_n454), .B(new_n455), .C1(new_n233), .C2(new_n406), .ZN(new_n456));
  AOI211_X1 g0256(.A(new_n446), .B(new_n449), .C1(new_n456), .C2(new_n300), .ZN(new_n457));
  INV_X1    g0257(.A(new_n272), .ZN(new_n458));
  INV_X1    g0258(.A(G45), .ZN(new_n459));
  NOR2_X1   g0259(.A1(new_n459), .A2(G1), .ZN(new_n460));
  AND2_X1   g0260(.A1(KEYINPUT5), .A2(G41), .ZN(new_n461));
  NOR2_X1   g0261(.A1(KEYINPUT5), .A2(G41), .ZN(new_n462));
  OAI21_X1  g0262(.A(new_n460), .B1(new_n461), .B2(new_n462), .ZN(new_n463));
  AND2_X1   g0263(.A1(new_n458), .A2(new_n463), .ZN(new_n464));
  NAND2_X1  g0264(.A1(new_n464), .A2(G257), .ZN(new_n465));
  OR2_X1    g0265(.A1(new_n463), .A2(new_n278), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  INV_X1    g0267(.A(KEYINPUT82), .ZN(new_n468));
  NOR2_X1   g0268(.A1(new_n468), .A2(KEYINPUT4), .ZN(new_n469));
  INV_X1    g0269(.A(G244), .ZN(new_n470));
  OAI21_X1  g0270(.A(new_n469), .B1(new_n318), .B2(new_n470), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n267), .A2(G250), .ZN(new_n472));
  INV_X1    g0272(.A(new_n469), .ZN(new_n473));
  NAND4_X1  g0273(.A1(new_n317), .A2(new_n473), .A3(G244), .A4(new_n266), .ZN(new_n474));
  NAND2_X1  g0274(.A1(G33), .A2(G283), .ZN(new_n475));
  NAND4_X1  g0275(.A1(new_n471), .A2(new_n472), .A3(new_n474), .A4(new_n475), .ZN(new_n476));
  AOI21_X1  g0276(.A(new_n467), .B1(new_n272), .B2(new_n476), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n477), .A2(G190), .ZN(new_n478));
  AND3_X1   g0278(.A1(new_n476), .A2(KEYINPUT83), .A3(new_n272), .ZN(new_n479));
  AOI21_X1  g0279(.A(KEYINPUT83), .B1(new_n476), .B2(new_n272), .ZN(new_n480));
  NOR3_X1   g0280(.A1(new_n479), .A2(new_n480), .A3(new_n467), .ZN(new_n481));
  OAI211_X1 g0281(.A(new_n457), .B(new_n478), .C1(new_n481), .C2(new_n346), .ZN(new_n482));
  OR2_X1    g0282(.A1(new_n477), .A2(G169), .ZN(new_n483));
  AOI21_X1  g0283(.A(new_n446), .B1(new_n456), .B2(new_n300), .ZN(new_n484));
  INV_X1    g0284(.A(new_n449), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n484), .A2(new_n485), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n476), .A2(new_n272), .ZN(new_n487));
  INV_X1    g0287(.A(KEYINPUT83), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n487), .A2(new_n488), .ZN(new_n489));
  INV_X1    g0289(.A(new_n467), .ZN(new_n490));
  NAND3_X1  g0290(.A1(new_n476), .A2(KEYINPUT83), .A3(new_n272), .ZN(new_n491));
  NAND4_X1  g0291(.A1(new_n489), .A2(new_n293), .A3(new_n490), .A4(new_n491), .ZN(new_n492));
  NAND3_X1  g0292(.A1(new_n483), .A2(new_n486), .A3(new_n492), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n482), .A2(new_n493), .ZN(new_n494));
  NAND2_X1  g0294(.A1(KEYINPUT23), .A2(G107), .ZN(new_n495));
  NAND2_X1  g0295(.A1(G33), .A2(G116), .ZN(new_n496));
  INV_X1    g0296(.A(KEYINPUT23), .ZN(new_n497));
  AOI21_X1  g0297(.A(G20), .B1(new_n496), .B2(new_n497), .ZN(new_n498));
  NOR2_X1   g0298(.A1(new_n224), .A2(KEYINPUT23), .ZN(new_n499));
  AOI21_X1  g0299(.A(new_n498), .B1(new_n499), .B2(new_n233), .ZN(new_n500));
  INV_X1    g0300(.A(KEYINPUT22), .ZN(new_n501));
  NOR2_X1   g0301(.A1(new_n263), .A2(new_n388), .ZN(new_n502));
  AOI21_X1  g0302(.A(new_n501), .B1(new_n502), .B2(G87), .ZN(new_n503));
  NAND3_X1  g0303(.A1(new_n224), .A2(new_n317), .A3(G87), .ZN(new_n504));
  NOR2_X1   g0304(.A1(new_n504), .A2(KEYINPUT22), .ZN(new_n505));
  OAI211_X1 g0305(.A(new_n495), .B(new_n500), .C1(new_n503), .C2(new_n505), .ZN(new_n506));
  INV_X1    g0306(.A(KEYINPUT90), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  XNOR2_X1  g0308(.A(new_n504), .B(KEYINPUT22), .ZN(new_n509));
  NAND4_X1  g0309(.A1(new_n509), .A2(KEYINPUT90), .A3(new_n495), .A4(new_n500), .ZN(new_n510));
  XNOR2_X1  g0310(.A(KEYINPUT89), .B(KEYINPUT24), .ZN(new_n511));
  NAND3_X1  g0311(.A1(new_n508), .A2(new_n510), .A3(new_n511), .ZN(new_n512));
  INV_X1    g0312(.A(new_n511), .ZN(new_n513));
  NAND3_X1  g0313(.A1(new_n506), .A2(new_n507), .A3(new_n513), .ZN(new_n514));
  NAND3_X1  g0314(.A1(new_n512), .A2(new_n300), .A3(new_n514), .ZN(new_n515));
  AOI22_X1  g0315(.A1(G250), .A2(new_n264), .B1(new_n267), .B2(G257), .ZN(new_n516));
  INV_X1    g0316(.A(G294), .ZN(new_n517));
  OAI21_X1  g0317(.A(new_n516), .B1(new_n314), .B2(new_n517), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n518), .A2(new_n272), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n464), .A2(G264), .ZN(new_n520));
  NAND4_X1  g0320(.A1(new_n519), .A2(G190), .A3(new_n466), .A4(new_n520), .ZN(new_n521));
  INV_X1    g0321(.A(new_n447), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n522), .A2(G107), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n306), .A2(new_n233), .ZN(new_n524));
  XOR2_X1   g0324(.A(new_n524), .B(KEYINPUT25), .Z(new_n525));
  NAND4_X1  g0325(.A1(new_n515), .A2(new_n521), .A3(new_n523), .A4(new_n525), .ZN(new_n526));
  INV_X1    g0326(.A(new_n526), .ZN(new_n527));
  AND2_X1   g0327(.A1(new_n519), .A2(new_n520), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n528), .A2(new_n466), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n529), .A2(G200), .ZN(new_n530));
  AOI21_X1  g0330(.A(new_n494), .B1(new_n527), .B2(new_n530), .ZN(new_n531));
  NAND3_X1  g0331(.A1(new_n515), .A2(new_n523), .A3(new_n525), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n529), .A2(new_n288), .ZN(new_n533));
  NAND3_X1  g0333(.A1(new_n528), .A2(new_n293), .A3(new_n466), .ZN(new_n534));
  NAND3_X1  g0334(.A1(new_n532), .A2(new_n533), .A3(new_n534), .ZN(new_n535));
  AND2_X1   g0335(.A1(new_n531), .A2(new_n535), .ZN(new_n536));
  INV_X1    g0336(.A(KEYINPUT85), .ZN(new_n537));
  AND2_X1   g0337(.A1(KEYINPUT84), .A2(KEYINPUT19), .ZN(new_n538));
  NOR2_X1   g0338(.A1(KEYINPUT84), .A2(KEYINPUT19), .ZN(new_n539));
  NOR3_X1   g0339(.A1(new_n538), .A2(new_n539), .A3(new_n269), .ZN(new_n540));
  OAI21_X1  g0340(.A(new_n537), .B1(new_n540), .B2(new_n388), .ZN(new_n541));
  INV_X1    g0341(.A(G87), .ZN(new_n542));
  NAND3_X1  g0342(.A1(new_n542), .A2(new_n448), .A3(new_n233), .ZN(new_n543));
  XNOR2_X1  g0343(.A(KEYINPUT84), .B(KEYINPUT19), .ZN(new_n544));
  OAI211_X1 g0344(.A(new_n224), .B(KEYINPUT85), .C1(new_n544), .C2(new_n269), .ZN(new_n545));
  NAND3_X1  g0345(.A1(new_n541), .A2(new_n543), .A3(new_n545), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n502), .A2(G68), .ZN(new_n547));
  OAI21_X1  g0347(.A(new_n544), .B1(new_n297), .B2(new_n448), .ZN(new_n548));
  NAND3_X1  g0348(.A1(new_n546), .A2(new_n547), .A3(new_n548), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n549), .A2(KEYINPUT86), .ZN(new_n550));
  INV_X1    g0350(.A(KEYINPUT86), .ZN(new_n551));
  NAND4_X1  g0351(.A1(new_n546), .A2(new_n551), .A3(new_n547), .A4(new_n548), .ZN(new_n552));
  NAND3_X1  g0352(.A1(new_n550), .A2(new_n300), .A3(new_n552), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n330), .A2(new_n306), .ZN(new_n554));
  INV_X1    g0354(.A(new_n330), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n522), .A2(new_n555), .ZN(new_n556));
  NAND3_X1  g0356(.A1(new_n553), .A2(new_n554), .A3(new_n556), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n557), .A2(KEYINPUT87), .ZN(new_n558));
  INV_X1    g0358(.A(KEYINPUT87), .ZN(new_n559));
  NAND4_X1  g0359(.A1(new_n553), .A2(new_n559), .A3(new_n554), .A4(new_n556), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n558), .A2(new_n560), .ZN(new_n561));
  INV_X1    g0361(.A(G238), .ZN(new_n562));
  OAI221_X1 g0362(.A(new_n496), .B1(new_n361), .B2(new_n470), .C1(new_n562), .C2(new_n318), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n563), .A2(new_n272), .ZN(new_n564));
  OAI211_X1 g0364(.A(new_n458), .B(G250), .C1(G1), .C2(new_n459), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n460), .A2(G274), .ZN(new_n566));
  NAND3_X1  g0366(.A1(new_n564), .A2(new_n565), .A3(new_n566), .ZN(new_n567));
  INV_X1    g0367(.A(new_n567), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n568), .A2(new_n293), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n567), .A2(new_n288), .ZN(new_n570));
  NAND3_X1  g0370(.A1(new_n561), .A2(new_n569), .A3(new_n570), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n553), .A2(new_n554), .ZN(new_n572));
  AOI21_X1  g0372(.A(new_n572), .B1(G87), .B2(new_n522), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n568), .A2(G190), .ZN(new_n574));
  OAI211_X1 g0374(.A(new_n573), .B(new_n574), .C1(new_n346), .C2(new_n568), .ZN(new_n575));
  AND2_X1   g0375(.A1(new_n571), .A2(new_n575), .ZN(new_n576));
  INV_X1    g0376(.A(G116), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n306), .A2(new_n577), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n522), .A2(G116), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n577), .A2(G20), .ZN(new_n580));
  AND3_X1   g0380(.A1(new_n300), .A2(KEYINPUT88), .A3(new_n580), .ZN(new_n581));
  AOI21_X1  g0381(.A(KEYINPUT88), .B1(new_n300), .B2(new_n580), .ZN(new_n582));
  OR2_X1    g0382(.A1(new_n581), .A2(new_n582), .ZN(new_n583));
  OAI211_X1 g0383(.A(new_n224), .B(new_n475), .C1(G33), .C2(new_n448), .ZN(new_n584));
  AOI21_X1  g0384(.A(KEYINPUT20), .B1(new_n583), .B2(new_n584), .ZN(new_n585));
  OAI211_X1 g0385(.A(new_n584), .B(KEYINPUT20), .C1(new_n581), .C2(new_n582), .ZN(new_n586));
  INV_X1    g0386(.A(new_n586), .ZN(new_n587));
  OAI211_X1 g0387(.A(new_n578), .B(new_n579), .C1(new_n585), .C2(new_n587), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n464), .A2(G270), .ZN(new_n589));
  INV_X1    g0389(.A(G303), .ZN(new_n590));
  OAI22_X1  g0390(.A1(new_n361), .A2(new_n234), .B1(new_n590), .B2(new_n317), .ZN(new_n591));
  AOI21_X1  g0391(.A(new_n591), .B1(G257), .B2(new_n264), .ZN(new_n592));
  OAI211_X1 g0392(.A(new_n466), .B(new_n589), .C1(new_n592), .C2(new_n458), .ZN(new_n593));
  NAND3_X1  g0393(.A1(new_n588), .A2(G169), .A3(new_n593), .ZN(new_n594));
  INV_X1    g0394(.A(KEYINPUT21), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n594), .A2(new_n595), .ZN(new_n596));
  NOR2_X1   g0396(.A1(new_n593), .A2(new_n293), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n597), .A2(new_n588), .ZN(new_n598));
  NAND4_X1  g0398(.A1(new_n588), .A2(new_n593), .A3(KEYINPUT21), .A4(G169), .ZN(new_n599));
  AND3_X1   g0399(.A1(new_n596), .A2(new_n598), .A3(new_n599), .ZN(new_n600));
  INV_X1    g0400(.A(new_n600), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n593), .A2(G200), .ZN(new_n602));
  INV_X1    g0402(.A(G190), .ZN(new_n603));
  OAI21_X1  g0403(.A(new_n602), .B1(new_n603), .B2(new_n593), .ZN(new_n604));
  NOR2_X1   g0404(.A1(new_n604), .A2(new_n588), .ZN(new_n605));
  NOR2_X1   g0405(.A1(new_n601), .A2(new_n605), .ZN(new_n606));
  NAND4_X1  g0406(.A1(new_n444), .A2(new_n536), .A3(new_n576), .A4(new_n606), .ZN(new_n607));
  XNOR2_X1  g0407(.A(new_n607), .B(KEYINPUT91), .ZN(G372));
  INV_X1    g0408(.A(new_n367), .ZN(new_n609));
  INV_X1    g0409(.A(new_n352), .ZN(new_n610));
  AOI21_X1  g0410(.A(new_n610), .B1(new_n312), .B2(new_n343), .ZN(new_n611));
  AND3_X1   g0411(.A1(new_n440), .A2(KEYINPUT80), .A3(new_n436), .ZN(new_n612));
  AOI21_X1  g0412(.A(KEYINPUT80), .B1(new_n440), .B2(new_n436), .ZN(new_n613));
  OAI21_X1  g0413(.A(new_n611), .B1(new_n612), .B2(new_n613), .ZN(new_n614));
  OR2_X1    g0414(.A1(new_n423), .A2(new_n425), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  INV_X1    g0416(.A(KEYINPUT94), .ZN(new_n617));
  XNOR2_X1  g0417(.A(new_n380), .B(new_n617), .ZN(new_n618));
  AOI21_X1  g0418(.A(new_n609), .B1(new_n616), .B2(new_n618), .ZN(new_n619));
  INV_X1    g0419(.A(new_n493), .ZN(new_n620));
  NAND3_X1  g0420(.A1(new_n571), .A2(new_n575), .A3(new_n620), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n621), .A2(KEYINPUT26), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n535), .A2(new_n600), .ZN(new_n623));
  OR2_X1    g0423(.A1(new_n570), .A2(KEYINPUT92), .ZN(new_n624));
  AOI22_X1  g0424(.A1(new_n570), .A2(KEYINPUT92), .B1(new_n568), .B2(new_n293), .ZN(new_n625));
  NAND3_X1  g0425(.A1(new_n561), .A2(new_n624), .A3(new_n625), .ZN(new_n626));
  NAND4_X1  g0426(.A1(new_n531), .A2(new_n575), .A3(new_n623), .A4(new_n626), .ZN(new_n627));
  INV_X1    g0427(.A(KEYINPUT93), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n626), .A2(new_n628), .ZN(new_n629));
  NAND4_X1  g0429(.A1(new_n561), .A2(KEYINPUT93), .A3(new_n624), .A4(new_n625), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  INV_X1    g0431(.A(KEYINPUT26), .ZN(new_n632));
  NAND4_X1  g0432(.A1(new_n626), .A2(new_n575), .A3(new_n632), .A4(new_n620), .ZN(new_n633));
  NAND4_X1  g0433(.A1(new_n622), .A2(new_n627), .A3(new_n631), .A4(new_n633), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n444), .A2(new_n634), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n619), .A2(new_n635), .ZN(G369));
  NOR2_X1   g0436(.A1(new_n388), .A2(new_n305), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n637), .A2(new_n276), .ZN(new_n638));
  OR2_X1    g0438(.A1(new_n638), .A2(KEYINPUT27), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n638), .A2(KEYINPUT27), .ZN(new_n640));
  NAND3_X1  g0440(.A1(new_n639), .A2(G213), .A3(new_n640), .ZN(new_n641));
  INV_X1    g0441(.A(G343), .ZN(new_n642));
  NOR2_X1   g0442(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n588), .A2(new_n643), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n606), .A2(new_n644), .ZN(new_n645));
  OAI21_X1  g0445(.A(new_n645), .B1(new_n600), .B2(new_n644), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n646), .A2(G330), .ZN(new_n647));
  INV_X1    g0447(.A(KEYINPUT95), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n532), .A2(new_n643), .ZN(new_n649));
  INV_X1    g0449(.A(new_n530), .ZN(new_n650));
  OAI21_X1  g0450(.A(new_n649), .B1(new_n650), .B2(new_n526), .ZN(new_n651));
  INV_X1    g0451(.A(new_n535), .ZN(new_n652));
  OAI21_X1  g0452(.A(new_n648), .B1(new_n651), .B2(new_n652), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n527), .A2(new_n530), .ZN(new_n654));
  NAND4_X1  g0454(.A1(new_n654), .A2(KEYINPUT95), .A3(new_n535), .A4(new_n649), .ZN(new_n655));
  INV_X1    g0455(.A(KEYINPUT96), .ZN(new_n656));
  NAND3_X1  g0456(.A1(new_n652), .A2(new_n656), .A3(new_n643), .ZN(new_n657));
  INV_X1    g0457(.A(new_n643), .ZN(new_n658));
  OAI21_X1  g0458(.A(KEYINPUT96), .B1(new_n535), .B2(new_n658), .ZN(new_n659));
  AOI22_X1  g0459(.A1(new_n653), .A2(new_n655), .B1(new_n657), .B2(new_n659), .ZN(new_n660));
  NOR2_X1   g0460(.A1(new_n647), .A2(new_n660), .ZN(new_n661));
  INV_X1    g0461(.A(new_n661), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n653), .A2(new_n655), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n657), .A2(new_n659), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  NOR2_X1   g0465(.A1(new_n600), .A2(new_n643), .ZN(new_n666));
  AOI22_X1  g0466(.A1(new_n665), .A2(new_n666), .B1(new_n652), .B2(new_n658), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n662), .A2(new_n667), .ZN(G399));
  INV_X1    g0468(.A(new_n227), .ZN(new_n669));
  NOR2_X1   g0469(.A1(new_n669), .A2(G41), .ZN(new_n670));
  INV_X1    g0470(.A(new_n670), .ZN(new_n671));
  NOR2_X1   g0471(.A1(new_n543), .A2(G116), .ZN(new_n672));
  NAND3_X1  g0472(.A1(new_n671), .A2(G1), .A3(new_n672), .ZN(new_n673));
  INV_X1    g0473(.A(new_n216), .ZN(new_n674));
  OAI21_X1  g0474(.A(new_n673), .B1(new_n674), .B2(new_n671), .ZN(new_n675));
  XNOR2_X1  g0475(.A(new_n675), .B(KEYINPUT28), .ZN(new_n676));
  NAND3_X1  g0476(.A1(new_n576), .A2(new_n632), .A3(new_n620), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n626), .A2(new_n575), .ZN(new_n678));
  OAI21_X1  g0478(.A(KEYINPUT26), .B1(new_n678), .B2(new_n493), .ZN(new_n679));
  NAND4_X1  g0479(.A1(new_n677), .A2(new_n631), .A3(new_n679), .A4(new_n627), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n680), .A2(new_n658), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n681), .A2(KEYINPUT29), .ZN(new_n682));
  INV_X1    g0482(.A(KEYINPUT29), .ZN(new_n683));
  NAND3_X1  g0483(.A1(new_n634), .A2(new_n683), .A3(new_n658), .ZN(new_n684));
  INV_X1    g0484(.A(G330), .ZN(new_n685));
  NAND4_X1  g0485(.A1(new_n536), .A2(new_n576), .A3(new_n606), .A4(new_n658), .ZN(new_n686));
  NAND4_X1  g0486(.A1(new_n597), .A2(new_n528), .A3(new_n477), .A4(new_n568), .ZN(new_n687));
  XOR2_X1   g0487(.A(new_n687), .B(KEYINPUT30), .Z(new_n688));
  INV_X1    g0488(.A(new_n529), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n593), .A2(new_n293), .ZN(new_n690));
  NOR4_X1   g0490(.A1(new_n689), .A2(new_n481), .A3(new_n568), .A4(new_n690), .ZN(new_n691));
  OAI21_X1  g0491(.A(new_n643), .B1(new_n688), .B2(new_n691), .ZN(new_n692));
  NAND3_X1  g0492(.A1(new_n686), .A2(KEYINPUT31), .A3(new_n692), .ZN(new_n693));
  OR2_X1    g0493(.A1(new_n692), .A2(KEYINPUT31), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  OAI211_X1 g0495(.A(new_n682), .B(new_n684), .C1(new_n685), .C2(new_n695), .ZN(new_n696));
  INV_X1    g0496(.A(new_n696), .ZN(new_n697));
  OAI21_X1  g0497(.A(new_n676), .B1(new_n697), .B2(G1), .ZN(G364));
  INV_X1    g0498(.A(new_n647), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n637), .A2(G45), .ZN(new_n700));
  NAND3_X1  g0500(.A1(new_n671), .A2(new_n700), .A3(G1), .ZN(new_n701));
  INV_X1    g0501(.A(new_n701), .ZN(new_n702));
  NOR2_X1   g0502(.A1(new_n699), .A2(new_n702), .ZN(new_n703));
  OAI21_X1  g0503(.A(new_n703), .B1(G330), .B2(new_n646), .ZN(new_n704));
  AOI21_X1  g0504(.A(new_n219), .B1(G20), .B2(new_n288), .ZN(new_n705));
  XNOR2_X1  g0505(.A(new_n705), .B(KEYINPUT97), .ZN(new_n706));
  NAND2_X1  g0506(.A1(new_n293), .A2(G200), .ZN(new_n707));
  XNOR2_X1  g0507(.A(new_n707), .B(KEYINPUT98), .ZN(new_n708));
  NAND3_X1  g0508(.A1(new_n708), .A2(G20), .A3(G190), .ZN(new_n709));
  OAI21_X1  g0509(.A(new_n263), .B1(new_n709), .B2(new_n590), .ZN(new_n710));
  NOR2_X1   g0510(.A1(new_n224), .A2(new_n293), .ZN(new_n711));
  NOR2_X1   g0511(.A1(G190), .A2(G200), .ZN(new_n712));
  AND2_X1   g0512(.A1(new_n711), .A2(new_n712), .ZN(new_n713));
  NOR2_X1   g0513(.A1(G179), .A2(G200), .ZN(new_n714));
  NAND3_X1  g0514(.A1(new_n388), .A2(new_n603), .A3(new_n714), .ZN(new_n715));
  INV_X1    g0515(.A(new_n715), .ZN(new_n716));
  AOI22_X1  g0516(.A1(new_n713), .A2(G311), .B1(G329), .B2(new_n716), .ZN(new_n717));
  INV_X1    g0517(.A(G283), .ZN(new_n718));
  NAND3_X1  g0518(.A1(new_n708), .A2(new_n603), .A3(new_n388), .ZN(new_n719));
  OAI21_X1  g0519(.A(new_n717), .B1(new_n718), .B2(new_n719), .ZN(new_n720));
  NAND2_X1  g0520(.A1(new_n711), .A2(G200), .ZN(new_n721));
  NOR2_X1   g0521(.A1(new_n721), .A2(new_n603), .ZN(new_n722));
  AOI211_X1 g0522(.A(new_n710), .B(new_n720), .C1(G326), .C2(new_n722), .ZN(new_n723));
  INV_X1    g0523(.A(G322), .ZN(new_n724));
  NAND3_X1  g0524(.A1(new_n711), .A2(G190), .A3(new_n346), .ZN(new_n725));
  NAND3_X1  g0525(.A1(new_n711), .A2(new_n603), .A3(G200), .ZN(new_n726));
  XOR2_X1   g0526(.A(KEYINPUT33), .B(G317), .Z(new_n727));
  OAI22_X1  g0527(.A1(new_n724), .A2(new_n725), .B1(new_n726), .B2(new_n727), .ZN(new_n728));
  XOR2_X1   g0528(.A(new_n728), .B(KEYINPUT100), .Z(new_n729));
  AOI21_X1  g0529(.A(new_n224), .B1(G190), .B2(new_n714), .ZN(new_n730));
  OAI211_X1 g0530(.A(new_n723), .B(new_n729), .C1(new_n517), .C2(new_n730), .ZN(new_n731));
  INV_X1    g0531(.A(new_n722), .ZN(new_n732));
  NOR2_X1   g0532(.A1(new_n732), .A2(new_n207), .ZN(new_n733));
  XOR2_X1   g0533(.A(new_n730), .B(KEYINPUT99), .Z(new_n734));
  NOR2_X1   g0534(.A1(new_n734), .A2(new_n448), .ZN(new_n735));
  INV_X1    g0535(.A(new_n726), .ZN(new_n736));
  AOI211_X1 g0536(.A(new_n733), .B(new_n735), .C1(G68), .C2(new_n736), .ZN(new_n737));
  NAND2_X1  g0537(.A1(new_n716), .A2(G159), .ZN(new_n738));
  AOI21_X1  g0538(.A(new_n263), .B1(new_n738), .B2(KEYINPUT32), .ZN(new_n739));
  NOR2_X1   g0539(.A1(new_n719), .A2(new_n233), .ZN(new_n740));
  INV_X1    g0540(.A(new_n713), .ZN(new_n741));
  OAI22_X1  g0541(.A1(new_n741), .A2(new_n211), .B1(new_n542), .B2(new_n709), .ZN(new_n742));
  INV_X1    g0542(.A(new_n725), .ZN(new_n743));
  AOI211_X1 g0543(.A(new_n740), .B(new_n742), .C1(G58), .C2(new_n743), .ZN(new_n744));
  NAND3_X1  g0544(.A1(new_n737), .A2(new_n739), .A3(new_n744), .ZN(new_n745));
  NOR2_X1   g0545(.A1(new_n738), .A2(KEYINPUT32), .ZN(new_n746));
  OAI21_X1  g0546(.A(new_n731), .B1(new_n745), .B2(new_n746), .ZN(new_n747));
  NAND3_X1  g0547(.A1(new_n317), .A2(G355), .A3(new_n227), .ZN(new_n748));
  AND2_X1   g0548(.A1(new_n255), .A2(G45), .ZN(new_n749));
  NOR2_X1   g0549(.A1(new_n381), .A2(new_n383), .ZN(new_n750));
  NOR2_X1   g0550(.A1(new_n750), .A2(new_n669), .ZN(new_n751));
  OAI21_X1  g0551(.A(new_n751), .B1(new_n218), .B2(G45), .ZN(new_n752));
  OAI221_X1 g0552(.A(new_n748), .B1(G116), .B2(new_n227), .C1(new_n749), .C2(new_n752), .ZN(new_n753));
  NOR2_X1   g0553(.A1(G13), .A2(G33), .ZN(new_n754));
  INV_X1    g0554(.A(new_n754), .ZN(new_n755));
  NOR2_X1   g0555(.A1(new_n755), .A2(G20), .ZN(new_n756));
  NOR2_X1   g0556(.A1(new_n706), .A2(new_n756), .ZN(new_n757));
  AOI22_X1  g0557(.A1(new_n706), .A2(new_n747), .B1(new_n753), .B2(new_n757), .ZN(new_n758));
  INV_X1    g0558(.A(new_n756), .ZN(new_n759));
  OAI21_X1  g0559(.A(new_n758), .B1(new_n646), .B2(new_n759), .ZN(new_n760));
  OAI21_X1  g0560(.A(new_n704), .B1(new_n701), .B2(new_n760), .ZN(G396));
  NAND2_X1  g0561(.A1(new_n634), .A2(new_n658), .ZN(new_n762));
  INV_X1    g0562(.A(KEYINPUT104), .ZN(new_n763));
  NAND2_X1  g0563(.A1(new_n343), .A2(new_n763), .ZN(new_n764));
  NAND2_X1  g0564(.A1(new_n643), .A2(new_n335), .ZN(new_n765));
  NAND2_X1  g0565(.A1(new_n764), .A2(new_n765), .ZN(new_n766));
  NAND2_X1  g0566(.A1(new_n343), .A2(new_n348), .ZN(new_n767));
  NAND4_X1  g0567(.A1(new_n343), .A2(new_n763), .A3(new_n335), .A4(new_n643), .ZN(new_n768));
  NAND3_X1  g0568(.A1(new_n766), .A2(new_n767), .A3(new_n768), .ZN(new_n769));
  NAND2_X1  g0569(.A1(new_n769), .A2(KEYINPUT105), .ZN(new_n770));
  INV_X1    g0570(.A(KEYINPUT105), .ZN(new_n771));
  NAND4_X1  g0571(.A1(new_n766), .A2(new_n771), .A3(new_n767), .A4(new_n768), .ZN(new_n772));
  NAND2_X1  g0572(.A1(new_n770), .A2(new_n772), .ZN(new_n773));
  XNOR2_X1  g0573(.A(new_n762), .B(new_n773), .ZN(new_n774));
  NOR2_X1   g0574(.A1(new_n695), .A2(new_n685), .ZN(new_n775));
  NAND2_X1  g0575(.A1(new_n774), .A2(new_n775), .ZN(new_n776));
  XNOR2_X1  g0576(.A(new_n776), .B(KEYINPUT106), .ZN(new_n777));
  NAND2_X1  g0577(.A1(new_n777), .A2(new_n701), .ZN(new_n778));
  INV_X1    g0578(.A(KEYINPUT107), .ZN(new_n779));
  NAND2_X1  g0579(.A1(new_n778), .A2(new_n779), .ZN(new_n780));
  OR2_X1    g0580(.A1(new_n774), .A2(new_n775), .ZN(new_n781));
  NAND3_X1  g0581(.A1(new_n777), .A2(KEYINPUT107), .A3(new_n701), .ZN(new_n782));
  NAND3_X1  g0582(.A1(new_n780), .A2(new_n781), .A3(new_n782), .ZN(new_n783));
  INV_X1    g0583(.A(G137), .ZN(new_n784));
  INV_X1    g0584(.A(G150), .ZN(new_n785));
  OAI22_X1  g0585(.A1(new_n732), .A2(new_n784), .B1(new_n785), .B2(new_n726), .ZN(new_n786));
  XNOR2_X1  g0586(.A(new_n786), .B(KEYINPUT102), .ZN(new_n787));
  INV_X1    g0587(.A(G143), .ZN(new_n788));
  INV_X1    g0588(.A(G159), .ZN(new_n789));
  OAI221_X1 g0589(.A(new_n787), .B1(new_n788), .B2(new_n725), .C1(new_n789), .C2(new_n741), .ZN(new_n790));
  XOR2_X1   g0590(.A(new_n790), .B(KEYINPUT103), .Z(new_n791));
  XNOR2_X1  g0591(.A(new_n791), .B(KEYINPUT34), .ZN(new_n792));
  INV_X1    g0592(.A(new_n750), .ZN(new_n793));
  INV_X1    g0593(.A(new_n719), .ZN(new_n794));
  NAND2_X1  g0594(.A1(new_n794), .A2(G68), .ZN(new_n795));
  OAI21_X1  g0595(.A(new_n795), .B1(new_n207), .B2(new_n709), .ZN(new_n796));
  AOI211_X1 g0596(.A(new_n793), .B(new_n796), .C1(G132), .C2(new_n716), .ZN(new_n797));
  OAI211_X1 g0597(.A(new_n792), .B(new_n797), .C1(new_n201), .C2(new_n730), .ZN(new_n798));
  NOR2_X1   g0598(.A1(new_n719), .A2(new_n542), .ZN(new_n799));
  XNOR2_X1  g0599(.A(KEYINPUT101), .B(G283), .ZN(new_n800));
  OAI22_X1  g0600(.A1(new_n732), .A2(new_n590), .B1(new_n726), .B2(new_n800), .ZN(new_n801));
  NOR2_X1   g0601(.A1(new_n735), .A2(new_n801), .ZN(new_n802));
  OAI22_X1  g0602(.A1(new_n741), .A2(new_n577), .B1(new_n233), .B2(new_n709), .ZN(new_n803));
  AOI21_X1  g0603(.A(new_n803), .B1(G294), .B2(new_n743), .ZN(new_n804));
  AOI21_X1  g0604(.A(new_n317), .B1(new_n716), .B2(G311), .ZN(new_n805));
  NAND3_X1  g0605(.A1(new_n802), .A2(new_n804), .A3(new_n805), .ZN(new_n806));
  OAI21_X1  g0606(.A(new_n798), .B1(new_n799), .B2(new_n806), .ZN(new_n807));
  NOR2_X1   g0607(.A1(new_n706), .A2(new_n754), .ZN(new_n808));
  AOI22_X1  g0608(.A1(new_n807), .A2(new_n706), .B1(new_n211), .B2(new_n808), .ZN(new_n809));
  OAI211_X1 g0609(.A(new_n809), .B(new_n702), .C1(new_n755), .C2(new_n773), .ZN(new_n810));
  NAND2_X1  g0610(.A1(new_n783), .A2(new_n810), .ZN(G384));
  INV_X1    g0611(.A(new_n684), .ZN(new_n812));
  AOI21_X1  g0612(.A(new_n683), .B1(new_n680), .B2(new_n658), .ZN(new_n813));
  OAI21_X1  g0613(.A(new_n444), .B1(new_n812), .B2(new_n813), .ZN(new_n814));
  NAND2_X1  g0614(.A1(new_n619), .A2(new_n814), .ZN(new_n815));
  XNOR2_X1  g0615(.A(new_n815), .B(KEYINPUT111), .ZN(new_n816));
  OR2_X1    g0616(.A1(new_n429), .A2(KEYINPUT16), .ZN(new_n817));
  AOI21_X1  g0617(.A(new_n411), .B1(new_n817), .B2(new_n430), .ZN(new_n818));
  OAI21_X1  g0618(.A(new_n439), .B1(new_n818), .B2(new_n641), .ZN(new_n819));
  NOR2_X1   g0619(.A1(new_n818), .A2(new_n421), .ZN(new_n820));
  OAI21_X1  g0620(.A(KEYINPUT37), .B1(new_n819), .B2(new_n820), .ZN(new_n821));
  INV_X1    g0621(.A(new_n439), .ZN(new_n822));
  AOI22_X1  g0622(.A1(new_n409), .A2(new_n412), .B1(new_n421), .B2(new_n641), .ZN(new_n823));
  OR2_X1    g0623(.A1(new_n822), .A2(new_n823), .ZN(new_n824));
  OAI21_X1  g0624(.A(new_n821), .B1(KEYINPUT37), .B2(new_n824), .ZN(new_n825));
  NAND2_X1  g0625(.A1(new_n402), .A2(new_n300), .ZN(new_n826));
  NOR2_X1   g0626(.A1(new_n429), .A2(KEYINPUT16), .ZN(new_n827));
  OAI21_X1  g0627(.A(new_n412), .B1(new_n826), .B2(new_n827), .ZN(new_n828));
  INV_X1    g0628(.A(new_n641), .ZN(new_n829));
  NAND2_X1  g0629(.A1(new_n828), .A2(new_n829), .ZN(new_n830));
  OAI211_X1 g0630(.A(KEYINPUT38), .B(new_n825), .C1(new_n442), .C2(new_n830), .ZN(new_n831));
  INV_X1    g0631(.A(KEYINPUT108), .ZN(new_n832));
  NAND2_X1  g0632(.A1(new_n831), .A2(new_n832), .ZN(new_n833));
  OAI21_X1  g0633(.A(new_n615), .B1(new_n612), .B2(new_n613), .ZN(new_n834));
  INV_X1    g0634(.A(new_n830), .ZN(new_n835));
  NAND2_X1  g0635(.A1(new_n834), .A2(new_n835), .ZN(new_n836));
  NAND4_X1  g0636(.A1(new_n836), .A2(KEYINPUT108), .A3(KEYINPUT38), .A4(new_n825), .ZN(new_n837));
  NAND2_X1  g0637(.A1(new_n833), .A2(new_n837), .ZN(new_n838));
  NAND2_X1  g0638(.A1(new_n836), .A2(new_n825), .ZN(new_n839));
  INV_X1    g0639(.A(KEYINPUT38), .ZN(new_n840));
  AOI21_X1  g0640(.A(KEYINPUT109), .B1(new_n839), .B2(new_n840), .ZN(new_n841));
  NOR3_X1   g0641(.A1(new_n822), .A2(new_n823), .A3(KEYINPUT37), .ZN(new_n842));
  NAND2_X1  g0642(.A1(new_n828), .A2(new_n422), .ZN(new_n843));
  NAND3_X1  g0643(.A1(new_n830), .A2(new_n843), .A3(new_n439), .ZN(new_n844));
  AOI21_X1  g0644(.A(new_n842), .B1(KEYINPUT37), .B2(new_n844), .ZN(new_n845));
  AOI21_X1  g0645(.A(new_n845), .B1(new_n834), .B2(new_n835), .ZN(new_n846));
  INV_X1    g0646(.A(KEYINPUT109), .ZN(new_n847));
  NOR3_X1   g0647(.A1(new_n846), .A2(new_n847), .A3(KEYINPUT38), .ZN(new_n848));
  OAI21_X1  g0648(.A(new_n838), .B1(new_n841), .B2(new_n848), .ZN(new_n849));
  NAND2_X1  g0649(.A1(new_n311), .A2(new_n643), .ZN(new_n850));
  NAND3_X1  g0650(.A1(new_n312), .A2(new_n352), .A3(new_n850), .ZN(new_n851));
  OAI211_X1 g0651(.A(new_n311), .B(new_n643), .C1(new_n610), .C2(new_n294), .ZN(new_n852));
  AND2_X1   g0652(.A1(new_n851), .A2(new_n852), .ZN(new_n853));
  NAND3_X1  g0653(.A1(new_n773), .A2(new_n634), .A3(new_n658), .ZN(new_n854));
  NAND2_X1  g0654(.A1(new_n344), .A2(new_n658), .ZN(new_n855));
  AOI21_X1  g0655(.A(new_n853), .B1(new_n854), .B2(new_n855), .ZN(new_n856));
  AOI22_X1  g0656(.A1(new_n849), .A2(new_n856), .B1(new_n426), .B2(new_n641), .ZN(new_n857));
  NOR2_X1   g0657(.A1(new_n431), .A2(new_n641), .ZN(new_n858));
  INV_X1    g0658(.A(new_n858), .ZN(new_n859));
  NAND2_X1  g0659(.A1(new_n440), .A2(new_n436), .ZN(new_n860));
  AOI21_X1  g0660(.A(new_n426), .B1(KEYINPUT110), .B2(new_n860), .ZN(new_n861));
  OR2_X1    g0661(.A1(new_n860), .A2(KEYINPUT110), .ZN(new_n862));
  AOI21_X1  g0662(.A(new_n859), .B1(new_n861), .B2(new_n862), .ZN(new_n863));
  AND2_X1   g0663(.A1(new_n824), .A2(KEYINPUT37), .ZN(new_n864));
  NOR2_X1   g0664(.A1(new_n864), .A2(new_n842), .ZN(new_n865));
  OAI21_X1  g0665(.A(new_n840), .B1(new_n863), .B2(new_n865), .ZN(new_n866));
  INV_X1    g0666(.A(KEYINPUT39), .ZN(new_n867));
  AND3_X1   g0667(.A1(new_n866), .A2(new_n867), .A3(new_n831), .ZN(new_n868));
  AOI21_X1  g0668(.A(new_n868), .B1(new_n849), .B2(KEYINPUT39), .ZN(new_n869));
  NAND3_X1  g0669(.A1(new_n294), .A2(new_n311), .A3(new_n658), .ZN(new_n870));
  OAI21_X1  g0670(.A(new_n857), .B1(new_n869), .B2(new_n870), .ZN(new_n871));
  XOR2_X1   g0671(.A(new_n816), .B(new_n871), .Z(new_n872));
  INV_X1    g0672(.A(KEYINPUT40), .ZN(new_n873));
  OAI21_X1  g0673(.A(new_n847), .B1(new_n846), .B2(KEYINPUT38), .ZN(new_n874));
  NOR2_X1   g0674(.A1(new_n442), .A2(new_n830), .ZN(new_n875));
  OAI211_X1 g0675(.A(KEYINPUT109), .B(new_n840), .C1(new_n875), .C2(new_n845), .ZN(new_n876));
  AOI22_X1  g0676(.A1(new_n874), .A2(new_n876), .B1(new_n833), .B2(new_n837), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n851), .A2(new_n852), .ZN(new_n878));
  NAND4_X1  g0678(.A1(new_n693), .A2(new_n694), .A3(new_n773), .A4(new_n878), .ZN(new_n879));
  OAI21_X1  g0679(.A(new_n873), .B1(new_n877), .B2(new_n879), .ZN(new_n880));
  INV_X1    g0680(.A(new_n879), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n866), .A2(new_n831), .ZN(new_n882));
  NAND3_X1  g0682(.A1(new_n881), .A2(KEYINPUT40), .A3(new_n882), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n880), .A2(new_n883), .ZN(new_n884));
  NOR3_X1   g0684(.A1(new_n695), .A2(new_n443), .A3(new_n368), .ZN(new_n885));
  XNOR2_X1  g0685(.A(new_n884), .B(new_n885), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n886), .A2(G330), .ZN(new_n887));
  XNOR2_X1  g0687(.A(new_n872), .B(new_n887), .ZN(new_n888));
  OAI21_X1  g0688(.A(new_n888), .B1(new_n276), .B2(new_n637), .ZN(new_n889));
  AOI21_X1  g0689(.A(new_n577), .B1(new_n452), .B2(KEYINPUT35), .ZN(new_n890));
  NOR2_X1   g0690(.A1(new_n224), .A2(new_n219), .ZN(new_n891));
  OAI211_X1 g0691(.A(new_n890), .B(new_n891), .C1(KEYINPUT35), .C2(new_n452), .ZN(new_n892));
  XNOR2_X1  g0692(.A(new_n892), .B(KEYINPUT36), .ZN(new_n893));
  NOR3_X1   g0693(.A1(new_n674), .A2(new_n211), .A3(new_n398), .ZN(new_n894));
  NOR2_X1   g0694(.A1(new_n202), .A2(G50), .ZN(new_n895));
  OAI211_X1 g0695(.A(G1), .B(new_n305), .C1(new_n894), .C2(new_n895), .ZN(new_n896));
  NAND3_X1  g0696(.A1(new_n889), .A2(new_n893), .A3(new_n896), .ZN(G367));
  NAND2_X1  g0697(.A1(new_n665), .A2(new_n666), .ZN(new_n898));
  OAI211_X1 g0698(.A(new_n482), .B(new_n493), .C1(new_n457), .C2(new_n658), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n620), .A2(new_n643), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n899), .A2(new_n900), .ZN(new_n901));
  INV_X1    g0701(.A(new_n901), .ZN(new_n902));
  OAI21_X1  g0702(.A(KEYINPUT42), .B1(new_n898), .B2(new_n902), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n652), .A2(new_n482), .ZN(new_n904));
  AOI21_X1  g0704(.A(new_n643), .B1(new_n904), .B2(new_n493), .ZN(new_n905));
  INV_X1    g0705(.A(new_n905), .ZN(new_n906));
  INV_X1    g0706(.A(new_n666), .ZN(new_n907));
  NOR2_X1   g0707(.A1(new_n660), .A2(new_n907), .ZN(new_n908));
  INV_X1    g0708(.A(KEYINPUT42), .ZN(new_n909));
  NAND3_X1  g0709(.A1(new_n908), .A2(new_n909), .A3(new_n901), .ZN(new_n910));
  NAND3_X1  g0710(.A1(new_n903), .A2(new_n906), .A3(new_n910), .ZN(new_n911));
  NOR2_X1   g0711(.A1(new_n573), .A2(new_n658), .ZN(new_n912));
  NAND3_X1  g0712(.A1(new_n629), .A2(new_n630), .A3(new_n912), .ZN(new_n913));
  OAI21_X1  g0713(.A(new_n913), .B1(new_n678), .B2(new_n912), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n914), .A2(KEYINPUT43), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n911), .A2(new_n915), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n661), .A2(new_n901), .ZN(new_n917));
  INV_X1    g0717(.A(new_n917), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n916), .A2(new_n918), .ZN(new_n919));
  NOR2_X1   g0719(.A1(new_n914), .A2(KEYINPUT43), .ZN(new_n920));
  NAND3_X1  g0720(.A1(new_n911), .A2(new_n917), .A3(new_n915), .ZN(new_n921));
  AND3_X1   g0721(.A1(new_n919), .A2(new_n920), .A3(new_n921), .ZN(new_n922));
  AOI21_X1  g0722(.A(new_n920), .B1(new_n919), .B2(new_n921), .ZN(new_n923));
  NOR2_X1   g0723(.A1(new_n922), .A2(new_n923), .ZN(new_n924));
  XNOR2_X1  g0724(.A(new_n670), .B(KEYINPUT41), .ZN(new_n925));
  INV_X1    g0725(.A(new_n925), .ZN(new_n926));
  NAND2_X1  g0726(.A1(new_n652), .A2(new_n658), .ZN(new_n927));
  OAI21_X1  g0727(.A(new_n927), .B1(new_n660), .B2(new_n907), .ZN(new_n928));
  AND3_X1   g0728(.A1(new_n928), .A2(KEYINPUT44), .A3(new_n902), .ZN(new_n929));
  AOI21_X1  g0729(.A(KEYINPUT44), .B1(new_n928), .B2(new_n902), .ZN(new_n930));
  NOR2_X1   g0730(.A1(new_n929), .A2(new_n930), .ZN(new_n931));
  OAI211_X1 g0731(.A(new_n927), .B(new_n901), .C1(new_n660), .C2(new_n907), .ZN(new_n932));
  XNOR2_X1  g0732(.A(new_n932), .B(KEYINPUT45), .ZN(new_n933));
  OAI211_X1 g0733(.A(KEYINPUT112), .B(new_n661), .C1(new_n931), .C2(new_n933), .ZN(new_n934));
  NOR2_X1   g0734(.A1(new_n665), .A2(new_n666), .ZN(new_n935));
  OAI21_X1  g0735(.A(new_n647), .B1(new_n935), .B2(new_n908), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n660), .A2(new_n907), .ZN(new_n937));
  NAND3_X1  g0737(.A1(new_n699), .A2(new_n898), .A3(new_n937), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n936), .A2(new_n938), .ZN(new_n939));
  NOR2_X1   g0739(.A1(new_n661), .A2(KEYINPUT112), .ZN(new_n940));
  NOR3_X1   g0740(.A1(new_n696), .A2(new_n939), .A3(new_n940), .ZN(new_n941));
  INV_X1    g0741(.A(KEYINPUT44), .ZN(new_n942));
  OAI21_X1  g0742(.A(new_n942), .B1(new_n667), .B2(new_n901), .ZN(new_n943));
  NAND3_X1  g0743(.A1(new_n928), .A2(KEYINPUT44), .A3(new_n902), .ZN(new_n944));
  NAND4_X1  g0744(.A1(new_n898), .A2(KEYINPUT45), .A3(new_n927), .A4(new_n901), .ZN(new_n945));
  INV_X1    g0745(.A(KEYINPUT45), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n932), .A2(new_n946), .ZN(new_n947));
  AOI22_X1  g0747(.A1(new_n943), .A2(new_n944), .B1(new_n945), .B2(new_n947), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n948), .A2(new_n662), .ZN(new_n949));
  NAND3_X1  g0749(.A1(new_n934), .A2(new_n941), .A3(new_n949), .ZN(new_n950));
  AOI21_X1  g0750(.A(new_n926), .B1(new_n950), .B2(new_n697), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n700), .A2(G1), .ZN(new_n952));
  OAI21_X1  g0752(.A(new_n924), .B1(new_n951), .B2(new_n952), .ZN(new_n953));
  NOR2_X1   g0753(.A1(new_n719), .A2(new_n211), .ZN(new_n954));
  AOI21_X1  g0754(.A(new_n954), .B1(G50), .B2(new_n713), .ZN(new_n955));
  OAI21_X1  g0755(.A(new_n955), .B1(new_n201), .B2(new_n709), .ZN(new_n956));
  AOI21_X1  g0756(.A(new_n956), .B1(G150), .B2(new_n743), .ZN(new_n957));
  OAI22_X1  g0757(.A1(new_n732), .A2(new_n788), .B1(new_n789), .B2(new_n726), .ZN(new_n958));
  AOI211_X1 g0758(.A(new_n263), .B(new_n958), .C1(G137), .C2(new_n716), .ZN(new_n959));
  INV_X1    g0759(.A(new_n734), .ZN(new_n960));
  NAND2_X1  g0760(.A1(new_n960), .A2(G68), .ZN(new_n961));
  NAND3_X1  g0761(.A1(new_n957), .A2(new_n959), .A3(new_n961), .ZN(new_n962));
  NOR2_X1   g0762(.A1(new_n725), .A2(new_n590), .ZN(new_n963));
  NOR2_X1   g0763(.A1(new_n719), .A2(new_n448), .ZN(new_n964));
  OAI221_X1 g0764(.A(new_n793), .B1(new_n730), .B2(new_n233), .C1(new_n726), .C2(new_n517), .ZN(new_n965));
  AOI211_X1 g0765(.A(new_n964), .B(new_n965), .C1(G311), .C2(new_n722), .ZN(new_n966));
  INV_X1    g0766(.A(G317), .ZN(new_n967));
  OAI22_X1  g0767(.A1(new_n741), .A2(new_n800), .B1(new_n967), .B2(new_n715), .ZN(new_n968));
  INV_X1    g0768(.A(KEYINPUT113), .ZN(new_n969));
  OAI21_X1  g0769(.A(new_n969), .B1(new_n709), .B2(new_n577), .ZN(new_n970));
  AOI21_X1  g0770(.A(new_n968), .B1(KEYINPUT46), .B2(new_n970), .ZN(new_n971));
  OAI211_X1 g0771(.A(new_n966), .B(new_n971), .C1(KEYINPUT46), .C2(new_n970), .ZN(new_n972));
  OAI21_X1  g0772(.A(new_n962), .B1(new_n963), .B2(new_n972), .ZN(new_n973));
  XNOR2_X1  g0773(.A(new_n973), .B(KEYINPUT47), .ZN(new_n974));
  AOI21_X1  g0774(.A(new_n701), .B1(new_n974), .B2(new_n706), .ZN(new_n975));
  INV_X1    g0775(.A(new_n751), .ZN(new_n976));
  OAI221_X1 g0776(.A(new_n757), .B1(new_n227), .B2(new_n330), .C1(new_n250), .C2(new_n976), .ZN(new_n977));
  OAI211_X1 g0777(.A(new_n975), .B(new_n977), .C1(new_n759), .C2(new_n914), .ZN(new_n978));
  NAND2_X1  g0778(.A1(new_n953), .A2(new_n978), .ZN(G387));
  INV_X1    g0779(.A(new_n939), .ZN(new_n980));
  NAND2_X1  g0780(.A1(new_n980), .A2(new_n952), .ZN(new_n981));
  AOI22_X1  g0781(.A1(new_n722), .A2(G322), .B1(G303), .B2(new_n713), .ZN(new_n982));
  INV_X1    g0782(.A(G311), .ZN(new_n983));
  OAI221_X1 g0783(.A(new_n982), .B1(new_n983), .B2(new_n726), .C1(new_n967), .C2(new_n725), .ZN(new_n984));
  XNOR2_X1  g0784(.A(new_n984), .B(KEYINPUT48), .ZN(new_n985));
  OAI221_X1 g0785(.A(new_n985), .B1(new_n517), .B2(new_n709), .C1(new_n730), .C2(new_n800), .ZN(new_n986));
  XNOR2_X1  g0786(.A(new_n986), .B(KEYINPUT49), .ZN(new_n987));
  AOI21_X1  g0787(.A(new_n750), .B1(G326), .B2(new_n716), .ZN(new_n988));
  OAI211_X1 g0788(.A(new_n987), .B(new_n988), .C1(new_n577), .C2(new_n719), .ZN(new_n989));
  OAI22_X1  g0789(.A1(new_n732), .A2(new_n789), .B1(new_n207), .B2(new_n725), .ZN(new_n990));
  NOR2_X1   g0790(.A1(new_n734), .A2(new_n330), .ZN(new_n991));
  INV_X1    g0791(.A(new_n991), .ZN(new_n992));
  OAI21_X1  g0792(.A(new_n992), .B1(new_n354), .B2(new_n726), .ZN(new_n993));
  INV_X1    g0793(.A(KEYINPUT115), .ZN(new_n994));
  NOR2_X1   g0794(.A1(new_n964), .A2(new_n793), .ZN(new_n995));
  INV_X1    g0795(.A(new_n709), .ZN(new_n996));
  NAND2_X1  g0796(.A1(new_n996), .A2(G77), .ZN(new_n997));
  OAI211_X1 g0797(.A(new_n995), .B(new_n997), .C1(new_n785), .C2(new_n715), .ZN(new_n998));
  AOI211_X1 g0798(.A(new_n990), .B(new_n993), .C1(new_n994), .C2(new_n998), .ZN(new_n999));
  OAI221_X1 g0799(.A(new_n999), .B1(new_n994), .B2(new_n998), .C1(new_n202), .C2(new_n741), .ZN(new_n1000));
  NAND2_X1  g0800(.A1(new_n989), .A2(new_n1000), .ZN(new_n1001));
  NOR2_X1   g0801(.A1(new_n247), .A2(new_n459), .ZN(new_n1002));
  INV_X1    g0802(.A(new_n1002), .ZN(new_n1003));
  OR2_X1    g0803(.A1(new_n1003), .A2(KEYINPUT114), .ZN(new_n1004));
  NAND2_X1  g0804(.A1(new_n1003), .A2(KEYINPUT114), .ZN(new_n1005));
  OR3_X1    g0805(.A1(new_n354), .A2(KEYINPUT50), .A3(G50), .ZN(new_n1006));
  AOI211_X1 g0806(.A(G116), .B(new_n543), .C1(G68), .C2(G77), .ZN(new_n1007));
  OAI21_X1  g0807(.A(KEYINPUT50), .B1(new_n354), .B2(G50), .ZN(new_n1008));
  NAND4_X1  g0808(.A1(new_n1006), .A2(new_n1007), .A3(new_n1008), .A4(new_n459), .ZN(new_n1009));
  NAND4_X1  g0809(.A1(new_n1004), .A2(new_n1005), .A3(new_n751), .A4(new_n1009), .ZN(new_n1010));
  NAND2_X1  g0810(.A1(new_n317), .A2(new_n227), .ZN(new_n1011));
  OAI221_X1 g0811(.A(new_n1010), .B1(G107), .B2(new_n227), .C1(new_n672), .C2(new_n1011), .ZN(new_n1012));
  AOI22_X1  g0812(.A1(new_n1001), .A2(new_n706), .B1(new_n757), .B2(new_n1012), .ZN(new_n1013));
  OAI211_X1 g0813(.A(new_n1013), .B(new_n702), .C1(new_n665), .C2(new_n759), .ZN(new_n1014));
  NAND2_X1  g0814(.A1(new_n697), .A2(new_n980), .ZN(new_n1015));
  INV_X1    g0815(.A(new_n1015), .ZN(new_n1016));
  OAI21_X1  g0816(.A(new_n670), .B1(new_n697), .B2(new_n980), .ZN(new_n1017));
  OAI211_X1 g0817(.A(new_n981), .B(new_n1014), .C1(new_n1016), .C2(new_n1017), .ZN(G393));
  OAI21_X1  g0818(.A(KEYINPUT116), .B1(new_n948), .B2(new_n662), .ZN(new_n1019));
  INV_X1    g0819(.A(KEYINPUT116), .ZN(new_n1020));
  OAI211_X1 g0820(.A(new_n1020), .B(new_n661), .C1(new_n931), .C2(new_n933), .ZN(new_n1021));
  NAND4_X1  g0821(.A1(new_n1019), .A2(new_n1021), .A3(new_n952), .A4(new_n949), .ZN(new_n1022));
  OAI22_X1  g0822(.A1(new_n732), .A2(new_n967), .B1(new_n983), .B2(new_n725), .ZN(new_n1023));
  XNOR2_X1  g0823(.A(new_n1023), .B(KEYINPUT52), .ZN(new_n1024));
  OAI22_X1  g0824(.A1(new_n709), .A2(new_n800), .B1(new_n715), .B2(new_n724), .ZN(new_n1025));
  NOR2_X1   g0825(.A1(new_n726), .A2(new_n590), .ZN(new_n1026));
  OAI21_X1  g0826(.A(new_n263), .B1(new_n730), .B2(new_n577), .ZN(new_n1027));
  NOR4_X1   g0827(.A1(new_n1025), .A2(new_n740), .A3(new_n1026), .A4(new_n1027), .ZN(new_n1028));
  OAI211_X1 g0828(.A(new_n1024), .B(new_n1028), .C1(new_n517), .C2(new_n741), .ZN(new_n1029));
  AOI22_X1  g0829(.A1(new_n996), .A2(G68), .B1(G143), .B2(new_n716), .ZN(new_n1030));
  OAI21_X1  g0830(.A(new_n1030), .B1(new_n354), .B2(new_n741), .ZN(new_n1031));
  AOI211_X1 g0831(.A(new_n799), .B(new_n1031), .C1(G50), .C2(new_n736), .ZN(new_n1032));
  NAND2_X1  g0832(.A1(new_n960), .A2(G77), .ZN(new_n1033));
  OAI22_X1  g0833(.A1(new_n732), .A2(new_n785), .B1(new_n789), .B2(new_n725), .ZN(new_n1034));
  XNOR2_X1  g0834(.A(new_n1034), .B(KEYINPUT51), .ZN(new_n1035));
  NAND3_X1  g0835(.A1(new_n1032), .A2(new_n1033), .A3(new_n1035), .ZN(new_n1036));
  OAI21_X1  g0836(.A(new_n1029), .B1(new_n1036), .B2(new_n793), .ZN(new_n1037));
  AOI21_X1  g0837(.A(new_n701), .B1(new_n1037), .B2(new_n706), .ZN(new_n1038));
  AOI22_X1  g0838(.A1(new_n259), .A2(new_n751), .B1(G97), .B2(new_n669), .ZN(new_n1039));
  NAND2_X1  g0839(.A1(new_n1039), .A2(new_n757), .ZN(new_n1040));
  OAI211_X1 g0840(.A(new_n1038), .B(new_n1040), .C1(new_n759), .C2(new_n901), .ZN(new_n1041));
  AND2_X1   g0841(.A1(new_n1022), .A2(new_n1041), .ZN(new_n1042));
  NAND3_X1  g0842(.A1(new_n1019), .A2(new_n949), .A3(new_n1021), .ZN(new_n1043));
  AND2_X1   g0843(.A1(new_n1043), .A2(new_n1015), .ZN(new_n1044));
  NAND2_X1  g0844(.A1(new_n950), .A2(new_n670), .ZN(new_n1045));
  OAI21_X1  g0845(.A(new_n1042), .B1(new_n1044), .B2(new_n1045), .ZN(G390));
  NAND2_X1  g0846(.A1(new_n854), .A2(new_n855), .ZN(new_n1047));
  NAND4_X1  g0847(.A1(new_n693), .A2(G330), .A3(new_n694), .A4(new_n773), .ZN(new_n1048));
  AND2_X1   g0848(.A1(new_n1048), .A2(new_n853), .ZN(new_n1049));
  NOR2_X1   g0849(.A1(new_n1048), .A2(new_n853), .ZN(new_n1050));
  OAI21_X1  g0850(.A(new_n1047), .B1(new_n1049), .B2(new_n1050), .ZN(new_n1051));
  OR2_X1    g0851(.A1(new_n1048), .A2(new_n853), .ZN(new_n1052));
  NAND3_X1  g0852(.A1(new_n680), .A2(new_n658), .A3(new_n773), .ZN(new_n1053));
  AND2_X1   g0853(.A1(new_n1053), .A2(new_n855), .ZN(new_n1054));
  NAND2_X1  g0854(.A1(new_n1048), .A2(new_n853), .ZN(new_n1055));
  NAND3_X1  g0855(.A1(new_n1052), .A2(new_n1054), .A3(new_n1055), .ZN(new_n1056));
  NAND2_X1  g0856(.A1(new_n1051), .A2(new_n1056), .ZN(new_n1057));
  NAND4_X1  g0857(.A1(new_n444), .A2(new_n693), .A3(G330), .A4(new_n694), .ZN(new_n1058));
  NAND3_X1  g0858(.A1(new_n619), .A2(new_n814), .A3(new_n1058), .ZN(new_n1059));
  INV_X1    g0859(.A(new_n1059), .ZN(new_n1060));
  NAND2_X1  g0860(.A1(new_n1057), .A2(new_n1060), .ZN(new_n1061));
  OAI211_X1 g0861(.A(new_n882), .B(new_n870), .C1(new_n1054), .C2(new_n853), .ZN(new_n1062));
  NAND3_X1  g0862(.A1(new_n866), .A2(new_n867), .A3(new_n831), .ZN(new_n1063));
  OAI21_X1  g0863(.A(new_n1063), .B1(new_n877), .B2(new_n867), .ZN(new_n1064));
  INV_X1    g0864(.A(new_n870), .ZN(new_n1065));
  NOR2_X1   g0865(.A1(new_n856), .A2(new_n1065), .ZN(new_n1066));
  OAI211_X1 g0866(.A(new_n1062), .B(new_n1052), .C1(new_n1064), .C2(new_n1066), .ZN(new_n1067));
  INV_X1    g0867(.A(new_n1067), .ZN(new_n1068));
  OAI221_X1 g0868(.A(new_n1063), .B1(new_n856), .B2(new_n1065), .C1(new_n877), .C2(new_n867), .ZN(new_n1069));
  AOI21_X1  g0869(.A(new_n1052), .B1(new_n1069), .B2(new_n1062), .ZN(new_n1070));
  OAI21_X1  g0870(.A(new_n1061), .B1(new_n1068), .B2(new_n1070), .ZN(new_n1071));
  OAI21_X1  g0871(.A(new_n1062), .B1(new_n1064), .B2(new_n1066), .ZN(new_n1072));
  NAND2_X1  g0872(.A1(new_n1072), .A2(new_n1050), .ZN(new_n1073));
  AOI21_X1  g0873(.A(new_n1059), .B1(new_n1051), .B2(new_n1056), .ZN(new_n1074));
  NAND3_X1  g0874(.A1(new_n1073), .A2(new_n1074), .A3(new_n1067), .ZN(new_n1075));
  NAND3_X1  g0875(.A1(new_n1071), .A2(new_n670), .A3(new_n1075), .ZN(new_n1076));
  NAND2_X1  g0876(.A1(new_n869), .A2(new_n754), .ZN(new_n1077));
  OAI221_X1 g0877(.A(new_n795), .B1(new_n517), .B2(new_n715), .C1(new_n577), .C2(new_n725), .ZN(new_n1078));
  AOI21_X1  g0878(.A(new_n1078), .B1(G97), .B2(new_n713), .ZN(new_n1079));
  OAI22_X1  g0879(.A1(new_n732), .A2(new_n718), .B1(new_n233), .B2(new_n726), .ZN(new_n1080));
  AOI21_X1  g0880(.A(new_n1080), .B1(G87), .B2(new_n996), .ZN(new_n1081));
  NAND4_X1  g0881(.A1(new_n1079), .A2(new_n263), .A3(new_n1033), .A4(new_n1081), .ZN(new_n1082));
  AOI22_X1  g0882(.A1(new_n960), .A2(G159), .B1(new_n736), .B2(G137), .ZN(new_n1083));
  XOR2_X1   g0883(.A(KEYINPUT54), .B(G143), .Z(new_n1084));
  NAND2_X1  g0884(.A1(new_n713), .A2(new_n1084), .ZN(new_n1085));
  AOI21_X1  g0885(.A(new_n263), .B1(new_n722), .B2(G128), .ZN(new_n1086));
  INV_X1    g0886(.A(G125), .ZN(new_n1087));
  OAI22_X1  g0887(.A1(new_n719), .A2(new_n207), .B1(new_n715), .B2(new_n1087), .ZN(new_n1088));
  NAND3_X1  g0888(.A1(new_n996), .A2(KEYINPUT53), .A3(G150), .ZN(new_n1089));
  INV_X1    g0889(.A(KEYINPUT53), .ZN(new_n1090));
  OAI21_X1  g0890(.A(new_n1090), .B1(new_n709), .B2(new_n785), .ZN(new_n1091));
  AOI21_X1  g0891(.A(new_n1088), .B1(new_n1089), .B2(new_n1091), .ZN(new_n1092));
  NAND4_X1  g0892(.A1(new_n1083), .A2(new_n1085), .A3(new_n1086), .A4(new_n1092), .ZN(new_n1093));
  INV_X1    g0893(.A(G132), .ZN(new_n1094));
  NOR2_X1   g0894(.A1(new_n725), .A2(new_n1094), .ZN(new_n1095));
  OAI21_X1  g0895(.A(new_n1082), .B1(new_n1093), .B2(new_n1095), .ZN(new_n1096));
  AOI22_X1  g0896(.A1(new_n1096), .A2(new_n706), .B1(new_n354), .B2(new_n808), .ZN(new_n1097));
  AND3_X1   g0897(.A1(new_n1077), .A2(new_n702), .A3(new_n1097), .ZN(new_n1098));
  NOR2_X1   g0898(.A1(new_n1068), .A2(new_n1070), .ZN(new_n1099));
  AOI21_X1  g0899(.A(new_n1098), .B1(new_n1099), .B2(new_n952), .ZN(new_n1100));
  NAND2_X1  g0900(.A1(new_n1076), .A2(new_n1100), .ZN(new_n1101));
  INV_X1    g0901(.A(KEYINPUT117), .ZN(new_n1102));
  NAND2_X1  g0902(.A1(new_n1101), .A2(new_n1102), .ZN(new_n1103));
  NAND3_X1  g0903(.A1(new_n1076), .A2(new_n1100), .A3(KEYINPUT117), .ZN(new_n1104));
  NAND2_X1  g0904(.A1(new_n1103), .A2(new_n1104), .ZN(G378));
  NAND2_X1  g0905(.A1(new_n1075), .A2(new_n1060), .ZN(new_n1106));
  AND3_X1   g0906(.A1(new_n880), .A2(G330), .A3(new_n883), .ZN(new_n1107));
  NAND2_X1  g0907(.A1(new_n1107), .A2(new_n871), .ZN(new_n1108));
  NOR2_X1   g0908(.A1(new_n369), .A2(new_n641), .ZN(new_n1109));
  INV_X1    g0909(.A(new_n1109), .ZN(new_n1110));
  NAND3_X1  g0910(.A1(new_n618), .A2(new_n367), .A3(new_n1110), .ZN(new_n1111));
  NOR2_X1   g0911(.A1(new_n380), .A2(new_n617), .ZN(new_n1112));
  AOI21_X1  g0912(.A(KEYINPUT94), .B1(new_n376), .B2(new_n379), .ZN(new_n1113));
  OAI21_X1  g0913(.A(new_n367), .B1(new_n1112), .B2(new_n1113), .ZN(new_n1114));
  NAND2_X1  g0914(.A1(new_n1114), .A2(new_n1109), .ZN(new_n1115));
  INV_X1    g0915(.A(KEYINPUT55), .ZN(new_n1116));
  AND3_X1   g0916(.A1(new_n1111), .A2(new_n1115), .A3(new_n1116), .ZN(new_n1117));
  AOI21_X1  g0917(.A(new_n1116), .B1(new_n1111), .B2(new_n1115), .ZN(new_n1118));
  INV_X1    g0918(.A(KEYINPUT56), .ZN(new_n1119));
  NOR3_X1   g0919(.A1(new_n1117), .A2(new_n1118), .A3(new_n1119), .ZN(new_n1120));
  NAND2_X1  g0920(.A1(new_n1111), .A2(new_n1115), .ZN(new_n1121));
  NAND2_X1  g0921(.A1(new_n1121), .A2(KEYINPUT55), .ZN(new_n1122));
  NAND3_X1  g0922(.A1(new_n1111), .A2(new_n1115), .A3(new_n1116), .ZN(new_n1123));
  AOI21_X1  g0923(.A(KEYINPUT56), .B1(new_n1122), .B2(new_n1123), .ZN(new_n1124));
  NOR2_X1   g0924(.A1(new_n1120), .A2(new_n1124), .ZN(new_n1125));
  NAND3_X1  g0925(.A1(new_n880), .A2(G330), .A3(new_n883), .ZN(new_n1126));
  NAND2_X1  g0926(.A1(new_n1064), .A2(new_n1065), .ZN(new_n1127));
  NAND3_X1  g0927(.A1(new_n1126), .A2(new_n1127), .A3(new_n857), .ZN(new_n1128));
  AND3_X1   g0928(.A1(new_n1108), .A2(new_n1125), .A3(new_n1128), .ZN(new_n1129));
  AOI21_X1  g0929(.A(new_n1125), .B1(new_n1108), .B2(new_n1128), .ZN(new_n1130));
  OAI21_X1  g0930(.A(new_n1106), .B1(new_n1129), .B2(new_n1130), .ZN(new_n1131));
  INV_X1    g0931(.A(KEYINPUT57), .ZN(new_n1132));
  NAND2_X1  g0932(.A1(new_n1131), .A2(new_n1132), .ZN(new_n1133));
  OR2_X1    g0933(.A1(new_n1120), .A2(new_n1124), .ZN(new_n1134));
  NOR2_X1   g0934(.A1(new_n1107), .A2(new_n871), .ZN(new_n1135));
  AOI21_X1  g0935(.A(new_n1126), .B1(new_n1127), .B2(new_n857), .ZN(new_n1136));
  OAI21_X1  g0936(.A(new_n1134), .B1(new_n1135), .B2(new_n1136), .ZN(new_n1137));
  NAND3_X1  g0937(.A1(new_n1108), .A2(new_n1125), .A3(new_n1128), .ZN(new_n1138));
  NAND2_X1  g0938(.A1(new_n1137), .A2(new_n1138), .ZN(new_n1139));
  NAND3_X1  g0939(.A1(new_n1139), .A2(KEYINPUT57), .A3(new_n1106), .ZN(new_n1140));
  NAND3_X1  g0940(.A1(new_n1133), .A2(new_n1140), .A3(new_n670), .ZN(new_n1141));
  NAND2_X1  g0941(.A1(new_n1125), .A2(new_n754), .ZN(new_n1142));
  AOI22_X1  g0942(.A1(new_n996), .A2(new_n1084), .B1(new_n743), .B2(G128), .ZN(new_n1143));
  XOR2_X1   g0943(.A(new_n1143), .B(KEYINPUT119), .Z(new_n1144));
  OAI22_X1  g0944(.A1(new_n732), .A2(new_n1087), .B1(new_n741), .B2(new_n784), .ZN(new_n1145));
  AOI21_X1  g0945(.A(new_n1145), .B1(G150), .B2(new_n960), .ZN(new_n1146));
  OAI211_X1 g0946(.A(new_n1144), .B(new_n1146), .C1(new_n1094), .C2(new_n726), .ZN(new_n1147));
  XOR2_X1   g0947(.A(new_n1147), .B(KEYINPUT120), .Z(new_n1148));
  XNOR2_X1  g0948(.A(new_n1148), .B(KEYINPUT59), .ZN(new_n1149));
  AOI21_X1  g0949(.A(G41), .B1(new_n794), .B2(G159), .ZN(new_n1150));
  AOI21_X1  g0950(.A(G33), .B1(new_n716), .B2(G124), .ZN(new_n1151));
  NAND3_X1  g0951(.A1(new_n1149), .A2(new_n1150), .A3(new_n1151), .ZN(new_n1152));
  NAND2_X1  g0952(.A1(new_n750), .A2(G33), .ZN(new_n1153));
  INV_X1    g0953(.A(G41), .ZN(new_n1154));
  AOI21_X1  g0954(.A(G50), .B1(new_n1153), .B2(new_n1154), .ZN(new_n1155));
  INV_X1    g0955(.A(KEYINPUT118), .ZN(new_n1156));
  NAND2_X1  g0956(.A1(new_n1155), .A2(new_n1156), .ZN(new_n1157));
  OAI22_X1  g0957(.A1(new_n741), .A2(new_n330), .B1(new_n233), .B2(new_n725), .ZN(new_n1158));
  AOI21_X1  g0958(.A(new_n1158), .B1(G283), .B2(new_n716), .ZN(new_n1159));
  NAND3_X1  g0959(.A1(new_n997), .A2(new_n1154), .A3(new_n793), .ZN(new_n1160));
  INV_X1    g0960(.A(new_n1160), .ZN(new_n1161));
  AOI22_X1  g0961(.A1(G116), .A2(new_n722), .B1(new_n736), .B2(G97), .ZN(new_n1162));
  NAND4_X1  g0962(.A1(new_n1159), .A2(new_n1161), .A3(new_n961), .A4(new_n1162), .ZN(new_n1163));
  NOR2_X1   g0963(.A1(new_n719), .A2(new_n201), .ZN(new_n1164));
  NOR2_X1   g0964(.A1(new_n1163), .A2(new_n1164), .ZN(new_n1165));
  OAI21_X1  g0965(.A(new_n1157), .B1(new_n1165), .B2(KEYINPUT58), .ZN(new_n1166));
  AOI21_X1  g0966(.A(new_n1166), .B1(KEYINPUT58), .B2(new_n1165), .ZN(new_n1167));
  OAI211_X1 g0967(.A(new_n1152), .B(new_n1167), .C1(new_n1156), .C2(new_n1155), .ZN(new_n1168));
  AOI22_X1  g0968(.A1(new_n1168), .A2(new_n706), .B1(new_n207), .B2(new_n808), .ZN(new_n1169));
  AND3_X1   g0969(.A1(new_n1142), .A2(new_n702), .A3(new_n1169), .ZN(new_n1170));
  AOI21_X1  g0970(.A(new_n1170), .B1(new_n1139), .B2(new_n952), .ZN(new_n1171));
  NAND2_X1  g0971(.A1(new_n1141), .A2(new_n1171), .ZN(new_n1172));
  NAND2_X1  g0972(.A1(new_n1172), .A2(KEYINPUT121), .ZN(new_n1173));
  INV_X1    g0973(.A(KEYINPUT121), .ZN(new_n1174));
  NAND3_X1  g0974(.A1(new_n1141), .A2(new_n1174), .A3(new_n1171), .ZN(new_n1175));
  NAND2_X1  g0975(.A1(new_n1173), .A2(new_n1175), .ZN(G375));
  NAND2_X1  g0976(.A1(new_n853), .A2(new_n754), .ZN(new_n1177));
  OAI22_X1  g0977(.A1(new_n734), .A2(new_n207), .B1(new_n732), .B2(new_n1094), .ZN(new_n1178));
  NOR2_X1   g0978(.A1(new_n1178), .A2(new_n1164), .ZN(new_n1179));
  NAND2_X1  g0979(.A1(new_n713), .A2(G150), .ZN(new_n1180));
  NAND2_X1  g0980(.A1(new_n716), .A2(G128), .ZN(new_n1181));
  OAI21_X1  g0981(.A(new_n1181), .B1(new_n709), .B2(new_n789), .ZN(new_n1182));
  AOI21_X1  g0982(.A(new_n1182), .B1(new_n743), .B2(G137), .ZN(new_n1183));
  AOI21_X1  g0983(.A(new_n793), .B1(new_n736), .B2(new_n1084), .ZN(new_n1184));
  NAND4_X1  g0984(.A1(new_n1179), .A2(new_n1180), .A3(new_n1183), .A4(new_n1184), .ZN(new_n1185));
  AOI22_X1  g0985(.A1(new_n743), .A2(G283), .B1(new_n713), .B2(G107), .ZN(new_n1186));
  OAI21_X1  g0986(.A(new_n1186), .B1(new_n590), .B2(new_n715), .ZN(new_n1187));
  AOI21_X1  g0987(.A(new_n1187), .B1(G97), .B2(new_n996), .ZN(new_n1188));
  NOR2_X1   g0988(.A1(new_n726), .A2(new_n577), .ZN(new_n1189));
  AOI211_X1 g0989(.A(new_n1189), .B(new_n954), .C1(G294), .C2(new_n722), .ZN(new_n1190));
  NAND3_X1  g0990(.A1(new_n1188), .A2(new_n992), .A3(new_n1190), .ZN(new_n1191));
  OAI21_X1  g0991(.A(new_n1185), .B1(new_n1191), .B2(new_n317), .ZN(new_n1192));
  AOI22_X1  g0992(.A1(new_n1192), .A2(new_n706), .B1(new_n202), .B2(new_n808), .ZN(new_n1193));
  AND3_X1   g0993(.A1(new_n1177), .A2(new_n702), .A3(new_n1193), .ZN(new_n1194));
  AOI21_X1  g0994(.A(new_n1194), .B1(new_n1057), .B2(new_n952), .ZN(new_n1195));
  NAND3_X1  g0995(.A1(new_n1051), .A2(new_n1056), .A3(new_n1059), .ZN(new_n1196));
  NAND2_X1  g0996(.A1(new_n1196), .A2(new_n925), .ZN(new_n1197));
  OAI21_X1  g0997(.A(new_n1195), .B1(new_n1197), .B2(new_n1074), .ZN(G381));
  INV_X1    g0998(.A(KEYINPUT123), .ZN(new_n1199));
  NAND2_X1  g0999(.A1(new_n1101), .A2(new_n1199), .ZN(new_n1200));
  NAND3_X1  g1000(.A1(new_n1076), .A2(new_n1100), .A3(KEYINPUT123), .ZN(new_n1201));
  NAND2_X1  g1001(.A1(new_n1200), .A2(new_n1201), .ZN(new_n1202));
  INV_X1    g1002(.A(new_n1202), .ZN(new_n1203));
  NOR2_X1   g1003(.A1(G375), .A2(new_n1203), .ZN(new_n1204));
  NOR2_X1   g1004(.A1(G390), .A2(G381), .ZN(new_n1205));
  AND2_X1   g1005(.A1(new_n783), .A2(new_n810), .ZN(new_n1206));
  NOR2_X1   g1006(.A1(G393), .A2(G396), .ZN(new_n1207));
  NAND2_X1  g1007(.A1(new_n1206), .A2(new_n1207), .ZN(new_n1208));
  XNOR2_X1  g1008(.A(new_n1208), .B(KEYINPUT122), .ZN(new_n1209));
  NOR2_X1   g1009(.A1(new_n1209), .A2(G387), .ZN(new_n1210));
  NAND3_X1  g1010(.A1(new_n1204), .A2(new_n1205), .A3(new_n1210), .ZN(G407));
  INV_X1    g1011(.A(G213), .ZN(new_n1212));
  AOI21_X1  g1012(.A(new_n1212), .B1(new_n1204), .B2(new_n642), .ZN(new_n1213));
  NAND2_X1  g1013(.A1(new_n1213), .A2(G407), .ZN(G409));
  INV_X1    g1014(.A(KEYINPUT126), .ZN(new_n1215));
  NAND2_X1  g1015(.A1(new_n1022), .A2(new_n1041), .ZN(new_n1216));
  INV_X1    g1016(.A(new_n1045), .ZN(new_n1217));
  NAND2_X1  g1017(.A1(new_n1043), .A2(new_n1015), .ZN(new_n1218));
  AOI21_X1  g1018(.A(new_n1216), .B1(new_n1217), .B2(new_n1218), .ZN(new_n1219));
  OAI21_X1  g1019(.A(new_n1215), .B1(G387), .B2(new_n1219), .ZN(new_n1220));
  INV_X1    g1020(.A(new_n1207), .ZN(new_n1221));
  NAND2_X1  g1021(.A1(G393), .A2(G396), .ZN(new_n1222));
  NAND3_X1  g1022(.A1(new_n1220), .A2(new_n1221), .A3(new_n1222), .ZN(new_n1223));
  NAND2_X1  g1023(.A1(G387), .A2(new_n1219), .ZN(new_n1224));
  NAND3_X1  g1024(.A1(G390), .A2(new_n978), .A3(new_n953), .ZN(new_n1225));
  NAND2_X1  g1025(.A1(new_n1224), .A2(new_n1225), .ZN(new_n1226));
  NOR2_X1   g1026(.A1(new_n1223), .A2(new_n1226), .ZN(new_n1227));
  AOI21_X1  g1027(.A(new_n1207), .B1(new_n1225), .B2(new_n1215), .ZN(new_n1228));
  AOI22_X1  g1028(.A1(new_n1228), .A2(new_n1222), .B1(new_n1225), .B2(new_n1224), .ZN(new_n1229));
  NOR2_X1   g1029(.A1(new_n1227), .A2(new_n1229), .ZN(new_n1230));
  INV_X1    g1030(.A(KEYINPUT61), .ZN(new_n1231));
  NOR2_X1   g1031(.A1(new_n1212), .A2(G343), .ZN(new_n1232));
  NAND3_X1  g1032(.A1(new_n1141), .A2(G378), .A3(new_n1171), .ZN(new_n1233));
  OAI211_X1 g1033(.A(new_n925), .B(new_n1106), .C1(new_n1129), .C2(new_n1130), .ZN(new_n1234));
  INV_X1    g1034(.A(KEYINPUT124), .ZN(new_n1235));
  NAND2_X1  g1035(.A1(new_n1234), .A2(new_n1235), .ZN(new_n1236));
  NAND4_X1  g1036(.A1(new_n1139), .A2(KEYINPUT124), .A3(new_n925), .A4(new_n1106), .ZN(new_n1237));
  NAND3_X1  g1037(.A1(new_n1236), .A2(new_n1171), .A3(new_n1237), .ZN(new_n1238));
  NAND2_X1  g1038(.A1(new_n1238), .A2(new_n1202), .ZN(new_n1239));
  AOI21_X1  g1039(.A(new_n1232), .B1(new_n1233), .B2(new_n1239), .ZN(new_n1240));
  INV_X1    g1040(.A(KEYINPUT60), .ZN(new_n1241));
  AOI21_X1  g1041(.A(new_n671), .B1(new_n1196), .B2(new_n1241), .ZN(new_n1242));
  OAI211_X1 g1042(.A(new_n1242), .B(new_n1061), .C1(new_n1241), .C2(new_n1196), .ZN(new_n1243));
  NAND2_X1  g1043(.A1(new_n1243), .A2(new_n1195), .ZN(new_n1244));
  NAND2_X1  g1044(.A1(new_n1206), .A2(new_n1244), .ZN(new_n1245));
  NAND3_X1  g1045(.A1(G384), .A2(new_n1195), .A3(new_n1243), .ZN(new_n1246));
  NAND2_X1  g1046(.A1(new_n1245), .A2(new_n1246), .ZN(new_n1247));
  NAND3_X1  g1047(.A1(new_n1247), .A2(G2897), .A3(new_n1232), .ZN(new_n1248));
  NAND2_X1  g1048(.A1(new_n1232), .A2(G2897), .ZN(new_n1249));
  NAND3_X1  g1049(.A1(new_n1245), .A2(new_n1246), .A3(new_n1249), .ZN(new_n1250));
  NAND2_X1  g1050(.A1(new_n1248), .A2(new_n1250), .ZN(new_n1251));
  OAI211_X1 g1051(.A(new_n1230), .B(new_n1231), .C1(new_n1240), .C2(new_n1251), .ZN(new_n1252));
  INV_X1    g1052(.A(new_n1252), .ZN(new_n1253));
  AOI211_X1 g1053(.A(new_n1232), .B(new_n1247), .C1(new_n1233), .C2(new_n1239), .ZN(new_n1254));
  OAI21_X1  g1054(.A(KEYINPUT125), .B1(new_n1254), .B2(KEYINPUT63), .ZN(new_n1255));
  INV_X1    g1055(.A(new_n1247), .ZN(new_n1256));
  NAND2_X1  g1056(.A1(new_n1240), .A2(new_n1256), .ZN(new_n1257));
  INV_X1    g1057(.A(KEYINPUT125), .ZN(new_n1258));
  INV_X1    g1058(.A(KEYINPUT63), .ZN(new_n1259));
  NAND3_X1  g1059(.A1(new_n1257), .A2(new_n1258), .A3(new_n1259), .ZN(new_n1260));
  NAND2_X1  g1060(.A1(new_n1254), .A2(KEYINPUT63), .ZN(new_n1261));
  NAND4_X1  g1061(.A1(new_n1253), .A2(new_n1255), .A3(new_n1260), .A4(new_n1261), .ZN(new_n1262));
  OR2_X1    g1062(.A1(new_n1227), .A2(new_n1229), .ZN(new_n1263));
  NAND2_X1  g1063(.A1(new_n1233), .A2(new_n1239), .ZN(new_n1264));
  INV_X1    g1064(.A(new_n1232), .ZN(new_n1265));
  XOR2_X1   g1065(.A(KEYINPUT127), .B(KEYINPUT62), .Z(new_n1266));
  NAND4_X1  g1066(.A1(new_n1264), .A2(new_n1265), .A3(new_n1256), .A4(new_n1266), .ZN(new_n1267));
  NAND2_X1  g1067(.A1(KEYINPUT127), .A2(KEYINPUT62), .ZN(new_n1268));
  OAI21_X1  g1068(.A(new_n1267), .B1(new_n1254), .B2(new_n1268), .ZN(new_n1269));
  OAI21_X1  g1069(.A(new_n1231), .B1(new_n1240), .B2(new_n1251), .ZN(new_n1270));
  OAI21_X1  g1070(.A(new_n1263), .B1(new_n1269), .B2(new_n1270), .ZN(new_n1271));
  NAND2_X1  g1071(.A1(new_n1262), .A2(new_n1271), .ZN(G405));
  NAND2_X1  g1072(.A1(G375), .A2(new_n1202), .ZN(new_n1273));
  AOI21_X1  g1073(.A(new_n1263), .B1(new_n1273), .B2(new_n1233), .ZN(new_n1274));
  AOI21_X1  g1074(.A(new_n1203), .B1(new_n1173), .B2(new_n1175), .ZN(new_n1275));
  INV_X1    g1075(.A(new_n1233), .ZN(new_n1276));
  NOR3_X1   g1076(.A1(new_n1275), .A2(new_n1230), .A3(new_n1276), .ZN(new_n1277));
  OAI21_X1  g1077(.A(new_n1247), .B1(new_n1274), .B2(new_n1277), .ZN(new_n1278));
  NAND3_X1  g1078(.A1(new_n1273), .A2(new_n1263), .A3(new_n1233), .ZN(new_n1279));
  OAI21_X1  g1079(.A(new_n1230), .B1(new_n1275), .B2(new_n1276), .ZN(new_n1280));
  NAND3_X1  g1080(.A1(new_n1279), .A2(new_n1280), .A3(new_n1256), .ZN(new_n1281));
  NAND2_X1  g1081(.A1(new_n1278), .A2(new_n1281), .ZN(G402));
endmodule


