//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 1 0 0 0 0 1 0 0 0 0 1 1 1 0 0 1 0 0 0 0 1 1 1 0 0 1 0 1 1 0 1 1 1 1 0 0 0 1 1 0 1 1 0 1 1 1 0 1 1 1 0 1 0 1 0 0 0 0 1 0 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:27:51 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n678,
    new_n679, new_n680, new_n681, new_n682, new_n683, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n692, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n733, new_n734, new_n735, new_n736, new_n737, new_n738,
    new_n739, new_n740, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n752, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n760, new_n761, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n769, new_n770, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n784, new_n785, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n821, new_n822, new_n823, new_n824,
    new_n825, new_n826, new_n827, new_n828, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n915, new_n916, new_n917,
    new_n918, new_n919, new_n920, new_n921, new_n922, new_n923, new_n924,
    new_n925, new_n926, new_n927, new_n928, new_n929, new_n930, new_n931,
    new_n932, new_n933, new_n934, new_n935, new_n936, new_n937, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n949, new_n950, new_n951, new_n952, new_n954, new_n955,
    new_n956, new_n957, new_n958, new_n959, new_n960, new_n961, new_n962,
    new_n963, new_n965, new_n966, new_n967, new_n968, new_n969, new_n970,
    new_n971, new_n972, new_n973, new_n974, new_n975, new_n976, new_n977,
    new_n978, new_n980, new_n981, new_n982, new_n983, new_n984, new_n985,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1017, new_n1018,
    new_n1019, new_n1020, new_n1021, new_n1022, new_n1023, new_n1024,
    new_n1025, new_n1026, new_n1028, new_n1029, new_n1030, new_n1031,
    new_n1032, new_n1033, new_n1034, new_n1035, new_n1036, new_n1037,
    new_n1038, new_n1039;
  NOR2_X1   g000(.A1(G237), .A2(G953), .ZN(new_n187));
  NAND2_X1  g001(.A1(new_n187), .A2(G210), .ZN(new_n188));
  XNOR2_X1  g002(.A(new_n188), .B(KEYINPUT27), .ZN(new_n189));
  XNOR2_X1  g003(.A(KEYINPUT26), .B(G101), .ZN(new_n190));
  XNOR2_X1  g004(.A(new_n189), .B(new_n190), .ZN(new_n191));
  INV_X1    g005(.A(KEYINPUT28), .ZN(new_n192));
  INV_X1    g006(.A(G146), .ZN(new_n193));
  OAI21_X1  g007(.A(KEYINPUT64), .B1(new_n193), .B2(G143), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n193), .A2(G143), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n194), .A2(new_n195), .ZN(new_n196));
  NAND3_X1  g010(.A1(new_n193), .A2(KEYINPUT64), .A3(G143), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n195), .A2(KEYINPUT1), .ZN(new_n198));
  AOI22_X1  g012(.A1(new_n196), .A2(new_n197), .B1(new_n198), .B2(G128), .ZN(new_n199));
  INV_X1    g013(.A(KEYINPUT1), .ZN(new_n200));
  INV_X1    g014(.A(G143), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n201), .A2(G146), .ZN(new_n202));
  AND4_X1   g016(.A1(new_n200), .A2(new_n195), .A3(new_n202), .A4(G128), .ZN(new_n203));
  OAI21_X1  g017(.A(KEYINPUT67), .B1(new_n199), .B2(new_n203), .ZN(new_n204));
  AND2_X1   g018(.A1(new_n195), .A2(new_n202), .ZN(new_n205));
  NAND3_X1  g019(.A1(new_n205), .A2(new_n200), .A3(G128), .ZN(new_n206));
  INV_X1    g020(.A(KEYINPUT67), .ZN(new_n207));
  INV_X1    g021(.A(new_n197), .ZN(new_n208));
  AOI21_X1  g022(.A(new_n208), .B1(new_n195), .B2(new_n194), .ZN(new_n209));
  INV_X1    g023(.A(G128), .ZN(new_n210));
  AOI21_X1  g024(.A(new_n210), .B1(new_n195), .B2(KEYINPUT1), .ZN(new_n211));
  OAI211_X1 g025(.A(new_n206), .B(new_n207), .C1(new_n209), .C2(new_n211), .ZN(new_n212));
  INV_X1    g026(.A(KEYINPUT65), .ZN(new_n213));
  INV_X1    g027(.A(G137), .ZN(new_n214));
  OAI21_X1  g028(.A(new_n213), .B1(new_n214), .B2(G134), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n214), .A2(G134), .ZN(new_n216));
  INV_X1    g030(.A(G134), .ZN(new_n217));
  NAND3_X1  g031(.A1(new_n217), .A2(KEYINPUT65), .A3(G137), .ZN(new_n218));
  NAND3_X1  g032(.A1(new_n215), .A2(new_n216), .A3(new_n218), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n219), .A2(G131), .ZN(new_n220));
  INV_X1    g034(.A(G131), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n217), .A2(G137), .ZN(new_n222));
  INV_X1    g036(.A(KEYINPUT11), .ZN(new_n223));
  AOI21_X1  g037(.A(new_n223), .B1(G134), .B2(new_n214), .ZN(new_n224));
  NOR3_X1   g038(.A1(new_n217), .A2(KEYINPUT11), .A3(G137), .ZN(new_n225));
  OAI211_X1 g039(.A(new_n221), .B(new_n222), .C1(new_n224), .C2(new_n225), .ZN(new_n226));
  AND3_X1   g040(.A1(new_n220), .A2(new_n226), .A3(KEYINPUT66), .ZN(new_n227));
  AOI21_X1  g041(.A(KEYINPUT66), .B1(new_n220), .B2(new_n226), .ZN(new_n228));
  OAI211_X1 g042(.A(new_n204), .B(new_n212), .C1(new_n227), .C2(new_n228), .ZN(new_n229));
  INV_X1    g043(.A(G119), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n230), .A2(G116), .ZN(new_n231));
  INV_X1    g045(.A(G116), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n232), .A2(G119), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n231), .A2(new_n233), .ZN(new_n234));
  INV_X1    g048(.A(new_n234), .ZN(new_n235));
  XNOR2_X1  g049(.A(KEYINPUT2), .B(G113), .ZN(new_n236));
  INV_X1    g050(.A(new_n236), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n235), .A2(new_n237), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n234), .A2(new_n236), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n238), .A2(new_n239), .ZN(new_n240));
  INV_X1    g054(.A(new_n240), .ZN(new_n241));
  OAI21_X1  g055(.A(new_n222), .B1(new_n224), .B2(new_n225), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n242), .A2(G131), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n243), .A2(new_n226), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n196), .A2(new_n197), .ZN(new_n245));
  AND2_X1   g059(.A1(KEYINPUT0), .A2(G128), .ZN(new_n246));
  NOR2_X1   g060(.A1(KEYINPUT0), .A2(G128), .ZN(new_n247));
  NOR2_X1   g061(.A1(new_n246), .A2(new_n247), .ZN(new_n248));
  AOI22_X1  g062(.A1(new_n245), .A2(new_n248), .B1(new_n246), .B2(new_n205), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n244), .A2(new_n249), .ZN(new_n250));
  NAND3_X1  g064(.A1(new_n229), .A2(new_n241), .A3(new_n250), .ZN(new_n251));
  OAI21_X1  g065(.A(new_n206), .B1(new_n209), .B2(new_n211), .ZN(new_n252));
  NAND3_X1  g066(.A1(new_n252), .A2(new_n226), .A3(new_n220), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n253), .A2(new_n250), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n254), .A2(new_n240), .ZN(new_n255));
  AOI21_X1  g069(.A(new_n192), .B1(new_n251), .B2(new_n255), .ZN(new_n256));
  INV_X1    g070(.A(new_n256), .ZN(new_n257));
  NAND3_X1  g071(.A1(new_n229), .A2(KEYINPUT70), .A3(new_n250), .ZN(new_n258));
  INV_X1    g072(.A(new_n258), .ZN(new_n259));
  AOI21_X1  g073(.A(KEYINPUT70), .B1(new_n229), .B2(new_n250), .ZN(new_n260));
  NOR3_X1   g074(.A1(new_n259), .A2(new_n260), .A3(new_n240), .ZN(new_n261));
  OAI211_X1 g075(.A(new_n191), .B(new_n257), .C1(new_n261), .C2(KEYINPUT28), .ZN(new_n262));
  INV_X1    g076(.A(KEYINPUT71), .ZN(new_n263));
  AOI21_X1  g077(.A(KEYINPUT29), .B1(new_n262), .B2(new_n263), .ZN(new_n264));
  INV_X1    g078(.A(new_n251), .ZN(new_n265));
  AOI21_X1  g079(.A(KEYINPUT30), .B1(new_n253), .B2(new_n250), .ZN(new_n266));
  NOR2_X1   g080(.A1(new_n266), .A2(new_n241), .ZN(new_n267));
  INV_X1    g081(.A(KEYINPUT30), .ZN(new_n268));
  AOI21_X1  g082(.A(new_n268), .B1(new_n244), .B2(new_n249), .ZN(new_n269));
  AND3_X1   g083(.A1(new_n229), .A2(KEYINPUT68), .A3(new_n269), .ZN(new_n270));
  AOI21_X1  g084(.A(KEYINPUT68), .B1(new_n229), .B2(new_n269), .ZN(new_n271));
  OAI21_X1  g085(.A(new_n267), .B1(new_n270), .B2(new_n271), .ZN(new_n272));
  INV_X1    g086(.A(KEYINPUT69), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n272), .A2(new_n273), .ZN(new_n274));
  OAI211_X1 g088(.A(new_n267), .B(KEYINPUT69), .C1(new_n270), .C2(new_n271), .ZN(new_n275));
  AOI211_X1 g089(.A(new_n191), .B(new_n265), .C1(new_n274), .C2(new_n275), .ZN(new_n276));
  INV_X1    g090(.A(new_n191), .ZN(new_n277));
  INV_X1    g091(.A(new_n260), .ZN(new_n278));
  NAND3_X1  g092(.A1(new_n278), .A2(new_n241), .A3(new_n258), .ZN(new_n279));
  AOI21_X1  g093(.A(new_n256), .B1(new_n279), .B2(new_n192), .ZN(new_n280));
  AOI21_X1  g094(.A(new_n277), .B1(new_n280), .B2(KEYINPUT71), .ZN(new_n281));
  OAI21_X1  g095(.A(new_n264), .B1(new_n276), .B2(new_n281), .ZN(new_n282));
  NOR2_X1   g096(.A1(new_n261), .A2(KEYINPUT28), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n229), .A2(new_n250), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n284), .A2(new_n240), .ZN(new_n285));
  AOI21_X1  g099(.A(new_n192), .B1(new_n285), .B2(new_n251), .ZN(new_n286));
  NOR2_X1   g100(.A1(new_n283), .A2(new_n286), .ZN(new_n287));
  AND2_X1   g101(.A1(new_n191), .A2(KEYINPUT29), .ZN(new_n288));
  AOI21_X1  g102(.A(G902), .B1(new_n287), .B2(new_n288), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n282), .A2(new_n289), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n290), .A2(G472), .ZN(new_n291));
  OAI21_X1  g105(.A(new_n277), .B1(new_n283), .B2(new_n256), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n274), .A2(new_n275), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n251), .A2(new_n191), .ZN(new_n294));
  INV_X1    g108(.A(new_n294), .ZN(new_n295));
  AOI21_X1  g109(.A(KEYINPUT31), .B1(new_n293), .B2(new_n295), .ZN(new_n296));
  INV_X1    g110(.A(KEYINPUT31), .ZN(new_n297));
  AOI211_X1 g111(.A(new_n297), .B(new_n294), .C1(new_n274), .C2(new_n275), .ZN(new_n298));
  OAI21_X1  g112(.A(new_n292), .B1(new_n296), .B2(new_n298), .ZN(new_n299));
  INV_X1    g113(.A(KEYINPUT32), .ZN(new_n300));
  NOR2_X1   g114(.A1(G472), .A2(G902), .ZN(new_n301));
  AND3_X1   g115(.A1(new_n299), .A2(new_n300), .A3(new_n301), .ZN(new_n302));
  AOI21_X1  g116(.A(new_n300), .B1(new_n299), .B2(new_n301), .ZN(new_n303));
  OAI21_X1  g117(.A(new_n291), .B1(new_n302), .B2(new_n303), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n304), .A2(KEYINPUT72), .ZN(new_n305));
  INV_X1    g119(.A(G902), .ZN(new_n306));
  XOR2_X1   g120(.A(KEYINPUT86), .B(G469), .Z(new_n307));
  INV_X1    g121(.A(G104), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n308), .A2(G107), .ZN(new_n309));
  INV_X1    g123(.A(new_n309), .ZN(new_n310));
  NOR2_X1   g124(.A1(new_n308), .A2(G107), .ZN(new_n311));
  OAI21_X1  g125(.A(G101), .B1(new_n310), .B2(new_n311), .ZN(new_n312));
  OAI21_X1  g126(.A(KEYINPUT3), .B1(new_n308), .B2(G107), .ZN(new_n313));
  INV_X1    g127(.A(KEYINPUT3), .ZN(new_n314));
  INV_X1    g128(.A(G107), .ZN(new_n315));
  NAND3_X1  g129(.A1(new_n314), .A2(new_n315), .A3(G104), .ZN(new_n316));
  INV_X1    g130(.A(G101), .ZN(new_n317));
  NAND4_X1  g131(.A1(new_n313), .A2(new_n316), .A3(new_n317), .A4(new_n309), .ZN(new_n318));
  AND3_X1   g132(.A1(new_n312), .A2(new_n318), .A3(KEYINPUT10), .ZN(new_n319));
  NAND3_X1  g133(.A1(new_n204), .A2(new_n212), .A3(new_n319), .ZN(new_n320));
  INV_X1    g134(.A(KEYINPUT83), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n320), .A2(new_n321), .ZN(new_n322));
  NAND4_X1  g136(.A1(new_n204), .A2(new_n212), .A3(KEYINPUT83), .A4(new_n319), .ZN(new_n323));
  NAND2_X1  g137(.A1(new_n322), .A2(new_n323), .ZN(new_n324));
  INV_X1    g138(.A(new_n244), .ZN(new_n325));
  NAND3_X1  g139(.A1(new_n313), .A2(new_n316), .A3(new_n309), .ZN(new_n326));
  INV_X1    g140(.A(KEYINPUT4), .ZN(new_n327));
  NAND3_X1  g141(.A1(new_n326), .A2(new_n327), .A3(G101), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n328), .A2(KEYINPUT81), .ZN(new_n329));
  INV_X1    g143(.A(KEYINPUT81), .ZN(new_n330));
  NAND4_X1  g144(.A1(new_n326), .A2(new_n330), .A3(new_n327), .A4(G101), .ZN(new_n331));
  AND2_X1   g145(.A1(new_n318), .A2(KEYINPUT4), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n326), .A2(G101), .ZN(new_n333));
  AOI22_X1  g147(.A1(new_n329), .A2(new_n331), .B1(new_n332), .B2(new_n333), .ZN(new_n334));
  OAI21_X1  g148(.A(new_n206), .B1(new_n205), .B2(new_n211), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n312), .A2(new_n318), .ZN(new_n336));
  INV_X1    g150(.A(new_n336), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n335), .A2(new_n337), .ZN(new_n338));
  XNOR2_X1  g152(.A(KEYINPUT82), .B(KEYINPUT10), .ZN(new_n339));
  AOI22_X1  g153(.A1(new_n334), .A2(new_n249), .B1(new_n338), .B2(new_n339), .ZN(new_n340));
  NAND3_X1  g154(.A1(new_n324), .A2(new_n325), .A3(new_n340), .ZN(new_n341));
  XNOR2_X1  g155(.A(G110), .B(G140), .ZN(new_n342));
  INV_X1    g156(.A(G953), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n343), .A2(G227), .ZN(new_n344));
  XOR2_X1   g158(.A(new_n342), .B(new_n344), .Z(new_n345));
  INV_X1    g159(.A(new_n345), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n341), .A2(new_n346), .ZN(new_n347));
  OAI21_X1  g161(.A(new_n338), .B1(new_n252), .B2(new_n337), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n348), .A2(new_n244), .ZN(new_n349));
  AOI21_X1  g163(.A(KEYINPUT12), .B1(new_n244), .B2(KEYINPUT84), .ZN(new_n350));
  INV_X1    g164(.A(new_n350), .ZN(new_n351));
  XNOR2_X1  g165(.A(new_n349), .B(new_n351), .ZN(new_n352));
  NOR2_X1   g166(.A1(new_n347), .A2(new_n352), .ZN(new_n353));
  NAND2_X1  g167(.A1(new_n324), .A2(new_n340), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n354), .A2(new_n244), .ZN(new_n355));
  AOI21_X1  g169(.A(new_n346), .B1(new_n355), .B2(new_n341), .ZN(new_n356));
  OAI211_X1 g170(.A(new_n306), .B(new_n307), .C1(new_n353), .C2(new_n356), .ZN(new_n357));
  INV_X1    g171(.A(KEYINPUT85), .ZN(new_n358));
  NAND2_X1  g172(.A1(new_n347), .A2(new_n358), .ZN(new_n359));
  NAND3_X1  g173(.A1(new_n341), .A2(KEYINPUT85), .A3(new_n346), .ZN(new_n360));
  NAND3_X1  g174(.A1(new_n359), .A2(new_n355), .A3(new_n360), .ZN(new_n361));
  XOR2_X1   g175(.A(new_n345), .B(KEYINPUT80), .Z(new_n362));
  INV_X1    g176(.A(new_n341), .ZN(new_n363));
  OAI21_X1  g177(.A(new_n362), .B1(new_n352), .B2(new_n363), .ZN(new_n364));
  AOI21_X1  g178(.A(G902), .B1(new_n361), .B2(new_n364), .ZN(new_n365));
  INV_X1    g179(.A(G469), .ZN(new_n366));
  OAI21_X1  g180(.A(new_n357), .B1(new_n365), .B2(new_n366), .ZN(new_n367));
  XNOR2_X1  g181(.A(KEYINPUT9), .B(G234), .ZN(new_n368));
  OAI21_X1  g182(.A(G221), .B1(new_n368), .B2(G902), .ZN(new_n369));
  AND2_X1   g183(.A1(new_n367), .A2(new_n369), .ZN(new_n370));
  INV_X1    g184(.A(G140), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n371), .A2(G125), .ZN(new_n372));
  INV_X1    g186(.A(G125), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n373), .A2(G140), .ZN(new_n374));
  INV_X1    g188(.A(KEYINPUT74), .ZN(new_n375));
  NAND3_X1  g189(.A1(new_n372), .A2(new_n374), .A3(new_n375), .ZN(new_n376));
  NAND3_X1  g190(.A1(new_n371), .A2(KEYINPUT74), .A3(G125), .ZN(new_n377));
  NAND3_X1  g191(.A1(new_n376), .A2(G146), .A3(new_n377), .ZN(new_n378));
  AND2_X1   g192(.A1(new_n372), .A2(new_n374), .ZN(new_n379));
  NAND2_X1  g193(.A1(new_n379), .A2(new_n193), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n378), .A2(new_n380), .ZN(new_n381));
  INV_X1    g195(.A(G237), .ZN(new_n382));
  AND4_X1   g196(.A1(G143), .A2(new_n382), .A3(new_n343), .A4(G214), .ZN(new_n383));
  AOI21_X1  g197(.A(G143), .B1(new_n187), .B2(G214), .ZN(new_n384));
  NOR2_X1   g198(.A1(new_n383), .A2(new_n384), .ZN(new_n385));
  NAND2_X1  g199(.A1(KEYINPUT18), .A2(G131), .ZN(new_n386));
  NAND2_X1  g200(.A1(new_n385), .A2(new_n386), .ZN(new_n387));
  NAND3_X1  g201(.A1(new_n382), .A2(new_n343), .A3(G214), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n388), .A2(new_n201), .ZN(new_n389));
  NAND3_X1  g203(.A1(new_n187), .A2(G143), .A3(G214), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n389), .A2(new_n390), .ZN(new_n391));
  INV_X1    g205(.A(new_n386), .ZN(new_n392));
  AOI21_X1  g206(.A(KEYINPUT92), .B1(new_n391), .B2(new_n392), .ZN(new_n393));
  INV_X1    g207(.A(KEYINPUT92), .ZN(new_n394));
  AOI211_X1 g208(.A(new_n394), .B(new_n386), .C1(new_n389), .C2(new_n390), .ZN(new_n395));
  OAI211_X1 g209(.A(new_n381), .B(new_n387), .C1(new_n393), .C2(new_n395), .ZN(new_n396));
  XNOR2_X1  g210(.A(G113), .B(G122), .ZN(new_n397));
  XNOR2_X1  g211(.A(new_n397), .B(new_n308), .ZN(new_n398));
  XOR2_X1   g212(.A(new_n398), .B(KEYINPUT95), .Z(new_n399));
  NAND3_X1  g213(.A1(new_n376), .A2(KEYINPUT16), .A3(new_n377), .ZN(new_n400));
  INV_X1    g214(.A(KEYINPUT16), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n372), .A2(new_n401), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n400), .A2(new_n402), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n403), .A2(G146), .ZN(new_n404));
  INV_X1    g218(.A(KEYINPUT75), .ZN(new_n405));
  NAND3_X1  g219(.A1(new_n400), .A2(new_n193), .A3(new_n402), .ZN(new_n406));
  NAND3_X1  g220(.A1(new_n404), .A2(new_n405), .A3(new_n406), .ZN(new_n407));
  NAND3_X1  g221(.A1(new_n403), .A2(KEYINPUT75), .A3(G146), .ZN(new_n408));
  AND2_X1   g222(.A1(new_n407), .A2(new_n408), .ZN(new_n409));
  INV_X1    g223(.A(KEYINPUT17), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n385), .A2(new_n221), .ZN(new_n411));
  INV_X1    g225(.A(KEYINPUT93), .ZN(new_n412));
  AOI21_X1  g226(.A(new_n412), .B1(new_n391), .B2(G131), .ZN(new_n413));
  AOI211_X1 g227(.A(KEYINPUT93), .B(new_n221), .C1(new_n389), .C2(new_n390), .ZN(new_n414));
  OAI211_X1 g228(.A(new_n410), .B(new_n411), .C1(new_n413), .C2(new_n414), .ZN(new_n415));
  OAI21_X1  g229(.A(G131), .B1(new_n383), .B2(new_n384), .ZN(new_n416));
  NAND2_X1  g230(.A1(new_n416), .A2(KEYINPUT93), .ZN(new_n417));
  NAND3_X1  g231(.A1(new_n391), .A2(new_n412), .A3(G131), .ZN(new_n418));
  NAND3_X1  g232(.A1(new_n417), .A2(KEYINPUT17), .A3(new_n418), .ZN(new_n419));
  NAND2_X1  g233(.A1(new_n415), .A2(new_n419), .ZN(new_n420));
  OAI211_X1 g234(.A(new_n396), .B(new_n399), .C1(new_n409), .C2(new_n420), .ZN(new_n421));
  AND2_X1   g235(.A1(new_n415), .A2(new_n419), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n407), .A2(new_n408), .ZN(new_n423));
  OR2_X1    g237(.A1(new_n393), .A2(new_n395), .ZN(new_n424));
  AND2_X1   g238(.A1(new_n381), .A2(new_n387), .ZN(new_n425));
  AOI22_X1  g239(.A1(new_n422), .A2(new_n423), .B1(new_n424), .B2(new_n425), .ZN(new_n426));
  OAI21_X1  g240(.A(new_n421), .B1(new_n426), .B2(new_n398), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n427), .A2(new_n306), .ZN(new_n428));
  XOR2_X1   g242(.A(KEYINPUT96), .B(G475), .Z(new_n429));
  INV_X1    g243(.A(new_n429), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n428), .A2(new_n430), .ZN(new_n431));
  INV_X1    g245(.A(KEYINPUT19), .ZN(new_n432));
  AOI21_X1  g246(.A(new_n432), .B1(new_n376), .B2(new_n377), .ZN(new_n433));
  NOR2_X1   g247(.A1(new_n379), .A2(KEYINPUT19), .ZN(new_n434));
  OAI21_X1  g248(.A(new_n193), .B1(new_n433), .B2(new_n434), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n404), .A2(new_n435), .ZN(new_n436));
  AOI22_X1  g250(.A1(new_n417), .A2(new_n418), .B1(new_n221), .B2(new_n385), .ZN(new_n437));
  OAI21_X1  g251(.A(new_n396), .B1(new_n436), .B2(new_n437), .ZN(new_n438));
  INV_X1    g252(.A(KEYINPUT94), .ZN(new_n439));
  INV_X1    g253(.A(new_n398), .ZN(new_n440));
  AND3_X1   g254(.A1(new_n438), .A2(new_n439), .A3(new_n440), .ZN(new_n441));
  AOI21_X1  g255(.A(new_n439), .B1(new_n438), .B2(new_n440), .ZN(new_n442));
  OAI21_X1  g256(.A(new_n421), .B1(new_n441), .B2(new_n442), .ZN(new_n443));
  INV_X1    g257(.A(KEYINPUT20), .ZN(new_n444));
  NOR2_X1   g258(.A1(G475), .A2(G902), .ZN(new_n445));
  AND3_X1   g259(.A1(new_n443), .A2(new_n444), .A3(new_n445), .ZN(new_n446));
  XOR2_X1   g260(.A(KEYINPUT91), .B(KEYINPUT20), .Z(new_n447));
  AOI21_X1  g261(.A(new_n447), .B1(new_n443), .B2(new_n445), .ZN(new_n448));
  OAI21_X1  g262(.A(new_n431), .B1(new_n446), .B2(new_n448), .ZN(new_n449));
  INV_X1    g263(.A(G478), .ZN(new_n450));
  NOR2_X1   g264(.A1(new_n450), .A2(KEYINPUT15), .ZN(new_n451));
  INV_X1    g265(.A(G122), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n452), .A2(G116), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n232), .A2(G122), .ZN(new_n454));
  NAND3_X1  g268(.A1(new_n453), .A2(new_n454), .A3(new_n315), .ZN(new_n455));
  NOR2_X1   g269(.A1(new_n201), .A2(G128), .ZN(new_n456));
  INV_X1    g270(.A(KEYINPUT97), .ZN(new_n457));
  NAND3_X1  g271(.A1(new_n457), .A2(new_n201), .A3(G128), .ZN(new_n458));
  OAI21_X1  g272(.A(KEYINPUT97), .B1(new_n210), .B2(G143), .ZN(new_n459));
  AOI211_X1 g273(.A(G134), .B(new_n456), .C1(new_n458), .C2(new_n459), .ZN(new_n460));
  NAND2_X1  g274(.A1(new_n459), .A2(new_n458), .ZN(new_n461));
  INV_X1    g275(.A(new_n456), .ZN(new_n462));
  AOI21_X1  g276(.A(new_n217), .B1(new_n461), .B2(new_n462), .ZN(new_n463));
  OAI21_X1  g277(.A(new_n455), .B1(new_n460), .B2(new_n463), .ZN(new_n464));
  OAI21_X1  g278(.A(KEYINPUT14), .B1(new_n452), .B2(G116), .ZN(new_n465));
  NAND2_X1  g279(.A1(new_n465), .A2(KEYINPUT98), .ZN(new_n466));
  INV_X1    g280(.A(KEYINPUT98), .ZN(new_n467));
  NAND3_X1  g281(.A1(new_n454), .A2(new_n467), .A3(KEYINPUT14), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n466), .A2(new_n468), .ZN(new_n469));
  NOR2_X1   g283(.A1(new_n232), .A2(G122), .ZN(new_n470));
  INV_X1    g284(.A(new_n454), .ZN(new_n471));
  INV_X1    g285(.A(KEYINPUT14), .ZN(new_n472));
  AOI21_X1  g286(.A(new_n470), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  AOI21_X1  g287(.A(new_n315), .B1(new_n469), .B2(new_n473), .ZN(new_n474));
  INV_X1    g288(.A(KEYINPUT13), .ZN(new_n475));
  AOI21_X1  g289(.A(new_n456), .B1(new_n461), .B2(new_n475), .ZN(new_n476));
  NAND3_X1  g290(.A1(new_n459), .A2(new_n458), .A3(KEYINPUT13), .ZN(new_n477));
  AOI21_X1  g291(.A(new_n217), .B1(new_n476), .B2(new_n477), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n453), .A2(new_n454), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n479), .A2(G107), .ZN(new_n480));
  NAND2_X1  g294(.A1(new_n480), .A2(new_n455), .ZN(new_n481));
  AOI21_X1  g295(.A(new_n456), .B1(new_n459), .B2(new_n458), .ZN(new_n482));
  NAND2_X1  g296(.A1(new_n482), .A2(new_n217), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n481), .A2(new_n483), .ZN(new_n484));
  OAI22_X1  g298(.A1(new_n464), .A2(new_n474), .B1(new_n478), .B2(new_n484), .ZN(new_n485));
  INV_X1    g299(.A(G217), .ZN(new_n486));
  NOR3_X1   g300(.A1(new_n368), .A2(new_n486), .A3(G953), .ZN(new_n487));
  INV_X1    g301(.A(new_n487), .ZN(new_n488));
  NAND2_X1  g302(.A1(new_n485), .A2(new_n488), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n461), .A2(new_n462), .ZN(new_n490));
  NAND2_X1  g304(.A1(new_n490), .A2(G134), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n491), .A2(new_n483), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n469), .A2(new_n473), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n493), .A2(G107), .ZN(new_n494));
  NAND3_X1  g308(.A1(new_n492), .A2(new_n494), .A3(new_n455), .ZN(new_n495));
  AOI22_X1  g309(.A1(new_n480), .A2(new_n455), .B1(new_n482), .B2(new_n217), .ZN(new_n496));
  AND3_X1   g310(.A1(new_n459), .A2(new_n458), .A3(KEYINPUT13), .ZN(new_n497));
  AOI21_X1  g311(.A(KEYINPUT13), .B1(new_n459), .B2(new_n458), .ZN(new_n498));
  NOR3_X1   g312(.A1(new_n497), .A2(new_n498), .A3(new_n456), .ZN(new_n499));
  OAI21_X1  g313(.A(new_n496), .B1(new_n499), .B2(new_n217), .ZN(new_n500));
  NAND4_X1  g314(.A1(new_n495), .A2(KEYINPUT99), .A3(new_n500), .A4(new_n487), .ZN(new_n501));
  NAND2_X1  g315(.A1(new_n489), .A2(new_n501), .ZN(new_n502));
  INV_X1    g316(.A(new_n455), .ZN(new_n503));
  AOI21_X1  g317(.A(new_n503), .B1(new_n491), .B2(new_n483), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n461), .A2(new_n475), .ZN(new_n505));
  NAND3_X1  g319(.A1(new_n505), .A2(new_n477), .A3(new_n462), .ZN(new_n506));
  NAND2_X1  g320(.A1(new_n506), .A2(G134), .ZN(new_n507));
  AOI22_X1  g321(.A1(new_n494), .A2(new_n504), .B1(new_n507), .B2(new_n496), .ZN(new_n508));
  AOI21_X1  g322(.A(KEYINPUT99), .B1(new_n508), .B2(new_n487), .ZN(new_n509));
  OAI21_X1  g323(.A(new_n306), .B1(new_n502), .B2(new_n509), .ZN(new_n510));
  NAND2_X1  g324(.A1(new_n510), .A2(KEYINPUT100), .ZN(new_n511));
  INV_X1    g325(.A(KEYINPUT100), .ZN(new_n512));
  OAI211_X1 g326(.A(new_n512), .B(new_n306), .C1(new_n502), .C2(new_n509), .ZN(new_n513));
  AOI21_X1  g327(.A(new_n451), .B1(new_n511), .B2(new_n513), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n513), .A2(new_n451), .ZN(new_n515));
  INV_X1    g329(.A(new_n515), .ZN(new_n516));
  OAI21_X1  g330(.A(KEYINPUT101), .B1(new_n514), .B2(new_n516), .ZN(new_n517));
  INV_X1    g331(.A(new_n451), .ZN(new_n518));
  INV_X1    g332(.A(new_n513), .ZN(new_n519));
  INV_X1    g333(.A(KEYINPUT99), .ZN(new_n520));
  OAI21_X1  g334(.A(new_n520), .B1(new_n485), .B2(new_n488), .ZN(new_n521));
  NAND3_X1  g335(.A1(new_n521), .A2(new_n489), .A3(new_n501), .ZN(new_n522));
  AOI21_X1  g336(.A(new_n512), .B1(new_n522), .B2(new_n306), .ZN(new_n523));
  OAI21_X1  g337(.A(new_n518), .B1(new_n519), .B2(new_n523), .ZN(new_n524));
  INV_X1    g338(.A(KEYINPUT101), .ZN(new_n525));
  NAND3_X1  g339(.A1(new_n524), .A2(new_n525), .A3(new_n515), .ZN(new_n526));
  AOI21_X1  g340(.A(new_n449), .B1(new_n517), .B2(new_n526), .ZN(new_n527));
  INV_X1    g341(.A(KEYINPUT6), .ZN(new_n528));
  AND3_X1   g342(.A1(new_n231), .A2(new_n233), .A3(KEYINPUT5), .ZN(new_n529));
  OAI21_X1  g343(.A(G113), .B1(new_n231), .B2(KEYINPUT5), .ZN(new_n530));
  OAI21_X1  g344(.A(new_n238), .B1(new_n529), .B2(new_n530), .ZN(new_n531));
  NOR2_X1   g345(.A1(new_n531), .A2(new_n336), .ZN(new_n532));
  AOI21_X1  g346(.A(new_n532), .B1(new_n334), .B2(new_n240), .ZN(new_n533));
  XNOR2_X1  g347(.A(G110), .B(G122), .ZN(new_n534));
  AOI21_X1  g348(.A(new_n528), .B1(new_n533), .B2(new_n534), .ZN(new_n535));
  INV_X1    g349(.A(new_n534), .ZN(new_n536));
  OAI21_X1  g350(.A(new_n536), .B1(new_n533), .B2(KEYINPUT87), .ZN(new_n537));
  NAND2_X1  g351(.A1(new_n329), .A2(new_n331), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n332), .A2(new_n333), .ZN(new_n539));
  NAND3_X1  g353(.A1(new_n538), .A2(new_n240), .A3(new_n539), .ZN(new_n540));
  INV_X1    g354(.A(new_n529), .ZN(new_n541));
  INV_X1    g355(.A(new_n530), .ZN(new_n542));
  AOI22_X1  g356(.A1(new_n541), .A2(new_n542), .B1(new_n237), .B2(new_n235), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n543), .A2(new_n337), .ZN(new_n544));
  NAND2_X1  g358(.A1(new_n540), .A2(new_n544), .ZN(new_n545));
  INV_X1    g359(.A(KEYINPUT87), .ZN(new_n546));
  NOR2_X1   g360(.A1(new_n545), .A2(new_n546), .ZN(new_n547));
  OAI21_X1  g361(.A(new_n535), .B1(new_n537), .B2(new_n547), .ZN(new_n548));
  AOI21_X1  g362(.A(new_n534), .B1(new_n545), .B2(new_n546), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n533), .A2(KEYINPUT87), .ZN(new_n550));
  NAND3_X1  g364(.A1(new_n549), .A2(new_n528), .A3(new_n550), .ZN(new_n551));
  OAI211_X1 g365(.A(new_n206), .B(new_n373), .C1(new_n209), .C2(new_n211), .ZN(new_n552));
  OAI21_X1  g366(.A(new_n552), .B1(new_n249), .B2(new_n373), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n553), .A2(KEYINPUT88), .ZN(new_n554));
  INV_X1    g368(.A(KEYINPUT88), .ZN(new_n555));
  OAI21_X1  g369(.A(new_n555), .B1(new_n249), .B2(new_n373), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n554), .A2(new_n556), .ZN(new_n557));
  INV_X1    g371(.A(G224), .ZN(new_n558));
  NOR2_X1   g372(.A1(new_n558), .A2(G953), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n557), .A2(new_n559), .ZN(new_n560));
  INV_X1    g374(.A(new_n559), .ZN(new_n561));
  NAND3_X1  g375(.A1(new_n554), .A2(new_n561), .A3(new_n556), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n560), .A2(new_n562), .ZN(new_n563));
  NAND3_X1  g377(.A1(new_n548), .A2(new_n551), .A3(new_n563), .ZN(new_n564));
  NAND4_X1  g378(.A1(new_n554), .A2(KEYINPUT7), .A3(new_n561), .A4(new_n556), .ZN(new_n565));
  OAI21_X1  g379(.A(KEYINPUT90), .B1(new_n531), .B2(new_n336), .ZN(new_n566));
  INV_X1    g380(.A(KEYINPUT90), .ZN(new_n567));
  NAND3_X1  g381(.A1(new_n543), .A2(new_n337), .A3(new_n567), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n531), .A2(new_n336), .ZN(new_n569));
  NAND3_X1  g383(.A1(new_n566), .A2(new_n568), .A3(new_n569), .ZN(new_n570));
  XNOR2_X1  g384(.A(new_n534), .B(KEYINPUT89), .ZN(new_n571));
  XOR2_X1   g385(.A(new_n571), .B(KEYINPUT8), .Z(new_n572));
  NAND2_X1  g386(.A1(new_n570), .A2(new_n572), .ZN(new_n573));
  NAND3_X1  g387(.A1(new_n540), .A2(new_n544), .A3(new_n534), .ZN(new_n574));
  INV_X1    g388(.A(KEYINPUT7), .ZN(new_n575));
  OAI21_X1  g389(.A(new_n553), .B1(new_n575), .B2(new_n559), .ZN(new_n576));
  NAND4_X1  g390(.A1(new_n565), .A2(new_n573), .A3(new_n574), .A4(new_n576), .ZN(new_n577));
  AND2_X1   g391(.A1(new_n577), .A2(new_n306), .ZN(new_n578));
  NAND2_X1  g392(.A1(new_n564), .A2(new_n578), .ZN(new_n579));
  OAI21_X1  g393(.A(G210), .B1(G237), .B2(G902), .ZN(new_n580));
  INV_X1    g394(.A(new_n580), .ZN(new_n581));
  NAND2_X1  g395(.A1(new_n579), .A2(new_n581), .ZN(new_n582));
  NAND3_X1  g396(.A1(new_n564), .A2(new_n578), .A3(new_n580), .ZN(new_n583));
  NAND2_X1  g397(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  OAI21_X1  g398(.A(G214), .B1(G237), .B2(G902), .ZN(new_n585));
  AND2_X1   g399(.A1(new_n343), .A2(G952), .ZN(new_n586));
  INV_X1    g400(.A(G234), .ZN(new_n587));
  OAI21_X1  g401(.A(new_n586), .B1(new_n587), .B2(new_n382), .ZN(new_n588));
  INV_X1    g402(.A(new_n588), .ZN(new_n589));
  AOI211_X1 g403(.A(new_n306), .B(new_n343), .C1(G234), .C2(G237), .ZN(new_n590));
  XNOR2_X1  g404(.A(KEYINPUT21), .B(G898), .ZN(new_n591));
  AOI21_X1  g405(.A(new_n589), .B1(new_n590), .B2(new_n591), .ZN(new_n592));
  INV_X1    g406(.A(new_n592), .ZN(new_n593));
  NAND3_X1  g407(.A1(new_n584), .A2(new_n585), .A3(new_n593), .ZN(new_n594));
  INV_X1    g408(.A(new_n594), .ZN(new_n595));
  AND3_X1   g409(.A1(new_n370), .A2(new_n527), .A3(new_n595), .ZN(new_n596));
  INV_X1    g410(.A(KEYINPUT23), .ZN(new_n597));
  OAI21_X1  g411(.A(new_n597), .B1(new_n230), .B2(G128), .ZN(new_n598));
  NAND3_X1  g412(.A1(new_n210), .A2(KEYINPUT23), .A3(G119), .ZN(new_n599));
  OAI211_X1 g413(.A(new_n598), .B(new_n599), .C1(G119), .C2(new_n210), .ZN(new_n600));
  NAND2_X1  g414(.A1(new_n600), .A2(G110), .ZN(new_n601));
  INV_X1    g415(.A(KEYINPUT73), .ZN(new_n602));
  XNOR2_X1  g416(.A(new_n601), .B(new_n602), .ZN(new_n603));
  XOR2_X1   g417(.A(G119), .B(G128), .Z(new_n604));
  XNOR2_X1  g418(.A(KEYINPUT24), .B(G110), .ZN(new_n605));
  OR2_X1    g419(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  NAND4_X1  g420(.A1(new_n407), .A2(new_n603), .A3(new_n408), .A4(new_n606), .ZN(new_n607));
  NOR2_X1   g421(.A1(new_n600), .A2(G110), .ZN(new_n608));
  AND2_X1   g422(.A1(new_n604), .A2(new_n605), .ZN(new_n609));
  OAI211_X1 g423(.A(new_n404), .B(new_n380), .C1(new_n608), .C2(new_n609), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n607), .A2(new_n610), .ZN(new_n611));
  NAND2_X1  g425(.A1(new_n611), .A2(KEYINPUT77), .ZN(new_n612));
  INV_X1    g426(.A(KEYINPUT77), .ZN(new_n613));
  NAND3_X1  g427(.A1(new_n607), .A2(new_n613), .A3(new_n610), .ZN(new_n614));
  NAND3_X1  g428(.A1(new_n343), .A2(G221), .A3(G234), .ZN(new_n615));
  XNOR2_X1  g429(.A(new_n615), .B(KEYINPUT76), .ZN(new_n616));
  XNOR2_X1  g430(.A(KEYINPUT22), .B(G137), .ZN(new_n617));
  XNOR2_X1  g431(.A(new_n616), .B(new_n617), .ZN(new_n618));
  INV_X1    g432(.A(new_n618), .ZN(new_n619));
  NAND3_X1  g433(.A1(new_n612), .A2(new_n614), .A3(new_n619), .ZN(new_n620));
  NAND3_X1  g434(.A1(new_n611), .A2(KEYINPUT77), .A3(new_n618), .ZN(new_n621));
  NAND2_X1  g435(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  NAND2_X1  g436(.A1(new_n622), .A2(new_n306), .ZN(new_n623));
  NAND3_X1  g437(.A1(new_n623), .A2(KEYINPUT78), .A3(KEYINPUT25), .ZN(new_n624));
  AOI21_X1  g438(.A(new_n486), .B1(G234), .B2(new_n306), .ZN(new_n625));
  INV_X1    g439(.A(KEYINPUT25), .ZN(new_n626));
  AOI21_X1  g440(.A(G902), .B1(new_n620), .B2(new_n621), .ZN(new_n627));
  INV_X1    g441(.A(KEYINPUT78), .ZN(new_n628));
  OAI21_X1  g442(.A(new_n626), .B1(new_n627), .B2(new_n628), .ZN(new_n629));
  NAND3_X1  g443(.A1(new_n624), .A2(new_n625), .A3(new_n629), .ZN(new_n630));
  NOR2_X1   g444(.A1(new_n625), .A2(G902), .ZN(new_n631));
  XOR2_X1   g445(.A(new_n631), .B(KEYINPUT79), .Z(new_n632));
  NAND2_X1  g446(.A1(new_n622), .A2(new_n632), .ZN(new_n633));
  NAND2_X1  g447(.A1(new_n630), .A2(new_n633), .ZN(new_n634));
  INV_X1    g448(.A(new_n634), .ZN(new_n635));
  INV_X1    g449(.A(KEYINPUT72), .ZN(new_n636));
  OAI211_X1 g450(.A(new_n291), .B(new_n636), .C1(new_n302), .C2(new_n303), .ZN(new_n637));
  NAND4_X1  g451(.A1(new_n305), .A2(new_n596), .A3(new_n635), .A4(new_n637), .ZN(new_n638));
  XNOR2_X1  g452(.A(new_n638), .B(G101), .ZN(G3));
  NAND2_X1  g453(.A1(new_n299), .A2(new_n306), .ZN(new_n640));
  NAND2_X1  g454(.A1(new_n640), .A2(G472), .ZN(new_n641));
  NAND2_X1  g455(.A1(new_n299), .A2(new_n301), .ZN(new_n642));
  NAND2_X1  g456(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  NOR2_X1   g457(.A1(new_n643), .A2(new_n634), .ZN(new_n644));
  AND3_X1   g458(.A1(new_n564), .A2(new_n578), .A3(new_n580), .ZN(new_n645));
  AOI21_X1  g459(.A(new_n580), .B1(new_n564), .B2(new_n578), .ZN(new_n646));
  OAI21_X1  g460(.A(new_n585), .B1(new_n645), .B2(new_n646), .ZN(new_n647));
  NAND2_X1  g461(.A1(new_n647), .A2(KEYINPUT102), .ZN(new_n648));
  INV_X1    g462(.A(KEYINPUT102), .ZN(new_n649));
  OAI211_X1 g463(.A(new_n649), .B(new_n585), .C1(new_n645), .C2(new_n646), .ZN(new_n650));
  NAND2_X1  g464(.A1(new_n648), .A2(new_n650), .ZN(new_n651));
  AOI21_X1  g465(.A(new_n429), .B1(new_n427), .B2(new_n306), .ZN(new_n652));
  INV_X1    g466(.A(new_n447), .ZN(new_n653));
  NAND2_X1  g467(.A1(new_n438), .A2(new_n440), .ZN(new_n654));
  NAND2_X1  g468(.A1(new_n654), .A2(KEYINPUT94), .ZN(new_n655));
  NAND3_X1  g469(.A1(new_n438), .A2(new_n439), .A3(new_n440), .ZN(new_n656));
  AOI22_X1  g470(.A1(new_n655), .A2(new_n656), .B1(new_n426), .B2(new_n399), .ZN(new_n657));
  INV_X1    g471(.A(new_n445), .ZN(new_n658));
  OAI21_X1  g472(.A(new_n653), .B1(new_n657), .B2(new_n658), .ZN(new_n659));
  NAND3_X1  g473(.A1(new_n443), .A2(new_n444), .A3(new_n445), .ZN(new_n660));
  AOI21_X1  g474(.A(new_n652), .B1(new_n659), .B2(new_n660), .ZN(new_n661));
  NOR2_X1   g475(.A1(new_n450), .A2(G902), .ZN(new_n662));
  INV_X1    g476(.A(new_n662), .ZN(new_n663));
  OR3_X1    g477(.A1(new_n502), .A2(new_n509), .A3(KEYINPUT33), .ZN(new_n664));
  NAND3_X1  g478(.A1(new_n508), .A2(KEYINPUT103), .A3(new_n487), .ZN(new_n665));
  NAND2_X1  g479(.A1(new_n665), .A2(new_n489), .ZN(new_n666));
  AOI21_X1  g480(.A(KEYINPUT103), .B1(new_n508), .B2(new_n487), .ZN(new_n667));
  OAI21_X1  g481(.A(KEYINPUT33), .B1(new_n666), .B2(new_n667), .ZN(new_n668));
  AOI21_X1  g482(.A(new_n663), .B1(new_n664), .B2(new_n668), .ZN(new_n669));
  AOI21_X1  g483(.A(G478), .B1(new_n522), .B2(new_n306), .ZN(new_n670));
  NOR2_X1   g484(.A1(new_n669), .A2(new_n670), .ZN(new_n671));
  NOR2_X1   g485(.A1(new_n661), .A2(new_n671), .ZN(new_n672));
  AND3_X1   g486(.A1(new_n651), .A2(new_n593), .A3(new_n672), .ZN(new_n673));
  NAND3_X1  g487(.A1(new_n644), .A2(new_n370), .A3(new_n673), .ZN(new_n674));
  XNOR2_X1  g488(.A(new_n674), .B(G104), .ZN(new_n675));
  XOR2_X1   g489(.A(KEYINPUT104), .B(KEYINPUT34), .Z(new_n676));
  XNOR2_X1  g490(.A(new_n675), .B(new_n676), .ZN(G6));
  NAND3_X1  g491(.A1(new_n443), .A2(new_n445), .A3(new_n447), .ZN(new_n678));
  AOI21_X1  g492(.A(new_n652), .B1(new_n659), .B2(new_n678), .ZN(new_n679));
  AND3_X1   g493(.A1(new_n517), .A2(new_n679), .A3(new_n526), .ZN(new_n680));
  AND3_X1   g494(.A1(new_n651), .A2(new_n593), .A3(new_n680), .ZN(new_n681));
  NAND3_X1  g495(.A1(new_n644), .A2(new_n370), .A3(new_n681), .ZN(new_n682));
  XOR2_X1   g496(.A(KEYINPUT35), .B(G107), .Z(new_n683));
  XNOR2_X1  g497(.A(new_n682), .B(new_n683), .ZN(G9));
  NOR2_X1   g498(.A1(new_n619), .A2(KEYINPUT36), .ZN(new_n685));
  XNOR2_X1  g499(.A(new_n611), .B(new_n685), .ZN(new_n686));
  NAND2_X1  g500(.A1(new_n686), .A2(new_n632), .ZN(new_n687));
  NAND2_X1  g501(.A1(new_n630), .A2(new_n687), .ZN(new_n688));
  INV_X1    g502(.A(new_n688), .ZN(new_n689));
  NOR2_X1   g503(.A1(new_n643), .A2(new_n689), .ZN(new_n690));
  NAND2_X1  g504(.A1(new_n690), .A2(new_n596), .ZN(new_n691));
  XOR2_X1   g505(.A(KEYINPUT37), .B(G110), .Z(new_n692));
  XNOR2_X1  g506(.A(new_n691), .B(new_n692), .ZN(G12));
  AOI21_X1  g507(.A(new_n649), .B1(new_n584), .B2(new_n585), .ZN(new_n694));
  INV_X1    g508(.A(new_n650), .ZN(new_n695));
  OAI21_X1  g509(.A(new_n688), .B1(new_n694), .B2(new_n695), .ZN(new_n696));
  INV_X1    g510(.A(G900), .ZN(new_n697));
  AOI21_X1  g511(.A(new_n589), .B1(new_n590), .B2(new_n697), .ZN(new_n698));
  INV_X1    g512(.A(new_n698), .ZN(new_n699));
  NAND4_X1  g513(.A1(new_n680), .A2(new_n369), .A3(new_n367), .A4(new_n699), .ZN(new_n700));
  NOR2_X1   g514(.A1(new_n696), .A2(new_n700), .ZN(new_n701));
  NAND3_X1  g515(.A1(new_n305), .A2(new_n637), .A3(new_n701), .ZN(new_n702));
  INV_X1    g516(.A(KEYINPUT105), .ZN(new_n703));
  NAND2_X1  g517(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  NAND4_X1  g518(.A1(new_n305), .A2(new_n701), .A3(KEYINPUT105), .A4(new_n637), .ZN(new_n705));
  NAND2_X1  g519(.A1(new_n704), .A2(new_n705), .ZN(new_n706));
  XNOR2_X1  g520(.A(new_n706), .B(G128), .ZN(G30));
  XOR2_X1   g521(.A(new_n698), .B(KEYINPUT39), .Z(new_n708));
  NAND2_X1  g522(.A1(new_n370), .A2(new_n708), .ZN(new_n709));
  INV_X1    g523(.A(KEYINPUT40), .ZN(new_n710));
  NAND2_X1  g524(.A1(new_n709), .A2(new_n710), .ZN(new_n711));
  NAND3_X1  g525(.A1(new_n370), .A2(KEYINPUT40), .A3(new_n708), .ZN(new_n712));
  NAND2_X1  g526(.A1(new_n711), .A2(new_n712), .ZN(new_n713));
  NAND2_X1  g527(.A1(new_n713), .A2(KEYINPUT108), .ZN(new_n714));
  AOI21_X1  g528(.A(new_n191), .B1(new_n285), .B2(new_n251), .ZN(new_n715));
  XNOR2_X1  g529(.A(new_n715), .B(KEYINPUT106), .ZN(new_n716));
  AOI21_X1  g530(.A(new_n294), .B1(new_n274), .B2(new_n275), .ZN(new_n717));
  OAI21_X1  g531(.A(new_n306), .B1(new_n716), .B2(new_n717), .ZN(new_n718));
  NAND2_X1  g532(.A1(new_n718), .A2(G472), .ZN(new_n719));
  OAI21_X1  g533(.A(new_n719), .B1(new_n302), .B2(new_n303), .ZN(new_n720));
  INV_X1    g534(.A(new_n720), .ZN(new_n721));
  INV_X1    g535(.A(KEYINPUT38), .ZN(new_n722));
  XNOR2_X1  g536(.A(new_n584), .B(new_n722), .ZN(new_n723));
  NOR2_X1   g537(.A1(new_n721), .A2(new_n723), .ZN(new_n724));
  INV_X1    g538(.A(KEYINPUT108), .ZN(new_n725));
  NAND3_X1  g539(.A1(new_n711), .A2(new_n725), .A3(new_n712), .ZN(new_n726));
  INV_X1    g540(.A(new_n585), .ZN(new_n727));
  NAND3_X1  g541(.A1(new_n517), .A2(new_n449), .A3(new_n526), .ZN(new_n728));
  NOR3_X1   g542(.A1(new_n688), .A2(new_n727), .A3(new_n728), .ZN(new_n729));
  XNOR2_X1  g543(.A(new_n729), .B(KEYINPUT107), .ZN(new_n730));
  NAND4_X1  g544(.A1(new_n714), .A2(new_n724), .A3(new_n726), .A4(new_n730), .ZN(new_n731));
  XNOR2_X1  g545(.A(new_n731), .B(G143), .ZN(G45));
  NOR3_X1   g546(.A1(new_n661), .A2(new_n671), .A3(new_n698), .ZN(new_n733));
  NAND3_X1  g547(.A1(new_n733), .A2(new_n367), .A3(new_n369), .ZN(new_n734));
  NOR2_X1   g548(.A1(new_n696), .A2(new_n734), .ZN(new_n735));
  NAND3_X1  g549(.A1(new_n305), .A2(new_n637), .A3(new_n735), .ZN(new_n736));
  NAND2_X1  g550(.A1(new_n736), .A2(KEYINPUT109), .ZN(new_n737));
  INV_X1    g551(.A(KEYINPUT109), .ZN(new_n738));
  NAND4_X1  g552(.A1(new_n305), .A2(new_n735), .A3(new_n738), .A4(new_n637), .ZN(new_n739));
  NAND2_X1  g553(.A1(new_n737), .A2(new_n739), .ZN(new_n740));
  XNOR2_X1  g554(.A(new_n740), .B(G146), .ZN(G48));
  NAND2_X1  g555(.A1(new_n355), .A2(new_n341), .ZN(new_n742));
  NAND2_X1  g556(.A1(new_n742), .A2(new_n345), .ZN(new_n743));
  XNOR2_X1  g557(.A(new_n349), .B(new_n350), .ZN(new_n744));
  NAND3_X1  g558(.A1(new_n744), .A2(new_n341), .A3(new_n346), .ZN(new_n745));
  AOI21_X1  g559(.A(G902), .B1(new_n743), .B2(new_n745), .ZN(new_n746));
  OAI211_X1 g560(.A(new_n357), .B(new_n369), .C1(new_n746), .C2(new_n366), .ZN(new_n747));
  NOR2_X1   g561(.A1(new_n634), .A2(new_n747), .ZN(new_n748));
  NAND4_X1  g562(.A1(new_n305), .A2(new_n637), .A3(new_n673), .A4(new_n748), .ZN(new_n749));
  XNOR2_X1  g563(.A(KEYINPUT41), .B(G113), .ZN(new_n750));
  XNOR2_X1  g564(.A(new_n749), .B(new_n750), .ZN(G15));
  NAND4_X1  g565(.A1(new_n305), .A2(new_n637), .A3(new_n681), .A4(new_n748), .ZN(new_n752));
  XNOR2_X1  g566(.A(new_n752), .B(G116), .ZN(G18));
  NOR2_X1   g567(.A1(new_n747), .A2(new_n592), .ZN(new_n754));
  NAND3_X1  g568(.A1(new_n754), .A2(new_n688), .A3(new_n527), .ZN(new_n755));
  INV_X1    g569(.A(new_n651), .ZN(new_n756));
  NOR2_X1   g570(.A1(new_n755), .A2(new_n756), .ZN(new_n757));
  NAND3_X1  g571(.A1(new_n305), .A2(new_n757), .A3(new_n637), .ZN(new_n758));
  XNOR2_X1  g572(.A(new_n758), .B(G119), .ZN(G21));
  OAI22_X1  g573(.A1(new_n296), .A2(new_n298), .B1(new_n287), .B2(new_n191), .ZN(new_n760));
  NAND2_X1  g574(.A1(new_n760), .A2(new_n301), .ZN(new_n761));
  AND4_X1   g575(.A1(new_n635), .A2(new_n641), .A3(new_n754), .A4(new_n761), .ZN(new_n762));
  INV_X1    g576(.A(new_n728), .ZN(new_n763));
  AOI21_X1  g577(.A(KEYINPUT110), .B1(new_n651), .B2(new_n763), .ZN(new_n764));
  INV_X1    g578(.A(KEYINPUT110), .ZN(new_n765));
  AOI211_X1 g579(.A(new_n765), .B(new_n728), .C1(new_n648), .C2(new_n650), .ZN(new_n766));
  OAI21_X1  g580(.A(new_n762), .B1(new_n764), .B2(new_n766), .ZN(new_n767));
  XNOR2_X1  g581(.A(new_n767), .B(G122), .ZN(G24));
  NAND4_X1  g582(.A1(new_n641), .A2(new_n688), .A3(new_n733), .A4(new_n761), .ZN(new_n769));
  NOR3_X1   g583(.A1(new_n769), .A2(new_n756), .A3(new_n747), .ZN(new_n770));
  XNOR2_X1  g584(.A(new_n770), .B(new_n373), .ZN(G27));
  NAND2_X1  g585(.A1(new_n367), .A2(new_n369), .ZN(new_n772));
  NOR2_X1   g586(.A1(new_n645), .A2(new_n646), .ZN(new_n773));
  NAND2_X1  g587(.A1(new_n773), .A2(new_n585), .ZN(new_n774));
  NOR2_X1   g588(.A1(new_n772), .A2(new_n774), .ZN(new_n775));
  NAND4_X1  g589(.A1(new_n304), .A2(new_n635), .A3(new_n775), .A4(new_n733), .ZN(new_n776));
  NAND2_X1  g590(.A1(new_n776), .A2(KEYINPUT42), .ZN(new_n777));
  NAND4_X1  g591(.A1(new_n305), .A2(new_n635), .A3(new_n637), .A4(new_n775), .ZN(new_n778));
  INV_X1    g592(.A(new_n733), .ZN(new_n779));
  NOR2_X1   g593(.A1(new_n779), .A2(KEYINPUT42), .ZN(new_n780));
  INV_X1    g594(.A(new_n780), .ZN(new_n781));
  OAI21_X1  g595(.A(new_n777), .B1(new_n778), .B2(new_n781), .ZN(new_n782));
  XNOR2_X1  g596(.A(new_n782), .B(new_n221), .ZN(G33));
  NAND2_X1  g597(.A1(new_n680), .A2(new_n699), .ZN(new_n784));
  OR2_X1    g598(.A1(new_n778), .A2(new_n784), .ZN(new_n785));
  XNOR2_X1  g599(.A(new_n785), .B(G134), .ZN(G36));
  OR3_X1    g600(.A1(new_n669), .A2(KEYINPUT112), .A3(new_n670), .ZN(new_n787));
  OAI21_X1  g601(.A(KEYINPUT112), .B1(new_n669), .B2(new_n670), .ZN(new_n788));
  NAND3_X1  g602(.A1(new_n787), .A2(new_n661), .A3(new_n788), .ZN(new_n789));
  INV_X1    g603(.A(KEYINPUT43), .ZN(new_n790));
  NAND2_X1  g604(.A1(new_n789), .A2(new_n790), .ZN(new_n791));
  INV_X1    g605(.A(KEYINPUT113), .ZN(new_n792));
  NOR2_X1   g606(.A1(new_n671), .A2(new_n790), .ZN(new_n793));
  AOI21_X1  g607(.A(new_n792), .B1(new_n793), .B2(new_n661), .ZN(new_n794));
  NOR4_X1   g608(.A1(new_n449), .A2(new_n671), .A3(KEYINPUT113), .A4(new_n790), .ZN(new_n795));
  OAI21_X1  g609(.A(new_n791), .B1(new_n794), .B2(new_n795), .ZN(new_n796));
  NAND4_X1  g610(.A1(new_n796), .A2(new_n643), .A3(KEYINPUT44), .A4(new_n688), .ZN(new_n797));
  INV_X1    g611(.A(KEYINPUT114), .ZN(new_n798));
  NAND2_X1  g612(.A1(new_n797), .A2(new_n798), .ZN(new_n799));
  INV_X1    g613(.A(new_n774), .ZN(new_n800));
  AOI21_X1  g614(.A(new_n689), .B1(new_n642), .B2(new_n641), .ZN(new_n801));
  NAND4_X1  g615(.A1(new_n801), .A2(KEYINPUT114), .A3(KEYINPUT44), .A4(new_n796), .ZN(new_n802));
  NAND3_X1  g616(.A1(new_n799), .A2(new_n800), .A3(new_n802), .ZN(new_n803));
  NAND2_X1  g617(.A1(new_n803), .A2(KEYINPUT115), .ZN(new_n804));
  NAND2_X1  g618(.A1(new_n361), .A2(new_n364), .ZN(new_n805));
  INV_X1    g619(.A(KEYINPUT45), .ZN(new_n806));
  AOI21_X1  g620(.A(new_n366), .B1(new_n805), .B2(new_n806), .ZN(new_n807));
  NAND3_X1  g621(.A1(new_n361), .A2(KEYINPUT45), .A3(new_n364), .ZN(new_n808));
  AOI22_X1  g622(.A1(new_n807), .A2(new_n808), .B1(G469), .B2(G902), .ZN(new_n809));
  AND2_X1   g623(.A1(new_n809), .A2(KEYINPUT46), .ZN(new_n810));
  OAI21_X1  g624(.A(new_n357), .B1(new_n809), .B2(KEYINPUT46), .ZN(new_n811));
  OAI211_X1 g625(.A(new_n369), .B(new_n708), .C1(new_n810), .C2(new_n811), .ZN(new_n812));
  INV_X1    g626(.A(KEYINPUT111), .ZN(new_n813));
  XNOR2_X1  g627(.A(new_n812), .B(new_n813), .ZN(new_n814));
  AND2_X1   g628(.A1(new_n801), .A2(new_n796), .ZN(new_n815));
  OR2_X1    g629(.A1(new_n815), .A2(KEYINPUT44), .ZN(new_n816));
  INV_X1    g630(.A(KEYINPUT115), .ZN(new_n817));
  NAND4_X1  g631(.A1(new_n799), .A2(new_n802), .A3(new_n817), .A4(new_n800), .ZN(new_n818));
  NAND4_X1  g632(.A1(new_n804), .A2(new_n814), .A3(new_n816), .A4(new_n818), .ZN(new_n819));
  XNOR2_X1  g633(.A(new_n819), .B(G137), .ZN(G39));
  OAI21_X1  g634(.A(new_n369), .B1(new_n810), .B2(new_n811), .ZN(new_n821));
  INV_X1    g635(.A(KEYINPUT47), .ZN(new_n822));
  NAND2_X1  g636(.A1(new_n821), .A2(new_n822), .ZN(new_n823));
  OAI211_X1 g637(.A(KEYINPUT47), .B(new_n369), .C1(new_n810), .C2(new_n811), .ZN(new_n824));
  NAND2_X1  g638(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  NAND3_X1  g639(.A1(new_n800), .A2(new_n634), .A3(new_n733), .ZN(new_n826));
  AOI21_X1  g640(.A(new_n826), .B1(new_n305), .B2(new_n637), .ZN(new_n827));
  NAND2_X1  g641(.A1(new_n825), .A2(new_n827), .ZN(new_n828));
  XNOR2_X1  g642(.A(new_n828), .B(G140), .ZN(G42));
  NAND2_X1  g643(.A1(new_n369), .A2(new_n585), .ZN(new_n830));
  NOR4_X1   g644(.A1(new_n634), .A2(new_n449), .A3(new_n671), .A4(new_n830), .ZN(new_n831));
  AND2_X1   g645(.A1(new_n721), .A2(new_n831), .ZN(new_n832));
  INV_X1    g646(.A(new_n723), .ZN(new_n833));
  NOR2_X1   g647(.A1(new_n746), .A2(new_n366), .ZN(new_n834));
  AOI21_X1  g648(.A(new_n834), .B1(new_n746), .B2(new_n307), .ZN(new_n835));
  XOR2_X1   g649(.A(new_n835), .B(KEYINPUT116), .Z(new_n836));
  INV_X1    g650(.A(new_n836), .ZN(new_n837));
  AOI21_X1  g651(.A(new_n833), .B1(new_n837), .B2(KEYINPUT49), .ZN(new_n838));
  OAI211_X1 g652(.A(new_n832), .B(new_n838), .C1(KEYINPUT49), .C2(new_n837), .ZN(new_n839));
  NAND4_X1  g653(.A1(new_n749), .A2(new_n752), .A3(new_n758), .A4(new_n767), .ZN(new_n840));
  INV_X1    g654(.A(KEYINPUT117), .ZN(new_n841));
  XNOR2_X1  g655(.A(new_n840), .B(new_n841), .ZN(new_n842));
  NOR2_X1   g656(.A1(new_n514), .A2(new_n516), .ZN(new_n843));
  NAND3_X1  g657(.A1(new_n679), .A2(new_n843), .A3(new_n699), .ZN(new_n844));
  NOR2_X1   g658(.A1(new_n689), .A2(new_n844), .ZN(new_n845));
  NAND4_X1  g659(.A1(new_n305), .A2(new_n637), .A3(new_n775), .A4(new_n845), .ZN(new_n846));
  INV_X1    g660(.A(new_n775), .ZN(new_n847));
  OAI221_X1 g661(.A(new_n846), .B1(new_n769), .B2(new_n847), .C1(new_n778), .C2(new_n784), .ZN(new_n848));
  NOR2_X1   g662(.A1(new_n449), .A2(new_n843), .ZN(new_n849));
  NOR2_X1   g663(.A1(new_n672), .A2(new_n849), .ZN(new_n850));
  NOR3_X1   g664(.A1(new_n850), .A2(new_n772), .A3(new_n594), .ZN(new_n851));
  AOI22_X1  g665(.A1(new_n596), .A2(new_n690), .B1(new_n644), .B2(new_n851), .ZN(new_n852));
  NAND2_X1  g666(.A1(new_n852), .A2(new_n638), .ZN(new_n853));
  NOR3_X1   g667(.A1(new_n848), .A2(new_n782), .A3(new_n853), .ZN(new_n854));
  AND2_X1   g668(.A1(new_n842), .A2(new_n854), .ZN(new_n855));
  AOI21_X1  g669(.A(new_n770), .B1(new_n704), .B2(new_n705), .ZN(new_n856));
  NOR2_X1   g670(.A1(new_n764), .A2(new_n766), .ZN(new_n857));
  NOR3_X1   g671(.A1(new_n772), .A2(new_n688), .A3(new_n698), .ZN(new_n858));
  NAND2_X1  g672(.A1(new_n858), .A2(new_n720), .ZN(new_n859));
  NOR2_X1   g673(.A1(new_n857), .A2(new_n859), .ZN(new_n860));
  AOI21_X1  g674(.A(new_n860), .B1(new_n737), .B2(new_n739), .ZN(new_n861));
  NAND2_X1  g675(.A1(new_n856), .A2(new_n861), .ZN(new_n862));
  INV_X1    g676(.A(KEYINPUT52), .ZN(new_n863));
  NAND2_X1  g677(.A1(new_n862), .A2(new_n863), .ZN(new_n864));
  OAI21_X1  g678(.A(KEYINPUT52), .B1(new_n857), .B2(new_n859), .ZN(new_n865));
  AOI21_X1  g679(.A(new_n865), .B1(new_n737), .B2(new_n739), .ZN(new_n866));
  AND3_X1   g680(.A1(new_n866), .A2(new_n856), .A3(KEYINPUT118), .ZN(new_n867));
  AOI21_X1  g681(.A(KEYINPUT118), .B1(new_n866), .B2(new_n856), .ZN(new_n868));
  OAI21_X1  g682(.A(new_n864), .B1(new_n867), .B2(new_n868), .ZN(new_n869));
  INV_X1    g683(.A(KEYINPUT53), .ZN(new_n870));
  NAND3_X1  g684(.A1(new_n855), .A2(new_n869), .A3(new_n870), .ZN(new_n871));
  NAND2_X1  g685(.A1(new_n866), .A2(new_n856), .ZN(new_n872));
  INV_X1    g686(.A(new_n872), .ZN(new_n873));
  AOI21_X1  g687(.A(KEYINPUT52), .B1(new_n856), .B2(new_n861), .ZN(new_n874));
  OAI211_X1 g688(.A(new_n842), .B(new_n854), .C1(new_n873), .C2(new_n874), .ZN(new_n875));
  NAND2_X1  g689(.A1(new_n875), .A2(KEYINPUT53), .ZN(new_n876));
  NAND3_X1  g690(.A1(new_n871), .A2(new_n876), .A3(KEYINPUT54), .ZN(new_n877));
  NAND2_X1  g691(.A1(new_n875), .A2(new_n870), .ZN(new_n878));
  NOR2_X1   g692(.A1(new_n840), .A2(new_n870), .ZN(new_n879));
  AND2_X1   g693(.A1(new_n854), .A2(new_n879), .ZN(new_n880));
  NAND2_X1  g694(.A1(new_n869), .A2(new_n880), .ZN(new_n881));
  XOR2_X1   g695(.A(KEYINPUT119), .B(KEYINPUT54), .Z(new_n882));
  NAND3_X1  g696(.A1(new_n878), .A2(new_n881), .A3(new_n882), .ZN(new_n883));
  NOR3_X1   g697(.A1(new_n774), .A2(new_n747), .A3(new_n588), .ZN(new_n884));
  AND2_X1   g698(.A1(new_n796), .A2(new_n884), .ZN(new_n885));
  AND2_X1   g699(.A1(new_n641), .A2(new_n761), .ZN(new_n886));
  NAND3_X1  g700(.A1(new_n885), .A2(new_n688), .A3(new_n886), .ZN(new_n887));
  AND2_X1   g701(.A1(new_n884), .A2(new_n635), .ZN(new_n888));
  NAND2_X1  g702(.A1(new_n888), .A2(new_n721), .ZN(new_n889));
  NAND2_X1  g703(.A1(new_n661), .A2(new_n671), .ZN(new_n890));
  OAI21_X1  g704(.A(new_n887), .B1(new_n889), .B2(new_n890), .ZN(new_n891));
  AND4_X1   g705(.A1(new_n635), .A2(new_n886), .A3(new_n589), .A4(new_n796), .ZN(new_n892));
  NOR3_X1   g706(.A1(new_n833), .A2(new_n585), .A3(new_n747), .ZN(new_n893));
  AND2_X1   g707(.A1(new_n892), .A2(new_n893), .ZN(new_n894));
  OR2_X1    g708(.A1(new_n894), .A2(KEYINPUT50), .ZN(new_n895));
  NAND2_X1  g709(.A1(new_n894), .A2(KEYINPUT50), .ZN(new_n896));
  AOI21_X1  g710(.A(new_n891), .B1(new_n895), .B2(new_n896), .ZN(new_n897));
  AOI21_X1  g711(.A(new_n369), .B1(new_n836), .B2(KEYINPUT120), .ZN(new_n898));
  OAI21_X1  g712(.A(new_n898), .B1(KEYINPUT120), .B2(new_n836), .ZN(new_n899));
  NAND3_X1  g713(.A1(new_n899), .A2(new_n823), .A3(new_n824), .ZN(new_n900));
  NAND3_X1  g714(.A1(new_n900), .A2(new_n800), .A3(new_n892), .ZN(new_n901));
  NAND3_X1  g715(.A1(new_n897), .A2(KEYINPUT51), .A3(new_n901), .ZN(new_n902));
  AOI21_X1  g716(.A(KEYINPUT51), .B1(new_n897), .B2(new_n901), .ZN(new_n903));
  AND2_X1   g717(.A1(new_n304), .A2(new_n635), .ZN(new_n904));
  NAND2_X1  g718(.A1(new_n885), .A2(new_n904), .ZN(new_n905));
  XOR2_X1   g719(.A(new_n905), .B(KEYINPUT48), .Z(new_n906));
  NAND4_X1  g720(.A1(new_n892), .A2(new_n369), .A3(new_n651), .A4(new_n835), .ZN(new_n907));
  NAND3_X1  g721(.A1(new_n888), .A2(new_n721), .A3(new_n672), .ZN(new_n908));
  NAND3_X1  g722(.A1(new_n907), .A2(new_n586), .A3(new_n908), .ZN(new_n909));
  NOR3_X1   g723(.A1(new_n903), .A2(new_n906), .A3(new_n909), .ZN(new_n910));
  AND4_X1   g724(.A1(new_n877), .A2(new_n883), .A3(new_n902), .A4(new_n910), .ZN(new_n911));
  NOR2_X1   g725(.A1(G952), .A2(G953), .ZN(new_n912));
  XOR2_X1   g726(.A(new_n912), .B(KEYINPUT121), .Z(new_n913));
  OAI21_X1  g727(.A(new_n839), .B1(new_n911), .B2(new_n913), .ZN(G75));
  NOR2_X1   g728(.A1(new_n343), .A2(G952), .ZN(new_n915));
  INV_X1    g729(.A(new_n915), .ZN(new_n916));
  AOI21_X1  g730(.A(new_n306), .B1(new_n878), .B2(new_n881), .ZN(new_n917));
  AOI21_X1  g731(.A(KEYINPUT56), .B1(new_n917), .B2(G210), .ZN(new_n918));
  AND2_X1   g732(.A1(new_n548), .A2(new_n551), .ZN(new_n919));
  XOR2_X1   g733(.A(new_n919), .B(new_n563), .Z(new_n920));
  XNOR2_X1  g734(.A(new_n920), .B(KEYINPUT55), .ZN(new_n921));
  OAI21_X1  g735(.A(new_n916), .B1(new_n918), .B2(new_n921), .ZN(new_n922));
  INV_X1    g736(.A(KEYINPUT122), .ZN(new_n923));
  AOI22_X1  g737(.A1(new_n870), .A2(new_n875), .B1(new_n869), .B2(new_n880), .ZN(new_n924));
  OAI21_X1  g738(.A(new_n923), .B1(new_n924), .B2(new_n306), .ZN(new_n925));
  NAND2_X1  g739(.A1(new_n864), .A2(new_n872), .ZN(new_n926));
  AOI21_X1  g740(.A(KEYINPUT53), .B1(new_n855), .B2(new_n926), .ZN(new_n927));
  NAND2_X1  g741(.A1(new_n854), .A2(new_n879), .ZN(new_n928));
  INV_X1    g742(.A(KEYINPUT118), .ZN(new_n929));
  NAND2_X1  g743(.A1(new_n872), .A2(new_n929), .ZN(new_n930));
  NAND3_X1  g744(.A1(new_n866), .A2(new_n856), .A3(KEYINPUT118), .ZN(new_n931));
  NAND2_X1  g745(.A1(new_n930), .A2(new_n931), .ZN(new_n932));
  AOI21_X1  g746(.A(new_n928), .B1(new_n932), .B2(new_n864), .ZN(new_n933));
  OAI211_X1 g747(.A(KEYINPUT122), .B(G902), .C1(new_n927), .C2(new_n933), .ZN(new_n934));
  NAND3_X1  g748(.A1(new_n925), .A2(new_n934), .A3(new_n581), .ZN(new_n935));
  INV_X1    g749(.A(KEYINPUT56), .ZN(new_n936));
  AND2_X1   g750(.A1(new_n921), .A2(new_n936), .ZN(new_n937));
  AOI21_X1  g751(.A(new_n922), .B1(new_n935), .B2(new_n937), .ZN(G51));
  NAND2_X1  g752(.A1(G469), .A2(G902), .ZN(new_n939));
  XNOR2_X1  g753(.A(new_n939), .B(KEYINPUT123), .ZN(new_n940));
  XNOR2_X1  g754(.A(new_n940), .B(KEYINPUT57), .ZN(new_n941));
  NOR2_X1   g755(.A1(new_n924), .A2(new_n882), .ZN(new_n942));
  INV_X1    g756(.A(new_n883), .ZN(new_n943));
  OAI21_X1  g757(.A(new_n941), .B1(new_n942), .B2(new_n943), .ZN(new_n944));
  NAND2_X1  g758(.A1(new_n743), .A2(new_n745), .ZN(new_n945));
  NAND2_X1  g759(.A1(new_n944), .A2(new_n945), .ZN(new_n946));
  NAND4_X1  g760(.A1(new_n925), .A2(new_n934), .A3(new_n808), .A4(new_n807), .ZN(new_n947));
  AOI21_X1  g761(.A(new_n915), .B1(new_n946), .B2(new_n947), .ZN(G54));
  AND2_X1   g762(.A1(KEYINPUT58), .A2(G475), .ZN(new_n949));
  NAND3_X1  g763(.A1(new_n925), .A2(new_n934), .A3(new_n949), .ZN(new_n950));
  NAND2_X1  g764(.A1(new_n950), .A2(new_n657), .ZN(new_n951));
  NAND4_X1  g765(.A1(new_n925), .A2(new_n934), .A3(new_n443), .A4(new_n949), .ZN(new_n952));
  AND3_X1   g766(.A1(new_n951), .A2(new_n916), .A3(new_n952), .ZN(G60));
  NAND2_X1  g767(.A1(G478), .A2(G902), .ZN(new_n954));
  XOR2_X1   g768(.A(new_n954), .B(KEYINPUT59), .Z(new_n955));
  AOI21_X1  g769(.A(new_n955), .B1(new_n877), .B2(new_n883), .ZN(new_n956));
  NAND2_X1  g770(.A1(new_n664), .A2(new_n668), .ZN(new_n957));
  OAI21_X1  g771(.A(new_n916), .B1(new_n956), .B2(new_n957), .ZN(new_n958));
  AOI21_X1  g772(.A(new_n955), .B1(new_n664), .B2(new_n668), .ZN(new_n959));
  OAI21_X1  g773(.A(new_n959), .B1(new_n942), .B2(new_n943), .ZN(new_n960));
  NAND2_X1  g774(.A1(new_n960), .A2(KEYINPUT124), .ZN(new_n961));
  INV_X1    g775(.A(KEYINPUT124), .ZN(new_n962));
  OAI211_X1 g776(.A(new_n962), .B(new_n959), .C1(new_n942), .C2(new_n943), .ZN(new_n963));
  AOI21_X1  g777(.A(new_n958), .B1(new_n961), .B2(new_n963), .ZN(G63));
  INV_X1    g778(.A(KEYINPUT125), .ZN(new_n965));
  INV_X1    g779(.A(KEYINPUT61), .ZN(new_n966));
  AOI21_X1  g780(.A(new_n915), .B1(KEYINPUT125), .B2(new_n966), .ZN(new_n967));
  NAND2_X1  g781(.A1(G217), .A2(G902), .ZN(new_n968));
  XNOR2_X1  g782(.A(new_n968), .B(KEYINPUT60), .ZN(new_n969));
  AOI21_X1  g783(.A(new_n969), .B1(new_n878), .B2(new_n881), .ZN(new_n970));
  OAI21_X1  g784(.A(new_n967), .B1(new_n970), .B2(new_n622), .ZN(new_n971));
  XOR2_X1   g785(.A(new_n611), .B(new_n685), .Z(new_n972));
  NOR3_X1   g786(.A1(new_n924), .A2(new_n972), .A3(new_n969), .ZN(new_n973));
  OAI211_X1 g787(.A(new_n965), .B(KEYINPUT61), .C1(new_n971), .C2(new_n973), .ZN(new_n974));
  OR2_X1    g788(.A1(new_n970), .A2(new_n622), .ZN(new_n975));
  NAND2_X1  g789(.A1(new_n965), .A2(KEYINPUT61), .ZN(new_n976));
  NAND2_X1  g790(.A1(new_n970), .A2(new_n686), .ZN(new_n977));
  NAND4_X1  g791(.A1(new_n975), .A2(new_n976), .A3(new_n977), .A4(new_n967), .ZN(new_n978));
  AND2_X1   g792(.A1(new_n974), .A2(new_n978), .ZN(G66));
  INV_X1    g793(.A(new_n591), .ZN(new_n980));
  AOI21_X1  g794(.A(new_n343), .B1(new_n980), .B2(G224), .ZN(new_n981));
  NAND3_X1  g795(.A1(new_n842), .A2(new_n638), .A3(new_n852), .ZN(new_n982));
  AOI21_X1  g796(.A(new_n981), .B1(new_n982), .B2(new_n343), .ZN(new_n983));
  INV_X1    g797(.A(G898), .ZN(new_n984));
  AOI21_X1  g798(.A(new_n919), .B1(new_n984), .B2(G953), .ZN(new_n985));
  XNOR2_X1  g799(.A(new_n983), .B(new_n985), .ZN(G69));
  AOI21_X1  g800(.A(new_n343), .B1(G227), .B2(G900), .ZN(new_n987));
  INV_X1    g801(.A(KEYINPUT126), .ZN(new_n988));
  NAND2_X1  g802(.A1(new_n305), .A2(new_n637), .ZN(new_n989));
  NOR2_X1   g803(.A1(new_n989), .A2(new_n634), .ZN(new_n990));
  NOR3_X1   g804(.A1(new_n709), .A2(new_n774), .A3(new_n850), .ZN(new_n991));
  AOI22_X1  g805(.A1(new_n825), .A2(new_n827), .B1(new_n990), .B2(new_n991), .ZN(new_n992));
  AND2_X1   g806(.A1(new_n819), .A2(new_n992), .ZN(new_n993));
  NAND3_X1  g807(.A1(new_n856), .A2(new_n731), .A3(new_n740), .ZN(new_n994));
  OR2_X1    g808(.A1(new_n994), .A2(KEYINPUT62), .ZN(new_n995));
  NAND2_X1  g809(.A1(new_n994), .A2(KEYINPUT62), .ZN(new_n996));
  NAND3_X1  g810(.A1(new_n993), .A2(new_n995), .A3(new_n996), .ZN(new_n997));
  NAND2_X1  g811(.A1(new_n997), .A2(new_n343), .ZN(new_n998));
  INV_X1    g812(.A(new_n266), .ZN(new_n999));
  OAI21_X1  g813(.A(new_n999), .B1(new_n270), .B2(new_n271), .ZN(new_n1000));
  OR2_X1    g814(.A1(new_n433), .A2(new_n434), .ZN(new_n1001));
  XNOR2_X1  g815(.A(new_n1000), .B(new_n1001), .ZN(new_n1002));
  AOI21_X1  g816(.A(new_n988), .B1(new_n998), .B2(new_n1002), .ZN(new_n1003));
  INV_X1    g817(.A(new_n1002), .ZN(new_n1004));
  AOI211_X1 g818(.A(KEYINPUT126), .B(new_n1004), .C1(new_n997), .C2(new_n343), .ZN(new_n1005));
  NOR2_X1   g819(.A1(new_n1003), .A2(new_n1005), .ZN(new_n1006));
  XNOR2_X1  g820(.A(new_n812), .B(KEYINPUT111), .ZN(new_n1007));
  OAI21_X1  g821(.A(new_n904), .B1(new_n764), .B2(new_n766), .ZN(new_n1008));
  OAI211_X1 g822(.A(new_n856), .B(new_n740), .C1(new_n1007), .C2(new_n1008), .ZN(new_n1009));
  OR2_X1    g823(.A1(new_n778), .A2(new_n781), .ZN(new_n1010));
  NAND4_X1  g824(.A1(new_n828), .A2(new_n1010), .A3(new_n777), .A4(new_n785), .ZN(new_n1011));
  NOR2_X1   g825(.A1(new_n1009), .A2(new_n1011), .ZN(new_n1012));
  AOI21_X1  g826(.A(G953), .B1(new_n1012), .B2(new_n819), .ZN(new_n1013));
  NOR2_X1   g827(.A1(new_n343), .A2(G900), .ZN(new_n1014));
  OAI21_X1  g828(.A(KEYINPUT127), .B1(new_n1013), .B2(new_n1014), .ZN(new_n1015));
  INV_X1    g829(.A(KEYINPUT127), .ZN(new_n1016));
  INV_X1    g830(.A(new_n1014), .ZN(new_n1017));
  INV_X1    g831(.A(new_n819), .ZN(new_n1018));
  NOR3_X1   g832(.A1(new_n1018), .A2(new_n1009), .A3(new_n1011), .ZN(new_n1019));
  OAI211_X1 g833(.A(new_n1016), .B(new_n1017), .C1(new_n1019), .C2(G953), .ZN(new_n1020));
  NAND3_X1  g834(.A1(new_n1015), .A2(new_n1020), .A3(new_n1004), .ZN(new_n1021));
  AOI21_X1  g835(.A(new_n987), .B1(new_n1006), .B2(new_n1021), .ZN(new_n1022));
  NAND2_X1  g836(.A1(new_n998), .A2(new_n1002), .ZN(new_n1023));
  NAND2_X1  g837(.A1(new_n1023), .A2(KEYINPUT126), .ZN(new_n1024));
  NAND3_X1  g838(.A1(new_n998), .A2(new_n988), .A3(new_n1002), .ZN(new_n1025));
  AND4_X1   g839(.A1(new_n1021), .A2(new_n1024), .A3(new_n1025), .A4(new_n987), .ZN(new_n1026));
  NOR2_X1   g840(.A1(new_n1022), .A2(new_n1026), .ZN(G72));
  NAND2_X1  g841(.A1(G472), .A2(G902), .ZN(new_n1028));
  XOR2_X1   g842(.A(new_n1028), .B(KEYINPUT63), .Z(new_n1029));
  INV_X1    g843(.A(new_n1019), .ZN(new_n1030));
  OAI21_X1  g844(.A(new_n1029), .B1(new_n1030), .B2(new_n982), .ZN(new_n1031));
  NAND2_X1  g845(.A1(new_n1031), .A2(new_n276), .ZN(new_n1032));
  INV_X1    g846(.A(new_n276), .ZN(new_n1033));
  NAND2_X1  g847(.A1(new_n1033), .A2(new_n1029), .ZN(new_n1034));
  AOI21_X1  g848(.A(new_n277), .B1(new_n293), .B2(new_n251), .ZN(new_n1035));
  NOR2_X1   g849(.A1(new_n1034), .A2(new_n1035), .ZN(new_n1036));
  NAND3_X1  g850(.A1(new_n871), .A2(new_n876), .A3(new_n1036), .ZN(new_n1037));
  NAND3_X1  g851(.A1(new_n1032), .A2(new_n916), .A3(new_n1037), .ZN(new_n1038));
  OAI21_X1  g852(.A(new_n1029), .B1(new_n997), .B2(new_n982), .ZN(new_n1039));
  AOI21_X1  g853(.A(new_n1038), .B1(new_n1039), .B2(new_n1035), .ZN(G57));
endmodule


