

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301,
         n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312,
         n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323,
         n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334,
         n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
         n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
         n588;

  XOR2_X1 U323 ( .A(KEYINPUT85), .B(G99GAT), .Z(n291) );
  XOR2_X1 U324 ( .A(n375), .B(n374), .Z(n292) );
  INV_X1 U325 ( .A(KEYINPUT65), .ZN(n379) );
  XNOR2_X1 U326 ( .A(n380), .B(n379), .ZN(n381) );
  NAND2_X1 U327 ( .A1(n555), .A2(n552), .ZN(n442) );
  XNOR2_X1 U328 ( .A(n382), .B(n381), .ZN(n383) );
  XOR2_X1 U329 ( .A(KEYINPUT38), .B(n468), .Z(n476) );
  XNOR2_X1 U330 ( .A(G1GAT), .B(KEYINPUT34), .ZN(n293) );
  XNOR2_X1 U331 ( .A(n293), .B(KEYINPUT101), .ZN(n294) );
  XOR2_X1 U332 ( .A(KEYINPUT100), .B(n294), .Z(n455) );
  XOR2_X1 U333 ( .A(KEYINPUT71), .B(KEYINPUT30), .Z(n296) );
  XNOR2_X1 U334 ( .A(KEYINPUT73), .B(KEYINPUT68), .ZN(n295) );
  XNOR2_X1 U335 ( .A(n296), .B(n295), .ZN(n314) );
  XOR2_X1 U336 ( .A(G22GAT), .B(G113GAT), .Z(n298) );
  XNOR2_X1 U337 ( .A(G50GAT), .B(G36GAT), .ZN(n297) );
  XNOR2_X1 U338 ( .A(n298), .B(n297), .ZN(n302) );
  XOR2_X1 U339 ( .A(KEYINPUT74), .B(KEYINPUT72), .Z(n300) );
  XNOR2_X1 U340 ( .A(G197GAT), .B(G141GAT), .ZN(n299) );
  XNOR2_X1 U341 ( .A(n300), .B(n299), .ZN(n301) );
  XOR2_X1 U342 ( .A(n302), .B(n301), .Z(n307) );
  XOR2_X1 U343 ( .A(KEYINPUT69), .B(KEYINPUT29), .Z(n304) );
  NAND2_X1 U344 ( .A1(G229GAT), .A2(G233GAT), .ZN(n303) );
  XNOR2_X1 U345 ( .A(n304), .B(n303), .ZN(n305) );
  XNOR2_X1 U346 ( .A(KEYINPUT70), .B(n305), .ZN(n306) );
  XNOR2_X1 U347 ( .A(n307), .B(n306), .ZN(n308) );
  XOR2_X1 U348 ( .A(G169GAT), .B(G8GAT), .Z(n418) );
  XOR2_X1 U349 ( .A(n308), .B(n418), .Z(n312) );
  XOR2_X1 U350 ( .A(G29GAT), .B(G43GAT), .Z(n310) );
  XNOR2_X1 U351 ( .A(KEYINPUT8), .B(KEYINPUT7), .ZN(n309) );
  XNOR2_X1 U352 ( .A(n310), .B(n309), .ZN(n347) );
  XOR2_X1 U353 ( .A(G15GAT), .B(G1GAT), .Z(n353) );
  XNOR2_X1 U354 ( .A(n347), .B(n353), .ZN(n311) );
  XNOR2_X1 U355 ( .A(n312), .B(n311), .ZN(n313) );
  XOR2_X2 U356 ( .A(n314), .B(n313), .Z(n572) );
  XOR2_X1 U357 ( .A(G120GAT), .B(G71GAT), .Z(n375) );
  XOR2_X1 U358 ( .A(G57GAT), .B(KEYINPUT13), .Z(n352) );
  XNOR2_X1 U359 ( .A(n375), .B(n352), .ZN(n329) );
  XOR2_X1 U360 ( .A(G92GAT), .B(KEYINPUT75), .Z(n316) );
  XNOR2_X1 U361 ( .A(G99GAT), .B(G85GAT), .ZN(n315) );
  XNOR2_X1 U362 ( .A(n316), .B(n315), .ZN(n346) );
  XOR2_X1 U363 ( .A(n346), .B(KEYINPUT31), .Z(n318) );
  NAND2_X1 U364 ( .A1(G230GAT), .A2(G233GAT), .ZN(n317) );
  XNOR2_X1 U365 ( .A(n318), .B(n317), .ZN(n322) );
  XOR2_X1 U366 ( .A(KEYINPUT76), .B(KEYINPUT32), .Z(n320) );
  XNOR2_X1 U367 ( .A(KEYINPUT77), .B(KEYINPUT33), .ZN(n319) );
  XNOR2_X1 U368 ( .A(n320), .B(n319), .ZN(n321) );
  XOR2_X1 U369 ( .A(n322), .B(n321), .Z(n327) );
  XNOR2_X1 U370 ( .A(G106GAT), .B(G78GAT), .ZN(n323) );
  XNOR2_X1 U371 ( .A(n323), .B(G148GAT), .ZN(n427) );
  XOR2_X1 U372 ( .A(KEYINPUT78), .B(G64GAT), .Z(n325) );
  XNOR2_X1 U373 ( .A(G176GAT), .B(G204GAT), .ZN(n324) );
  XNOR2_X1 U374 ( .A(n325), .B(n324), .ZN(n405) );
  XNOR2_X1 U375 ( .A(n427), .B(n405), .ZN(n326) );
  XNOR2_X1 U376 ( .A(n327), .B(n326), .ZN(n328) );
  XNOR2_X1 U377 ( .A(n329), .B(n328), .ZN(n577) );
  NAND2_X1 U378 ( .A1(n572), .A2(n577), .ZN(n467) );
  XOR2_X1 U379 ( .A(KEYINPUT80), .B(KEYINPUT10), .Z(n331) );
  XNOR2_X1 U380 ( .A(G106GAT), .B(KEYINPUT79), .ZN(n330) );
  XNOR2_X1 U381 ( .A(n331), .B(n330), .ZN(n339) );
  XOR2_X1 U382 ( .A(G36GAT), .B(G190GAT), .Z(n406) );
  INV_X1 U383 ( .A(n406), .ZN(n332) );
  NAND2_X1 U384 ( .A1(KEYINPUT9), .A2(n332), .ZN(n335) );
  INV_X1 U385 ( .A(KEYINPUT9), .ZN(n333) );
  NAND2_X1 U386 ( .A1(n333), .A2(n406), .ZN(n334) );
  NAND2_X1 U387 ( .A1(n335), .A2(n334), .ZN(n337) );
  XOR2_X1 U388 ( .A(G50GAT), .B(G162GAT), .Z(n437) );
  XNOR2_X1 U389 ( .A(G218GAT), .B(n437), .ZN(n336) );
  XNOR2_X1 U390 ( .A(n337), .B(n336), .ZN(n338) );
  XOR2_X1 U391 ( .A(n339), .B(n338), .Z(n341) );
  NAND2_X1 U392 ( .A1(G232GAT), .A2(G233GAT), .ZN(n340) );
  XNOR2_X1 U393 ( .A(n341), .B(n340), .ZN(n345) );
  XOR2_X1 U394 ( .A(KEYINPUT67), .B(KEYINPUT11), .Z(n343) );
  XNOR2_X1 U395 ( .A(G134GAT), .B(KEYINPUT66), .ZN(n342) );
  XNOR2_X1 U396 ( .A(n343), .B(n342), .ZN(n344) );
  XOR2_X1 U397 ( .A(n345), .B(n344), .Z(n349) );
  XNOR2_X1 U398 ( .A(n347), .B(n346), .ZN(n348) );
  XNOR2_X1 U399 ( .A(n349), .B(n348), .ZN(n566) );
  XOR2_X1 U400 ( .A(G78GAT), .B(G211GAT), .Z(n351) );
  XNOR2_X1 U401 ( .A(G127GAT), .B(G71GAT), .ZN(n350) );
  XNOR2_X1 U402 ( .A(n351), .B(n350), .ZN(n366) );
  XOR2_X1 U403 ( .A(G183GAT), .B(KEYINPUT81), .Z(n413) );
  XOR2_X1 U404 ( .A(n413), .B(n352), .Z(n355) );
  XOR2_X1 U405 ( .A(G22GAT), .B(G155GAT), .Z(n436) );
  XNOR2_X1 U406 ( .A(n353), .B(n436), .ZN(n354) );
  XNOR2_X1 U407 ( .A(n355), .B(n354), .ZN(n359) );
  XOR2_X1 U408 ( .A(G64GAT), .B(KEYINPUT14), .Z(n357) );
  NAND2_X1 U409 ( .A1(G231GAT), .A2(G233GAT), .ZN(n356) );
  XNOR2_X1 U410 ( .A(n357), .B(n356), .ZN(n358) );
  XOR2_X1 U411 ( .A(n359), .B(n358), .Z(n364) );
  XOR2_X1 U412 ( .A(KEYINPUT15), .B(KEYINPUT83), .Z(n361) );
  XNOR2_X1 U413 ( .A(KEYINPUT12), .B(KEYINPUT82), .ZN(n360) );
  XNOR2_X1 U414 ( .A(n361), .B(n360), .ZN(n362) );
  XNOR2_X1 U415 ( .A(G8GAT), .B(n362), .ZN(n363) );
  XNOR2_X1 U416 ( .A(n364), .B(n363), .ZN(n365) );
  XNOR2_X1 U417 ( .A(n366), .B(n365), .ZN(n582) );
  INV_X1 U418 ( .A(n582), .ZN(n510) );
  NOR2_X1 U419 ( .A1(n566), .A2(n510), .ZN(n367) );
  XNOR2_X1 U420 ( .A(n367), .B(KEYINPUT16), .ZN(n453) );
  XOR2_X1 U421 ( .A(KEYINPUT0), .B(G134GAT), .Z(n369) );
  XNOR2_X1 U422 ( .A(KEYINPUT84), .B(G127GAT), .ZN(n368) );
  XNOR2_X1 U423 ( .A(n369), .B(n368), .ZN(n370) );
  XOR2_X1 U424 ( .A(G113GAT), .B(n370), .Z(n404) );
  XOR2_X1 U425 ( .A(G176GAT), .B(G183GAT), .Z(n372) );
  XNOR2_X1 U426 ( .A(G169GAT), .B(G15GAT), .ZN(n371) );
  XNOR2_X1 U427 ( .A(n372), .B(n371), .ZN(n384) );
  XNOR2_X1 U428 ( .A(G43GAT), .B(G190GAT), .ZN(n373) );
  XNOR2_X1 U429 ( .A(n291), .B(n373), .ZN(n374) );
  NAND2_X1 U430 ( .A1(G227GAT), .A2(G233GAT), .ZN(n376) );
  XNOR2_X1 U431 ( .A(n292), .B(n376), .ZN(n382) );
  XOR2_X1 U432 ( .A(KEYINPUT19), .B(KEYINPUT86), .Z(n378) );
  XNOR2_X1 U433 ( .A(KEYINPUT17), .B(KEYINPUT18), .ZN(n377) );
  XNOR2_X1 U434 ( .A(n378), .B(n377), .ZN(n410) );
  XNOR2_X1 U435 ( .A(n410), .B(KEYINPUT20), .ZN(n380) );
  XOR2_X1 U436 ( .A(n384), .B(n383), .Z(n385) );
  XNOR2_X1 U437 ( .A(n404), .B(n385), .ZN(n519) );
  INV_X1 U438 ( .A(n519), .ZN(n555) );
  XNOR2_X1 U439 ( .A(G141GAT), .B(KEYINPUT2), .ZN(n386) );
  XNOR2_X1 U440 ( .A(n386), .B(KEYINPUT3), .ZN(n434) );
  XOR2_X1 U441 ( .A(G85GAT), .B(n434), .Z(n388) );
  XNOR2_X1 U442 ( .A(G120GAT), .B(G162GAT), .ZN(n387) );
  XNOR2_X1 U443 ( .A(n388), .B(n387), .ZN(n389) );
  XNOR2_X1 U444 ( .A(G29GAT), .B(n389), .ZN(n402) );
  XOR2_X1 U445 ( .A(G57GAT), .B(G155GAT), .Z(n391) );
  XNOR2_X1 U446 ( .A(G1GAT), .B(G148GAT), .ZN(n390) );
  XNOR2_X1 U447 ( .A(n391), .B(n390), .ZN(n395) );
  XOR2_X1 U448 ( .A(KEYINPUT1), .B(KEYINPUT6), .Z(n393) );
  XNOR2_X1 U449 ( .A(KEYINPUT5), .B(KEYINPUT93), .ZN(n392) );
  XNOR2_X1 U450 ( .A(n393), .B(n392), .ZN(n394) );
  XOR2_X1 U451 ( .A(n395), .B(n394), .Z(n400) );
  XOR2_X1 U452 ( .A(KEYINPUT94), .B(KEYINPUT95), .Z(n397) );
  NAND2_X1 U453 ( .A1(G225GAT), .A2(G233GAT), .ZN(n396) );
  XNOR2_X1 U454 ( .A(n397), .B(n396), .ZN(n398) );
  XNOR2_X1 U455 ( .A(KEYINPUT4), .B(n398), .ZN(n399) );
  XNOR2_X1 U456 ( .A(n400), .B(n399), .ZN(n401) );
  XNOR2_X1 U457 ( .A(n402), .B(n401), .ZN(n403) );
  XNOR2_X1 U458 ( .A(n404), .B(n403), .ZN(n550) );
  XOR2_X1 U459 ( .A(n406), .B(n405), .Z(n408) );
  NAND2_X1 U460 ( .A1(G226GAT), .A2(G233GAT), .ZN(n407) );
  XNOR2_X1 U461 ( .A(n408), .B(n407), .ZN(n409) );
  XOR2_X1 U462 ( .A(n409), .B(KEYINPUT96), .Z(n412) );
  XNOR2_X1 U463 ( .A(n410), .B(G92GAT), .ZN(n411) );
  XNOR2_X1 U464 ( .A(n412), .B(n411), .ZN(n414) );
  XOR2_X1 U465 ( .A(n414), .B(n413), .Z(n420) );
  XOR2_X1 U466 ( .A(KEYINPUT88), .B(G218GAT), .Z(n416) );
  XNOR2_X1 U467 ( .A(KEYINPUT21), .B(G211GAT), .ZN(n415) );
  XNOR2_X1 U468 ( .A(n416), .B(n415), .ZN(n417) );
  XOR2_X1 U469 ( .A(G197GAT), .B(n417), .Z(n431) );
  XNOR2_X1 U470 ( .A(n418), .B(n431), .ZN(n419) );
  XNOR2_X1 U471 ( .A(n420), .B(n419), .ZN(n547) );
  XNOR2_X1 U472 ( .A(n547), .B(KEYINPUT27), .ZN(n443) );
  OR2_X1 U473 ( .A1(n550), .A2(n443), .ZN(n518) );
  XOR2_X1 U474 ( .A(KEYINPUT92), .B(KEYINPUT90), .Z(n422) );
  XNOR2_X1 U475 ( .A(KEYINPUT91), .B(KEYINPUT22), .ZN(n421) );
  XNOR2_X1 U476 ( .A(n422), .B(n421), .ZN(n426) );
  XOR2_X1 U477 ( .A(G204GAT), .B(KEYINPUT23), .Z(n424) );
  XNOR2_X1 U478 ( .A(KEYINPUT24), .B(KEYINPUT89), .ZN(n423) );
  XNOR2_X1 U479 ( .A(n424), .B(n423), .ZN(n425) );
  XOR2_X1 U480 ( .A(n426), .B(n425), .Z(n433) );
  XOR2_X1 U481 ( .A(n427), .B(KEYINPUT87), .Z(n429) );
  NAND2_X1 U482 ( .A1(G228GAT), .A2(G233GAT), .ZN(n428) );
  XNOR2_X1 U483 ( .A(n429), .B(n428), .ZN(n430) );
  XNOR2_X1 U484 ( .A(n431), .B(n430), .ZN(n432) );
  XNOR2_X1 U485 ( .A(n433), .B(n432), .ZN(n435) );
  XOR2_X1 U486 ( .A(n435), .B(n434), .Z(n439) );
  XNOR2_X1 U487 ( .A(n437), .B(n436), .ZN(n438) );
  XNOR2_X1 U488 ( .A(n439), .B(n438), .ZN(n552) );
  XNOR2_X1 U489 ( .A(n552), .B(KEYINPUT28), .ZN(n522) );
  NOR2_X1 U490 ( .A1(n518), .A2(n522), .ZN(n440) );
  NAND2_X1 U491 ( .A1(n555), .A2(n440), .ZN(n451) );
  XOR2_X1 U492 ( .A(KEYINPUT97), .B(KEYINPUT26), .Z(n441) );
  XNOR2_X1 U493 ( .A(n442), .B(n441), .ZN(n571) );
  OR2_X1 U494 ( .A1(n571), .A2(n443), .ZN(n444) );
  XNOR2_X1 U495 ( .A(n444), .B(KEYINPUT98), .ZN(n448) );
  NOR2_X1 U496 ( .A1(n555), .A2(n547), .ZN(n445) );
  NOR2_X1 U497 ( .A1(n552), .A2(n445), .ZN(n446) );
  XNOR2_X1 U498 ( .A(KEYINPUT25), .B(n446), .ZN(n447) );
  NAND2_X1 U499 ( .A1(n448), .A2(n447), .ZN(n449) );
  NAND2_X1 U500 ( .A1(n449), .A2(n550), .ZN(n450) );
  NAND2_X1 U501 ( .A1(n451), .A2(n450), .ZN(n452) );
  XOR2_X1 U502 ( .A(KEYINPUT99), .B(n452), .Z(n463) );
  NAND2_X1 U503 ( .A1(n453), .A2(n463), .ZN(n482) );
  NOR2_X1 U504 ( .A1(n467), .A2(n482), .ZN(n461) );
  INV_X1 U505 ( .A(n550), .ZN(n494) );
  NAND2_X1 U506 ( .A1(n461), .A2(n494), .ZN(n454) );
  XNOR2_X1 U507 ( .A(n455), .B(n454), .ZN(G1324GAT) );
  INV_X1 U508 ( .A(n547), .ZN(n497) );
  NAND2_X1 U509 ( .A1(n497), .A2(n461), .ZN(n456) );
  XNOR2_X1 U510 ( .A(n456), .B(KEYINPUT102), .ZN(n457) );
  XNOR2_X1 U511 ( .A(G8GAT), .B(n457), .ZN(G1325GAT) );
  XOR2_X1 U512 ( .A(KEYINPUT35), .B(KEYINPUT103), .Z(n459) );
  NAND2_X1 U513 ( .A1(n461), .A2(n519), .ZN(n458) );
  XNOR2_X1 U514 ( .A(n459), .B(n458), .ZN(n460) );
  XOR2_X1 U515 ( .A(G15GAT), .B(n460), .Z(G1326GAT) );
  NAND2_X1 U516 ( .A1(n522), .A2(n461), .ZN(n462) );
  XNOR2_X1 U517 ( .A(n462), .B(G22GAT), .ZN(G1327GAT) );
  NAND2_X1 U518 ( .A1(n510), .A2(n463), .ZN(n465) );
  XNOR2_X1 U519 ( .A(KEYINPUT36), .B(KEYINPUT104), .ZN(n464) );
  XOR2_X1 U520 ( .A(n464), .B(n566), .Z(n585) );
  NOR2_X1 U521 ( .A1(n465), .A2(n585), .ZN(n466) );
  XNOR2_X1 U522 ( .A(n466), .B(KEYINPUT37), .ZN(n493) );
  NOR2_X1 U523 ( .A1(n493), .A2(n467), .ZN(n468) );
  NOR2_X1 U524 ( .A1(n476), .A2(n550), .ZN(n469) );
  XNOR2_X1 U525 ( .A(n469), .B(KEYINPUT39), .ZN(n470) );
  XNOR2_X1 U526 ( .A(G29GAT), .B(n470), .ZN(G1328GAT) );
  XNOR2_X1 U527 ( .A(G36GAT), .B(KEYINPUT105), .ZN(n472) );
  NOR2_X1 U528 ( .A1(n547), .A2(n476), .ZN(n471) );
  XNOR2_X1 U529 ( .A(n472), .B(n471), .ZN(G1329GAT) );
  XNOR2_X1 U530 ( .A(KEYINPUT106), .B(KEYINPUT40), .ZN(n474) );
  NOR2_X1 U531 ( .A1(n555), .A2(n476), .ZN(n473) );
  XNOR2_X1 U532 ( .A(n474), .B(n473), .ZN(n475) );
  XOR2_X1 U533 ( .A(n475), .B(G43GAT), .Z(G1330GAT) );
  INV_X1 U534 ( .A(n522), .ZN(n477) );
  NOR2_X1 U535 ( .A1(n477), .A2(n476), .ZN(n478) );
  XOR2_X1 U536 ( .A(G50GAT), .B(n478), .Z(G1331GAT) );
  XOR2_X1 U537 ( .A(KEYINPUT108), .B(KEYINPUT42), .Z(n484) );
  XNOR2_X1 U538 ( .A(n577), .B(KEYINPUT41), .ZN(n503) );
  INV_X1 U539 ( .A(n503), .ZN(n479) );
  INV_X1 U540 ( .A(n479), .ZN(n560) );
  INV_X1 U541 ( .A(n572), .ZN(n480) );
  NAND2_X1 U542 ( .A1(n560), .A2(n480), .ZN(n481) );
  XOR2_X1 U543 ( .A(KEYINPUT107), .B(n481), .Z(n492) );
  NOR2_X1 U544 ( .A1(n492), .A2(n482), .ZN(n488) );
  NAND2_X1 U545 ( .A1(n488), .A2(n494), .ZN(n483) );
  XNOR2_X1 U546 ( .A(n484), .B(n483), .ZN(n485) );
  XOR2_X1 U547 ( .A(G57GAT), .B(n485), .Z(G1332GAT) );
  NAND2_X1 U548 ( .A1(n497), .A2(n488), .ZN(n486) );
  XNOR2_X1 U549 ( .A(n486), .B(G64GAT), .ZN(G1333GAT) );
  NAND2_X1 U550 ( .A1(n519), .A2(n488), .ZN(n487) );
  XNOR2_X1 U551 ( .A(n487), .B(G71GAT), .ZN(G1334GAT) );
  XOR2_X1 U552 ( .A(KEYINPUT43), .B(KEYINPUT109), .Z(n490) );
  NAND2_X1 U553 ( .A1(n488), .A2(n522), .ZN(n489) );
  XNOR2_X1 U554 ( .A(n490), .B(n489), .ZN(n491) );
  XOR2_X1 U555 ( .A(G78GAT), .B(n491), .Z(G1335GAT) );
  NOR2_X1 U556 ( .A1(n493), .A2(n492), .ZN(n500) );
  NAND2_X1 U557 ( .A1(n500), .A2(n494), .ZN(n495) );
  XNOR2_X1 U558 ( .A(n495), .B(KEYINPUT110), .ZN(n496) );
  XNOR2_X1 U559 ( .A(G85GAT), .B(n496), .ZN(G1336GAT) );
  NAND2_X1 U560 ( .A1(n497), .A2(n500), .ZN(n498) );
  XNOR2_X1 U561 ( .A(n498), .B(G92GAT), .ZN(G1337GAT) );
  NAND2_X1 U562 ( .A1(n519), .A2(n500), .ZN(n499) );
  XNOR2_X1 U563 ( .A(n499), .B(G99GAT), .ZN(G1338GAT) );
  NAND2_X1 U564 ( .A1(n522), .A2(n500), .ZN(n501) );
  XNOR2_X1 U565 ( .A(n501), .B(KEYINPUT44), .ZN(n502) );
  XNOR2_X1 U566 ( .A(G106GAT), .B(n502), .ZN(G1339GAT) );
  XNOR2_X1 U567 ( .A(G113GAT), .B(KEYINPUT114), .ZN(n524) );
  XOR2_X1 U568 ( .A(KEYINPUT111), .B(KEYINPUT46), .Z(n505) );
  NAND2_X1 U569 ( .A1(n572), .A2(n503), .ZN(n504) );
  XNOR2_X1 U570 ( .A(n505), .B(n504), .ZN(n507) );
  NOR2_X1 U571 ( .A1(n582), .A2(n566), .ZN(n506) );
  NAND2_X1 U572 ( .A1(n507), .A2(n506), .ZN(n508) );
  XNOR2_X1 U573 ( .A(KEYINPUT112), .B(n508), .ZN(n509) );
  XNOR2_X1 U574 ( .A(n509), .B(KEYINPUT47), .ZN(n515) );
  NOR2_X1 U575 ( .A1(n510), .A2(n585), .ZN(n511) );
  XNOR2_X1 U576 ( .A(KEYINPUT45), .B(n511), .ZN(n512) );
  NAND2_X1 U577 ( .A1(n512), .A2(n577), .ZN(n513) );
  NOR2_X1 U578 ( .A1(n513), .A2(n572), .ZN(n514) );
  NOR2_X1 U579 ( .A1(n515), .A2(n514), .ZN(n516) );
  XNOR2_X1 U580 ( .A(n516), .B(KEYINPUT64), .ZN(n517) );
  XNOR2_X1 U581 ( .A(n517), .B(KEYINPUT48), .ZN(n548) );
  NOR2_X1 U582 ( .A1(n548), .A2(n518), .ZN(n535) );
  NAND2_X1 U583 ( .A1(n535), .A2(n519), .ZN(n520) );
  XOR2_X1 U584 ( .A(KEYINPUT113), .B(n520), .Z(n521) );
  NOR2_X1 U585 ( .A1(n522), .A2(n521), .ZN(n532) );
  NAND2_X1 U586 ( .A1(n572), .A2(n532), .ZN(n523) );
  XNOR2_X1 U587 ( .A(n524), .B(n523), .ZN(G1340GAT) );
  XOR2_X1 U588 ( .A(KEYINPUT49), .B(KEYINPUT116), .Z(n526) );
  NAND2_X1 U589 ( .A1(n532), .A2(n560), .ZN(n525) );
  XNOR2_X1 U590 ( .A(n526), .B(n525), .ZN(n528) );
  XOR2_X1 U591 ( .A(G120GAT), .B(KEYINPUT115), .Z(n527) );
  XNOR2_X1 U592 ( .A(n528), .B(n527), .ZN(G1341GAT) );
  XOR2_X1 U593 ( .A(KEYINPUT50), .B(KEYINPUT117), .Z(n530) );
  NAND2_X1 U594 ( .A1(n532), .A2(n582), .ZN(n529) );
  XNOR2_X1 U595 ( .A(n530), .B(n529), .ZN(n531) );
  XNOR2_X1 U596 ( .A(G127GAT), .B(n531), .ZN(G1342GAT) );
  XOR2_X1 U597 ( .A(G134GAT), .B(KEYINPUT51), .Z(n534) );
  NAND2_X1 U598 ( .A1(n532), .A2(n566), .ZN(n533) );
  XNOR2_X1 U599 ( .A(n534), .B(n533), .ZN(G1343GAT) );
  INV_X1 U600 ( .A(n571), .ZN(n536) );
  NAND2_X1 U601 ( .A1(n536), .A2(n535), .ZN(n537) );
  XOR2_X1 U602 ( .A(KEYINPUT118), .B(n537), .Z(n545) );
  NAND2_X1 U603 ( .A1(n545), .A2(n572), .ZN(n538) );
  XNOR2_X1 U604 ( .A(n538), .B(G141GAT), .ZN(G1344GAT) );
  XOR2_X1 U605 ( .A(KEYINPUT52), .B(KEYINPUT53), .Z(n540) );
  NAND2_X1 U606 ( .A1(n545), .A2(n560), .ZN(n539) );
  XNOR2_X1 U607 ( .A(n540), .B(n539), .ZN(n542) );
  XOR2_X1 U608 ( .A(G148GAT), .B(KEYINPUT119), .Z(n541) );
  XNOR2_X1 U609 ( .A(n542), .B(n541), .ZN(G1345GAT) );
  NAND2_X1 U610 ( .A1(n545), .A2(n582), .ZN(n543) );
  XNOR2_X1 U611 ( .A(n543), .B(KEYINPUT120), .ZN(n544) );
  XNOR2_X1 U612 ( .A(G155GAT), .B(n544), .ZN(G1346GAT) );
  NAND2_X1 U613 ( .A1(n545), .A2(n566), .ZN(n546) );
  XNOR2_X1 U614 ( .A(n546), .B(G162GAT), .ZN(G1347GAT) );
  NOR2_X1 U615 ( .A1(n548), .A2(n547), .ZN(n549) );
  XNOR2_X1 U616 ( .A(n549), .B(KEYINPUT54), .ZN(n551) );
  NAND2_X1 U617 ( .A1(n551), .A2(n550), .ZN(n570) );
  NOR2_X1 U618 ( .A1(n552), .A2(n570), .ZN(n553) );
  XNOR2_X1 U619 ( .A(n553), .B(KEYINPUT55), .ZN(n554) );
  NOR2_X1 U620 ( .A1(n555), .A2(n554), .ZN(n567) );
  NAND2_X1 U621 ( .A1(n572), .A2(n567), .ZN(n556) );
  XNOR2_X1 U622 ( .A(G169GAT), .B(n556), .ZN(G1348GAT) );
  XOR2_X1 U623 ( .A(KEYINPUT57), .B(KEYINPUT122), .Z(n558) );
  XNOR2_X1 U624 ( .A(G176GAT), .B(KEYINPUT56), .ZN(n557) );
  XNOR2_X1 U625 ( .A(n558), .B(n557), .ZN(n559) );
  XOR2_X1 U626 ( .A(KEYINPUT121), .B(n559), .Z(n562) );
  NAND2_X1 U627 ( .A1(n567), .A2(n560), .ZN(n561) );
  XNOR2_X1 U628 ( .A(n562), .B(n561), .ZN(G1349GAT) );
  XOR2_X1 U629 ( .A(KEYINPUT123), .B(KEYINPUT124), .Z(n564) );
  NAND2_X1 U630 ( .A1(n567), .A2(n582), .ZN(n563) );
  XNOR2_X1 U631 ( .A(n564), .B(n563), .ZN(n565) );
  XNOR2_X1 U632 ( .A(G183GAT), .B(n565), .ZN(G1350GAT) );
  NAND2_X1 U633 ( .A1(n567), .A2(n566), .ZN(n568) );
  XNOR2_X1 U634 ( .A(n568), .B(KEYINPUT58), .ZN(n569) );
  XNOR2_X1 U635 ( .A(G190GAT), .B(n569), .ZN(G1351GAT) );
  XOR2_X1 U636 ( .A(G197GAT), .B(KEYINPUT60), .Z(n574) );
  NOR2_X1 U637 ( .A1(n571), .A2(n570), .ZN(n581) );
  NAND2_X1 U638 ( .A1(n581), .A2(n572), .ZN(n573) );
  XNOR2_X1 U639 ( .A(n574), .B(n573), .ZN(n576) );
  XOR2_X1 U640 ( .A(KEYINPUT125), .B(KEYINPUT59), .Z(n575) );
  XNOR2_X1 U641 ( .A(n576), .B(n575), .ZN(G1352GAT) );
  XOR2_X1 U642 ( .A(KEYINPUT126), .B(KEYINPUT61), .Z(n579) );
  INV_X1 U643 ( .A(n581), .ZN(n584) );
  OR2_X1 U644 ( .A1(n584), .A2(n577), .ZN(n578) );
  XNOR2_X1 U645 ( .A(n579), .B(n578), .ZN(n580) );
  XNOR2_X1 U646 ( .A(G204GAT), .B(n580), .ZN(G1353GAT) );
  NAND2_X1 U647 ( .A1(n582), .A2(n581), .ZN(n583) );
  XNOR2_X1 U648 ( .A(n583), .B(G211GAT), .ZN(G1354GAT) );
  NOR2_X1 U649 ( .A1(n585), .A2(n584), .ZN(n587) );
  XNOR2_X1 U650 ( .A(KEYINPUT62), .B(KEYINPUT127), .ZN(n586) );
  XNOR2_X1 U651 ( .A(n587), .B(n586), .ZN(n588) );
  XNOR2_X1 U652 ( .A(G218GAT), .B(n588), .ZN(G1355GAT) );
endmodule

