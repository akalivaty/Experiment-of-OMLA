

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
         n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
         n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590,
         n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601,
         n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612,
         n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623,
         n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634,
         n635, n636, n637, n638, n639, n640, n641, n642, n643, n644, n645,
         n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, n656,
         n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n667,
         n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678,
         n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689,
         n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700,
         n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711,
         n712, n713, n714, n715, n716, n717, n718, n719, n720, n721, n722,
         n723, n724, n725, n726, n727, n728, n729, n730, n731, n732, n733,
         n734, n735, n736, n737, n738, n739, n740, n741, n742, n743, n744,
         n745, n746, n747, n748, n749, n750, n751, n752, n753, n754, n755,
         n756, n757, n758, n759, n760, n761, n762, n763, n764, n765, n766,
         n767, n768, n769, n770, n771, n772, n773, n774, n775, n776, n777,
         n778, n779, n780, n781, n782, n783, n784, n785, n786, n787, n788,
         n789, n790, n791, n792, n793, n794, n795, n796, n797, n798, n799,
         n800, n801, n802, n803, n804, n805, n806, n807, n808, n809, n810,
         n811, n812, n813, n814, n815, n816, n817, n818, n819, n820, n821,
         n822, n823, n824, n825, n826, n827, n828, n829, n830, n831, n832,
         n833, n834, n835, n836, n837, n838, n839, n840, n841, n842, n843,
         n844, n845, n846, n847, n848, n849, n850, n851, n852, n853, n854,
         n855, n856, n857, n858, n859, n860, n861, n862, n863, n864, n865,
         n866, n867, n868, n869, n870, n871, n872, n873, n874, n875, n876,
         n877, n878, n879, n880, n881, n882, n883, n884, n885, n886, n887,
         n888, n889, n890, n891, n892, n893, n894, n895, n896, n897, n898,
         n899, n900, n901, n902, n903, n904, n905, n906, n907, n908, n909,
         n910, n911, n912, n913, n914, n915, n916, n917, n918, n919, n920,
         n921, n922, n923, n924, n925, n926, n927, n928, n929, n930, n931,
         n932, n933, n934, n935, n936, n937, n938, n939, n940, n941, n942,
         n943, n944, n945, n946, n947, n948, n949, n950, n951, n952, n953,
         n954, n955, n956, n957, n958, n959, n960, n961, n962, n963, n964,
         n965, n966, n967, n968, n969, n970, n971, n972, n973, n974, n975,
         n976, n977, n978, n979, n980, n981, n982, n983, n984, n985, n986,
         n987, n988, n989, n990, n991, n992, n993, n994, n995, n996, n997,
         n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007,
         n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017,
         n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  AND2_X1 U556 ( .A1(n753), .A2(n521), .ZN(n754) );
  AND2_X1 U557 ( .A1(n540), .A2(G2104), .ZN(n879) );
  NOR2_X1 U558 ( .A1(n752), .A2(n751), .ZN(n521) );
  XNOR2_X1 U559 ( .A(n722), .B(KEYINPUT30), .ZN(n723) );
  INV_X1 U560 ( .A(n1004), .ZN(n751) );
  NOR2_X2 U561 ( .A1(n687), .A2(n686), .ZN(n716) );
  INV_X1 U562 ( .A(n716), .ZN(n732) );
  NOR2_X1 U563 ( .A1(G651), .A2(n634), .ZN(n640) );
  INV_X1 U564 ( .A(KEYINPUT64), .ZN(n545) );
  XNOR2_X1 U565 ( .A(n545), .B(KEYINPUT23), .ZN(n546) );
  XNOR2_X1 U566 ( .A(n547), .B(n546), .ZN(n553) );
  NOR2_X1 U567 ( .A1(G651), .A2(G543), .ZN(n647) );
  NAND2_X1 U568 ( .A1(G89), .A2(n647), .ZN(n522) );
  XNOR2_X1 U569 ( .A(n522), .B(KEYINPUT76), .ZN(n523) );
  XNOR2_X1 U570 ( .A(n523), .B(KEYINPUT4), .ZN(n525) );
  XOR2_X1 U571 ( .A(KEYINPUT0), .B(G543), .Z(n634) );
  INV_X1 U572 ( .A(G651), .ZN(n527) );
  NOR2_X1 U573 ( .A1(n634), .A2(n527), .ZN(n642) );
  NAND2_X1 U574 ( .A1(G76), .A2(n642), .ZN(n524) );
  NAND2_X1 U575 ( .A1(n525), .A2(n524), .ZN(n526) );
  XNOR2_X1 U576 ( .A(KEYINPUT5), .B(n526), .ZN(n534) );
  XNOR2_X1 U577 ( .A(KEYINPUT77), .B(KEYINPUT6), .ZN(n532) );
  NOR2_X1 U578 ( .A1(G543), .A2(n527), .ZN(n528) );
  XOR2_X1 U579 ( .A(KEYINPUT1), .B(n528), .Z(n644) );
  NAND2_X1 U580 ( .A1(G63), .A2(n644), .ZN(n530) );
  NAND2_X1 U581 ( .A1(G51), .A2(n640), .ZN(n529) );
  NAND2_X1 U582 ( .A1(n530), .A2(n529), .ZN(n531) );
  XNOR2_X1 U583 ( .A(n532), .B(n531), .ZN(n533) );
  NAND2_X1 U584 ( .A1(n534), .A2(n533), .ZN(n535) );
  XNOR2_X1 U585 ( .A(KEYINPUT7), .B(n535), .ZN(G168) );
  XNOR2_X1 U586 ( .A(KEYINPUT17), .B(KEYINPUT65), .ZN(n537) );
  NOR2_X1 U587 ( .A1(G2104), .A2(G2105), .ZN(n536) );
  XNOR2_X2 U588 ( .A(n537), .B(n536), .ZN(n878) );
  NAND2_X1 U589 ( .A1(G138), .A2(n878), .ZN(n539) );
  INV_X1 U590 ( .A(G2105), .ZN(n540) );
  NAND2_X1 U591 ( .A1(G102), .A2(n879), .ZN(n538) );
  NAND2_X1 U592 ( .A1(n539), .A2(n538), .ZN(n544) );
  NOR2_X1 U593 ( .A1(G2104), .A2(n540), .ZN(n885) );
  NAND2_X1 U594 ( .A1(G126), .A2(n885), .ZN(n542) );
  AND2_X1 U595 ( .A1(G2104), .A2(G2105), .ZN(n883) );
  NAND2_X1 U596 ( .A1(G114), .A2(n883), .ZN(n541) );
  NAND2_X1 U597 ( .A1(n542), .A2(n541), .ZN(n543) );
  NOR2_X1 U598 ( .A1(n544), .A2(n543), .ZN(G164) );
  NAND2_X1 U599 ( .A1(G101), .A2(n879), .ZN(n547) );
  AND2_X1 U600 ( .A1(G125), .A2(n885), .ZN(n551) );
  NAND2_X1 U601 ( .A1(G113), .A2(n883), .ZN(n549) );
  NAND2_X1 U602 ( .A1(G137), .A2(n878), .ZN(n548) );
  NAND2_X1 U603 ( .A1(n549), .A2(n548), .ZN(n550) );
  NOR2_X1 U604 ( .A1(n551), .A2(n550), .ZN(n552) );
  AND2_X1 U605 ( .A1(n553), .A2(n552), .ZN(G160) );
  NAND2_X1 U606 ( .A1(G90), .A2(n647), .ZN(n555) );
  NAND2_X1 U607 ( .A1(G77), .A2(n642), .ZN(n554) );
  NAND2_X1 U608 ( .A1(n555), .A2(n554), .ZN(n556) );
  XNOR2_X1 U609 ( .A(n556), .B(KEYINPUT9), .ZN(n558) );
  NAND2_X1 U610 ( .A1(G64), .A2(n644), .ZN(n557) );
  NAND2_X1 U611 ( .A1(n558), .A2(n557), .ZN(n561) );
  NAND2_X1 U612 ( .A1(G52), .A2(n640), .ZN(n559) );
  XNOR2_X1 U613 ( .A(KEYINPUT67), .B(n559), .ZN(n560) );
  NOR2_X1 U614 ( .A1(n561), .A2(n560), .ZN(G171) );
  AND2_X1 U615 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U616 ( .A(G132), .ZN(G219) );
  INV_X1 U617 ( .A(G82), .ZN(G220) );
  INV_X1 U618 ( .A(G57), .ZN(G237) );
  NAND2_X1 U619 ( .A1(n644), .A2(G62), .ZN(n564) );
  NAND2_X1 U620 ( .A1(G50), .A2(n640), .ZN(n562) );
  XOR2_X1 U621 ( .A(KEYINPUT83), .B(n562), .Z(n563) );
  NAND2_X1 U622 ( .A1(n564), .A2(n563), .ZN(n568) );
  NAND2_X1 U623 ( .A1(G88), .A2(n647), .ZN(n566) );
  NAND2_X1 U624 ( .A1(G75), .A2(n642), .ZN(n565) );
  NAND2_X1 U625 ( .A1(n566), .A2(n565), .ZN(n567) );
  NOR2_X1 U626 ( .A1(n568), .A2(n567), .ZN(G166) );
  NAND2_X1 U627 ( .A1(G7), .A2(G661), .ZN(n569) );
  XNOR2_X1 U628 ( .A(n569), .B(KEYINPUT10), .ZN(G223) );
  XNOR2_X1 U629 ( .A(G223), .B(KEYINPUT71), .ZN(n820) );
  NAND2_X1 U630 ( .A1(n820), .A2(G567), .ZN(n570) );
  XOR2_X1 U631 ( .A(KEYINPUT11), .B(n570), .Z(G234) );
  XOR2_X1 U632 ( .A(KEYINPUT14), .B(KEYINPUT72), .Z(n572) );
  NAND2_X1 U633 ( .A1(G56), .A2(n644), .ZN(n571) );
  XNOR2_X1 U634 ( .A(n572), .B(n571), .ZN(n578) );
  NAND2_X1 U635 ( .A1(n647), .A2(G81), .ZN(n573) );
  XNOR2_X1 U636 ( .A(n573), .B(KEYINPUT12), .ZN(n575) );
  NAND2_X1 U637 ( .A1(G68), .A2(n642), .ZN(n574) );
  NAND2_X1 U638 ( .A1(n575), .A2(n574), .ZN(n576) );
  XOR2_X1 U639 ( .A(KEYINPUT13), .B(n576), .Z(n577) );
  NOR2_X1 U640 ( .A1(n578), .A2(n577), .ZN(n580) );
  NAND2_X1 U641 ( .A1(n640), .A2(G43), .ZN(n579) );
  NAND2_X1 U642 ( .A1(n580), .A2(n579), .ZN(n996) );
  XNOR2_X1 U643 ( .A(G860), .B(KEYINPUT73), .ZN(n604) );
  OR2_X1 U644 ( .A1(n996), .A2(n604), .ZN(G153) );
  XOR2_X1 U645 ( .A(G171), .B(KEYINPUT74), .Z(G301) );
  NAND2_X1 U646 ( .A1(G868), .A2(G301), .ZN(n590) );
  NAND2_X1 U647 ( .A1(G54), .A2(n640), .ZN(n587) );
  NAND2_X1 U648 ( .A1(G79), .A2(n642), .ZN(n582) );
  NAND2_X1 U649 ( .A1(G66), .A2(n644), .ZN(n581) );
  NAND2_X1 U650 ( .A1(n582), .A2(n581), .ZN(n585) );
  NAND2_X1 U651 ( .A1(G92), .A2(n647), .ZN(n583) );
  XNOR2_X1 U652 ( .A(KEYINPUT75), .B(n583), .ZN(n584) );
  NOR2_X1 U653 ( .A1(n585), .A2(n584), .ZN(n586) );
  NAND2_X1 U654 ( .A1(n587), .A2(n586), .ZN(n588) );
  XOR2_X1 U655 ( .A(n588), .B(KEYINPUT15), .Z(n999) );
  INV_X1 U656 ( .A(G868), .ZN(n665) );
  NAND2_X1 U657 ( .A1(n999), .A2(n665), .ZN(n589) );
  NAND2_X1 U658 ( .A1(n590), .A2(n589), .ZN(G284) );
  NAND2_X1 U659 ( .A1(G91), .A2(n647), .ZN(n591) );
  XNOR2_X1 U660 ( .A(n591), .B(KEYINPUT68), .ZN(n599) );
  NAND2_X1 U661 ( .A1(G53), .A2(n640), .ZN(n592) );
  XNOR2_X1 U662 ( .A(n592), .B(KEYINPUT70), .ZN(n594) );
  NAND2_X1 U663 ( .A1(n644), .A2(G65), .ZN(n593) );
  NAND2_X1 U664 ( .A1(n594), .A2(n593), .ZN(n597) );
  NAND2_X1 U665 ( .A1(G78), .A2(n642), .ZN(n595) );
  XNOR2_X1 U666 ( .A(KEYINPUT69), .B(n595), .ZN(n596) );
  NOR2_X1 U667 ( .A1(n597), .A2(n596), .ZN(n598) );
  NAND2_X1 U668 ( .A1(n599), .A2(n598), .ZN(G299) );
  XOR2_X1 U669 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NOR2_X1 U670 ( .A1(G868), .A2(G299), .ZN(n600) );
  XNOR2_X1 U671 ( .A(n600), .B(KEYINPUT78), .ZN(n602) );
  NOR2_X1 U672 ( .A1(n665), .A2(G286), .ZN(n601) );
  NOR2_X1 U673 ( .A1(n602), .A2(n601), .ZN(n603) );
  XOR2_X1 U674 ( .A(KEYINPUT79), .B(n603), .Z(G297) );
  NAND2_X1 U675 ( .A1(n604), .A2(G559), .ZN(n605) );
  INV_X1 U676 ( .A(n999), .ZN(n898) );
  NAND2_X1 U677 ( .A1(n605), .A2(n898), .ZN(n606) );
  XNOR2_X1 U678 ( .A(n606), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U679 ( .A1(G868), .A2(n996), .ZN(n609) );
  NAND2_X1 U680 ( .A1(G868), .A2(n898), .ZN(n607) );
  NOR2_X1 U681 ( .A1(G559), .A2(n607), .ZN(n608) );
  NOR2_X1 U682 ( .A1(n609), .A2(n608), .ZN(G282) );
  NAND2_X1 U683 ( .A1(n885), .A2(G123), .ZN(n610) );
  XNOR2_X1 U684 ( .A(n610), .B(KEYINPUT18), .ZN(n612) );
  NAND2_X1 U685 ( .A1(G135), .A2(n878), .ZN(n611) );
  NAND2_X1 U686 ( .A1(n612), .A2(n611), .ZN(n613) );
  XNOR2_X1 U687 ( .A(KEYINPUT80), .B(n613), .ZN(n617) );
  NAND2_X1 U688 ( .A1(G111), .A2(n883), .ZN(n615) );
  NAND2_X1 U689 ( .A1(G99), .A2(n879), .ZN(n614) );
  NAND2_X1 U690 ( .A1(n615), .A2(n614), .ZN(n616) );
  NOR2_X1 U691 ( .A1(n617), .A2(n616), .ZN(n920) );
  XNOR2_X1 U692 ( .A(n920), .B(G2096), .ZN(n618) );
  INV_X1 U693 ( .A(G2100), .ZN(n830) );
  NAND2_X1 U694 ( .A1(n618), .A2(n830), .ZN(G156) );
  NAND2_X1 U695 ( .A1(n898), .A2(G559), .ZN(n660) );
  XNOR2_X1 U696 ( .A(n996), .B(n660), .ZN(n619) );
  NOR2_X1 U697 ( .A1(n619), .A2(G860), .ZN(n626) );
  NAND2_X1 U698 ( .A1(G93), .A2(n647), .ZN(n621) );
  NAND2_X1 U699 ( .A1(G67), .A2(n644), .ZN(n620) );
  NAND2_X1 U700 ( .A1(n621), .A2(n620), .ZN(n625) );
  NAND2_X1 U701 ( .A1(G80), .A2(n642), .ZN(n623) );
  NAND2_X1 U702 ( .A1(G55), .A2(n640), .ZN(n622) );
  NAND2_X1 U703 ( .A1(n623), .A2(n622), .ZN(n624) );
  OR2_X1 U704 ( .A1(n625), .A2(n624), .ZN(n664) );
  XOR2_X1 U705 ( .A(n626), .B(n664), .Z(G145) );
  NAND2_X1 U706 ( .A1(G85), .A2(n647), .ZN(n628) );
  NAND2_X1 U707 ( .A1(G72), .A2(n642), .ZN(n627) );
  NAND2_X1 U708 ( .A1(n628), .A2(n627), .ZN(n629) );
  XOR2_X1 U709 ( .A(KEYINPUT66), .B(n629), .Z(n633) );
  NAND2_X1 U710 ( .A1(G60), .A2(n644), .ZN(n631) );
  NAND2_X1 U711 ( .A1(G47), .A2(n640), .ZN(n630) );
  AND2_X1 U712 ( .A1(n631), .A2(n630), .ZN(n632) );
  NAND2_X1 U713 ( .A1(n633), .A2(n632), .ZN(G290) );
  NAND2_X1 U714 ( .A1(G49), .A2(n640), .ZN(n636) );
  NAND2_X1 U715 ( .A1(G87), .A2(n634), .ZN(n635) );
  NAND2_X1 U716 ( .A1(n636), .A2(n635), .ZN(n637) );
  NOR2_X1 U717 ( .A1(n644), .A2(n637), .ZN(n639) );
  NAND2_X1 U718 ( .A1(G651), .A2(G74), .ZN(n638) );
  NAND2_X1 U719 ( .A1(n639), .A2(n638), .ZN(G288) );
  NAND2_X1 U720 ( .A1(G48), .A2(n640), .ZN(n641) );
  XNOR2_X1 U721 ( .A(n641), .B(KEYINPUT82), .ZN(n652) );
  NAND2_X1 U722 ( .A1(n642), .A2(G73), .ZN(n643) );
  XNOR2_X1 U723 ( .A(n643), .B(KEYINPUT2), .ZN(n646) );
  NAND2_X1 U724 ( .A1(G61), .A2(n644), .ZN(n645) );
  NAND2_X1 U725 ( .A1(n646), .A2(n645), .ZN(n650) );
  NAND2_X1 U726 ( .A1(G86), .A2(n647), .ZN(n648) );
  XNOR2_X1 U727 ( .A(KEYINPUT81), .B(n648), .ZN(n649) );
  NOR2_X1 U728 ( .A1(n650), .A2(n649), .ZN(n651) );
  NAND2_X1 U729 ( .A1(n652), .A2(n651), .ZN(G305) );
  XNOR2_X1 U730 ( .A(KEYINPUT19), .B(G290), .ZN(n653) );
  XNOR2_X1 U731 ( .A(n653), .B(G288), .ZN(n654) );
  XNOR2_X1 U732 ( .A(KEYINPUT84), .B(n654), .ZN(n656) );
  XOR2_X1 U733 ( .A(G305), .B(G299), .Z(n655) );
  XNOR2_X1 U734 ( .A(n656), .B(n655), .ZN(n657) );
  XOR2_X1 U735 ( .A(n664), .B(n657), .Z(n658) );
  XOR2_X1 U736 ( .A(n658), .B(G166), .Z(n659) );
  XNOR2_X1 U737 ( .A(n996), .B(n659), .ZN(n899) );
  XNOR2_X1 U738 ( .A(n899), .B(KEYINPUT85), .ZN(n661) );
  XNOR2_X1 U739 ( .A(n661), .B(n660), .ZN(n662) );
  NAND2_X1 U740 ( .A1(n662), .A2(G868), .ZN(n663) );
  XNOR2_X1 U741 ( .A(n663), .B(KEYINPUT86), .ZN(n667) );
  NAND2_X1 U742 ( .A1(n665), .A2(n664), .ZN(n666) );
  NAND2_X1 U743 ( .A1(n667), .A2(n666), .ZN(G295) );
  NAND2_X1 U744 ( .A1(G2084), .A2(G2078), .ZN(n670) );
  XNOR2_X1 U745 ( .A(KEYINPUT87), .B(KEYINPUT20), .ZN(n668) );
  XNOR2_X1 U746 ( .A(n668), .B(KEYINPUT88), .ZN(n669) );
  XNOR2_X1 U747 ( .A(n670), .B(n669), .ZN(n671) );
  NAND2_X1 U748 ( .A1(n671), .A2(G2090), .ZN(n672) );
  XNOR2_X1 U749 ( .A(KEYINPUT21), .B(n672), .ZN(n673) );
  NAND2_X1 U750 ( .A1(n673), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U751 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NAND2_X1 U752 ( .A1(G69), .A2(G120), .ZN(n674) );
  NOR2_X1 U753 ( .A1(G237), .A2(n674), .ZN(n675) );
  NAND2_X1 U754 ( .A1(G108), .A2(n675), .ZN(n827) );
  NAND2_X1 U755 ( .A1(G567), .A2(n827), .ZN(n676) );
  XOR2_X1 U756 ( .A(KEYINPUT89), .B(n676), .Z(n681) );
  NOR2_X1 U757 ( .A1(G220), .A2(G219), .ZN(n677) );
  XOR2_X1 U758 ( .A(KEYINPUT22), .B(n677), .Z(n678) );
  NOR2_X1 U759 ( .A1(G218), .A2(n678), .ZN(n679) );
  NAND2_X1 U760 ( .A1(G96), .A2(n679), .ZN(n828) );
  NAND2_X1 U761 ( .A1(G2106), .A2(n828), .ZN(n680) );
  NAND2_X1 U762 ( .A1(n681), .A2(n680), .ZN(n829) );
  NAND2_X1 U763 ( .A1(G483), .A2(G661), .ZN(n682) );
  NOR2_X1 U764 ( .A1(n829), .A2(n682), .ZN(n826) );
  NAND2_X1 U765 ( .A1(n826), .A2(G36), .ZN(G176) );
  INV_X1 U766 ( .A(G166), .ZN(G303) );
  XNOR2_X1 U767 ( .A(G1986), .B(G290), .ZN(n1003) );
  NAND2_X1 U768 ( .A1(G160), .A2(G40), .ZN(n686) );
  NOR2_X1 U769 ( .A1(G164), .A2(G1384), .ZN(n685) );
  NOR2_X1 U770 ( .A1(n686), .A2(n685), .ZN(n683) );
  XNOR2_X1 U771 ( .A(n683), .B(KEYINPUT90), .ZN(n815) );
  NAND2_X1 U772 ( .A1(n1003), .A2(n815), .ZN(n803) );
  XNOR2_X1 U773 ( .A(G1981), .B(KEYINPUT101), .ZN(n684) );
  XNOR2_X1 U774 ( .A(n684), .B(G305), .ZN(n993) );
  INV_X1 U775 ( .A(n685), .ZN(n687) );
  NAND2_X1 U776 ( .A1(G8), .A2(n732), .ZN(n752) );
  INV_X1 U777 ( .A(n752), .ZN(n768) );
  NOR2_X1 U778 ( .A1(G1976), .A2(G288), .ZN(n688) );
  XNOR2_X1 U779 ( .A(KEYINPUT100), .B(n688), .ZN(n750) );
  AND2_X1 U780 ( .A1(n768), .A2(n750), .ZN(n689) );
  NAND2_X1 U781 ( .A1(KEYINPUT33), .A2(n689), .ZN(n690) );
  NAND2_X1 U782 ( .A1(n993), .A2(n690), .ZN(n756) );
  INV_X1 U783 ( .A(KEYINPUT97), .ZN(n695) );
  NAND2_X1 U784 ( .A1(G1996), .A2(n716), .ZN(n691) );
  XNOR2_X1 U785 ( .A(n691), .B(KEYINPUT26), .ZN(n693) );
  NAND2_X1 U786 ( .A1(G1341), .A2(n732), .ZN(n692) );
  NAND2_X1 U787 ( .A1(n693), .A2(n692), .ZN(n694) );
  XNOR2_X1 U788 ( .A(n695), .B(n694), .ZN(n696) );
  NOR2_X1 U789 ( .A1(n696), .A2(n996), .ZN(n697) );
  OR2_X1 U790 ( .A1(n898), .A2(n697), .ZN(n703) );
  NAND2_X1 U791 ( .A1(n697), .A2(n898), .ZN(n701) );
  NOR2_X1 U792 ( .A1(n716), .A2(G1348), .ZN(n699) );
  NOR2_X1 U793 ( .A1(G2067), .A2(n732), .ZN(n698) );
  NOR2_X1 U794 ( .A1(n699), .A2(n698), .ZN(n700) );
  NAND2_X1 U795 ( .A1(n701), .A2(n700), .ZN(n702) );
  NAND2_X1 U796 ( .A1(n703), .A2(n702), .ZN(n708) );
  INV_X1 U797 ( .A(G299), .ZN(n710) );
  NAND2_X1 U798 ( .A1(n716), .A2(G2072), .ZN(n704) );
  XNOR2_X1 U799 ( .A(n704), .B(KEYINPUT27), .ZN(n706) );
  AND2_X1 U800 ( .A1(G1956), .A2(n732), .ZN(n705) );
  NOR2_X1 U801 ( .A1(n706), .A2(n705), .ZN(n709) );
  NAND2_X1 U802 ( .A1(n710), .A2(n709), .ZN(n707) );
  NAND2_X1 U803 ( .A1(n708), .A2(n707), .ZN(n713) );
  NOR2_X1 U804 ( .A1(n710), .A2(n709), .ZN(n711) );
  XOR2_X1 U805 ( .A(n711), .B(KEYINPUT28), .Z(n712) );
  NAND2_X1 U806 ( .A1(n713), .A2(n712), .ZN(n714) );
  XOR2_X1 U807 ( .A(KEYINPUT29), .B(n714), .Z(n720) );
  NOR2_X1 U808 ( .A1(n716), .A2(G1961), .ZN(n715) );
  XOR2_X1 U809 ( .A(KEYINPUT96), .B(n715), .Z(n718) );
  XNOR2_X1 U810 ( .A(G2078), .B(KEYINPUT25), .ZN(n946) );
  NAND2_X1 U811 ( .A1(n716), .A2(n946), .ZN(n717) );
  NAND2_X1 U812 ( .A1(n718), .A2(n717), .ZN(n724) );
  NAND2_X1 U813 ( .A1(n724), .A2(G171), .ZN(n719) );
  NAND2_X1 U814 ( .A1(n720), .A2(n719), .ZN(n731) );
  NOR2_X1 U815 ( .A1(G1966), .A2(n752), .ZN(n744) );
  NOR2_X1 U816 ( .A1(G2084), .A2(n732), .ZN(n741) );
  NOR2_X1 U817 ( .A1(n744), .A2(n741), .ZN(n721) );
  NAND2_X1 U818 ( .A1(G8), .A2(n721), .ZN(n722) );
  NOR2_X1 U819 ( .A1(n723), .A2(G168), .ZN(n726) );
  NOR2_X1 U820 ( .A1(G171), .A2(n724), .ZN(n725) );
  NOR2_X1 U821 ( .A1(n726), .A2(n725), .ZN(n728) );
  INV_X1 U822 ( .A(KEYINPUT31), .ZN(n727) );
  XNOR2_X1 U823 ( .A(n728), .B(n727), .ZN(n729) );
  XNOR2_X1 U824 ( .A(KEYINPUT98), .B(n729), .ZN(n730) );
  NAND2_X1 U825 ( .A1(n731), .A2(n730), .ZN(n742) );
  NAND2_X1 U826 ( .A1(n742), .A2(G286), .ZN(n738) );
  NOR2_X1 U827 ( .A1(G2090), .A2(n732), .ZN(n733) );
  XNOR2_X1 U828 ( .A(KEYINPUT99), .B(n733), .ZN(n736) );
  NOR2_X1 U829 ( .A1(G1971), .A2(n752), .ZN(n734) );
  NOR2_X1 U830 ( .A1(G166), .A2(n734), .ZN(n735) );
  NAND2_X1 U831 ( .A1(n736), .A2(n735), .ZN(n737) );
  NAND2_X1 U832 ( .A1(n738), .A2(n737), .ZN(n739) );
  NAND2_X1 U833 ( .A1(n739), .A2(G8), .ZN(n740) );
  XNOR2_X1 U834 ( .A(n740), .B(KEYINPUT32), .ZN(n748) );
  NAND2_X1 U835 ( .A1(G8), .A2(n741), .ZN(n746) );
  INV_X1 U836 ( .A(n742), .ZN(n743) );
  NOR2_X1 U837 ( .A1(n744), .A2(n743), .ZN(n745) );
  NAND2_X1 U838 ( .A1(n746), .A2(n745), .ZN(n747) );
  NAND2_X1 U839 ( .A1(n748), .A2(n747), .ZN(n757) );
  NOR2_X1 U840 ( .A1(G1971), .A2(G303), .ZN(n749) );
  NOR2_X1 U841 ( .A1(n750), .A2(n749), .ZN(n998) );
  NAND2_X1 U842 ( .A1(n757), .A2(n998), .ZN(n753) );
  NAND2_X1 U843 ( .A1(G1976), .A2(G288), .ZN(n1004) );
  NOR2_X1 U844 ( .A1(KEYINPUT33), .A2(n754), .ZN(n755) );
  NOR2_X1 U845 ( .A1(n756), .A2(n755), .ZN(n763) );
  INV_X1 U846 ( .A(n757), .ZN(n760) );
  NAND2_X1 U847 ( .A1(G8), .A2(G166), .ZN(n758) );
  NOR2_X1 U848 ( .A1(G2090), .A2(n758), .ZN(n759) );
  NOR2_X1 U849 ( .A1(n760), .A2(n759), .ZN(n761) );
  NOR2_X1 U850 ( .A1(n768), .A2(n761), .ZN(n762) );
  NOR2_X1 U851 ( .A1(n763), .A2(n762), .ZN(n764) );
  XNOR2_X1 U852 ( .A(n764), .B(KEYINPUT102), .ZN(n771) );
  NOR2_X1 U853 ( .A1(G1981), .A2(G305), .ZN(n767) );
  XOR2_X1 U854 ( .A(KEYINPUT24), .B(KEYINPUT95), .Z(n765) );
  XNOR2_X1 U855 ( .A(KEYINPUT94), .B(n765), .ZN(n766) );
  XNOR2_X1 U856 ( .A(n767), .B(n766), .ZN(n769) );
  NAND2_X1 U857 ( .A1(n769), .A2(n768), .ZN(n770) );
  AND2_X1 U858 ( .A1(n771), .A2(n770), .ZN(n801) );
  NAND2_X1 U859 ( .A1(n885), .A2(G119), .ZN(n772) );
  XOR2_X1 U860 ( .A(KEYINPUT91), .B(n772), .Z(n774) );
  NAND2_X1 U861 ( .A1(n883), .A2(G107), .ZN(n773) );
  NAND2_X1 U862 ( .A1(n774), .A2(n773), .ZN(n775) );
  XOR2_X1 U863 ( .A(KEYINPUT92), .B(n775), .Z(n779) );
  NAND2_X1 U864 ( .A1(G131), .A2(n878), .ZN(n777) );
  NAND2_X1 U865 ( .A1(G95), .A2(n879), .ZN(n776) );
  AND2_X1 U866 ( .A1(n777), .A2(n776), .ZN(n778) );
  NAND2_X1 U867 ( .A1(n779), .A2(n778), .ZN(n860) );
  AND2_X1 U868 ( .A1(n860), .A2(G1991), .ZN(n789) );
  NAND2_X1 U869 ( .A1(G105), .A2(n879), .ZN(n780) );
  XOR2_X1 U870 ( .A(KEYINPUT38), .B(n780), .Z(n785) );
  NAND2_X1 U871 ( .A1(G129), .A2(n885), .ZN(n782) );
  NAND2_X1 U872 ( .A1(G117), .A2(n883), .ZN(n781) );
  NAND2_X1 U873 ( .A1(n782), .A2(n781), .ZN(n783) );
  XOR2_X1 U874 ( .A(KEYINPUT93), .B(n783), .Z(n784) );
  NOR2_X1 U875 ( .A1(n785), .A2(n784), .ZN(n787) );
  NAND2_X1 U876 ( .A1(n878), .A2(G141), .ZN(n786) );
  NAND2_X1 U877 ( .A1(n787), .A2(n786), .ZN(n861) );
  AND2_X1 U878 ( .A1(n861), .A2(G1996), .ZN(n788) );
  NOR2_X1 U879 ( .A1(n789), .A2(n788), .ZN(n922) );
  INV_X1 U880 ( .A(n922), .ZN(n790) );
  NAND2_X1 U881 ( .A1(n815), .A2(n790), .ZN(n804) );
  XNOR2_X1 U882 ( .A(KEYINPUT37), .B(G2067), .ZN(n813) );
  NAND2_X1 U883 ( .A1(G140), .A2(n878), .ZN(n792) );
  NAND2_X1 U884 ( .A1(G104), .A2(n879), .ZN(n791) );
  NAND2_X1 U885 ( .A1(n792), .A2(n791), .ZN(n793) );
  XNOR2_X1 U886 ( .A(KEYINPUT34), .B(n793), .ZN(n798) );
  NAND2_X1 U887 ( .A1(G128), .A2(n885), .ZN(n795) );
  NAND2_X1 U888 ( .A1(G116), .A2(n883), .ZN(n794) );
  NAND2_X1 U889 ( .A1(n795), .A2(n794), .ZN(n796) );
  XOR2_X1 U890 ( .A(KEYINPUT35), .B(n796), .Z(n797) );
  NOR2_X1 U891 ( .A1(n798), .A2(n797), .ZN(n799) );
  XNOR2_X1 U892 ( .A(KEYINPUT36), .B(n799), .ZN(n895) );
  NOR2_X1 U893 ( .A1(n813), .A2(n895), .ZN(n940) );
  NAND2_X1 U894 ( .A1(n940), .A2(n815), .ZN(n811) );
  NAND2_X1 U895 ( .A1(n804), .A2(n811), .ZN(n800) );
  NOR2_X1 U896 ( .A1(n801), .A2(n800), .ZN(n802) );
  NAND2_X1 U897 ( .A1(n803), .A2(n802), .ZN(n818) );
  NOR2_X1 U898 ( .A1(G1996), .A2(n861), .ZN(n935) );
  INV_X1 U899 ( .A(n804), .ZN(n808) );
  NOR2_X1 U900 ( .A1(G1986), .A2(G290), .ZN(n806) );
  NOR2_X1 U901 ( .A1(G1991), .A2(n860), .ZN(n805) );
  XOR2_X1 U902 ( .A(KEYINPUT103), .B(n805), .Z(n924) );
  NOR2_X1 U903 ( .A1(n806), .A2(n924), .ZN(n807) );
  NOR2_X1 U904 ( .A1(n808), .A2(n807), .ZN(n809) );
  NOR2_X1 U905 ( .A1(n935), .A2(n809), .ZN(n810) );
  XNOR2_X1 U906 ( .A(KEYINPUT39), .B(n810), .ZN(n812) );
  NAND2_X1 U907 ( .A1(n812), .A2(n811), .ZN(n814) );
  NAND2_X1 U908 ( .A1(n813), .A2(n895), .ZN(n925) );
  NAND2_X1 U909 ( .A1(n814), .A2(n925), .ZN(n816) );
  NAND2_X1 U910 ( .A1(n816), .A2(n815), .ZN(n817) );
  NAND2_X1 U911 ( .A1(n818), .A2(n817), .ZN(n819) );
  XNOR2_X1 U912 ( .A(KEYINPUT40), .B(n819), .ZN(G329) );
  NAND2_X1 U913 ( .A1(n820), .A2(G2106), .ZN(n821) );
  XOR2_X1 U914 ( .A(KEYINPUT105), .B(n821), .Z(G217) );
  INV_X1 U915 ( .A(G661), .ZN(n823) );
  NAND2_X1 U916 ( .A1(G2), .A2(G15), .ZN(n822) );
  NOR2_X1 U917 ( .A1(n823), .A2(n822), .ZN(n824) );
  XOR2_X1 U918 ( .A(KEYINPUT106), .B(n824), .Z(G259) );
  NAND2_X1 U919 ( .A1(G3), .A2(G1), .ZN(n825) );
  NAND2_X1 U920 ( .A1(n826), .A2(n825), .ZN(G188) );
  INV_X1 U922 ( .A(G120), .ZN(G236) );
  INV_X1 U923 ( .A(G96), .ZN(G221) );
  INV_X1 U924 ( .A(G69), .ZN(G235) );
  NOR2_X1 U925 ( .A1(n828), .A2(n827), .ZN(G325) );
  INV_X1 U926 ( .A(G325), .ZN(G261) );
  XNOR2_X1 U927 ( .A(KEYINPUT107), .B(n829), .ZN(G319) );
  XOR2_X1 U928 ( .A(KEYINPUT43), .B(KEYINPUT110), .Z(n832) );
  XOR2_X1 U929 ( .A(G2678), .B(n830), .Z(n831) );
  XNOR2_X1 U930 ( .A(n832), .B(n831), .ZN(n833) );
  XOR2_X1 U931 ( .A(n833), .B(KEYINPUT42), .Z(n835) );
  XNOR2_X1 U932 ( .A(G2078), .B(G2072), .ZN(n834) );
  XNOR2_X1 U933 ( .A(n835), .B(n834), .ZN(n839) );
  XOR2_X1 U934 ( .A(G2096), .B(G2084), .Z(n837) );
  XNOR2_X1 U935 ( .A(G2067), .B(G2090), .ZN(n836) );
  XNOR2_X1 U936 ( .A(n837), .B(n836), .ZN(n838) );
  XOR2_X1 U937 ( .A(n839), .B(n838), .Z(n841) );
  XNOR2_X1 U938 ( .A(KEYINPUT108), .B(KEYINPUT109), .ZN(n840) );
  XNOR2_X1 U939 ( .A(n841), .B(n840), .ZN(G227) );
  XOR2_X1 U940 ( .A(G1976), .B(G1971), .Z(n843) );
  XNOR2_X1 U941 ( .A(G1986), .B(G1961), .ZN(n842) );
  XNOR2_X1 U942 ( .A(n843), .B(n842), .ZN(n847) );
  XOR2_X1 U943 ( .A(G1966), .B(G1981), .Z(n845) );
  XNOR2_X1 U944 ( .A(G1996), .B(G1991), .ZN(n844) );
  XNOR2_X1 U945 ( .A(n845), .B(n844), .ZN(n846) );
  XOR2_X1 U946 ( .A(n847), .B(n846), .Z(n849) );
  XNOR2_X1 U947 ( .A(G2474), .B(KEYINPUT111), .ZN(n848) );
  XNOR2_X1 U948 ( .A(n849), .B(n848), .ZN(n850) );
  XNOR2_X1 U949 ( .A(KEYINPUT41), .B(n850), .ZN(n851) );
  XOR2_X1 U950 ( .A(n851), .B(G1956), .Z(G229) );
  NAND2_X1 U951 ( .A1(G112), .A2(n883), .ZN(n853) );
  NAND2_X1 U952 ( .A1(G100), .A2(n879), .ZN(n852) );
  NAND2_X1 U953 ( .A1(n853), .A2(n852), .ZN(n854) );
  XNOR2_X1 U954 ( .A(KEYINPUT112), .B(n854), .ZN(n859) );
  NAND2_X1 U955 ( .A1(n885), .A2(G124), .ZN(n855) );
  XNOR2_X1 U956 ( .A(n855), .B(KEYINPUT44), .ZN(n857) );
  NAND2_X1 U957 ( .A1(G136), .A2(n878), .ZN(n856) );
  NAND2_X1 U958 ( .A1(n857), .A2(n856), .ZN(n858) );
  NOR2_X1 U959 ( .A1(n859), .A2(n858), .ZN(G162) );
  XNOR2_X1 U960 ( .A(n861), .B(n860), .ZN(n868) );
  XOR2_X1 U961 ( .A(KEYINPUT117), .B(KEYINPUT46), .Z(n863) );
  XNOR2_X1 U962 ( .A(KEYINPUT48), .B(KEYINPUT118), .ZN(n862) );
  XNOR2_X1 U963 ( .A(n863), .B(n862), .ZN(n864) );
  XOR2_X1 U964 ( .A(n864), .B(G162), .Z(n866) );
  XNOR2_X1 U965 ( .A(G164), .B(G160), .ZN(n865) );
  XNOR2_X1 U966 ( .A(n866), .B(n865), .ZN(n867) );
  XNOR2_X1 U967 ( .A(n868), .B(n867), .ZN(n877) );
  NAND2_X1 U968 ( .A1(G130), .A2(n885), .ZN(n870) );
  NAND2_X1 U969 ( .A1(G118), .A2(n883), .ZN(n869) );
  NAND2_X1 U970 ( .A1(n870), .A2(n869), .ZN(n875) );
  NAND2_X1 U971 ( .A1(G142), .A2(n878), .ZN(n872) );
  NAND2_X1 U972 ( .A1(G106), .A2(n879), .ZN(n871) );
  NAND2_X1 U973 ( .A1(n872), .A2(n871), .ZN(n873) );
  XOR2_X1 U974 ( .A(KEYINPUT45), .B(n873), .Z(n874) );
  NOR2_X1 U975 ( .A1(n875), .A2(n874), .ZN(n876) );
  XOR2_X1 U976 ( .A(n877), .B(n876), .Z(n894) );
  NAND2_X1 U977 ( .A1(G139), .A2(n878), .ZN(n881) );
  NAND2_X1 U978 ( .A1(G103), .A2(n879), .ZN(n880) );
  NAND2_X1 U979 ( .A1(n881), .A2(n880), .ZN(n882) );
  XNOR2_X1 U980 ( .A(KEYINPUT113), .B(n882), .ZN(n891) );
  NAND2_X1 U981 ( .A1(n883), .A2(G115), .ZN(n884) );
  XNOR2_X1 U982 ( .A(n884), .B(KEYINPUT114), .ZN(n887) );
  NAND2_X1 U983 ( .A1(G127), .A2(n885), .ZN(n886) );
  NAND2_X1 U984 ( .A1(n887), .A2(n886), .ZN(n889) );
  XOR2_X1 U985 ( .A(KEYINPUT47), .B(KEYINPUT115), .Z(n888) );
  XNOR2_X1 U986 ( .A(n889), .B(n888), .ZN(n890) );
  NAND2_X1 U987 ( .A1(n891), .A2(n890), .ZN(n892) );
  XNOR2_X1 U988 ( .A(KEYINPUT116), .B(n892), .ZN(n927) );
  XNOR2_X1 U989 ( .A(n927), .B(n920), .ZN(n893) );
  XNOR2_X1 U990 ( .A(n894), .B(n893), .ZN(n896) );
  XOR2_X1 U991 ( .A(n896), .B(n895), .Z(n897) );
  NOR2_X1 U992 ( .A1(G37), .A2(n897), .ZN(G395) );
  XOR2_X1 U993 ( .A(G286), .B(n898), .Z(n900) );
  XNOR2_X1 U994 ( .A(n900), .B(n899), .ZN(n901) );
  XOR2_X1 U995 ( .A(G171), .B(n901), .Z(n902) );
  NOR2_X1 U996 ( .A1(G37), .A2(n902), .ZN(G397) );
  XOR2_X1 U997 ( .A(G2438), .B(KEYINPUT104), .Z(n904) );
  XNOR2_X1 U998 ( .A(G2443), .B(G2430), .ZN(n903) );
  XNOR2_X1 U999 ( .A(n904), .B(n903), .ZN(n905) );
  XOR2_X1 U1000 ( .A(n905), .B(G2435), .Z(n907) );
  XNOR2_X1 U1001 ( .A(G1348), .B(G1341), .ZN(n906) );
  XNOR2_X1 U1002 ( .A(n907), .B(n906), .ZN(n911) );
  XOR2_X1 U1003 ( .A(G2451), .B(G2427), .Z(n909) );
  XNOR2_X1 U1004 ( .A(G2454), .B(G2446), .ZN(n908) );
  XNOR2_X1 U1005 ( .A(n909), .B(n908), .ZN(n910) );
  XOR2_X1 U1006 ( .A(n911), .B(n910), .Z(n912) );
  NAND2_X1 U1007 ( .A1(G14), .A2(n912), .ZN(n918) );
  NAND2_X1 U1008 ( .A1(G319), .A2(n918), .ZN(n915) );
  NOR2_X1 U1009 ( .A1(G227), .A2(G229), .ZN(n913) );
  XNOR2_X1 U1010 ( .A(KEYINPUT49), .B(n913), .ZN(n914) );
  NOR2_X1 U1011 ( .A1(n915), .A2(n914), .ZN(n917) );
  NOR2_X1 U1012 ( .A1(G395), .A2(G397), .ZN(n916) );
  NAND2_X1 U1013 ( .A1(n917), .A2(n916), .ZN(G225) );
  INV_X1 U1014 ( .A(G225), .ZN(G308) );
  INV_X1 U1015 ( .A(G108), .ZN(G238) );
  INV_X1 U1016 ( .A(n918), .ZN(G401) );
  INV_X1 U1017 ( .A(KEYINPUT55), .ZN(n965) );
  XNOR2_X1 U1018 ( .A(KEYINPUT120), .B(KEYINPUT52), .ZN(n942) );
  XOR2_X1 U1019 ( .A(G2084), .B(G160), .Z(n919) );
  NOR2_X1 U1020 ( .A1(n920), .A2(n919), .ZN(n921) );
  NAND2_X1 U1021 ( .A1(n922), .A2(n921), .ZN(n923) );
  NOR2_X1 U1022 ( .A1(n924), .A2(n923), .ZN(n926) );
  NAND2_X1 U1023 ( .A1(n926), .A2(n925), .ZN(n932) );
  XOR2_X1 U1024 ( .A(G164), .B(G2078), .Z(n929) );
  XNOR2_X1 U1025 ( .A(G2072), .B(n927), .ZN(n928) );
  NOR2_X1 U1026 ( .A1(n929), .A2(n928), .ZN(n930) );
  XOR2_X1 U1027 ( .A(KEYINPUT50), .B(n930), .Z(n931) );
  NOR2_X1 U1028 ( .A1(n932), .A2(n931), .ZN(n938) );
  XNOR2_X1 U1029 ( .A(G2090), .B(G162), .ZN(n933) );
  XNOR2_X1 U1030 ( .A(n933), .B(KEYINPUT119), .ZN(n934) );
  NOR2_X1 U1031 ( .A1(n935), .A2(n934), .ZN(n936) );
  XOR2_X1 U1032 ( .A(KEYINPUT51), .B(n936), .Z(n937) );
  NAND2_X1 U1033 ( .A1(n938), .A2(n937), .ZN(n939) );
  NOR2_X1 U1034 ( .A1(n940), .A2(n939), .ZN(n941) );
  XNOR2_X1 U1035 ( .A(n942), .B(n941), .ZN(n943) );
  NAND2_X1 U1036 ( .A1(n965), .A2(n943), .ZN(n944) );
  NAND2_X1 U1037 ( .A1(n944), .A2(G29), .ZN(n1018) );
  XNOR2_X1 U1038 ( .A(G2084), .B(G34), .ZN(n945) );
  XNOR2_X1 U1039 ( .A(n945), .B(KEYINPUT54), .ZN(n963) );
  XNOR2_X1 U1040 ( .A(G2090), .B(G35), .ZN(n960) );
  XOR2_X1 U1041 ( .A(n946), .B(G27), .Z(n948) );
  XNOR2_X1 U1042 ( .A(G1996), .B(G32), .ZN(n947) );
  NOR2_X1 U1043 ( .A1(n948), .A2(n947), .ZN(n949) );
  XNOR2_X1 U1044 ( .A(KEYINPUT122), .B(n949), .ZN(n955) );
  XOR2_X1 U1045 ( .A(G2072), .B(G33), .Z(n950) );
  NAND2_X1 U1046 ( .A1(n950), .A2(G28), .ZN(n953) );
  XOR2_X1 U1047 ( .A(G25), .B(G1991), .Z(n951) );
  XNOR2_X1 U1048 ( .A(KEYINPUT121), .B(n951), .ZN(n952) );
  NOR2_X1 U1049 ( .A1(n953), .A2(n952), .ZN(n954) );
  NAND2_X1 U1050 ( .A1(n955), .A2(n954), .ZN(n957) );
  XNOR2_X1 U1051 ( .A(G26), .B(G2067), .ZN(n956) );
  NOR2_X1 U1052 ( .A1(n957), .A2(n956), .ZN(n958) );
  XNOR2_X1 U1053 ( .A(KEYINPUT53), .B(n958), .ZN(n959) );
  NOR2_X1 U1054 ( .A1(n960), .A2(n959), .ZN(n961) );
  XNOR2_X1 U1055 ( .A(n961), .B(KEYINPUT123), .ZN(n962) );
  NOR2_X1 U1056 ( .A1(n963), .A2(n962), .ZN(n964) );
  XNOR2_X1 U1057 ( .A(n965), .B(n964), .ZN(n966) );
  NOR2_X1 U1058 ( .A1(G29), .A2(n966), .ZN(n967) );
  XNOR2_X1 U1059 ( .A(KEYINPUT124), .B(n967), .ZN(n1016) );
  XOR2_X1 U1060 ( .A(G1961), .B(G5), .Z(n980) );
  XOR2_X1 U1061 ( .A(G20), .B(G1956), .Z(n971) );
  XNOR2_X1 U1062 ( .A(G1981), .B(G6), .ZN(n969) );
  XNOR2_X1 U1063 ( .A(G1341), .B(G19), .ZN(n968) );
  NOR2_X1 U1064 ( .A1(n969), .A2(n968), .ZN(n970) );
  NAND2_X1 U1065 ( .A1(n971), .A2(n970), .ZN(n974) );
  XOR2_X1 U1066 ( .A(KEYINPUT59), .B(G1348), .Z(n972) );
  XNOR2_X1 U1067 ( .A(G4), .B(n972), .ZN(n973) );
  NOR2_X1 U1068 ( .A1(n974), .A2(n973), .ZN(n975) );
  XOR2_X1 U1069 ( .A(KEYINPUT60), .B(n975), .Z(n977) );
  XNOR2_X1 U1070 ( .A(G1966), .B(G21), .ZN(n976) );
  NOR2_X1 U1071 ( .A1(n977), .A2(n976), .ZN(n978) );
  XNOR2_X1 U1072 ( .A(KEYINPUT126), .B(n978), .ZN(n979) );
  NAND2_X1 U1073 ( .A1(n980), .A2(n979), .ZN(n988) );
  XOR2_X1 U1074 ( .A(G1986), .B(G24), .Z(n984) );
  XNOR2_X1 U1075 ( .A(G1971), .B(G22), .ZN(n982) );
  XNOR2_X1 U1076 ( .A(G23), .B(G1976), .ZN(n981) );
  NOR2_X1 U1077 ( .A1(n982), .A2(n981), .ZN(n983) );
  NAND2_X1 U1078 ( .A1(n984), .A2(n983), .ZN(n985) );
  XOR2_X1 U1079 ( .A(KEYINPUT58), .B(n985), .Z(n986) );
  XNOR2_X1 U1080 ( .A(KEYINPUT127), .B(n986), .ZN(n987) );
  NOR2_X1 U1081 ( .A1(n988), .A2(n987), .ZN(n989) );
  XNOR2_X1 U1082 ( .A(n989), .B(KEYINPUT61), .ZN(n1013) );
  XOR2_X1 U1083 ( .A(G299), .B(G1956), .Z(n991) );
  XNOR2_X1 U1084 ( .A(G171), .B(G1961), .ZN(n990) );
  NAND2_X1 U1085 ( .A1(n991), .A2(n990), .ZN(n1011) );
  XOR2_X1 U1086 ( .A(G1966), .B(G168), .Z(n992) );
  XNOR2_X1 U1087 ( .A(KEYINPUT125), .B(n992), .ZN(n994) );
  NAND2_X1 U1088 ( .A1(n994), .A2(n993), .ZN(n995) );
  XNOR2_X1 U1089 ( .A(n995), .B(KEYINPUT57), .ZN(n1009) );
  XOR2_X1 U1090 ( .A(G1341), .B(n996), .Z(n997) );
  NAND2_X1 U1091 ( .A1(n998), .A2(n997), .ZN(n1007) );
  XOR2_X1 U1092 ( .A(n999), .B(G1348), .Z(n1001) );
  NAND2_X1 U1093 ( .A1(G1971), .A2(G303), .ZN(n1000) );
  NAND2_X1 U1094 ( .A1(n1001), .A2(n1000), .ZN(n1002) );
  NOR2_X1 U1095 ( .A1(n1003), .A2(n1002), .ZN(n1005) );
  NAND2_X1 U1096 ( .A1(n1005), .A2(n1004), .ZN(n1006) );
  NOR2_X1 U1097 ( .A1(n1007), .A2(n1006), .ZN(n1008) );
  NAND2_X1 U1098 ( .A1(n1009), .A2(n1008), .ZN(n1010) );
  NOR2_X1 U1099 ( .A1(n1011), .A2(n1010), .ZN(n1019) );
  NOR2_X1 U1100 ( .A1(KEYINPUT56), .A2(n1019), .ZN(n1012) );
  NOR2_X1 U1101 ( .A1(n1013), .A2(n1012), .ZN(n1014) );
  NOR2_X1 U1102 ( .A1(G16), .A2(n1014), .ZN(n1015) );
  NOR2_X1 U1103 ( .A1(n1016), .A2(n1015), .ZN(n1017) );
  NAND2_X1 U1104 ( .A1(n1018), .A2(n1017), .ZN(n1024) );
  INV_X1 U1105 ( .A(G16), .ZN(n1020) );
  NOR2_X1 U1106 ( .A1(n1020), .A2(n1019), .ZN(n1021) );
  NAND2_X1 U1107 ( .A1(KEYINPUT56), .A2(n1021), .ZN(n1022) );
  NAND2_X1 U1108 ( .A1(G11), .A2(n1022), .ZN(n1023) );
  NOR2_X1 U1109 ( .A1(n1024), .A2(n1023), .ZN(n1025) );
  XOR2_X1 U1110 ( .A(n1025), .B(KEYINPUT62), .Z(G150) );
  INV_X1 U1111 ( .A(G150), .ZN(G311) );
endmodule

