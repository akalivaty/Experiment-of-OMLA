

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301,
         n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312,
         n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323,
         n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334,
         n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
         n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583;

  XNOR2_X1 U323 ( .A(n330), .B(n329), .ZN(n331) );
  INV_X1 U324 ( .A(G50GAT), .ZN(n329) );
  NOR2_X1 U325 ( .A1(n523), .A2(n479), .ZN(n480) );
  XNOR2_X1 U326 ( .A(n388), .B(n387), .ZN(n526) );
  AND2_X1 U327 ( .A1(G226GAT), .A2(G233GAT), .ZN(n291) );
  XOR2_X1 U328 ( .A(n317), .B(n316), .Z(n292) );
  XOR2_X1 U329 ( .A(KEYINPUT94), .B(KEYINPUT92), .Z(n293) );
  XOR2_X1 U330 ( .A(KEYINPUT40), .B(n508), .Z(n294) );
  XNOR2_X1 U331 ( .A(n318), .B(n292), .ZN(n319) );
  XNOR2_X1 U332 ( .A(n320), .B(n319), .ZN(n326) );
  XNOR2_X1 U333 ( .A(n332), .B(n331), .ZN(n337) );
  XNOR2_X1 U334 ( .A(n379), .B(n291), .ZN(n380) );
  XNOR2_X1 U335 ( .A(n433), .B(n380), .ZN(n382) );
  XNOR2_X1 U336 ( .A(KEYINPUT37), .B(n502), .ZN(n522) );
  XOR2_X1 U337 ( .A(KEYINPUT122), .B(n457), .Z(n564) );
  XNOR2_X1 U338 ( .A(n346), .B(n345), .ZN(n568) );
  XNOR2_X1 U339 ( .A(n504), .B(KEYINPUT38), .ZN(n509) );
  XNOR2_X1 U340 ( .A(n463), .B(n462), .ZN(n464) );
  XNOR2_X1 U341 ( .A(n465), .B(n464), .ZN(G1351GAT) );
  XOR2_X1 U342 ( .A(G57GAT), .B(KEYINPUT13), .Z(n310) );
  XOR2_X1 U343 ( .A(G22GAT), .B(G155GAT), .Z(n428) );
  XOR2_X1 U344 ( .A(n310), .B(n428), .Z(n296) );
  XOR2_X1 U345 ( .A(KEYINPUT70), .B(G1GAT), .Z(n328) );
  XOR2_X1 U346 ( .A(G15GAT), .B(G127GAT), .Z(n436) );
  XNOR2_X1 U347 ( .A(n328), .B(n436), .ZN(n295) );
  XNOR2_X1 U348 ( .A(n296), .B(n295), .ZN(n309) );
  XOR2_X1 U349 ( .A(KEYINPUT80), .B(KEYINPUT12), .Z(n298) );
  NAND2_X1 U350 ( .A1(G231GAT), .A2(G233GAT), .ZN(n297) );
  XNOR2_X1 U351 ( .A(n298), .B(n297), .ZN(n299) );
  XOR2_X1 U352 ( .A(n299), .B(KEYINPUT15), .Z(n307) );
  XOR2_X1 U353 ( .A(G78GAT), .B(G211GAT), .Z(n301) );
  XNOR2_X1 U354 ( .A(G183GAT), .B(G71GAT), .ZN(n300) );
  XNOR2_X1 U355 ( .A(n301), .B(n300), .ZN(n305) );
  XOR2_X1 U356 ( .A(KEYINPUT79), .B(KEYINPUT14), .Z(n303) );
  XNOR2_X1 U357 ( .A(G8GAT), .B(G64GAT), .ZN(n302) );
  XNOR2_X1 U358 ( .A(n303), .B(n302), .ZN(n304) );
  XNOR2_X1 U359 ( .A(n305), .B(n304), .ZN(n306) );
  XNOR2_X1 U360 ( .A(n307), .B(n306), .ZN(n308) );
  XOR2_X1 U361 ( .A(n309), .B(n308), .Z(n577) );
  XNOR2_X1 U362 ( .A(KEYINPUT41), .B(KEYINPUT64), .ZN(n327) );
  XOR2_X1 U363 ( .A(G99GAT), .B(G85GAT), .Z(n352) );
  XOR2_X1 U364 ( .A(n310), .B(n352), .Z(n312) );
  NAND2_X1 U365 ( .A1(G230GAT), .A2(G233GAT), .ZN(n311) );
  XNOR2_X1 U366 ( .A(n312), .B(n311), .ZN(n320) );
  XOR2_X1 U367 ( .A(G120GAT), .B(G71GAT), .Z(n435) );
  XOR2_X1 U368 ( .A(KEYINPUT76), .B(KEYINPUT31), .Z(n314) );
  XNOR2_X1 U369 ( .A(KEYINPUT73), .B(KEYINPUT74), .ZN(n313) );
  XNOR2_X1 U370 ( .A(n314), .B(n313), .ZN(n315) );
  XNOR2_X1 U371 ( .A(n435), .B(n315), .ZN(n318) );
  XOR2_X1 U372 ( .A(KEYINPUT72), .B(KEYINPUT32), .Z(n317) );
  XNOR2_X1 U373 ( .A(KEYINPUT77), .B(KEYINPUT33), .ZN(n316) );
  XOR2_X1 U374 ( .A(G78GAT), .B(G148GAT), .Z(n322) );
  XNOR2_X1 U375 ( .A(G106GAT), .B(KEYINPUT75), .ZN(n321) );
  XNOR2_X1 U376 ( .A(n322), .B(n321), .ZN(n420) );
  XOR2_X1 U377 ( .A(G64GAT), .B(G92GAT), .Z(n324) );
  XNOR2_X1 U378 ( .A(G176GAT), .B(G204GAT), .ZN(n323) );
  XNOR2_X1 U379 ( .A(n324), .B(n323), .ZN(n381) );
  XOR2_X1 U380 ( .A(n420), .B(n381), .Z(n325) );
  XNOR2_X1 U381 ( .A(n326), .B(n325), .ZN(n369) );
  XOR2_X1 U382 ( .A(n327), .B(n369), .Z(n511) );
  XOR2_X1 U383 ( .A(G169GAT), .B(G8GAT), .Z(n386) );
  XNOR2_X1 U384 ( .A(n386), .B(n328), .ZN(n332) );
  XOR2_X1 U385 ( .A(G113GAT), .B(G15GAT), .Z(n330) );
  XOR2_X1 U386 ( .A(KEYINPUT29), .B(G197GAT), .Z(n334) );
  XNOR2_X1 U387 ( .A(G141GAT), .B(G22GAT), .ZN(n333) );
  XNOR2_X1 U388 ( .A(n334), .B(n333), .ZN(n335) );
  XNOR2_X1 U389 ( .A(n335), .B(G36GAT), .ZN(n336) );
  XNOR2_X1 U390 ( .A(n337), .B(n336), .ZN(n341) );
  XOR2_X1 U391 ( .A(KEYINPUT68), .B(KEYINPUT30), .Z(n339) );
  NAND2_X1 U392 ( .A1(G229GAT), .A2(G233GAT), .ZN(n338) );
  XNOR2_X1 U393 ( .A(n339), .B(n338), .ZN(n340) );
  XOR2_X1 U394 ( .A(n341), .B(n340), .Z(n346) );
  XOR2_X1 U395 ( .A(KEYINPUT8), .B(KEYINPUT69), .Z(n343) );
  XNOR2_X1 U396 ( .A(G43GAT), .B(G29GAT), .ZN(n342) );
  XNOR2_X1 U397 ( .A(n343), .B(n342), .ZN(n344) );
  XOR2_X1 U398 ( .A(KEYINPUT7), .B(n344), .Z(n365) );
  XNOR2_X1 U399 ( .A(n365), .B(KEYINPUT71), .ZN(n345) );
  INV_X1 U400 ( .A(n568), .ZN(n347) );
  OR2_X1 U401 ( .A1(n511), .A2(n347), .ZN(n349) );
  XNOR2_X1 U402 ( .A(KEYINPUT113), .B(KEYINPUT46), .ZN(n348) );
  XNOR2_X1 U403 ( .A(n349), .B(n348), .ZN(n350) );
  NOR2_X1 U404 ( .A1(n577), .A2(n350), .ZN(n351) );
  XNOR2_X1 U405 ( .A(n351), .B(KEYINPUT114), .ZN(n366) );
  XOR2_X1 U406 ( .A(G36GAT), .B(G190GAT), .Z(n379) );
  XOR2_X1 U407 ( .A(n352), .B(n379), .Z(n354) );
  NAND2_X1 U408 ( .A1(G232GAT), .A2(G233GAT), .ZN(n353) );
  XNOR2_X1 U409 ( .A(n354), .B(n353), .ZN(n358) );
  XOR2_X1 U410 ( .A(KEYINPUT10), .B(G92GAT), .Z(n356) );
  XNOR2_X1 U411 ( .A(G134GAT), .B(G106GAT), .ZN(n355) );
  XNOR2_X1 U412 ( .A(n356), .B(n355), .ZN(n357) );
  XOR2_X1 U413 ( .A(n358), .B(n357), .Z(n363) );
  XOR2_X1 U414 ( .A(G50GAT), .B(G162GAT), .Z(n429) );
  XOR2_X1 U415 ( .A(KEYINPUT11), .B(KEYINPUT67), .Z(n360) );
  XNOR2_X1 U416 ( .A(G218GAT), .B(KEYINPUT9), .ZN(n359) );
  XNOR2_X1 U417 ( .A(n360), .B(n359), .ZN(n361) );
  XNOR2_X1 U418 ( .A(n429), .B(n361), .ZN(n362) );
  XNOR2_X1 U419 ( .A(n363), .B(n362), .ZN(n364) );
  XNOR2_X1 U420 ( .A(n365), .B(n364), .ZN(n485) );
  NAND2_X1 U421 ( .A1(n366), .A2(n485), .ZN(n367) );
  XNOR2_X1 U422 ( .A(n367), .B(KEYINPUT47), .ZN(n373) );
  XNOR2_X1 U423 ( .A(KEYINPUT36), .B(n485), .ZN(n581) );
  INV_X1 U424 ( .A(n577), .ZN(n500) );
  NOR2_X1 U425 ( .A1(n581), .A2(n500), .ZN(n368) );
  XNOR2_X1 U426 ( .A(n368), .B(KEYINPUT45), .ZN(n370) );
  NAND2_X1 U427 ( .A1(n370), .A2(n369), .ZN(n371) );
  NOR2_X1 U428 ( .A1(n568), .A2(n371), .ZN(n372) );
  NOR2_X1 U429 ( .A1(n373), .A2(n372), .ZN(n374) );
  XNOR2_X1 U430 ( .A(KEYINPUT48), .B(n374), .ZN(n534) );
  XNOR2_X1 U431 ( .A(G218GAT), .B(KEYINPUT93), .ZN(n375) );
  XNOR2_X1 U432 ( .A(n293), .B(n375), .ZN(n376) );
  XOR2_X1 U433 ( .A(n376), .B(KEYINPUT21), .Z(n378) );
  XNOR2_X1 U434 ( .A(G197GAT), .B(G211GAT), .ZN(n377) );
  XNOR2_X1 U435 ( .A(n378), .B(n377), .ZN(n433) );
  XOR2_X1 U436 ( .A(n382), .B(n381), .Z(n388) );
  XOR2_X1 U437 ( .A(KEYINPUT18), .B(KEYINPUT19), .Z(n384) );
  XNOR2_X1 U438 ( .A(KEYINPUT87), .B(G183GAT), .ZN(n383) );
  XNOR2_X1 U439 ( .A(n384), .B(n383), .ZN(n385) );
  XOR2_X1 U440 ( .A(KEYINPUT17), .B(n385), .Z(n453) );
  XNOR2_X1 U441 ( .A(n386), .B(n453), .ZN(n387) );
  XOR2_X1 U442 ( .A(KEYINPUT121), .B(n526), .Z(n389) );
  NOR2_X1 U443 ( .A1(n534), .A2(n389), .ZN(n390) );
  XNOR2_X1 U444 ( .A(n390), .B(KEYINPUT54), .ZN(n415) );
  NAND2_X1 U445 ( .A1(G225GAT), .A2(G233GAT), .ZN(n396) );
  XOR2_X1 U446 ( .A(G85GAT), .B(G155GAT), .Z(n392) );
  XNOR2_X1 U447 ( .A(G127GAT), .B(G120GAT), .ZN(n391) );
  XNOR2_X1 U448 ( .A(n392), .B(n391), .ZN(n394) );
  XOR2_X1 U449 ( .A(G29GAT), .B(G162GAT), .Z(n393) );
  XNOR2_X1 U450 ( .A(n394), .B(n393), .ZN(n395) );
  XNOR2_X1 U451 ( .A(n396), .B(n395), .ZN(n414) );
  XOR2_X1 U452 ( .A(KEYINPUT100), .B(KEYINPUT98), .Z(n398) );
  XNOR2_X1 U453 ( .A(KEYINPUT6), .B(KEYINPUT99), .ZN(n397) );
  XNOR2_X1 U454 ( .A(n398), .B(n397), .ZN(n412) );
  XOR2_X1 U455 ( .A(KEYINPUT101), .B(G57GAT), .Z(n400) );
  XNOR2_X1 U456 ( .A(G1GAT), .B(G148GAT), .ZN(n399) );
  XNOR2_X1 U457 ( .A(n400), .B(n399), .ZN(n404) );
  XOR2_X1 U458 ( .A(KEYINPUT1), .B(KEYINPUT4), .Z(n402) );
  XNOR2_X1 U459 ( .A(KEYINPUT97), .B(KEYINPUT5), .ZN(n401) );
  XNOR2_X1 U460 ( .A(n402), .B(n401), .ZN(n403) );
  XOR2_X1 U461 ( .A(n404), .B(n403), .Z(n410) );
  XOR2_X1 U462 ( .A(KEYINPUT0), .B(KEYINPUT82), .Z(n406) );
  XNOR2_X1 U463 ( .A(G113GAT), .B(G134GAT), .ZN(n405) );
  XNOR2_X1 U464 ( .A(n406), .B(n405), .ZN(n440) );
  XOR2_X1 U465 ( .A(KEYINPUT2), .B(KEYINPUT3), .Z(n408) );
  XNOR2_X1 U466 ( .A(G141GAT), .B(KEYINPUT95), .ZN(n407) );
  XNOR2_X1 U467 ( .A(n408), .B(n407), .ZN(n421) );
  XNOR2_X1 U468 ( .A(n440), .B(n421), .ZN(n409) );
  XNOR2_X1 U469 ( .A(n410), .B(n409), .ZN(n411) );
  XOR2_X1 U470 ( .A(n412), .B(n411), .Z(n413) );
  XNOR2_X1 U471 ( .A(n414), .B(n413), .ZN(n523) );
  NAND2_X1 U472 ( .A1(n415), .A2(n523), .ZN(n416) );
  XNOR2_X1 U473 ( .A(n416), .B(KEYINPUT65), .ZN(n567) );
  XOR2_X1 U474 ( .A(KEYINPUT91), .B(G204GAT), .Z(n418) );
  NAND2_X1 U475 ( .A1(G228GAT), .A2(G233GAT), .ZN(n417) );
  XNOR2_X1 U476 ( .A(n418), .B(n417), .ZN(n419) );
  XOR2_X1 U477 ( .A(n419), .B(KEYINPUT22), .Z(n423) );
  XNOR2_X1 U478 ( .A(n421), .B(n420), .ZN(n422) );
  XNOR2_X1 U479 ( .A(n423), .B(n422), .ZN(n427) );
  XOR2_X1 U480 ( .A(KEYINPUT90), .B(KEYINPUT24), .Z(n425) );
  XNOR2_X1 U481 ( .A(KEYINPUT23), .B(KEYINPUT96), .ZN(n424) );
  XNOR2_X1 U482 ( .A(n425), .B(n424), .ZN(n426) );
  XOR2_X1 U483 ( .A(n427), .B(n426), .Z(n431) );
  XNOR2_X1 U484 ( .A(n429), .B(n428), .ZN(n430) );
  XNOR2_X1 U485 ( .A(n431), .B(n430), .ZN(n432) );
  XOR2_X1 U486 ( .A(n433), .B(n432), .Z(n481) );
  NAND2_X1 U487 ( .A1(n567), .A2(n481), .ZN(n434) );
  XNOR2_X1 U488 ( .A(n434), .B(KEYINPUT55), .ZN(n456) );
  XOR2_X1 U489 ( .A(KEYINPUT86), .B(G99GAT), .Z(n438) );
  XNOR2_X1 U490 ( .A(n436), .B(n435), .ZN(n437) );
  XNOR2_X1 U491 ( .A(n438), .B(n437), .ZN(n439) );
  XOR2_X1 U492 ( .A(n439), .B(G190GAT), .Z(n445) );
  XOR2_X1 U493 ( .A(n440), .B(G176GAT), .Z(n442) );
  NAND2_X1 U494 ( .A1(G227GAT), .A2(G233GAT), .ZN(n441) );
  XNOR2_X1 U495 ( .A(n442), .B(n441), .ZN(n443) );
  XNOR2_X1 U496 ( .A(G43GAT), .B(n443), .ZN(n444) );
  XNOR2_X1 U497 ( .A(n445), .B(n444), .ZN(n449) );
  XOR2_X1 U498 ( .A(KEYINPUT89), .B(KEYINPUT66), .Z(n447) );
  XNOR2_X1 U499 ( .A(G169GAT), .B(KEYINPUT20), .ZN(n446) );
  XNOR2_X1 U500 ( .A(n447), .B(n446), .ZN(n448) );
  XOR2_X1 U501 ( .A(n449), .B(n448), .Z(n455) );
  XOR2_X1 U502 ( .A(KEYINPUT88), .B(KEYINPUT84), .Z(n451) );
  XNOR2_X1 U503 ( .A(KEYINPUT83), .B(KEYINPUT85), .ZN(n450) );
  XNOR2_X1 U504 ( .A(n451), .B(n450), .ZN(n452) );
  XNOR2_X1 U505 ( .A(n453), .B(n452), .ZN(n454) );
  XNOR2_X1 U506 ( .A(n455), .B(n454), .ZN(n482) );
  NAND2_X1 U507 ( .A1(n456), .A2(n482), .ZN(n457) );
  INV_X1 U508 ( .A(n511), .ZN(n553) );
  NAND2_X1 U509 ( .A1(n564), .A2(n553), .ZN(n461) );
  XOR2_X1 U510 ( .A(KEYINPUT57), .B(KEYINPUT123), .Z(n459) );
  XOR2_X1 U511 ( .A(G176GAT), .B(KEYINPUT56), .Z(n458) );
  XNOR2_X1 U512 ( .A(n459), .B(n458), .ZN(n460) );
  XNOR2_X1 U513 ( .A(n461), .B(n460), .ZN(G1349GAT) );
  INV_X1 U514 ( .A(n485), .ZN(n559) );
  NAND2_X1 U515 ( .A1(n559), .A2(n564), .ZN(n465) );
  XOR2_X1 U516 ( .A(KEYINPUT124), .B(KEYINPUT58), .Z(n463) );
  INV_X1 U517 ( .A(G190GAT), .ZN(n462) );
  INV_X1 U518 ( .A(n482), .ZN(n535) );
  NOR2_X1 U519 ( .A1(n526), .A2(n535), .ZN(n466) );
  XNOR2_X1 U520 ( .A(KEYINPUT105), .B(n466), .ZN(n467) );
  NAND2_X1 U521 ( .A1(n467), .A2(n481), .ZN(n469) );
  XOR2_X1 U522 ( .A(KEYINPUT106), .B(KEYINPUT107), .Z(n468) );
  XNOR2_X1 U523 ( .A(n469), .B(n468), .ZN(n470) );
  XNOR2_X1 U524 ( .A(n470), .B(KEYINPUT25), .ZN(n476) );
  XNOR2_X1 U525 ( .A(KEYINPUT104), .B(KEYINPUT26), .ZN(n472) );
  NOR2_X1 U526 ( .A1(n482), .A2(n481), .ZN(n471) );
  XNOR2_X1 U527 ( .A(n472), .B(n471), .ZN(n566) );
  INV_X1 U528 ( .A(n566), .ZN(n474) );
  XNOR2_X1 U529 ( .A(n526), .B(KEYINPUT102), .ZN(n473) );
  XNOR2_X1 U530 ( .A(n473), .B(KEYINPUT27), .ZN(n479) );
  NOR2_X1 U531 ( .A1(n474), .A2(n479), .ZN(n475) );
  NOR2_X1 U532 ( .A1(n476), .A2(n475), .ZN(n478) );
  INV_X1 U533 ( .A(n523), .ZN(n477) );
  NOR2_X1 U534 ( .A1(n478), .A2(n477), .ZN(n484) );
  XOR2_X1 U535 ( .A(KEYINPUT103), .B(n480), .Z(n549) );
  XNOR2_X1 U536 ( .A(n481), .B(KEYINPUT28), .ZN(n531) );
  NAND2_X1 U537 ( .A1(n549), .A2(n531), .ZN(n537) );
  NOR2_X1 U538 ( .A1(n482), .A2(n537), .ZN(n483) );
  NOR2_X1 U539 ( .A1(n484), .A2(n483), .ZN(n499) );
  XOR2_X1 U540 ( .A(KEYINPUT81), .B(KEYINPUT16), .Z(n487) );
  NAND2_X1 U541 ( .A1(n577), .A2(n485), .ZN(n486) );
  XNOR2_X1 U542 ( .A(n487), .B(n486), .ZN(n488) );
  NOR2_X1 U543 ( .A1(n499), .A2(n488), .ZN(n512) );
  NAND2_X1 U544 ( .A1(n369), .A2(n568), .ZN(n489) );
  XOR2_X1 U545 ( .A(KEYINPUT78), .B(n489), .Z(n503) );
  NAND2_X1 U546 ( .A1(n512), .A2(n503), .ZN(n497) );
  NOR2_X1 U547 ( .A1(n523), .A2(n497), .ZN(n491) );
  XNOR2_X1 U548 ( .A(KEYINPUT34), .B(KEYINPUT108), .ZN(n490) );
  XNOR2_X1 U549 ( .A(n491), .B(n490), .ZN(n492) );
  XOR2_X1 U550 ( .A(G1GAT), .B(n492), .Z(G1324GAT) );
  NOR2_X1 U551 ( .A1(n526), .A2(n497), .ZN(n493) );
  XOR2_X1 U552 ( .A(G8GAT), .B(n493), .Z(G1325GAT) );
  NOR2_X1 U553 ( .A1(n535), .A2(n497), .ZN(n495) );
  XNOR2_X1 U554 ( .A(KEYINPUT109), .B(KEYINPUT35), .ZN(n494) );
  XNOR2_X1 U555 ( .A(n495), .B(n494), .ZN(n496) );
  XOR2_X1 U556 ( .A(G15GAT), .B(n496), .Z(G1326GAT) );
  NOR2_X1 U557 ( .A1(n531), .A2(n497), .ZN(n498) );
  XOR2_X1 U558 ( .A(G22GAT), .B(n498), .Z(G1327GAT) );
  XNOR2_X1 U559 ( .A(G29GAT), .B(KEYINPUT39), .ZN(n506) );
  NOR2_X1 U560 ( .A1(n581), .A2(n499), .ZN(n501) );
  NAND2_X1 U561 ( .A1(n501), .A2(n500), .ZN(n502) );
  NAND2_X1 U562 ( .A1(n503), .A2(n522), .ZN(n504) );
  NOR2_X1 U563 ( .A1(n523), .A2(n509), .ZN(n505) );
  XNOR2_X1 U564 ( .A(n506), .B(n505), .ZN(G1328GAT) );
  NOR2_X1 U565 ( .A1(n509), .A2(n526), .ZN(n507) );
  XOR2_X1 U566 ( .A(G36GAT), .B(n507), .Z(G1329GAT) );
  NOR2_X1 U567 ( .A1(n509), .A2(n535), .ZN(n508) );
  XNOR2_X1 U568 ( .A(G43GAT), .B(n294), .ZN(G1330GAT) );
  NOR2_X1 U569 ( .A1(n509), .A2(n531), .ZN(n510) );
  XOR2_X1 U570 ( .A(G50GAT), .B(n510), .Z(G1331GAT) );
  NOR2_X1 U571 ( .A1(n568), .A2(n511), .ZN(n521) );
  NAND2_X1 U572 ( .A1(n521), .A2(n512), .ZN(n518) );
  NOR2_X1 U573 ( .A1(n523), .A2(n518), .ZN(n514) );
  XNOR2_X1 U574 ( .A(KEYINPUT110), .B(KEYINPUT42), .ZN(n513) );
  XNOR2_X1 U575 ( .A(n514), .B(n513), .ZN(n515) );
  XOR2_X1 U576 ( .A(G57GAT), .B(n515), .Z(G1332GAT) );
  NOR2_X1 U577 ( .A1(n526), .A2(n518), .ZN(n516) );
  XOR2_X1 U578 ( .A(G64GAT), .B(n516), .Z(G1333GAT) );
  NOR2_X1 U579 ( .A1(n535), .A2(n518), .ZN(n517) );
  XOR2_X1 U580 ( .A(G71GAT), .B(n517), .Z(G1334GAT) );
  NOR2_X1 U581 ( .A1(n531), .A2(n518), .ZN(n520) );
  XNOR2_X1 U582 ( .A(G78GAT), .B(KEYINPUT43), .ZN(n519) );
  XNOR2_X1 U583 ( .A(n520), .B(n519), .ZN(G1335GAT) );
  NAND2_X1 U584 ( .A1(n522), .A2(n521), .ZN(n530) );
  NOR2_X1 U585 ( .A1(n523), .A2(n530), .ZN(n525) );
  XNOR2_X1 U586 ( .A(G85GAT), .B(KEYINPUT111), .ZN(n524) );
  XNOR2_X1 U587 ( .A(n525), .B(n524), .ZN(G1336GAT) );
  NOR2_X1 U588 ( .A1(n526), .A2(n530), .ZN(n527) );
  XOR2_X1 U589 ( .A(G92GAT), .B(n527), .Z(G1337GAT) );
  NOR2_X1 U590 ( .A1(n535), .A2(n530), .ZN(n528) );
  XOR2_X1 U591 ( .A(KEYINPUT112), .B(n528), .Z(n529) );
  XNOR2_X1 U592 ( .A(G99GAT), .B(n529), .ZN(G1338GAT) );
  NOR2_X1 U593 ( .A1(n531), .A2(n530), .ZN(n532) );
  XOR2_X1 U594 ( .A(KEYINPUT44), .B(n532), .Z(n533) );
  XNOR2_X1 U595 ( .A(G106GAT), .B(n533), .ZN(G1339GAT) );
  OR2_X1 U596 ( .A1(n535), .A2(n534), .ZN(n536) );
  NOR2_X1 U597 ( .A1(n537), .A2(n536), .ZN(n545) );
  NAND2_X1 U598 ( .A1(n568), .A2(n545), .ZN(n538) );
  XNOR2_X1 U599 ( .A(G113GAT), .B(n538), .ZN(G1340GAT) );
  XOR2_X1 U600 ( .A(G120GAT), .B(KEYINPUT49), .Z(n540) );
  NAND2_X1 U601 ( .A1(n545), .A2(n553), .ZN(n539) );
  XNOR2_X1 U602 ( .A(n540), .B(n539), .ZN(G1341GAT) );
  XNOR2_X1 U603 ( .A(G127GAT), .B(KEYINPUT115), .ZN(n544) );
  XOR2_X1 U604 ( .A(KEYINPUT116), .B(KEYINPUT50), .Z(n542) );
  NAND2_X1 U605 ( .A1(n545), .A2(n577), .ZN(n541) );
  XNOR2_X1 U606 ( .A(n542), .B(n541), .ZN(n543) );
  XNOR2_X1 U607 ( .A(n544), .B(n543), .ZN(G1342GAT) );
  XOR2_X1 U608 ( .A(KEYINPUT117), .B(KEYINPUT51), .Z(n547) );
  NAND2_X1 U609 ( .A1(n545), .A2(n559), .ZN(n546) );
  XNOR2_X1 U610 ( .A(n547), .B(n546), .ZN(n548) );
  XOR2_X1 U611 ( .A(G134GAT), .B(n548), .Z(G1343GAT) );
  NAND2_X1 U612 ( .A1(n566), .A2(n549), .ZN(n550) );
  NOR2_X1 U613 ( .A1(n550), .A2(n534), .ZN(n551) );
  XNOR2_X1 U614 ( .A(n551), .B(KEYINPUT118), .ZN(n560) );
  NAND2_X1 U615 ( .A1(n568), .A2(n560), .ZN(n552) );
  XNOR2_X1 U616 ( .A(G141GAT), .B(n552), .ZN(G1344GAT) );
  XOR2_X1 U617 ( .A(KEYINPUT52), .B(KEYINPUT119), .Z(n555) );
  NAND2_X1 U618 ( .A1(n560), .A2(n553), .ZN(n554) );
  XNOR2_X1 U619 ( .A(n555), .B(n554), .ZN(n557) );
  XOR2_X1 U620 ( .A(G148GAT), .B(KEYINPUT53), .Z(n556) );
  XNOR2_X1 U621 ( .A(n557), .B(n556), .ZN(G1345GAT) );
  NAND2_X1 U622 ( .A1(n560), .A2(n577), .ZN(n558) );
  XNOR2_X1 U623 ( .A(n558), .B(G155GAT), .ZN(G1346GAT) );
  NAND2_X1 U624 ( .A1(n560), .A2(n559), .ZN(n561) );
  XNOR2_X1 U625 ( .A(n561), .B(KEYINPUT120), .ZN(n562) );
  XNOR2_X1 U626 ( .A(G162GAT), .B(n562), .ZN(G1347GAT) );
  NAND2_X1 U627 ( .A1(n568), .A2(n564), .ZN(n563) );
  XNOR2_X1 U628 ( .A(G169GAT), .B(n563), .ZN(G1348GAT) );
  NAND2_X1 U629 ( .A1(n564), .A2(n577), .ZN(n565) );
  XNOR2_X1 U630 ( .A(n565), .B(G183GAT), .ZN(G1350GAT) );
  XOR2_X1 U631 ( .A(KEYINPUT126), .B(KEYINPUT60), .Z(n570) );
  NAND2_X1 U632 ( .A1(n567), .A2(n566), .ZN(n580) );
  INV_X1 U633 ( .A(n580), .ZN(n578) );
  NAND2_X1 U634 ( .A1(n578), .A2(n568), .ZN(n569) );
  XNOR2_X1 U635 ( .A(n570), .B(n569), .ZN(n571) );
  XOR2_X1 U636 ( .A(n571), .B(KEYINPUT59), .Z(n573) );
  XNOR2_X1 U637 ( .A(G197GAT), .B(KEYINPUT125), .ZN(n572) );
  XNOR2_X1 U638 ( .A(n573), .B(n572), .ZN(G1352GAT) );
  XOR2_X1 U639 ( .A(KEYINPUT127), .B(KEYINPUT61), .Z(n575) );
  OR2_X1 U640 ( .A1(n580), .A2(n369), .ZN(n574) );
  XNOR2_X1 U641 ( .A(n575), .B(n574), .ZN(n576) );
  XOR2_X1 U642 ( .A(G204GAT), .B(n576), .Z(G1353GAT) );
  NAND2_X1 U643 ( .A1(n578), .A2(n577), .ZN(n579) );
  XNOR2_X1 U644 ( .A(n579), .B(G211GAT), .ZN(G1354GAT) );
  NOR2_X1 U645 ( .A1(n581), .A2(n580), .ZN(n582) );
  XOR2_X1 U646 ( .A(KEYINPUT62), .B(n582), .Z(n583) );
  XNOR2_X1 U647 ( .A(G218GAT), .B(n583), .ZN(G1355GAT) );
endmodule

