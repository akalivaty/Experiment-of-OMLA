//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 0 0 0 1 1 0 0 0 1 0 1 0 1 1 1 1 0 0 1 1 0 0 0 0 1 1 0 1 1 1 0 1 0 1 0 1 0 0 1 1 0 0 0 0 0 1 1 0 0 1 0 0 0 1 0 1 1 0 0 0 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:39:03 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n205, new_n206, new_n207, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n241, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1108, new_n1109, new_n1110, new_n1111, new_n1112,
    new_n1113, new_n1114, new_n1115, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1186, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1251, new_n1252,
    new_n1253, new_n1254, new_n1255, new_n1256, new_n1257, new_n1258,
    new_n1259, new_n1260, new_n1261, new_n1262, new_n1263, new_n1264,
    new_n1265, new_n1266, new_n1267, new_n1268, new_n1269, new_n1270,
    new_n1271, new_n1272, new_n1273, new_n1275, new_n1276, new_n1277,
    new_n1278, new_n1279, new_n1280, new_n1281, new_n1282, new_n1283,
    new_n1284, new_n1285, new_n1286, new_n1287, new_n1288, new_n1289,
    new_n1290, new_n1291, new_n1292, new_n1293, new_n1294, new_n1295,
    new_n1297, new_n1298, new_n1299, new_n1300, new_n1301, new_n1302,
    new_n1303, new_n1304, new_n1305, new_n1306, new_n1307, new_n1308,
    new_n1310, new_n1311, new_n1312, new_n1313, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1346,
    new_n1347, new_n1348, new_n1349, new_n1350, new_n1351, new_n1352,
    new_n1353, new_n1354, new_n1355, new_n1356, new_n1357, new_n1358,
    new_n1359, new_n1360, new_n1361, new_n1362, new_n1363, new_n1364,
    new_n1365, new_n1366, new_n1367, new_n1369, new_n1370, new_n1371,
    new_n1372;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  INV_X1    g0004(.A(G97), .ZN(new_n205));
  INV_X1    g0005(.A(G107), .ZN(new_n206));
  NAND2_X1  g0006(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  NAND2_X1  g0007(.A1(new_n207), .A2(G87), .ZN(G355));
  INV_X1    g0008(.A(G1), .ZN(new_n209));
  INV_X1    g0009(.A(G20), .ZN(new_n210));
  NOR2_X1   g0010(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  INV_X1    g0011(.A(new_n211), .ZN(new_n212));
  NOR2_X1   g0012(.A1(new_n212), .A2(G13), .ZN(new_n213));
  OAI211_X1 g0013(.A(new_n213), .B(G250), .C1(G257), .C2(G264), .ZN(new_n214));
  XNOR2_X1  g0014(.A(new_n214), .B(KEYINPUT0), .ZN(new_n215));
  INV_X1    g0015(.A(new_n201), .ZN(new_n216));
  NAND2_X1  g0016(.A1(new_n216), .A2(G50), .ZN(new_n217));
  INV_X1    g0017(.A(new_n217), .ZN(new_n218));
  NAND2_X1  g0018(.A1(G1), .A2(G13), .ZN(new_n219));
  INV_X1    g0019(.A(new_n219), .ZN(new_n220));
  NAND3_X1  g0020(.A1(new_n218), .A2(G20), .A3(new_n220), .ZN(new_n221));
  XNOR2_X1  g0021(.A(KEYINPUT64), .B(G68), .ZN(new_n222));
  INV_X1    g0022(.A(G238), .ZN(new_n223));
  NOR2_X1   g0023(.A1(new_n222), .A2(new_n223), .ZN(new_n224));
  AOI22_X1  g0024(.A1(G107), .A2(G264), .B1(G116), .B2(G270), .ZN(new_n225));
  AOI22_X1  g0025(.A1(G50), .A2(G226), .B1(G77), .B2(G244), .ZN(new_n226));
  AOI22_X1  g0026(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n227));
  NAND2_X1  g0027(.A1(G58), .A2(G232), .ZN(new_n228));
  NAND4_X1  g0028(.A1(new_n225), .A2(new_n226), .A3(new_n227), .A4(new_n228), .ZN(new_n229));
  OAI21_X1  g0029(.A(new_n212), .B1(new_n224), .B2(new_n229), .ZN(new_n230));
  OAI211_X1 g0030(.A(new_n215), .B(new_n221), .C1(KEYINPUT1), .C2(new_n230), .ZN(new_n231));
  AOI21_X1  g0031(.A(new_n231), .B1(KEYINPUT1), .B2(new_n230), .ZN(G361));
  XNOR2_X1  g0032(.A(G238), .B(G244), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n233), .B(G232), .ZN(new_n234));
  XNOR2_X1  g0034(.A(KEYINPUT2), .B(G226), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XOR2_X1   g0036(.A(G264), .B(G270), .Z(new_n237));
  XNOR2_X1  g0037(.A(G250), .B(G257), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n236), .B(new_n239), .ZN(G358));
  XOR2_X1   g0040(.A(G87), .B(G97), .Z(new_n241));
  XNOR2_X1  g0041(.A(new_n241), .B(KEYINPUT65), .ZN(new_n242));
  XNOR2_X1  g0042(.A(G107), .B(G116), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XNOR2_X1  g0044(.A(G50), .B(G68), .ZN(new_n245));
  XNOR2_X1  g0045(.A(G58), .B(G77), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n245), .B(new_n246), .ZN(new_n247));
  XOR2_X1   g0047(.A(new_n244), .B(new_n247), .Z(G351));
  AND2_X1   g0048(.A1(KEYINPUT3), .A2(G33), .ZN(new_n249));
  NOR2_X1   g0049(.A1(KEYINPUT3), .A2(G33), .ZN(new_n250));
  NOR2_X1   g0050(.A1(new_n249), .A2(new_n250), .ZN(new_n251));
  NOR2_X1   g0051(.A1(new_n251), .A2(G1698), .ZN(new_n252));
  NAND2_X1  g0052(.A1(new_n252), .A2(G222), .ZN(new_n253));
  INV_X1    g0053(.A(G77), .ZN(new_n254));
  XNOR2_X1  g0054(.A(KEYINPUT3), .B(G33), .ZN(new_n255));
  INV_X1    g0055(.A(G223), .ZN(new_n256));
  NAND2_X1  g0056(.A1(new_n255), .A2(G1698), .ZN(new_n257));
  OAI221_X1 g0057(.A(new_n253), .B1(new_n254), .B2(new_n255), .C1(new_n256), .C2(new_n257), .ZN(new_n258));
  NAND2_X1  g0058(.A1(G33), .A2(G41), .ZN(new_n259));
  NAND3_X1  g0059(.A1(new_n259), .A2(G1), .A3(G13), .ZN(new_n260));
  INV_X1    g0060(.A(new_n260), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n258), .A2(new_n261), .ZN(new_n262));
  INV_X1    g0062(.A(G41), .ZN(new_n263));
  INV_X1    g0063(.A(G45), .ZN(new_n264));
  AOI21_X1  g0064(.A(G1), .B1(new_n263), .B2(new_n264), .ZN(new_n265));
  NAND3_X1  g0065(.A1(new_n265), .A2(new_n260), .A3(G274), .ZN(new_n266));
  INV_X1    g0066(.A(KEYINPUT66), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n266), .A2(new_n267), .ZN(new_n268));
  INV_X1    g0068(.A(G274), .ZN(new_n269));
  AOI21_X1  g0069(.A(new_n269), .B1(new_n220), .B2(new_n259), .ZN(new_n270));
  NAND3_X1  g0070(.A1(new_n270), .A2(KEYINPUT66), .A3(new_n265), .ZN(new_n271));
  NOR2_X1   g0071(.A1(new_n261), .A2(new_n265), .ZN(new_n272));
  AOI22_X1  g0072(.A1(new_n268), .A2(new_n271), .B1(new_n272), .B2(G226), .ZN(new_n273));
  NAND2_X1  g0073(.A1(new_n262), .A2(new_n273), .ZN(new_n274));
  INV_X1    g0074(.A(new_n274), .ZN(new_n275));
  NOR2_X1   g0075(.A1(new_n275), .A2(G169), .ZN(new_n276));
  INV_X1    g0076(.A(G13), .ZN(new_n277));
  NOR3_X1   g0077(.A1(new_n277), .A2(new_n210), .A3(G1), .ZN(new_n278));
  INV_X1    g0078(.A(new_n278), .ZN(new_n279));
  NAND2_X1  g0079(.A1(new_n279), .A2(new_n202), .ZN(new_n280));
  NAND3_X1  g0080(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n281));
  NAND2_X1  g0081(.A1(new_n281), .A2(new_n219), .ZN(new_n282));
  AOI21_X1  g0082(.A(new_n282), .B1(new_n209), .B2(G20), .ZN(new_n283));
  OAI21_X1  g0083(.A(new_n280), .B1(new_n283), .B2(new_n202), .ZN(new_n284));
  XNOR2_X1  g0084(.A(new_n284), .B(KEYINPUT68), .ZN(new_n285));
  INV_X1    g0085(.A(new_n282), .ZN(new_n286));
  NOR2_X1   g0086(.A1(KEYINPUT8), .A2(G58), .ZN(new_n287));
  INV_X1    g0087(.A(G58), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n288), .A2(KEYINPUT67), .ZN(new_n289));
  INV_X1    g0089(.A(KEYINPUT67), .ZN(new_n290));
  NAND2_X1  g0090(.A1(new_n290), .A2(G58), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n289), .A2(new_n291), .ZN(new_n292));
  AOI21_X1  g0092(.A(new_n287), .B1(new_n292), .B2(KEYINPUT8), .ZN(new_n293));
  NAND3_X1  g0093(.A1(new_n293), .A2(new_n210), .A3(G33), .ZN(new_n294));
  NOR2_X1   g0094(.A1(G20), .A2(G33), .ZN(new_n295));
  AOI22_X1  g0095(.A1(new_n203), .A2(G20), .B1(G150), .B2(new_n295), .ZN(new_n296));
  AOI21_X1  g0096(.A(new_n286), .B1(new_n294), .B2(new_n296), .ZN(new_n297));
  NOR2_X1   g0097(.A1(new_n285), .A2(new_n297), .ZN(new_n298));
  OAI21_X1  g0098(.A(KEYINPUT69), .B1(new_n276), .B2(new_n298), .ZN(new_n299));
  INV_X1    g0099(.A(new_n298), .ZN(new_n300));
  INV_X1    g0100(.A(KEYINPUT69), .ZN(new_n301));
  OAI211_X1 g0101(.A(new_n300), .B(new_n301), .C1(new_n275), .C2(G169), .ZN(new_n302));
  INV_X1    g0102(.A(G179), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n275), .A2(new_n303), .ZN(new_n304));
  AND3_X1   g0104(.A1(new_n299), .A2(new_n302), .A3(new_n304), .ZN(new_n305));
  INV_X1    g0105(.A(G190), .ZN(new_n306));
  NOR2_X1   g0106(.A1(new_n274), .A2(new_n306), .ZN(new_n307));
  AOI21_X1  g0107(.A(new_n307), .B1(G200), .B2(new_n274), .ZN(new_n308));
  INV_X1    g0108(.A(KEYINPUT9), .ZN(new_n309));
  XNOR2_X1  g0109(.A(new_n298), .B(new_n309), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n308), .A2(new_n310), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n311), .A2(KEYINPUT10), .ZN(new_n312));
  INV_X1    g0112(.A(KEYINPUT10), .ZN(new_n313));
  NAND3_X1  g0113(.A1(new_n308), .A2(new_n310), .A3(new_n313), .ZN(new_n314));
  AOI21_X1  g0114(.A(new_n305), .B1(new_n312), .B2(new_n314), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n295), .A2(G50), .ZN(new_n316));
  XNOR2_X1  g0116(.A(new_n316), .B(KEYINPUT71), .ZN(new_n317));
  INV_X1    g0117(.A(G68), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n318), .A2(KEYINPUT64), .ZN(new_n319));
  INV_X1    g0119(.A(KEYINPUT64), .ZN(new_n320));
  NAND2_X1  g0120(.A1(new_n320), .A2(G68), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n319), .A2(new_n321), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n210), .A2(G33), .ZN(new_n323));
  OAI22_X1  g0123(.A1(new_n322), .A2(new_n210), .B1(new_n254), .B2(new_n323), .ZN(new_n324));
  OAI21_X1  g0124(.A(new_n282), .B1(new_n317), .B2(new_n324), .ZN(new_n325));
  XNOR2_X1  g0125(.A(new_n325), .B(KEYINPUT11), .ZN(new_n326));
  INV_X1    g0126(.A(KEYINPUT72), .ZN(new_n327));
  INV_X1    g0127(.A(new_n283), .ZN(new_n328));
  OAI21_X1  g0128(.A(new_n327), .B1(new_n328), .B2(new_n318), .ZN(new_n329));
  NAND3_X1  g0129(.A1(new_n283), .A2(KEYINPUT72), .A3(G68), .ZN(new_n330));
  INV_X1    g0130(.A(KEYINPUT12), .ZN(new_n331));
  AOI21_X1  g0131(.A(new_n331), .B1(new_n222), .B2(new_n278), .ZN(new_n332));
  NAND3_X1  g0132(.A1(new_n278), .A2(new_n331), .A3(new_n318), .ZN(new_n333));
  AOI21_X1  g0133(.A(new_n332), .B1(KEYINPUT73), .B2(new_n333), .ZN(new_n334));
  OR2_X1    g0134(.A1(new_n333), .A2(KEYINPUT73), .ZN(new_n335));
  AOI22_X1  g0135(.A1(new_n329), .A2(new_n330), .B1(new_n334), .B2(new_n335), .ZN(new_n336));
  AND2_X1   g0136(.A1(new_n326), .A2(new_n336), .ZN(new_n337));
  INV_X1    g0137(.A(new_n337), .ZN(new_n338));
  INV_X1    g0138(.A(KEYINPUT14), .ZN(new_n339));
  OAI211_X1 g0139(.A(G232), .B(G1698), .C1(new_n249), .C2(new_n250), .ZN(new_n340));
  XNOR2_X1  g0140(.A(new_n340), .B(KEYINPUT70), .ZN(new_n341));
  AOI22_X1  g0141(.A1(new_n252), .A2(G226), .B1(G33), .B2(G97), .ZN(new_n342));
  AOI21_X1  g0142(.A(new_n260), .B1(new_n341), .B2(new_n342), .ZN(new_n343));
  NAND2_X1  g0143(.A1(new_n268), .A2(new_n271), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n272), .A2(G238), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n344), .A2(new_n345), .ZN(new_n346));
  NOR3_X1   g0146(.A1(new_n343), .A2(KEYINPUT13), .A3(new_n346), .ZN(new_n347));
  INV_X1    g0147(.A(KEYINPUT13), .ZN(new_n348));
  INV_X1    g0148(.A(KEYINPUT70), .ZN(new_n349));
  XNOR2_X1  g0149(.A(new_n340), .B(new_n349), .ZN(new_n350));
  NAND2_X1  g0150(.A1(G33), .A2(G97), .ZN(new_n351));
  INV_X1    g0151(.A(G1698), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n255), .A2(new_n352), .ZN(new_n353));
  INV_X1    g0153(.A(G226), .ZN(new_n354));
  OAI21_X1  g0154(.A(new_n351), .B1(new_n353), .B2(new_n354), .ZN(new_n355));
  OAI21_X1  g0155(.A(new_n261), .B1(new_n350), .B2(new_n355), .ZN(new_n356));
  AND2_X1   g0156(.A1(new_n344), .A2(new_n345), .ZN(new_n357));
  AOI21_X1  g0157(.A(new_n348), .B1(new_n356), .B2(new_n357), .ZN(new_n358));
  OAI211_X1 g0158(.A(new_n339), .B(G169), .C1(new_n347), .C2(new_n358), .ZN(new_n359));
  OAI21_X1  g0159(.A(KEYINPUT13), .B1(new_n343), .B2(new_n346), .ZN(new_n360));
  NAND3_X1  g0160(.A1(new_n356), .A2(new_n357), .A3(new_n348), .ZN(new_n361));
  NAND3_X1  g0161(.A1(new_n360), .A2(G179), .A3(new_n361), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n359), .A2(new_n362), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n360), .A2(new_n361), .ZN(new_n364));
  AOI21_X1  g0164(.A(new_n339), .B1(new_n364), .B2(G169), .ZN(new_n365));
  OAI21_X1  g0165(.A(new_n338), .B1(new_n363), .B2(new_n365), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n252), .A2(G232), .ZN(new_n367));
  OAI221_X1 g0167(.A(new_n367), .B1(new_n206), .B2(new_n255), .C1(new_n223), .C2(new_n257), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n368), .A2(new_n261), .ZN(new_n369));
  AOI22_X1  g0169(.A1(new_n268), .A2(new_n271), .B1(new_n272), .B2(G244), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n369), .A2(new_n370), .ZN(new_n371));
  NOR2_X1   g0171(.A1(new_n371), .A2(G179), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n278), .A2(new_n254), .ZN(new_n373));
  OAI21_X1  g0173(.A(new_n373), .B1(new_n328), .B2(new_n254), .ZN(new_n374));
  XOR2_X1   g0174(.A(KEYINPUT8), .B(G58), .Z(new_n375));
  AOI22_X1  g0175(.A1(new_n375), .A2(new_n295), .B1(G20), .B2(G77), .ZN(new_n376));
  XNOR2_X1  g0176(.A(KEYINPUT15), .B(G87), .ZN(new_n377));
  OAI21_X1  g0177(.A(new_n376), .B1(new_n323), .B2(new_n377), .ZN(new_n378));
  AOI21_X1  g0178(.A(new_n374), .B1(new_n282), .B2(new_n378), .ZN(new_n379));
  AOI21_X1  g0179(.A(G169), .B1(new_n369), .B2(new_n370), .ZN(new_n380));
  NOR3_X1   g0180(.A1(new_n372), .A2(new_n379), .A3(new_n380), .ZN(new_n381));
  INV_X1    g0181(.A(new_n381), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n371), .A2(G200), .ZN(new_n383));
  OAI211_X1 g0183(.A(new_n383), .B(new_n379), .C1(new_n306), .C2(new_n371), .ZN(new_n384));
  OAI21_X1  g0184(.A(G200), .B1(new_n347), .B2(new_n358), .ZN(new_n385));
  NAND3_X1  g0185(.A1(new_n360), .A2(G190), .A3(new_n361), .ZN(new_n386));
  NAND3_X1  g0186(.A1(new_n385), .A2(new_n337), .A3(new_n386), .ZN(new_n387));
  AND3_X1   g0187(.A1(new_n382), .A2(new_n384), .A3(new_n387), .ZN(new_n388));
  AND3_X1   g0188(.A1(new_n315), .A2(new_n366), .A3(new_n388), .ZN(new_n389));
  INV_X1    g0189(.A(KEYINPUT17), .ZN(new_n390));
  NAND2_X1  g0190(.A1(new_n328), .A2(new_n293), .ZN(new_n391));
  OAI21_X1  g0191(.A(new_n391), .B1(new_n278), .B2(new_n293), .ZN(new_n392));
  INV_X1    g0192(.A(new_n392), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n295), .A2(G159), .ZN(new_n394));
  INV_X1    g0194(.A(new_n394), .ZN(new_n395));
  XNOR2_X1  g0195(.A(KEYINPUT67), .B(G58), .ZN(new_n396));
  OAI21_X1  g0196(.A(new_n216), .B1(new_n222), .B2(new_n396), .ZN(new_n397));
  AOI21_X1  g0197(.A(new_n395), .B1(new_n397), .B2(G20), .ZN(new_n398));
  AOI21_X1  g0198(.A(G20), .B1(KEYINPUT3), .B2(G33), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n399), .A2(KEYINPUT7), .ZN(new_n400));
  AND2_X1   g0200(.A1(KEYINPUT74), .A2(G33), .ZN(new_n401));
  NOR2_X1   g0201(.A1(KEYINPUT74), .A2(G33), .ZN(new_n402));
  NOR2_X1   g0202(.A1(new_n401), .A2(new_n402), .ZN(new_n403));
  INV_X1    g0203(.A(KEYINPUT3), .ZN(new_n404));
  AOI21_X1  g0204(.A(new_n400), .B1(new_n403), .B2(new_n404), .ZN(new_n405));
  INV_X1    g0205(.A(new_n250), .ZN(new_n406));
  AOI21_X1  g0206(.A(KEYINPUT7), .B1(new_n406), .B2(new_n399), .ZN(new_n407));
  OAI21_X1  g0207(.A(new_n322), .B1(new_n405), .B2(new_n407), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n398), .A2(new_n408), .ZN(new_n409));
  INV_X1    g0209(.A(KEYINPUT16), .ZN(new_n410));
  AOI21_X1  g0210(.A(new_n286), .B1(new_n409), .B2(new_n410), .ZN(new_n411));
  INV_X1    g0211(.A(KEYINPUT7), .ZN(new_n412));
  INV_X1    g0212(.A(KEYINPUT74), .ZN(new_n413));
  INV_X1    g0213(.A(G33), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n413), .A2(new_n414), .ZN(new_n415));
  NAND2_X1  g0215(.A1(KEYINPUT74), .A2(G33), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n415), .A2(new_n416), .ZN(new_n417));
  AOI21_X1  g0217(.A(new_n250), .B1(new_n417), .B2(KEYINPUT3), .ZN(new_n418));
  AOI21_X1  g0218(.A(new_n412), .B1(new_n418), .B2(new_n210), .ZN(new_n419));
  OAI21_X1  g0219(.A(KEYINPUT3), .B1(new_n401), .B2(new_n402), .ZN(new_n420));
  NAND4_X1  g0220(.A1(new_n420), .A2(new_n412), .A3(new_n210), .A4(new_n406), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n421), .A2(G68), .ZN(new_n422));
  OAI211_X1 g0222(.A(new_n398), .B(KEYINPUT16), .C1(new_n419), .C2(new_n422), .ZN(new_n423));
  AOI21_X1  g0223(.A(new_n393), .B1(new_n411), .B2(new_n423), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n272), .A2(G232), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n344), .A2(new_n425), .ZN(new_n426));
  AOI21_X1  g0226(.A(new_n352), .B1(new_n420), .B2(new_n406), .ZN(new_n427));
  AOI22_X1  g0227(.A1(new_n427), .A2(G226), .B1(G33), .B2(G87), .ZN(new_n428));
  AOI21_X1  g0228(.A(new_n404), .B1(new_n415), .B2(new_n416), .ZN(new_n429));
  OAI211_X1 g0229(.A(G223), .B(new_n352), .C1(new_n429), .C2(new_n250), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n430), .A2(KEYINPUT75), .ZN(new_n431));
  AOI21_X1  g0231(.A(G1698), .B1(new_n420), .B2(new_n406), .ZN(new_n432));
  INV_X1    g0232(.A(KEYINPUT75), .ZN(new_n433));
  NAND3_X1  g0233(.A1(new_n432), .A2(new_n433), .A3(G223), .ZN(new_n434));
  NAND3_X1  g0234(.A1(new_n428), .A2(new_n431), .A3(new_n434), .ZN(new_n435));
  AOI21_X1  g0235(.A(new_n426), .B1(new_n435), .B2(new_n261), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n436), .A2(G190), .ZN(new_n437));
  NAND2_X1  g0237(.A1(new_n424), .A2(new_n437), .ZN(new_n438));
  INV_X1    g0238(.A(G200), .ZN(new_n439));
  NOR2_X1   g0239(.A1(new_n436), .A2(new_n439), .ZN(new_n440));
  OAI211_X1 g0240(.A(KEYINPUT76), .B(new_n390), .C1(new_n438), .C2(new_n440), .ZN(new_n441));
  OAI211_X1 g0241(.A(KEYINPUT7), .B(new_n399), .C1(new_n417), .C2(KEYINPUT3), .ZN(new_n442));
  INV_X1    g0242(.A(new_n407), .ZN(new_n443));
  AOI21_X1  g0243(.A(new_n222), .B1(new_n442), .B2(new_n443), .ZN(new_n444));
  AOI21_X1  g0244(.A(new_n201), .B1(new_n322), .B2(new_n292), .ZN(new_n445));
  OAI21_X1  g0245(.A(new_n394), .B1(new_n445), .B2(new_n210), .ZN(new_n446));
  OAI21_X1  g0246(.A(new_n410), .B1(new_n444), .B2(new_n446), .ZN(new_n447));
  NAND3_X1  g0247(.A1(new_n447), .A2(new_n423), .A3(new_n282), .ZN(new_n448));
  NAND2_X1  g0248(.A1(new_n448), .A2(new_n392), .ZN(new_n449));
  AOI211_X1 g0249(.A(new_n306), .B(new_n426), .C1(new_n435), .C2(new_n261), .ZN(new_n450));
  NOR2_X1   g0250(.A1(new_n449), .A2(new_n450), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n390), .A2(KEYINPUT76), .ZN(new_n452));
  OR2_X1    g0252(.A1(new_n390), .A2(KEYINPUT76), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n435), .A2(new_n261), .ZN(new_n454));
  INV_X1    g0254(.A(new_n426), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n454), .A2(new_n455), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n456), .A2(G200), .ZN(new_n457));
  NAND4_X1  g0257(.A1(new_n451), .A2(new_n452), .A3(new_n453), .A4(new_n457), .ZN(new_n458));
  INV_X1    g0258(.A(G169), .ZN(new_n459));
  NOR2_X1   g0259(.A1(new_n436), .A2(new_n459), .ZN(new_n460));
  AOI211_X1 g0260(.A(new_n303), .B(new_n426), .C1(new_n435), .C2(new_n261), .ZN(new_n461));
  OAI21_X1  g0261(.A(new_n449), .B1(new_n460), .B2(new_n461), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n462), .A2(KEYINPUT18), .ZN(new_n463));
  INV_X1    g0263(.A(KEYINPUT18), .ZN(new_n464));
  OAI211_X1 g0264(.A(new_n464), .B(new_n449), .C1(new_n460), .C2(new_n461), .ZN(new_n465));
  NAND4_X1  g0265(.A1(new_n441), .A2(new_n458), .A3(new_n463), .A4(new_n465), .ZN(new_n466));
  INV_X1    g0266(.A(new_n466), .ZN(new_n467));
  OR2_X1    g0267(.A1(new_n467), .A2(KEYINPUT77), .ZN(new_n468));
  NAND2_X1  g0268(.A1(new_n467), .A2(KEYINPUT77), .ZN(new_n469));
  NAND3_X1  g0269(.A1(new_n389), .A2(new_n468), .A3(new_n469), .ZN(new_n470));
  INV_X1    g0270(.A(new_n470), .ZN(new_n471));
  NOR2_X1   g0271(.A1(new_n264), .A2(G1), .ZN(new_n472));
  XNOR2_X1  g0272(.A(KEYINPUT5), .B(G41), .ZN(new_n473));
  AOI21_X1  g0273(.A(new_n261), .B1(new_n472), .B2(new_n473), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n474), .A2(G257), .ZN(new_n475));
  NAND3_X1  g0275(.A1(new_n270), .A2(new_n472), .A3(new_n473), .ZN(new_n476));
  INV_X1    g0276(.A(KEYINPUT4), .ZN(new_n477));
  INV_X1    g0277(.A(G244), .ZN(new_n478));
  NOR2_X1   g0278(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  OAI211_X1 g0279(.A(new_n479), .B(new_n352), .C1(new_n250), .C2(new_n249), .ZN(new_n480));
  NAND2_X1  g0280(.A1(G33), .A2(G283), .ZN(new_n481));
  OAI211_X1 g0281(.A(G250), .B(G1698), .C1(new_n249), .C2(new_n250), .ZN(new_n482));
  NAND3_X1  g0282(.A1(new_n480), .A2(new_n481), .A3(new_n482), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n420), .A2(new_n406), .ZN(new_n484));
  NAND3_X1  g0284(.A1(new_n484), .A2(G244), .A3(new_n352), .ZN(new_n485));
  AOI21_X1  g0285(.A(new_n483), .B1(new_n485), .B2(new_n477), .ZN(new_n486));
  OAI211_X1 g0286(.A(new_n475), .B(new_n476), .C1(new_n486), .C2(new_n260), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n487), .A2(G200), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n278), .A2(new_n205), .ZN(new_n489));
  OAI211_X1 g0289(.A(new_n279), .B(new_n286), .C1(G1), .C2(new_n414), .ZN(new_n490));
  OAI21_X1  g0290(.A(new_n489), .B1(new_n490), .B2(new_n205), .ZN(new_n491));
  OAI21_X1  g0291(.A(G107), .B1(new_n405), .B2(new_n407), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n295), .A2(G77), .ZN(new_n493));
  NAND2_X1  g0293(.A1(G97), .A2(G107), .ZN(new_n494));
  AOI21_X1  g0294(.A(KEYINPUT6), .B1(new_n207), .B2(new_n494), .ZN(new_n495));
  AND3_X1   g0295(.A1(new_n206), .A2(KEYINPUT6), .A3(G97), .ZN(new_n496));
  OAI21_X1  g0296(.A(G20), .B1(new_n495), .B2(new_n496), .ZN(new_n497));
  NAND3_X1  g0297(.A1(new_n492), .A2(new_n493), .A3(new_n497), .ZN(new_n498));
  AOI21_X1  g0298(.A(new_n491), .B1(new_n498), .B2(new_n282), .ZN(new_n499));
  OAI211_X1 g0299(.A(new_n488), .B(new_n499), .C1(new_n306), .C2(new_n487), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n487), .A2(new_n459), .ZN(new_n501));
  INV_X1    g0301(.A(new_n499), .ZN(new_n502));
  AOI21_X1  g0302(.A(KEYINPUT4), .B1(new_n432), .B2(G244), .ZN(new_n503));
  OAI21_X1  g0303(.A(new_n261), .B1(new_n503), .B2(new_n483), .ZN(new_n504));
  NAND4_X1  g0304(.A1(new_n504), .A2(new_n303), .A3(new_n475), .A4(new_n476), .ZN(new_n505));
  NAND3_X1  g0305(.A1(new_n501), .A2(new_n502), .A3(new_n505), .ZN(new_n506));
  AND2_X1   g0306(.A1(new_n500), .A2(new_n506), .ZN(new_n507));
  INV_X1    g0307(.A(KEYINPUT79), .ZN(new_n508));
  NAND3_X1  g0308(.A1(new_n484), .A2(G244), .A3(G1698), .ZN(new_n509));
  INV_X1    g0309(.A(G116), .ZN(new_n510));
  NOR2_X1   g0310(.A1(new_n403), .A2(new_n510), .ZN(new_n511));
  INV_X1    g0311(.A(new_n511), .ZN(new_n512));
  OAI211_X1 g0312(.A(G238), .B(new_n352), .C1(new_n429), .C2(new_n250), .ZN(new_n513));
  NAND3_X1  g0313(.A1(new_n509), .A2(new_n512), .A3(new_n513), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n514), .A2(new_n261), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n270), .A2(new_n472), .ZN(new_n516));
  INV_X1    g0316(.A(G250), .ZN(new_n517));
  AOI21_X1  g0317(.A(new_n517), .B1(new_n209), .B2(G45), .ZN(new_n518));
  INV_X1    g0318(.A(KEYINPUT78), .ZN(new_n519));
  NAND3_X1  g0319(.A1(new_n518), .A2(new_n260), .A3(new_n519), .ZN(new_n520));
  INV_X1    g0320(.A(new_n520), .ZN(new_n521));
  AOI21_X1  g0321(.A(new_n519), .B1(new_n518), .B2(new_n260), .ZN(new_n522));
  OAI21_X1  g0322(.A(new_n516), .B1(new_n521), .B2(new_n522), .ZN(new_n523));
  INV_X1    g0323(.A(new_n523), .ZN(new_n524));
  NAND3_X1  g0324(.A1(new_n515), .A2(G190), .A3(new_n524), .ZN(new_n525));
  NOR3_X1   g0325(.A1(G87), .A2(G97), .A3(G107), .ZN(new_n526));
  AOI21_X1  g0326(.A(new_n526), .B1(new_n210), .B2(new_n351), .ZN(new_n527));
  INV_X1    g0327(.A(KEYINPUT19), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n528), .A2(G97), .ZN(new_n529));
  OAI22_X1  g0329(.A1(new_n527), .A2(new_n528), .B1(new_n323), .B2(new_n529), .ZN(new_n530));
  NAND3_X1  g0330(.A1(new_n484), .A2(new_n210), .A3(G68), .ZN(new_n531));
  AOI21_X1  g0331(.A(new_n286), .B1(new_n530), .B2(new_n531), .ZN(new_n532));
  INV_X1    g0332(.A(new_n377), .ZN(new_n533));
  NOR2_X1   g0333(.A1(new_n533), .A2(new_n279), .ZN(new_n534));
  INV_X1    g0334(.A(G87), .ZN(new_n535));
  NOR2_X1   g0335(.A1(new_n490), .A2(new_n535), .ZN(new_n536));
  NOR3_X1   g0336(.A1(new_n532), .A2(new_n534), .A3(new_n536), .ZN(new_n537));
  AOI21_X1  g0337(.A(new_n523), .B1(new_n514), .B2(new_n261), .ZN(new_n538));
  OAI211_X1 g0338(.A(new_n525), .B(new_n537), .C1(new_n439), .C2(new_n538), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n538), .A2(new_n303), .ZN(new_n540));
  AOI21_X1  g0340(.A(new_n511), .B1(new_n432), .B2(G238), .ZN(new_n541));
  AOI21_X1  g0341(.A(new_n260), .B1(new_n541), .B2(new_n509), .ZN(new_n542));
  OAI21_X1  g0342(.A(new_n459), .B1(new_n542), .B2(new_n523), .ZN(new_n543));
  INV_X1    g0343(.A(new_n534), .ZN(new_n544));
  INV_X1    g0344(.A(new_n490), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n545), .A2(new_n533), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n530), .A2(new_n531), .ZN(new_n547));
  INV_X1    g0347(.A(new_n547), .ZN(new_n548));
  OAI211_X1 g0348(.A(new_n544), .B(new_n546), .C1(new_n548), .C2(new_n286), .ZN(new_n549));
  NAND3_X1  g0349(.A1(new_n540), .A2(new_n543), .A3(new_n549), .ZN(new_n550));
  AND2_X1   g0350(.A1(new_n539), .A2(new_n550), .ZN(new_n551));
  NAND3_X1  g0351(.A1(new_n507), .A2(new_n508), .A3(new_n551), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n500), .A2(new_n506), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n539), .A2(new_n550), .ZN(new_n554));
  OAI21_X1  g0354(.A(KEYINPUT79), .B1(new_n553), .B2(new_n554), .ZN(new_n555));
  XNOR2_X1  g0355(.A(KEYINPUT81), .B(KEYINPUT24), .ZN(new_n556));
  NAND4_X1  g0356(.A1(new_n484), .A2(KEYINPUT22), .A3(new_n210), .A4(G87), .ZN(new_n557));
  INV_X1    g0357(.A(new_n557), .ZN(new_n558));
  INV_X1    g0358(.A(KEYINPUT22), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n210), .A2(G87), .ZN(new_n560));
  OAI21_X1  g0360(.A(new_n559), .B1(new_n251), .B2(new_n560), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n206), .A2(G20), .ZN(new_n562));
  INV_X1    g0362(.A(KEYINPUT23), .ZN(new_n563));
  XNOR2_X1  g0363(.A(new_n562), .B(new_n563), .ZN(new_n564));
  NAND3_X1  g0364(.A1(new_n417), .A2(new_n210), .A3(G116), .ZN(new_n565));
  NAND3_X1  g0365(.A1(new_n561), .A2(new_n564), .A3(new_n565), .ZN(new_n566));
  OAI21_X1  g0366(.A(new_n556), .B1(new_n558), .B2(new_n566), .ZN(new_n567));
  AND2_X1   g0367(.A1(new_n564), .A2(new_n565), .ZN(new_n568));
  INV_X1    g0368(.A(new_n556), .ZN(new_n569));
  NAND4_X1  g0369(.A1(new_n568), .A2(new_n557), .A3(new_n561), .A4(new_n569), .ZN(new_n570));
  AOI21_X1  g0370(.A(new_n286), .B1(new_n567), .B2(new_n570), .ZN(new_n571));
  AND2_X1   g0371(.A1(KEYINPUT82), .A2(KEYINPUT25), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n278), .A2(new_n206), .ZN(new_n573));
  NOR2_X1   g0373(.A1(KEYINPUT82), .A2(KEYINPUT25), .ZN(new_n574));
  AOI21_X1  g0374(.A(new_n572), .B1(new_n573), .B2(new_n574), .ZN(new_n575));
  OAI21_X1  g0375(.A(new_n575), .B1(new_n574), .B2(new_n573), .ZN(new_n576));
  OAI21_X1  g0376(.A(new_n576), .B1(new_n206), .B2(new_n490), .ZN(new_n577));
  NOR2_X1   g0377(.A1(new_n571), .A2(new_n577), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n473), .A2(new_n472), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n579), .A2(new_n260), .ZN(new_n580));
  INV_X1    g0380(.A(G264), .ZN(new_n581));
  OAI21_X1  g0381(.A(new_n476), .B1(new_n580), .B2(new_n581), .ZN(new_n582));
  OAI211_X1 g0382(.A(G257), .B(G1698), .C1(new_n429), .C2(new_n250), .ZN(new_n583));
  OAI211_X1 g0383(.A(G250), .B(new_n352), .C1(new_n429), .C2(new_n250), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n417), .A2(G294), .ZN(new_n585));
  NAND3_X1  g0385(.A1(new_n583), .A2(new_n584), .A3(new_n585), .ZN(new_n586));
  AOI21_X1  g0386(.A(new_n582), .B1(new_n586), .B2(new_n261), .ZN(new_n587));
  AND2_X1   g0387(.A1(new_n587), .A2(new_n306), .ZN(new_n588));
  NOR2_X1   g0388(.A1(new_n587), .A2(G200), .ZN(new_n589));
  OAI21_X1  g0389(.A(new_n578), .B1(new_n588), .B2(new_n589), .ZN(new_n590));
  AND2_X1   g0390(.A1(new_n587), .A2(G179), .ZN(new_n591));
  NOR2_X1   g0391(.A1(new_n587), .A2(new_n459), .ZN(new_n592));
  OAI22_X1  g0392(.A1(new_n591), .A2(new_n592), .B1(new_n571), .B2(new_n577), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n590), .A2(new_n593), .ZN(new_n594));
  INV_X1    g0394(.A(G270), .ZN(new_n595));
  OAI21_X1  g0395(.A(new_n476), .B1(new_n580), .B2(new_n595), .ZN(new_n596));
  NAND3_X1  g0396(.A1(new_n484), .A2(G257), .A3(new_n352), .ZN(new_n597));
  NAND3_X1  g0397(.A1(new_n484), .A2(G264), .A3(G1698), .ZN(new_n598));
  INV_X1    g0398(.A(G303), .ZN(new_n599));
  OAI211_X1 g0399(.A(new_n597), .B(new_n598), .C1(new_n599), .C2(new_n255), .ZN(new_n600));
  AOI21_X1  g0400(.A(new_n596), .B1(new_n600), .B2(new_n261), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n601), .A2(G190), .ZN(new_n602));
  AOI22_X1  g0402(.A1(new_n281), .A2(new_n219), .B1(G20), .B2(new_n510), .ZN(new_n603));
  AOI21_X1  g0403(.A(G20), .B1(G33), .B2(G283), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n414), .A2(G97), .ZN(new_n605));
  INV_X1    g0405(.A(KEYINPUT80), .ZN(new_n606));
  AND3_X1   g0406(.A1(new_n604), .A2(new_n605), .A3(new_n606), .ZN(new_n607));
  AOI21_X1  g0407(.A(new_n606), .B1(new_n604), .B2(new_n605), .ZN(new_n608));
  OAI21_X1  g0408(.A(new_n603), .B1(new_n607), .B2(new_n608), .ZN(new_n609));
  INV_X1    g0409(.A(KEYINPUT20), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n609), .A2(new_n610), .ZN(new_n611));
  OAI211_X1 g0411(.A(KEYINPUT20), .B(new_n603), .C1(new_n607), .C2(new_n608), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n611), .A2(new_n612), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n545), .A2(G116), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n278), .A2(new_n510), .ZN(new_n615));
  NAND3_X1  g0415(.A1(new_n613), .A2(new_n614), .A3(new_n615), .ZN(new_n616));
  INV_X1    g0416(.A(new_n616), .ZN(new_n617));
  OAI211_X1 g0417(.A(new_n602), .B(new_n617), .C1(new_n439), .C2(new_n601), .ZN(new_n618));
  INV_X1    g0418(.A(KEYINPUT21), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n616), .A2(G169), .ZN(new_n620));
  OAI21_X1  g0420(.A(new_n619), .B1(new_n620), .B2(new_n601), .ZN(new_n621));
  AOI211_X1 g0421(.A(new_n303), .B(new_n596), .C1(new_n600), .C2(new_n261), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n622), .A2(new_n616), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n600), .A2(new_n261), .ZN(new_n624));
  INV_X1    g0424(.A(new_n596), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  NAND4_X1  g0426(.A1(new_n626), .A2(KEYINPUT21), .A3(G169), .A4(new_n616), .ZN(new_n627));
  NAND4_X1  g0427(.A1(new_n618), .A2(new_n621), .A3(new_n623), .A4(new_n627), .ZN(new_n628));
  NOR2_X1   g0428(.A1(new_n594), .A2(new_n628), .ZN(new_n629));
  AND4_X1   g0429(.A1(new_n471), .A2(new_n552), .A3(new_n555), .A4(new_n629), .ZN(G372));
  INV_X1    g0430(.A(new_n550), .ZN(new_n631));
  INV_X1    g0431(.A(KEYINPUT26), .ZN(new_n632));
  OAI21_X1  g0432(.A(new_n632), .B1(new_n554), .B2(new_n506), .ZN(new_n633));
  AND3_X1   g0433(.A1(new_n501), .A2(new_n502), .A3(new_n505), .ZN(new_n634));
  NAND4_X1  g0434(.A1(new_n634), .A2(KEYINPUT26), .A3(new_n550), .A4(new_n539), .ZN(new_n635));
  AOI21_X1  g0435(.A(new_n631), .B1(new_n633), .B2(new_n635), .ZN(new_n636));
  NAND4_X1  g0436(.A1(new_n593), .A2(new_n621), .A3(new_n623), .A4(new_n627), .ZN(new_n637));
  NAND4_X1  g0437(.A1(new_n507), .A2(new_n637), .A3(new_n551), .A4(new_n590), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n636), .A2(new_n638), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n471), .A2(new_n639), .ZN(new_n640));
  XOR2_X1   g0440(.A(new_n640), .B(KEYINPUT83), .Z(new_n641));
  AND2_X1   g0441(.A1(new_n463), .A2(new_n465), .ZN(new_n642));
  AND2_X1   g0442(.A1(new_n441), .A2(new_n458), .ZN(new_n643));
  INV_X1    g0443(.A(new_n643), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n381), .A2(new_n387), .ZN(new_n645));
  AND2_X1   g0445(.A1(new_n366), .A2(new_n645), .ZN(new_n646));
  OAI21_X1  g0446(.A(new_n642), .B1(new_n644), .B2(new_n646), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n312), .A2(new_n314), .ZN(new_n648));
  AOI21_X1  g0448(.A(new_n305), .B1(new_n647), .B2(new_n648), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n641), .A2(new_n649), .ZN(G369));
  NAND3_X1  g0450(.A1(new_n621), .A2(new_n623), .A3(new_n627), .ZN(new_n651));
  NAND3_X1  g0451(.A1(new_n209), .A2(new_n210), .A3(G13), .ZN(new_n652));
  XNOR2_X1  g0452(.A(new_n652), .B(KEYINPUT84), .ZN(new_n653));
  OR2_X1    g0453(.A1(new_n653), .A2(KEYINPUT27), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n653), .A2(KEYINPUT27), .ZN(new_n655));
  NAND3_X1  g0455(.A1(new_n654), .A2(G213), .A3(new_n655), .ZN(new_n656));
  INV_X1    g0456(.A(G343), .ZN(new_n657));
  NOR2_X1   g0457(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  INV_X1    g0458(.A(new_n658), .ZN(new_n659));
  NOR2_X1   g0459(.A1(new_n659), .A2(new_n617), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n651), .A2(new_n660), .ZN(new_n661));
  OAI21_X1  g0461(.A(new_n661), .B1(new_n628), .B2(new_n660), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n662), .A2(KEYINPUT85), .ZN(new_n663));
  INV_X1    g0463(.A(new_n663), .ZN(new_n664));
  NOR2_X1   g0464(.A1(new_n662), .A2(KEYINPUT85), .ZN(new_n665));
  OAI21_X1  g0465(.A(G330), .B1(new_n664), .B2(new_n665), .ZN(new_n666));
  INV_X1    g0466(.A(new_n666), .ZN(new_n667));
  INV_X1    g0467(.A(new_n593), .ZN(new_n668));
  NAND3_X1  g0468(.A1(new_n668), .A2(KEYINPUT86), .A3(new_n658), .ZN(new_n669));
  INV_X1    g0469(.A(KEYINPUT86), .ZN(new_n670));
  OAI21_X1  g0470(.A(new_n670), .B1(new_n593), .B2(new_n659), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n669), .A2(new_n671), .ZN(new_n672));
  OAI211_X1 g0472(.A(new_n590), .B(new_n593), .C1(new_n578), .C2(new_n659), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n667), .A2(new_n674), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n651), .A2(new_n659), .ZN(new_n676));
  AOI21_X1  g0476(.A(new_n676), .B1(new_n672), .B2(new_n673), .ZN(new_n677));
  XNOR2_X1  g0477(.A(new_n658), .B(KEYINPUT87), .ZN(new_n678));
  INV_X1    g0478(.A(new_n678), .ZN(new_n679));
  NOR2_X1   g0479(.A1(new_n679), .A2(new_n593), .ZN(new_n680));
  NOR2_X1   g0480(.A1(new_n677), .A2(new_n680), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n675), .A2(new_n681), .ZN(G399));
  INV_X1    g0482(.A(new_n213), .ZN(new_n683));
  NOR2_X1   g0483(.A1(new_n683), .A2(G41), .ZN(new_n684));
  INV_X1    g0484(.A(new_n684), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n526), .A2(new_n510), .ZN(new_n686));
  INV_X1    g0486(.A(new_n686), .ZN(new_n687));
  NAND3_X1  g0487(.A1(new_n685), .A2(G1), .A3(new_n687), .ZN(new_n688));
  OAI22_X1  g0488(.A1(new_n688), .A2(KEYINPUT88), .B1(new_n217), .B2(new_n685), .ZN(new_n689));
  AOI21_X1  g0489(.A(new_n689), .B1(KEYINPUT88), .B2(new_n688), .ZN(new_n690));
  XOR2_X1   g0490(.A(new_n690), .B(KEYINPUT28), .Z(new_n691));
  INV_X1    g0491(.A(KEYINPUT31), .ZN(new_n692));
  AND4_X1   g0492(.A1(new_n504), .A2(new_n515), .A3(new_n475), .A4(new_n524), .ZN(new_n693));
  INV_X1    g0493(.A(KEYINPUT30), .ZN(new_n694));
  NAND4_X1  g0494(.A1(new_n693), .A2(new_n694), .A3(new_n587), .A4(new_n622), .ZN(new_n695));
  NAND4_X1  g0495(.A1(new_n538), .A2(new_n587), .A3(new_n504), .A4(new_n475), .ZN(new_n696));
  NAND3_X1  g0496(.A1(new_n624), .A2(G179), .A3(new_n625), .ZN(new_n697));
  OAI21_X1  g0497(.A(KEYINPUT30), .B1(new_n696), .B2(new_n697), .ZN(new_n698));
  OAI21_X1  g0498(.A(new_n303), .B1(new_n542), .B2(new_n523), .ZN(new_n699));
  NOR3_X1   g0499(.A1(new_n699), .A2(new_n587), .A3(new_n601), .ZN(new_n700));
  AOI22_X1  g0500(.A1(new_n695), .A2(new_n698), .B1(new_n700), .B2(new_n487), .ZN(new_n701));
  INV_X1    g0501(.A(KEYINPUT89), .ZN(new_n702));
  OAI21_X1  g0502(.A(new_n658), .B1(new_n701), .B2(new_n702), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n695), .A2(new_n698), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n700), .A2(new_n487), .ZN(new_n705));
  AND3_X1   g0505(.A1(new_n704), .A2(new_n702), .A3(new_n705), .ZN(new_n706));
  OAI21_X1  g0506(.A(new_n692), .B1(new_n703), .B2(new_n706), .ZN(new_n707));
  NAND4_X1  g0507(.A1(new_n629), .A2(new_n552), .A3(new_n555), .A4(new_n678), .ZN(new_n708));
  INV_X1    g0508(.A(new_n475), .ZN(new_n709));
  AND3_X1   g0509(.A1(new_n480), .A2(new_n481), .A3(new_n482), .ZN(new_n710));
  AOI211_X1 g0510(.A(new_n478), .B(G1698), .C1(new_n420), .C2(new_n406), .ZN(new_n711));
  OAI21_X1  g0511(.A(new_n710), .B1(new_n711), .B2(KEYINPUT4), .ZN(new_n712));
  AOI21_X1  g0512(.A(new_n709), .B1(new_n712), .B2(new_n261), .ZN(new_n713));
  AND3_X1   g0513(.A1(new_n713), .A2(new_n538), .A3(new_n587), .ZN(new_n714));
  AOI21_X1  g0514(.A(new_n694), .B1(new_n714), .B2(new_n622), .ZN(new_n715));
  NOR3_X1   g0515(.A1(new_n696), .A2(new_n697), .A3(KEYINPUT30), .ZN(new_n716));
  OAI21_X1  g0516(.A(new_n705), .B1(new_n715), .B2(new_n716), .ZN(new_n717));
  NAND3_X1  g0517(.A1(new_n717), .A2(KEYINPUT31), .A3(new_n679), .ZN(new_n718));
  NAND3_X1  g0518(.A1(new_n707), .A2(new_n708), .A3(new_n718), .ZN(new_n719));
  AND3_X1   g0519(.A1(new_n719), .A2(KEYINPUT90), .A3(G330), .ZN(new_n720));
  AOI21_X1  g0520(.A(KEYINPUT90), .B1(new_n719), .B2(G330), .ZN(new_n721));
  NOR2_X1   g0521(.A1(new_n720), .A2(new_n721), .ZN(new_n722));
  INV_X1    g0522(.A(KEYINPUT93), .ZN(new_n723));
  NAND2_X1  g0523(.A1(new_n637), .A2(new_n723), .ZN(new_n724));
  AND2_X1   g0524(.A1(new_n627), .A2(new_n623), .ZN(new_n725));
  NAND4_X1  g0525(.A1(new_n725), .A2(KEYINPUT93), .A3(new_n593), .A4(new_n621), .ZN(new_n726));
  NOR2_X1   g0526(.A1(new_n553), .A2(new_n554), .ZN(new_n727));
  NAND4_X1  g0527(.A1(new_n724), .A2(new_n726), .A3(new_n727), .A4(new_n590), .ZN(new_n728));
  AOI21_X1  g0528(.A(KEYINPUT26), .B1(new_n551), .B2(new_n634), .ZN(new_n729));
  INV_X1    g0529(.A(KEYINPUT92), .ZN(new_n730));
  NOR2_X1   g0530(.A1(new_n730), .A2(KEYINPUT26), .ZN(new_n731));
  AOI21_X1  g0531(.A(new_n631), .B1(new_n729), .B2(new_n731), .ZN(new_n732));
  NAND3_X1  g0532(.A1(new_n633), .A2(new_n635), .A3(new_n730), .ZN(new_n733));
  NAND3_X1  g0533(.A1(new_n728), .A2(new_n732), .A3(new_n733), .ZN(new_n734));
  NAND3_X1  g0534(.A1(new_n734), .A2(KEYINPUT29), .A3(new_n659), .ZN(new_n735));
  AOI21_X1  g0535(.A(new_n679), .B1(new_n636), .B2(new_n638), .ZN(new_n736));
  XNOR2_X1  g0536(.A(KEYINPUT91), .B(KEYINPUT29), .ZN(new_n737));
  OAI21_X1  g0537(.A(new_n735), .B1(new_n736), .B2(new_n737), .ZN(new_n738));
  NAND2_X1  g0538(.A1(new_n722), .A2(new_n738), .ZN(new_n739));
  INV_X1    g0539(.A(new_n739), .ZN(new_n740));
  OAI21_X1  g0540(.A(new_n691), .B1(new_n740), .B2(G1), .ZN(G364));
  NOR2_X1   g0541(.A1(new_n277), .A2(G20), .ZN(new_n742));
  AOI21_X1  g0542(.A(new_n209), .B1(new_n742), .B2(G45), .ZN(new_n743));
  INV_X1    g0543(.A(new_n743), .ZN(new_n744));
  NOR2_X1   g0544(.A1(new_n684), .A2(new_n744), .ZN(new_n745));
  INV_X1    g0545(.A(new_n745), .ZN(new_n746));
  OR3_X1    g0546(.A1(new_n664), .A2(G330), .A3(new_n665), .ZN(new_n747));
  NAND3_X1  g0547(.A1(new_n666), .A2(new_n746), .A3(new_n747), .ZN(new_n748));
  NOR2_X1   g0548(.A1(new_n683), .A2(new_n251), .ZN(new_n749));
  NAND2_X1  g0549(.A1(new_n749), .A2(G355), .ZN(new_n750));
  OAI21_X1  g0550(.A(new_n750), .B1(G116), .B2(new_n213), .ZN(new_n751));
  NOR2_X1   g0551(.A1(new_n683), .A2(new_n484), .ZN(new_n752));
  INV_X1    g0552(.A(new_n752), .ZN(new_n753));
  AOI21_X1  g0553(.A(new_n753), .B1(new_n264), .B2(new_n218), .ZN(new_n754));
  NAND2_X1  g0554(.A1(new_n247), .A2(G45), .ZN(new_n755));
  AOI21_X1  g0555(.A(new_n751), .B1(new_n754), .B2(new_n755), .ZN(new_n756));
  NOR2_X1   g0556(.A1(G13), .A2(G33), .ZN(new_n757));
  INV_X1    g0557(.A(new_n757), .ZN(new_n758));
  NOR2_X1   g0558(.A1(new_n758), .A2(G20), .ZN(new_n759));
  AOI21_X1  g0559(.A(new_n219), .B1(G20), .B2(new_n459), .ZN(new_n760));
  NOR2_X1   g0560(.A1(new_n759), .A2(new_n760), .ZN(new_n761));
  INV_X1    g0561(.A(new_n761), .ZN(new_n762));
  OAI21_X1  g0562(.A(new_n745), .B1(new_n756), .B2(new_n762), .ZN(new_n763));
  NOR2_X1   g0563(.A1(new_n210), .A2(G179), .ZN(new_n764));
  NOR2_X1   g0564(.A1(G190), .A2(G200), .ZN(new_n765));
  NAND2_X1  g0565(.A1(new_n764), .A2(new_n765), .ZN(new_n766));
  INV_X1    g0566(.A(G159), .ZN(new_n767));
  NOR3_X1   g0567(.A1(new_n766), .A2(KEYINPUT32), .A3(new_n767), .ZN(new_n768));
  NAND3_X1  g0568(.A1(new_n764), .A2(G190), .A3(G200), .ZN(new_n769));
  INV_X1    g0569(.A(new_n769), .ZN(new_n770));
  AOI21_X1  g0570(.A(new_n768), .B1(G87), .B2(new_n770), .ZN(new_n771));
  NAND3_X1  g0571(.A1(new_n764), .A2(new_n306), .A3(G200), .ZN(new_n772));
  INV_X1    g0572(.A(new_n772), .ZN(new_n773));
  NAND2_X1  g0573(.A1(new_n773), .A2(G107), .ZN(new_n774));
  OAI21_X1  g0574(.A(KEYINPUT32), .B1(new_n766), .B2(new_n767), .ZN(new_n775));
  NAND3_X1  g0575(.A1(new_n771), .A2(new_n774), .A3(new_n775), .ZN(new_n776));
  NOR2_X1   g0576(.A1(new_n210), .A2(new_n303), .ZN(new_n777));
  INV_X1    g0577(.A(new_n777), .ZN(new_n778));
  OR3_X1    g0578(.A1(new_n778), .A2(KEYINPUT95), .A3(new_n439), .ZN(new_n779));
  OAI21_X1  g0579(.A(KEYINPUT95), .B1(new_n778), .B2(new_n439), .ZN(new_n780));
  NAND3_X1  g0580(.A1(new_n779), .A2(G190), .A3(new_n780), .ZN(new_n781));
  NAND3_X1  g0581(.A1(new_n779), .A2(new_n306), .A3(new_n780), .ZN(new_n782));
  OAI22_X1  g0582(.A1(new_n202), .A2(new_n781), .B1(new_n782), .B2(new_n318), .ZN(new_n783));
  AND3_X1   g0583(.A1(new_n777), .A2(KEYINPUT94), .A3(new_n765), .ZN(new_n784));
  AOI21_X1  g0584(.A(KEYINPUT94), .B1(new_n777), .B2(new_n765), .ZN(new_n785));
  OR2_X1    g0585(.A1(new_n784), .A2(new_n785), .ZN(new_n786));
  INV_X1    g0586(.A(new_n786), .ZN(new_n787));
  NOR2_X1   g0587(.A1(new_n787), .A2(new_n254), .ZN(new_n788));
  NOR3_X1   g0588(.A1(new_n306), .A2(G179), .A3(G200), .ZN(new_n789));
  NOR2_X1   g0589(.A1(new_n789), .A2(new_n210), .ZN(new_n790));
  NOR3_X1   g0590(.A1(new_n778), .A2(new_n306), .A3(G200), .ZN(new_n791));
  INV_X1    g0591(.A(new_n791), .ZN(new_n792));
  OAI221_X1 g0592(.A(new_n255), .B1(new_n205), .B2(new_n790), .C1(new_n792), .C2(new_n396), .ZN(new_n793));
  OR4_X1    g0593(.A1(new_n776), .A2(new_n783), .A3(new_n788), .A4(new_n793), .ZN(new_n794));
  INV_X1    g0594(.A(new_n781), .ZN(new_n795));
  NAND2_X1  g0595(.A1(new_n795), .A2(G326), .ZN(new_n796));
  INV_X1    g0596(.A(new_n782), .ZN(new_n797));
  XNOR2_X1  g0597(.A(KEYINPUT33), .B(G317), .ZN(new_n798));
  NAND2_X1  g0598(.A1(new_n797), .A2(new_n798), .ZN(new_n799));
  NAND2_X1  g0599(.A1(new_n777), .A2(new_n765), .ZN(new_n800));
  INV_X1    g0600(.A(G311), .ZN(new_n801));
  INV_X1    g0601(.A(G329), .ZN(new_n802));
  OAI22_X1  g0602(.A1(new_n800), .A2(new_n801), .B1(new_n766), .B2(new_n802), .ZN(new_n803));
  AOI211_X1 g0603(.A(new_n255), .B(new_n803), .C1(G322), .C2(new_n791), .ZN(new_n804));
  INV_X1    g0604(.A(G283), .ZN(new_n805));
  OAI22_X1  g0605(.A1(new_n805), .A2(new_n772), .B1(new_n769), .B2(new_n599), .ZN(new_n806));
  INV_X1    g0606(.A(new_n790), .ZN(new_n807));
  AOI21_X1  g0607(.A(new_n806), .B1(G294), .B2(new_n807), .ZN(new_n808));
  NAND4_X1  g0608(.A1(new_n796), .A2(new_n799), .A3(new_n804), .A4(new_n808), .ZN(new_n809));
  NAND2_X1  g0609(.A1(new_n794), .A2(new_n809), .ZN(new_n810));
  AOI21_X1  g0610(.A(new_n763), .B1(new_n810), .B2(new_n760), .ZN(new_n811));
  INV_X1    g0611(.A(new_n759), .ZN(new_n812));
  OAI21_X1  g0612(.A(new_n811), .B1(new_n662), .B2(new_n812), .ZN(new_n813));
  AND2_X1   g0613(.A1(new_n748), .A2(new_n813), .ZN(new_n814));
  INV_X1    g0614(.A(new_n814), .ZN(G396));
  INV_X1    g0615(.A(KEYINPUT98), .ZN(new_n816));
  NAND2_X1  g0616(.A1(new_n639), .A2(new_n678), .ZN(new_n817));
  NOR4_X1   g0617(.A1(new_n372), .A2(new_n380), .A3(new_n379), .A4(new_n658), .ZN(new_n818));
  OAI21_X1  g0618(.A(new_n384), .B1(new_n379), .B2(new_n659), .ZN(new_n819));
  AOI21_X1  g0619(.A(new_n818), .B1(new_n819), .B2(new_n382), .ZN(new_n820));
  INV_X1    g0620(.A(new_n820), .ZN(new_n821));
  OAI21_X1  g0621(.A(new_n816), .B1(new_n817), .B2(new_n821), .ZN(new_n822));
  NAND3_X1  g0622(.A1(new_n736), .A2(KEYINPUT98), .A3(new_n820), .ZN(new_n823));
  AOI22_X1  g0623(.A1(new_n822), .A2(new_n823), .B1(new_n817), .B2(new_n821), .ZN(new_n824));
  OAI21_X1  g0624(.A(new_n824), .B1(new_n721), .B2(new_n720), .ZN(new_n825));
  NAND2_X1  g0625(.A1(new_n825), .A2(new_n746), .ZN(new_n826));
  INV_X1    g0626(.A(new_n824), .ZN(new_n827));
  AOI22_X1  g0627(.A1(new_n826), .A2(KEYINPUT99), .B1(new_n722), .B2(new_n827), .ZN(new_n828));
  OAI21_X1  g0628(.A(new_n828), .B1(KEYINPUT99), .B2(new_n826), .ZN(new_n829));
  NOR2_X1   g0629(.A1(new_n760), .A2(new_n757), .ZN(new_n830));
  XNOR2_X1  g0630(.A(new_n830), .B(KEYINPUT96), .ZN(new_n831));
  OAI21_X1  g0631(.A(new_n745), .B1(new_n831), .B2(G77), .ZN(new_n832));
  XOR2_X1   g0632(.A(new_n832), .B(KEYINPUT97), .Z(new_n833));
  INV_X1    g0633(.A(new_n760), .ZN(new_n834));
  OAI22_X1  g0634(.A1(new_n805), .A2(new_n782), .B1(new_n781), .B2(new_n599), .ZN(new_n835));
  NOR2_X1   g0635(.A1(new_n787), .A2(new_n510), .ZN(new_n836));
  INV_X1    g0636(.A(G294), .ZN(new_n837));
  OAI221_X1 g0637(.A(new_n251), .B1(new_n766), .B2(new_n801), .C1(new_n792), .C2(new_n837), .ZN(new_n838));
  NAND2_X1  g0638(.A1(new_n773), .A2(G87), .ZN(new_n839));
  OAI221_X1 g0639(.A(new_n839), .B1(new_n206), .B2(new_n769), .C1(new_n205), .C2(new_n790), .ZN(new_n840));
  NOR4_X1   g0640(.A1(new_n835), .A2(new_n836), .A3(new_n838), .A4(new_n840), .ZN(new_n841));
  AOI22_X1  g0641(.A1(new_n786), .A2(G159), .B1(G143), .B2(new_n791), .ZN(new_n842));
  INV_X1    g0642(.A(G137), .ZN(new_n843));
  INV_X1    g0643(.A(G150), .ZN(new_n844));
  OAI221_X1 g0644(.A(new_n842), .B1(new_n843), .B2(new_n781), .C1(new_n844), .C2(new_n782), .ZN(new_n845));
  XNOR2_X1  g0645(.A(new_n845), .B(KEYINPUT34), .ZN(new_n846));
  OAI22_X1  g0646(.A1(new_n790), .A2(new_n396), .B1(new_n772), .B2(new_n318), .ZN(new_n847));
  INV_X1    g0647(.A(G132), .ZN(new_n848));
  OAI21_X1  g0648(.A(new_n484), .B1(new_n848), .B2(new_n766), .ZN(new_n849));
  AOI211_X1 g0649(.A(new_n847), .B(new_n849), .C1(G50), .C2(new_n770), .ZN(new_n850));
  AOI21_X1  g0650(.A(new_n841), .B1(new_n846), .B2(new_n850), .ZN(new_n851));
  OAI221_X1 g0651(.A(new_n833), .B1(new_n834), .B2(new_n851), .C1(new_n820), .C2(new_n758), .ZN(new_n852));
  NAND2_X1  g0652(.A1(new_n829), .A2(new_n852), .ZN(G384));
  NOR3_X1   g0653(.A1(new_n219), .A2(new_n210), .A3(new_n510), .ZN(new_n854));
  NOR2_X1   g0654(.A1(new_n495), .A2(new_n496), .ZN(new_n855));
  XNOR2_X1  g0655(.A(new_n855), .B(KEYINPUT100), .ZN(new_n856));
  INV_X1    g0656(.A(new_n856), .ZN(new_n857));
  INV_X1    g0657(.A(KEYINPUT35), .ZN(new_n858));
  OAI21_X1  g0658(.A(new_n854), .B1(new_n857), .B2(new_n858), .ZN(new_n859));
  AOI21_X1  g0659(.A(new_n859), .B1(new_n858), .B2(new_n857), .ZN(new_n860));
  XNOR2_X1  g0660(.A(new_n860), .B(KEYINPUT36), .ZN(new_n861));
  OAI211_X1 g0661(.A(new_n218), .B(G77), .C1(new_n222), .C2(new_n396), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n202), .A2(G68), .ZN(new_n863));
  AOI211_X1 g0663(.A(new_n209), .B(G13), .C1(new_n862), .C2(new_n863), .ZN(new_n864));
  NOR2_X1   g0664(.A1(new_n861), .A2(new_n864), .ZN(new_n865));
  INV_X1    g0665(.A(G330), .ZN(new_n866));
  NAND3_X1  g0666(.A1(new_n457), .A2(new_n424), .A3(new_n437), .ZN(new_n867));
  INV_X1    g0667(.A(KEYINPUT37), .ZN(new_n868));
  INV_X1    g0668(.A(new_n656), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n449), .A2(new_n869), .ZN(new_n870));
  NAND4_X1  g0670(.A1(new_n867), .A2(new_n462), .A3(new_n868), .A4(new_n870), .ZN(new_n871));
  INV_X1    g0671(.A(KEYINPUT103), .ZN(new_n872));
  NAND3_X1  g0672(.A1(new_n420), .A2(new_n210), .A3(new_n406), .ZN(new_n873));
  NAND2_X1  g0673(.A1(new_n873), .A2(KEYINPUT7), .ZN(new_n874));
  NAND3_X1  g0674(.A1(new_n874), .A2(G68), .A3(new_n421), .ZN(new_n875));
  AOI21_X1  g0675(.A(KEYINPUT16), .B1(new_n875), .B2(new_n398), .ZN(new_n876));
  OAI21_X1  g0676(.A(new_n872), .B1(new_n876), .B2(new_n286), .ZN(new_n877));
  AND2_X1   g0677(.A1(new_n421), .A2(G68), .ZN(new_n878));
  AOI21_X1  g0678(.A(new_n446), .B1(new_n878), .B2(new_n874), .ZN(new_n879));
  OAI211_X1 g0679(.A(KEYINPUT103), .B(new_n282), .C1(new_n879), .C2(KEYINPUT16), .ZN(new_n880));
  NAND3_X1  g0680(.A1(new_n877), .A2(new_n880), .A3(new_n423), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n456), .A2(G169), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n436), .A2(G179), .ZN(new_n883));
  AOI22_X1  g0683(.A1(new_n881), .A2(new_n392), .B1(new_n882), .B2(new_n883), .ZN(new_n884));
  AOI21_X1  g0684(.A(new_n656), .B1(new_n881), .B2(new_n392), .ZN(new_n885));
  NOR3_X1   g0685(.A1(new_n440), .A2(new_n449), .A3(new_n450), .ZN(new_n886));
  NOR3_X1   g0686(.A1(new_n884), .A2(new_n885), .A3(new_n886), .ZN(new_n887));
  OAI21_X1  g0687(.A(new_n871), .B1(new_n887), .B2(new_n868), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n466), .A2(new_n885), .ZN(new_n889));
  NAND3_X1  g0689(.A1(new_n888), .A2(KEYINPUT38), .A3(new_n889), .ZN(new_n890));
  INV_X1    g0690(.A(KEYINPUT104), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n890), .A2(new_n891), .ZN(new_n892));
  NAND4_X1  g0692(.A1(new_n888), .A2(KEYINPUT104), .A3(KEYINPUT38), .A4(new_n889), .ZN(new_n893));
  INV_X1    g0693(.A(KEYINPUT38), .ZN(new_n894));
  OAI21_X1  g0694(.A(new_n398), .B1(new_n419), .B2(new_n422), .ZN(new_n895));
  AOI21_X1  g0695(.A(new_n286), .B1(new_n895), .B2(new_n410), .ZN(new_n896));
  OAI21_X1  g0696(.A(new_n423), .B1(new_n896), .B2(KEYINPUT103), .ZN(new_n897));
  NOR3_X1   g0697(.A1(new_n876), .A2(new_n872), .A3(new_n286), .ZN(new_n898));
  OAI21_X1  g0698(.A(new_n392), .B1(new_n897), .B2(new_n898), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n899), .A2(new_n869), .ZN(new_n900));
  AOI21_X1  g0700(.A(new_n900), .B1(new_n643), .B2(new_n642), .ZN(new_n901));
  AND4_X1   g0701(.A1(new_n868), .A2(new_n867), .A3(new_n462), .A4(new_n870), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n882), .A2(new_n883), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n899), .A2(new_n903), .ZN(new_n904));
  NAND3_X1  g0704(.A1(new_n904), .A2(new_n900), .A3(new_n867), .ZN(new_n905));
  AOI21_X1  g0705(.A(new_n902), .B1(new_n905), .B2(KEYINPUT37), .ZN(new_n906));
  OAI21_X1  g0706(.A(new_n894), .B1(new_n901), .B2(new_n906), .ZN(new_n907));
  NAND3_X1  g0707(.A1(new_n892), .A2(new_n893), .A3(new_n907), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n717), .A2(KEYINPUT89), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n701), .A2(new_n702), .ZN(new_n910));
  NAND4_X1  g0710(.A1(new_n909), .A2(KEYINPUT31), .A3(new_n910), .A4(new_n658), .ZN(new_n911));
  NAND3_X1  g0711(.A1(new_n707), .A2(new_n708), .A3(new_n911), .ZN(new_n912));
  INV_X1    g0712(.A(KEYINPUT101), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n366), .A2(new_n913), .ZN(new_n914));
  OAI211_X1 g0714(.A(KEYINPUT101), .B(new_n338), .C1(new_n363), .C2(new_n365), .ZN(new_n915));
  NOR2_X1   g0715(.A1(new_n337), .A2(new_n659), .ZN(new_n916));
  INV_X1    g0716(.A(new_n916), .ZN(new_n917));
  AND2_X1   g0717(.A1(new_n917), .A2(new_n387), .ZN(new_n918));
  NAND3_X1  g0718(.A1(new_n914), .A2(new_n915), .A3(new_n918), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n364), .A2(G169), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n920), .A2(KEYINPUT14), .ZN(new_n921));
  NAND4_X1  g0721(.A1(new_n387), .A2(new_n921), .A3(new_n362), .A4(new_n359), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n922), .A2(new_n916), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n923), .A2(KEYINPUT102), .ZN(new_n924));
  INV_X1    g0724(.A(KEYINPUT102), .ZN(new_n925));
  NAND3_X1  g0725(.A1(new_n922), .A2(new_n925), .A3(new_n916), .ZN(new_n926));
  NAND3_X1  g0726(.A1(new_n919), .A2(new_n924), .A3(new_n926), .ZN(new_n927));
  AND3_X1   g0727(.A1(new_n912), .A2(new_n820), .A3(new_n927), .ZN(new_n928));
  AOI21_X1  g0728(.A(KEYINPUT40), .B1(new_n908), .B2(new_n928), .ZN(new_n929));
  INV_X1    g0729(.A(KEYINPUT40), .ZN(new_n930));
  INV_X1    g0730(.A(new_n870), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n466), .A2(new_n931), .ZN(new_n932));
  NAND3_X1  g0732(.A1(new_n867), .A2(new_n462), .A3(new_n870), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n933), .A2(KEYINPUT37), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n934), .A2(new_n871), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n932), .A2(new_n935), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n936), .A2(new_n894), .ZN(new_n937));
  AOI21_X1  g0737(.A(new_n930), .B1(new_n937), .B2(new_n890), .ZN(new_n938));
  AOI21_X1  g0738(.A(new_n929), .B1(new_n928), .B2(new_n938), .ZN(new_n939));
  AND2_X1   g0739(.A1(new_n471), .A2(new_n912), .ZN(new_n940));
  AOI21_X1  g0740(.A(new_n866), .B1(new_n939), .B2(new_n940), .ZN(new_n941));
  OAI21_X1  g0741(.A(new_n941), .B1(new_n939), .B2(new_n940), .ZN(new_n942));
  INV_X1    g0742(.A(new_n818), .ZN(new_n943));
  AND4_X1   g0743(.A1(KEYINPUT98), .A2(new_n639), .A3(new_n820), .A4(new_n678), .ZN(new_n944));
  AOI21_X1  g0744(.A(KEYINPUT98), .B1(new_n736), .B2(new_n820), .ZN(new_n945));
  OAI21_X1  g0745(.A(new_n943), .B1(new_n944), .B2(new_n945), .ZN(new_n946));
  NAND3_X1  g0746(.A1(new_n908), .A2(new_n946), .A3(new_n927), .ZN(new_n947));
  OR2_X1    g0747(.A1(new_n642), .A2(new_n869), .ZN(new_n948));
  INV_X1    g0748(.A(KEYINPUT39), .ZN(new_n949));
  AND3_X1   g0749(.A1(new_n937), .A2(new_n949), .A3(new_n890), .ZN(new_n950));
  AOI21_X1  g0750(.A(new_n950), .B1(new_n908), .B2(KEYINPUT39), .ZN(new_n951));
  AOI21_X1  g0751(.A(new_n658), .B1(new_n914), .B2(new_n915), .ZN(new_n952));
  INV_X1    g0752(.A(new_n952), .ZN(new_n953));
  OAI211_X1 g0753(.A(new_n947), .B(new_n948), .C1(new_n951), .C2(new_n953), .ZN(new_n954));
  OR2_X1    g0754(.A1(new_n470), .A2(new_n738), .ZN(new_n955));
  NAND2_X1  g0755(.A1(new_n955), .A2(new_n649), .ZN(new_n956));
  XNOR2_X1  g0756(.A(new_n954), .B(new_n956), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n942), .A2(new_n957), .ZN(new_n958));
  OAI21_X1  g0758(.A(new_n958), .B1(new_n209), .B2(new_n742), .ZN(new_n959));
  NOR2_X1   g0759(.A1(new_n942), .A2(new_n957), .ZN(new_n960));
  OAI21_X1  g0760(.A(new_n865), .B1(new_n959), .B2(new_n960), .ZN(new_n961));
  XNOR2_X1  g0761(.A(new_n961), .B(KEYINPUT105), .ZN(G367));
  NOR2_X1   g0762(.A1(new_n659), .A2(new_n537), .ZN(new_n963));
  NAND2_X1  g0763(.A1(new_n963), .A2(new_n550), .ZN(new_n964));
  OAI21_X1  g0764(.A(new_n964), .B1(new_n551), .B2(new_n963), .ZN(new_n965));
  XOR2_X1   g0765(.A(new_n965), .B(KEYINPUT106), .Z(new_n966));
  NAND2_X1  g0766(.A1(new_n966), .A2(new_n759), .ZN(new_n967));
  OAI221_X1 g0767(.A(new_n761), .B1(new_n213), .B2(new_n377), .C1(new_n753), .C2(new_n239), .ZN(new_n968));
  NAND2_X1  g0768(.A1(new_n968), .A2(new_n745), .ZN(new_n969));
  AOI22_X1  g0769(.A1(G143), .A2(new_n795), .B1(new_n797), .B2(G159), .ZN(new_n970));
  NOR2_X1   g0770(.A1(new_n772), .A2(new_n254), .ZN(new_n971));
  NOR2_X1   g0771(.A1(new_n790), .A2(new_n318), .ZN(new_n972));
  AOI211_X1 g0772(.A(new_n971), .B(new_n972), .C1(new_n292), .C2(new_n770), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n786), .A2(G50), .ZN(new_n974));
  OAI21_X1  g0774(.A(new_n255), .B1(new_n766), .B2(new_n843), .ZN(new_n975));
  AOI21_X1  g0775(.A(new_n975), .B1(new_n791), .B2(G150), .ZN(new_n976));
  NAND4_X1  g0776(.A1(new_n970), .A2(new_n973), .A3(new_n974), .A4(new_n976), .ZN(new_n977));
  INV_X1    g0777(.A(G317), .ZN(new_n978));
  OAI21_X1  g0778(.A(new_n418), .B1(new_n978), .B2(new_n766), .ZN(new_n979));
  OAI22_X1  g0779(.A1(new_n790), .A2(new_n206), .B1(new_n772), .B2(new_n205), .ZN(new_n980));
  AOI211_X1 g0780(.A(new_n979), .B(new_n980), .C1(new_n797), .C2(G294), .ZN(new_n981));
  OAI22_X1  g0781(.A1(new_n781), .A2(new_n801), .B1(new_n599), .B2(new_n792), .ZN(new_n982));
  INV_X1    g0782(.A(KEYINPUT109), .ZN(new_n983));
  NAND2_X1  g0783(.A1(new_n982), .A2(new_n983), .ZN(new_n984));
  NOR2_X1   g0784(.A1(new_n769), .A2(new_n510), .ZN(new_n985));
  XNOR2_X1  g0785(.A(new_n985), .B(KEYINPUT46), .ZN(new_n986));
  AOI21_X1  g0786(.A(new_n986), .B1(G283), .B2(new_n786), .ZN(new_n987));
  NAND3_X1  g0787(.A1(new_n981), .A2(new_n984), .A3(new_n987), .ZN(new_n988));
  NOR2_X1   g0788(.A1(new_n982), .A2(new_n983), .ZN(new_n989));
  OAI21_X1  g0789(.A(new_n977), .B1(new_n988), .B2(new_n989), .ZN(new_n990));
  XOR2_X1   g0790(.A(KEYINPUT110), .B(KEYINPUT47), .Z(new_n991));
  XNOR2_X1  g0791(.A(new_n990), .B(new_n991), .ZN(new_n992));
  AOI21_X1  g0792(.A(new_n969), .B1(new_n992), .B2(new_n760), .ZN(new_n993));
  NAND2_X1  g0793(.A1(new_n967), .A2(new_n993), .ZN(new_n994));
  INV_X1    g0794(.A(KEYINPUT107), .ZN(new_n995));
  INV_X1    g0795(.A(new_n676), .ZN(new_n996));
  NAND2_X1  g0796(.A1(new_n674), .A2(new_n996), .ZN(new_n997));
  OAI21_X1  g0797(.A(new_n507), .B1(new_n499), .B2(new_n678), .ZN(new_n998));
  NAND2_X1  g0798(.A1(new_n679), .A2(new_n634), .ZN(new_n999));
  NAND2_X1  g0799(.A1(new_n998), .A2(new_n999), .ZN(new_n1000));
  INV_X1    g0800(.A(new_n1000), .ZN(new_n1001));
  OAI21_X1  g0801(.A(new_n995), .B1(new_n997), .B2(new_n1001), .ZN(new_n1002));
  NAND3_X1  g0802(.A1(new_n677), .A2(KEYINPUT107), .A3(new_n1000), .ZN(new_n1003));
  NAND2_X1  g0803(.A1(new_n1002), .A2(new_n1003), .ZN(new_n1004));
  OR2_X1    g0804(.A1(new_n1004), .A2(KEYINPUT42), .ZN(new_n1005));
  OAI21_X1  g0805(.A(new_n506), .B1(new_n998), .B2(new_n593), .ZN(new_n1006));
  NAND2_X1  g0806(.A1(new_n1006), .A2(new_n678), .ZN(new_n1007));
  NAND2_X1  g0807(.A1(new_n1004), .A2(KEYINPUT42), .ZN(new_n1008));
  NAND3_X1  g0808(.A1(new_n1005), .A2(new_n1007), .A3(new_n1008), .ZN(new_n1009));
  INV_X1    g0809(.A(KEYINPUT43), .ZN(new_n1010));
  NAND2_X1  g0810(.A1(new_n966), .A2(new_n1010), .ZN(new_n1011));
  OR2_X1    g0811(.A1(new_n966), .A2(new_n1010), .ZN(new_n1012));
  NAND3_X1  g0812(.A1(new_n1009), .A2(new_n1011), .A3(new_n1012), .ZN(new_n1013));
  AND2_X1   g0813(.A1(new_n1008), .A2(new_n1007), .ZN(new_n1014));
  NAND4_X1  g0814(.A1(new_n1014), .A2(new_n1010), .A3(new_n966), .A4(new_n1005), .ZN(new_n1015));
  NAND2_X1  g0815(.A1(new_n1013), .A2(new_n1015), .ZN(new_n1016));
  OAI21_X1  g0816(.A(new_n1016), .B1(new_n675), .B2(new_n1001), .ZN(new_n1017));
  INV_X1    g0817(.A(new_n675), .ZN(new_n1018));
  NAND4_X1  g0818(.A1(new_n1013), .A2(new_n1015), .A3(new_n1018), .A4(new_n1000), .ZN(new_n1019));
  NAND2_X1  g0819(.A1(new_n1017), .A2(new_n1019), .ZN(new_n1020));
  INV_X1    g0820(.A(KEYINPUT45), .ZN(new_n1021));
  INV_X1    g0821(.A(new_n680), .ZN(new_n1022));
  NAND2_X1  g0822(.A1(new_n997), .A2(new_n1022), .ZN(new_n1023));
  OAI21_X1  g0823(.A(new_n1021), .B1(new_n1023), .B2(new_n1001), .ZN(new_n1024));
  NAND3_X1  g0824(.A1(new_n681), .A2(KEYINPUT45), .A3(new_n1000), .ZN(new_n1025));
  NAND2_X1  g0825(.A1(new_n1024), .A2(new_n1025), .ZN(new_n1026));
  NAND3_X1  g0826(.A1(new_n1023), .A2(KEYINPUT44), .A3(new_n1001), .ZN(new_n1027));
  INV_X1    g0827(.A(KEYINPUT44), .ZN(new_n1028));
  OAI21_X1  g0828(.A(new_n1028), .B1(new_n681), .B2(new_n1000), .ZN(new_n1029));
  NAND2_X1  g0829(.A1(new_n1027), .A2(new_n1029), .ZN(new_n1030));
  NAND2_X1  g0830(.A1(new_n1026), .A2(new_n1030), .ZN(new_n1031));
  NAND2_X1  g0831(.A1(new_n1031), .A2(new_n1018), .ZN(new_n1032));
  NAND3_X1  g0832(.A1(new_n1026), .A2(new_n1030), .A3(new_n675), .ZN(new_n1033));
  NAND2_X1  g0833(.A1(new_n1032), .A2(new_n1033), .ZN(new_n1034));
  INV_X1    g0834(.A(KEYINPUT108), .ZN(new_n1035));
  NAND2_X1  g0835(.A1(new_n666), .A2(new_n1035), .ZN(new_n1036));
  NOR2_X1   g0836(.A1(new_n674), .A2(new_n996), .ZN(new_n1037));
  NOR2_X1   g0837(.A1(new_n1037), .A2(new_n677), .ZN(new_n1038));
  INV_X1    g0838(.A(new_n1038), .ZN(new_n1039));
  NAND2_X1  g0839(.A1(new_n1036), .A2(new_n1039), .ZN(new_n1040));
  NAND3_X1  g0840(.A1(new_n666), .A2(new_n1038), .A3(new_n1035), .ZN(new_n1041));
  NAND2_X1  g0841(.A1(new_n1040), .A2(new_n1041), .ZN(new_n1042));
  INV_X1    g0842(.A(new_n1042), .ZN(new_n1043));
  OAI21_X1  g0843(.A(new_n740), .B1(new_n1034), .B2(new_n1043), .ZN(new_n1044));
  XOR2_X1   g0844(.A(new_n684), .B(KEYINPUT41), .Z(new_n1045));
  INV_X1    g0845(.A(new_n1045), .ZN(new_n1046));
  AOI21_X1  g0846(.A(new_n744), .B1(new_n1044), .B2(new_n1046), .ZN(new_n1047));
  OAI21_X1  g0847(.A(new_n994), .B1(new_n1020), .B2(new_n1047), .ZN(new_n1048));
  INV_X1    g0848(.A(KEYINPUT111), .ZN(new_n1049));
  XNOR2_X1  g0849(.A(new_n1048), .B(new_n1049), .ZN(new_n1050));
  INV_X1    g0850(.A(new_n1050), .ZN(G387));
  NAND2_X1  g0851(.A1(new_n1043), .A2(new_n739), .ZN(new_n1052));
  NAND3_X1  g0852(.A1(new_n1042), .A2(new_n722), .A3(new_n738), .ZN(new_n1053));
  NAND3_X1  g0853(.A1(new_n1052), .A2(new_n684), .A3(new_n1053), .ZN(new_n1054));
  AOI22_X1  g0854(.A1(new_n749), .A2(new_n686), .B1(new_n206), .B2(new_n683), .ZN(new_n1055));
  NOR2_X1   g0855(.A1(new_n236), .A2(new_n264), .ZN(new_n1056));
  NAND2_X1  g0856(.A1(new_n375), .A2(new_n202), .ZN(new_n1057));
  XNOR2_X1  g0857(.A(new_n1057), .B(KEYINPUT50), .ZN(new_n1058));
  OAI211_X1 g0858(.A(new_n687), .B(new_n264), .C1(new_n318), .C2(new_n254), .ZN(new_n1059));
  OAI21_X1  g0859(.A(new_n752), .B1(new_n1058), .B2(new_n1059), .ZN(new_n1060));
  OAI21_X1  g0860(.A(new_n1055), .B1(new_n1056), .B2(new_n1060), .ZN(new_n1061));
  NAND2_X1  g0861(.A1(new_n1061), .A2(new_n761), .ZN(new_n1062));
  NAND2_X1  g0862(.A1(new_n1062), .A2(new_n745), .ZN(new_n1063));
  NOR2_X1   g0863(.A1(new_n674), .A2(new_n812), .ZN(new_n1064));
  AOI22_X1  g0864(.A1(G159), .A2(new_n795), .B1(new_n797), .B2(new_n293), .ZN(new_n1065));
  OAI22_X1  g0865(.A1(new_n792), .A2(new_n202), .B1(new_n800), .B2(new_n318), .ZN(new_n1066));
  INV_X1    g0866(.A(new_n766), .ZN(new_n1067));
  AOI21_X1  g0867(.A(new_n1066), .B1(G150), .B2(new_n1067), .ZN(new_n1068));
  NOR2_X1   g0868(.A1(new_n790), .A2(new_n377), .ZN(new_n1069));
  OAI21_X1  g0869(.A(new_n484), .B1(new_n205), .B2(new_n772), .ZN(new_n1070));
  AOI211_X1 g0870(.A(new_n1069), .B(new_n1070), .C1(G77), .C2(new_n770), .ZN(new_n1071));
  NAND3_X1  g0871(.A1(new_n1065), .A2(new_n1068), .A3(new_n1071), .ZN(new_n1072));
  AOI21_X1  g0872(.A(new_n484), .B1(G326), .B2(new_n1067), .ZN(new_n1073));
  OAI22_X1  g0873(.A1(new_n790), .A2(new_n805), .B1(new_n769), .B2(new_n837), .ZN(new_n1074));
  AOI22_X1  g0874(.A1(new_n786), .A2(G303), .B1(G317), .B2(new_n791), .ZN(new_n1075));
  INV_X1    g0875(.A(G322), .ZN(new_n1076));
  OAI221_X1 g0876(.A(new_n1075), .B1(new_n801), .B2(new_n782), .C1(new_n1076), .C2(new_n781), .ZN(new_n1077));
  INV_X1    g0877(.A(KEYINPUT48), .ZN(new_n1078));
  AOI21_X1  g0878(.A(new_n1074), .B1(new_n1077), .B2(new_n1078), .ZN(new_n1079));
  OAI21_X1  g0879(.A(new_n1079), .B1(new_n1078), .B2(new_n1077), .ZN(new_n1080));
  INV_X1    g0880(.A(KEYINPUT49), .ZN(new_n1081));
  OAI221_X1 g0881(.A(new_n1073), .B1(new_n510), .B2(new_n772), .C1(new_n1080), .C2(new_n1081), .ZN(new_n1082));
  AND2_X1   g0882(.A1(new_n1080), .A2(new_n1081), .ZN(new_n1083));
  OAI21_X1  g0883(.A(new_n1072), .B1(new_n1082), .B2(new_n1083), .ZN(new_n1084));
  AOI211_X1 g0884(.A(new_n1063), .B(new_n1064), .C1(new_n760), .C2(new_n1084), .ZN(new_n1085));
  AOI21_X1  g0885(.A(new_n1085), .B1(new_n1042), .B2(new_n744), .ZN(new_n1086));
  NAND2_X1  g0886(.A1(new_n1054), .A2(new_n1086), .ZN(G393));
  INV_X1    g0887(.A(new_n1033), .ZN(new_n1088));
  AOI21_X1  g0888(.A(new_n675), .B1(new_n1026), .B2(new_n1030), .ZN(new_n1089));
  NOR2_X1   g0889(.A1(new_n1088), .A2(new_n1089), .ZN(new_n1090));
  NAND2_X1  g0890(.A1(new_n1001), .A2(new_n759), .ZN(new_n1091));
  NOR2_X1   g0891(.A1(new_n244), .A2(new_n753), .ZN(new_n1092));
  OAI21_X1  g0892(.A(new_n761), .B1(new_n205), .B2(new_n213), .ZN(new_n1093));
  OAI21_X1  g0893(.A(new_n745), .B1(new_n1092), .B2(new_n1093), .ZN(new_n1094));
  OAI22_X1  g0894(.A1(new_n781), .A2(new_n844), .B1(new_n767), .B2(new_n792), .ZN(new_n1095));
  XNOR2_X1  g0895(.A(new_n1095), .B(KEYINPUT51), .ZN(new_n1096));
  INV_X1    g0896(.A(G143), .ZN(new_n1097));
  OAI21_X1  g0897(.A(new_n484), .B1(new_n1097), .B2(new_n766), .ZN(new_n1098));
  OAI221_X1 g0898(.A(new_n839), .B1(new_n222), .B2(new_n769), .C1(new_n254), .C2(new_n790), .ZN(new_n1099));
  AOI211_X1 g0899(.A(new_n1098), .B(new_n1099), .C1(new_n375), .C2(new_n786), .ZN(new_n1100));
  OAI211_X1 g0900(.A(new_n1096), .B(new_n1100), .C1(new_n202), .C2(new_n782), .ZN(new_n1101));
  INV_X1    g0901(.A(KEYINPUT112), .ZN(new_n1102));
  OR2_X1    g0902(.A1(new_n1101), .A2(new_n1102), .ZN(new_n1103));
  OAI22_X1  g0903(.A1(new_n781), .A2(new_n978), .B1(new_n801), .B2(new_n792), .ZN(new_n1104));
  XNOR2_X1  g0904(.A(new_n1104), .B(KEYINPUT52), .ZN(new_n1105));
  OAI221_X1 g0905(.A(new_n251), .B1(new_n766), .B2(new_n1076), .C1(new_n837), .C2(new_n800), .ZN(new_n1106));
  OAI221_X1 g0906(.A(new_n774), .B1(new_n805), .B2(new_n769), .C1(new_n510), .C2(new_n790), .ZN(new_n1107));
  AOI211_X1 g0907(.A(new_n1106), .B(new_n1107), .C1(G303), .C2(new_n797), .ZN(new_n1108));
  NAND2_X1  g0908(.A1(new_n1105), .A2(new_n1108), .ZN(new_n1109));
  NAND2_X1  g0909(.A1(new_n1101), .A2(new_n1102), .ZN(new_n1110));
  NAND3_X1  g0910(.A1(new_n1103), .A2(new_n1109), .A3(new_n1110), .ZN(new_n1111));
  AOI21_X1  g0911(.A(new_n1094), .B1(new_n1111), .B2(new_n760), .ZN(new_n1112));
  AOI22_X1  g0912(.A1(new_n1090), .A2(new_n744), .B1(new_n1091), .B2(new_n1112), .ZN(new_n1113));
  AND2_X1   g0913(.A1(new_n1034), .A2(new_n1053), .ZN(new_n1114));
  OAI21_X1  g0914(.A(new_n684), .B1(new_n1034), .B2(new_n1053), .ZN(new_n1115));
  OAI21_X1  g0915(.A(new_n1113), .B1(new_n1114), .B2(new_n1115), .ZN(G390));
  NAND2_X1  g0916(.A1(new_n937), .A2(new_n890), .ZN(new_n1117));
  NAND2_X1  g0917(.A1(new_n819), .A2(new_n382), .ZN(new_n1118));
  NAND3_X1  g0918(.A1(new_n734), .A2(new_n659), .A3(new_n1118), .ZN(new_n1119));
  AND2_X1   g0919(.A1(new_n1119), .A2(new_n943), .ZN(new_n1120));
  INV_X1    g0920(.A(new_n927), .ZN(new_n1121));
  OAI211_X1 g0921(.A(new_n953), .B(new_n1117), .C1(new_n1120), .C2(new_n1121), .ZN(new_n1122));
  NAND2_X1  g0922(.A1(new_n907), .A2(new_n893), .ZN(new_n1123));
  NAND2_X1  g0923(.A1(new_n905), .A2(KEYINPUT37), .ZN(new_n1124));
  AOI22_X1  g0924(.A1(new_n1124), .A2(new_n871), .B1(new_n466), .B2(new_n885), .ZN(new_n1125));
  AOI21_X1  g0925(.A(KEYINPUT104), .B1(new_n1125), .B2(KEYINPUT38), .ZN(new_n1126));
  OAI21_X1  g0926(.A(KEYINPUT39), .B1(new_n1123), .B2(new_n1126), .ZN(new_n1127));
  NAND3_X1  g0927(.A1(new_n937), .A2(new_n949), .A3(new_n890), .ZN(new_n1128));
  NAND2_X1  g0928(.A1(new_n1127), .A2(new_n1128), .ZN(new_n1129));
  AOI21_X1  g0929(.A(new_n952), .B1(new_n946), .B2(new_n927), .ZN(new_n1130));
  OAI21_X1  g0930(.A(new_n1122), .B1(new_n1129), .B2(new_n1130), .ZN(new_n1131));
  AND2_X1   g0931(.A1(new_n927), .A2(new_n820), .ZN(new_n1132));
  AND3_X1   g0932(.A1(new_n1132), .A2(G330), .A3(new_n912), .ZN(new_n1133));
  NAND2_X1  g0933(.A1(new_n1131), .A2(new_n1133), .ZN(new_n1134));
  OAI211_X1 g0934(.A(new_n820), .B(new_n927), .C1(new_n720), .C2(new_n721), .ZN(new_n1135));
  OAI211_X1 g0935(.A(new_n1122), .B(new_n1135), .C1(new_n1129), .C2(new_n1130), .ZN(new_n1136));
  NAND3_X1  g0936(.A1(new_n1134), .A2(new_n744), .A3(new_n1136), .ZN(new_n1137));
  OAI21_X1  g0937(.A(new_n745), .B1(new_n831), .B2(new_n293), .ZN(new_n1138));
  AOI22_X1  g0938(.A1(new_n795), .A2(G283), .B1(G97), .B2(new_n786), .ZN(new_n1139));
  OAI21_X1  g0939(.A(new_n1139), .B1(new_n206), .B2(new_n782), .ZN(new_n1140));
  XNOR2_X1  g0940(.A(new_n1140), .B(KEYINPUT115), .ZN(new_n1141));
  OAI21_X1  g0941(.A(new_n251), .B1(new_n766), .B2(new_n837), .ZN(new_n1142));
  AOI21_X1  g0942(.A(new_n1142), .B1(new_n791), .B2(G116), .ZN(new_n1143));
  AOI22_X1  g0943(.A1(new_n770), .A2(G87), .B1(new_n773), .B2(G68), .ZN(new_n1144));
  OAI211_X1 g0944(.A(new_n1143), .B(new_n1144), .C1(new_n254), .C2(new_n790), .ZN(new_n1145));
  NOR2_X1   g0945(.A1(new_n769), .A2(new_n844), .ZN(new_n1146));
  XNOR2_X1  g0946(.A(new_n1146), .B(KEYINPUT53), .ZN(new_n1147));
  XNOR2_X1  g0947(.A(KEYINPUT54), .B(G143), .ZN(new_n1148));
  OAI21_X1  g0948(.A(new_n1147), .B1(new_n787), .B2(new_n1148), .ZN(new_n1149));
  OAI22_X1  g0949(.A1(new_n790), .A2(new_n767), .B1(new_n772), .B2(new_n202), .ZN(new_n1150));
  OAI21_X1  g0950(.A(new_n255), .B1(new_n792), .B2(new_n848), .ZN(new_n1151));
  AOI211_X1 g0951(.A(new_n1150), .B(new_n1151), .C1(G125), .C2(new_n1067), .ZN(new_n1152));
  NAND2_X1  g0952(.A1(new_n795), .A2(G128), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n797), .A2(G137), .ZN(new_n1154));
  NAND3_X1  g0954(.A1(new_n1152), .A2(new_n1153), .A3(new_n1154), .ZN(new_n1155));
  OAI22_X1  g0955(.A1(new_n1141), .A2(new_n1145), .B1(new_n1149), .B2(new_n1155), .ZN(new_n1156));
  OR2_X1    g0956(.A1(new_n1156), .A2(KEYINPUT116), .ZN(new_n1157));
  AOI21_X1  g0957(.A(new_n834), .B1(new_n1156), .B2(KEYINPUT116), .ZN(new_n1158));
  AOI21_X1  g0958(.A(new_n1138), .B1(new_n1157), .B2(new_n1158), .ZN(new_n1159));
  OAI21_X1  g0959(.A(new_n1159), .B1(new_n1129), .B2(new_n758), .ZN(new_n1160));
  NAND3_X1  g0960(.A1(new_n912), .A2(G330), .A3(new_n820), .ZN(new_n1161));
  NAND2_X1  g0961(.A1(new_n1161), .A2(new_n1121), .ZN(new_n1162));
  NAND2_X1  g0962(.A1(new_n1162), .A2(KEYINPUT113), .ZN(new_n1163));
  INV_X1    g0963(.A(KEYINPUT113), .ZN(new_n1164));
  NAND3_X1  g0964(.A1(new_n1161), .A2(new_n1164), .A3(new_n1121), .ZN(new_n1165));
  NAND4_X1  g0965(.A1(new_n1135), .A2(new_n1120), .A3(new_n1163), .A4(new_n1165), .ZN(new_n1166));
  OAI21_X1  g0966(.A(new_n820), .B1(new_n720), .B2(new_n721), .ZN(new_n1167));
  AOI21_X1  g0967(.A(new_n1133), .B1(new_n1167), .B2(new_n1121), .ZN(new_n1168));
  AOI21_X1  g0968(.A(new_n818), .B1(new_n822), .B2(new_n823), .ZN(new_n1169));
  OAI21_X1  g0969(.A(new_n1166), .B1(new_n1168), .B2(new_n1169), .ZN(new_n1170));
  NAND3_X1  g0970(.A1(new_n471), .A2(G330), .A3(new_n912), .ZN(new_n1171));
  AND3_X1   g0971(.A1(new_n1171), .A2(new_n649), .A3(new_n955), .ZN(new_n1172));
  NAND2_X1  g0972(.A1(new_n1170), .A2(new_n1172), .ZN(new_n1173));
  AOI21_X1  g0973(.A(new_n1121), .B1(new_n1119), .B2(new_n943), .ZN(new_n1174));
  NAND2_X1  g0974(.A1(new_n1117), .A2(new_n953), .ZN(new_n1175));
  NOR2_X1   g0975(.A1(new_n1174), .A2(new_n1175), .ZN(new_n1176));
  OAI21_X1  g0976(.A(new_n953), .B1(new_n1169), .B2(new_n1121), .ZN(new_n1177));
  AOI21_X1  g0977(.A(new_n1176), .B1(new_n1177), .B2(new_n951), .ZN(new_n1178));
  NAND3_X1  g0978(.A1(new_n1132), .A2(G330), .A3(new_n912), .ZN(new_n1179));
  OAI21_X1  g0979(.A(new_n1136), .B1(new_n1178), .B2(new_n1179), .ZN(new_n1180));
  NAND2_X1  g0980(.A1(new_n1173), .A2(new_n1180), .ZN(new_n1181));
  NAND4_X1  g0981(.A1(new_n1170), .A2(new_n1134), .A3(new_n1136), .A4(new_n1172), .ZN(new_n1182));
  NAND2_X1  g0982(.A1(new_n1182), .A2(new_n684), .ZN(new_n1183));
  INV_X1    g0983(.A(KEYINPUT114), .ZN(new_n1184));
  OAI21_X1  g0984(.A(new_n1181), .B1(new_n1183), .B2(new_n1184), .ZN(new_n1185));
  AOI21_X1  g0985(.A(KEYINPUT114), .B1(new_n1182), .B2(new_n684), .ZN(new_n1186));
  OAI211_X1 g0986(.A(new_n1137), .B(new_n1160), .C1(new_n1185), .C2(new_n1186), .ZN(G378));
  AOI21_X1  g0987(.A(new_n746), .B1(new_n202), .B2(new_n830), .ZN(new_n1188));
  NAND2_X1  g0988(.A1(new_n418), .A2(new_n263), .ZN(new_n1189));
  OAI22_X1  g0989(.A1(new_n792), .A2(new_n206), .B1(new_n377), .B2(new_n800), .ZN(new_n1190));
  AOI211_X1 g0990(.A(new_n1189), .B(new_n1190), .C1(G283), .C2(new_n1067), .ZN(new_n1191));
  NOR2_X1   g0991(.A1(new_n772), .A2(new_n396), .ZN(new_n1192));
  AOI211_X1 g0992(.A(new_n1192), .B(new_n972), .C1(G77), .C2(new_n770), .ZN(new_n1193));
  AOI22_X1  g0993(.A1(G97), .A2(new_n797), .B1(new_n795), .B2(G116), .ZN(new_n1194));
  NAND3_X1  g0994(.A1(new_n1191), .A2(new_n1193), .A3(new_n1194), .ZN(new_n1195));
  XNOR2_X1  g0995(.A(new_n1195), .B(KEYINPUT117), .ZN(new_n1196));
  OR2_X1    g0996(.A1(new_n1196), .A2(KEYINPUT58), .ZN(new_n1197));
  NAND2_X1  g0997(.A1(new_n791), .A2(G128), .ZN(new_n1198));
  OAI221_X1 g0998(.A(new_n1198), .B1(new_n800), .B2(new_n843), .C1(new_n790), .C2(new_n844), .ZN(new_n1199));
  INV_X1    g0999(.A(new_n1148), .ZN(new_n1200));
  AOI21_X1  g1000(.A(new_n1199), .B1(new_n770), .B2(new_n1200), .ZN(new_n1201));
  NAND2_X1  g1001(.A1(new_n795), .A2(G125), .ZN(new_n1202));
  OAI211_X1 g1002(.A(new_n1201), .B(new_n1202), .C1(new_n848), .C2(new_n782), .ZN(new_n1203));
  OR2_X1    g1003(.A1(new_n1203), .A2(KEYINPUT59), .ZN(new_n1204));
  NAND2_X1  g1004(.A1(new_n1203), .A2(KEYINPUT59), .ZN(new_n1205));
  NAND2_X1  g1005(.A1(new_n773), .A2(G159), .ZN(new_n1206));
  AOI211_X1 g1006(.A(G33), .B(G41), .C1(new_n1067), .C2(G124), .ZN(new_n1207));
  NAND4_X1  g1007(.A1(new_n1204), .A2(new_n1205), .A3(new_n1206), .A4(new_n1207), .ZN(new_n1208));
  OAI211_X1 g1008(.A(new_n1189), .B(new_n202), .C1(G33), .C2(G41), .ZN(new_n1209));
  NAND2_X1  g1009(.A1(new_n1196), .A2(KEYINPUT58), .ZN(new_n1210));
  AND4_X1   g1010(.A1(new_n1197), .A2(new_n1208), .A3(new_n1209), .A4(new_n1210), .ZN(new_n1211));
  OAI21_X1  g1011(.A(new_n1188), .B1(new_n1211), .B2(new_n834), .ZN(new_n1212));
  INV_X1    g1012(.A(new_n305), .ZN(new_n1213));
  NAND2_X1  g1013(.A1(new_n648), .A2(new_n1213), .ZN(new_n1214));
  NOR2_X1   g1014(.A1(new_n298), .A2(new_n656), .ZN(new_n1215));
  NAND2_X1  g1015(.A1(new_n1214), .A2(new_n1215), .ZN(new_n1216));
  OAI211_X1 g1016(.A(new_n648), .B(new_n1213), .C1(new_n298), .C2(new_n656), .ZN(new_n1217));
  XNOR2_X1  g1017(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1218));
  AND3_X1   g1018(.A1(new_n1216), .A2(new_n1217), .A3(new_n1218), .ZN(new_n1219));
  AOI21_X1  g1019(.A(new_n1218), .B1(new_n1216), .B2(new_n1217), .ZN(new_n1220));
  NOR2_X1   g1020(.A1(new_n1219), .A2(new_n1220), .ZN(new_n1221));
  AOI21_X1  g1021(.A(new_n1212), .B1(new_n1221), .B2(new_n757), .ZN(new_n1222));
  AOI21_X1  g1022(.A(new_n866), .B1(new_n928), .B2(new_n938), .ZN(new_n1223));
  NAND3_X1  g1023(.A1(new_n912), .A2(new_n927), .A3(new_n820), .ZN(new_n1224));
  AND2_X1   g1024(.A1(new_n907), .A2(new_n893), .ZN(new_n1225));
  AOI21_X1  g1025(.A(new_n1224), .B1(new_n1225), .B2(new_n892), .ZN(new_n1226));
  OAI211_X1 g1026(.A(new_n1223), .B(new_n1221), .C1(new_n1226), .C2(KEYINPUT40), .ZN(new_n1227));
  OR2_X1    g1027(.A1(new_n1219), .A2(new_n1220), .ZN(new_n1228));
  AND3_X1   g1028(.A1(new_n888), .A2(KEYINPUT38), .A3(new_n889), .ZN(new_n1229));
  AOI21_X1  g1029(.A(KEYINPUT38), .B1(new_n932), .B2(new_n935), .ZN(new_n1230));
  OAI21_X1  g1030(.A(KEYINPUT40), .B1(new_n1229), .B2(new_n1230), .ZN(new_n1231));
  OAI21_X1  g1031(.A(G330), .B1(new_n1231), .B2(new_n1224), .ZN(new_n1232));
  OAI21_X1  g1032(.A(new_n1228), .B1(new_n929), .B2(new_n1232), .ZN(new_n1233));
  NAND3_X1  g1033(.A1(new_n954), .A2(new_n1227), .A3(new_n1233), .ZN(new_n1234));
  INV_X1    g1034(.A(KEYINPUT118), .ZN(new_n1235));
  AND2_X1   g1035(.A1(new_n1234), .A2(new_n1235), .ZN(new_n1236));
  NAND2_X1  g1036(.A1(new_n1233), .A2(new_n1227), .ZN(new_n1237));
  NAND2_X1  g1037(.A1(new_n947), .A2(new_n948), .ZN(new_n1238));
  AOI21_X1  g1038(.A(new_n953), .B1(new_n1127), .B2(new_n1128), .ZN(new_n1239));
  NOR2_X1   g1039(.A1(new_n1238), .A2(new_n1239), .ZN(new_n1240));
  NAND2_X1  g1040(.A1(new_n1237), .A2(new_n1240), .ZN(new_n1241));
  NAND2_X1  g1041(.A1(new_n1241), .A2(KEYINPUT119), .ZN(new_n1242));
  INV_X1    g1042(.A(KEYINPUT119), .ZN(new_n1243));
  NAND3_X1  g1043(.A1(new_n1237), .A2(new_n1243), .A3(new_n1240), .ZN(new_n1244));
  NAND3_X1  g1044(.A1(new_n1236), .A2(new_n1242), .A3(new_n1244), .ZN(new_n1245));
  NAND2_X1  g1045(.A1(new_n1234), .A2(new_n1235), .ZN(new_n1246));
  AND3_X1   g1046(.A1(new_n1237), .A2(new_n1243), .A3(new_n1240), .ZN(new_n1247));
  AOI21_X1  g1047(.A(new_n1243), .B1(new_n1237), .B2(new_n1240), .ZN(new_n1248));
  OAI21_X1  g1048(.A(new_n1246), .B1(new_n1247), .B2(new_n1248), .ZN(new_n1249));
  NAND2_X1  g1049(.A1(new_n1245), .A2(new_n1249), .ZN(new_n1250));
  AOI21_X1  g1050(.A(new_n1222), .B1(new_n1250), .B2(new_n744), .ZN(new_n1251));
  NAND2_X1  g1051(.A1(new_n1241), .A2(new_n1234), .ZN(new_n1252));
  AND2_X1   g1052(.A1(new_n1252), .A2(KEYINPUT57), .ZN(new_n1253));
  NAND2_X1  g1053(.A1(new_n719), .A2(G330), .ZN(new_n1254));
  INV_X1    g1054(.A(KEYINPUT90), .ZN(new_n1255));
  NAND2_X1  g1055(.A1(new_n1254), .A2(new_n1255), .ZN(new_n1256));
  NAND3_X1  g1056(.A1(new_n719), .A2(KEYINPUT90), .A3(G330), .ZN(new_n1257));
  AOI21_X1  g1057(.A(new_n821), .B1(new_n1256), .B2(new_n1257), .ZN(new_n1258));
  OAI21_X1  g1058(.A(new_n1179), .B1(new_n1258), .B2(new_n927), .ZN(new_n1259));
  NAND2_X1  g1059(.A1(new_n1165), .A2(new_n1120), .ZN(new_n1260));
  AOI21_X1  g1060(.A(new_n1164), .B1(new_n1161), .B2(new_n1121), .ZN(new_n1261));
  NOR2_X1   g1061(.A1(new_n1260), .A2(new_n1261), .ZN(new_n1262));
  AOI22_X1  g1062(.A1(new_n946), .A2(new_n1259), .B1(new_n1262), .B2(new_n1135), .ZN(new_n1263));
  OAI211_X1 g1063(.A(KEYINPUT120), .B(new_n1172), .C1(new_n1180), .C2(new_n1263), .ZN(new_n1264));
  INV_X1    g1064(.A(new_n1264), .ZN(new_n1265));
  AOI21_X1  g1065(.A(KEYINPUT120), .B1(new_n1182), .B2(new_n1172), .ZN(new_n1266));
  OAI21_X1  g1066(.A(new_n1253), .B1(new_n1265), .B2(new_n1266), .ZN(new_n1267));
  NAND2_X1  g1067(.A1(new_n1267), .A2(new_n684), .ZN(new_n1268));
  OAI21_X1  g1068(.A(new_n1172), .B1(new_n1180), .B2(new_n1263), .ZN(new_n1269));
  INV_X1    g1069(.A(KEYINPUT120), .ZN(new_n1270));
  NAND2_X1  g1070(.A1(new_n1269), .A2(new_n1270), .ZN(new_n1271));
  NAND2_X1  g1071(.A1(new_n1271), .A2(new_n1264), .ZN(new_n1272));
  AOI21_X1  g1072(.A(KEYINPUT57), .B1(new_n1250), .B2(new_n1272), .ZN(new_n1273));
  OAI21_X1  g1073(.A(new_n1251), .B1(new_n1268), .B2(new_n1273), .ZN(G375));
  INV_X1    g1074(.A(new_n1172), .ZN(new_n1275));
  NAND2_X1  g1075(.A1(new_n1263), .A2(new_n1275), .ZN(new_n1276));
  NAND3_X1  g1076(.A1(new_n1276), .A2(new_n1046), .A3(new_n1173), .ZN(new_n1277));
  NAND2_X1  g1077(.A1(new_n1121), .A2(new_n757), .ZN(new_n1278));
  OAI21_X1  g1078(.A(new_n745), .B1(new_n831), .B2(G68), .ZN(new_n1279));
  OAI21_X1  g1079(.A(new_n251), .B1(new_n792), .B2(new_n805), .ZN(new_n1280));
  AOI21_X1  g1080(.A(new_n1280), .B1(G303), .B2(new_n1067), .ZN(new_n1281));
  NAND2_X1  g1081(.A1(new_n770), .A2(G97), .ZN(new_n1282));
  NOR2_X1   g1082(.A1(new_n1069), .A2(new_n971), .ZN(new_n1283));
  NAND2_X1  g1083(.A1(new_n786), .A2(G107), .ZN(new_n1284));
  NAND4_X1  g1084(.A1(new_n1281), .A2(new_n1282), .A3(new_n1283), .A4(new_n1284), .ZN(new_n1285));
  OAI22_X1  g1085(.A1(new_n510), .A2(new_n782), .B1(new_n781), .B2(new_n837), .ZN(new_n1286));
  OAI22_X1  g1086(.A1(new_n792), .A2(new_n843), .B1(new_n800), .B2(new_n844), .ZN(new_n1287));
  AOI21_X1  g1087(.A(new_n1287), .B1(G128), .B2(new_n1067), .ZN(new_n1288));
  NOR2_X1   g1088(.A1(new_n1192), .A2(new_n418), .ZN(new_n1289));
  AOI22_X1  g1089(.A1(new_n807), .A2(G50), .B1(new_n770), .B2(G159), .ZN(new_n1290));
  NAND3_X1  g1090(.A1(new_n1288), .A2(new_n1289), .A3(new_n1290), .ZN(new_n1291));
  OAI22_X1  g1091(.A1(new_n848), .A2(new_n781), .B1(new_n782), .B2(new_n1148), .ZN(new_n1292));
  OAI22_X1  g1092(.A1(new_n1285), .A2(new_n1286), .B1(new_n1291), .B2(new_n1292), .ZN(new_n1293));
  AOI21_X1  g1093(.A(new_n1279), .B1(new_n1293), .B2(new_n760), .ZN(new_n1294));
  AOI22_X1  g1094(.A1(new_n1170), .A2(new_n744), .B1(new_n1278), .B2(new_n1294), .ZN(new_n1295));
  NAND2_X1  g1095(.A1(new_n1277), .A2(new_n1295), .ZN(G381));
  INV_X1    g1096(.A(G384), .ZN(new_n1297));
  NAND3_X1  g1097(.A1(new_n1054), .A2(new_n814), .A3(new_n1086), .ZN(new_n1298));
  INV_X1    g1098(.A(new_n1298), .ZN(new_n1299));
  NAND2_X1  g1099(.A1(new_n1297), .A2(new_n1299), .ZN(new_n1300));
  XNOR2_X1  g1100(.A(new_n1300), .B(KEYINPUT121), .ZN(new_n1301));
  NOR4_X1   g1101(.A1(G387), .A2(new_n1301), .A3(G390), .A4(G381), .ZN(new_n1302));
  NAND2_X1  g1102(.A1(new_n1137), .A2(new_n1160), .ZN(new_n1303));
  INV_X1    g1103(.A(new_n1185), .ZN(new_n1304));
  INV_X1    g1104(.A(new_n1186), .ZN(new_n1305));
  AOI21_X1  g1105(.A(new_n1303), .B1(new_n1304), .B2(new_n1305), .ZN(new_n1306));
  NAND2_X1  g1106(.A1(G375), .A2(KEYINPUT122), .ZN(new_n1307));
  OR2_X1    g1107(.A1(G375), .A2(KEYINPUT122), .ZN(new_n1308));
  NAND4_X1  g1108(.A1(new_n1302), .A2(new_n1306), .A3(new_n1307), .A4(new_n1308), .ZN(G407));
  NAND2_X1  g1109(.A1(new_n657), .A2(G213), .ZN(new_n1310));
  INV_X1    g1110(.A(new_n1310), .ZN(new_n1311));
  NAND4_X1  g1111(.A1(new_n1308), .A2(new_n1306), .A3(new_n1307), .A4(new_n1311), .ZN(new_n1312));
  NAND3_X1  g1112(.A1(G407), .A2(new_n1312), .A3(G213), .ZN(new_n1313));
  XOR2_X1   g1113(.A(new_n1313), .B(KEYINPUT123), .Z(G409));
  INV_X1    g1114(.A(KEYINPUT126), .ZN(new_n1315));
  AOI21_X1  g1115(.A(new_n814), .B1(new_n1054), .B2(new_n1086), .ZN(new_n1316));
  OAI21_X1  g1116(.A(G390), .B1(new_n1299), .B2(new_n1316), .ZN(new_n1317));
  NAND2_X1  g1117(.A1(G393), .A2(G396), .ZN(new_n1318));
  AOI21_X1  g1118(.A(new_n1049), .B1(new_n1318), .B2(new_n1298), .ZN(new_n1319));
  OAI21_X1  g1119(.A(new_n1317), .B1(new_n1319), .B2(G390), .ZN(new_n1320));
  INV_X1    g1120(.A(new_n1048), .ZN(new_n1321));
  NAND2_X1  g1121(.A1(new_n1320), .A2(new_n1321), .ZN(new_n1322));
  OAI211_X1 g1122(.A(new_n1048), .B(new_n1317), .C1(G390), .C2(new_n1319), .ZN(new_n1323));
  AND2_X1   g1123(.A1(new_n1322), .A2(new_n1323), .ZN(new_n1324));
  XOR2_X1   g1124(.A(new_n1324), .B(KEYINPUT125), .Z(new_n1325));
  INV_X1    g1125(.A(KEYINPUT62), .ZN(new_n1326));
  OAI211_X1 g1126(.A(G378), .B(new_n1251), .C1(new_n1268), .C2(new_n1273), .ZN(new_n1327));
  NAND3_X1  g1127(.A1(new_n1250), .A2(new_n1272), .A3(new_n1046), .ZN(new_n1328));
  AOI21_X1  g1128(.A(new_n1222), .B1(new_n1252), .B2(new_n744), .ZN(new_n1329));
  NAND2_X1  g1129(.A1(new_n1328), .A2(new_n1329), .ZN(new_n1330));
  NAND2_X1  g1130(.A1(new_n1330), .A2(new_n1306), .ZN(new_n1331));
  NAND2_X1  g1131(.A1(new_n1327), .A2(new_n1331), .ZN(new_n1332));
  NAND2_X1  g1132(.A1(new_n1173), .A2(KEYINPUT60), .ZN(new_n1333));
  NAND2_X1  g1133(.A1(new_n1333), .A2(new_n1276), .ZN(new_n1334));
  NAND3_X1  g1134(.A1(new_n1263), .A2(new_n1275), .A3(KEYINPUT60), .ZN(new_n1335));
  NAND3_X1  g1135(.A1(new_n1334), .A2(new_n684), .A3(new_n1335), .ZN(new_n1336));
  NAND3_X1  g1136(.A1(new_n1336), .A2(G384), .A3(new_n1295), .ZN(new_n1337));
  INV_X1    g1137(.A(new_n1337), .ZN(new_n1338));
  AOI21_X1  g1138(.A(G384), .B1(new_n1336), .B2(new_n1295), .ZN(new_n1339));
  NOR2_X1   g1139(.A1(new_n1338), .A2(new_n1339), .ZN(new_n1340));
  AND4_X1   g1140(.A1(new_n1326), .A2(new_n1332), .A3(new_n1310), .A4(new_n1340), .ZN(new_n1341));
  INV_X1    g1141(.A(KEYINPUT61), .ZN(new_n1342));
  AOI21_X1  g1142(.A(new_n1311), .B1(new_n1327), .B2(new_n1331), .ZN(new_n1343));
  NAND2_X1  g1143(.A1(new_n1311), .A2(G2897), .ZN(new_n1344));
  INV_X1    g1144(.A(new_n1344), .ZN(new_n1345));
  OAI21_X1  g1145(.A(new_n1345), .B1(new_n1338), .B2(new_n1339), .ZN(new_n1346));
  INV_X1    g1146(.A(new_n1339), .ZN(new_n1347));
  NAND3_X1  g1147(.A1(new_n1347), .A2(new_n1337), .A3(new_n1344), .ZN(new_n1348));
  NAND2_X1  g1148(.A1(new_n1346), .A2(new_n1348), .ZN(new_n1349));
  OAI21_X1  g1149(.A(new_n1342), .B1(new_n1343), .B2(new_n1349), .ZN(new_n1350));
  NOR2_X1   g1150(.A1(new_n1341), .A2(new_n1350), .ZN(new_n1351));
  AOI21_X1  g1151(.A(new_n1326), .B1(new_n1343), .B2(new_n1340), .ZN(new_n1352));
  INV_X1    g1152(.A(new_n1352), .ZN(new_n1353));
  AOI21_X1  g1153(.A(new_n1325), .B1(new_n1351), .B2(new_n1353), .ZN(new_n1354));
  NAND3_X1  g1154(.A1(new_n1322), .A2(new_n1323), .A3(new_n1342), .ZN(new_n1355));
  XNOR2_X1  g1155(.A(new_n1355), .B(KEYINPUT124), .ZN(new_n1356));
  OAI21_X1  g1156(.A(new_n1356), .B1(new_n1343), .B2(new_n1349), .ZN(new_n1357));
  NAND3_X1  g1157(.A1(new_n1343), .A2(KEYINPUT63), .A3(new_n1340), .ZN(new_n1358));
  INV_X1    g1158(.A(new_n1358), .ZN(new_n1359));
  AOI21_X1  g1159(.A(KEYINPUT63), .B1(new_n1343), .B2(new_n1340), .ZN(new_n1360));
  NOR3_X1   g1160(.A1(new_n1357), .A2(new_n1359), .A3(new_n1360), .ZN(new_n1361));
  OAI21_X1  g1161(.A(new_n1315), .B1(new_n1354), .B2(new_n1361), .ZN(new_n1362));
  INV_X1    g1162(.A(new_n1360), .ZN(new_n1363));
  OR2_X1    g1163(.A1(new_n1343), .A2(new_n1349), .ZN(new_n1364));
  NAND4_X1  g1164(.A1(new_n1363), .A2(new_n1364), .A3(new_n1358), .A4(new_n1356), .ZN(new_n1365));
  NOR3_X1   g1165(.A1(new_n1341), .A2(new_n1350), .A3(new_n1352), .ZN(new_n1366));
  OAI211_X1 g1166(.A(new_n1365), .B(KEYINPUT126), .C1(new_n1366), .C2(new_n1325), .ZN(new_n1367));
  NAND2_X1  g1167(.A1(new_n1362), .A2(new_n1367), .ZN(G405));
  NAND2_X1  g1168(.A1(G375), .A2(new_n1306), .ZN(new_n1369));
  NAND2_X1  g1169(.A1(new_n1369), .A2(new_n1327), .ZN(new_n1370));
  NAND2_X1  g1170(.A1(new_n1340), .A2(KEYINPUT127), .ZN(new_n1371));
  XNOR2_X1  g1171(.A(new_n1370), .B(new_n1371), .ZN(new_n1372));
  XNOR2_X1  g1172(.A(new_n1372), .B(new_n1324), .ZN(G402));
endmodule


