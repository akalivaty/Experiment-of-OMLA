

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n511, n512, n513, n514,
         n515, n516, n517, n518, n519, n520, n521, n522, n523, n524, n525,
         n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536,
         n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547,
         n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558,
         n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569,
         n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580,
         n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591,
         n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602,
         n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, n613,
         n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624,
         n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635,
         n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, n646,
         n647, n648, n649, n650, n651, n652, n653, n654, n655, n656, n657,
         n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668,
         n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679,
         n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690,
         n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701,
         n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712,
         n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723,
         n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, n734,
         n735, n736, n737, n738, n739, n740, n741, n742, n743, n744, n745,
         n746, n747, n748, n749, n750, n751, n752, n753, n754, n755, n756,
         n757, n758, n759, n760, n761, n762, n763, n764, n765, n766, n767,
         n768, n769, n770, n771, n772, n773, n774, n775, n776, n777, n778,
         n779, n780, n781, n782, n783, n784, n785, n786, n787, n788, n789,
         n790, n791, n792, n793, n794, n795, n796, n797, n798, n799, n800,
         n801, n802, n803, n804, n805, n806, n807, n808, n809, n810, n811,
         n812, n813, n814, n815, n816, n817, n818, n819, n820, n821, n822,
         n823, n824, n825, n826, n827, n828, n829, n830, n831, n832, n833,
         n834, n835, n836, n837, n838, n839, n840, n841, n842, n843, n844,
         n845, n846, n847, n848, n849, n850, n851, n852, n853, n854, n855,
         n856, n857, n858, n859, n860, n861, n862, n863, n864, n865, n866,
         n867, n868, n869, n870, n871, n872, n873, n874, n875, n876, n877,
         n878, n879, n880, n881, n882, n883, n884, n885, n886, n887, n888,
         n889, n890, n891, n892, n893, n894, n895, n896, n897, n898, n899,
         n900, n901, n902, n903, n904, n905, n906, n907, n908, n909, n910,
         n911, n912, n913, n914, n915, n916, n917, n918, n919, n920, n921,
         n922, n923, n924, n925, n926, n927, n928, n929, n930, n931, n932,
         n933, n934, n935, n936, n937, n938, n939, n940, n941, n942, n943,
         n944, n945, n946, n947, n948, n949, n950, n951, n952, n953, n954,
         n955, n956, n957, n958, n959, n960, n961, n962, n963, n964, n965,
         n966, n967, n968, n969, n970, n971, n972, n973, n974, n975, n976,
         n977, n978, n979, n980, n981, n982, n983, n984, n985, n986, n987,
         n988, n989, n990, n991, n992, n993, n994, n995, n996, n997, n998,
         n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008,
         n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018,
         n1019, n1020, n1021, n1022, n1023;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NOR2_X1 U547 ( .A1(n686), .A2(n685), .ZN(n779) );
  XOR2_X1 U548 ( .A(G543), .B(KEYINPUT0), .Z(n511) );
  NAND2_X1 U549 ( .A1(n779), .A2(n781), .ZN(n730) );
  INV_X1 U550 ( .A(KEYINPUT98), .ZN(n740) );
  XNOR2_X1 U551 ( .A(n767), .B(KEYINPUT100), .ZN(n769) );
  INV_X1 U552 ( .A(n1013), .ZN(n768) );
  AND2_X1 U553 ( .A1(n551), .A2(G2104), .ZN(n872) );
  NAND2_X1 U554 ( .A1(n873), .A2(G137), .ZN(n557) );
  OR2_X1 U555 ( .A1(n776), .A2(n775), .ZN(n512) );
  AND2_X1 U556 ( .A1(n777), .A2(n512), .ZN(n513) );
  AND2_X1 U557 ( .A1(n698), .A2(n697), .ZN(n514) );
  XOR2_X1 U558 ( .A(KEYINPUT96), .B(n706), .Z(n515) );
  AND2_X1 U559 ( .A1(n514), .A2(n701), .ZN(n702) );
  AND2_X1 U560 ( .A1(n781), .A2(n779), .ZN(n716) );
  OR2_X1 U561 ( .A1(n722), .A2(n721), .ZN(n745) );
  XNOR2_X1 U562 ( .A(n741), .B(n740), .ZN(n742) );
  INV_X1 U563 ( .A(KEYINPUT17), .ZN(n547) );
  XNOR2_X1 U564 ( .A(n548), .B(n547), .ZN(n873) );
  XNOR2_X1 U565 ( .A(KEYINPUT65), .B(KEYINPUT23), .ZN(n560) );
  NOR2_X1 U566 ( .A1(n523), .A2(n645), .ZN(n655) );
  XNOR2_X1 U567 ( .A(n561), .B(n560), .ZN(n563) );
  NAND2_X1 U568 ( .A1(n585), .A2(n584), .ZN(n1009) );
  NOR2_X1 U569 ( .A1(G651), .A2(G543), .ZN(n648) );
  NAND2_X1 U570 ( .A1(n648), .A2(G90), .ZN(n516) );
  XNOR2_X1 U571 ( .A(n516), .B(KEYINPUT72), .ZN(n518) );
  INV_X1 U572 ( .A(G651), .ZN(n523) );
  XNOR2_X1 U573 ( .A(KEYINPUT68), .B(n511), .ZN(n645) );
  NAND2_X1 U574 ( .A1(G77), .A2(n655), .ZN(n517) );
  NAND2_X1 U575 ( .A1(n518), .A2(n517), .ZN(n519) );
  XNOR2_X1 U576 ( .A(n519), .B(KEYINPUT9), .ZN(n522) );
  NOR2_X1 U577 ( .A1(G651), .A2(n645), .ZN(n520) );
  XNOR2_X1 U578 ( .A(KEYINPUT64), .B(n520), .ZN(n588) );
  NAND2_X1 U579 ( .A1(G52), .A2(n588), .ZN(n521) );
  NAND2_X1 U580 ( .A1(n522), .A2(n521), .ZN(n528) );
  NOR2_X1 U581 ( .A1(G543), .A2(n523), .ZN(n525) );
  XNOR2_X1 U582 ( .A(KEYINPUT1), .B(KEYINPUT69), .ZN(n524) );
  XNOR2_X1 U583 ( .A(n525), .B(n524), .ZN(n649) );
  NAND2_X1 U584 ( .A1(G64), .A2(n649), .ZN(n526) );
  XNOR2_X1 U585 ( .A(KEYINPUT71), .B(n526), .ZN(n527) );
  NOR2_X1 U586 ( .A1(n528), .A2(n527), .ZN(G171) );
  XOR2_X1 U587 ( .A(KEYINPUT102), .B(G2446), .Z(n530) );
  XNOR2_X1 U588 ( .A(KEYINPUT103), .B(G2451), .ZN(n529) );
  XNOR2_X1 U589 ( .A(n530), .B(n529), .ZN(n534) );
  XOR2_X1 U590 ( .A(KEYINPUT104), .B(G2438), .Z(n532) );
  XNOR2_X1 U591 ( .A(G2435), .B(G2454), .ZN(n531) );
  XNOR2_X1 U592 ( .A(n532), .B(n531), .ZN(n533) );
  XOR2_X1 U593 ( .A(n534), .B(n533), .Z(n536) );
  XNOR2_X1 U594 ( .A(G2443), .B(G2427), .ZN(n535) );
  XNOR2_X1 U595 ( .A(n536), .B(n535), .ZN(n539) );
  XNOR2_X1 U596 ( .A(G1348), .B(G2430), .ZN(n537) );
  INV_X1 U597 ( .A(G1341), .ZN(n694) );
  XNOR2_X1 U598 ( .A(n537), .B(n694), .ZN(n538) );
  XOR2_X1 U599 ( .A(n539), .B(n538), .Z(n540) );
  AND2_X1 U600 ( .A1(G14), .A2(n540), .ZN(G401) );
  AND2_X1 U601 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U602 ( .A(G57), .ZN(G237) );
  INV_X1 U603 ( .A(G132), .ZN(G219) );
  INV_X1 U604 ( .A(G82), .ZN(G220) );
  NAND2_X1 U605 ( .A1(G88), .A2(n648), .ZN(n542) );
  NAND2_X1 U606 ( .A1(G75), .A2(n655), .ZN(n541) );
  NAND2_X1 U607 ( .A1(n542), .A2(n541), .ZN(n546) );
  NAND2_X1 U608 ( .A1(G62), .A2(n649), .ZN(n544) );
  NAND2_X1 U609 ( .A1(G50), .A2(n588), .ZN(n543) );
  NAND2_X1 U610 ( .A1(n544), .A2(n543), .ZN(n545) );
  NOR2_X1 U611 ( .A1(n546), .A2(n545), .ZN(G166) );
  INV_X1 U612 ( .A(G2105), .ZN(n551) );
  NAND2_X1 U613 ( .A1(G102), .A2(n872), .ZN(n550) );
  NOR2_X1 U614 ( .A1(G2104), .A2(G2105), .ZN(n548) );
  NAND2_X1 U615 ( .A1(G138), .A2(n873), .ZN(n549) );
  NAND2_X1 U616 ( .A1(n550), .A2(n549), .ZN(n555) );
  AND2_X1 U617 ( .A1(G2104), .A2(G2105), .ZN(n876) );
  NAND2_X1 U618 ( .A1(G114), .A2(n876), .ZN(n553) );
  NOR2_X1 U619 ( .A1(G2104), .A2(n551), .ZN(n877) );
  NAND2_X1 U620 ( .A1(G126), .A2(n877), .ZN(n552) );
  NAND2_X1 U621 ( .A1(n553), .A2(n552), .ZN(n554) );
  NOR2_X1 U622 ( .A1(n555), .A2(n554), .ZN(G164) );
  NAND2_X1 U623 ( .A1(G113), .A2(n876), .ZN(n556) );
  XNOR2_X1 U624 ( .A(n556), .B(KEYINPUT66), .ZN(n559) );
  XOR2_X1 U625 ( .A(KEYINPUT67), .B(n557), .Z(n558) );
  NAND2_X1 U626 ( .A1(n559), .A2(n558), .ZN(n685) );
  NAND2_X1 U627 ( .A1(G101), .A2(n872), .ZN(n561) );
  NAND2_X1 U628 ( .A1(G125), .A2(n877), .ZN(n562) );
  NAND2_X1 U629 ( .A1(n563), .A2(n562), .ZN(n683) );
  NOR2_X1 U630 ( .A1(n685), .A2(n683), .ZN(G160) );
  NAND2_X1 U631 ( .A1(n648), .A2(G89), .ZN(n564) );
  XNOR2_X1 U632 ( .A(n564), .B(KEYINPUT4), .ZN(n566) );
  NAND2_X1 U633 ( .A1(G76), .A2(n655), .ZN(n565) );
  NAND2_X1 U634 ( .A1(n566), .A2(n565), .ZN(n567) );
  XNOR2_X1 U635 ( .A(n567), .B(KEYINPUT5), .ZN(n572) );
  NAND2_X1 U636 ( .A1(G63), .A2(n649), .ZN(n569) );
  NAND2_X1 U637 ( .A1(G51), .A2(n588), .ZN(n568) );
  NAND2_X1 U638 ( .A1(n569), .A2(n568), .ZN(n570) );
  XOR2_X1 U639 ( .A(KEYINPUT6), .B(n570), .Z(n571) );
  NAND2_X1 U640 ( .A1(n572), .A2(n571), .ZN(n573) );
  XNOR2_X1 U641 ( .A(n573), .B(KEYINPUT7), .ZN(G168) );
  XOR2_X1 U642 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U643 ( .A1(G7), .A2(G661), .ZN(n574) );
  XNOR2_X1 U644 ( .A(n574), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U645 ( .A(G223), .ZN(n831) );
  NAND2_X1 U646 ( .A1(n831), .A2(G567), .ZN(n575) );
  XOR2_X1 U647 ( .A(KEYINPUT11), .B(n575), .Z(G234) );
  NAND2_X1 U648 ( .A1(G68), .A2(n655), .ZN(n578) );
  NAND2_X1 U649 ( .A1(n648), .A2(G81), .ZN(n576) );
  XNOR2_X1 U650 ( .A(n576), .B(KEYINPUT12), .ZN(n577) );
  NAND2_X1 U651 ( .A1(n578), .A2(n577), .ZN(n580) );
  XOR2_X1 U652 ( .A(KEYINPUT13), .B(KEYINPUT76), .Z(n579) );
  XNOR2_X1 U653 ( .A(n580), .B(n579), .ZN(n583) );
  NAND2_X1 U654 ( .A1(n649), .A2(G56), .ZN(n581) );
  XOR2_X1 U655 ( .A(KEYINPUT14), .B(n581), .Z(n582) );
  NOR2_X1 U656 ( .A1(n583), .A2(n582), .ZN(n585) );
  NAND2_X1 U657 ( .A1(G43), .A2(n588), .ZN(n584) );
  INV_X1 U658 ( .A(G860), .ZN(n608) );
  OR2_X1 U659 ( .A1(n1009), .A2(n608), .ZN(G153) );
  XNOR2_X1 U660 ( .A(G171), .B(KEYINPUT77), .ZN(G301) );
  NAND2_X1 U661 ( .A1(G868), .A2(G301), .ZN(n597) );
  INV_X1 U662 ( .A(KEYINPUT78), .ZN(n595) );
  NAND2_X1 U663 ( .A1(G92), .A2(n648), .ZN(n587) );
  NAND2_X1 U664 ( .A1(G79), .A2(n655), .ZN(n586) );
  NAND2_X1 U665 ( .A1(n587), .A2(n586), .ZN(n592) );
  NAND2_X1 U666 ( .A1(G66), .A2(n649), .ZN(n590) );
  NAND2_X1 U667 ( .A1(G54), .A2(n588), .ZN(n589) );
  NAND2_X1 U668 ( .A1(n590), .A2(n589), .ZN(n591) );
  NOR2_X1 U669 ( .A1(n592), .A2(n591), .ZN(n593) );
  XNOR2_X1 U670 ( .A(KEYINPUT15), .B(n593), .ZN(n594) );
  XNOR2_X1 U671 ( .A(n595), .B(n594), .ZN(n691) );
  BUF_X1 U672 ( .A(n691), .Z(n994) );
  OR2_X1 U673 ( .A1(n994), .A2(G868), .ZN(n596) );
  NAND2_X1 U674 ( .A1(n597), .A2(n596), .ZN(G284) );
  NAND2_X1 U675 ( .A1(G78), .A2(n655), .ZN(n598) );
  XNOR2_X1 U676 ( .A(n598), .B(KEYINPUT74), .ZN(n601) );
  NAND2_X1 U677 ( .A1(G91), .A2(n648), .ZN(n599) );
  XOR2_X1 U678 ( .A(KEYINPUT73), .B(n599), .Z(n600) );
  NAND2_X1 U679 ( .A1(n601), .A2(n600), .ZN(n605) );
  NAND2_X1 U680 ( .A1(G65), .A2(n649), .ZN(n603) );
  NAND2_X1 U681 ( .A1(G53), .A2(n588), .ZN(n602) );
  NAND2_X1 U682 ( .A1(n603), .A2(n602), .ZN(n604) );
  NOR2_X1 U683 ( .A1(n605), .A2(n604), .ZN(n1001) );
  XNOR2_X1 U684 ( .A(n1001), .B(KEYINPUT75), .ZN(G299) );
  NAND2_X1 U685 ( .A1(G286), .A2(G868), .ZN(n607) );
  INV_X1 U686 ( .A(G868), .ZN(n666) );
  NAND2_X1 U687 ( .A1(G299), .A2(n666), .ZN(n606) );
  NAND2_X1 U688 ( .A1(n607), .A2(n606), .ZN(G297) );
  NAND2_X1 U689 ( .A1(n608), .A2(G559), .ZN(n609) );
  NAND2_X1 U690 ( .A1(n609), .A2(n994), .ZN(n610) );
  XNOR2_X1 U691 ( .A(n610), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U692 ( .A1(G868), .A2(n1009), .ZN(n613) );
  NAND2_X1 U693 ( .A1(n994), .A2(G868), .ZN(n611) );
  NOR2_X1 U694 ( .A1(G559), .A2(n611), .ZN(n612) );
  NOR2_X1 U695 ( .A1(n613), .A2(n612), .ZN(G282) );
  XOR2_X1 U696 ( .A(G2100), .B(KEYINPUT80), .Z(n623) );
  NAND2_X1 U697 ( .A1(G99), .A2(n872), .ZN(n615) );
  NAND2_X1 U698 ( .A1(G111), .A2(n876), .ZN(n614) );
  NAND2_X1 U699 ( .A1(n615), .A2(n614), .ZN(n616) );
  XNOR2_X1 U700 ( .A(n616), .B(KEYINPUT79), .ZN(n618) );
  NAND2_X1 U701 ( .A1(G135), .A2(n873), .ZN(n617) );
  NAND2_X1 U702 ( .A1(n618), .A2(n617), .ZN(n621) );
  NAND2_X1 U703 ( .A1(n877), .A2(G123), .ZN(n619) );
  XOR2_X1 U704 ( .A(KEYINPUT18), .B(n619), .Z(n620) );
  NOR2_X1 U705 ( .A1(n621), .A2(n620), .ZN(n959) );
  XNOR2_X1 U706 ( .A(G2096), .B(n959), .ZN(n622) );
  NAND2_X1 U707 ( .A1(n623), .A2(n622), .ZN(G156) );
  NAND2_X1 U708 ( .A1(G67), .A2(n649), .ZN(n625) );
  NAND2_X1 U709 ( .A1(G55), .A2(n588), .ZN(n624) );
  NAND2_X1 U710 ( .A1(n625), .A2(n624), .ZN(n626) );
  XNOR2_X1 U711 ( .A(KEYINPUT82), .B(n626), .ZN(n630) );
  NAND2_X1 U712 ( .A1(G93), .A2(n648), .ZN(n628) );
  NAND2_X1 U713 ( .A1(G80), .A2(n655), .ZN(n627) );
  NAND2_X1 U714 ( .A1(n628), .A2(n627), .ZN(n629) );
  OR2_X1 U715 ( .A1(n630), .A2(n629), .ZN(n665) );
  NAND2_X1 U716 ( .A1(n994), .A2(G559), .ZN(n631) );
  XOR2_X1 U717 ( .A(n1009), .B(n631), .Z(n663) );
  XNOR2_X1 U718 ( .A(KEYINPUT81), .B(n663), .ZN(n632) );
  NOR2_X1 U719 ( .A1(G860), .A2(n632), .ZN(n633) );
  XOR2_X1 U720 ( .A(n665), .B(n633), .Z(G145) );
  NAND2_X1 U721 ( .A1(G73), .A2(n655), .ZN(n634) );
  XOR2_X1 U722 ( .A(KEYINPUT2), .B(n634), .Z(n639) );
  NAND2_X1 U723 ( .A1(G86), .A2(n648), .ZN(n636) );
  NAND2_X1 U724 ( .A1(G61), .A2(n649), .ZN(n635) );
  NAND2_X1 U725 ( .A1(n636), .A2(n635), .ZN(n637) );
  XOR2_X1 U726 ( .A(KEYINPUT83), .B(n637), .Z(n638) );
  NOR2_X1 U727 ( .A1(n639), .A2(n638), .ZN(n641) );
  NAND2_X1 U728 ( .A1(G48), .A2(n588), .ZN(n640) );
  NAND2_X1 U729 ( .A1(n641), .A2(n640), .ZN(G305) );
  NAND2_X1 U730 ( .A1(G651), .A2(G74), .ZN(n643) );
  NAND2_X1 U731 ( .A1(G49), .A2(n588), .ZN(n642) );
  NAND2_X1 U732 ( .A1(n643), .A2(n642), .ZN(n644) );
  NOR2_X1 U733 ( .A1(n649), .A2(n644), .ZN(n647) );
  NAND2_X1 U734 ( .A1(G87), .A2(n645), .ZN(n646) );
  NAND2_X1 U735 ( .A1(n647), .A2(n646), .ZN(G288) );
  NAND2_X1 U736 ( .A1(G85), .A2(n648), .ZN(n651) );
  NAND2_X1 U737 ( .A1(G60), .A2(n649), .ZN(n650) );
  NAND2_X1 U738 ( .A1(n651), .A2(n650), .ZN(n654) );
  NAND2_X1 U739 ( .A1(n588), .A2(G47), .ZN(n652) );
  XOR2_X1 U740 ( .A(KEYINPUT70), .B(n652), .Z(n653) );
  NOR2_X1 U741 ( .A1(n654), .A2(n653), .ZN(n657) );
  NAND2_X1 U742 ( .A1(n655), .A2(G72), .ZN(n656) );
  NAND2_X1 U743 ( .A1(n657), .A2(n656), .ZN(G290) );
  XOR2_X1 U744 ( .A(n665), .B(G305), .Z(n658) );
  XNOR2_X1 U745 ( .A(n658), .B(G288), .ZN(n659) );
  XNOR2_X1 U746 ( .A(KEYINPUT19), .B(n659), .ZN(n661) );
  XNOR2_X1 U747 ( .A(G290), .B(G166), .ZN(n660) );
  XNOR2_X1 U748 ( .A(n661), .B(n660), .ZN(n662) );
  XNOR2_X1 U749 ( .A(n662), .B(G299), .ZN(n895) );
  XNOR2_X1 U750 ( .A(n663), .B(n895), .ZN(n664) );
  NAND2_X1 U751 ( .A1(n664), .A2(G868), .ZN(n668) );
  NAND2_X1 U752 ( .A1(n666), .A2(n665), .ZN(n667) );
  NAND2_X1 U753 ( .A1(n668), .A2(n667), .ZN(G295) );
  NAND2_X1 U754 ( .A1(G2078), .A2(G2084), .ZN(n669) );
  XOR2_X1 U755 ( .A(KEYINPUT20), .B(n669), .Z(n670) );
  NAND2_X1 U756 ( .A1(G2090), .A2(n670), .ZN(n672) );
  XNOR2_X1 U757 ( .A(KEYINPUT21), .B(KEYINPUT84), .ZN(n671) );
  XNOR2_X1 U758 ( .A(n672), .B(n671), .ZN(n673) );
  NAND2_X1 U759 ( .A1(G2072), .A2(n673), .ZN(G158) );
  XNOR2_X1 U760 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U761 ( .A1(G220), .A2(G219), .ZN(n674) );
  XOR2_X1 U762 ( .A(KEYINPUT22), .B(n674), .Z(n675) );
  NOR2_X1 U763 ( .A1(G218), .A2(n675), .ZN(n676) );
  XOR2_X1 U764 ( .A(KEYINPUT85), .B(n676), .Z(n677) );
  NAND2_X1 U765 ( .A1(G96), .A2(n677), .ZN(n907) );
  NAND2_X1 U766 ( .A1(n907), .A2(G2106), .ZN(n681) );
  NAND2_X1 U767 ( .A1(G69), .A2(G120), .ZN(n678) );
  NOR2_X1 U768 ( .A1(G237), .A2(n678), .ZN(n679) );
  NAND2_X1 U769 ( .A1(G108), .A2(n679), .ZN(n908) );
  NAND2_X1 U770 ( .A1(n908), .A2(G567), .ZN(n680) );
  NAND2_X1 U771 ( .A1(n681), .A2(n680), .ZN(n835) );
  NAND2_X1 U772 ( .A1(G661), .A2(G483), .ZN(n682) );
  NOR2_X1 U773 ( .A1(n835), .A2(n682), .ZN(n834) );
  NAND2_X1 U774 ( .A1(n834), .A2(G36), .ZN(G176) );
  INV_X1 U775 ( .A(G166), .ZN(G303) );
  NOR2_X1 U776 ( .A1(G164), .A2(G1384), .ZN(n781) );
  INV_X1 U777 ( .A(n683), .ZN(n684) );
  NAND2_X1 U778 ( .A1(G40), .A2(n684), .ZN(n686) );
  NAND2_X1 U779 ( .A1(n716), .A2(G2067), .ZN(n688) );
  NAND2_X1 U780 ( .A1(G1348), .A2(n730), .ZN(n687) );
  NAND2_X1 U781 ( .A1(n688), .A2(n687), .ZN(n689) );
  XNOR2_X1 U782 ( .A(n689), .B(KEYINPUT95), .ZN(n690) );
  NAND2_X1 U783 ( .A1(n690), .A2(n691), .ZN(n705) );
  INV_X1 U784 ( .A(n690), .ZN(n693) );
  INV_X1 U785 ( .A(n691), .ZN(n692) );
  NAND2_X1 U786 ( .A1(n693), .A2(n692), .ZN(n703) );
  XNOR2_X1 U787 ( .A(KEYINPUT26), .B(KEYINPUT94), .ZN(n699) );
  NAND2_X1 U788 ( .A1(n694), .A2(n699), .ZN(n695) );
  NAND2_X1 U789 ( .A1(n695), .A2(n730), .ZN(n698) );
  AND2_X1 U790 ( .A1(n716), .A2(G1996), .ZN(n696) );
  NAND2_X1 U791 ( .A1(n696), .A2(n699), .ZN(n697) );
  NOR2_X1 U792 ( .A1(G1996), .A2(n699), .ZN(n700) );
  NOR2_X1 U793 ( .A1(n700), .A2(n1009), .ZN(n701) );
  NAND2_X1 U794 ( .A1(n703), .A2(n702), .ZN(n704) );
  NAND2_X1 U795 ( .A1(n705), .A2(n704), .ZN(n706) );
  NAND2_X1 U796 ( .A1(n716), .A2(G2072), .ZN(n707) );
  XNOR2_X1 U797 ( .A(n707), .B(KEYINPUT27), .ZN(n709) );
  AND2_X1 U798 ( .A1(G1956), .A2(n730), .ZN(n708) );
  NOR2_X1 U799 ( .A1(n709), .A2(n708), .ZN(n711) );
  NAND2_X1 U800 ( .A1(n711), .A2(n1001), .ZN(n710) );
  NAND2_X1 U801 ( .A1(n515), .A2(n710), .ZN(n714) );
  NOR2_X1 U802 ( .A1(n711), .A2(n1001), .ZN(n712) );
  XOR2_X1 U803 ( .A(n712), .B(KEYINPUT28), .Z(n713) );
  NAND2_X1 U804 ( .A1(n714), .A2(n713), .ZN(n715) );
  XNOR2_X1 U805 ( .A(n715), .B(KEYINPUT29), .ZN(n722) );
  XOR2_X1 U806 ( .A(G2078), .B(KEYINPUT25), .Z(n942) );
  NAND2_X1 U807 ( .A1(n716), .A2(n942), .ZN(n718) );
  NAND2_X1 U808 ( .A1(G1961), .A2(n730), .ZN(n717) );
  NAND2_X1 U809 ( .A1(n718), .A2(n717), .ZN(n719) );
  XOR2_X1 U810 ( .A(KEYINPUT92), .B(n719), .Z(n726) );
  NAND2_X1 U811 ( .A1(G171), .A2(n726), .ZN(n720) );
  XNOR2_X1 U812 ( .A(KEYINPUT93), .B(n720), .ZN(n721) );
  NAND2_X1 U813 ( .A1(G8), .A2(n730), .ZN(n776) );
  NOR2_X1 U814 ( .A1(G1966), .A2(n776), .ZN(n748) );
  NOR2_X1 U815 ( .A1(G2084), .A2(n730), .ZN(n744) );
  NOR2_X1 U816 ( .A1(n748), .A2(n744), .ZN(n723) );
  NAND2_X1 U817 ( .A1(G8), .A2(n723), .ZN(n724) );
  XNOR2_X1 U818 ( .A(KEYINPUT30), .B(n724), .ZN(n725) );
  NOR2_X1 U819 ( .A1(G168), .A2(n725), .ZN(n728) );
  NOR2_X1 U820 ( .A1(G171), .A2(n726), .ZN(n727) );
  NOR2_X1 U821 ( .A1(n728), .A2(n727), .ZN(n729) );
  XOR2_X1 U822 ( .A(KEYINPUT31), .B(n729), .Z(n746) );
  NOR2_X1 U823 ( .A1(G2090), .A2(n730), .ZN(n731) );
  XOR2_X1 U824 ( .A(KEYINPUT97), .B(n731), .Z(n733) );
  NOR2_X1 U825 ( .A1(G1971), .A2(n776), .ZN(n732) );
  NOR2_X1 U826 ( .A1(n733), .A2(n732), .ZN(n734) );
  NAND2_X1 U827 ( .A1(n734), .A2(G303), .ZN(n736) );
  AND2_X1 U828 ( .A1(n746), .A2(n736), .ZN(n735) );
  NAND2_X1 U829 ( .A1(n745), .A2(n735), .ZN(n739) );
  INV_X1 U830 ( .A(n736), .ZN(n737) );
  OR2_X1 U831 ( .A1(n737), .A2(G286), .ZN(n738) );
  NAND2_X1 U832 ( .A1(n739), .A2(n738), .ZN(n741) );
  NAND2_X1 U833 ( .A1(n742), .A2(G8), .ZN(n743) );
  XNOR2_X1 U834 ( .A(n743), .B(KEYINPUT32), .ZN(n752) );
  NAND2_X1 U835 ( .A1(G8), .A2(n744), .ZN(n750) );
  AND2_X1 U836 ( .A1(n746), .A2(n745), .ZN(n747) );
  NOR2_X1 U837 ( .A1(n748), .A2(n747), .ZN(n749) );
  NAND2_X1 U838 ( .A1(n750), .A2(n749), .ZN(n751) );
  NAND2_X1 U839 ( .A1(n752), .A2(n751), .ZN(n754) );
  INV_X1 U840 ( .A(KEYINPUT99), .ZN(n753) );
  XNOR2_X1 U841 ( .A(n754), .B(n753), .ZN(n772) );
  NOR2_X1 U842 ( .A1(G1976), .A2(G288), .ZN(n997) );
  NOR2_X1 U843 ( .A1(G1971), .A2(G303), .ZN(n755) );
  NOR2_X1 U844 ( .A1(n997), .A2(n755), .ZN(n757) );
  INV_X1 U845 ( .A(n776), .ZN(n761) );
  NAND2_X1 U846 ( .A1(n997), .A2(n761), .ZN(n756) );
  NAND2_X1 U847 ( .A1(n756), .A2(KEYINPUT33), .ZN(n759) );
  AND2_X1 U848 ( .A1(n757), .A2(n759), .ZN(n758) );
  NAND2_X1 U849 ( .A1(n772), .A2(n758), .ZN(n766) );
  INV_X1 U850 ( .A(n759), .ZN(n764) );
  INV_X1 U851 ( .A(KEYINPUT33), .ZN(n760) );
  NAND2_X1 U852 ( .A1(G1976), .A2(G288), .ZN(n999) );
  AND2_X1 U853 ( .A1(n760), .A2(n999), .ZN(n762) );
  AND2_X1 U854 ( .A1(n762), .A2(n761), .ZN(n763) );
  OR2_X1 U855 ( .A1(n764), .A2(n763), .ZN(n765) );
  AND2_X1 U856 ( .A1(n766), .A2(n765), .ZN(n767) );
  XNOR2_X1 U857 ( .A(G1981), .B(G305), .ZN(n1013) );
  NAND2_X1 U858 ( .A1(n769), .A2(n768), .ZN(n778) );
  NOR2_X1 U859 ( .A1(G2090), .A2(G303), .ZN(n770) );
  NAND2_X1 U860 ( .A1(G8), .A2(n770), .ZN(n771) );
  NAND2_X1 U861 ( .A1(n772), .A2(n771), .ZN(n773) );
  NAND2_X1 U862 ( .A1(n773), .A2(n776), .ZN(n777) );
  NOR2_X1 U863 ( .A1(G1981), .A2(G305), .ZN(n774) );
  XOR2_X1 U864 ( .A(n774), .B(KEYINPUT24), .Z(n775) );
  NAND2_X1 U865 ( .A1(n778), .A2(n513), .ZN(n815) );
  XNOR2_X1 U866 ( .A(G1986), .B(G290), .ZN(n996) );
  INV_X1 U867 ( .A(n779), .ZN(n780) );
  NOR2_X1 U868 ( .A1(n781), .A2(n780), .ZN(n826) );
  NAND2_X1 U869 ( .A1(n996), .A2(n826), .ZN(n813) );
  NAND2_X1 U870 ( .A1(G117), .A2(n876), .ZN(n783) );
  NAND2_X1 U871 ( .A1(G129), .A2(n877), .ZN(n782) );
  NAND2_X1 U872 ( .A1(n783), .A2(n782), .ZN(n786) );
  NAND2_X1 U873 ( .A1(n872), .A2(G105), .ZN(n784) );
  XOR2_X1 U874 ( .A(KEYINPUT38), .B(n784), .Z(n785) );
  NOR2_X1 U875 ( .A1(n786), .A2(n785), .ZN(n787) );
  XOR2_X1 U876 ( .A(KEYINPUT89), .B(n787), .Z(n789) );
  NAND2_X1 U877 ( .A1(n873), .A2(G141), .ZN(n788) );
  NAND2_X1 U878 ( .A1(n789), .A2(n788), .ZN(n884) );
  NAND2_X1 U879 ( .A1(G1996), .A2(n884), .ZN(n798) );
  NAND2_X1 U880 ( .A1(G95), .A2(n872), .ZN(n791) );
  NAND2_X1 U881 ( .A1(G131), .A2(n873), .ZN(n790) );
  NAND2_X1 U882 ( .A1(n791), .A2(n790), .ZN(n795) );
  NAND2_X1 U883 ( .A1(G107), .A2(n876), .ZN(n793) );
  NAND2_X1 U884 ( .A1(G119), .A2(n877), .ZN(n792) );
  NAND2_X1 U885 ( .A1(n793), .A2(n792), .ZN(n794) );
  NOR2_X1 U886 ( .A1(n795), .A2(n794), .ZN(n887) );
  XNOR2_X1 U887 ( .A(KEYINPUT87), .B(G1991), .ZN(n941) );
  NOR2_X1 U888 ( .A1(n887), .A2(n941), .ZN(n796) );
  XOR2_X1 U889 ( .A(KEYINPUT88), .B(n796), .Z(n797) );
  NAND2_X1 U890 ( .A1(n798), .A2(n797), .ZN(n799) );
  XOR2_X1 U891 ( .A(KEYINPUT90), .B(n799), .Z(n972) );
  XNOR2_X1 U892 ( .A(n826), .B(KEYINPUT91), .ZN(n800) );
  NOR2_X1 U893 ( .A1(n972), .A2(n800), .ZN(n818) );
  INV_X1 U894 ( .A(n818), .ZN(n811) );
  XNOR2_X1 U895 ( .A(KEYINPUT86), .B(KEYINPUT34), .ZN(n804) );
  NAND2_X1 U896 ( .A1(G104), .A2(n872), .ZN(n802) );
  NAND2_X1 U897 ( .A1(G140), .A2(n873), .ZN(n801) );
  NAND2_X1 U898 ( .A1(n802), .A2(n801), .ZN(n803) );
  XNOR2_X1 U899 ( .A(n804), .B(n803), .ZN(n809) );
  NAND2_X1 U900 ( .A1(G116), .A2(n876), .ZN(n806) );
  NAND2_X1 U901 ( .A1(G128), .A2(n877), .ZN(n805) );
  NAND2_X1 U902 ( .A1(n806), .A2(n805), .ZN(n807) );
  XOR2_X1 U903 ( .A(KEYINPUT35), .B(n807), .Z(n808) );
  NOR2_X1 U904 ( .A1(n809), .A2(n808), .ZN(n810) );
  XNOR2_X1 U905 ( .A(KEYINPUT36), .B(n810), .ZN(n891) );
  XNOR2_X1 U906 ( .A(G2067), .B(KEYINPUT37), .ZN(n824) );
  NOR2_X1 U907 ( .A1(n891), .A2(n824), .ZN(n971) );
  NAND2_X1 U908 ( .A1(n826), .A2(n971), .ZN(n821) );
  AND2_X1 U909 ( .A1(n811), .A2(n821), .ZN(n812) );
  AND2_X1 U910 ( .A1(n813), .A2(n812), .ZN(n814) );
  NAND2_X1 U911 ( .A1(n815), .A2(n814), .ZN(n829) );
  NOR2_X1 U912 ( .A1(G1996), .A2(n884), .ZN(n965) );
  NOR2_X1 U913 ( .A1(G1986), .A2(G290), .ZN(n816) );
  AND2_X1 U914 ( .A1(n941), .A2(n887), .ZN(n960) );
  NOR2_X1 U915 ( .A1(n816), .A2(n960), .ZN(n817) );
  NOR2_X1 U916 ( .A1(n818), .A2(n817), .ZN(n819) );
  NOR2_X1 U917 ( .A1(n965), .A2(n819), .ZN(n820) );
  XNOR2_X1 U918 ( .A(n820), .B(KEYINPUT39), .ZN(n822) );
  NAND2_X1 U919 ( .A1(n822), .A2(n821), .ZN(n823) );
  XOR2_X1 U920 ( .A(KEYINPUT101), .B(n823), .Z(n825) );
  NAND2_X1 U921 ( .A1(n891), .A2(n824), .ZN(n975) );
  NAND2_X1 U922 ( .A1(n825), .A2(n975), .ZN(n827) );
  NAND2_X1 U923 ( .A1(n827), .A2(n826), .ZN(n828) );
  NAND2_X1 U924 ( .A1(n829), .A2(n828), .ZN(n830) );
  XNOR2_X1 U925 ( .A(KEYINPUT40), .B(n830), .ZN(G329) );
  NAND2_X1 U926 ( .A1(G2106), .A2(n831), .ZN(G217) );
  AND2_X1 U927 ( .A1(G15), .A2(G2), .ZN(n832) );
  NAND2_X1 U928 ( .A1(G661), .A2(n832), .ZN(G259) );
  NAND2_X1 U929 ( .A1(G3), .A2(G1), .ZN(n833) );
  NAND2_X1 U930 ( .A1(n834), .A2(n833), .ZN(G188) );
  INV_X1 U931 ( .A(n835), .ZN(G319) );
  XOR2_X1 U932 ( .A(G2096), .B(G2100), .Z(n837) );
  XNOR2_X1 U933 ( .A(KEYINPUT42), .B(G2678), .ZN(n836) );
  XNOR2_X1 U934 ( .A(n837), .B(n836), .ZN(n841) );
  XOR2_X1 U935 ( .A(KEYINPUT43), .B(G2072), .Z(n839) );
  XNOR2_X1 U936 ( .A(G2067), .B(G2090), .ZN(n838) );
  XNOR2_X1 U937 ( .A(n839), .B(n838), .ZN(n840) );
  XOR2_X1 U938 ( .A(n841), .B(n840), .Z(n843) );
  XNOR2_X1 U939 ( .A(G2078), .B(G2084), .ZN(n842) );
  XNOR2_X1 U940 ( .A(n843), .B(n842), .ZN(G227) );
  XOR2_X1 U941 ( .A(KEYINPUT106), .B(G1976), .Z(n845) );
  XNOR2_X1 U942 ( .A(G1961), .B(G1956), .ZN(n844) );
  XNOR2_X1 U943 ( .A(n845), .B(n844), .ZN(n846) );
  XOR2_X1 U944 ( .A(n846), .B(KEYINPUT41), .Z(n848) );
  XNOR2_X1 U945 ( .A(G1996), .B(G1991), .ZN(n847) );
  XNOR2_X1 U946 ( .A(n848), .B(n847), .ZN(n852) );
  XOR2_X1 U947 ( .A(G1981), .B(G1971), .Z(n850) );
  XNOR2_X1 U948 ( .A(G1986), .B(G1966), .ZN(n849) );
  XNOR2_X1 U949 ( .A(n850), .B(n849), .ZN(n851) );
  XOR2_X1 U950 ( .A(n852), .B(n851), .Z(n854) );
  XNOR2_X1 U951 ( .A(KEYINPUT105), .B(G2474), .ZN(n853) );
  XNOR2_X1 U952 ( .A(n854), .B(n853), .ZN(G229) );
  NAND2_X1 U953 ( .A1(G124), .A2(n877), .ZN(n855) );
  XNOR2_X1 U954 ( .A(n855), .B(KEYINPUT44), .ZN(n857) );
  NAND2_X1 U955 ( .A1(n872), .A2(G100), .ZN(n856) );
  NAND2_X1 U956 ( .A1(n857), .A2(n856), .ZN(n861) );
  NAND2_X1 U957 ( .A1(G112), .A2(n876), .ZN(n859) );
  NAND2_X1 U958 ( .A1(G136), .A2(n873), .ZN(n858) );
  NAND2_X1 U959 ( .A1(n859), .A2(n858), .ZN(n860) );
  NOR2_X1 U960 ( .A1(n861), .A2(n860), .ZN(G162) );
  XNOR2_X1 U961 ( .A(G164), .B(G162), .ZN(n870) );
  NAND2_X1 U962 ( .A1(G118), .A2(n876), .ZN(n863) );
  NAND2_X1 U963 ( .A1(G130), .A2(n877), .ZN(n862) );
  NAND2_X1 U964 ( .A1(n863), .A2(n862), .ZN(n868) );
  NAND2_X1 U965 ( .A1(G106), .A2(n872), .ZN(n865) );
  NAND2_X1 U966 ( .A1(G142), .A2(n873), .ZN(n864) );
  NAND2_X1 U967 ( .A1(n865), .A2(n864), .ZN(n866) );
  XOR2_X1 U968 ( .A(KEYINPUT45), .B(n866), .Z(n867) );
  NOR2_X1 U969 ( .A1(n868), .A2(n867), .ZN(n869) );
  XNOR2_X1 U970 ( .A(n870), .B(n869), .ZN(n871) );
  XNOR2_X1 U971 ( .A(n959), .B(n871), .ZN(n886) );
  NAND2_X1 U972 ( .A1(G103), .A2(n872), .ZN(n875) );
  NAND2_X1 U973 ( .A1(G139), .A2(n873), .ZN(n874) );
  NAND2_X1 U974 ( .A1(n875), .A2(n874), .ZN(n883) );
  NAND2_X1 U975 ( .A1(G115), .A2(n876), .ZN(n879) );
  NAND2_X1 U976 ( .A1(G127), .A2(n877), .ZN(n878) );
  NAND2_X1 U977 ( .A1(n879), .A2(n878), .ZN(n880) );
  XNOR2_X1 U978 ( .A(KEYINPUT107), .B(n880), .ZN(n881) );
  XNOR2_X1 U979 ( .A(KEYINPUT47), .B(n881), .ZN(n882) );
  NOR2_X1 U980 ( .A1(n883), .A2(n882), .ZN(n978) );
  XNOR2_X1 U981 ( .A(n884), .B(n978), .ZN(n885) );
  XNOR2_X1 U982 ( .A(n886), .B(n885), .ZN(n893) );
  XOR2_X1 U983 ( .A(KEYINPUT46), .B(KEYINPUT48), .Z(n889) );
  XNOR2_X1 U984 ( .A(n887), .B(G160), .ZN(n888) );
  XNOR2_X1 U985 ( .A(n889), .B(n888), .ZN(n890) );
  XNOR2_X1 U986 ( .A(n891), .B(n890), .ZN(n892) );
  XNOR2_X1 U987 ( .A(n893), .B(n892), .ZN(n894) );
  NOR2_X1 U988 ( .A1(G37), .A2(n894), .ZN(G395) );
  XNOR2_X1 U989 ( .A(n895), .B(KEYINPUT108), .ZN(n897) );
  XNOR2_X1 U990 ( .A(n1009), .B(G286), .ZN(n896) );
  XNOR2_X1 U991 ( .A(n897), .B(n896), .ZN(n899) );
  XNOR2_X1 U992 ( .A(n994), .B(G171), .ZN(n898) );
  XNOR2_X1 U993 ( .A(n899), .B(n898), .ZN(n900) );
  NOR2_X1 U994 ( .A1(G37), .A2(n900), .ZN(G397) );
  NOR2_X1 U995 ( .A1(G227), .A2(G229), .ZN(n901) );
  XOR2_X1 U996 ( .A(KEYINPUT49), .B(n901), .Z(n902) );
  NAND2_X1 U997 ( .A1(G319), .A2(n902), .ZN(n903) );
  NOR2_X1 U998 ( .A1(G401), .A2(n903), .ZN(n906) );
  NOR2_X1 U999 ( .A1(G395), .A2(G397), .ZN(n904) );
  XOR2_X1 U1000 ( .A(KEYINPUT109), .B(n904), .Z(n905) );
  NAND2_X1 U1001 ( .A1(n906), .A2(n905), .ZN(G225) );
  XOR2_X1 U1002 ( .A(KEYINPUT110), .B(G225), .Z(G308) );
  INV_X1 U1004 ( .A(G120), .ZN(G236) );
  INV_X1 U1005 ( .A(G96), .ZN(G221) );
  INV_X1 U1006 ( .A(G69), .ZN(G235) );
  NOR2_X1 U1007 ( .A1(n908), .A2(n907), .ZN(G325) );
  INV_X1 U1008 ( .A(G325), .ZN(G261) );
  INV_X1 U1009 ( .A(G108), .ZN(G238) );
  XNOR2_X1 U1010 ( .A(G1971), .B(G22), .ZN(n910) );
  XNOR2_X1 U1011 ( .A(G23), .B(G1976), .ZN(n909) );
  NOR2_X1 U1012 ( .A1(n910), .A2(n909), .ZN(n912) );
  XOR2_X1 U1013 ( .A(G1986), .B(G24), .Z(n911) );
  NAND2_X1 U1014 ( .A1(n912), .A2(n911), .ZN(n914) );
  XNOR2_X1 U1015 ( .A(KEYINPUT127), .B(KEYINPUT58), .ZN(n913) );
  XNOR2_X1 U1016 ( .A(n914), .B(n913), .ZN(n917) );
  XNOR2_X1 U1017 ( .A(G1961), .B(KEYINPUT123), .ZN(n915) );
  XNOR2_X1 U1018 ( .A(n915), .B(G5), .ZN(n916) );
  NAND2_X1 U1019 ( .A1(n917), .A2(n916), .ZN(n932) );
  XOR2_X1 U1020 ( .A(G4), .B(KEYINPUT125), .Z(n919) );
  XNOR2_X1 U1021 ( .A(G1348), .B(KEYINPUT59), .ZN(n918) );
  XNOR2_X1 U1022 ( .A(n919), .B(n918), .ZN(n923) );
  XNOR2_X1 U1023 ( .A(G1956), .B(G20), .ZN(n921) );
  XNOR2_X1 U1024 ( .A(G19), .B(G1341), .ZN(n920) );
  NOR2_X1 U1025 ( .A1(n921), .A2(n920), .ZN(n922) );
  NAND2_X1 U1026 ( .A1(n923), .A2(n922), .ZN(n926) );
  XNOR2_X1 U1027 ( .A(KEYINPUT124), .B(G1981), .ZN(n924) );
  XNOR2_X1 U1028 ( .A(G6), .B(n924), .ZN(n925) );
  NOR2_X1 U1029 ( .A1(n926), .A2(n925), .ZN(n927) );
  XOR2_X1 U1030 ( .A(KEYINPUT60), .B(n927), .Z(n929) );
  XNOR2_X1 U1031 ( .A(G1966), .B(G21), .ZN(n928) );
  NOR2_X1 U1032 ( .A1(n929), .A2(n928), .ZN(n930) );
  XOR2_X1 U1033 ( .A(KEYINPUT126), .B(n930), .Z(n931) );
  NOR2_X1 U1034 ( .A1(n932), .A2(n931), .ZN(n933) );
  XOR2_X1 U1035 ( .A(KEYINPUT61), .B(n933), .Z(n934) );
  NOR2_X1 U1036 ( .A1(G16), .A2(n934), .ZN(n958) );
  XNOR2_X1 U1037 ( .A(KEYINPUT55), .B(KEYINPUT117), .ZN(n987) );
  XNOR2_X1 U1038 ( .A(G2067), .B(G26), .ZN(n936) );
  XNOR2_X1 U1039 ( .A(G33), .B(G2072), .ZN(n935) );
  NOR2_X1 U1040 ( .A1(n936), .A2(n935), .ZN(n937) );
  NAND2_X1 U1041 ( .A1(G28), .A2(n937), .ZN(n940) );
  XOR2_X1 U1042 ( .A(KEYINPUT119), .B(G1996), .Z(n938) );
  XNOR2_X1 U1043 ( .A(G32), .B(n938), .ZN(n939) );
  NOR2_X1 U1044 ( .A1(n940), .A2(n939), .ZN(n946) );
  XOR2_X1 U1045 ( .A(n941), .B(G25), .Z(n944) );
  XNOR2_X1 U1046 ( .A(G27), .B(n942), .ZN(n943) );
  NOR2_X1 U1047 ( .A1(n944), .A2(n943), .ZN(n945) );
  NAND2_X1 U1048 ( .A1(n946), .A2(n945), .ZN(n947) );
  XNOR2_X1 U1049 ( .A(n947), .B(KEYINPUT53), .ZN(n950) );
  XOR2_X1 U1050 ( .A(G2084), .B(G34), .Z(n948) );
  XNOR2_X1 U1051 ( .A(KEYINPUT54), .B(n948), .ZN(n949) );
  NAND2_X1 U1052 ( .A1(n950), .A2(n949), .ZN(n952) );
  XNOR2_X1 U1053 ( .A(G35), .B(G2090), .ZN(n951) );
  NOR2_X1 U1054 ( .A1(n952), .A2(n951), .ZN(n953) );
  XOR2_X1 U1055 ( .A(n987), .B(n953), .Z(n955) );
  INV_X1 U1056 ( .A(G29), .ZN(n954) );
  NAND2_X1 U1057 ( .A1(n955), .A2(n954), .ZN(n956) );
  NAND2_X1 U1058 ( .A1(n956), .A2(G11), .ZN(n957) );
  NOR2_X1 U1059 ( .A1(n958), .A2(n957), .ZN(n992) );
  XNOR2_X1 U1060 ( .A(G160), .B(G2084), .ZN(n962) );
  NOR2_X1 U1061 ( .A1(n960), .A2(n959), .ZN(n961) );
  NAND2_X1 U1062 ( .A1(n962), .A2(n961), .ZN(n963) );
  XNOR2_X1 U1063 ( .A(KEYINPUT111), .B(n963), .ZN(n969) );
  XOR2_X1 U1064 ( .A(G2090), .B(G162), .Z(n964) );
  XNOR2_X1 U1065 ( .A(KEYINPUT112), .B(n964), .ZN(n966) );
  NOR2_X1 U1066 ( .A1(n966), .A2(n965), .ZN(n967) );
  XOR2_X1 U1067 ( .A(KEYINPUT51), .B(n967), .Z(n968) );
  NAND2_X1 U1068 ( .A1(n969), .A2(n968), .ZN(n970) );
  NOR2_X1 U1069 ( .A1(n971), .A2(n970), .ZN(n973) );
  NAND2_X1 U1070 ( .A1(n973), .A2(n972), .ZN(n974) );
  XNOR2_X1 U1071 ( .A(n974), .B(KEYINPUT113), .ZN(n976) );
  NAND2_X1 U1072 ( .A1(n976), .A2(n975), .ZN(n977) );
  XNOR2_X1 U1073 ( .A(KEYINPUT114), .B(n977), .ZN(n985) );
  XOR2_X1 U1074 ( .A(n978), .B(KEYINPUT115), .Z(n979) );
  XOR2_X1 U1075 ( .A(G2072), .B(n979), .Z(n981) );
  XOR2_X1 U1076 ( .A(G164), .B(G2078), .Z(n980) );
  NOR2_X1 U1077 ( .A1(n981), .A2(n980), .ZN(n982) );
  XOR2_X1 U1078 ( .A(KEYINPUT50), .B(n982), .Z(n983) );
  XNOR2_X1 U1079 ( .A(KEYINPUT116), .B(n983), .ZN(n984) );
  NOR2_X1 U1080 ( .A1(n985), .A2(n984), .ZN(n986) );
  XNOR2_X1 U1081 ( .A(n986), .B(KEYINPUT52), .ZN(n988) );
  NAND2_X1 U1082 ( .A1(n988), .A2(n987), .ZN(n989) );
  XNOR2_X1 U1083 ( .A(KEYINPUT118), .B(n989), .ZN(n990) );
  NAND2_X1 U1084 ( .A1(n990), .A2(G29), .ZN(n991) );
  NAND2_X1 U1085 ( .A1(n992), .A2(n991), .ZN(n1022) );
  XOR2_X1 U1086 ( .A(G16), .B(KEYINPUT56), .Z(n993) );
  XNOR2_X1 U1087 ( .A(KEYINPUT120), .B(n993), .ZN(n1020) );
  XOR2_X1 U1088 ( .A(G1348), .B(n994), .Z(n995) );
  NOR2_X1 U1089 ( .A1(n996), .A2(n995), .ZN(n1007) );
  INV_X1 U1090 ( .A(n997), .ZN(n998) );
  NAND2_X1 U1091 ( .A1(n999), .A2(n998), .ZN(n1000) );
  XNOR2_X1 U1092 ( .A(n1000), .B(KEYINPUT122), .ZN(n1005) );
  XNOR2_X1 U1093 ( .A(G1956), .B(n1001), .ZN(n1003) );
  XNOR2_X1 U1094 ( .A(G166), .B(G1971), .ZN(n1002) );
  NAND2_X1 U1095 ( .A1(n1003), .A2(n1002), .ZN(n1004) );
  NOR2_X1 U1096 ( .A1(n1005), .A2(n1004), .ZN(n1006) );
  NAND2_X1 U1097 ( .A1(n1007), .A2(n1006), .ZN(n1018) );
  XNOR2_X1 U1098 ( .A(G171), .B(G1961), .ZN(n1008) );
  XNOR2_X1 U1099 ( .A(n1008), .B(KEYINPUT121), .ZN(n1011) );
  XNOR2_X1 U1100 ( .A(G1341), .B(n1009), .ZN(n1010) );
  NOR2_X1 U1101 ( .A1(n1011), .A2(n1010), .ZN(n1016) );
  XOR2_X1 U1102 ( .A(G168), .B(G1966), .Z(n1012) );
  NOR2_X1 U1103 ( .A1(n1013), .A2(n1012), .ZN(n1014) );
  XOR2_X1 U1104 ( .A(KEYINPUT57), .B(n1014), .Z(n1015) );
  NAND2_X1 U1105 ( .A1(n1016), .A2(n1015), .ZN(n1017) );
  NOR2_X1 U1106 ( .A1(n1018), .A2(n1017), .ZN(n1019) );
  NOR2_X1 U1107 ( .A1(n1020), .A2(n1019), .ZN(n1021) );
  NOR2_X1 U1108 ( .A1(n1022), .A2(n1021), .ZN(n1023) );
  XNOR2_X1 U1109 ( .A(n1023), .B(KEYINPUT62), .ZN(G311) );
  INV_X1 U1110 ( .A(G311), .ZN(G150) );
endmodule

