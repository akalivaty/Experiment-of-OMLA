//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 1 1 0 0 1 0 1 1 0 1 0 1 1 1 1 1 1 0 0 0 0 0 1 1 0 0 1 0 1 0 1 1 1 1 0 0 0 1 0 0 0 1 0 1 0 0 1 1 0 0 0 1 0 1 0 1 1 1 1 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:15:28 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n685,
    new_n686, new_n687, new_n688, new_n689, new_n690, new_n692, new_n693,
    new_n694, new_n696, new_n697, new_n698, new_n699, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n725, new_n726, new_n727, new_n728, new_n729, new_n730, new_n731,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n755,
    new_n756, new_n757, new_n758, new_n760, new_n761, new_n762, new_n764,
    new_n765, new_n766, new_n768, new_n770, new_n771, new_n772, new_n773,
    new_n774, new_n775, new_n776, new_n777, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n786, new_n787, new_n788, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n837, new_n838, new_n840, new_n841, new_n843,
    new_n844, new_n845, new_n846, new_n847, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n904, new_n905, new_n906, new_n908, new_n909, new_n910,
    new_n911, new_n912, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n922, new_n923, new_n924, new_n926, new_n927,
    new_n928, new_n929, new_n930, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n938, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n949, new_n950, new_n951,
    new_n952, new_n954, new_n955, new_n956, new_n957, new_n958, new_n959,
    new_n961, new_n962;
  XNOR2_X1  g000(.A(G113gat), .B(G141gat), .ZN(new_n202));
  XNOR2_X1  g001(.A(KEYINPUT90), .B(KEYINPUT11), .ZN(new_n203));
  XNOR2_X1  g002(.A(new_n202), .B(new_n203), .ZN(new_n204));
  XNOR2_X1  g003(.A(G169gat), .B(G197gat), .ZN(new_n205));
  XNOR2_X1  g004(.A(new_n204), .B(new_n205), .ZN(new_n206));
  XNOR2_X1  g005(.A(new_n206), .B(KEYINPUT12), .ZN(new_n207));
  XOR2_X1   g006(.A(G43gat), .B(G50gat), .Z(new_n208));
  INV_X1    g007(.A(KEYINPUT15), .ZN(new_n209));
  AOI22_X1  g008(.A1(new_n208), .A2(new_n209), .B1(G29gat), .B2(G36gat), .ZN(new_n210));
  INV_X1    g009(.A(KEYINPUT91), .ZN(new_n211));
  OAI21_X1  g010(.A(new_n211), .B1(G29gat), .B2(G36gat), .ZN(new_n212));
  OAI21_X1  g011(.A(new_n210), .B1(KEYINPUT14), .B2(new_n212), .ZN(new_n213));
  NOR2_X1   g012(.A1(new_n208), .A2(new_n209), .ZN(new_n214));
  INV_X1    g013(.A(G29gat), .ZN(new_n215));
  INV_X1    g014(.A(G36gat), .ZN(new_n216));
  NAND3_X1  g015(.A1(new_n215), .A2(new_n216), .A3(KEYINPUT91), .ZN(new_n217));
  AND3_X1   g016(.A1(new_n217), .A2(new_n212), .A3(KEYINPUT14), .ZN(new_n218));
  OR3_X1    g017(.A1(new_n213), .A2(new_n214), .A3(new_n218), .ZN(new_n219));
  OAI21_X1  g018(.A(new_n214), .B1(new_n213), .B2(new_n218), .ZN(new_n220));
  NAND2_X1  g019(.A1(new_n219), .A2(new_n220), .ZN(new_n221));
  INV_X1    g020(.A(KEYINPUT17), .ZN(new_n222));
  NAND2_X1  g021(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  XNOR2_X1  g022(.A(G15gat), .B(G22gat), .ZN(new_n224));
  INV_X1    g023(.A(KEYINPUT92), .ZN(new_n225));
  XNOR2_X1  g024(.A(new_n224), .B(new_n225), .ZN(new_n226));
  INV_X1    g025(.A(G1gat), .ZN(new_n227));
  NAND2_X1  g026(.A1(new_n226), .A2(new_n227), .ZN(new_n228));
  AND2_X1   g027(.A1(new_n227), .A2(KEYINPUT16), .ZN(new_n229));
  OAI21_X1  g028(.A(new_n228), .B1(new_n229), .B2(new_n226), .ZN(new_n230));
  INV_X1    g029(.A(G8gat), .ZN(new_n231));
  XNOR2_X1  g030(.A(new_n230), .B(new_n231), .ZN(new_n232));
  NAND3_X1  g031(.A1(new_n219), .A2(KEYINPUT17), .A3(new_n220), .ZN(new_n233));
  NAND3_X1  g032(.A1(new_n223), .A2(new_n232), .A3(new_n233), .ZN(new_n234));
  NAND2_X1  g033(.A1(G229gat), .A2(G233gat), .ZN(new_n235));
  XNOR2_X1  g034(.A(new_n230), .B(G8gat), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n236), .A2(new_n221), .ZN(new_n237));
  NAND3_X1  g036(.A1(new_n234), .A2(new_n235), .A3(new_n237), .ZN(new_n238));
  INV_X1    g037(.A(KEYINPUT18), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n238), .A2(new_n239), .ZN(new_n240));
  AOI21_X1  g039(.A(new_n207), .B1(new_n240), .B2(KEYINPUT93), .ZN(new_n241));
  NAND3_X1  g040(.A1(new_n232), .A2(new_n220), .A3(new_n219), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n242), .A2(new_n237), .ZN(new_n243));
  XOR2_X1   g042(.A(new_n235), .B(KEYINPUT13), .Z(new_n244));
  NAND2_X1  g043(.A1(new_n243), .A2(new_n244), .ZN(new_n245));
  NAND4_X1  g044(.A1(new_n234), .A2(KEYINPUT18), .A3(new_n235), .A4(new_n237), .ZN(new_n246));
  NAND3_X1  g045(.A1(new_n240), .A2(new_n245), .A3(new_n246), .ZN(new_n247));
  NAND2_X1  g046(.A1(new_n241), .A2(new_n247), .ZN(new_n248));
  AOI22_X1  g047(.A1(new_n238), .A2(new_n239), .B1(new_n243), .B2(new_n244), .ZN(new_n249));
  INV_X1    g048(.A(KEYINPUT93), .ZN(new_n250));
  AOI21_X1  g049(.A(new_n250), .B1(new_n238), .B2(new_n239), .ZN(new_n251));
  OAI211_X1 g050(.A(new_n249), .B(new_n246), .C1(new_n251), .C2(new_n207), .ZN(new_n252));
  NAND2_X1  g051(.A1(new_n248), .A2(new_n252), .ZN(new_n253));
  INV_X1    g052(.A(KEYINPUT94), .ZN(new_n254));
  NAND2_X1  g053(.A1(new_n253), .A2(new_n254), .ZN(new_n255));
  NAND3_X1  g054(.A1(new_n248), .A2(new_n252), .A3(KEYINPUT94), .ZN(new_n256));
  NAND2_X1  g055(.A1(new_n255), .A2(new_n256), .ZN(new_n257));
  XNOR2_X1  g056(.A(KEYINPUT79), .B(KEYINPUT31), .ZN(new_n258));
  INV_X1    g057(.A(new_n258), .ZN(new_n259));
  XNOR2_X1  g058(.A(G78gat), .B(G106gat), .ZN(new_n260));
  INV_X1    g059(.A(G50gat), .ZN(new_n261));
  XNOR2_X1  g060(.A(new_n260), .B(new_n261), .ZN(new_n262));
  INV_X1    g061(.A(new_n262), .ZN(new_n263));
  INV_X1    g062(.A(G22gat), .ZN(new_n264));
  INV_X1    g063(.A(G228gat), .ZN(new_n265));
  INV_X1    g064(.A(G233gat), .ZN(new_n266));
  INV_X1    g065(.A(KEYINPUT3), .ZN(new_n267));
  XOR2_X1   g066(.A(G211gat), .B(G218gat), .Z(new_n268));
  NAND2_X1  g067(.A1(new_n268), .A2(KEYINPUT70), .ZN(new_n269));
  XNOR2_X1  g068(.A(G197gat), .B(G204gat), .ZN(new_n270));
  INV_X1    g069(.A(KEYINPUT22), .ZN(new_n271));
  INV_X1    g070(.A(G211gat), .ZN(new_n272));
  INV_X1    g071(.A(G218gat), .ZN(new_n273));
  OAI21_X1  g072(.A(new_n271), .B1(new_n272), .B2(new_n273), .ZN(new_n274));
  NAND2_X1  g073(.A1(new_n270), .A2(new_n274), .ZN(new_n275));
  XNOR2_X1  g074(.A(new_n269), .B(new_n275), .ZN(new_n276));
  OAI21_X1  g075(.A(new_n267), .B1(new_n276), .B2(KEYINPUT29), .ZN(new_n277));
  INV_X1    g076(.A(KEYINPUT2), .ZN(new_n278));
  INV_X1    g077(.A(G155gat), .ZN(new_n279));
  INV_X1    g078(.A(G162gat), .ZN(new_n280));
  NAND3_X1  g079(.A1(new_n278), .A2(new_n279), .A3(new_n280), .ZN(new_n281));
  NAND2_X1  g080(.A1(G155gat), .A2(G162gat), .ZN(new_n282));
  NAND2_X1  g081(.A1(new_n281), .A2(new_n282), .ZN(new_n283));
  INV_X1    g082(.A(G141gat), .ZN(new_n284));
  NAND2_X1  g083(.A1(new_n284), .A2(G148gat), .ZN(new_n285));
  INV_X1    g084(.A(G148gat), .ZN(new_n286));
  NAND2_X1  g085(.A1(new_n286), .A2(G141gat), .ZN(new_n287));
  NAND3_X1  g086(.A1(new_n285), .A2(new_n287), .A3(KEYINPUT73), .ZN(new_n288));
  OAI211_X1 g087(.A(new_n283), .B(new_n288), .C1(KEYINPUT73), .C2(new_n285), .ZN(new_n289));
  NOR2_X1   g088(.A1(new_n286), .A2(G141gat), .ZN(new_n290));
  NOR2_X1   g089(.A1(new_n284), .A2(G148gat), .ZN(new_n291));
  OAI21_X1  g090(.A(new_n278), .B1(new_n290), .B2(new_n291), .ZN(new_n292));
  XOR2_X1   g091(.A(G155gat), .B(G162gat), .Z(new_n293));
  NAND2_X1  g092(.A1(new_n292), .A2(new_n293), .ZN(new_n294));
  NAND2_X1  g093(.A1(new_n289), .A2(new_n294), .ZN(new_n295));
  AOI211_X1 g094(.A(new_n265), .B(new_n266), .C1(new_n277), .C2(new_n295), .ZN(new_n296));
  INV_X1    g095(.A(KEYINPUT74), .ZN(new_n297));
  OAI21_X1  g096(.A(new_n297), .B1(new_n295), .B2(KEYINPUT3), .ZN(new_n298));
  INV_X1    g097(.A(KEYINPUT73), .ZN(new_n299));
  AOI22_X1  g098(.A1(new_n281), .A2(new_n282), .B1(new_n290), .B2(new_n299), .ZN(new_n300));
  AOI22_X1  g099(.A1(new_n300), .A2(new_n288), .B1(new_n292), .B2(new_n293), .ZN(new_n301));
  NAND3_X1  g100(.A1(new_n301), .A2(KEYINPUT74), .A3(new_n267), .ZN(new_n302));
  AOI21_X1  g101(.A(KEYINPUT29), .B1(new_n298), .B2(new_n302), .ZN(new_n303));
  AND2_X1   g102(.A1(new_n303), .A2(KEYINPUT80), .ZN(new_n304));
  OAI21_X1  g103(.A(new_n276), .B1(new_n303), .B2(KEYINPUT80), .ZN(new_n305));
  OAI21_X1  g104(.A(new_n296), .B1(new_n304), .B2(new_n305), .ZN(new_n306));
  INV_X1    g105(.A(new_n275), .ZN(new_n307));
  AND2_X1   g106(.A1(new_n307), .A2(new_n268), .ZN(new_n308));
  INV_X1    g107(.A(KEYINPUT29), .ZN(new_n309));
  OAI21_X1  g108(.A(new_n309), .B1(new_n307), .B2(new_n268), .ZN(new_n310));
  OAI21_X1  g109(.A(new_n267), .B1(new_n308), .B2(new_n310), .ZN(new_n311));
  NAND2_X1  g110(.A1(new_n311), .A2(new_n295), .ZN(new_n312));
  INV_X1    g111(.A(new_n276), .ZN(new_n313));
  OAI21_X1  g112(.A(new_n312), .B1(new_n303), .B2(new_n313), .ZN(new_n314));
  OAI21_X1  g113(.A(new_n314), .B1(new_n265), .B2(new_n266), .ZN(new_n315));
  AOI21_X1  g114(.A(new_n264), .B1(new_n306), .B2(new_n315), .ZN(new_n316));
  INV_X1    g115(.A(new_n316), .ZN(new_n317));
  NAND3_X1  g116(.A1(new_n306), .A2(new_n264), .A3(new_n315), .ZN(new_n318));
  AOI21_X1  g117(.A(new_n263), .B1(new_n317), .B2(new_n318), .ZN(new_n319));
  INV_X1    g118(.A(new_n318), .ZN(new_n320));
  NOR3_X1   g119(.A1(new_n320), .A2(new_n262), .A3(new_n316), .ZN(new_n321));
  OAI21_X1  g120(.A(new_n259), .B1(new_n319), .B2(new_n321), .ZN(new_n322));
  OAI21_X1  g121(.A(new_n262), .B1(new_n320), .B2(new_n316), .ZN(new_n323));
  NAND3_X1  g122(.A1(new_n317), .A2(new_n263), .A3(new_n318), .ZN(new_n324));
  NAND3_X1  g123(.A1(new_n323), .A2(new_n324), .A3(new_n258), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n322), .A2(new_n325), .ZN(new_n326));
  AND2_X1   g125(.A1(G227gat), .A2(G233gat), .ZN(new_n327));
  INV_X1    g126(.A(KEYINPUT69), .ZN(new_n328));
  OAI21_X1  g127(.A(KEYINPUT34), .B1(new_n327), .B2(new_n328), .ZN(new_n329));
  XNOR2_X1  g128(.A(G15gat), .B(G43gat), .ZN(new_n330));
  XNOR2_X1  g129(.A(new_n330), .B(KEYINPUT68), .ZN(new_n331));
  INV_X1    g130(.A(G71gat), .ZN(new_n332));
  XNOR2_X1  g131(.A(new_n331), .B(new_n332), .ZN(new_n333));
  XNOR2_X1  g132(.A(new_n333), .B(G99gat), .ZN(new_n334));
  INV_X1    g133(.A(G183gat), .ZN(new_n335));
  NOR2_X1   g134(.A1(new_n335), .A2(KEYINPUT24), .ZN(new_n336));
  NAND2_X1  g135(.A1(G183gat), .A2(G190gat), .ZN(new_n337));
  AOI22_X1  g136(.A1(new_n336), .A2(G190gat), .B1(KEYINPUT24), .B2(new_n337), .ZN(new_n338));
  NOR2_X1   g137(.A1(G183gat), .A2(G190gat), .ZN(new_n339));
  OAI21_X1  g138(.A(KEYINPUT65), .B1(new_n338), .B2(new_n339), .ZN(new_n340));
  NOR2_X1   g139(.A1(G169gat), .A2(G176gat), .ZN(new_n341));
  NAND2_X1  g140(.A1(new_n341), .A2(KEYINPUT23), .ZN(new_n342));
  INV_X1    g141(.A(KEYINPUT23), .ZN(new_n343));
  AOI21_X1  g142(.A(new_n343), .B1(G169gat), .B2(G176gat), .ZN(new_n344));
  OAI211_X1 g143(.A(KEYINPUT25), .B(new_n342), .C1(new_n344), .C2(new_n341), .ZN(new_n345));
  INV_X1    g144(.A(new_n345), .ZN(new_n346));
  NAND2_X1  g145(.A1(new_n337), .A2(KEYINPUT24), .ZN(new_n347));
  INV_X1    g146(.A(KEYINPUT24), .ZN(new_n348));
  NAND3_X1  g147(.A1(new_n348), .A2(G183gat), .A3(G190gat), .ZN(new_n349));
  NAND2_X1  g148(.A1(new_n347), .A2(new_n349), .ZN(new_n350));
  INV_X1    g149(.A(KEYINPUT65), .ZN(new_n351));
  INV_X1    g150(.A(new_n339), .ZN(new_n352));
  NAND3_X1  g151(.A1(new_n350), .A2(new_n351), .A3(new_n352), .ZN(new_n353));
  NAND3_X1  g152(.A1(new_n340), .A2(new_n346), .A3(new_n353), .ZN(new_n354));
  INV_X1    g153(.A(KEYINPUT25), .ZN(new_n355));
  INV_X1    g154(.A(KEYINPUT64), .ZN(new_n356));
  NAND2_X1  g155(.A1(new_n339), .A2(new_n356), .ZN(new_n357));
  OAI21_X1  g156(.A(KEYINPUT64), .B1(G183gat), .B2(G190gat), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n357), .A2(new_n358), .ZN(new_n359));
  NOR2_X1   g158(.A1(new_n338), .A2(new_n359), .ZN(new_n360));
  OAI21_X1  g159(.A(new_n342), .B1(new_n344), .B2(new_n341), .ZN(new_n361));
  OAI21_X1  g160(.A(new_n355), .B1(new_n360), .B2(new_n361), .ZN(new_n362));
  NAND2_X1  g161(.A1(new_n335), .A2(KEYINPUT27), .ZN(new_n363));
  INV_X1    g162(.A(KEYINPUT27), .ZN(new_n364));
  NAND2_X1  g163(.A1(new_n364), .A2(G183gat), .ZN(new_n365));
  INV_X1    g164(.A(G190gat), .ZN(new_n366));
  NAND3_X1  g165(.A1(new_n363), .A2(new_n365), .A3(new_n366), .ZN(new_n367));
  NAND3_X1  g166(.A1(new_n367), .A2(KEYINPUT66), .A3(KEYINPUT28), .ZN(new_n368));
  AOI21_X1  g167(.A(KEYINPUT28), .B1(new_n367), .B2(KEYINPUT66), .ZN(new_n369));
  INV_X1    g168(.A(KEYINPUT26), .ZN(new_n370));
  INV_X1    g169(.A(G169gat), .ZN(new_n371));
  INV_X1    g170(.A(G176gat), .ZN(new_n372));
  NAND3_X1  g171(.A1(new_n370), .A2(new_n371), .A3(new_n372), .ZN(new_n373));
  NAND2_X1  g172(.A1(G169gat), .A2(G176gat), .ZN(new_n374));
  OAI21_X1  g173(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n375));
  NAND3_X1  g174(.A1(new_n373), .A2(new_n374), .A3(new_n375), .ZN(new_n376));
  NAND2_X1  g175(.A1(new_n376), .A2(new_n337), .ZN(new_n377));
  NOR2_X1   g176(.A1(new_n369), .A2(new_n377), .ZN(new_n378));
  AOI22_X1  g177(.A1(new_n354), .A2(new_n362), .B1(new_n368), .B2(new_n378), .ZN(new_n379));
  INV_X1    g178(.A(KEYINPUT1), .ZN(new_n380));
  AND2_X1   g179(.A1(G113gat), .A2(G120gat), .ZN(new_n381));
  NOR2_X1   g180(.A1(G113gat), .A2(G120gat), .ZN(new_n382));
  NOR2_X1   g181(.A1(new_n381), .A2(new_n382), .ZN(new_n383));
  AND2_X1   g182(.A1(G127gat), .A2(G134gat), .ZN(new_n384));
  NOR2_X1   g183(.A1(G127gat), .A2(G134gat), .ZN(new_n385));
  NOR2_X1   g184(.A1(new_n384), .A2(new_n385), .ZN(new_n386));
  INV_X1    g185(.A(KEYINPUT67), .ZN(new_n387));
  OAI211_X1 g186(.A(new_n380), .B(new_n383), .C1(new_n386), .C2(new_n387), .ZN(new_n388));
  INV_X1    g187(.A(G113gat), .ZN(new_n389));
  INV_X1    g188(.A(G120gat), .ZN(new_n390));
  NAND2_X1  g189(.A1(new_n389), .A2(new_n390), .ZN(new_n391));
  NAND2_X1  g190(.A1(G113gat), .A2(G120gat), .ZN(new_n392));
  NAND3_X1  g191(.A1(new_n391), .A2(new_n380), .A3(new_n392), .ZN(new_n393));
  NAND3_X1  g192(.A1(new_n391), .A2(new_n387), .A3(new_n392), .ZN(new_n394));
  XNOR2_X1  g193(.A(G127gat), .B(G134gat), .ZN(new_n395));
  NAND3_X1  g194(.A1(new_n393), .A2(new_n394), .A3(new_n395), .ZN(new_n396));
  AND2_X1   g195(.A1(new_n388), .A2(new_n396), .ZN(new_n397));
  NAND2_X1  g196(.A1(new_n379), .A2(new_n397), .ZN(new_n398));
  NAND2_X1  g197(.A1(new_n367), .A2(KEYINPUT66), .ZN(new_n399));
  INV_X1    g198(.A(KEYINPUT28), .ZN(new_n400));
  NAND2_X1  g199(.A1(new_n399), .A2(new_n400), .ZN(new_n401));
  NAND4_X1  g200(.A1(new_n401), .A2(new_n337), .A3(new_n368), .A4(new_n376), .ZN(new_n402));
  AOI21_X1  g201(.A(new_n351), .B1(new_n350), .B2(new_n352), .ZN(new_n403));
  AOI211_X1 g202(.A(KEYINPUT65), .B(new_n339), .C1(new_n347), .C2(new_n349), .ZN(new_n404));
  NOR3_X1   g203(.A1(new_n403), .A2(new_n404), .A3(new_n345), .ZN(new_n405));
  INV_X1    g204(.A(new_n361), .ZN(new_n406));
  NAND3_X1  g205(.A1(new_n350), .A2(new_n358), .A3(new_n357), .ZN(new_n407));
  AOI21_X1  g206(.A(KEYINPUT25), .B1(new_n406), .B2(new_n407), .ZN(new_n408));
  OAI21_X1  g207(.A(new_n402), .B1(new_n405), .B2(new_n408), .ZN(new_n409));
  NAND2_X1  g208(.A1(new_n388), .A2(new_n396), .ZN(new_n410));
  NAND2_X1  g209(.A1(new_n409), .A2(new_n410), .ZN(new_n411));
  NAND3_X1  g210(.A1(new_n398), .A2(new_n411), .A3(new_n327), .ZN(new_n412));
  INV_X1    g211(.A(KEYINPUT33), .ZN(new_n413));
  AOI21_X1  g212(.A(new_n334), .B1(new_n412), .B2(new_n413), .ZN(new_n414));
  NAND2_X1  g213(.A1(new_n412), .A2(KEYINPUT32), .ZN(new_n415));
  NAND2_X1  g214(.A1(new_n414), .A2(new_n415), .ZN(new_n416));
  AND2_X1   g215(.A1(new_n398), .A2(new_n411), .ZN(new_n417));
  NOR2_X1   g216(.A1(new_n417), .A2(new_n327), .ZN(new_n418));
  INV_X1    g217(.A(new_n418), .ZN(new_n419));
  OAI211_X1 g218(.A(KEYINPUT32), .B(new_n412), .C1(new_n334), .C2(new_n413), .ZN(new_n420));
  NAND3_X1  g219(.A1(new_n416), .A2(new_n419), .A3(new_n420), .ZN(new_n421));
  INV_X1    g220(.A(new_n421), .ZN(new_n422));
  AOI21_X1  g221(.A(new_n419), .B1(new_n416), .B2(new_n420), .ZN(new_n423));
  OAI21_X1  g222(.A(new_n329), .B1(new_n422), .B2(new_n423), .ZN(new_n424));
  INV_X1    g223(.A(new_n423), .ZN(new_n425));
  INV_X1    g224(.A(new_n329), .ZN(new_n426));
  NAND3_X1  g225(.A1(new_n425), .A2(new_n426), .A3(new_n421), .ZN(new_n427));
  NAND2_X1  g226(.A1(new_n424), .A2(new_n427), .ZN(new_n428));
  NOR2_X1   g227(.A1(new_n326), .A2(new_n428), .ZN(new_n429));
  NAND2_X1  g228(.A1(G226gat), .A2(G233gat), .ZN(new_n430));
  INV_X1    g229(.A(new_n430), .ZN(new_n431));
  AOI21_X1  g230(.A(new_n431), .B1(new_n409), .B2(new_n309), .ZN(new_n432));
  NOR2_X1   g231(.A1(new_n379), .A2(new_n430), .ZN(new_n433));
  OAI21_X1  g232(.A(new_n276), .B1(new_n432), .B2(new_n433), .ZN(new_n434));
  OAI21_X1  g233(.A(new_n430), .B1(new_n379), .B2(KEYINPUT29), .ZN(new_n435));
  NAND2_X1  g234(.A1(new_n409), .A2(new_n431), .ZN(new_n436));
  NAND3_X1  g235(.A1(new_n435), .A2(new_n313), .A3(new_n436), .ZN(new_n437));
  XNOR2_X1  g236(.A(G8gat), .B(G36gat), .ZN(new_n438));
  XNOR2_X1  g237(.A(new_n438), .B(KEYINPUT71), .ZN(new_n439));
  XNOR2_X1  g238(.A(G64gat), .B(G92gat), .ZN(new_n440));
  XNOR2_X1  g239(.A(new_n439), .B(new_n440), .ZN(new_n441));
  NAND3_X1  g240(.A1(new_n434), .A2(new_n437), .A3(new_n441), .ZN(new_n442));
  INV_X1    g241(.A(KEYINPUT30), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  NAND4_X1  g243(.A1(new_n434), .A2(new_n437), .A3(KEYINPUT30), .A4(new_n441), .ZN(new_n445));
  INV_X1    g244(.A(new_n441), .ZN(new_n446));
  NOR3_X1   g245(.A1(new_n432), .A2(new_n433), .A3(new_n276), .ZN(new_n447));
  AOI21_X1  g246(.A(new_n313), .B1(new_n435), .B2(new_n436), .ZN(new_n448));
  OAI21_X1  g247(.A(new_n446), .B1(new_n447), .B2(new_n448), .ZN(new_n449));
  NAND4_X1  g248(.A1(new_n444), .A2(KEYINPUT72), .A3(new_n445), .A4(new_n449), .ZN(new_n450));
  INV_X1    g249(.A(KEYINPUT81), .ZN(new_n451));
  OR2_X1    g250(.A1(new_n445), .A2(KEYINPUT72), .ZN(new_n452));
  NAND3_X1  g251(.A1(new_n450), .A2(new_n451), .A3(new_n452), .ZN(new_n453));
  INV_X1    g252(.A(new_n453), .ZN(new_n454));
  AOI21_X1  g253(.A(new_n451), .B1(new_n450), .B2(new_n452), .ZN(new_n455));
  NOR2_X1   g254(.A1(new_n454), .A2(new_n455), .ZN(new_n456));
  INV_X1    g255(.A(new_n456), .ZN(new_n457));
  XNOR2_X1  g256(.A(G1gat), .B(G29gat), .ZN(new_n458));
  XNOR2_X1  g257(.A(new_n458), .B(KEYINPUT0), .ZN(new_n459));
  XNOR2_X1  g258(.A(G57gat), .B(G85gat), .ZN(new_n460));
  XOR2_X1   g259(.A(new_n459), .B(new_n460), .Z(new_n461));
  INV_X1    g260(.A(new_n461), .ZN(new_n462));
  NAND2_X1  g261(.A1(G225gat), .A2(G233gat), .ZN(new_n463));
  INV_X1    g262(.A(new_n463), .ZN(new_n464));
  NAND2_X1  g263(.A1(new_n298), .A2(new_n302), .ZN(new_n465));
  AOI21_X1  g264(.A(new_n410), .B1(new_n295), .B2(KEYINPUT3), .ZN(new_n466));
  AOI21_X1  g265(.A(new_n464), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  AND3_X1   g266(.A1(new_n301), .A2(new_n410), .A3(KEYINPUT75), .ZN(new_n468));
  AOI21_X1  g267(.A(KEYINPUT75), .B1(new_n301), .B2(new_n410), .ZN(new_n469));
  NOR2_X1   g268(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  INV_X1    g269(.A(KEYINPUT4), .ZN(new_n471));
  NAND2_X1  g270(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  NAND3_X1  g271(.A1(new_n301), .A2(new_n410), .A3(KEYINPUT4), .ZN(new_n473));
  NAND3_X1  g272(.A1(new_n467), .A2(new_n472), .A3(new_n473), .ZN(new_n474));
  INV_X1    g273(.A(new_n474), .ZN(new_n475));
  INV_X1    g274(.A(KEYINPUT5), .ZN(new_n476));
  INV_X1    g275(.A(KEYINPUT75), .ZN(new_n477));
  OAI21_X1  g276(.A(new_n477), .B1(new_n397), .B2(new_n295), .ZN(new_n478));
  NAND3_X1  g277(.A1(new_n301), .A2(new_n410), .A3(KEYINPUT75), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n397), .A2(new_n295), .ZN(new_n480));
  NAND3_X1  g279(.A1(new_n478), .A2(new_n479), .A3(new_n480), .ZN(new_n481));
  AOI21_X1  g280(.A(new_n476), .B1(new_n481), .B2(new_n464), .ZN(new_n482));
  INV_X1    g281(.A(KEYINPUT76), .ZN(new_n483));
  OR2_X1    g282(.A1(new_n482), .A2(new_n483), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n482), .A2(new_n483), .ZN(new_n485));
  AOI21_X1  g284(.A(new_n475), .B1(new_n484), .B2(new_n485), .ZN(new_n486));
  NAND2_X1  g285(.A1(new_n467), .A2(new_n476), .ZN(new_n487));
  OAI21_X1  g286(.A(KEYINPUT4), .B1(new_n468), .B2(new_n469), .ZN(new_n488));
  OAI21_X1  g287(.A(new_n471), .B1(new_n397), .B2(new_n295), .ZN(new_n489));
  NAND2_X1  g288(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  NOR2_X1   g289(.A1(new_n487), .A2(new_n490), .ZN(new_n491));
  OAI21_X1  g290(.A(new_n462), .B1(new_n486), .B2(new_n491), .ZN(new_n492));
  XOR2_X1   g291(.A(KEYINPUT78), .B(KEYINPUT6), .Z(new_n493));
  NOR3_X1   g292(.A1(new_n492), .A2(KEYINPUT86), .A3(new_n493), .ZN(new_n494));
  INV_X1    g293(.A(KEYINPUT86), .ZN(new_n495));
  AND2_X1   g294(.A1(new_n482), .A2(new_n483), .ZN(new_n496));
  NOR2_X1   g295(.A1(new_n482), .A2(new_n483), .ZN(new_n497));
  OAI21_X1  g296(.A(new_n474), .B1(new_n496), .B2(new_n497), .ZN(new_n498));
  INV_X1    g297(.A(new_n491), .ZN(new_n499));
  AOI21_X1  g298(.A(new_n461), .B1(new_n498), .B2(new_n499), .ZN(new_n500));
  INV_X1    g299(.A(new_n493), .ZN(new_n501));
  AOI21_X1  g300(.A(new_n495), .B1(new_n500), .B2(new_n501), .ZN(new_n502));
  NOR2_X1   g301(.A1(new_n494), .A2(new_n502), .ZN(new_n503));
  NAND3_X1  g302(.A1(new_n498), .A2(new_n461), .A3(new_n499), .ZN(new_n504));
  NAND2_X1  g303(.A1(new_n504), .A2(KEYINPUT77), .ZN(new_n505));
  INV_X1    g304(.A(KEYINPUT77), .ZN(new_n506));
  NAND4_X1  g305(.A1(new_n498), .A2(new_n506), .A3(new_n461), .A4(new_n499), .ZN(new_n507));
  NAND2_X1  g306(.A1(new_n505), .A2(new_n507), .ZN(new_n508));
  NAND3_X1  g307(.A1(new_n508), .A2(new_n492), .A3(new_n493), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n503), .A2(new_n509), .ZN(new_n510));
  XOR2_X1   g309(.A(KEYINPUT88), .B(KEYINPUT35), .Z(new_n511));
  NAND4_X1  g310(.A1(new_n429), .A2(new_n457), .A3(new_n510), .A4(new_n511), .ZN(new_n512));
  NAND3_X1  g311(.A1(new_n449), .A2(KEYINPUT72), .A3(new_n445), .ZN(new_n513));
  AND2_X1   g312(.A1(new_n442), .A2(new_n443), .ZN(new_n514));
  OAI21_X1  g313(.A(new_n452), .B1(new_n513), .B2(new_n514), .ZN(new_n515));
  AOI211_X1 g314(.A(new_n500), .B(new_n501), .C1(new_n505), .C2(new_n507), .ZN(new_n516));
  NOR2_X1   g315(.A1(new_n492), .A2(new_n493), .ZN(new_n517));
  OAI21_X1  g316(.A(new_n515), .B1(new_n516), .B2(new_n517), .ZN(new_n518));
  AND2_X1   g317(.A1(new_n322), .A2(new_n325), .ZN(new_n519));
  INV_X1    g318(.A(new_n428), .ZN(new_n520));
  NAND3_X1  g319(.A1(new_n519), .A2(new_n520), .A3(KEYINPUT89), .ZN(new_n521));
  INV_X1    g320(.A(KEYINPUT89), .ZN(new_n522));
  OAI21_X1  g321(.A(new_n522), .B1(new_n326), .B2(new_n428), .ZN(new_n523));
  AOI21_X1  g322(.A(new_n518), .B1(new_n521), .B2(new_n523), .ZN(new_n524));
  INV_X1    g323(.A(KEYINPUT35), .ZN(new_n525));
  OAI21_X1  g324(.A(new_n512), .B1(new_n524), .B2(new_n525), .ZN(new_n526));
  INV_X1    g325(.A(KEYINPUT40), .ZN(new_n527));
  AOI21_X1  g326(.A(KEYINPUT74), .B1(new_n301), .B2(new_n267), .ZN(new_n528));
  AND4_X1   g327(.A1(KEYINPUT74), .A2(new_n289), .A3(new_n267), .A4(new_n294), .ZN(new_n529));
  OAI21_X1  g328(.A(new_n466), .B1(new_n528), .B2(new_n529), .ZN(new_n530));
  NAND3_X1  g329(.A1(new_n488), .A2(new_n530), .A3(new_n489), .ZN(new_n531));
  AND3_X1   g330(.A1(new_n531), .A2(KEYINPUT82), .A3(new_n464), .ZN(new_n532));
  AOI21_X1  g331(.A(KEYINPUT82), .B1(new_n531), .B2(new_n464), .ZN(new_n533));
  NOR2_X1   g332(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  NAND3_X1  g333(.A1(new_n470), .A2(new_n463), .A3(new_n480), .ZN(new_n535));
  AND2_X1   g334(.A1(new_n535), .A2(KEYINPUT84), .ZN(new_n536));
  NOR2_X1   g335(.A1(new_n535), .A2(KEYINPUT84), .ZN(new_n537));
  INV_X1    g336(.A(KEYINPUT39), .ZN(new_n538));
  NOR3_X1   g337(.A1(new_n536), .A2(new_n537), .A3(new_n538), .ZN(new_n539));
  AOI21_X1  g338(.A(new_n527), .B1(new_n534), .B2(new_n539), .ZN(new_n540));
  OAI21_X1  g339(.A(new_n538), .B1(new_n532), .B2(new_n533), .ZN(new_n541));
  INV_X1    g340(.A(KEYINPUT83), .ZN(new_n542));
  AND3_X1   g341(.A1(new_n541), .A2(new_n542), .A3(new_n461), .ZN(new_n543));
  AOI21_X1  g342(.A(new_n542), .B1(new_n541), .B2(new_n461), .ZN(new_n544));
  OAI21_X1  g343(.A(new_n540), .B1(new_n543), .B2(new_n544), .ZN(new_n545));
  NAND2_X1  g344(.A1(new_n515), .A2(KEYINPUT81), .ZN(new_n546));
  NAND4_X1  g345(.A1(new_n545), .A2(new_n492), .A3(new_n546), .A4(new_n453), .ZN(new_n547));
  NAND2_X1  g346(.A1(new_n531), .A2(new_n464), .ZN(new_n548));
  INV_X1    g347(.A(KEYINPUT82), .ZN(new_n549));
  NAND2_X1  g348(.A1(new_n548), .A2(new_n549), .ZN(new_n550));
  NAND3_X1  g349(.A1(new_n531), .A2(KEYINPUT82), .A3(new_n464), .ZN(new_n551));
  AOI21_X1  g350(.A(KEYINPUT39), .B1(new_n550), .B2(new_n551), .ZN(new_n552));
  OAI21_X1  g351(.A(KEYINPUT83), .B1(new_n552), .B2(new_n462), .ZN(new_n553));
  NAND3_X1  g352(.A1(new_n541), .A2(new_n542), .A3(new_n461), .ZN(new_n554));
  NAND2_X1  g353(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  NAND2_X1  g354(.A1(new_n534), .A2(new_n539), .ZN(new_n556));
  AOI21_X1  g355(.A(KEYINPUT40), .B1(new_n555), .B2(new_n556), .ZN(new_n557));
  OAI21_X1  g356(.A(KEYINPUT85), .B1(new_n547), .B2(new_n557), .ZN(new_n558));
  OAI21_X1  g357(.A(new_n556), .B1(new_n543), .B2(new_n544), .ZN(new_n559));
  NAND2_X1  g358(.A1(new_n559), .A2(new_n527), .ZN(new_n560));
  AOI21_X1  g359(.A(new_n500), .B1(new_n555), .B2(new_n540), .ZN(new_n561));
  INV_X1    g360(.A(KEYINPUT85), .ZN(new_n562));
  NAND4_X1  g361(.A1(new_n456), .A2(new_n560), .A3(new_n561), .A4(new_n562), .ZN(new_n563));
  NAND2_X1  g362(.A1(new_n434), .A2(new_n437), .ZN(new_n564));
  OR2_X1    g363(.A1(new_n564), .A2(KEYINPUT37), .ZN(new_n565));
  INV_X1    g364(.A(KEYINPUT38), .ZN(new_n566));
  AOI21_X1  g365(.A(new_n441), .B1(new_n564), .B2(KEYINPUT37), .ZN(new_n567));
  NAND3_X1  g366(.A1(new_n565), .A2(new_n566), .A3(new_n567), .ZN(new_n568));
  NAND2_X1  g367(.A1(new_n568), .A2(new_n442), .ZN(new_n569));
  OR2_X1    g368(.A1(new_n567), .A2(KEYINPUT87), .ZN(new_n570));
  NAND2_X1  g369(.A1(new_n567), .A2(KEYINPUT87), .ZN(new_n571));
  NAND3_X1  g370(.A1(new_n570), .A2(new_n571), .A3(new_n565), .ZN(new_n572));
  AOI21_X1  g371(.A(new_n569), .B1(new_n572), .B2(KEYINPUT38), .ZN(new_n573));
  NAND3_X1  g372(.A1(new_n503), .A2(new_n573), .A3(new_n509), .ZN(new_n574));
  NAND4_X1  g373(.A1(new_n558), .A2(new_n563), .A3(new_n519), .A4(new_n574), .ZN(new_n575));
  INV_X1    g374(.A(KEYINPUT36), .ZN(new_n576));
  NAND2_X1  g375(.A1(new_n428), .A2(new_n576), .ZN(new_n577));
  NAND3_X1  g376(.A1(new_n424), .A2(new_n427), .A3(KEYINPUT36), .ZN(new_n578));
  AOI22_X1  g377(.A1(new_n518), .A2(new_n326), .B1(new_n577), .B2(new_n578), .ZN(new_n579));
  NAND2_X1  g378(.A1(new_n575), .A2(new_n579), .ZN(new_n580));
  AOI21_X1  g379(.A(new_n257), .B1(new_n526), .B2(new_n580), .ZN(new_n581));
  XNOR2_X1  g380(.A(G134gat), .B(G162gat), .ZN(new_n582));
  INV_X1    g381(.A(KEYINPUT41), .ZN(new_n583));
  INV_X1    g382(.A(G232gat), .ZN(new_n584));
  OAI21_X1  g383(.A(new_n583), .B1(new_n584), .B2(new_n266), .ZN(new_n585));
  XOR2_X1   g384(.A(new_n582), .B(new_n585), .Z(new_n586));
  INV_X1    g385(.A(new_n586), .ZN(new_n587));
  XNOR2_X1  g386(.A(KEYINPUT97), .B(KEYINPUT7), .ZN(new_n588));
  INV_X1    g387(.A(G85gat), .ZN(new_n589));
  INV_X1    g388(.A(G92gat), .ZN(new_n590));
  NOR2_X1   g389(.A1(new_n589), .A2(new_n590), .ZN(new_n591));
  OR2_X1    g390(.A1(new_n588), .A2(new_n591), .ZN(new_n592));
  NAND2_X1  g391(.A1(new_n588), .A2(new_n591), .ZN(new_n593));
  NAND2_X1  g392(.A1(G99gat), .A2(G106gat), .ZN(new_n594));
  AOI22_X1  g393(.A1(KEYINPUT8), .A2(new_n594), .B1(new_n589), .B2(new_n590), .ZN(new_n595));
  NAND3_X1  g394(.A1(new_n592), .A2(new_n593), .A3(new_n595), .ZN(new_n596));
  XOR2_X1   g395(.A(G99gat), .B(G106gat), .Z(new_n597));
  OR2_X1    g396(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  NAND2_X1  g397(.A1(new_n596), .A2(new_n597), .ZN(new_n599));
  AND2_X1   g398(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  AOI21_X1  g399(.A(new_n600), .B1(new_n221), .B2(new_n222), .ZN(new_n601));
  NAND2_X1  g400(.A1(new_n601), .A2(new_n233), .ZN(new_n602));
  NAND2_X1  g401(.A1(new_n602), .A2(KEYINPUT98), .ZN(new_n603));
  INV_X1    g402(.A(KEYINPUT98), .ZN(new_n604));
  NAND3_X1  g403(.A1(new_n601), .A2(new_n604), .A3(new_n233), .ZN(new_n605));
  NAND2_X1  g404(.A1(new_n603), .A2(new_n605), .ZN(new_n606));
  XNOR2_X1  g405(.A(G190gat), .B(G218gat), .ZN(new_n607));
  INV_X1    g406(.A(new_n607), .ZN(new_n608));
  AND2_X1   g407(.A1(new_n608), .A2(KEYINPUT99), .ZN(new_n609));
  XNOR2_X1  g408(.A(new_n609), .B(KEYINPUT100), .ZN(new_n610));
  INV_X1    g409(.A(new_n610), .ZN(new_n611));
  NAND3_X1  g410(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n612));
  OAI21_X1  g411(.A(new_n612), .B1(new_n608), .B2(KEYINPUT99), .ZN(new_n613));
  AOI21_X1  g412(.A(new_n613), .B1(new_n221), .B2(new_n600), .ZN(new_n614));
  AND3_X1   g413(.A1(new_n606), .A2(new_n611), .A3(new_n614), .ZN(new_n615));
  AOI21_X1  g414(.A(new_n611), .B1(new_n606), .B2(new_n614), .ZN(new_n616));
  OAI21_X1  g415(.A(new_n587), .B1(new_n615), .B2(new_n616), .ZN(new_n617));
  NAND2_X1  g416(.A1(new_n606), .A2(new_n614), .ZN(new_n618));
  NAND2_X1  g417(.A1(new_n618), .A2(new_n610), .ZN(new_n619));
  NAND3_X1  g418(.A1(new_n606), .A2(new_n611), .A3(new_n614), .ZN(new_n620));
  NAND3_X1  g419(.A1(new_n619), .A2(new_n586), .A3(new_n620), .ZN(new_n621));
  NAND2_X1  g420(.A1(new_n617), .A2(new_n621), .ZN(new_n622));
  INV_X1    g421(.A(new_n622), .ZN(new_n623));
  NAND2_X1  g422(.A1(G71gat), .A2(G78gat), .ZN(new_n624));
  NOR2_X1   g423(.A1(G71gat), .A2(G78gat), .ZN(new_n625));
  OAI21_X1  g424(.A(new_n624), .B1(new_n625), .B2(KEYINPUT95), .ZN(new_n626));
  XNOR2_X1  g425(.A(G57gat), .B(G64gat), .ZN(new_n627));
  INV_X1    g426(.A(KEYINPUT9), .ZN(new_n628));
  OAI21_X1  g427(.A(new_n626), .B1(new_n627), .B2(new_n628), .ZN(new_n629));
  AOI21_X1  g428(.A(new_n624), .B1(new_n627), .B2(KEYINPUT95), .ZN(new_n630));
  OR2_X1    g429(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  NAND2_X1  g430(.A1(new_n625), .A2(KEYINPUT9), .ZN(new_n632));
  AOI22_X1  g431(.A1(new_n627), .A2(KEYINPUT96), .B1(new_n632), .B2(new_n624), .ZN(new_n633));
  OAI21_X1  g432(.A(new_n633), .B1(KEYINPUT96), .B2(new_n627), .ZN(new_n634));
  NAND2_X1  g433(.A1(new_n631), .A2(new_n634), .ZN(new_n635));
  INV_X1    g434(.A(KEYINPUT21), .ZN(new_n636));
  NAND2_X1  g435(.A1(new_n635), .A2(new_n636), .ZN(new_n637));
  NAND2_X1  g436(.A1(G231gat), .A2(G233gat), .ZN(new_n638));
  XNOR2_X1  g437(.A(new_n637), .B(new_n638), .ZN(new_n639));
  XNOR2_X1  g438(.A(new_n639), .B(G127gat), .ZN(new_n640));
  OAI21_X1  g439(.A(new_n232), .B1(new_n636), .B2(new_n635), .ZN(new_n641));
  XNOR2_X1  g440(.A(new_n640), .B(new_n641), .ZN(new_n642));
  XNOR2_X1  g441(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n643));
  XNOR2_X1  g442(.A(new_n643), .B(new_n279), .ZN(new_n644));
  XOR2_X1   g443(.A(G183gat), .B(G211gat), .Z(new_n645));
  XNOR2_X1  g444(.A(new_n644), .B(new_n645), .ZN(new_n646));
  INV_X1    g445(.A(new_n646), .ZN(new_n647));
  OR2_X1    g446(.A1(new_n642), .A2(new_n647), .ZN(new_n648));
  NAND2_X1  g447(.A1(new_n642), .A2(new_n647), .ZN(new_n649));
  NAND2_X1  g448(.A1(new_n648), .A2(new_n649), .ZN(new_n650));
  NAND4_X1  g449(.A1(new_n598), .A2(new_n631), .A3(new_n634), .A4(new_n599), .ZN(new_n651));
  INV_X1    g450(.A(new_n651), .ZN(new_n652));
  INV_X1    g451(.A(KEYINPUT101), .ZN(new_n653));
  NAND3_X1  g452(.A1(new_n652), .A2(new_n653), .A3(KEYINPUT10), .ZN(new_n654));
  NAND2_X1  g453(.A1(new_n598), .A2(new_n599), .ZN(new_n655));
  NAND2_X1  g454(.A1(new_n655), .A2(new_n635), .ZN(new_n656));
  INV_X1    g455(.A(KEYINPUT10), .ZN(new_n657));
  NAND3_X1  g456(.A1(new_n656), .A2(new_n657), .A3(new_n651), .ZN(new_n658));
  OAI21_X1  g457(.A(KEYINPUT101), .B1(new_n651), .B2(new_n657), .ZN(new_n659));
  NAND3_X1  g458(.A1(new_n654), .A2(new_n658), .A3(new_n659), .ZN(new_n660));
  NAND2_X1  g459(.A1(G230gat), .A2(G233gat), .ZN(new_n661));
  XNOR2_X1  g460(.A(new_n661), .B(KEYINPUT102), .ZN(new_n662));
  INV_X1    g461(.A(new_n662), .ZN(new_n663));
  NAND2_X1  g462(.A1(new_n660), .A2(new_n663), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n656), .A2(new_n651), .ZN(new_n665));
  NAND2_X1  g464(.A1(new_n665), .A2(new_n662), .ZN(new_n666));
  NAND2_X1  g465(.A1(new_n664), .A2(new_n666), .ZN(new_n667));
  XNOR2_X1  g466(.A(G120gat), .B(G148gat), .ZN(new_n668));
  XNOR2_X1  g467(.A(G176gat), .B(G204gat), .ZN(new_n669));
  XOR2_X1   g468(.A(new_n668), .B(new_n669), .Z(new_n670));
  INV_X1    g469(.A(new_n670), .ZN(new_n671));
  NAND2_X1  g470(.A1(new_n667), .A2(new_n671), .ZN(new_n672));
  NAND3_X1  g471(.A1(new_n664), .A2(new_n666), .A3(new_n670), .ZN(new_n673));
  AND2_X1   g472(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  NAND3_X1  g473(.A1(new_n623), .A2(new_n650), .A3(new_n674), .ZN(new_n675));
  OR2_X1    g474(.A1(new_n675), .A2(KEYINPUT103), .ZN(new_n676));
  NAND2_X1  g475(.A1(new_n675), .A2(KEYINPUT103), .ZN(new_n677));
  NAND2_X1  g476(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  INV_X1    g477(.A(new_n678), .ZN(new_n679));
  NAND2_X1  g478(.A1(new_n581), .A2(new_n679), .ZN(new_n680));
  NOR2_X1   g479(.A1(new_n516), .A2(new_n517), .ZN(new_n681));
  INV_X1    g480(.A(new_n681), .ZN(new_n682));
  NOR2_X1   g481(.A1(new_n680), .A2(new_n682), .ZN(new_n683));
  XNOR2_X1  g482(.A(new_n683), .B(new_n227), .ZN(G1324gat));
  NAND3_X1  g483(.A1(new_n581), .A2(new_n456), .A3(new_n679), .ZN(new_n685));
  XNOR2_X1  g484(.A(KEYINPUT16), .B(G8gat), .ZN(new_n686));
  NOR2_X1   g485(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  NOR2_X1   g486(.A1(new_n687), .A2(KEYINPUT42), .ZN(new_n688));
  AOI21_X1  g487(.A(new_n688), .B1(G8gat), .B2(new_n685), .ZN(new_n689));
  NAND2_X1  g488(.A1(new_n687), .A2(KEYINPUT42), .ZN(new_n690));
  NAND2_X1  g489(.A1(new_n689), .A2(new_n690), .ZN(G1325gat));
  NAND2_X1  g490(.A1(new_n577), .A2(new_n578), .ZN(new_n692));
  OAI21_X1  g491(.A(G15gat), .B1(new_n680), .B2(new_n692), .ZN(new_n693));
  OR2_X1    g492(.A1(new_n428), .A2(G15gat), .ZN(new_n694));
  OAI21_X1  g493(.A(new_n693), .B1(new_n680), .B2(new_n694), .ZN(G1326gat));
  NOR2_X1   g494(.A1(new_n680), .A2(new_n519), .ZN(new_n696));
  XOR2_X1   g495(.A(KEYINPUT43), .B(G22gat), .Z(new_n697));
  XNOR2_X1  g496(.A(new_n696), .B(new_n697), .ZN(new_n698));
  XNOR2_X1  g497(.A(KEYINPUT104), .B(KEYINPUT105), .ZN(new_n699));
  XNOR2_X1  g498(.A(new_n698), .B(new_n699), .ZN(G1327gat));
  NAND2_X1  g499(.A1(new_n526), .A2(new_n580), .ZN(new_n701));
  INV_X1    g500(.A(new_n257), .ZN(new_n702));
  INV_X1    g501(.A(new_n674), .ZN(new_n703));
  NOR2_X1   g502(.A1(new_n650), .A2(new_n703), .ZN(new_n704));
  AND4_X1   g503(.A1(new_n701), .A2(new_n702), .A3(new_n622), .A4(new_n704), .ZN(new_n705));
  NAND3_X1  g504(.A1(new_n705), .A2(new_n215), .A3(new_n681), .ZN(new_n706));
  XNOR2_X1  g505(.A(new_n706), .B(KEYINPUT45), .ZN(new_n707));
  NAND2_X1  g506(.A1(new_n701), .A2(new_n622), .ZN(new_n708));
  NAND2_X1  g507(.A1(new_n708), .A2(KEYINPUT44), .ZN(new_n709));
  AND3_X1   g508(.A1(new_n575), .A2(KEYINPUT106), .A3(new_n579), .ZN(new_n710));
  AOI21_X1  g509(.A(KEYINPUT106), .B1(new_n575), .B2(new_n579), .ZN(new_n711));
  OAI21_X1  g510(.A(new_n526), .B1(new_n710), .B2(new_n711), .ZN(new_n712));
  INV_X1    g511(.A(KEYINPUT107), .ZN(new_n713));
  NOR2_X1   g512(.A1(new_n623), .A2(KEYINPUT44), .ZN(new_n714));
  AND3_X1   g513(.A1(new_n712), .A2(new_n713), .A3(new_n714), .ZN(new_n715));
  AOI21_X1  g514(.A(new_n713), .B1(new_n712), .B2(new_n714), .ZN(new_n716));
  OAI21_X1  g515(.A(new_n709), .B1(new_n715), .B2(new_n716), .ZN(new_n717));
  INV_X1    g516(.A(new_n717), .ZN(new_n718));
  INV_X1    g517(.A(new_n704), .ZN(new_n719));
  INV_X1    g518(.A(new_n253), .ZN(new_n720));
  NOR2_X1   g519(.A1(new_n719), .A2(new_n720), .ZN(new_n721));
  INV_X1    g520(.A(new_n721), .ZN(new_n722));
  NOR3_X1   g521(.A1(new_n718), .A2(new_n682), .A3(new_n722), .ZN(new_n723));
  OAI21_X1  g522(.A(new_n707), .B1(new_n723), .B2(new_n215), .ZN(G1328gat));
  NAND3_X1  g523(.A1(new_n705), .A2(new_n216), .A3(new_n456), .ZN(new_n725));
  XOR2_X1   g524(.A(new_n725), .B(KEYINPUT46), .Z(new_n726));
  NOR3_X1   g525(.A1(new_n718), .A2(new_n457), .A3(new_n722), .ZN(new_n727));
  OAI21_X1  g526(.A(new_n726), .B1(new_n727), .B2(new_n216), .ZN(new_n728));
  INV_X1    g527(.A(KEYINPUT108), .ZN(new_n729));
  NAND2_X1  g528(.A1(new_n728), .A2(new_n729), .ZN(new_n730));
  OAI211_X1 g529(.A(new_n726), .B(KEYINPUT108), .C1(new_n727), .C2(new_n216), .ZN(new_n731));
  NAND2_X1  g530(.A1(new_n730), .A2(new_n731), .ZN(G1329gat));
  INV_X1    g531(.A(new_n692), .ZN(new_n733));
  NAND3_X1  g532(.A1(new_n717), .A2(new_n733), .A3(new_n721), .ZN(new_n734));
  NAND2_X1  g533(.A1(new_n734), .A2(G43gat), .ZN(new_n735));
  INV_X1    g534(.A(G43gat), .ZN(new_n736));
  NAND3_X1  g535(.A1(new_n705), .A2(new_n736), .A3(new_n520), .ZN(new_n737));
  NAND3_X1  g536(.A1(new_n735), .A2(KEYINPUT47), .A3(new_n737), .ZN(new_n738));
  INV_X1    g537(.A(KEYINPUT110), .ZN(new_n739));
  AND3_X1   g538(.A1(new_n734), .A2(new_n739), .A3(G43gat), .ZN(new_n740));
  AOI21_X1  g539(.A(new_n739), .B1(new_n734), .B2(G43gat), .ZN(new_n741));
  INV_X1    g540(.A(new_n737), .ZN(new_n742));
  NOR3_X1   g541(.A1(new_n740), .A2(new_n741), .A3(new_n742), .ZN(new_n743));
  XNOR2_X1  g542(.A(KEYINPUT109), .B(KEYINPUT47), .ZN(new_n744));
  OAI21_X1  g543(.A(new_n738), .B1(new_n743), .B2(new_n744), .ZN(G1330gat));
  NAND2_X1  g544(.A1(new_n326), .A2(new_n261), .ZN(new_n746));
  XNOR2_X1  g545(.A(new_n746), .B(KEYINPUT111), .ZN(new_n747));
  NAND2_X1  g546(.A1(new_n705), .A2(new_n747), .ZN(new_n748));
  NOR3_X1   g547(.A1(new_n718), .A2(new_n519), .A3(new_n722), .ZN(new_n749));
  OAI21_X1  g548(.A(new_n748), .B1(new_n749), .B2(new_n261), .ZN(new_n750));
  INV_X1    g549(.A(KEYINPUT48), .ZN(new_n751));
  NAND2_X1  g550(.A1(new_n750), .A2(new_n751), .ZN(new_n752));
  OAI211_X1 g551(.A(KEYINPUT48), .B(new_n748), .C1(new_n749), .C2(new_n261), .ZN(new_n753));
  NAND2_X1  g552(.A1(new_n752), .A2(new_n753), .ZN(G1331gat));
  INV_X1    g553(.A(new_n650), .ZN(new_n755));
  NOR4_X1   g554(.A1(new_n755), .A2(new_n253), .A3(new_n622), .A4(new_n674), .ZN(new_n756));
  AND2_X1   g555(.A1(new_n712), .A2(new_n756), .ZN(new_n757));
  NAND2_X1  g556(.A1(new_n757), .A2(new_n681), .ZN(new_n758));
  XNOR2_X1  g557(.A(new_n758), .B(G57gat), .ZN(G1332gat));
  NAND2_X1  g558(.A1(new_n757), .A2(new_n456), .ZN(new_n760));
  OAI21_X1  g559(.A(new_n760), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n761));
  XOR2_X1   g560(.A(KEYINPUT49), .B(G64gat), .Z(new_n762));
  OAI21_X1  g561(.A(new_n761), .B1(new_n760), .B2(new_n762), .ZN(G1333gat));
  AOI21_X1  g562(.A(new_n332), .B1(new_n757), .B2(new_n733), .ZN(new_n764));
  NOR2_X1   g563(.A1(new_n428), .A2(G71gat), .ZN(new_n765));
  AOI21_X1  g564(.A(new_n764), .B1(new_n757), .B2(new_n765), .ZN(new_n766));
  XNOR2_X1  g565(.A(new_n766), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g566(.A1(new_n757), .A2(new_n326), .ZN(new_n768));
  XNOR2_X1  g567(.A(new_n768), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g568(.A1(new_n650), .A2(new_n253), .ZN(new_n770));
  NAND3_X1  g569(.A1(new_n712), .A2(new_n622), .A3(new_n770), .ZN(new_n771));
  INV_X1    g570(.A(KEYINPUT51), .ZN(new_n772));
  XNOR2_X1  g571(.A(new_n771), .B(new_n772), .ZN(new_n773));
  NAND4_X1  g572(.A1(new_n773), .A2(new_n589), .A3(new_n681), .A4(new_n703), .ZN(new_n774));
  NAND2_X1  g573(.A1(new_n770), .A2(new_n703), .ZN(new_n775));
  XNOR2_X1  g574(.A(new_n775), .B(KEYINPUT112), .ZN(new_n776));
  NOR3_X1   g575(.A1(new_n718), .A2(new_n682), .A3(new_n776), .ZN(new_n777));
  OAI21_X1  g576(.A(new_n774), .B1(new_n777), .B2(new_n589), .ZN(G1336gat));
  NAND4_X1  g577(.A1(new_n773), .A2(new_n590), .A3(new_n456), .A4(new_n703), .ZN(new_n779));
  NOR3_X1   g578(.A1(new_n718), .A2(new_n457), .A3(new_n776), .ZN(new_n780));
  OAI21_X1  g579(.A(new_n779), .B1(new_n780), .B2(new_n590), .ZN(new_n781));
  NAND2_X1  g580(.A1(new_n781), .A2(KEYINPUT52), .ZN(new_n782));
  INV_X1    g581(.A(KEYINPUT52), .ZN(new_n783));
  OAI211_X1 g582(.A(new_n783), .B(new_n779), .C1(new_n780), .C2(new_n590), .ZN(new_n784));
  NAND2_X1  g583(.A1(new_n782), .A2(new_n784), .ZN(G1337gat));
  INV_X1    g584(.A(G99gat), .ZN(new_n786));
  NAND4_X1  g585(.A1(new_n773), .A2(new_n786), .A3(new_n520), .A4(new_n703), .ZN(new_n787));
  NOR3_X1   g586(.A1(new_n718), .A2(new_n692), .A3(new_n776), .ZN(new_n788));
  OAI21_X1  g587(.A(new_n787), .B1(new_n788), .B2(new_n786), .ZN(G1338gat));
  INV_X1    g588(.A(G106gat), .ZN(new_n790));
  NAND4_X1  g589(.A1(new_n773), .A2(new_n790), .A3(new_n326), .A4(new_n703), .ZN(new_n791));
  NOR3_X1   g590(.A1(new_n718), .A2(new_n519), .A3(new_n776), .ZN(new_n792));
  OAI21_X1  g591(.A(new_n791), .B1(new_n792), .B2(new_n790), .ZN(new_n793));
  INV_X1    g592(.A(KEYINPUT53), .ZN(new_n794));
  INV_X1    g593(.A(KEYINPUT113), .ZN(new_n795));
  AOI21_X1  g594(.A(new_n794), .B1(new_n791), .B2(new_n795), .ZN(new_n796));
  NAND2_X1  g595(.A1(new_n793), .A2(new_n796), .ZN(new_n797));
  OAI221_X1 g596(.A(new_n791), .B1(new_n795), .B2(new_n794), .C1(new_n792), .C2(new_n790), .ZN(new_n798));
  NAND2_X1  g597(.A1(new_n797), .A2(new_n798), .ZN(G1339gat));
  INV_X1    g598(.A(KEYINPUT54), .ZN(new_n800));
  NAND3_X1  g599(.A1(new_n660), .A2(new_n800), .A3(new_n663), .ZN(new_n801));
  AND2_X1   g600(.A1(new_n801), .A2(new_n671), .ZN(new_n802));
  NAND4_X1  g601(.A1(new_n654), .A2(new_n658), .A3(new_n662), .A4(new_n659), .ZN(new_n803));
  NAND3_X1  g602(.A1(new_n664), .A2(KEYINPUT54), .A3(new_n803), .ZN(new_n804));
  NAND2_X1  g603(.A1(new_n802), .A2(new_n804), .ZN(new_n805));
  INV_X1    g604(.A(KEYINPUT55), .ZN(new_n806));
  NAND2_X1  g605(.A1(new_n805), .A2(new_n806), .ZN(new_n807));
  NAND4_X1  g606(.A1(new_n804), .A2(KEYINPUT55), .A3(new_n671), .A4(new_n801), .ZN(new_n808));
  NAND2_X1  g607(.A1(new_n808), .A2(new_n673), .ZN(new_n809));
  NOR2_X1   g608(.A1(new_n809), .A2(KEYINPUT114), .ZN(new_n810));
  INV_X1    g609(.A(KEYINPUT114), .ZN(new_n811));
  AOI21_X1  g610(.A(new_n811), .B1(new_n808), .B2(new_n673), .ZN(new_n812));
  OAI211_X1 g611(.A(new_n253), .B(new_n807), .C1(new_n810), .C2(new_n812), .ZN(new_n813));
  NAND3_X1  g612(.A1(new_n249), .A2(new_n207), .A3(new_n246), .ZN(new_n814));
  NOR2_X1   g613(.A1(new_n243), .A2(new_n244), .ZN(new_n815));
  AOI21_X1  g614(.A(new_n235), .B1(new_n234), .B2(new_n237), .ZN(new_n816));
  OAI21_X1  g615(.A(new_n206), .B1(new_n815), .B2(new_n816), .ZN(new_n817));
  NAND2_X1  g616(.A1(new_n814), .A2(new_n817), .ZN(new_n818));
  OR2_X1    g617(.A1(new_n818), .A2(new_n674), .ZN(new_n819));
  AOI21_X1  g618(.A(new_n622), .B1(new_n813), .B2(new_n819), .ZN(new_n820));
  AOI21_X1  g619(.A(new_n818), .B1(new_n617), .B2(new_n621), .ZN(new_n821));
  OAI211_X1 g620(.A(new_n821), .B(new_n807), .C1(new_n812), .C2(new_n810), .ZN(new_n822));
  INV_X1    g621(.A(new_n822), .ZN(new_n823));
  OAI21_X1  g622(.A(new_n755), .B1(new_n820), .B2(new_n823), .ZN(new_n824));
  OR2_X1    g623(.A1(new_n675), .A2(new_n253), .ZN(new_n825));
  AOI21_X1  g624(.A(new_n326), .B1(new_n824), .B2(new_n825), .ZN(new_n826));
  NOR2_X1   g625(.A1(new_n682), .A2(new_n456), .ZN(new_n827));
  NAND3_X1  g626(.A1(new_n826), .A2(new_n520), .A3(new_n827), .ZN(new_n828));
  NOR3_X1   g627(.A1(new_n828), .A2(new_n389), .A3(new_n257), .ZN(new_n829));
  NAND2_X1  g628(.A1(new_n824), .A2(new_n825), .ZN(new_n830));
  AND2_X1   g629(.A1(new_n830), .A2(new_n827), .ZN(new_n831));
  NAND2_X1  g630(.A1(new_n521), .A2(new_n523), .ZN(new_n832));
  NAND2_X1  g631(.A1(new_n831), .A2(new_n832), .ZN(new_n833));
  INV_X1    g632(.A(new_n833), .ZN(new_n834));
  NAND2_X1  g633(.A1(new_n834), .A2(new_n253), .ZN(new_n835));
  AOI21_X1  g634(.A(new_n829), .B1(new_n835), .B2(new_n389), .ZN(G1340gat));
  NOR3_X1   g635(.A1(new_n828), .A2(new_n390), .A3(new_n674), .ZN(new_n837));
  NAND2_X1  g636(.A1(new_n834), .A2(new_n703), .ZN(new_n838));
  AOI21_X1  g637(.A(new_n837), .B1(new_n838), .B2(new_n390), .ZN(G1341gat));
  OAI21_X1  g638(.A(G127gat), .B1(new_n828), .B2(new_n755), .ZN(new_n840));
  OR2_X1    g639(.A1(new_n755), .A2(G127gat), .ZN(new_n841));
  OAI21_X1  g640(.A(new_n840), .B1(new_n833), .B2(new_n841), .ZN(G1342gat));
  NOR3_X1   g641(.A1(new_n833), .A2(G134gat), .A3(new_n623), .ZN(new_n843));
  INV_X1    g642(.A(new_n843), .ZN(new_n844));
  OR2_X1    g643(.A1(new_n844), .A2(KEYINPUT56), .ZN(new_n845));
  OAI21_X1  g644(.A(G134gat), .B1(new_n828), .B2(new_n623), .ZN(new_n846));
  NAND2_X1  g645(.A1(new_n844), .A2(KEYINPUT56), .ZN(new_n847));
  NAND3_X1  g646(.A1(new_n845), .A2(new_n846), .A3(new_n847), .ZN(G1343gat));
  NAND2_X1  g647(.A1(new_n692), .A2(new_n326), .ZN(new_n849));
  INV_X1    g648(.A(new_n849), .ZN(new_n850));
  NAND2_X1  g649(.A1(new_n831), .A2(new_n850), .ZN(new_n851));
  INV_X1    g650(.A(new_n851), .ZN(new_n852));
  NAND3_X1  g651(.A1(new_n852), .A2(new_n284), .A3(new_n702), .ZN(new_n853));
  INV_X1    g652(.A(KEYINPUT117), .ZN(new_n854));
  OAI21_X1  g653(.A(new_n853), .B1(new_n854), .B2(KEYINPUT58), .ZN(new_n855));
  NAND2_X1  g654(.A1(new_n827), .A2(new_n692), .ZN(new_n856));
  INV_X1    g655(.A(new_n856), .ZN(new_n857));
  NAND2_X1  g656(.A1(new_n326), .A2(KEYINPUT57), .ZN(new_n858));
  NAND4_X1  g657(.A1(new_n807), .A2(KEYINPUT115), .A3(new_n673), .A4(new_n808), .ZN(new_n859));
  INV_X1    g658(.A(KEYINPUT115), .ZN(new_n860));
  AOI21_X1  g659(.A(KEYINPUT55), .B1(new_n802), .B2(new_n804), .ZN(new_n861));
  OAI21_X1  g660(.A(new_n860), .B1(new_n809), .B2(new_n861), .ZN(new_n862));
  NAND4_X1  g661(.A1(new_n859), .A2(new_n862), .A3(new_n255), .A4(new_n256), .ZN(new_n863));
  AOI21_X1  g662(.A(new_n622), .B1(new_n863), .B2(new_n819), .ZN(new_n864));
  OAI21_X1  g663(.A(new_n755), .B1(new_n864), .B2(new_n823), .ZN(new_n865));
  AOI21_X1  g664(.A(new_n858), .B1(new_n865), .B2(new_n825), .ZN(new_n866));
  INV_X1    g665(.A(KEYINPUT116), .ZN(new_n867));
  AOI21_X1  g666(.A(new_n519), .B1(new_n824), .B2(new_n825), .ZN(new_n868));
  OAI22_X1  g667(.A1(new_n866), .A2(new_n867), .B1(new_n868), .B2(KEYINPUT57), .ZN(new_n869));
  AND2_X1   g668(.A1(new_n866), .A2(new_n867), .ZN(new_n870));
  OAI21_X1  g669(.A(new_n857), .B1(new_n869), .B2(new_n870), .ZN(new_n871));
  INV_X1    g670(.A(new_n871), .ZN(new_n872));
  NAND2_X1  g671(.A1(new_n872), .A2(new_n253), .ZN(new_n873));
  INV_X1    g672(.A(KEYINPUT58), .ZN(new_n874));
  NOR2_X1   g673(.A1(new_n874), .A2(new_n284), .ZN(new_n875));
  AOI21_X1  g674(.A(new_n855), .B1(new_n873), .B2(new_n875), .ZN(new_n876));
  OAI21_X1  g675(.A(G141gat), .B1(new_n871), .B2(new_n257), .ZN(new_n877));
  OAI21_X1  g676(.A(new_n877), .B1(new_n854), .B2(new_n853), .ZN(new_n878));
  AOI21_X1  g677(.A(new_n876), .B1(new_n874), .B2(new_n878), .ZN(G1344gat));
  INV_X1    g678(.A(KEYINPUT59), .ZN(new_n880));
  NAND2_X1  g679(.A1(new_n830), .A2(new_n326), .ZN(new_n881));
  NAND2_X1  g680(.A1(new_n881), .A2(KEYINPUT57), .ZN(new_n882));
  OAI21_X1  g681(.A(new_n865), .B1(new_n678), .B2(new_n702), .ZN(new_n883));
  INV_X1    g682(.A(KEYINPUT57), .ZN(new_n884));
  NAND3_X1  g683(.A1(new_n883), .A2(new_n884), .A3(new_n326), .ZN(new_n885));
  NAND4_X1  g684(.A1(new_n882), .A2(new_n885), .A3(new_n703), .A4(new_n857), .ZN(new_n886));
  AOI21_X1  g685(.A(new_n880), .B1(new_n886), .B2(G148gat), .ZN(new_n887));
  OAI211_X1 g686(.A(new_n703), .B(new_n857), .C1(new_n869), .C2(new_n870), .ZN(new_n888));
  NOR2_X1   g687(.A1(new_n286), .A2(KEYINPUT59), .ZN(new_n889));
  NAND2_X1  g688(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  INV_X1    g689(.A(KEYINPUT118), .ZN(new_n891));
  NAND2_X1  g690(.A1(new_n890), .A2(new_n891), .ZN(new_n892));
  NAND3_X1  g691(.A1(new_n888), .A2(KEYINPUT118), .A3(new_n889), .ZN(new_n893));
  AOI21_X1  g692(.A(new_n887), .B1(new_n892), .B2(new_n893), .ZN(new_n894));
  NOR3_X1   g693(.A1(new_n851), .A2(G148gat), .A3(new_n674), .ZN(new_n895));
  OAI21_X1  g694(.A(KEYINPUT119), .B1(new_n894), .B2(new_n895), .ZN(new_n896));
  INV_X1    g695(.A(KEYINPUT119), .ZN(new_n897));
  INV_X1    g696(.A(new_n895), .ZN(new_n898));
  AND3_X1   g697(.A1(new_n888), .A2(KEYINPUT118), .A3(new_n889), .ZN(new_n899));
  AOI21_X1  g698(.A(KEYINPUT118), .B1(new_n888), .B2(new_n889), .ZN(new_n900));
  NOR2_X1   g699(.A1(new_n899), .A2(new_n900), .ZN(new_n901));
  OAI211_X1 g700(.A(new_n897), .B(new_n898), .C1(new_n901), .C2(new_n887), .ZN(new_n902));
  NAND2_X1  g701(.A1(new_n896), .A2(new_n902), .ZN(G1345gat));
  AOI21_X1  g702(.A(G155gat), .B1(new_n852), .B2(new_n650), .ZN(new_n904));
  NAND2_X1  g703(.A1(new_n650), .A2(G155gat), .ZN(new_n905));
  XNOR2_X1  g704(.A(new_n905), .B(KEYINPUT120), .ZN(new_n906));
  AOI21_X1  g705(.A(new_n904), .B1(new_n872), .B2(new_n906), .ZN(G1346gat));
  NAND3_X1  g706(.A1(new_n852), .A2(new_n280), .A3(new_n622), .ZN(new_n908));
  INV_X1    g707(.A(KEYINPUT121), .ZN(new_n909));
  OAI21_X1  g708(.A(new_n909), .B1(new_n871), .B2(new_n623), .ZN(new_n910));
  NAND2_X1  g709(.A1(new_n910), .A2(G162gat), .ZN(new_n911));
  NOR3_X1   g710(.A1(new_n871), .A2(new_n909), .A3(new_n623), .ZN(new_n912));
  OAI21_X1  g711(.A(new_n908), .B1(new_n911), .B2(new_n912), .ZN(G1347gat));
  NAND4_X1  g712(.A1(new_n826), .A2(new_n682), .A3(new_n456), .A4(new_n520), .ZN(new_n914));
  NOR3_X1   g713(.A1(new_n914), .A2(new_n371), .A3(new_n257), .ZN(new_n915));
  AOI21_X1  g714(.A(new_n681), .B1(new_n824), .B2(new_n825), .ZN(new_n916));
  NAND3_X1  g715(.A1(new_n916), .A2(new_n456), .A3(new_n832), .ZN(new_n917));
  XNOR2_X1  g716(.A(new_n917), .B(KEYINPUT122), .ZN(new_n918));
  INV_X1    g717(.A(new_n918), .ZN(new_n919));
  NAND2_X1  g718(.A1(new_n919), .A2(new_n253), .ZN(new_n920));
  AOI21_X1  g719(.A(new_n915), .B1(new_n920), .B2(new_n371), .ZN(G1348gat));
  AOI21_X1  g720(.A(G176gat), .B1(new_n919), .B2(new_n703), .ZN(new_n922));
  NOR3_X1   g721(.A1(new_n914), .A2(new_n372), .A3(new_n674), .ZN(new_n923));
  XNOR2_X1  g722(.A(new_n923), .B(KEYINPUT123), .ZN(new_n924));
  NOR2_X1   g723(.A1(new_n922), .A2(new_n924), .ZN(G1349gat));
  OAI21_X1  g724(.A(G183gat), .B1(new_n914), .B2(new_n755), .ZN(new_n926));
  NAND3_X1  g725(.A1(new_n650), .A2(new_n363), .A3(new_n365), .ZN(new_n927));
  OAI21_X1  g726(.A(new_n926), .B1(new_n917), .B2(new_n927), .ZN(new_n928));
  OAI21_X1  g727(.A(new_n928), .B1(KEYINPUT124), .B2(KEYINPUT60), .ZN(new_n929));
  NAND2_X1  g728(.A1(KEYINPUT124), .A2(KEYINPUT60), .ZN(new_n930));
  XNOR2_X1  g729(.A(new_n929), .B(new_n930), .ZN(G1350gat));
  OAI21_X1  g730(.A(G190gat), .B1(new_n914), .B2(new_n623), .ZN(new_n932));
  OR2_X1    g731(.A1(new_n932), .A2(KEYINPUT125), .ZN(new_n933));
  NAND2_X1  g732(.A1(new_n932), .A2(KEYINPUT125), .ZN(new_n934));
  NAND3_X1  g733(.A1(new_n933), .A2(KEYINPUT61), .A3(new_n934), .ZN(new_n935));
  NAND3_X1  g734(.A1(new_n919), .A2(new_n366), .A3(new_n622), .ZN(new_n936));
  OAI211_X1 g735(.A(new_n935), .B(new_n936), .C1(KEYINPUT61), .C2(new_n934), .ZN(G1351gat));
  NAND3_X1  g736(.A1(new_n850), .A2(KEYINPUT126), .A3(new_n456), .ZN(new_n938));
  INV_X1    g737(.A(KEYINPUT126), .ZN(new_n939));
  OAI21_X1  g738(.A(new_n939), .B1(new_n849), .B2(new_n457), .ZN(new_n940));
  NAND3_X1  g739(.A1(new_n916), .A2(new_n938), .A3(new_n940), .ZN(new_n941));
  INV_X1    g740(.A(new_n941), .ZN(new_n942));
  AOI21_X1  g741(.A(G197gat), .B1(new_n942), .B2(new_n253), .ZN(new_n943));
  NAND2_X1  g742(.A1(new_n882), .A2(new_n885), .ZN(new_n944));
  NAND3_X1  g743(.A1(new_n682), .A2(new_n692), .A3(new_n456), .ZN(new_n945));
  NOR2_X1   g744(.A1(new_n944), .A2(new_n945), .ZN(new_n946));
  AND2_X1   g745(.A1(new_n702), .A2(G197gat), .ZN(new_n947));
  AOI21_X1  g746(.A(new_n943), .B1(new_n946), .B2(new_n947), .ZN(G1352gat));
  NOR3_X1   g747(.A1(new_n941), .A2(G204gat), .A3(new_n674), .ZN(new_n949));
  XNOR2_X1  g748(.A(new_n949), .B(KEYINPUT62), .ZN(new_n950));
  INV_X1    g749(.A(G204gat), .ZN(new_n951));
  NOR3_X1   g750(.A1(new_n944), .A2(new_n674), .A3(new_n945), .ZN(new_n952));
  OAI21_X1  g751(.A(new_n950), .B1(new_n951), .B2(new_n952), .ZN(G1353gat));
  OAI21_X1  g752(.A(G211gat), .B1(KEYINPUT127), .B2(KEYINPUT63), .ZN(new_n954));
  AOI21_X1  g753(.A(new_n954), .B1(new_n946), .B2(new_n650), .ZN(new_n955));
  NAND2_X1  g754(.A1(KEYINPUT127), .A2(KEYINPUT63), .ZN(new_n956));
  OR2_X1    g755(.A1(new_n955), .A2(new_n956), .ZN(new_n957));
  NAND2_X1  g756(.A1(new_n955), .A2(new_n956), .ZN(new_n958));
  NAND3_X1  g757(.A1(new_n942), .A2(new_n272), .A3(new_n650), .ZN(new_n959));
  NAND3_X1  g758(.A1(new_n957), .A2(new_n958), .A3(new_n959), .ZN(G1354gat));
  NAND3_X1  g759(.A1(new_n942), .A2(new_n273), .A3(new_n622), .ZN(new_n961));
  NOR3_X1   g760(.A1(new_n944), .A2(new_n623), .A3(new_n945), .ZN(new_n962));
  OAI21_X1  g761(.A(new_n961), .B1(new_n962), .B2(new_n273), .ZN(G1355gat));
endmodule


