//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 0 0 0 0 0 0 0 1 0 0 0 1 0 0 0 0 1 0 1 1 0 0 1 0 0 1 1 1 1 1 0 1 0 1 1 1 1 0 0 1 1 0 1 1 0 0 1 0 1 1 1 1 1 0 0 0 1 0 1 0 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:33:15 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n442, new_n444, new_n448, new_n449, new_n451, new_n454, new_n455,
    new_n456, new_n457, new_n458, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n525,
    new_n526, new_n527, new_n528, new_n529, new_n530, new_n532, new_n533,
    new_n534, new_n535, new_n536, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n548, new_n549, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n569, new_n570,
    new_n571, new_n572, new_n573, new_n574, new_n575, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n599, new_n600, new_n603, new_n605,
    new_n607, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n639, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n819, new_n820, new_n821, new_n822, new_n823, new_n824,
    new_n825, new_n826, new_n827, new_n828, new_n829, new_n830, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n896, new_n897, new_n898,
    new_n899, new_n900, new_n901, new_n902, new_n903, new_n904, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1144, new_n1145, new_n1146;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  XNOR2_X1  g009(.A(KEYINPUT64), .B(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  AND2_X1   g016(.A1(G2072), .A2(G2078), .ZN(new_n442));
  NAND3_X1  g017(.A1(new_n442), .A2(G2084), .A3(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(new_n444));
  XOR2_X1   g019(.A(new_n444), .B(KEYINPUT65), .Z(G259));
  BUF_X1    g020(.A(G452), .Z(G391));
  AND2_X1   g021(.A1(G94), .A2(G452), .ZN(G173));
  XNOR2_X1  g022(.A(KEYINPUT66), .B(KEYINPUT1), .ZN(new_n448));
  NAND2_X1  g023(.A1(G7), .A2(G661), .ZN(new_n449));
  XNOR2_X1  g024(.A(new_n448), .B(new_n449), .ZN(G223));
  INV_X1    g025(.A(new_n449), .ZN(new_n451));
  NAND2_X1  g026(.A1(new_n451), .A2(G567), .ZN(G234));
  NAND2_X1  g027(.A1(new_n451), .A2(G2106), .ZN(G217));
  NOR4_X1   g028(.A1(G219), .A2(G220), .A3(G218), .A4(G221), .ZN(new_n454));
  XOR2_X1   g029(.A(new_n454), .B(KEYINPUT2), .Z(new_n455));
  NOR4_X1   g030(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n456));
  INV_X1    g031(.A(new_n456), .ZN(new_n457));
  OR2_X1    g032(.A1(new_n455), .A2(new_n457), .ZN(new_n458));
  XOR2_X1   g033(.A(new_n458), .B(KEYINPUT67), .Z(G261));
  INV_X1    g034(.A(G261), .ZN(G325));
  AOI22_X1  g035(.A1(new_n455), .A2(G2106), .B1(G567), .B2(new_n457), .ZN(G319));
  INV_X1    g036(.A(G2104), .ZN(new_n462));
  NOR2_X1   g037(.A1(new_n462), .A2(G2105), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n463), .A2(G101), .ZN(new_n464));
  INV_X1    g039(.A(KEYINPUT70), .ZN(new_n465));
  XNOR2_X1  g040(.A(new_n464), .B(new_n465), .ZN(new_n466));
  NAND2_X1  g041(.A1(G113), .A2(G2104), .ZN(new_n467));
  XNOR2_X1  g042(.A(new_n467), .B(KEYINPUT68), .ZN(new_n468));
  INV_X1    g043(.A(G125), .ZN(new_n469));
  INV_X1    g044(.A(KEYINPUT3), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n470), .A2(new_n462), .ZN(new_n471));
  NAND2_X1  g046(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n472));
  AOI21_X1  g047(.A(new_n469), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  OAI21_X1  g048(.A(G2105), .B1(new_n468), .B2(new_n473), .ZN(new_n474));
  OAI21_X1  g049(.A(new_n470), .B1(new_n462), .B2(KEYINPUT69), .ZN(new_n475));
  INV_X1    g050(.A(KEYINPUT69), .ZN(new_n476));
  NAND3_X1  g051(.A1(new_n476), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n477));
  AOI21_X1  g052(.A(G2105), .B1(new_n475), .B2(new_n477), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n478), .A2(G137), .ZN(new_n479));
  AND3_X1   g054(.A1(new_n466), .A2(new_n474), .A3(new_n479), .ZN(G160));
  NAND2_X1  g055(.A1(new_n478), .A2(G136), .ZN(new_n481));
  INV_X1    g056(.A(G2105), .ZN(new_n482));
  NOR2_X1   g057(.A1(new_n482), .A2(G112), .ZN(new_n483));
  OAI21_X1  g058(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n484));
  OAI21_X1  g059(.A(new_n481), .B1(new_n483), .B2(new_n484), .ZN(new_n485));
  AOI21_X1  g060(.A(new_n482), .B1(new_n475), .B2(new_n477), .ZN(new_n486));
  XOR2_X1   g061(.A(new_n486), .B(KEYINPUT71), .Z(new_n487));
  AOI21_X1  g062(.A(new_n485), .B1(new_n487), .B2(G124), .ZN(G162));
  NAND2_X1  g063(.A1(new_n482), .A2(G138), .ZN(new_n489));
  INV_X1    g064(.A(new_n489), .ZN(new_n490));
  AND3_X1   g065(.A1(new_n476), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n491));
  AOI21_X1  g066(.A(KEYINPUT3), .B1(new_n476), .B2(G2104), .ZN(new_n492));
  OAI21_X1  g067(.A(new_n490), .B1(new_n491), .B2(new_n492), .ZN(new_n493));
  INV_X1    g068(.A(KEYINPUT72), .ZN(new_n494));
  NAND3_X1  g069(.A1(new_n493), .A2(new_n494), .A3(KEYINPUT4), .ZN(new_n495));
  AOI21_X1  g070(.A(new_n489), .B1(new_n475), .B2(new_n477), .ZN(new_n496));
  INV_X1    g071(.A(KEYINPUT4), .ZN(new_n497));
  OAI21_X1  g072(.A(KEYINPUT72), .B1(new_n496), .B2(new_n497), .ZN(new_n498));
  NAND2_X1  g073(.A1(new_n471), .A2(new_n472), .ZN(new_n499));
  NAND3_X1  g074(.A1(new_n499), .A2(new_n497), .A3(new_n490), .ZN(new_n500));
  NAND3_X1  g075(.A1(new_n495), .A2(new_n498), .A3(new_n500), .ZN(new_n501));
  OAI21_X1  g076(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n502));
  INV_X1    g077(.A(G114), .ZN(new_n503));
  AOI21_X1  g078(.A(new_n502), .B1(new_n503), .B2(G2105), .ZN(new_n504));
  AOI21_X1  g079(.A(new_n504), .B1(new_n486), .B2(G126), .ZN(new_n505));
  NAND2_X1  g080(.A1(new_n501), .A2(new_n505), .ZN(new_n506));
  INV_X1    g081(.A(new_n506), .ZN(G164));
  AND2_X1   g082(.A1(KEYINPUT6), .A2(G651), .ZN(new_n508));
  NOR2_X1   g083(.A1(KEYINPUT6), .A2(G651), .ZN(new_n509));
  OR2_X1    g084(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  NAND2_X1  g085(.A1(KEYINPUT73), .A2(KEYINPUT5), .ZN(new_n511));
  INV_X1    g086(.A(G543), .ZN(new_n512));
  NAND2_X1  g087(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  NAND3_X1  g088(.A1(KEYINPUT73), .A2(KEYINPUT5), .A3(G543), .ZN(new_n514));
  NAND2_X1  g089(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  AND2_X1   g090(.A1(new_n510), .A2(new_n515), .ZN(new_n516));
  NAND2_X1  g091(.A1(new_n516), .A2(G88), .ZN(new_n517));
  INV_X1    g092(.A(G50), .ZN(new_n518));
  NAND2_X1  g093(.A1(new_n510), .A2(G543), .ZN(new_n519));
  OAI21_X1  g094(.A(new_n517), .B1(new_n518), .B2(new_n519), .ZN(new_n520));
  AOI22_X1  g095(.A1(new_n515), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n521));
  INV_X1    g096(.A(G651), .ZN(new_n522));
  NOR2_X1   g097(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  NOR2_X1   g098(.A1(new_n520), .A2(new_n523), .ZN(G166));
  AND2_X1   g099(.A1(new_n516), .A2(G89), .ZN(new_n525));
  NAND3_X1  g100(.A1(new_n515), .A2(G63), .A3(G651), .ZN(new_n526));
  NAND3_X1  g101(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n527));
  XNOR2_X1  g102(.A(new_n527), .B(KEYINPUT7), .ZN(new_n528));
  INV_X1    g103(.A(G51), .ZN(new_n529));
  OAI211_X1 g104(.A(new_n526), .B(new_n528), .C1(new_n519), .C2(new_n529), .ZN(new_n530));
  NOR2_X1   g105(.A1(new_n525), .A2(new_n530), .ZN(G168));
  NAND2_X1  g106(.A1(new_n516), .A2(G90), .ZN(new_n532));
  INV_X1    g107(.A(G52), .ZN(new_n533));
  OAI21_X1  g108(.A(new_n532), .B1(new_n533), .B2(new_n519), .ZN(new_n534));
  AOI22_X1  g109(.A1(new_n515), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n535));
  NOR2_X1   g110(.A1(new_n535), .A2(new_n522), .ZN(new_n536));
  NOR2_X1   g111(.A1(new_n534), .A2(new_n536), .ZN(G171));
  INV_X1    g112(.A(new_n519), .ZN(new_n538));
  AOI22_X1  g113(.A1(G43), .A2(new_n538), .B1(new_n516), .B2(G81), .ZN(new_n539));
  AND2_X1   g114(.A1(G68), .A2(G543), .ZN(new_n540));
  AOI21_X1  g115(.A(new_n540), .B1(new_n515), .B2(G56), .ZN(new_n541));
  OR3_X1    g116(.A1(new_n541), .A2(KEYINPUT74), .A3(new_n522), .ZN(new_n542));
  OAI21_X1  g117(.A(KEYINPUT74), .B1(new_n541), .B2(new_n522), .ZN(new_n543));
  NAND3_X1  g118(.A1(new_n539), .A2(new_n542), .A3(new_n543), .ZN(new_n544));
  XNOR2_X1  g119(.A(new_n544), .B(KEYINPUT75), .ZN(new_n545));
  NAND2_X1  g120(.A1(new_n545), .A2(G860), .ZN(G153));
  NAND4_X1  g121(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g122(.A1(G1), .A2(G3), .ZN(new_n548));
  XNOR2_X1  g123(.A(new_n548), .B(KEYINPUT8), .ZN(new_n549));
  NAND4_X1  g124(.A1(G319), .A2(G483), .A3(G661), .A4(new_n549), .ZN(G188));
  NAND2_X1  g125(.A1(new_n538), .A2(G53), .ZN(new_n551));
  XOR2_X1   g126(.A(new_n551), .B(KEYINPUT9), .Z(new_n552));
  NAND2_X1  g127(.A1(new_n516), .A2(G91), .ZN(new_n553));
  XOR2_X1   g128(.A(KEYINPUT76), .B(G65), .Z(new_n554));
  AOI22_X1  g129(.A1(new_n554), .A2(new_n515), .B1(G78), .B2(G543), .ZN(new_n555));
  OAI21_X1  g130(.A(new_n553), .B1(new_n522), .B2(new_n555), .ZN(new_n556));
  OR2_X1    g131(.A1(new_n552), .A2(new_n556), .ZN(G299));
  INV_X1    g132(.A(G171), .ZN(G301));
  INV_X1    g133(.A(G168), .ZN(G286));
  INV_X1    g134(.A(G166), .ZN(G303));
  INV_X1    g135(.A(KEYINPUT77), .ZN(new_n561));
  NAND3_X1  g136(.A1(new_n538), .A2(new_n561), .A3(G49), .ZN(new_n562));
  INV_X1    g137(.A(G49), .ZN(new_n563));
  OAI21_X1  g138(.A(KEYINPUT77), .B1(new_n519), .B2(new_n563), .ZN(new_n564));
  NAND2_X1  g139(.A1(new_n562), .A2(new_n564), .ZN(new_n565));
  OR2_X1    g140(.A1(new_n515), .A2(G74), .ZN(new_n566));
  AOI22_X1  g141(.A1(G87), .A2(new_n516), .B1(new_n566), .B2(G651), .ZN(new_n567));
  NAND2_X1  g142(.A1(new_n565), .A2(new_n567), .ZN(G288));
  INV_X1    g143(.A(G61), .ZN(new_n569));
  AOI21_X1  g144(.A(new_n569), .B1(new_n513), .B2(new_n514), .ZN(new_n570));
  NAND2_X1  g145(.A1(G73), .A2(G543), .ZN(new_n571));
  INV_X1    g146(.A(new_n571), .ZN(new_n572));
  OAI21_X1  g147(.A(G651), .B1(new_n570), .B2(new_n572), .ZN(new_n573));
  NAND3_X1  g148(.A1(new_n510), .A2(G86), .A3(new_n515), .ZN(new_n574));
  NAND3_X1  g149(.A1(new_n510), .A2(G48), .A3(G543), .ZN(new_n575));
  NAND3_X1  g150(.A1(new_n573), .A2(new_n574), .A3(new_n575), .ZN(G305));
  XOR2_X1   g151(.A(KEYINPUT79), .B(G47), .Z(new_n577));
  AOI22_X1  g152(.A1(new_n538), .A2(new_n577), .B1(new_n516), .B2(G85), .ZN(new_n578));
  INV_X1    g153(.A(KEYINPUT78), .ZN(new_n579));
  NAND2_X1  g154(.A1(new_n515), .A2(G60), .ZN(new_n580));
  NAND2_X1  g155(.A1(G72), .A2(G543), .ZN(new_n581));
  AOI21_X1  g156(.A(new_n522), .B1(new_n580), .B2(new_n581), .ZN(new_n582));
  OAI21_X1  g157(.A(new_n578), .B1(new_n579), .B2(new_n582), .ZN(new_n583));
  AND2_X1   g158(.A1(new_n582), .A2(new_n579), .ZN(new_n584));
  NOR2_X1   g159(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  INV_X1    g160(.A(new_n585), .ZN(G290));
  NAND2_X1  g161(.A1(G301), .A2(G868), .ZN(new_n587));
  AOI22_X1  g162(.A1(new_n515), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n588));
  INV_X1    g163(.A(G54), .ZN(new_n589));
  OAI22_X1  g164(.A1(new_n588), .A2(new_n522), .B1(new_n519), .B2(new_n589), .ZN(new_n590));
  XNOR2_X1  g165(.A(new_n590), .B(KEYINPUT80), .ZN(new_n591));
  NAND2_X1  g166(.A1(new_n516), .A2(G92), .ZN(new_n592));
  INV_X1    g167(.A(KEYINPUT10), .ZN(new_n593));
  XNOR2_X1  g168(.A(new_n592), .B(new_n593), .ZN(new_n594));
  NAND2_X1  g169(.A1(new_n591), .A2(new_n594), .ZN(new_n595));
  INV_X1    g170(.A(new_n595), .ZN(new_n596));
  OAI21_X1  g171(.A(new_n587), .B1(new_n596), .B2(G868), .ZN(G284));
  OAI21_X1  g172(.A(new_n587), .B1(new_n596), .B2(G868), .ZN(G321));
  NAND2_X1  g173(.A1(G286), .A2(G868), .ZN(new_n599));
  NOR2_X1   g174(.A1(new_n552), .A2(new_n556), .ZN(new_n600));
  OAI21_X1  g175(.A(new_n599), .B1(new_n600), .B2(G868), .ZN(G297));
  XOR2_X1   g176(.A(G297), .B(KEYINPUT81), .Z(G280));
  INV_X1    g177(.A(G559), .ZN(new_n603));
  OAI21_X1  g178(.A(new_n596), .B1(new_n603), .B2(G860), .ZN(G148));
  OAI21_X1  g179(.A(G868), .B1(new_n595), .B2(G559), .ZN(new_n605));
  OAI21_X1  g180(.A(new_n605), .B1(G868), .B2(new_n545), .ZN(G323));
  XNOR2_X1  g181(.A(KEYINPUT82), .B(KEYINPUT11), .ZN(new_n607));
  XNOR2_X1  g182(.A(G323), .B(new_n607), .ZN(G282));
  NAND2_X1  g183(.A1(new_n499), .A2(new_n463), .ZN(new_n609));
  XOR2_X1   g184(.A(KEYINPUT83), .B(KEYINPUT12), .Z(new_n610));
  XNOR2_X1  g185(.A(new_n609), .B(new_n610), .ZN(new_n611));
  XNOR2_X1  g186(.A(new_n611), .B(KEYINPUT13), .ZN(new_n612));
  XNOR2_X1  g187(.A(new_n612), .B(G2100), .ZN(new_n613));
  NAND2_X1  g188(.A1(new_n487), .A2(G123), .ZN(new_n614));
  OAI21_X1  g189(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n615));
  INV_X1    g190(.A(G111), .ZN(new_n616));
  AOI21_X1  g191(.A(new_n615), .B1(new_n616), .B2(G2105), .ZN(new_n617));
  AOI21_X1  g192(.A(new_n617), .B1(new_n478), .B2(G135), .ZN(new_n618));
  NAND2_X1  g193(.A1(new_n614), .A2(new_n618), .ZN(new_n619));
  XOR2_X1   g194(.A(KEYINPUT84), .B(G2096), .Z(new_n620));
  XNOR2_X1  g195(.A(new_n619), .B(new_n620), .ZN(new_n621));
  NAND2_X1  g196(.A1(new_n613), .A2(new_n621), .ZN(G156));
  XOR2_X1   g197(.A(G2451), .B(G2454), .Z(new_n623));
  XNOR2_X1  g198(.A(new_n623), .B(KEYINPUT16), .ZN(new_n624));
  XNOR2_X1  g199(.A(G1341), .B(G1348), .ZN(new_n625));
  XNOR2_X1  g200(.A(new_n624), .B(new_n625), .ZN(new_n626));
  INV_X1    g201(.A(KEYINPUT14), .ZN(new_n627));
  XNOR2_X1  g202(.A(G2427), .B(G2438), .ZN(new_n628));
  XNOR2_X1  g203(.A(new_n628), .B(G2430), .ZN(new_n629));
  XNOR2_X1  g204(.A(KEYINPUT15), .B(G2435), .ZN(new_n630));
  AOI21_X1  g205(.A(new_n627), .B1(new_n629), .B2(new_n630), .ZN(new_n631));
  OAI21_X1  g206(.A(new_n631), .B1(new_n630), .B2(new_n629), .ZN(new_n632));
  XOR2_X1   g207(.A(new_n626), .B(new_n632), .Z(new_n633));
  INV_X1    g208(.A(new_n633), .ZN(new_n634));
  XNOR2_X1  g209(.A(G2443), .B(G2446), .ZN(new_n635));
  INV_X1    g210(.A(new_n635), .ZN(new_n636));
  OAI21_X1  g211(.A(G14), .B1(new_n634), .B2(new_n636), .ZN(new_n637));
  AOI21_X1  g212(.A(new_n637), .B1(new_n636), .B2(new_n634), .ZN(G401));
  XOR2_X1   g213(.A(G2067), .B(G2678), .Z(new_n639));
  XNOR2_X1  g214(.A(new_n639), .B(KEYINPUT85), .ZN(new_n640));
  NOR2_X1   g215(.A1(G2072), .A2(G2078), .ZN(new_n641));
  NOR2_X1   g216(.A1(new_n442), .A2(new_n641), .ZN(new_n642));
  XOR2_X1   g217(.A(G2084), .B(G2090), .Z(new_n643));
  INV_X1    g218(.A(new_n643), .ZN(new_n644));
  NOR3_X1   g219(.A1(new_n640), .A2(new_n642), .A3(new_n644), .ZN(new_n645));
  XNOR2_X1  g220(.A(new_n645), .B(KEYINPUT18), .ZN(new_n646));
  NAND2_X1  g221(.A1(new_n640), .A2(new_n642), .ZN(new_n647));
  XNOR2_X1  g222(.A(new_n642), .B(KEYINPUT17), .ZN(new_n648));
  OAI211_X1 g223(.A(new_n647), .B(new_n644), .C1(new_n640), .C2(new_n648), .ZN(new_n649));
  NAND3_X1  g224(.A1(new_n640), .A2(new_n648), .A3(new_n643), .ZN(new_n650));
  NAND3_X1  g225(.A1(new_n646), .A2(new_n649), .A3(new_n650), .ZN(new_n651));
  XNOR2_X1  g226(.A(G2096), .B(G2100), .ZN(new_n652));
  XNOR2_X1  g227(.A(new_n652), .B(KEYINPUT86), .ZN(new_n653));
  XOR2_X1   g228(.A(new_n653), .B(KEYINPUT87), .Z(new_n654));
  XNOR2_X1  g229(.A(new_n651), .B(new_n654), .ZN(G227));
  XOR2_X1   g230(.A(G1971), .B(G1976), .Z(new_n656));
  XNOR2_X1  g231(.A(new_n656), .B(KEYINPUT19), .ZN(new_n657));
  XNOR2_X1  g232(.A(G1956), .B(G2474), .ZN(new_n658));
  XNOR2_X1  g233(.A(G1961), .B(G1966), .ZN(new_n659));
  NOR2_X1   g234(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  AND2_X1   g235(.A1(new_n658), .A2(new_n659), .ZN(new_n661));
  NOR3_X1   g236(.A1(new_n657), .A2(new_n660), .A3(new_n661), .ZN(new_n662));
  NAND2_X1  g237(.A1(new_n657), .A2(new_n660), .ZN(new_n663));
  XOR2_X1   g238(.A(new_n663), .B(KEYINPUT20), .Z(new_n664));
  AOI211_X1 g239(.A(new_n662), .B(new_n664), .C1(new_n657), .C2(new_n661), .ZN(new_n665));
  XOR2_X1   g240(.A(G1991), .B(G1996), .Z(new_n666));
  XNOR2_X1  g241(.A(new_n665), .B(new_n666), .ZN(new_n667));
  XOR2_X1   g242(.A(G1981), .B(G1986), .Z(new_n668));
  XNOR2_X1  g243(.A(new_n668), .B(KEYINPUT88), .ZN(new_n669));
  XOR2_X1   g244(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n670));
  XNOR2_X1  g245(.A(new_n669), .B(new_n670), .ZN(new_n671));
  XNOR2_X1  g246(.A(new_n667), .B(new_n671), .ZN(G229));
  INV_X1    g247(.A(G16), .ZN(new_n673));
  NAND2_X1  g248(.A1(new_n673), .A2(G20), .ZN(new_n674));
  XOR2_X1   g249(.A(new_n674), .B(KEYINPUT23), .Z(new_n675));
  AOI21_X1  g250(.A(new_n675), .B1(G299), .B2(G16), .ZN(new_n676));
  XNOR2_X1  g251(.A(new_n676), .B(G1956), .ZN(new_n677));
  INV_X1    g252(.A(G29), .ZN(new_n678));
  NAND2_X1  g253(.A1(new_n678), .A2(G26), .ZN(new_n679));
  XNOR2_X1  g254(.A(new_n679), .B(KEYINPUT28), .ZN(new_n680));
  OR2_X1    g255(.A1(G104), .A2(G2105), .ZN(new_n681));
  OAI211_X1 g256(.A(new_n681), .B(G2104), .C1(G116), .C2(new_n482), .ZN(new_n682));
  XNOR2_X1  g257(.A(new_n682), .B(KEYINPUT91), .ZN(new_n683));
  NAND2_X1  g258(.A1(new_n478), .A2(G140), .ZN(new_n684));
  NAND2_X1  g259(.A1(new_n683), .A2(new_n684), .ZN(new_n685));
  AOI21_X1  g260(.A(new_n685), .B1(G128), .B2(new_n487), .ZN(new_n686));
  OAI21_X1  g261(.A(new_n680), .B1(new_n686), .B2(new_n678), .ZN(new_n687));
  INV_X1    g262(.A(G2067), .ZN(new_n688));
  XNOR2_X1  g263(.A(new_n687), .B(new_n688), .ZN(new_n689));
  INV_X1    g264(.A(G2078), .ZN(new_n690));
  NOR2_X1   g265(.A1(G164), .A2(new_n678), .ZN(new_n691));
  AOI21_X1  g266(.A(new_n691), .B1(G27), .B2(new_n678), .ZN(new_n692));
  OAI211_X1 g267(.A(new_n677), .B(new_n689), .C1(new_n690), .C2(new_n692), .ZN(new_n693));
  INV_X1    g268(.A(KEYINPUT95), .ZN(new_n694));
  OR3_X1    g269(.A1(new_n694), .A2(G5), .A3(G16), .ZN(new_n695));
  OAI21_X1  g270(.A(new_n694), .B1(G5), .B2(G16), .ZN(new_n696));
  OAI211_X1 g271(.A(new_n695), .B(new_n696), .C1(G301), .C2(new_n673), .ZN(new_n697));
  XNOR2_X1  g272(.A(new_n697), .B(G1961), .ZN(new_n698));
  INV_X1    g273(.A(G34), .ZN(new_n699));
  AND2_X1   g274(.A1(new_n699), .A2(KEYINPUT24), .ZN(new_n700));
  NOR2_X1   g275(.A1(new_n699), .A2(KEYINPUT24), .ZN(new_n701));
  OAI21_X1  g276(.A(new_n678), .B1(new_n700), .B2(new_n701), .ZN(new_n702));
  OAI21_X1  g277(.A(new_n702), .B1(G160), .B2(new_n678), .ZN(new_n703));
  XOR2_X1   g278(.A(KEYINPUT93), .B(G2084), .Z(new_n704));
  XNOR2_X1  g279(.A(new_n703), .B(new_n704), .ZN(new_n705));
  NAND2_X1  g280(.A1(new_n678), .A2(G33), .ZN(new_n706));
  XNOR2_X1  g281(.A(KEYINPUT92), .B(KEYINPUT25), .ZN(new_n707));
  NAND3_X1  g282(.A1(new_n482), .A2(G103), .A3(G2104), .ZN(new_n708));
  XNOR2_X1  g283(.A(new_n707), .B(new_n708), .ZN(new_n709));
  AOI22_X1  g284(.A1(new_n499), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n710));
  NOR2_X1   g285(.A1(new_n710), .A2(new_n482), .ZN(new_n711));
  AOI211_X1 g286(.A(new_n709), .B(new_n711), .C1(G139), .C2(new_n478), .ZN(new_n712));
  OAI21_X1  g287(.A(new_n706), .B1(new_n712), .B2(new_n678), .ZN(new_n713));
  NAND2_X1  g288(.A1(new_n713), .A2(G2072), .ZN(new_n714));
  INV_X1    g289(.A(KEYINPUT30), .ZN(new_n715));
  AND2_X1   g290(.A1(new_n715), .A2(G28), .ZN(new_n716));
  OAI21_X1  g291(.A(new_n678), .B1(new_n715), .B2(G28), .ZN(new_n717));
  AND2_X1   g292(.A1(KEYINPUT31), .A2(G11), .ZN(new_n718));
  NOR2_X1   g293(.A1(KEYINPUT31), .A2(G11), .ZN(new_n719));
  OAI22_X1  g294(.A1(new_n716), .A2(new_n717), .B1(new_n718), .B2(new_n719), .ZN(new_n720));
  INV_X1    g295(.A(new_n619), .ZN(new_n721));
  AOI21_X1  g296(.A(new_n720), .B1(new_n721), .B2(G29), .ZN(new_n722));
  NAND4_X1  g297(.A1(new_n698), .A2(new_n705), .A3(new_n714), .A4(new_n722), .ZN(new_n723));
  NAND2_X1  g298(.A1(new_n692), .A2(new_n690), .ZN(new_n724));
  NAND2_X1  g299(.A1(new_n673), .A2(G21), .ZN(new_n725));
  OAI21_X1  g300(.A(new_n725), .B1(G168), .B2(new_n673), .ZN(new_n726));
  INV_X1    g301(.A(G1966), .ZN(new_n727));
  XNOR2_X1  g302(.A(new_n726), .B(new_n727), .ZN(new_n728));
  OAI211_X1 g303(.A(new_n724), .B(new_n728), .C1(G2072), .C2(new_n713), .ZN(new_n729));
  NOR3_X1   g304(.A1(new_n693), .A2(new_n723), .A3(new_n729), .ZN(new_n730));
  NAND2_X1  g305(.A1(new_n678), .A2(G35), .ZN(new_n731));
  XOR2_X1   g306(.A(new_n731), .B(KEYINPUT96), .Z(new_n732));
  OAI21_X1  g307(.A(new_n732), .B1(G162), .B2(new_n678), .ZN(new_n733));
  XOR2_X1   g308(.A(new_n733), .B(KEYINPUT29), .Z(new_n734));
  INV_X1    g309(.A(G2090), .ZN(new_n735));
  NOR2_X1   g310(.A1(new_n734), .A2(new_n735), .ZN(new_n736));
  XOR2_X1   g311(.A(new_n736), .B(KEYINPUT97), .Z(new_n737));
  NAND2_X1  g312(.A1(new_n678), .A2(G32), .ZN(new_n738));
  NAND2_X1  g313(.A1(new_n487), .A2(G129), .ZN(new_n739));
  NAND3_X1  g314(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n740));
  INV_X1    g315(.A(KEYINPUT26), .ZN(new_n741));
  OR2_X1    g316(.A1(new_n740), .A2(new_n741), .ZN(new_n742));
  NAND2_X1  g317(.A1(new_n740), .A2(new_n741), .ZN(new_n743));
  AOI22_X1  g318(.A1(new_n742), .A2(new_n743), .B1(G105), .B2(new_n463), .ZN(new_n744));
  NAND2_X1  g319(.A1(new_n478), .A2(G141), .ZN(new_n745));
  AND2_X1   g320(.A1(new_n744), .A2(new_n745), .ZN(new_n746));
  AND2_X1   g321(.A1(new_n739), .A2(new_n746), .ZN(new_n747));
  XNOR2_X1  g322(.A(new_n747), .B(KEYINPUT94), .ZN(new_n748));
  OAI21_X1  g323(.A(new_n738), .B1(new_n748), .B2(new_n678), .ZN(new_n749));
  XOR2_X1   g324(.A(KEYINPUT27), .B(G1996), .Z(new_n750));
  XNOR2_X1  g325(.A(new_n749), .B(new_n750), .ZN(new_n751));
  AOI21_X1  g326(.A(new_n751), .B1(new_n735), .B2(new_n734), .ZN(new_n752));
  NAND3_X1  g327(.A1(new_n730), .A2(new_n737), .A3(new_n752), .ZN(new_n753));
  NAND2_X1  g328(.A1(new_n673), .A2(G19), .ZN(new_n754));
  OAI21_X1  g329(.A(new_n754), .B1(new_n545), .B2(new_n673), .ZN(new_n755));
  NOR2_X1   g330(.A1(new_n755), .A2(G1341), .ZN(new_n756));
  NOR2_X1   g331(.A1(G4), .A2(G16), .ZN(new_n757));
  AOI21_X1  g332(.A(new_n757), .B1(new_n596), .B2(G16), .ZN(new_n758));
  XNOR2_X1  g333(.A(new_n758), .B(G1348), .ZN(new_n759));
  AND2_X1   g334(.A1(new_n755), .A2(G1341), .ZN(new_n760));
  NOR4_X1   g335(.A1(new_n753), .A2(new_n756), .A3(new_n759), .A4(new_n760), .ZN(new_n761));
  NAND2_X1  g336(.A1(new_n673), .A2(G23), .ZN(new_n762));
  INV_X1    g337(.A(G288), .ZN(new_n763));
  OAI21_X1  g338(.A(new_n762), .B1(new_n763), .B2(new_n673), .ZN(new_n764));
  XNOR2_X1  g339(.A(KEYINPUT33), .B(G1976), .ZN(new_n765));
  XNOR2_X1  g340(.A(new_n764), .B(new_n765), .ZN(new_n766));
  NAND2_X1  g341(.A1(new_n673), .A2(G22), .ZN(new_n767));
  OAI21_X1  g342(.A(new_n767), .B1(G166), .B2(new_n673), .ZN(new_n768));
  INV_X1    g343(.A(G1971), .ZN(new_n769));
  XNOR2_X1  g344(.A(new_n768), .B(new_n769), .ZN(new_n770));
  NOR2_X1   g345(.A1(G6), .A2(G16), .ZN(new_n771));
  INV_X1    g346(.A(G305), .ZN(new_n772));
  AOI21_X1  g347(.A(new_n771), .B1(new_n772), .B2(G16), .ZN(new_n773));
  XOR2_X1   g348(.A(KEYINPUT32), .B(G1981), .Z(new_n774));
  XNOR2_X1  g349(.A(new_n773), .B(new_n774), .ZN(new_n775));
  NAND3_X1  g350(.A1(new_n766), .A2(new_n770), .A3(new_n775), .ZN(new_n776));
  XOR2_X1   g351(.A(new_n776), .B(KEYINPUT34), .Z(new_n777));
  AOI21_X1  g352(.A(new_n673), .B1(G290), .B2(KEYINPUT90), .ZN(new_n778));
  OAI21_X1  g353(.A(new_n778), .B1(KEYINPUT90), .B2(G290), .ZN(new_n779));
  INV_X1    g354(.A(G24), .ZN(new_n780));
  OAI21_X1  g355(.A(new_n779), .B1(G16), .B2(new_n780), .ZN(new_n781));
  NAND2_X1  g356(.A1(new_n781), .A2(G1986), .ZN(new_n782));
  OR2_X1    g357(.A1(new_n781), .A2(G1986), .ZN(new_n783));
  NAND2_X1  g358(.A1(new_n678), .A2(G25), .ZN(new_n784));
  AND2_X1   g359(.A1(new_n478), .A2(G131), .ZN(new_n785));
  OAI21_X1  g360(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n786));
  INV_X1    g361(.A(G107), .ZN(new_n787));
  AOI21_X1  g362(.A(new_n786), .B1(new_n787), .B2(G2105), .ZN(new_n788));
  AOI211_X1 g363(.A(new_n785), .B(new_n788), .C1(new_n487), .C2(G119), .ZN(new_n789));
  OAI21_X1  g364(.A(new_n784), .B1(new_n789), .B2(new_n678), .ZN(new_n790));
  XOR2_X1   g365(.A(KEYINPUT35), .B(G1991), .Z(new_n791));
  XOR2_X1   g366(.A(new_n790), .B(new_n791), .Z(new_n792));
  XNOR2_X1  g367(.A(new_n792), .B(KEYINPUT89), .ZN(new_n793));
  NAND4_X1  g368(.A1(new_n777), .A2(new_n782), .A3(new_n783), .A4(new_n793), .ZN(new_n794));
  XNOR2_X1  g369(.A(new_n794), .B(KEYINPUT36), .ZN(new_n795));
  NAND2_X1  g370(.A1(new_n761), .A2(new_n795), .ZN(new_n796));
  INV_X1    g371(.A(new_n796), .ZN(G311));
  XOR2_X1   g372(.A(new_n796), .B(KEYINPUT98), .Z(G150));
  AOI22_X1  g373(.A1(G55), .A2(new_n538), .B1(new_n516), .B2(G93), .ZN(new_n799));
  NAND2_X1  g374(.A1(new_n515), .A2(G67), .ZN(new_n800));
  NAND2_X1  g375(.A1(G80), .A2(G543), .ZN(new_n801));
  AOI21_X1  g376(.A(new_n522), .B1(new_n800), .B2(new_n801), .ZN(new_n802));
  OAI21_X1  g377(.A(new_n799), .B1(KEYINPUT99), .B2(new_n802), .ZN(new_n803));
  AND2_X1   g378(.A1(new_n802), .A2(KEYINPUT99), .ZN(new_n804));
  NOR2_X1   g379(.A1(new_n803), .A2(new_n804), .ZN(new_n805));
  INV_X1    g380(.A(G860), .ZN(new_n806));
  NOR2_X1   g381(.A1(new_n805), .A2(new_n806), .ZN(new_n807));
  XNOR2_X1  g382(.A(new_n807), .B(KEYINPUT37), .ZN(new_n808));
  NOR2_X1   g383(.A1(new_n545), .A2(new_n805), .ZN(new_n809));
  NOR3_X1   g384(.A1(new_n803), .A2(new_n544), .A3(new_n804), .ZN(new_n810));
  NOR2_X1   g385(.A1(new_n809), .A2(new_n810), .ZN(new_n811));
  XNOR2_X1  g386(.A(new_n811), .B(KEYINPUT38), .ZN(new_n812));
  NAND2_X1  g387(.A1(new_n596), .A2(G559), .ZN(new_n813));
  XNOR2_X1  g388(.A(new_n812), .B(new_n813), .ZN(new_n814));
  NAND2_X1  g389(.A1(new_n814), .A2(KEYINPUT39), .ZN(new_n815));
  XOR2_X1   g390(.A(new_n815), .B(KEYINPUT100), .Z(new_n816));
  OAI21_X1  g391(.A(new_n806), .B1(new_n814), .B2(KEYINPUT39), .ZN(new_n817));
  OAI21_X1  g392(.A(new_n808), .B1(new_n816), .B2(new_n817), .ZN(G145));
  XNOR2_X1  g393(.A(new_n686), .B(G164), .ZN(new_n819));
  NAND2_X1  g394(.A1(new_n478), .A2(G142), .ZN(new_n820));
  NOR2_X1   g395(.A1(new_n482), .A2(G118), .ZN(new_n821));
  OAI21_X1  g396(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n822));
  OAI21_X1  g397(.A(new_n820), .B1(new_n821), .B2(new_n822), .ZN(new_n823));
  AOI21_X1  g398(.A(new_n823), .B1(new_n487), .B2(G130), .ZN(new_n824));
  XNOR2_X1  g399(.A(new_n819), .B(new_n824), .ZN(new_n825));
  XOR2_X1   g400(.A(new_n789), .B(new_n611), .Z(new_n826));
  XNOR2_X1  g401(.A(new_n825), .B(new_n826), .ZN(new_n827));
  INV_X1    g402(.A(new_n748), .ZN(new_n828));
  NAND2_X1  g403(.A1(new_n828), .A2(new_n712), .ZN(new_n829));
  INV_X1    g404(.A(new_n747), .ZN(new_n830));
  OAI21_X1  g405(.A(new_n829), .B1(new_n830), .B2(new_n712), .ZN(new_n831));
  XNOR2_X1  g406(.A(new_n827), .B(new_n831), .ZN(new_n832));
  XNOR2_X1  g407(.A(new_n619), .B(G162), .ZN(new_n833));
  XNOR2_X1  g408(.A(new_n833), .B(G160), .ZN(new_n834));
  AOI21_X1  g409(.A(G37), .B1(new_n832), .B2(new_n834), .ZN(new_n835));
  OAI21_X1  g410(.A(new_n835), .B1(new_n834), .B2(new_n832), .ZN(new_n836));
  XNOR2_X1  g411(.A(new_n836), .B(KEYINPUT40), .ZN(G395));
  NOR2_X1   g412(.A1(new_n595), .A2(G559), .ZN(new_n838));
  XNOR2_X1  g413(.A(new_n811), .B(new_n838), .ZN(new_n839));
  NOR2_X1   g414(.A1(G299), .A2(new_n596), .ZN(new_n840));
  NOR2_X1   g415(.A1(new_n600), .A2(new_n595), .ZN(new_n841));
  NOR2_X1   g416(.A1(new_n840), .A2(new_n841), .ZN(new_n842));
  INV_X1    g417(.A(new_n842), .ZN(new_n843));
  NAND2_X1  g418(.A1(new_n839), .A2(new_n843), .ZN(new_n844));
  INV_X1    g419(.A(KEYINPUT41), .ZN(new_n845));
  OR2_X1    g420(.A1(new_n840), .A2(KEYINPUT101), .ZN(new_n846));
  NAND2_X1  g421(.A1(new_n840), .A2(KEYINPUT101), .ZN(new_n847));
  NAND2_X1  g422(.A1(new_n846), .A2(new_n847), .ZN(new_n848));
  OAI21_X1  g423(.A(new_n845), .B1(new_n848), .B2(new_n841), .ZN(new_n849));
  NOR2_X1   g424(.A1(new_n841), .A2(new_n845), .ZN(new_n850));
  OAI21_X1  g425(.A(new_n850), .B1(G299), .B2(new_n596), .ZN(new_n851));
  AND2_X1   g426(.A1(new_n849), .A2(new_n851), .ZN(new_n852));
  OAI21_X1  g427(.A(new_n844), .B1(new_n852), .B2(new_n839), .ZN(new_n853));
  OR2_X1    g428(.A1(new_n853), .A2(KEYINPUT42), .ZN(new_n854));
  XNOR2_X1  g429(.A(G166), .B(KEYINPUT102), .ZN(new_n855));
  XNOR2_X1  g430(.A(new_n855), .B(new_n585), .ZN(new_n856));
  XNOR2_X1  g431(.A(G288), .B(G305), .ZN(new_n857));
  XNOR2_X1  g432(.A(new_n856), .B(new_n857), .ZN(new_n858));
  NAND2_X1  g433(.A1(new_n853), .A2(KEYINPUT42), .ZN(new_n859));
  AND3_X1   g434(.A1(new_n854), .A2(new_n858), .A3(new_n859), .ZN(new_n860));
  AOI21_X1  g435(.A(new_n858), .B1(new_n854), .B2(new_n859), .ZN(new_n861));
  OAI21_X1  g436(.A(G868), .B1(new_n860), .B2(new_n861), .ZN(new_n862));
  OAI21_X1  g437(.A(new_n862), .B1(G868), .B2(new_n805), .ZN(G295));
  OAI21_X1  g438(.A(new_n862), .B1(G868), .B2(new_n805), .ZN(G331));
  XNOR2_X1  g439(.A(G171), .B(G168), .ZN(new_n865));
  OR3_X1    g440(.A1(new_n809), .A2(new_n810), .A3(new_n865), .ZN(new_n866));
  INV_X1    g441(.A(KEYINPUT103), .ZN(new_n867));
  OAI21_X1  g442(.A(new_n865), .B1(new_n809), .B2(new_n810), .ZN(new_n868));
  NAND3_X1  g443(.A1(new_n866), .A2(new_n867), .A3(new_n868), .ZN(new_n869));
  OR2_X1    g444(.A1(new_n868), .A2(new_n867), .ZN(new_n870));
  AOI21_X1  g445(.A(new_n842), .B1(new_n869), .B2(new_n870), .ZN(new_n871));
  INV_X1    g446(.A(KEYINPUT104), .ZN(new_n872));
  OR2_X1    g447(.A1(new_n871), .A2(new_n872), .ZN(new_n873));
  NAND2_X1  g448(.A1(new_n849), .A2(new_n851), .ZN(new_n874));
  NAND2_X1  g449(.A1(new_n866), .A2(new_n868), .ZN(new_n875));
  NAND2_X1  g450(.A1(new_n874), .A2(new_n875), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n871), .A2(new_n872), .ZN(new_n877));
  NAND3_X1  g452(.A1(new_n873), .A2(new_n876), .A3(new_n877), .ZN(new_n878));
  INV_X1    g453(.A(new_n858), .ZN(new_n879));
  AOI21_X1  g454(.A(G37), .B1(new_n878), .B2(new_n879), .ZN(new_n880));
  NAND4_X1  g455(.A1(new_n873), .A2(new_n876), .A3(new_n858), .A4(new_n877), .ZN(new_n881));
  AOI21_X1  g456(.A(KEYINPUT43), .B1(new_n880), .B2(new_n881), .ZN(new_n882));
  AND2_X1   g457(.A1(new_n846), .A2(new_n847), .ZN(new_n883));
  AOI22_X1  g458(.A1(new_n883), .A2(new_n850), .B1(new_n845), .B2(new_n843), .ZN(new_n884));
  NAND2_X1  g459(.A1(new_n869), .A2(new_n870), .ZN(new_n885));
  OAI22_X1  g460(.A1(new_n884), .A2(new_n885), .B1(new_n842), .B2(new_n875), .ZN(new_n886));
  AOI21_X1  g461(.A(G37), .B1(new_n886), .B2(new_n879), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n887), .A2(new_n881), .ZN(new_n888));
  INV_X1    g463(.A(KEYINPUT43), .ZN(new_n889));
  NOR2_X1   g464(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  OAI21_X1  g465(.A(KEYINPUT44), .B1(new_n882), .B2(new_n890), .ZN(new_n891));
  AOI21_X1  g466(.A(new_n889), .B1(new_n880), .B2(new_n881), .ZN(new_n892));
  NOR2_X1   g467(.A1(new_n888), .A2(KEYINPUT43), .ZN(new_n893));
  NOR2_X1   g468(.A1(new_n892), .A2(new_n893), .ZN(new_n894));
  OAI21_X1  g469(.A(new_n891), .B1(new_n894), .B2(KEYINPUT44), .ZN(G397));
  AOI21_X1  g470(.A(G1384), .B1(new_n501), .B2(new_n505), .ZN(new_n896));
  NOR2_X1   g471(.A1(new_n896), .A2(KEYINPUT45), .ZN(new_n897));
  AND4_X1   g472(.A1(G40), .A2(new_n466), .A3(new_n474), .A4(new_n479), .ZN(new_n898));
  NAND2_X1  g473(.A1(new_n897), .A2(new_n898), .ZN(new_n899));
  INV_X1    g474(.A(new_n899), .ZN(new_n900));
  XNOR2_X1  g475(.A(new_n686), .B(G2067), .ZN(new_n901));
  INV_X1    g476(.A(new_n901), .ZN(new_n902));
  OAI21_X1  g477(.A(new_n900), .B1(new_n902), .B2(new_n830), .ZN(new_n903));
  NOR2_X1   g478(.A1(new_n899), .A2(G1996), .ZN(new_n904));
  INV_X1    g479(.A(new_n904), .ZN(new_n905));
  AND2_X1   g480(.A1(new_n905), .A2(KEYINPUT46), .ZN(new_n906));
  NOR2_X1   g481(.A1(new_n905), .A2(KEYINPUT46), .ZN(new_n907));
  OAI21_X1  g482(.A(new_n903), .B1(new_n906), .B2(new_n907), .ZN(new_n908));
  XNOR2_X1  g483(.A(new_n908), .B(KEYINPUT47), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n748), .A2(new_n904), .ZN(new_n910));
  AND2_X1   g485(.A1(new_n910), .A2(KEYINPUT105), .ZN(new_n911));
  NOR2_X1   g486(.A1(new_n910), .A2(KEYINPUT105), .ZN(new_n912));
  AOI21_X1  g487(.A(new_n902), .B1(G1996), .B2(new_n830), .ZN(new_n913));
  OAI22_X1  g488(.A1(new_n911), .A2(new_n912), .B1(new_n899), .B2(new_n913), .ZN(new_n914));
  XOR2_X1   g489(.A(new_n914), .B(KEYINPUT106), .Z(new_n915));
  XOR2_X1   g490(.A(new_n789), .B(new_n791), .Z(new_n916));
  OAI21_X1  g491(.A(new_n915), .B1(new_n899), .B2(new_n916), .ZN(new_n917));
  NOR3_X1   g492(.A1(new_n899), .A2(G290), .A3(G1986), .ZN(new_n918));
  XNOR2_X1  g493(.A(new_n918), .B(KEYINPUT48), .ZN(new_n919));
  OAI21_X1  g494(.A(new_n909), .B1(new_n917), .B2(new_n919), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n789), .A2(new_n791), .ZN(new_n921));
  XOR2_X1   g496(.A(new_n921), .B(KEYINPUT127), .Z(new_n922));
  NAND2_X1  g497(.A1(new_n915), .A2(new_n922), .ZN(new_n923));
  NAND2_X1  g498(.A1(new_n686), .A2(new_n688), .ZN(new_n924));
  AOI21_X1  g499(.A(new_n899), .B1(new_n923), .B2(new_n924), .ZN(new_n925));
  NOR2_X1   g500(.A1(new_n920), .A2(new_n925), .ZN(new_n926));
  INV_X1    g501(.A(KEYINPUT116), .ZN(new_n927));
  INV_X1    g502(.A(G8), .ZN(new_n928));
  NOR2_X1   g503(.A1(G166), .A2(new_n928), .ZN(new_n929));
  XNOR2_X1  g504(.A(KEYINPUT109), .B(KEYINPUT55), .ZN(new_n930));
  NAND2_X1  g505(.A1(new_n929), .A2(new_n930), .ZN(new_n931));
  NAND2_X1  g506(.A1(KEYINPUT109), .A2(KEYINPUT55), .ZN(new_n932));
  OAI21_X1  g507(.A(new_n932), .B1(G166), .B2(new_n928), .ZN(new_n933));
  NAND2_X1  g508(.A1(new_n931), .A2(new_n933), .ZN(new_n934));
  AOI21_X1  g509(.A(KEYINPUT107), .B1(new_n896), .B2(KEYINPUT45), .ZN(new_n935));
  OAI21_X1  g510(.A(new_n898), .B1(new_n935), .B2(new_n897), .ZN(new_n936));
  NOR3_X1   g511(.A1(new_n896), .A2(KEYINPUT107), .A3(KEYINPUT45), .ZN(new_n937));
  OAI21_X1  g512(.A(new_n769), .B1(new_n936), .B2(new_n937), .ZN(new_n938));
  NAND2_X1  g513(.A1(G160), .A2(G40), .ZN(new_n939));
  INV_X1    g514(.A(KEYINPUT50), .ZN(new_n940));
  AOI21_X1  g515(.A(new_n939), .B1(new_n896), .B2(new_n940), .ZN(new_n941));
  INV_X1    g516(.A(G1384), .ZN(new_n942));
  NAND2_X1  g517(.A1(new_n506), .A2(new_n942), .ZN(new_n943));
  NAND2_X1  g518(.A1(new_n943), .A2(KEYINPUT50), .ZN(new_n944));
  NAND3_X1  g519(.A1(new_n941), .A2(new_n735), .A3(new_n944), .ZN(new_n945));
  NAND2_X1  g520(.A1(new_n938), .A2(new_n945), .ZN(new_n946));
  INV_X1    g521(.A(KEYINPUT114), .ZN(new_n947));
  AOI21_X1  g522(.A(new_n928), .B1(new_n946), .B2(new_n947), .ZN(new_n948));
  INV_X1    g523(.A(new_n945), .ZN(new_n949));
  NAND2_X1  g524(.A1(new_n896), .A2(KEYINPUT45), .ZN(new_n950));
  INV_X1    g525(.A(KEYINPUT107), .ZN(new_n951));
  NAND2_X1  g526(.A1(new_n950), .A2(new_n951), .ZN(new_n952));
  INV_X1    g527(.A(KEYINPUT45), .ZN(new_n953));
  NAND2_X1  g528(.A1(new_n943), .A2(new_n953), .ZN(new_n954));
  NAND2_X1  g529(.A1(new_n952), .A2(new_n954), .ZN(new_n955));
  INV_X1    g530(.A(new_n937), .ZN(new_n956));
  NAND3_X1  g531(.A1(new_n955), .A2(new_n956), .A3(new_n898), .ZN(new_n957));
  AOI21_X1  g532(.A(new_n949), .B1(new_n957), .B2(new_n769), .ZN(new_n958));
  NAND2_X1  g533(.A1(new_n958), .A2(KEYINPUT114), .ZN(new_n959));
  AOI21_X1  g534(.A(new_n934), .B1(new_n948), .B2(new_n959), .ZN(new_n960));
  OAI21_X1  g535(.A(new_n898), .B1(new_n943), .B2(KEYINPUT50), .ZN(new_n961));
  OAI21_X1  g536(.A(KEYINPUT108), .B1(new_n896), .B2(new_n940), .ZN(new_n962));
  INV_X1    g537(.A(KEYINPUT108), .ZN(new_n963));
  NAND3_X1  g538(.A1(new_n943), .A2(new_n963), .A3(KEYINPUT50), .ZN(new_n964));
  AOI21_X1  g539(.A(new_n961), .B1(new_n962), .B2(new_n964), .ZN(new_n965));
  NAND2_X1  g540(.A1(new_n965), .A2(new_n735), .ZN(new_n966));
  NAND2_X1  g541(.A1(new_n966), .A2(new_n938), .ZN(new_n967));
  NAND3_X1  g542(.A1(new_n967), .A2(G8), .A3(new_n934), .ZN(new_n968));
  NAND2_X1  g543(.A1(new_n763), .A2(G1976), .ZN(new_n969));
  AOI21_X1  g544(.A(new_n928), .B1(new_n896), .B2(new_n898), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n969), .A2(new_n970), .ZN(new_n971));
  NAND2_X1  g546(.A1(new_n971), .A2(KEYINPUT52), .ZN(new_n972));
  INV_X1    g547(.A(KEYINPUT49), .ZN(new_n973));
  INV_X1    g548(.A(G1981), .ZN(new_n974));
  NAND4_X1  g549(.A1(new_n573), .A2(new_n574), .A3(new_n974), .A4(new_n575), .ZN(new_n975));
  INV_X1    g550(.A(KEYINPUT111), .ZN(new_n976));
  AOI21_X1  g551(.A(new_n973), .B1(new_n975), .B2(new_n976), .ZN(new_n977));
  INV_X1    g552(.A(new_n977), .ZN(new_n978));
  NAND3_X1  g553(.A1(new_n975), .A2(new_n976), .A3(new_n973), .ZN(new_n979));
  OAI211_X1 g554(.A(new_n978), .B(new_n979), .C1(new_n974), .C2(new_n772), .ZN(new_n980));
  INV_X1    g555(.A(new_n979), .ZN(new_n981));
  OAI211_X1 g556(.A(G1981), .B(G305), .C1(new_n981), .C2(new_n977), .ZN(new_n982));
  NAND3_X1  g557(.A1(new_n980), .A2(new_n982), .A3(new_n970), .ZN(new_n983));
  NAND2_X1  g558(.A1(new_n972), .A2(new_n983), .ZN(new_n984));
  INV_X1    g559(.A(G1976), .ZN(new_n985));
  AOI21_X1  g560(.A(KEYINPUT52), .B1(G288), .B2(new_n985), .ZN(new_n986));
  NAND3_X1  g561(.A1(new_n969), .A2(new_n970), .A3(new_n986), .ZN(new_n987));
  INV_X1    g562(.A(KEYINPUT110), .ZN(new_n988));
  NAND2_X1  g563(.A1(new_n987), .A2(new_n988), .ZN(new_n989));
  OR2_X1    g564(.A1(new_n987), .A2(new_n988), .ZN(new_n990));
  AOI21_X1  g565(.A(new_n984), .B1(new_n989), .B2(new_n990), .ZN(new_n991));
  NAND2_X1  g566(.A1(new_n968), .A2(new_n991), .ZN(new_n992));
  NAND3_X1  g567(.A1(new_n896), .A2(KEYINPUT115), .A3(KEYINPUT45), .ZN(new_n993));
  NAND3_X1  g568(.A1(new_n954), .A2(new_n898), .A3(new_n993), .ZN(new_n994));
  AOI21_X1  g569(.A(KEYINPUT115), .B1(new_n896), .B2(KEYINPUT45), .ZN(new_n995));
  OAI21_X1  g570(.A(new_n727), .B1(new_n994), .B2(new_n995), .ZN(new_n996));
  NAND2_X1  g571(.A1(new_n964), .A2(new_n962), .ZN(new_n997));
  INV_X1    g572(.A(G2084), .ZN(new_n998));
  NAND3_X1  g573(.A1(new_n997), .A2(new_n998), .A3(new_n941), .ZN(new_n999));
  AOI211_X1 g574(.A(new_n928), .B(G286), .C1(new_n996), .C2(new_n999), .ZN(new_n1000));
  INV_X1    g575(.A(new_n1000), .ZN(new_n1001));
  NOR3_X1   g576(.A1(new_n960), .A2(new_n992), .A3(new_n1001), .ZN(new_n1002));
  OAI21_X1  g577(.A(new_n927), .B1(new_n1002), .B2(KEYINPUT63), .ZN(new_n1003));
  INV_X1    g578(.A(new_n992), .ZN(new_n1004));
  INV_X1    g579(.A(new_n934), .ZN(new_n1005));
  OAI21_X1  g580(.A(G8), .B1(new_n958), .B2(KEYINPUT114), .ZN(new_n1006));
  NOR2_X1   g581(.A1(new_n946), .A2(new_n947), .ZN(new_n1007));
  OAI21_X1  g582(.A(new_n1005), .B1(new_n1006), .B2(new_n1007), .ZN(new_n1008));
  NAND3_X1  g583(.A1(new_n1004), .A2(new_n1008), .A3(new_n1000), .ZN(new_n1009));
  INV_X1    g584(.A(KEYINPUT63), .ZN(new_n1010));
  NAND3_X1  g585(.A1(new_n1009), .A2(KEYINPUT116), .A3(new_n1010), .ZN(new_n1011));
  NOR2_X1   g586(.A1(new_n1001), .A2(new_n1010), .ZN(new_n1012));
  AOI21_X1  g587(.A(new_n928), .B1(new_n966), .B2(new_n938), .ZN(new_n1013));
  OAI211_X1 g588(.A(new_n1004), .B(new_n1012), .C1(new_n1013), .C2(new_n934), .ZN(new_n1014));
  NAND3_X1  g589(.A1(new_n1003), .A2(new_n1011), .A3(new_n1014), .ZN(new_n1015));
  NAND3_X1  g590(.A1(new_n996), .A2(G168), .A3(new_n999), .ZN(new_n1016));
  NAND2_X1  g591(.A1(new_n1016), .A2(G8), .ZN(new_n1017));
  AOI21_X1  g592(.A(G168), .B1(new_n996), .B2(new_n999), .ZN(new_n1018));
  OAI21_X1  g593(.A(KEYINPUT51), .B1(new_n1017), .B2(new_n1018), .ZN(new_n1019));
  INV_X1    g594(.A(KEYINPUT62), .ZN(new_n1020));
  INV_X1    g595(.A(KEYINPUT51), .ZN(new_n1021));
  NAND3_X1  g596(.A1(new_n1016), .A2(new_n1021), .A3(G8), .ZN(new_n1022));
  AND3_X1   g597(.A1(new_n1019), .A2(new_n1020), .A3(new_n1022), .ZN(new_n1023));
  AOI21_X1  g598(.A(new_n1020), .B1(new_n1019), .B2(new_n1022), .ZN(new_n1024));
  NOR2_X1   g599(.A1(new_n1023), .A2(new_n1024), .ZN(new_n1025));
  INV_X1    g600(.A(KEYINPUT124), .ZN(new_n1026));
  NOR2_X1   g601(.A1(new_n897), .A2(new_n939), .ZN(new_n1027));
  INV_X1    g602(.A(new_n995), .ZN(new_n1028));
  INV_X1    g603(.A(KEYINPUT53), .ZN(new_n1029));
  NOR2_X1   g604(.A1(new_n1029), .A2(G2078), .ZN(new_n1030));
  NAND4_X1  g605(.A1(new_n1027), .A2(new_n1028), .A3(new_n993), .A4(new_n1030), .ZN(new_n1031));
  INV_X1    g606(.A(new_n1031), .ZN(new_n1032));
  AOI21_X1  g607(.A(G1961), .B1(new_n997), .B2(new_n941), .ZN(new_n1033));
  OAI21_X1  g608(.A(new_n1026), .B1(new_n1032), .B2(new_n1033), .ZN(new_n1034));
  NAND2_X1  g609(.A1(new_n997), .A2(new_n941), .ZN(new_n1035));
  INV_X1    g610(.A(G1961), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n1035), .A2(new_n1036), .ZN(new_n1037));
  NAND3_X1  g612(.A1(new_n1037), .A2(KEYINPUT124), .A3(new_n1031), .ZN(new_n1038));
  NAND2_X1  g613(.A1(new_n1034), .A2(new_n1038), .ZN(new_n1039));
  NOR2_X1   g614(.A1(new_n936), .A2(new_n937), .ZN(new_n1040));
  AOI21_X1  g615(.A(KEYINPUT53), .B1(new_n1040), .B2(new_n690), .ZN(new_n1041));
  INV_X1    g616(.A(new_n1041), .ZN(new_n1042));
  AOI21_X1  g617(.A(G301), .B1(new_n1039), .B2(new_n1042), .ZN(new_n1043));
  AND3_X1   g618(.A1(new_n1004), .A2(new_n1008), .A3(new_n1043), .ZN(new_n1044));
  NAND3_X1  g619(.A1(new_n983), .A2(new_n985), .A3(new_n763), .ZN(new_n1045));
  NAND2_X1  g620(.A1(new_n1045), .A2(new_n975), .ZN(new_n1046));
  INV_X1    g621(.A(KEYINPUT112), .ZN(new_n1047));
  NAND2_X1  g622(.A1(new_n1046), .A2(new_n1047), .ZN(new_n1048));
  NAND3_X1  g623(.A1(new_n1045), .A2(KEYINPUT112), .A3(new_n975), .ZN(new_n1049));
  NAND3_X1  g624(.A1(new_n1048), .A2(new_n970), .A3(new_n1049), .ZN(new_n1050));
  NAND3_X1  g625(.A1(new_n991), .A2(new_n1013), .A3(new_n934), .ZN(new_n1051));
  NAND2_X1  g626(.A1(new_n1050), .A2(new_n1051), .ZN(new_n1052));
  NAND2_X1  g627(.A1(new_n1052), .A2(KEYINPUT113), .ZN(new_n1053));
  INV_X1    g628(.A(KEYINPUT113), .ZN(new_n1054));
  NAND3_X1  g629(.A1(new_n1050), .A2(new_n1051), .A3(new_n1054), .ZN(new_n1055));
  AOI22_X1  g630(.A1(new_n1025), .A2(new_n1044), .B1(new_n1053), .B2(new_n1055), .ZN(new_n1056));
  AOI21_X1  g631(.A(KEYINPUT57), .B1(G299), .B2(KEYINPUT117), .ZN(new_n1057));
  INV_X1    g632(.A(KEYINPUT117), .ZN(new_n1058));
  INV_X1    g633(.A(KEYINPUT57), .ZN(new_n1059));
  NOR3_X1   g634(.A1(new_n600), .A2(new_n1058), .A3(new_n1059), .ZN(new_n1060));
  NOR2_X1   g635(.A1(new_n1057), .A2(new_n1060), .ZN(new_n1061));
  XNOR2_X1  g636(.A(KEYINPUT56), .B(G2072), .ZN(new_n1062));
  XOR2_X1   g637(.A(new_n1062), .B(KEYINPUT118), .Z(new_n1063));
  INV_X1    g638(.A(new_n1063), .ZN(new_n1064));
  NAND4_X1  g639(.A1(new_n955), .A2(new_n956), .A3(new_n898), .A4(new_n1064), .ZN(new_n1065));
  NAND2_X1  g640(.A1(new_n1065), .A2(KEYINPUT119), .ZN(new_n1066));
  NAND2_X1  g641(.A1(new_n941), .A2(new_n944), .ZN(new_n1067));
  INV_X1    g642(.A(G1956), .ZN(new_n1068));
  NAND2_X1  g643(.A1(new_n1067), .A2(new_n1068), .ZN(new_n1069));
  INV_X1    g644(.A(new_n936), .ZN(new_n1070));
  INV_X1    g645(.A(KEYINPUT119), .ZN(new_n1071));
  NAND4_X1  g646(.A1(new_n1070), .A2(new_n1071), .A3(new_n956), .A4(new_n1064), .ZN(new_n1072));
  AND4_X1   g647(.A1(new_n1061), .A2(new_n1066), .A3(new_n1069), .A4(new_n1072), .ZN(new_n1073));
  NAND2_X1  g648(.A1(new_n1072), .A2(new_n1069), .ZN(new_n1074));
  NOR3_X1   g649(.A1(new_n936), .A2(new_n937), .A3(new_n1063), .ZN(new_n1075));
  NOR2_X1   g650(.A1(new_n1075), .A2(new_n1071), .ZN(new_n1076));
  OAI22_X1  g651(.A1(new_n1074), .A2(new_n1076), .B1(new_n1057), .B2(new_n1060), .ZN(new_n1077));
  NAND2_X1  g652(.A1(new_n896), .A2(new_n898), .ZN(new_n1078));
  OAI22_X1  g653(.A1(new_n965), .A2(G1348), .B1(G2067), .B2(new_n1078), .ZN(new_n1079));
  NAND2_X1  g654(.A1(new_n1079), .A2(new_n596), .ZN(new_n1080));
  AOI21_X1  g655(.A(new_n1073), .B1(new_n1077), .B2(new_n1080), .ZN(new_n1081));
  INV_X1    g656(.A(KEYINPUT61), .ZN(new_n1082));
  AOI22_X1  g657(.A1(new_n1075), .A2(new_n1071), .B1(new_n1068), .B2(new_n1067), .ZN(new_n1083));
  AOI21_X1  g658(.A(new_n1061), .B1(new_n1083), .B2(new_n1066), .ZN(new_n1084));
  OAI21_X1  g659(.A(new_n1082), .B1(new_n1084), .B2(new_n1073), .ZN(new_n1085));
  INV_X1    g660(.A(KEYINPUT60), .ZN(new_n1086));
  AOI21_X1  g661(.A(new_n595), .B1(new_n1079), .B2(new_n1086), .ZN(new_n1087));
  INV_X1    g662(.A(KEYINPUT123), .ZN(new_n1088));
  NOR2_X1   g663(.A1(new_n1078), .A2(G2067), .ZN(new_n1089));
  INV_X1    g664(.A(G1348), .ZN(new_n1090));
  AOI21_X1  g665(.A(new_n1089), .B1(new_n1035), .B2(new_n1090), .ZN(new_n1091));
  AOI21_X1  g666(.A(new_n1088), .B1(new_n1091), .B2(KEYINPUT60), .ZN(new_n1092));
  AOI21_X1  g667(.A(G1348), .B1(new_n997), .B2(new_n941), .ZN(new_n1093));
  NOR4_X1   g668(.A1(new_n1093), .A2(KEYINPUT123), .A3(new_n1086), .A4(new_n1089), .ZN(new_n1094));
  OAI21_X1  g669(.A(new_n1087), .B1(new_n1092), .B2(new_n1094), .ZN(new_n1095));
  OAI21_X1  g670(.A(KEYINPUT123), .B1(new_n1079), .B2(new_n1086), .ZN(new_n1096));
  OAI21_X1  g671(.A(new_n596), .B1(new_n1091), .B2(KEYINPUT60), .ZN(new_n1097));
  NAND3_X1  g672(.A1(new_n1091), .A2(new_n1088), .A3(KEYINPUT60), .ZN(new_n1098));
  NAND3_X1  g673(.A1(new_n1096), .A2(new_n1097), .A3(new_n1098), .ZN(new_n1099));
  NAND2_X1  g674(.A1(new_n1095), .A2(new_n1099), .ZN(new_n1100));
  INV_X1    g675(.A(new_n545), .ZN(new_n1101));
  NOR2_X1   g676(.A1(new_n1101), .A2(KEYINPUT121), .ZN(new_n1102));
  NOR2_X1   g677(.A1(new_n957), .A2(G1996), .ZN(new_n1103));
  INV_X1    g678(.A(new_n1078), .ZN(new_n1104));
  XOR2_X1   g679(.A(KEYINPUT120), .B(KEYINPUT58), .Z(new_n1105));
  XNOR2_X1  g680(.A(new_n1105), .B(G1341), .ZN(new_n1106));
  NOR2_X1   g681(.A1(new_n1104), .A2(new_n1106), .ZN(new_n1107));
  OAI21_X1  g682(.A(new_n1102), .B1(new_n1103), .B2(new_n1107), .ZN(new_n1108));
  NAND2_X1  g683(.A1(new_n1108), .A2(KEYINPUT59), .ZN(new_n1109));
  INV_X1    g684(.A(KEYINPUT59), .ZN(new_n1110));
  OAI211_X1 g685(.A(new_n1110), .B(new_n1102), .C1(new_n1103), .C2(new_n1107), .ZN(new_n1111));
  NAND2_X1  g686(.A1(new_n1109), .A2(new_n1111), .ZN(new_n1112));
  AND3_X1   g687(.A1(new_n1085), .A2(new_n1100), .A3(new_n1112), .ZN(new_n1113));
  NAND3_X1  g688(.A1(new_n1083), .A2(new_n1061), .A3(new_n1066), .ZN(new_n1114));
  NAND3_X1  g689(.A1(new_n1077), .A2(new_n1114), .A3(KEYINPUT61), .ZN(new_n1115));
  NAND2_X1  g690(.A1(new_n1115), .A2(KEYINPUT122), .ZN(new_n1116));
  INV_X1    g691(.A(KEYINPUT122), .ZN(new_n1117));
  NAND4_X1  g692(.A1(new_n1077), .A2(new_n1114), .A3(new_n1117), .A4(KEYINPUT61), .ZN(new_n1118));
  NAND2_X1  g693(.A1(new_n1116), .A2(new_n1118), .ZN(new_n1119));
  AOI21_X1  g694(.A(new_n1081), .B1(new_n1113), .B2(new_n1119), .ZN(new_n1120));
  INV_X1    g695(.A(KEYINPUT125), .ZN(new_n1121));
  AOI211_X1 g696(.A(G171), .B(new_n1041), .C1(new_n1034), .C2(new_n1038), .ZN(new_n1122));
  NAND3_X1  g697(.A1(new_n1027), .A2(new_n950), .A3(new_n1030), .ZN(new_n1123));
  NAND2_X1  g698(.A1(new_n1037), .A2(new_n1123), .ZN(new_n1124));
  OAI21_X1  g699(.A(G171), .B1(new_n1124), .B2(new_n1041), .ZN(new_n1125));
  NAND2_X1  g700(.A1(new_n1125), .A2(KEYINPUT54), .ZN(new_n1126));
  OAI21_X1  g701(.A(new_n1121), .B1(new_n1122), .B2(new_n1126), .ZN(new_n1127));
  NAND3_X1  g702(.A1(new_n1039), .A2(G301), .A3(new_n1042), .ZN(new_n1128));
  NAND4_X1  g703(.A1(new_n1128), .A2(KEYINPUT125), .A3(KEYINPUT54), .A4(new_n1125), .ZN(new_n1129));
  NAND2_X1  g704(.A1(new_n1127), .A2(new_n1129), .ZN(new_n1130));
  NAND2_X1  g705(.A1(new_n1019), .A2(new_n1022), .ZN(new_n1131));
  AND3_X1   g706(.A1(new_n1131), .A2(new_n1008), .A3(new_n1004), .ZN(new_n1132));
  INV_X1    g707(.A(KEYINPUT54), .ZN(new_n1133));
  NOR3_X1   g708(.A1(new_n1124), .A2(new_n1041), .A3(G171), .ZN(new_n1134));
  OAI21_X1  g709(.A(new_n1133), .B1(new_n1043), .B2(new_n1134), .ZN(new_n1135));
  NAND3_X1  g710(.A1(new_n1130), .A2(new_n1132), .A3(new_n1135), .ZN(new_n1136));
  OAI211_X1 g711(.A(new_n1015), .B(new_n1056), .C1(new_n1120), .C2(new_n1136), .ZN(new_n1137));
  XOR2_X1   g712(.A(new_n585), .B(G1986), .Z(new_n1138));
  AOI21_X1  g713(.A(new_n917), .B1(new_n900), .B2(new_n1138), .ZN(new_n1139));
  AND3_X1   g714(.A1(new_n1137), .A2(KEYINPUT126), .A3(new_n1139), .ZN(new_n1140));
  AOI21_X1  g715(.A(KEYINPUT126), .B1(new_n1137), .B2(new_n1139), .ZN(new_n1141));
  OAI21_X1  g716(.A(new_n926), .B1(new_n1140), .B2(new_n1141), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g717(.A(G319), .ZN(new_n1144));
  NOR4_X1   g718(.A1(G229), .A2(G401), .A3(new_n1144), .A4(G227), .ZN(new_n1145));
  NAND2_X1  g719(.A1(new_n836), .A2(new_n1145), .ZN(new_n1146));
  NOR2_X1   g720(.A1(new_n894), .A2(new_n1146), .ZN(G308));
  OR2_X1    g721(.A1(new_n894), .A2(new_n1146), .ZN(G225));
endmodule


