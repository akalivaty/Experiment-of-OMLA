

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301,
         n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312,
         n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323,
         n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334,
         n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
         n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578;

  XNOR2_X1 U323 ( .A(n337), .B(KEYINPUT46), .ZN(n338) );
  XNOR2_X1 U324 ( .A(n339), .B(n338), .ZN(n377) );
  INV_X1 U325 ( .A(n343), .ZN(n330) );
  XNOR2_X1 U326 ( .A(n331), .B(n330), .ZN(n332) );
  XNOR2_X1 U327 ( .A(n333), .B(n332), .ZN(n334) );
  XOR2_X1 U328 ( .A(n322), .B(n321), .Z(n508) );
  XNOR2_X1 U329 ( .A(KEYINPUT118), .B(G169GAT), .ZN(n447) );
  XNOR2_X1 U330 ( .A(n448), .B(n447), .ZN(G1348GAT) );
  XOR2_X1 U331 ( .A(G29GAT), .B(G43GAT), .Z(n292) );
  XNOR2_X1 U332 ( .A(KEYINPUT8), .B(KEYINPUT7), .ZN(n291) );
  XNOR2_X1 U333 ( .A(n292), .B(n291), .ZN(n345) );
  XNOR2_X1 U334 ( .A(G50GAT), .B(G22GAT), .ZN(n293) );
  XNOR2_X1 U335 ( .A(n293), .B(G141GAT), .ZN(n415) );
  XNOR2_X1 U336 ( .A(n345), .B(n415), .ZN(n307) );
  XOR2_X1 U337 ( .A(G15GAT), .B(G1GAT), .Z(n358) );
  XNOR2_X1 U338 ( .A(G169GAT), .B(G36GAT), .ZN(n294) );
  XNOR2_X1 U339 ( .A(n294), .B(G8GAT), .ZN(n322) );
  XOR2_X1 U340 ( .A(n358), .B(n322), .Z(n296) );
  XNOR2_X1 U341 ( .A(G113GAT), .B(G197GAT), .ZN(n295) );
  XNOR2_X1 U342 ( .A(n296), .B(n295), .ZN(n300) );
  XOR2_X1 U343 ( .A(KEYINPUT71), .B(KEYINPUT70), .Z(n298) );
  NAND2_X1 U344 ( .A1(G229GAT), .A2(G233GAT), .ZN(n297) );
  XNOR2_X1 U345 ( .A(n298), .B(n297), .ZN(n299) );
  XOR2_X1 U346 ( .A(n300), .B(n299), .Z(n305) );
  XOR2_X1 U347 ( .A(KEYINPUT29), .B(KEYINPUT68), .Z(n302) );
  XNOR2_X1 U348 ( .A(KEYINPUT72), .B(KEYINPUT69), .ZN(n301) );
  XNOR2_X1 U349 ( .A(n302), .B(n301), .ZN(n303) );
  XNOR2_X1 U350 ( .A(n303), .B(KEYINPUT30), .ZN(n304) );
  XNOR2_X1 U351 ( .A(n305), .B(n304), .ZN(n306) );
  XNOR2_X1 U352 ( .A(n307), .B(n306), .ZN(n564) );
  XNOR2_X1 U353 ( .A(n564), .B(KEYINPUT73), .ZN(n518) );
  XOR2_X1 U354 ( .A(G190GAT), .B(KEYINPUT77), .Z(n344) );
  XOR2_X1 U355 ( .A(KEYINPUT93), .B(n344), .Z(n309) );
  NAND2_X1 U356 ( .A1(G226GAT), .A2(G233GAT), .ZN(n308) );
  XNOR2_X1 U357 ( .A(n309), .B(n308), .ZN(n314) );
  INV_X1 U358 ( .A(G204GAT), .ZN(n313) );
  XOR2_X1 U359 ( .A(G176GAT), .B(KEYINPUT76), .Z(n311) );
  XNOR2_X1 U360 ( .A(G92GAT), .B(G64GAT), .ZN(n310) );
  XNOR2_X1 U361 ( .A(n311), .B(n310), .ZN(n312) );
  XNOR2_X1 U362 ( .A(n313), .B(n312), .ZN(n326) );
  XOR2_X1 U363 ( .A(n314), .B(n326), .Z(n320) );
  XOR2_X1 U364 ( .A(G183GAT), .B(KEYINPUT18), .Z(n316) );
  XNOR2_X1 U365 ( .A(KEYINPUT19), .B(KEYINPUT17), .ZN(n315) );
  XNOR2_X1 U366 ( .A(n316), .B(n315), .ZN(n438) );
  XOR2_X1 U367 ( .A(G211GAT), .B(KEYINPUT21), .Z(n318) );
  XNOR2_X1 U368 ( .A(G197GAT), .B(G218GAT), .ZN(n317) );
  XNOR2_X1 U369 ( .A(n318), .B(n317), .ZN(n423) );
  XNOR2_X1 U370 ( .A(n438), .B(n423), .ZN(n319) );
  XNOR2_X1 U371 ( .A(n320), .B(n319), .ZN(n321) );
  INV_X1 U372 ( .A(n508), .ZN(n387) );
  XOR2_X1 U373 ( .A(KEYINPUT31), .B(KEYINPUT74), .Z(n324) );
  NAND2_X1 U374 ( .A1(G230GAT), .A2(G233GAT), .ZN(n323) );
  XNOR2_X1 U375 ( .A(n324), .B(n323), .ZN(n325) );
  XNOR2_X1 U376 ( .A(KEYINPUT75), .B(n325), .ZN(n335) );
  XOR2_X1 U377 ( .A(G57GAT), .B(KEYINPUT13), .Z(n357) );
  XOR2_X1 U378 ( .A(n357), .B(KEYINPUT33), .Z(n328) );
  XNOR2_X1 U379 ( .A(n326), .B(KEYINPUT32), .ZN(n327) );
  XNOR2_X1 U380 ( .A(n328), .B(n327), .ZN(n333) );
  XOR2_X1 U381 ( .A(G120GAT), .B(G71GAT), .Z(n434) );
  XNOR2_X1 U382 ( .A(G106GAT), .B(G78GAT), .ZN(n329) );
  XOR2_X1 U383 ( .A(n329), .B(G148GAT), .Z(n414) );
  XOR2_X1 U384 ( .A(n434), .B(n414), .Z(n331) );
  XOR2_X1 U385 ( .A(G99GAT), .B(G85GAT), .Z(n343) );
  XNOR2_X1 U386 ( .A(n335), .B(n334), .ZN(n381) );
  XOR2_X1 U387 ( .A(KEYINPUT64), .B(KEYINPUT41), .Z(n336) );
  XNOR2_X1 U388 ( .A(n381), .B(n336), .ZN(n540) );
  NOR2_X1 U389 ( .A1(n540), .A2(n564), .ZN(n339) );
  INV_X1 U390 ( .A(KEYINPUT108), .ZN(n337) );
  XOR2_X1 U391 ( .A(G92GAT), .B(G106GAT), .Z(n341) );
  XNOR2_X1 U392 ( .A(G50GAT), .B(G36GAT), .ZN(n340) );
  XNOR2_X1 U393 ( .A(n341), .B(n340), .ZN(n342) );
  XOR2_X1 U394 ( .A(n343), .B(n342), .Z(n347) );
  XNOR2_X1 U395 ( .A(n345), .B(n344), .ZN(n346) );
  XNOR2_X1 U396 ( .A(n347), .B(n346), .ZN(n351) );
  XOR2_X1 U397 ( .A(KEYINPUT66), .B(KEYINPUT10), .Z(n349) );
  NAND2_X1 U398 ( .A1(G232GAT), .A2(G233GAT), .ZN(n348) );
  XNOR2_X1 U399 ( .A(n349), .B(n348), .ZN(n350) );
  XOR2_X1 U400 ( .A(n351), .B(n350), .Z(n356) );
  XOR2_X1 U401 ( .A(KEYINPUT11), .B(G162GAT), .Z(n353) );
  XNOR2_X1 U402 ( .A(G134GAT), .B(G218GAT), .ZN(n352) );
  XNOR2_X1 U403 ( .A(n353), .B(n352), .ZN(n354) );
  XNOR2_X1 U404 ( .A(n354), .B(KEYINPUT9), .ZN(n355) );
  XOR2_X1 U405 ( .A(n356), .B(n355), .Z(n555) );
  XOR2_X1 U406 ( .A(n357), .B(G71GAT), .Z(n360) );
  XNOR2_X1 U407 ( .A(n358), .B(G127GAT), .ZN(n359) );
  XNOR2_X1 U408 ( .A(n360), .B(n359), .ZN(n364) );
  XOR2_X1 U409 ( .A(KEYINPUT78), .B(KEYINPUT14), .Z(n362) );
  XNOR2_X1 U410 ( .A(G8GAT), .B(KEYINPUT12), .ZN(n361) );
  XNOR2_X1 U411 ( .A(n362), .B(n361), .ZN(n363) );
  XOR2_X1 U412 ( .A(n364), .B(n363), .Z(n366) );
  XNOR2_X1 U413 ( .A(G22GAT), .B(G183GAT), .ZN(n365) );
  XNOR2_X1 U414 ( .A(n366), .B(n365), .ZN(n370) );
  XOR2_X1 U415 ( .A(KEYINPUT15), .B(KEYINPUT80), .Z(n368) );
  NAND2_X1 U416 ( .A1(G231GAT), .A2(G233GAT), .ZN(n367) );
  XNOR2_X1 U417 ( .A(n368), .B(n367), .ZN(n369) );
  XOR2_X1 U418 ( .A(n370), .B(n369), .Z(n375) );
  XOR2_X1 U419 ( .A(G64GAT), .B(G155GAT), .Z(n372) );
  XNOR2_X1 U420 ( .A(G78GAT), .B(G211GAT), .ZN(n371) );
  XNOR2_X1 U421 ( .A(n372), .B(n371), .ZN(n373) );
  XNOR2_X1 U422 ( .A(n373), .B(KEYINPUT79), .ZN(n374) );
  XOR2_X1 U423 ( .A(n375), .B(n374), .Z(n569) );
  INV_X1 U424 ( .A(n569), .ZN(n552) );
  NOR2_X1 U425 ( .A1(n555), .A2(n552), .ZN(n376) );
  NAND2_X1 U426 ( .A1(n377), .A2(n376), .ZN(n379) );
  XOR2_X1 U427 ( .A(KEYINPUT109), .B(KEYINPUT47), .Z(n378) );
  XNOR2_X1 U428 ( .A(n379), .B(n378), .ZN(n385) );
  XOR2_X1 U429 ( .A(n555), .B(KEYINPUT36), .Z(n575) );
  NOR2_X1 U430 ( .A1(n569), .A2(n575), .ZN(n380) );
  XNOR2_X1 U431 ( .A(KEYINPUT45), .B(n380), .ZN(n382) );
  NAND2_X1 U432 ( .A1(n382), .A2(n381), .ZN(n383) );
  NOR2_X1 U433 ( .A1(n518), .A2(n383), .ZN(n384) );
  NOR2_X1 U434 ( .A1(n385), .A2(n384), .ZN(n386) );
  XNOR2_X1 U435 ( .A(KEYINPUT48), .B(n386), .ZN(n533) );
  NOR2_X1 U436 ( .A1(n387), .A2(n533), .ZN(n388) );
  XNOR2_X1 U437 ( .A(n388), .B(KEYINPUT54), .ZN(n412) );
  XOR2_X1 U438 ( .A(KEYINPUT90), .B(KEYINPUT91), .Z(n390) );
  XNOR2_X1 U439 ( .A(G1GAT), .B(KEYINPUT92), .ZN(n389) );
  XNOR2_X1 U440 ( .A(n390), .B(n389), .ZN(n399) );
  XOR2_X1 U441 ( .A(KEYINPUT1), .B(KEYINPUT4), .Z(n397) );
  XOR2_X1 U442 ( .A(KEYINPUT82), .B(G134GAT), .Z(n392) );
  XNOR2_X1 U443 ( .A(KEYINPUT0), .B(G127GAT), .ZN(n391) );
  XNOR2_X1 U444 ( .A(n392), .B(n391), .ZN(n393) );
  XNOR2_X1 U445 ( .A(G113GAT), .B(n393), .ZN(n443) );
  XOR2_X1 U446 ( .A(G155GAT), .B(KEYINPUT2), .Z(n395) );
  XNOR2_X1 U447 ( .A(G162GAT), .B(KEYINPUT3), .ZN(n394) );
  XNOR2_X1 U448 ( .A(n395), .B(n394), .ZN(n422) );
  XOR2_X1 U449 ( .A(n443), .B(n422), .Z(n396) );
  XNOR2_X1 U450 ( .A(n397), .B(n396), .ZN(n398) );
  XNOR2_X1 U451 ( .A(n399), .B(n398), .ZN(n411) );
  NAND2_X1 U452 ( .A1(G225GAT), .A2(G233GAT), .ZN(n405) );
  XOR2_X1 U453 ( .A(KEYINPUT6), .B(G148GAT), .Z(n401) );
  XNOR2_X1 U454 ( .A(G141GAT), .B(G120GAT), .ZN(n400) );
  XNOR2_X1 U455 ( .A(n401), .B(n400), .ZN(n403) );
  XOR2_X1 U456 ( .A(G29GAT), .B(G85GAT), .Z(n402) );
  XNOR2_X1 U457 ( .A(n403), .B(n402), .ZN(n404) );
  XNOR2_X1 U458 ( .A(n405), .B(n404), .ZN(n409) );
  XOR2_X1 U459 ( .A(G57GAT), .B(KEYINPUT89), .Z(n407) );
  XNOR2_X1 U460 ( .A(KEYINPUT88), .B(KEYINPUT5), .ZN(n406) );
  XNOR2_X1 U461 ( .A(n407), .B(n406), .ZN(n408) );
  XNOR2_X1 U462 ( .A(n409), .B(n408), .ZN(n410) );
  XOR2_X1 U463 ( .A(n411), .B(n410), .Z(n469) );
  AND2_X1 U464 ( .A1(n412), .A2(n469), .ZN(n413) );
  XOR2_X1 U465 ( .A(KEYINPUT65), .B(n413), .Z(n563) );
  XNOR2_X1 U466 ( .A(n415), .B(n414), .ZN(n427) );
  XOR2_X1 U467 ( .A(KEYINPUT22), .B(KEYINPUT86), .Z(n417) );
  XNOR2_X1 U468 ( .A(KEYINPUT23), .B(KEYINPUT24), .ZN(n416) );
  XNOR2_X1 U469 ( .A(n417), .B(n416), .ZN(n421) );
  XOR2_X1 U470 ( .A(G204GAT), .B(KEYINPUT87), .Z(n419) );
  NAND2_X1 U471 ( .A1(G228GAT), .A2(G233GAT), .ZN(n418) );
  XNOR2_X1 U472 ( .A(n419), .B(n418), .ZN(n420) );
  XOR2_X1 U473 ( .A(n421), .B(n420), .Z(n425) );
  XNOR2_X1 U474 ( .A(n423), .B(n422), .ZN(n424) );
  XNOR2_X1 U475 ( .A(n425), .B(n424), .ZN(n426) );
  XNOR2_X1 U476 ( .A(n427), .B(n426), .ZN(n461) );
  NAND2_X1 U477 ( .A1(n563), .A2(n461), .ZN(n428) );
  XNOR2_X1 U478 ( .A(n428), .B(KEYINPUT55), .ZN(n445) );
  XOR2_X1 U479 ( .A(KEYINPUT85), .B(KEYINPUT20), .Z(n430) );
  XNOR2_X1 U480 ( .A(G15GAT), .B(KEYINPUT83), .ZN(n429) );
  XNOR2_X1 U481 ( .A(n430), .B(n429), .ZN(n442) );
  XOR2_X1 U482 ( .A(KEYINPUT84), .B(G99GAT), .Z(n432) );
  XNOR2_X1 U483 ( .A(G43GAT), .B(G190GAT), .ZN(n431) );
  XNOR2_X1 U484 ( .A(n432), .B(n431), .ZN(n433) );
  XOR2_X1 U485 ( .A(n434), .B(n433), .Z(n436) );
  NAND2_X1 U486 ( .A1(G227GAT), .A2(G233GAT), .ZN(n435) );
  XNOR2_X1 U487 ( .A(n436), .B(n435), .ZN(n437) );
  XOR2_X1 U488 ( .A(n437), .B(G176GAT), .Z(n440) );
  XNOR2_X1 U489 ( .A(G169GAT), .B(n438), .ZN(n439) );
  XNOR2_X1 U490 ( .A(n440), .B(n439), .ZN(n441) );
  XNOR2_X1 U491 ( .A(n442), .B(n441), .ZN(n444) );
  XNOR2_X1 U492 ( .A(n444), .B(n443), .ZN(n515) );
  NAND2_X1 U493 ( .A1(n445), .A2(n515), .ZN(n446) );
  XNOR2_X2 U494 ( .A(n446), .B(KEYINPUT117), .ZN(n556) );
  NAND2_X1 U495 ( .A1(n518), .A2(n556), .ZN(n448) );
  NAND2_X1 U496 ( .A1(n381), .A2(n518), .ZN(n481) );
  INV_X1 U497 ( .A(n555), .ZN(n545) );
  NAND2_X1 U498 ( .A1(n552), .A2(n545), .ZN(n449) );
  XNOR2_X1 U499 ( .A(n449), .B(KEYINPUT81), .ZN(n450) );
  XNOR2_X1 U500 ( .A(n450), .B(KEYINPUT16), .ZN(n468) );
  XNOR2_X1 U501 ( .A(KEYINPUT27), .B(KEYINPUT94), .ZN(n451) );
  XOR2_X1 U502 ( .A(n451), .B(n508), .Z(n463) );
  INV_X1 U503 ( .A(n463), .ZN(n454) );
  NOR2_X1 U504 ( .A1(n515), .A2(n461), .ZN(n452) );
  XOR2_X1 U505 ( .A(KEYINPUT26), .B(n452), .Z(n453) );
  XNOR2_X1 U506 ( .A(KEYINPUT97), .B(n453), .ZN(n562) );
  NAND2_X1 U507 ( .A1(n454), .A2(n562), .ZN(n532) );
  NAND2_X1 U508 ( .A1(n515), .A2(n508), .ZN(n455) );
  NAND2_X1 U509 ( .A1(n455), .A2(n461), .ZN(n456) );
  XNOR2_X1 U510 ( .A(n456), .B(KEYINPUT98), .ZN(n457) );
  XOR2_X1 U511 ( .A(KEYINPUT25), .B(n457), .Z(n458) );
  NAND2_X1 U512 ( .A1(n532), .A2(n458), .ZN(n459) );
  NAND2_X1 U513 ( .A1(n459), .A2(n469), .ZN(n467) );
  XOR2_X1 U514 ( .A(KEYINPUT28), .B(KEYINPUT67), .Z(n460) );
  XOR2_X1 U515 ( .A(n461), .B(n460), .Z(n512) );
  OR2_X1 U516 ( .A1(n469), .A2(n512), .ZN(n462) );
  NOR2_X1 U517 ( .A1(n463), .A2(n462), .ZN(n516) );
  XNOR2_X1 U518 ( .A(KEYINPUT95), .B(n516), .ZN(n464) );
  NOR2_X1 U519 ( .A1(n515), .A2(n464), .ZN(n465) );
  XOR2_X1 U520 ( .A(KEYINPUT96), .B(n465), .Z(n466) );
  NAND2_X1 U521 ( .A1(n467), .A2(n466), .ZN(n478) );
  NAND2_X1 U522 ( .A1(n468), .A2(n478), .ZN(n495) );
  NOR2_X1 U523 ( .A1(n481), .A2(n495), .ZN(n476) );
  INV_X1 U524 ( .A(n469), .ZN(n535) );
  NAND2_X1 U525 ( .A1(n476), .A2(n535), .ZN(n470) );
  XNOR2_X1 U526 ( .A(n470), .B(KEYINPUT34), .ZN(n471) );
  XNOR2_X1 U527 ( .A(G1GAT), .B(n471), .ZN(G1324GAT) );
  NAND2_X1 U528 ( .A1(n476), .A2(n508), .ZN(n472) );
  XNOR2_X1 U529 ( .A(n472), .B(G8GAT), .ZN(G1325GAT) );
  XOR2_X1 U530 ( .A(KEYINPUT99), .B(KEYINPUT35), .Z(n474) );
  NAND2_X1 U531 ( .A1(n476), .A2(n515), .ZN(n473) );
  XNOR2_X1 U532 ( .A(n474), .B(n473), .ZN(n475) );
  XOR2_X1 U533 ( .A(G15GAT), .B(n475), .Z(G1326GAT) );
  NAND2_X1 U534 ( .A1(n512), .A2(n476), .ZN(n477) );
  XNOR2_X1 U535 ( .A(n477), .B(G22GAT), .ZN(G1327GAT) );
  XOR2_X1 U536 ( .A(KEYINPUT39), .B(KEYINPUT101), .Z(n485) );
  NAND2_X1 U537 ( .A1(n569), .A2(n478), .ZN(n479) );
  NOR2_X1 U538 ( .A1(n479), .A2(n575), .ZN(n480) );
  XNOR2_X1 U539 ( .A(n480), .B(KEYINPUT37), .ZN(n505) );
  NOR2_X1 U540 ( .A1(n505), .A2(n481), .ZN(n483) );
  XNOR2_X1 U541 ( .A(KEYINPUT38), .B(KEYINPUT100), .ZN(n482) );
  XNOR2_X1 U542 ( .A(n483), .B(n482), .ZN(n492) );
  NAND2_X1 U543 ( .A1(n492), .A2(n535), .ZN(n484) );
  XNOR2_X1 U544 ( .A(n485), .B(n484), .ZN(n486) );
  XOR2_X1 U545 ( .A(G29GAT), .B(n486), .Z(G1328GAT) );
  XOR2_X1 U546 ( .A(KEYINPUT102), .B(KEYINPUT103), .Z(n488) );
  NAND2_X1 U547 ( .A1(n492), .A2(n508), .ZN(n487) );
  XNOR2_X1 U548 ( .A(n488), .B(n487), .ZN(n489) );
  XNOR2_X1 U549 ( .A(G36GAT), .B(n489), .ZN(G1329GAT) );
  NAND2_X1 U550 ( .A1(n515), .A2(n492), .ZN(n490) );
  XNOR2_X1 U551 ( .A(n490), .B(KEYINPUT40), .ZN(n491) );
  XNOR2_X1 U552 ( .A(G43GAT), .B(n491), .ZN(G1330GAT) );
  NAND2_X1 U553 ( .A1(n512), .A2(n492), .ZN(n493) );
  XNOR2_X1 U554 ( .A(n493), .B(KEYINPUT104), .ZN(n494) );
  XNOR2_X1 U555 ( .A(G50GAT), .B(n494), .ZN(G1331GAT) );
  XNOR2_X1 U556 ( .A(G57GAT), .B(KEYINPUT42), .ZN(n497) );
  XNOR2_X1 U557 ( .A(KEYINPUT105), .B(n540), .ZN(n547) );
  NAND2_X1 U558 ( .A1(n564), .A2(n547), .ZN(n504) );
  NOR2_X1 U559 ( .A1(n504), .A2(n495), .ZN(n500) );
  NAND2_X1 U560 ( .A1(n535), .A2(n500), .ZN(n496) );
  XNOR2_X1 U561 ( .A(n497), .B(n496), .ZN(G1332GAT) );
  NAND2_X1 U562 ( .A1(n500), .A2(n508), .ZN(n498) );
  XNOR2_X1 U563 ( .A(n498), .B(G64GAT), .ZN(G1333GAT) );
  NAND2_X1 U564 ( .A1(n515), .A2(n500), .ZN(n499) );
  XNOR2_X1 U565 ( .A(n499), .B(G71GAT), .ZN(G1334GAT) );
  XOR2_X1 U566 ( .A(KEYINPUT106), .B(KEYINPUT43), .Z(n502) );
  NAND2_X1 U567 ( .A1(n500), .A2(n512), .ZN(n501) );
  XNOR2_X1 U568 ( .A(n502), .B(n501), .ZN(n503) );
  XNOR2_X1 U569 ( .A(G78GAT), .B(n503), .ZN(G1335GAT) );
  XOR2_X1 U570 ( .A(G85GAT), .B(KEYINPUT107), .Z(n507) );
  NOR2_X1 U571 ( .A1(n505), .A2(n504), .ZN(n511) );
  NAND2_X1 U572 ( .A1(n511), .A2(n535), .ZN(n506) );
  XNOR2_X1 U573 ( .A(n507), .B(n506), .ZN(G1336GAT) );
  NAND2_X1 U574 ( .A1(n511), .A2(n508), .ZN(n509) );
  XNOR2_X1 U575 ( .A(n509), .B(G92GAT), .ZN(G1337GAT) );
  NAND2_X1 U576 ( .A1(n515), .A2(n511), .ZN(n510) );
  XNOR2_X1 U577 ( .A(n510), .B(G99GAT), .ZN(G1338GAT) );
  NAND2_X1 U578 ( .A1(n512), .A2(n511), .ZN(n513) );
  XNOR2_X1 U579 ( .A(n513), .B(KEYINPUT44), .ZN(n514) );
  XNOR2_X1 U580 ( .A(G106GAT), .B(n514), .ZN(G1339GAT) );
  NAND2_X1 U581 ( .A1(n516), .A2(n515), .ZN(n517) );
  NOR2_X1 U582 ( .A1(n533), .A2(n517), .ZN(n529) );
  NAND2_X1 U583 ( .A1(n518), .A2(n529), .ZN(n519) );
  XNOR2_X1 U584 ( .A(n519), .B(KEYINPUT110), .ZN(n520) );
  XNOR2_X1 U585 ( .A(G113GAT), .B(n520), .ZN(G1340GAT) );
  XOR2_X1 U586 ( .A(KEYINPUT111), .B(KEYINPUT49), .Z(n522) );
  NAND2_X1 U587 ( .A1(n529), .A2(n547), .ZN(n521) );
  XNOR2_X1 U588 ( .A(n522), .B(n521), .ZN(n523) );
  XOR2_X1 U589 ( .A(G120GAT), .B(n523), .Z(G1341GAT) );
  NAND2_X1 U590 ( .A1(n529), .A2(n552), .ZN(n524) );
  XNOR2_X1 U591 ( .A(n524), .B(KEYINPUT50), .ZN(n525) );
  XNOR2_X1 U592 ( .A(G127GAT), .B(n525), .ZN(G1342GAT) );
  XOR2_X1 U593 ( .A(KEYINPUT113), .B(KEYINPUT114), .Z(n527) );
  XNOR2_X1 U594 ( .A(G134GAT), .B(KEYINPUT51), .ZN(n526) );
  XNOR2_X1 U595 ( .A(n527), .B(n526), .ZN(n528) );
  XOR2_X1 U596 ( .A(KEYINPUT112), .B(n528), .Z(n531) );
  NAND2_X1 U597 ( .A1(n529), .A2(n555), .ZN(n530) );
  XNOR2_X1 U598 ( .A(n531), .B(n530), .ZN(G1343GAT) );
  NOR2_X1 U599 ( .A1(n533), .A2(n532), .ZN(n534) );
  NAND2_X1 U600 ( .A1(n535), .A2(n534), .ZN(n544) );
  NOR2_X1 U601 ( .A1(n564), .A2(n544), .ZN(n537) );
  XNOR2_X1 U602 ( .A(G141GAT), .B(KEYINPUT115), .ZN(n536) );
  XNOR2_X1 U603 ( .A(n537), .B(n536), .ZN(G1344GAT) );
  XOR2_X1 U604 ( .A(KEYINPUT52), .B(KEYINPUT116), .Z(n539) );
  XNOR2_X1 U605 ( .A(G148GAT), .B(KEYINPUT53), .ZN(n538) );
  XNOR2_X1 U606 ( .A(n539), .B(n538), .ZN(n542) );
  NOR2_X1 U607 ( .A1(n540), .A2(n544), .ZN(n541) );
  XOR2_X1 U608 ( .A(n542), .B(n541), .Z(G1345GAT) );
  NOR2_X1 U609 ( .A1(n569), .A2(n544), .ZN(n543) );
  XOR2_X1 U610 ( .A(G155GAT), .B(n543), .Z(G1346GAT) );
  NOR2_X1 U611 ( .A1(n545), .A2(n544), .ZN(n546) );
  XOR2_X1 U612 ( .A(G162GAT), .B(n546), .Z(G1347GAT) );
  NAND2_X1 U613 ( .A1(n547), .A2(n556), .ZN(n549) );
  XOR2_X1 U614 ( .A(G176GAT), .B(KEYINPUT119), .Z(n548) );
  XNOR2_X1 U615 ( .A(n549), .B(n548), .ZN(n551) );
  XOR2_X1 U616 ( .A(KEYINPUT56), .B(KEYINPUT57), .Z(n550) );
  XNOR2_X1 U617 ( .A(n551), .B(n550), .ZN(G1349GAT) );
  NAND2_X1 U618 ( .A1(n556), .A2(n552), .ZN(n553) );
  XNOR2_X1 U619 ( .A(n553), .B(KEYINPUT120), .ZN(n554) );
  XNOR2_X1 U620 ( .A(G183GAT), .B(n554), .ZN(G1350GAT) );
  NAND2_X1 U621 ( .A1(n556), .A2(n555), .ZN(n558) );
  XOR2_X1 U622 ( .A(KEYINPUT121), .B(KEYINPUT58), .Z(n557) );
  XNOR2_X1 U623 ( .A(n558), .B(n557), .ZN(n559) );
  XNOR2_X1 U624 ( .A(n559), .B(G190GAT), .ZN(G1351GAT) );
  XOR2_X1 U625 ( .A(KEYINPUT122), .B(KEYINPUT59), .Z(n561) );
  XNOR2_X1 U626 ( .A(G197GAT), .B(KEYINPUT60), .ZN(n560) );
  XNOR2_X1 U627 ( .A(n561), .B(n560), .ZN(n566) );
  NAND2_X1 U628 ( .A1(n563), .A2(n562), .ZN(n574) );
  NOR2_X1 U629 ( .A1(n564), .A2(n574), .ZN(n565) );
  XOR2_X1 U630 ( .A(n566), .B(n565), .Z(G1352GAT) );
  NOR2_X1 U631 ( .A1(n381), .A2(n574), .ZN(n568) );
  XNOR2_X1 U632 ( .A(G204GAT), .B(KEYINPUT61), .ZN(n567) );
  XNOR2_X1 U633 ( .A(n568), .B(n567), .ZN(G1353GAT) );
  NOR2_X1 U634 ( .A1(n569), .A2(n574), .ZN(n571) );
  XNOR2_X1 U635 ( .A(G211GAT), .B(KEYINPUT123), .ZN(n570) );
  XNOR2_X1 U636 ( .A(n571), .B(n570), .ZN(G1354GAT) );
  XOR2_X1 U637 ( .A(KEYINPUT62), .B(KEYINPUT126), .Z(n573) );
  XNOR2_X1 U638 ( .A(G218GAT), .B(KEYINPUT125), .ZN(n572) );
  XNOR2_X1 U639 ( .A(n573), .B(n572), .ZN(n577) );
  NOR2_X1 U640 ( .A1(n575), .A2(n574), .ZN(n576) );
  XOR2_X1 U641 ( .A(n577), .B(n576), .Z(n578) );
  XNOR2_X1 U642 ( .A(KEYINPUT124), .B(n578), .ZN(G1355GAT) );
endmodule

