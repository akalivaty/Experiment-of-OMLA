

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, n371,
         n372, n373, n374, n375, n376, n377, n378, n379, n380, n381, n382,
         n383, n384, n385, n386, n387, n388, n389, n390, n391, n392, n393,
         n394, n395, n396, n397, n398, n399, n400, n401, n402, n403, n404,
         n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, n415,
         n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426,
         n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437,
         n438, n439, n440, n441, n442, n443, n444, n445, n446, n447, n448,
         n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, n459,
         n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, n470,
         n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481,
         n482, n483, n484, n485, n486, n487, n488, n489, n490, n491, n492,
         n493, n494, n495, n496, n497, n498, n499, n500, n501, n502, n503,
         n504, n505, n506, n507, n508, n509, n510, n511, n512, n513, n514,
         n515, n516, n517, n518, n519, n520, n521, n522, n523, n524, n525,
         n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536,
         n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547,
         n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558,
         n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569,
         n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580,
         n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591,
         n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602,
         n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, n613,
         n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624,
         n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635,
         n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, n646,
         n647, n648, n649, n650, n651, n652, n653, n654, n655, n656, n657,
         n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668,
         n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679,
         n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690,
         n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701,
         n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712,
         n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723,
         n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, n734,
         n735, n736, n737, n738, n739, n740, n741, n742, n743, n744, n745,
         n746, n747, n748, n749, n750, n751, n752, n753, n754, n755, n756,
         n757, n758, n759, n760, n761, n762, n763, n764, n765, n766, n767,
         n768, n769, n770, n771, n772, n773, n774, n775, n776, n777, n778,
         n779, n780, n781, n782, n783, n784, n785, n786, n787, n788, n789,
         n790, n791, n792, n793, n794, n795, n796, n797, n798, n799, n800,
         n801, n802, n803, n804;

  NOR2_X2 U383 ( .A1(G953), .A2(G237), .ZN(n541) );
  INV_X1 U384 ( .A(KEYINPUT8), .ZN(n451) );
  XNOR2_X1 U385 ( .A(n395), .B(n394), .ZN(n460) );
  XNOR2_X1 U386 ( .A(KEYINPUT100), .B(KEYINPUT99), .ZN(n445) );
  XOR2_X1 U387 ( .A(n696), .B(KEYINPUT88), .Z(n361) );
  XNOR2_X2 U388 ( .A(n609), .B(n608), .ZN(n803) );
  NAND2_X2 U389 ( .A1(n791), .A2(n778), .ZN(n691) );
  XNOR2_X2 U390 ( .A(n666), .B(KEYINPUT45), .ZN(n778) );
  XNOR2_X1 U391 ( .A(n607), .B(n606), .ZN(n640) );
  XNOR2_X1 U392 ( .A(n439), .B(n438), .ZN(n605) );
  INV_X2 U393 ( .A(G146), .ZN(n488) );
  NOR2_X2 U394 ( .A1(n648), .A2(n707), .ZN(n650) );
  INV_X2 U395 ( .A(KEYINPUT67), .ZN(n412) );
  NOR2_X1 U396 ( .A1(n611), .A2(n610), .ZN(n612) );
  BUF_X1 U397 ( .A(G146), .Z(n411) );
  AND2_X1 U398 ( .A1(n461), .A2(n463), .ZN(n363) );
  OR2_X1 U399 ( .A1(n656), .A2(n655), .ZN(n661) );
  NAND2_X1 U400 ( .A1(n640), .A2(n758), .ZN(n609) );
  OR2_X1 U401 ( .A1(n580), .A2(n578), .ZN(n653) );
  NOR2_X1 U402 ( .A1(n580), .A2(n579), .ZN(n581) );
  XNOR2_X1 U403 ( .A(n404), .B(KEYINPUT104), .ZN(n642) );
  NOR2_X1 U404 ( .A1(n768), .A2(G902), .ZN(n408) );
  INV_X1 U405 ( .A(KEYINPUT19), .ZN(n413) );
  XOR2_X1 U406 ( .A(G116), .B(KEYINPUT5), .Z(n499) );
  NAND2_X1 U407 ( .A1(n419), .A2(n417), .ZN(n734) );
  AND2_X1 U408 ( .A1(n421), .A2(n374), .ZN(n419) );
  NAND2_X1 U409 ( .A1(n695), .A2(n694), .ZN(n696) );
  XNOR2_X1 U410 ( .A(n693), .B(n692), .ZN(n695) );
  AND2_X1 U411 ( .A1(n386), .A2(n385), .ZN(n384) );
  AND2_X1 U412 ( .A1(n427), .A2(n426), .ZN(n425) );
  AND2_X1 U413 ( .A1(n392), .A2(n391), .ZN(n390) );
  NAND2_X1 U414 ( .A1(n661), .A2(KEYINPUT44), .ZN(n431) );
  XNOR2_X1 U415 ( .A(n581), .B(KEYINPUT32), .ZN(n656) );
  AND2_X1 U416 ( .A1(n638), .A2(n470), .ZN(n766) );
  XNOR2_X1 U417 ( .A(n616), .B(KEYINPUT42), .ZN(n802) );
  AND2_X2 U418 ( .A1(n619), .A2(n618), .ZN(n754) );
  XNOR2_X1 U419 ( .A(n408), .B(G478), .ZN(n588) );
  AND2_X1 U420 ( .A1(n381), .A2(n380), .ZN(n379) );
  XNOR2_X1 U421 ( .A(n499), .B(n500), .ZN(n403) );
  XNOR2_X1 U422 ( .A(G119), .B(KEYINPUT23), .ZN(n446) );
  XNOR2_X1 U423 ( .A(G902), .B(KEYINPUT15), .ZN(n521) );
  XNOR2_X1 U424 ( .A(G119), .B(G113), .ZN(n501) );
  NAND2_X1 U425 ( .A1(n428), .A2(n371), .ZN(n424) );
  BUF_X1 U426 ( .A(n592), .Z(n362) );
  XNOR2_X1 U427 ( .A(n497), .B(n496), .ZN(n584) );
  AND2_X1 U428 ( .A1(n550), .A2(G221), .ZN(n449) );
  NAND2_X1 U429 ( .A1(n461), .A2(n463), .ZN(n468) );
  NOR2_X1 U430 ( .A1(n574), .A2(n593), .ZN(n636) );
  XNOR2_X1 U431 ( .A(n484), .B(n483), .ZN(n585) );
  NOR2_X1 U432 ( .A1(n745), .A2(G902), .ZN(n484) );
  NAND2_X1 U433 ( .A1(n363), .A2(n383), .ZN(n382) );
  BUF_X1 U434 ( .A(n640), .Z(n364) );
  BUF_X1 U435 ( .A(n745), .Z(n365) );
  XNOR2_X1 U436 ( .A(n790), .B(n481), .ZN(n745) );
  NAND2_X1 U437 ( .A1(n410), .A2(n369), .ZN(n366) );
  NAND2_X1 U438 ( .A1(n366), .A2(n367), .ZN(n373) );
  OR2_X1 U439 ( .A1(n368), .A2(n759), .ZN(n367) );
  INV_X1 U440 ( .A(n634), .ZN(n368) );
  AND2_X1 U441 ( .A1(KEYINPUT84), .A2(n634), .ZN(n369) );
  INV_X1 U442 ( .A(n389), .ZN(n370) );
  XNOR2_X1 U443 ( .A(n696), .B(KEYINPUT88), .ZN(n423) );
  NAND2_X1 U444 ( .A1(n605), .A2(n698), .ZN(n607) );
  BUF_X1 U445 ( .A(n585), .Z(n614) );
  XNOR2_X2 U446 ( .A(n535), .B(n473), .ZN(n474) );
  INV_X1 U447 ( .A(KEYINPUT48), .ZN(n394) );
  NAND2_X1 U448 ( .A1(n384), .A2(n382), .ZN(n397) );
  INV_X1 U449 ( .A(G134), .ZN(n473) );
  INV_X1 U450 ( .A(n766), .ZN(n469) );
  INV_X1 U451 ( .A(KEYINPUT46), .ZN(n393) );
  NAND2_X1 U452 ( .A1(n802), .A2(n393), .ZN(n391) );
  NAND2_X1 U453 ( .A1(G237), .A2(G234), .ZN(n528) );
  NAND2_X1 U454 ( .A1(n378), .A2(n521), .ZN(n377) );
  NAND2_X1 U455 ( .A1(n456), .A2(n455), .ZN(n454) );
  INV_X1 U456 ( .A(KEYINPUT89), .ZN(n455) );
  INV_X1 U457 ( .A(n639), .ZN(n456) );
  AND2_X1 U458 ( .A1(n639), .A2(KEYINPUT89), .ZN(n458) );
  XNOR2_X1 U459 ( .A(G122), .B(G104), .ZN(n537) );
  XNOR2_X1 U460 ( .A(n635), .B(KEYINPUT38), .ZN(n698) );
  INV_X1 U461 ( .A(KEYINPUT79), .ZN(n441) );
  XNOR2_X1 U462 ( .A(n482), .B(G469), .ZN(n483) );
  XNOR2_X1 U463 ( .A(n565), .B(n375), .ZN(n566) );
  XNOR2_X1 U464 ( .A(n403), .B(n498), .ZN(n505) );
  OR2_X1 U465 ( .A1(n732), .A2(KEYINPUT119), .ZN(n420) );
  NOR2_X1 U466 ( .A1(n466), .A2(KEYINPUT69), .ZN(n383) );
  NOR2_X1 U467 ( .A1(n802), .A2(n393), .ZN(n388) );
  NOR2_X1 U468 ( .A1(n571), .A2(n570), .ZN(n586) );
  INV_X1 U469 ( .A(G237), .ZN(n522) );
  INV_X1 U470 ( .A(KEYINPUT10), .ZN(n489) );
  XNOR2_X1 U471 ( .A(n450), .B(n487), .ZN(n550) );
  XNOR2_X1 U472 ( .A(n451), .B(KEYINPUT66), .ZN(n450) );
  XOR2_X1 U473 ( .A(G113), .B(KEYINPUT11), .Z(n543) );
  XNOR2_X1 U474 ( .A(G140), .B(G143), .ZN(n538) );
  XNOR2_X1 U475 ( .A(KEYINPUT17), .B(KEYINPUT18), .ZN(n514) );
  NOR2_X1 U476 ( .A1(n435), .A2(n706), .ZN(n723) );
  INV_X1 U477 ( .A(n728), .ZN(n437) );
  OR2_X1 U478 ( .A1(n711), .A2(n594), .ZN(n595) );
  XNOR2_X1 U479 ( .A(KEYINPUT30), .B(KEYINPUT110), .ZN(n407) );
  NAND2_X1 U480 ( .A1(n525), .A2(n670), .ZN(n380) );
  INV_X1 U481 ( .A(G902), .ZN(n523) );
  XNOR2_X1 U482 ( .A(n717), .B(KEYINPUT6), .ZN(n593) );
  INV_X1 U483 ( .A(KEYINPUT72), .ZN(n502) );
  AND2_X1 U484 ( .A1(n804), .A2(n454), .ZN(n453) );
  XNOR2_X1 U485 ( .A(G140), .B(KEYINPUT68), .ZN(n475) );
  XNOR2_X1 U486 ( .A(n446), .B(n445), .ZN(n444) );
  XOR2_X1 U487 ( .A(G134), .B(G122), .Z(n552) );
  NAND2_X1 U488 ( .A1(n671), .A2(KEYINPUT2), .ZN(n694) );
  XNOR2_X1 U489 ( .A(n411), .B(G101), .ZN(n476) );
  XOR2_X1 U490 ( .A(G104), .B(G107), .Z(n477) );
  XNOR2_X1 U491 ( .A(n547), .B(G475), .ZN(n548) );
  NAND2_X1 U492 ( .A1(n624), .A2(n532), .ZN(n534) );
  NAND2_X1 U493 ( .A1(n566), .A2(n593), .ZN(n580) );
  XNOR2_X1 U494 ( .A(n676), .B(n678), .ZN(n679) );
  XNOR2_X1 U495 ( .A(n399), .B(n736), .ZN(n738) );
  INV_X1 U496 ( .A(KEYINPUT119), .ZN(n418) );
  INV_X1 U497 ( .A(n711), .ZN(n470) );
  XNOR2_X1 U498 ( .A(n637), .B(n409), .ZN(n638) );
  XNOR2_X1 U499 ( .A(KEYINPUT36), .B(KEYINPUT93), .ZN(n409) );
  AND2_X1 U500 ( .A1(n600), .A2(n590), .ZN(n591) );
  XNOR2_X1 U501 ( .A(n685), .B(KEYINPUT62), .ZN(n686) );
  NAND2_X1 U502 ( .A1(n361), .A2(n418), .ZN(n417) );
  AND2_X1 U503 ( .A1(n434), .A2(KEYINPUT92), .ZN(n371) );
  INV_X2 U504 ( .A(G953), .ZN(n793) );
  XOR2_X1 U505 ( .A(n587), .B(n407), .Z(n372) );
  AND2_X1 U506 ( .A1(n420), .A2(n793), .ZN(n374) );
  XOR2_X1 U507 ( .A(KEYINPUT64), .B(KEYINPUT22), .Z(n375) );
  NOR2_X2 U508 ( .A1(n635), .A2(n527), .ZN(n414) );
  NAND2_X2 U509 ( .A1(n379), .A2(n376), .ZN(n635) );
  OR2_X1 U510 ( .A1(n737), .A2(n377), .ZN(n376) );
  INV_X1 U511 ( .A(n525), .ZN(n378) );
  NAND2_X1 U512 ( .A1(n737), .A2(n525), .ZN(n381) );
  XNOR2_X1 U513 ( .A(n520), .B(n784), .ZN(n737) );
  NAND2_X1 U514 ( .A1(n466), .A2(KEYINPUT69), .ZN(n385) );
  NAND2_X1 U515 ( .A1(n468), .A2(KEYINPUT69), .ZN(n386) );
  NAND2_X1 U516 ( .A1(n390), .A2(n387), .ZN(n396) );
  NAND2_X1 U517 ( .A1(n389), .A2(n388), .ZN(n387) );
  INV_X1 U518 ( .A(n803), .ZN(n389) );
  NAND2_X1 U519 ( .A1(n803), .A2(n393), .ZN(n392) );
  NAND2_X1 U520 ( .A1(n397), .A2(n396), .ZN(n395) );
  BUF_X1 U521 ( .A(n619), .Z(n398) );
  BUF_X1 U522 ( .A(n737), .Z(n399) );
  INV_X1 U523 ( .A(n584), .ZN(n400) );
  INV_X1 U524 ( .A(n400), .ZN(n401) );
  BUF_X1 U525 ( .A(n790), .Z(n402) );
  NAND2_X1 U526 ( .A1(n658), .A2(n429), .ZN(n426) );
  NAND2_X1 U527 ( .A1(n592), .A2(n585), .ZN(n404) );
  XNOR2_X1 U528 ( .A(n491), .B(n405), .ZN(n772) );
  XNOR2_X1 U529 ( .A(n443), .B(n449), .ZN(n405) );
  XNOR2_X1 U530 ( .A(n406), .B(n518), .ZN(n520) );
  XNOR2_X1 U531 ( .A(n519), .B(n517), .ZN(n406) );
  XNOR2_X2 U532 ( .A(n414), .B(n413), .ZN(n624) );
  INV_X1 U533 ( .A(n434), .ZN(n430) );
  AND2_X2 U534 ( .A1(n675), .A2(n694), .ZN(n773) );
  NOR2_X2 U535 ( .A1(n619), .A2(n618), .ZN(n758) );
  NAND2_X1 U536 ( .A1(n465), .A2(KEYINPUT76), .ZN(n467) );
  XNOR2_X1 U537 ( .A(n507), .B(n506), .ZN(n685) );
  NAND2_X1 U538 ( .A1(n550), .A2(G217), .ZN(n551) );
  NAND2_X1 U539 ( .A1(n469), .A2(n467), .ZN(n466) );
  NAND2_X1 U540 ( .A1(n410), .A2(KEYINPUT84), .ZN(n631) );
  XNOR2_X1 U541 ( .A(n630), .B(KEYINPUT77), .ZN(n410) );
  XNOR2_X2 U542 ( .A(n549), .B(n548), .ZN(n619) );
  NOR2_X2 U543 ( .A1(n452), .A2(n459), .ZN(n791) );
  XNOR2_X2 U544 ( .A(n412), .B(G131), .ZN(n535) );
  NAND2_X1 U545 ( .A1(n415), .A2(n362), .ZN(n594) );
  INV_X1 U546 ( .A(n593), .ZN(n415) );
  XNOR2_X2 U547 ( .A(n416), .B(G472), .ZN(n717) );
  NAND2_X1 U548 ( .A1(n685), .A2(n523), .ZN(n416) );
  NAND2_X1 U549 ( .A1(n423), .A2(n422), .ZN(n421) );
  AND2_X1 U550 ( .A1(n732), .A2(KEYINPUT119), .ZN(n422) );
  AND2_X2 U551 ( .A1(n653), .A2(n654), .ZN(n434) );
  NAND2_X1 U552 ( .A1(n425), .A2(n424), .ZN(n432) );
  NAND2_X1 U553 ( .A1(n430), .A2(n433), .ZN(n427) );
  NAND2_X1 U554 ( .A1(n658), .A2(KEYINPUT44), .ZN(n428) );
  AND2_X1 U555 ( .A1(n433), .A2(KEYINPUT44), .ZN(n429) );
  NAND2_X1 U556 ( .A1(n432), .A2(n431), .ZN(n657) );
  INV_X1 U557 ( .A(KEYINPUT92), .ZN(n433) );
  NAND2_X1 U558 ( .A1(n436), .A2(n643), .ZN(n599) );
  INV_X1 U559 ( .A(n436), .ZN(n435) );
  AND2_X1 U560 ( .A1(n436), .A2(n437), .ZN(n729) );
  XNOR2_X2 U561 ( .A(n595), .B(KEYINPUT33), .ZN(n436) );
  XNOR2_X2 U562 ( .A(n553), .B(KEYINPUT4), .ZN(n519) );
  INV_X1 U563 ( .A(KEYINPUT78), .ZN(n438) );
  NAND2_X1 U564 ( .A1(n440), .A2(n372), .ZN(n439) );
  XNOR2_X1 U565 ( .A(n442), .B(n441), .ZN(n440) );
  NOR2_X2 U566 ( .A1(n642), .A2(n586), .ZN(n442) );
  XNOR2_X1 U567 ( .A(n447), .B(n444), .ZN(n443) );
  XNOR2_X1 U568 ( .A(n486), .B(n448), .ZN(n447) );
  XNOR2_X2 U569 ( .A(G128), .B(G110), .ZN(n448) );
  NAND2_X1 U570 ( .A1(n457), .A2(n453), .ZN(n452) );
  NAND2_X1 U571 ( .A1(n460), .A2(n458), .ZN(n457) );
  NOR2_X1 U572 ( .A1(n460), .A2(KEYINPUT89), .ZN(n459) );
  NAND2_X1 U573 ( .A1(n471), .A2(n462), .ZN(n461) );
  AND2_X1 U574 ( .A1(n633), .A2(n373), .ZN(n462) );
  NAND2_X1 U575 ( .A1(n464), .A2(KEYINPUT76), .ZN(n463) );
  INV_X1 U576 ( .A(n471), .ZN(n464) );
  NAND2_X1 U577 ( .A1(n633), .A2(n632), .ZN(n465) );
  XNOR2_X1 U578 ( .A(n617), .B(KEYINPUT86), .ZN(n471) );
  NOR2_X2 U579 ( .A1(n758), .A2(n754), .ZN(n620) );
  OR2_X1 U580 ( .A1(n759), .A2(n627), .ZN(n472) );
  INV_X1 U581 ( .A(KEYINPUT76), .ZN(n634) );
  NOR2_X1 U582 ( .A1(n761), .A2(n610), .ZN(n573) );
  XNOR2_X1 U583 ( .A(KEYINPUT90), .B(KEYINPUT39), .ZN(n606) );
  BUF_X1 U584 ( .A(n772), .Z(n775) );
  XNOR2_X1 U585 ( .A(KEYINPUT40), .B(KEYINPUT111), .ZN(n608) );
  AND2_X1 U586 ( .A1(n681), .A2(G953), .ZN(n777) );
  NAND2_X1 U587 ( .A1(n605), .A2(n591), .ZN(n617) );
  XNOR2_X2 U588 ( .A(G143), .B(G128), .ZN(n553) );
  XNOR2_X2 U589 ( .A(n474), .B(n519), .ZN(n506) );
  XNOR2_X1 U590 ( .A(n475), .B(G137), .ZN(n490) );
  XNOR2_X2 U591 ( .A(n506), .B(n490), .ZN(n790) );
  XNOR2_X1 U592 ( .A(n477), .B(n476), .ZN(n480) );
  XNOR2_X1 U593 ( .A(KEYINPUT73), .B(G110), .ZN(n515) );
  NAND2_X1 U594 ( .A1(G227), .A2(n793), .ZN(n478) );
  XNOR2_X1 U595 ( .A(n515), .B(n478), .ZN(n479) );
  XNOR2_X1 U596 ( .A(n480), .B(n479), .ZN(n481) );
  XNOR2_X1 U597 ( .A(KEYINPUT71), .B(KEYINPUT70), .ZN(n482) );
  INV_X1 U598 ( .A(KEYINPUT1), .ZN(n485) );
  XNOR2_X2 U599 ( .A(n614), .B(n485), .ZN(n711) );
  XNOR2_X1 U600 ( .A(KEYINPUT24), .B(KEYINPUT98), .ZN(n486) );
  NAND2_X1 U601 ( .A1(G234), .A2(n793), .ZN(n487) );
  XNOR2_X2 U602 ( .A(n488), .B(G125), .ZN(n516) );
  XNOR2_X2 U603 ( .A(n516), .B(n489), .ZN(n536) );
  XNOR2_X1 U604 ( .A(n536), .B(n490), .ZN(n491) );
  NOR2_X1 U605 ( .A1(n772), .A2(G902), .ZN(n497) );
  XOR2_X1 U606 ( .A(KEYINPUT20), .B(KEYINPUT101), .Z(n493) );
  NAND2_X1 U607 ( .A1(G234), .A2(n521), .ZN(n492) );
  XNOR2_X1 U608 ( .A(n493), .B(n492), .ZN(n559) );
  NAND2_X1 U609 ( .A1(n559), .A2(G217), .ZN(n495) );
  XOR2_X1 U610 ( .A(KEYINPUT25), .B(KEYINPUT80), .Z(n494) );
  XNOR2_X1 U611 ( .A(n495), .B(n494), .ZN(n496) );
  XNOR2_X1 U612 ( .A(G137), .B(n411), .ZN(n498) );
  NAND2_X1 U613 ( .A1(n541), .A2(G210), .ZN(n500) );
  XNOR2_X1 U614 ( .A(n501), .B(KEYINPUT3), .ZN(n504) );
  XNOR2_X1 U615 ( .A(n502), .B(G101), .ZN(n503) );
  XNOR2_X1 U616 ( .A(n504), .B(n503), .ZN(n511) );
  XNOR2_X1 U617 ( .A(n505), .B(n511), .ZN(n507) );
  INV_X1 U618 ( .A(n717), .ZN(n611) );
  AND2_X1 U619 ( .A1(n401), .A2(n611), .ZN(n508) );
  AND2_X1 U620 ( .A1(n711), .A2(n508), .ZN(n567) );
  XNOR2_X2 U621 ( .A(G116), .B(G107), .ZN(n554) );
  XNOR2_X1 U622 ( .A(KEYINPUT75), .B(KEYINPUT16), .ZN(n509) );
  XNOR2_X1 U623 ( .A(n554), .B(n509), .ZN(n510) );
  XNOR2_X1 U624 ( .A(n510), .B(n537), .ZN(n512) );
  XNOR2_X1 U625 ( .A(n512), .B(n511), .ZN(n784) );
  NAND2_X1 U626 ( .A1(n793), .A2(G224), .ZN(n513) );
  XNOR2_X1 U627 ( .A(n514), .B(n513), .ZN(n518) );
  XNOR2_X1 U628 ( .A(n516), .B(n515), .ZN(n517) );
  INV_X1 U629 ( .A(n521), .ZN(n670) );
  NAND2_X1 U630 ( .A1(n523), .A2(n522), .ZN(n526) );
  NAND2_X1 U631 ( .A1(n526), .A2(G210), .ZN(n524) );
  XNOR2_X1 U632 ( .A(n524), .B(KEYINPUT96), .ZN(n525) );
  NAND2_X1 U633 ( .A1(n526), .A2(G214), .ZN(n697) );
  INV_X1 U634 ( .A(n697), .ZN(n527) );
  XOR2_X1 U635 ( .A(KEYINPUT14), .B(KEYINPUT97), .Z(n529) );
  XNOR2_X1 U636 ( .A(n529), .B(n528), .ZN(n530) );
  NAND2_X1 U637 ( .A1(n530), .A2(G952), .ZN(n727) );
  NOR2_X1 U638 ( .A1(n727), .A2(G953), .ZN(n571) );
  NAND2_X1 U639 ( .A1(n530), .A2(G902), .ZN(n568) );
  INV_X1 U640 ( .A(G898), .ZN(n781) );
  NAND2_X1 U641 ( .A1(G953), .A2(n781), .ZN(n785) );
  NOR2_X1 U642 ( .A1(n568), .A2(n785), .ZN(n531) );
  OR2_X1 U643 ( .A1(n571), .A2(n531), .ZN(n532) );
  INV_X1 U644 ( .A(KEYINPUT0), .ZN(n533) );
  XNOR2_X2 U645 ( .A(n534), .B(n533), .ZN(n643) );
  XNOR2_X1 U646 ( .A(n536), .B(n535), .ZN(n540) );
  XOR2_X1 U647 ( .A(n538), .B(n537), .Z(n539) );
  XNOR2_X1 U648 ( .A(n540), .B(n539), .ZN(n546) );
  NAND2_X1 U649 ( .A1(G214), .A2(n541), .ZN(n542) );
  XNOR2_X1 U650 ( .A(n543), .B(n542), .ZN(n544) );
  XOR2_X1 U651 ( .A(n544), .B(KEYINPUT12), .Z(n545) );
  XNOR2_X1 U652 ( .A(n546), .B(n545), .ZN(n676) );
  NOR2_X1 U653 ( .A1(G902), .A2(n676), .ZN(n549) );
  XNOR2_X1 U654 ( .A(KEYINPUT107), .B(KEYINPUT13), .ZN(n547) );
  XNOR2_X1 U655 ( .A(n552), .B(n551), .ZN(n558) );
  XNOR2_X1 U656 ( .A(n553), .B(n554), .ZN(n556) );
  XOR2_X1 U657 ( .A(KEYINPUT7), .B(KEYINPUT9), .Z(n555) );
  XNOR2_X1 U658 ( .A(n556), .B(n555), .ZN(n557) );
  XNOR2_X1 U659 ( .A(n558), .B(n557), .ZN(n768) );
  NAND2_X1 U660 ( .A1(n398), .A2(n588), .ZN(n701) );
  NAND2_X1 U661 ( .A1(n559), .A2(G221), .ZN(n563) );
  XOR2_X1 U662 ( .A(KEYINPUT102), .B(KEYINPUT103), .Z(n561) );
  INV_X1 U663 ( .A(KEYINPUT21), .ZN(n560) );
  XNOR2_X1 U664 ( .A(n561), .B(n560), .ZN(n562) );
  XNOR2_X1 U665 ( .A(n563), .B(n562), .ZN(n708) );
  INV_X1 U666 ( .A(n708), .ZN(n583) );
  NOR2_X1 U667 ( .A1(n701), .A2(n583), .ZN(n564) );
  NAND2_X1 U668 ( .A1(n643), .A2(n564), .ZN(n565) );
  AND2_X1 U669 ( .A1(n567), .A2(n566), .ZN(n655) );
  XOR2_X1 U670 ( .A(G110), .B(n655), .Z(G12) );
  INV_X1 U671 ( .A(n588), .ZN(n618) );
  INV_X1 U672 ( .A(n758), .ZN(n761) );
  OR2_X1 U673 ( .A1(n793), .A2(n568), .ZN(n569) );
  NOR2_X1 U674 ( .A1(G900), .A2(n569), .ZN(n570) );
  NOR2_X1 U675 ( .A1(n586), .A2(n583), .ZN(n572) );
  NAND2_X1 U676 ( .A1(n401), .A2(n572), .ZN(n610) );
  NAND2_X1 U677 ( .A1(n573), .A2(n697), .ZN(n574) );
  NAND2_X1 U678 ( .A1(n636), .A2(n711), .ZN(n575) );
  XNOR2_X1 U679 ( .A(KEYINPUT43), .B(n575), .ZN(n576) );
  NAND2_X1 U680 ( .A1(n576), .A2(n635), .ZN(n639) );
  XNOR2_X1 U681 ( .A(G140), .B(KEYINPUT114), .ZN(n577) );
  XNOR2_X1 U682 ( .A(n639), .B(n577), .ZN(G42) );
  NAND2_X1 U683 ( .A1(n711), .A2(n400), .ZN(n578) );
  XNOR2_X1 U684 ( .A(n653), .B(G101), .ZN(G3) );
  OR2_X1 U685 ( .A1(n711), .A2(n400), .ZN(n579) );
  XNOR2_X1 U686 ( .A(G119), .B(KEYINPUT125), .ZN(n582) );
  XNOR2_X1 U687 ( .A(n656), .B(n582), .ZN(G21) );
  NOR2_X2 U688 ( .A1(n584), .A2(n583), .ZN(n592) );
  NAND2_X1 U689 ( .A1(n697), .A2(n717), .ZN(n587) );
  OR2_X1 U690 ( .A1(n398), .A2(n588), .ZN(n589) );
  XNOR2_X1 U691 ( .A(n589), .B(KEYINPUT109), .ZN(n600) );
  INV_X1 U692 ( .A(n635), .ZN(n590) );
  XNOR2_X1 U693 ( .A(n617), .B(G143), .ZN(G45) );
  INV_X1 U694 ( .A(n362), .ZN(n710) );
  INV_X1 U695 ( .A(n643), .ZN(n648) );
  XNOR2_X1 U696 ( .A(KEYINPUT82), .B(KEYINPUT34), .ZN(n597) );
  INV_X1 U697 ( .A(KEYINPUT74), .ZN(n596) );
  XNOR2_X1 U698 ( .A(n597), .B(n596), .ZN(n598) );
  XNOR2_X1 U699 ( .A(n599), .B(n598), .ZN(n601) );
  NAND2_X1 U700 ( .A1(n601), .A2(n600), .ZN(n604) );
  INV_X1 U701 ( .A(KEYINPUT81), .ZN(n602) );
  XNOR2_X1 U702 ( .A(n602), .B(KEYINPUT35), .ZN(n603) );
  XNOR2_X2 U703 ( .A(n604), .B(n603), .ZN(n658) );
  XOR2_X1 U704 ( .A(n658), .B(G122), .Z(G24) );
  XNOR2_X1 U705 ( .A(n612), .B(KEYINPUT28), .ZN(n613) );
  NAND2_X1 U706 ( .A1(n614), .A2(n613), .ZN(n626) );
  NAND2_X1 U707 ( .A1(n698), .A2(n697), .ZN(n702) );
  NOR2_X1 U708 ( .A1(n701), .A2(n702), .ZN(n615) );
  XNOR2_X1 U709 ( .A(n615), .B(KEYINPUT41), .ZN(n728) );
  NOR2_X1 U710 ( .A1(n626), .A2(n728), .ZN(n616) );
  NOR2_X1 U711 ( .A1(KEYINPUT84), .A2(KEYINPUT47), .ZN(n623) );
  XNOR2_X2 U712 ( .A(n620), .B(KEYINPUT108), .ZN(n703) );
  NAND2_X1 U713 ( .A1(n703), .A2(KEYINPUT47), .ZN(n621) );
  XNOR2_X1 U714 ( .A(n621), .B(KEYINPUT85), .ZN(n622) );
  NOR2_X1 U715 ( .A1(n623), .A2(n622), .ZN(n628) );
  INV_X1 U716 ( .A(n624), .ZN(n625) );
  NOR2_X2 U717 ( .A1(n626), .A2(n625), .ZN(n759) );
  NAND2_X1 U718 ( .A1(KEYINPUT47), .A2(KEYINPUT84), .ZN(n627) );
  AND2_X1 U719 ( .A1(n628), .A2(n472), .ZN(n633) );
  XOR2_X1 U720 ( .A(KEYINPUT47), .B(KEYINPUT65), .Z(n629) );
  NOR2_X1 U721 ( .A1(n703), .A2(n629), .ZN(n630) );
  NAND2_X1 U722 ( .A1(n631), .A2(n759), .ZN(n632) );
  NAND2_X1 U723 ( .A1(n636), .A2(n590), .ZN(n637) );
  NAND2_X1 U724 ( .A1(n364), .A2(n754), .ZN(n641) );
  XNOR2_X1 U725 ( .A(n641), .B(KEYINPUT112), .ZN(n804) );
  NOR2_X1 U726 ( .A1(n642), .A2(n717), .ZN(n644) );
  NAND2_X1 U727 ( .A1(n644), .A2(n643), .ZN(n646) );
  INV_X1 U728 ( .A(KEYINPUT105), .ZN(n645) );
  XNOR2_X1 U729 ( .A(n646), .B(n645), .ZN(n750) );
  NAND2_X1 U730 ( .A1(n717), .A2(n362), .ZN(n647) );
  OR2_X1 U731 ( .A1(n711), .A2(n647), .ZN(n707) );
  XNOR2_X1 U732 ( .A(KEYINPUT106), .B(KEYINPUT31), .ZN(n649) );
  XNOR2_X1 U733 ( .A(n650), .B(n649), .ZN(n764) );
  NAND2_X1 U734 ( .A1(n750), .A2(n764), .ZN(n652) );
  INV_X1 U735 ( .A(n703), .ZN(n651) );
  NAND2_X1 U736 ( .A1(n652), .A2(n651), .ZN(n654) );
  XNOR2_X1 U737 ( .A(n657), .B(KEYINPUT91), .ZN(n665) );
  INV_X1 U738 ( .A(n658), .ZN(n660) );
  INV_X1 U739 ( .A(KEYINPUT44), .ZN(n659) );
  AND2_X1 U740 ( .A1(n660), .A2(n659), .ZN(n663) );
  INV_X1 U741 ( .A(n661), .ZN(n662) );
  NAND2_X1 U742 ( .A1(n663), .A2(n662), .ZN(n664) );
  NAND2_X1 U743 ( .A1(n665), .A2(n664), .ZN(n666) );
  OR2_X1 U744 ( .A1(KEYINPUT87), .A2(n521), .ZN(n667) );
  NOR2_X1 U745 ( .A1(n691), .A2(n667), .ZN(n669) );
  AND2_X1 U746 ( .A1(n670), .A2(KEYINPUT2), .ZN(n668) );
  NOR2_X1 U747 ( .A1(n669), .A2(n668), .ZN(n674) );
  INV_X1 U748 ( .A(n691), .ZN(n671) );
  NAND2_X1 U749 ( .A1(n671), .A2(n670), .ZN(n672) );
  NAND2_X1 U750 ( .A1(n672), .A2(KEYINPUT87), .ZN(n673) );
  NAND2_X1 U751 ( .A1(n673), .A2(n674), .ZN(n675) );
  NAND2_X1 U752 ( .A1(n773), .A2(G475), .ZN(n680) );
  XNOR2_X1 U753 ( .A(KEYINPUT95), .B(KEYINPUT121), .ZN(n677) );
  XNOR2_X1 U754 ( .A(n677), .B(KEYINPUT59), .ZN(n678) );
  XNOR2_X1 U755 ( .A(n680), .B(n679), .ZN(n682) );
  INV_X1 U756 ( .A(G952), .ZN(n681) );
  INV_X1 U757 ( .A(n777), .ZN(n740) );
  NAND2_X1 U758 ( .A1(n682), .A2(n740), .ZN(n684) );
  INV_X1 U759 ( .A(KEYINPUT60), .ZN(n683) );
  XNOR2_X1 U760 ( .A(n684), .B(n683), .ZN(G60) );
  NAND2_X1 U761 ( .A1(n773), .A2(G472), .ZN(n687) );
  XNOR2_X1 U762 ( .A(n687), .B(n686), .ZN(n688) );
  NAND2_X1 U763 ( .A1(n688), .A2(n740), .ZN(n689) );
  XNOR2_X1 U764 ( .A(n689), .B(KEYINPUT63), .ZN(G57) );
  INV_X1 U765 ( .A(KEYINPUT2), .ZN(n690) );
  NAND2_X1 U766 ( .A1(n691), .A2(n690), .ZN(n693) );
  INV_X1 U767 ( .A(KEYINPUT83), .ZN(n692) );
  NOR2_X1 U768 ( .A1(n698), .A2(n697), .ZN(n699) );
  XNOR2_X1 U769 ( .A(n699), .B(KEYINPUT116), .ZN(n700) );
  NOR2_X1 U770 ( .A1(n701), .A2(n700), .ZN(n705) );
  NOR2_X1 U771 ( .A1(n703), .A2(n702), .ZN(n704) );
  NOR2_X1 U772 ( .A1(n705), .A2(n704), .ZN(n706) );
  INV_X1 U773 ( .A(n707), .ZN(n719) );
  NOR2_X1 U774 ( .A1(n400), .A2(n708), .ZN(n709) );
  XNOR2_X1 U775 ( .A(KEYINPUT49), .B(n709), .ZN(n715) );
  XOR2_X1 U776 ( .A(KEYINPUT50), .B(KEYINPUT115), .Z(n713) );
  NAND2_X1 U777 ( .A1(n711), .A2(n710), .ZN(n712) );
  XNOR2_X1 U778 ( .A(n713), .B(n712), .ZN(n714) );
  NAND2_X1 U779 ( .A1(n715), .A2(n714), .ZN(n716) );
  NOR2_X1 U780 ( .A1(n717), .A2(n716), .ZN(n718) );
  NOR2_X1 U781 ( .A1(n719), .A2(n718), .ZN(n720) );
  XOR2_X1 U782 ( .A(KEYINPUT51), .B(n720), .Z(n721) );
  NOR2_X1 U783 ( .A1(n728), .A2(n721), .ZN(n722) );
  NOR2_X1 U784 ( .A1(n723), .A2(n722), .ZN(n724) );
  XOR2_X1 U785 ( .A(KEYINPUT52), .B(n724), .Z(n725) );
  XNOR2_X1 U786 ( .A(n725), .B(KEYINPUT117), .ZN(n726) );
  NOR2_X1 U787 ( .A1(n727), .A2(n726), .ZN(n730) );
  NOR2_X1 U788 ( .A1(n730), .A2(n729), .ZN(n731) );
  XNOR2_X1 U789 ( .A(n731), .B(KEYINPUT118), .ZN(n732) );
  XOR2_X1 U790 ( .A(KEYINPUT120), .B(KEYINPUT53), .Z(n733) );
  XNOR2_X1 U791 ( .A(n734), .B(n733), .ZN(G75) );
  NAND2_X1 U792 ( .A1(n773), .A2(G210), .ZN(n739) );
  XNOR2_X1 U793 ( .A(KEYINPUT94), .B(KEYINPUT54), .ZN(n735) );
  XNOR2_X1 U794 ( .A(n735), .B(KEYINPUT55), .ZN(n736) );
  XNOR2_X1 U795 ( .A(n739), .B(n738), .ZN(n741) );
  NAND2_X1 U796 ( .A1(n741), .A2(n740), .ZN(n743) );
  INV_X1 U797 ( .A(KEYINPUT56), .ZN(n742) );
  XNOR2_X1 U798 ( .A(n743), .B(n742), .ZN(G51) );
  NAND2_X1 U799 ( .A1(n773), .A2(G469), .ZN(n747) );
  XOR2_X1 U800 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n744) );
  XNOR2_X1 U801 ( .A(n365), .B(n744), .ZN(n746) );
  XNOR2_X1 U802 ( .A(n747), .B(n746), .ZN(n748) );
  NOR2_X1 U803 ( .A1(n748), .A2(n777), .ZN(G54) );
  NOR2_X1 U804 ( .A1(n761), .A2(n750), .ZN(n749) );
  XOR2_X1 U805 ( .A(G104), .B(n749), .Z(G6) );
  INV_X1 U806 ( .A(n754), .ZN(n763) );
  NOR2_X1 U807 ( .A1(n763), .A2(n750), .ZN(n752) );
  XNOR2_X1 U808 ( .A(KEYINPUT27), .B(KEYINPUT26), .ZN(n751) );
  XNOR2_X1 U809 ( .A(n752), .B(n751), .ZN(n753) );
  XNOR2_X1 U810 ( .A(G107), .B(n753), .ZN(G9) );
  XOR2_X1 U811 ( .A(KEYINPUT29), .B(KEYINPUT113), .Z(n756) );
  NAND2_X1 U812 ( .A1(n759), .A2(n754), .ZN(n755) );
  XNOR2_X1 U813 ( .A(n756), .B(n755), .ZN(n757) );
  XOR2_X1 U814 ( .A(G128), .B(n757), .Z(G30) );
  NAND2_X1 U815 ( .A1(n759), .A2(n758), .ZN(n760) );
  XNOR2_X1 U816 ( .A(n760), .B(n411), .ZN(G48) );
  NOR2_X1 U817 ( .A1(n764), .A2(n761), .ZN(n762) );
  XOR2_X1 U818 ( .A(G113), .B(n762), .Z(G15) );
  NOR2_X1 U819 ( .A1(n764), .A2(n763), .ZN(n765) );
  XOR2_X1 U820 ( .A(G116), .B(n765), .Z(G18) );
  XNOR2_X1 U821 ( .A(G125), .B(n766), .ZN(n767) );
  XNOR2_X1 U822 ( .A(n767), .B(KEYINPUT37), .ZN(G27) );
  NAND2_X1 U823 ( .A1(n773), .A2(G478), .ZN(n770) );
  XNOR2_X1 U824 ( .A(n768), .B(KEYINPUT122), .ZN(n769) );
  XNOR2_X1 U825 ( .A(n770), .B(n769), .ZN(n771) );
  NOR2_X1 U826 ( .A1(n777), .A2(n771), .ZN(G63) );
  NAND2_X1 U827 ( .A1(n773), .A2(G217), .ZN(n774) );
  XNOR2_X1 U828 ( .A(n775), .B(n774), .ZN(n776) );
  NOR2_X1 U829 ( .A1(n777), .A2(n776), .ZN(G66) );
  AND2_X1 U830 ( .A1(n778), .A2(n793), .ZN(n783) );
  NAND2_X1 U831 ( .A1(G953), .A2(G224), .ZN(n779) );
  XOR2_X1 U832 ( .A(KEYINPUT61), .B(n779), .Z(n780) );
  NOR2_X1 U833 ( .A1(n781), .A2(n780), .ZN(n782) );
  NOR2_X1 U834 ( .A1(n783), .A2(n782), .ZN(n789) );
  XOR2_X1 U835 ( .A(G110), .B(n784), .Z(n786) );
  NAND2_X1 U836 ( .A1(n786), .A2(n785), .ZN(n787) );
  XNOR2_X1 U837 ( .A(n787), .B(KEYINPUT123), .ZN(n788) );
  XOR2_X1 U838 ( .A(n789), .B(n788), .Z(G69) );
  XNOR2_X1 U839 ( .A(n536), .B(n402), .ZN(n796) );
  INV_X1 U840 ( .A(n791), .ZN(n792) );
  XNOR2_X1 U841 ( .A(n796), .B(n792), .ZN(n794) );
  NAND2_X1 U842 ( .A1(n794), .A2(n793), .ZN(n795) );
  XNOR2_X1 U843 ( .A(n795), .B(KEYINPUT124), .ZN(n800) );
  XNOR2_X1 U844 ( .A(G227), .B(n796), .ZN(n797) );
  NAND2_X1 U845 ( .A1(n797), .A2(G900), .ZN(n798) );
  NAND2_X1 U846 ( .A1(G953), .A2(n798), .ZN(n799) );
  NAND2_X1 U847 ( .A1(n800), .A2(n799), .ZN(G72) );
  XOR2_X1 U848 ( .A(G137), .B(KEYINPUT126), .Z(n801) );
  XNOR2_X1 U849 ( .A(n802), .B(n801), .ZN(G39) );
  XOR2_X1 U850 ( .A(n370), .B(G131), .Z(G33) );
  XNOR2_X1 U851 ( .A(G134), .B(n804), .ZN(G36) );
endmodule

