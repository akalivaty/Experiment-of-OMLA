

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588,
         n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599,
         n600, n601, n602, n603, n604, n605, n606, n607, n608, n609, n610,
         n611, n612, n613, n614, n615, n616, n617, n618, n619, n620, n621,
         n622, n623, n624, n625, n626, n627, n628, n629, n630, n631, n632,
         n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, n643,
         n644, n645, n646, n647, n648, n649, n650, n651, n652, n653, n654,
         n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, n665,
         n666, n667, n668, n669, n670, n671, n672, n673, n674, n675, n676,
         n677, n678, n679, n680, n681, n682, n683, n684, n685, n686, n687,
         n688, n689, n690, n691, n692, n693, n694, n695, n696, n697, n698,
         n699, n700, n701, n702, n703, n704, n705, n706, n707, n708, n709,
         n710, n711, n712, n713, n714, n715, n716, n717, n718, n719, n720,
         n721, n722, n723, n724, n725, n726, n727, n728, n729, n730, n731,
         n732, n733, n734, n735, n736, n737, n738, n739, n740, n741, n742,
         n743, n744, n745, n746, n747, n748, n749, n750, n751, n752, n753,
         n754, n755, n756, n757, n758, n759, n760, n761, n762, n763, n764,
         n765, n766, n767, n768, n769, n770, n771, n772, n773, n774, n775,
         n776, n777, n778, n779, n780, n781, n782, n783, n784, n785, n786,
         n787, n788, n789, n790, n791, n792, n793, n794, n795, n796, n797,
         n798, n799, n800, n801, n802, n803, n804, n805, n806, n807, n808,
         n809, n810, n811, n812, n813, n814, n815, n816, n817, n818, n819,
         n820, n821, n822, n823, n824, n825, n826, n827, n828, n829, n830,
         n831, n832, n833, n834, n835, n836, n837, n838, n839, n840, n841,
         n842, n843, n844, n845, n846, n847, n848, n849, n850, n851, n852,
         n853, n854, n855, n856, n857, n858, n859, n860, n861, n862, n863,
         n864, n865, n866, n867, n868, n869, n870, n871, n872, n873, n874,
         n875, n876, n877, n878, n879, n880, n881, n882, n883, n884, n885,
         n886, n887, n888, n889, n890, n891, n892, n893, n894, n895, n896,
         n897, n898, n899, n900, n901, n902, n903, n904, n905, n906, n907,
         n908, n909, n910, n911, n912, n913, n914, n915, n916, n917, n918,
         n919, n920, n921, n922, n923, n924, n925, n926, n927, n928, n929,
         n930, n931, n932, n933, n934, n935, n936, n937, n938, n939, n940,
         n941, n942, n943, n944, n945, n946, n947, n948, n949, n950, n951,
         n952, n953, n954, n955, n956, n957, n958, n959, n960, n961, n962,
         n963, n964, n965, n966, n967, n968, n969, n970, n971, n972, n973,
         n974, n975, n976, n977, n978, n979, n980, n981, n982, n983, n984,
         n985, n986, n987, n988, n989, n990, n991, n992, n993, n994, n995,
         n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005,
         n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015,
         n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025,
         n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NOR2_X2 U554 ( .A1(n755), .A2(n757), .ZN(n760) );
  INV_X1 U555 ( .A(n773), .ZN(n748) );
  XNOR2_X1 U556 ( .A(KEYINPUT15), .B(n588), .ZN(n965) );
  NOR2_X2 U557 ( .A1(n580), .A2(n579), .ZN(n962) );
  NOR2_X1 U558 ( .A1(G164), .A2(G1384), .ZN(n718) );
  AND2_X1 U559 ( .A1(n533), .A2(n532), .ZN(G164) );
  XNOR2_X1 U560 ( .A(n814), .B(KEYINPUT99), .ZN(n818) );
  XOR2_X1 U561 ( .A(n765), .B(n764), .Z(n519) );
  NOR2_X1 U562 ( .A1(n794), .A2(n793), .ZN(n520) );
  OR2_X1 U563 ( .A1(n817), .A2(n816), .ZN(n521) );
  AND2_X1 U564 ( .A1(n885), .A2(G114), .ZN(n522) );
  INV_X1 U565 ( .A(KEYINPUT95), .ZN(n761) );
  XNOR2_X1 U566 ( .A(KEYINPUT90), .B(KEYINPUT27), .ZN(n733) );
  XNOR2_X1 U567 ( .A(n734), .B(n733), .ZN(n736) );
  AND2_X1 U568 ( .A1(n818), .A2(n521), .ZN(n822) );
  NOR2_X1 U569 ( .A1(n822), .A2(n821), .ZN(n823) );
  AND2_X2 U570 ( .A1(n525), .A2(G2104), .ZN(n881) );
  INV_X1 U571 ( .A(KEYINPUT101), .ZN(n827) );
  NOR2_X2 U572 ( .A1(n623), .A2(n544), .ZN(n644) );
  XNOR2_X1 U573 ( .A(n828), .B(n827), .ZN(n829) );
  XOR2_X1 U574 ( .A(KEYINPUT0), .B(G543), .Z(n623) );
  INV_X1 U575 ( .A(G2105), .ZN(n525) );
  NOR2_X4 U576 ( .A1(G2104), .A2(n525), .ZN(n886) );
  NAND2_X1 U577 ( .A1(G126), .A2(n886), .ZN(n523) );
  XNOR2_X1 U578 ( .A(KEYINPUT83), .B(n523), .ZN(n524) );
  AND2_X1 U579 ( .A1(G2105), .A2(G2104), .ZN(n885) );
  NOR2_X1 U580 ( .A1(n524), .A2(n522), .ZN(n533) );
  NAND2_X1 U581 ( .A1(G102), .A2(n881), .ZN(n529) );
  XNOR2_X1 U582 ( .A(KEYINPUT65), .B(KEYINPUT17), .ZN(n527) );
  NOR2_X1 U583 ( .A1(G2105), .A2(G2104), .ZN(n526) );
  XNOR2_X1 U584 ( .A(n527), .B(n526), .ZN(n534) );
  NAND2_X1 U585 ( .A1(G138), .A2(n534), .ZN(n528) );
  NAND2_X1 U586 ( .A1(n529), .A2(n528), .ZN(n531) );
  INV_X1 U587 ( .A(KEYINPUT84), .ZN(n530) );
  XNOR2_X1 U588 ( .A(n531), .B(n530), .ZN(n532) );
  BUF_X1 U589 ( .A(n534), .Z(n882) );
  NAND2_X1 U590 ( .A1(n882), .A2(G137), .ZN(n537) );
  NAND2_X1 U591 ( .A1(G101), .A2(n881), .ZN(n535) );
  XOR2_X1 U592 ( .A(KEYINPUT23), .B(n535), .Z(n536) );
  AND2_X1 U593 ( .A1(n537), .A2(n536), .ZN(n687) );
  NAND2_X1 U594 ( .A1(G113), .A2(n885), .ZN(n539) );
  NAND2_X1 U595 ( .A1(G125), .A2(n886), .ZN(n538) );
  AND2_X1 U596 ( .A1(n539), .A2(n538), .ZN(n686) );
  AND2_X1 U597 ( .A1(n687), .A2(n686), .ZN(G160) );
  AND2_X1 U598 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U599 ( .A(G651), .ZN(n544) );
  NOR2_X1 U600 ( .A1(G543), .A2(n544), .ZN(n540) );
  XOR2_X1 U601 ( .A(KEYINPUT1), .B(n540), .Z(n647) );
  NAND2_X1 U602 ( .A1(G65), .A2(n647), .ZN(n543) );
  NOR2_X1 U603 ( .A1(G651), .A2(n623), .ZN(n541) );
  XNOR2_X2 U604 ( .A(KEYINPUT64), .B(n541), .ZN(n649) );
  NAND2_X1 U605 ( .A1(G53), .A2(n649), .ZN(n542) );
  NAND2_X1 U606 ( .A1(n543), .A2(n542), .ZN(n548) );
  NOR2_X1 U607 ( .A1(G651), .A2(G543), .ZN(n643) );
  NAND2_X1 U608 ( .A1(G91), .A2(n643), .ZN(n546) );
  NAND2_X1 U609 ( .A1(G78), .A2(n644), .ZN(n545) );
  NAND2_X1 U610 ( .A1(n546), .A2(n545), .ZN(n547) );
  NOR2_X1 U611 ( .A1(n548), .A2(n547), .ZN(n739) );
  INV_X1 U612 ( .A(n739), .ZN(G299) );
  INV_X1 U613 ( .A(G57), .ZN(G237) );
  INV_X1 U614 ( .A(G132), .ZN(G219) );
  INV_X1 U615 ( .A(G82), .ZN(G220) );
  NAND2_X1 U616 ( .A1(G64), .A2(n647), .ZN(n550) );
  NAND2_X1 U617 ( .A1(G52), .A2(n649), .ZN(n549) );
  NAND2_X1 U618 ( .A1(n550), .A2(n549), .ZN(n551) );
  XNOR2_X1 U619 ( .A(KEYINPUT68), .B(n551), .ZN(n557) );
  NAND2_X1 U620 ( .A1(G90), .A2(n643), .ZN(n553) );
  NAND2_X1 U621 ( .A1(G77), .A2(n644), .ZN(n552) );
  NAND2_X1 U622 ( .A1(n553), .A2(n552), .ZN(n554) );
  XNOR2_X1 U623 ( .A(KEYINPUT69), .B(n554), .ZN(n555) );
  XNOR2_X1 U624 ( .A(KEYINPUT9), .B(n555), .ZN(n556) );
  NOR2_X1 U625 ( .A1(n557), .A2(n556), .ZN(G171) );
  NAND2_X1 U626 ( .A1(n643), .A2(G89), .ZN(n558) );
  XNOR2_X1 U627 ( .A(n558), .B(KEYINPUT4), .ZN(n560) );
  NAND2_X1 U628 ( .A1(G76), .A2(n644), .ZN(n559) );
  NAND2_X1 U629 ( .A1(n560), .A2(n559), .ZN(n561) );
  XNOR2_X1 U630 ( .A(n561), .B(KEYINPUT5), .ZN(n566) );
  NAND2_X1 U631 ( .A1(G63), .A2(n647), .ZN(n563) );
  NAND2_X1 U632 ( .A1(G51), .A2(n649), .ZN(n562) );
  NAND2_X1 U633 ( .A1(n563), .A2(n562), .ZN(n564) );
  XOR2_X1 U634 ( .A(KEYINPUT6), .B(n564), .Z(n565) );
  NAND2_X1 U635 ( .A1(n566), .A2(n565), .ZN(n567) );
  XNOR2_X1 U636 ( .A(n567), .B(KEYINPUT7), .ZN(G168) );
  XOR2_X1 U637 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U638 ( .A1(G7), .A2(G661), .ZN(n568) );
  XOR2_X1 U639 ( .A(n568), .B(KEYINPUT10), .Z(n832) );
  NAND2_X1 U640 ( .A1(n832), .A2(G567), .ZN(n569) );
  XOR2_X1 U641 ( .A(KEYINPUT11), .B(n569), .Z(G234) );
  XNOR2_X1 U642 ( .A(G860), .B(KEYINPUT72), .ZN(n593) );
  XOR2_X1 U643 ( .A(KEYINPUT70), .B(KEYINPUT14), .Z(n571) );
  NAND2_X1 U644 ( .A1(G56), .A2(n647), .ZN(n570) );
  XNOR2_X1 U645 ( .A(n571), .B(n570), .ZN(n580) );
  NAND2_X1 U646 ( .A1(n643), .A2(G81), .ZN(n572) );
  XNOR2_X1 U647 ( .A(KEYINPUT12), .B(n572), .ZN(n575) );
  NAND2_X1 U648 ( .A1(n644), .A2(G68), .ZN(n573) );
  XOR2_X1 U649 ( .A(KEYINPUT71), .B(n573), .Z(n574) );
  NAND2_X1 U650 ( .A1(n575), .A2(n574), .ZN(n576) );
  XNOR2_X1 U651 ( .A(n576), .B(KEYINPUT13), .ZN(n578) );
  NAND2_X1 U652 ( .A1(G43), .A2(n649), .ZN(n577) );
  NAND2_X1 U653 ( .A1(n578), .A2(n577), .ZN(n579) );
  NAND2_X1 U654 ( .A1(n593), .A2(n962), .ZN(n581) );
  XOR2_X1 U655 ( .A(KEYINPUT73), .B(n581), .Z(G153) );
  INV_X1 U656 ( .A(G171), .ZN(G301) );
  NAND2_X1 U657 ( .A1(G868), .A2(G301), .ZN(n590) );
  NAND2_X1 U658 ( .A1(G92), .A2(n643), .ZN(n583) );
  NAND2_X1 U659 ( .A1(G66), .A2(n647), .ZN(n582) );
  NAND2_X1 U660 ( .A1(n583), .A2(n582), .ZN(n587) );
  NAND2_X1 U661 ( .A1(G79), .A2(n644), .ZN(n585) );
  NAND2_X1 U662 ( .A1(G54), .A2(n649), .ZN(n584) );
  NAND2_X1 U663 ( .A1(n585), .A2(n584), .ZN(n586) );
  NOR2_X1 U664 ( .A1(n587), .A2(n586), .ZN(n588) );
  INV_X1 U665 ( .A(G868), .ZN(n663) );
  NAND2_X1 U666 ( .A1(n965), .A2(n663), .ZN(n589) );
  NAND2_X1 U667 ( .A1(n590), .A2(n589), .ZN(G284) );
  NOR2_X1 U668 ( .A1(G286), .A2(n663), .ZN(n592) );
  NOR2_X1 U669 ( .A1(G868), .A2(G299), .ZN(n591) );
  NOR2_X1 U670 ( .A1(n592), .A2(n591), .ZN(G297) );
  INV_X1 U671 ( .A(G559), .ZN(n594) );
  NOR2_X1 U672 ( .A1(n594), .A2(n593), .ZN(n595) );
  NOR2_X1 U673 ( .A1(n965), .A2(n595), .ZN(n596) );
  XOR2_X1 U674 ( .A(KEYINPUT16), .B(n596), .Z(G148) );
  NOR2_X1 U675 ( .A1(n965), .A2(n663), .ZN(n597) );
  XNOR2_X1 U676 ( .A(n597), .B(KEYINPUT75), .ZN(n598) );
  NOR2_X1 U677 ( .A1(G559), .A2(n598), .ZN(n601) );
  NAND2_X1 U678 ( .A1(n962), .A2(n663), .ZN(n599) );
  XOR2_X1 U679 ( .A(KEYINPUT74), .B(n599), .Z(n600) );
  NOR2_X1 U680 ( .A1(n601), .A2(n600), .ZN(G282) );
  NAND2_X1 U681 ( .A1(G135), .A2(n882), .ZN(n603) );
  NAND2_X1 U682 ( .A1(G111), .A2(n885), .ZN(n602) );
  NAND2_X1 U683 ( .A1(n603), .A2(n602), .ZN(n606) );
  NAND2_X1 U684 ( .A1(n886), .A2(G123), .ZN(n604) );
  XOR2_X1 U685 ( .A(KEYINPUT18), .B(n604), .Z(n605) );
  NOR2_X1 U686 ( .A1(n606), .A2(n605), .ZN(n608) );
  NAND2_X1 U687 ( .A1(n881), .A2(G99), .ZN(n607) );
  NAND2_X1 U688 ( .A1(n608), .A2(n607), .ZN(n928) );
  XNOR2_X1 U689 ( .A(G2096), .B(n928), .ZN(n609) );
  NOR2_X1 U690 ( .A1(G2100), .A2(n609), .ZN(n610) );
  XOR2_X1 U691 ( .A(KEYINPUT76), .B(n610), .Z(G156) );
  INV_X1 U692 ( .A(n965), .ZN(n724) );
  NAND2_X1 U693 ( .A1(G559), .A2(n724), .ZN(n611) );
  XOR2_X1 U694 ( .A(n611), .B(n962), .Z(n661) );
  NOR2_X1 U695 ( .A1(n661), .A2(G860), .ZN(n619) );
  NAND2_X1 U696 ( .A1(G67), .A2(n647), .ZN(n613) );
  NAND2_X1 U697 ( .A1(G55), .A2(n649), .ZN(n612) );
  NAND2_X1 U698 ( .A1(n613), .A2(n612), .ZN(n618) );
  NAND2_X1 U699 ( .A1(G93), .A2(n643), .ZN(n615) );
  NAND2_X1 U700 ( .A1(G80), .A2(n644), .ZN(n614) );
  NAND2_X1 U701 ( .A1(n615), .A2(n614), .ZN(n616) );
  XOR2_X1 U702 ( .A(KEYINPUT77), .B(n616), .Z(n617) );
  OR2_X1 U703 ( .A1(n618), .A2(n617), .ZN(n664) );
  XOR2_X1 U704 ( .A(n619), .B(n664), .Z(G145) );
  NAND2_X1 U705 ( .A1(G651), .A2(G74), .ZN(n621) );
  NAND2_X1 U706 ( .A1(G49), .A2(n649), .ZN(n620) );
  NAND2_X1 U707 ( .A1(n621), .A2(n620), .ZN(n622) );
  NOR2_X1 U708 ( .A1(n647), .A2(n622), .ZN(n625) );
  NAND2_X1 U709 ( .A1(n623), .A2(G87), .ZN(n624) );
  NAND2_X1 U710 ( .A1(n625), .A2(n624), .ZN(G288) );
  XOR2_X1 U711 ( .A(KEYINPUT79), .B(KEYINPUT2), .Z(n627) );
  NAND2_X1 U712 ( .A1(G73), .A2(n644), .ZN(n626) );
  XNOR2_X1 U713 ( .A(n627), .B(n626), .ZN(n634) );
  NAND2_X1 U714 ( .A1(G86), .A2(n643), .ZN(n629) );
  NAND2_X1 U715 ( .A1(G48), .A2(n649), .ZN(n628) );
  NAND2_X1 U716 ( .A1(n629), .A2(n628), .ZN(n632) );
  NAND2_X1 U717 ( .A1(n647), .A2(G61), .ZN(n630) );
  XOR2_X1 U718 ( .A(KEYINPUT78), .B(n630), .Z(n631) );
  NOR2_X1 U719 ( .A1(n632), .A2(n631), .ZN(n633) );
  NAND2_X1 U720 ( .A1(n634), .A2(n633), .ZN(G305) );
  NAND2_X1 U721 ( .A1(G85), .A2(n643), .ZN(n635) );
  XNOR2_X1 U722 ( .A(n635), .B(KEYINPUT66), .ZN(n637) );
  NAND2_X1 U723 ( .A1(n647), .A2(G60), .ZN(n636) );
  NAND2_X1 U724 ( .A1(n637), .A2(n636), .ZN(n640) );
  NAND2_X1 U725 ( .A1(G72), .A2(n644), .ZN(n638) );
  XNOR2_X1 U726 ( .A(KEYINPUT67), .B(n638), .ZN(n639) );
  NOR2_X1 U727 ( .A1(n640), .A2(n639), .ZN(n642) );
  NAND2_X1 U728 ( .A1(G47), .A2(n649), .ZN(n641) );
  NAND2_X1 U729 ( .A1(n642), .A2(n641), .ZN(G290) );
  NAND2_X1 U730 ( .A1(G88), .A2(n643), .ZN(n646) );
  NAND2_X1 U731 ( .A1(G75), .A2(n644), .ZN(n645) );
  NAND2_X1 U732 ( .A1(n646), .A2(n645), .ZN(n653) );
  NAND2_X1 U733 ( .A1(n647), .A2(G62), .ZN(n648) );
  XNOR2_X1 U734 ( .A(n648), .B(KEYINPUT80), .ZN(n651) );
  NAND2_X1 U735 ( .A1(G50), .A2(n649), .ZN(n650) );
  NAND2_X1 U736 ( .A1(n651), .A2(n650), .ZN(n652) );
  NOR2_X1 U737 ( .A1(n653), .A2(n652), .ZN(G166) );
  INV_X1 U738 ( .A(G166), .ZN(G303) );
  XNOR2_X1 U739 ( .A(KEYINPUT19), .B(KEYINPUT82), .ZN(n655) );
  XNOR2_X1 U740 ( .A(G288), .B(KEYINPUT81), .ZN(n654) );
  XNOR2_X1 U741 ( .A(n655), .B(n654), .ZN(n658) );
  XOR2_X1 U742 ( .A(n664), .B(G305), .Z(n656) );
  XOR2_X1 U743 ( .A(n656), .B(n739), .Z(n657) );
  XNOR2_X1 U744 ( .A(n658), .B(n657), .ZN(n660) );
  XOR2_X1 U745 ( .A(G290), .B(G303), .Z(n659) );
  XNOR2_X1 U746 ( .A(n660), .B(n659), .ZN(n903) );
  XNOR2_X1 U747 ( .A(n903), .B(n661), .ZN(n662) );
  NOR2_X1 U748 ( .A1(n663), .A2(n662), .ZN(n666) );
  NOR2_X1 U749 ( .A1(G868), .A2(n664), .ZN(n665) );
  NOR2_X1 U750 ( .A1(n666), .A2(n665), .ZN(G295) );
  NAND2_X1 U751 ( .A1(G2078), .A2(G2084), .ZN(n667) );
  XOR2_X1 U752 ( .A(KEYINPUT20), .B(n667), .Z(n668) );
  NAND2_X1 U753 ( .A1(G2090), .A2(n668), .ZN(n669) );
  XNOR2_X1 U754 ( .A(KEYINPUT21), .B(n669), .ZN(n670) );
  NAND2_X1 U755 ( .A1(n670), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U756 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U757 ( .A1(G220), .A2(G219), .ZN(n671) );
  XOR2_X1 U758 ( .A(KEYINPUT22), .B(n671), .Z(n672) );
  NOR2_X1 U759 ( .A1(G218), .A2(n672), .ZN(n673) );
  NAND2_X1 U760 ( .A1(G96), .A2(n673), .ZN(n925) );
  NAND2_X1 U761 ( .A1(G2106), .A2(n925), .ZN(n677) );
  NAND2_X1 U762 ( .A1(G69), .A2(G120), .ZN(n674) );
  NOR2_X1 U763 ( .A1(G237), .A2(n674), .ZN(n675) );
  NAND2_X1 U764 ( .A1(G108), .A2(n675), .ZN(n926) );
  NAND2_X1 U765 ( .A1(G567), .A2(n926), .ZN(n676) );
  NAND2_X1 U766 ( .A1(n677), .A2(n676), .ZN(n838) );
  NAND2_X1 U767 ( .A1(G483), .A2(G661), .ZN(n678) );
  NOR2_X1 U768 ( .A1(n838), .A2(n678), .ZN(n837) );
  NAND2_X1 U769 ( .A1(n837), .A2(G36), .ZN(G176) );
  NAND2_X1 U770 ( .A1(G141), .A2(n882), .ZN(n680) );
  NAND2_X1 U771 ( .A1(G117), .A2(n885), .ZN(n679) );
  NAND2_X1 U772 ( .A1(n680), .A2(n679), .ZN(n683) );
  NAND2_X1 U773 ( .A1(n881), .A2(G105), .ZN(n681) );
  XOR2_X1 U774 ( .A(KEYINPUT38), .B(n681), .Z(n682) );
  NOR2_X1 U775 ( .A1(n683), .A2(n682), .ZN(n685) );
  NAND2_X1 U776 ( .A1(n886), .A2(G129), .ZN(n684) );
  NAND2_X1 U777 ( .A1(n685), .A2(n684), .ZN(n878) );
  NOR2_X1 U778 ( .A1(G1996), .A2(n878), .ZN(n939) );
  AND2_X1 U779 ( .A1(G40), .A2(n686), .ZN(n688) );
  NAND2_X1 U780 ( .A1(n688), .A2(n687), .ZN(n755) );
  NOR2_X1 U781 ( .A1(n718), .A2(n755), .ZN(n824) );
  NAND2_X1 U782 ( .A1(G95), .A2(n881), .ZN(n690) );
  NAND2_X1 U783 ( .A1(G131), .A2(n882), .ZN(n689) );
  NAND2_X1 U784 ( .A1(n690), .A2(n689), .ZN(n691) );
  XOR2_X1 U785 ( .A(KEYINPUT86), .B(n691), .Z(n695) );
  NAND2_X1 U786 ( .A1(G107), .A2(n885), .ZN(n693) );
  NAND2_X1 U787 ( .A1(G119), .A2(n886), .ZN(n692) );
  AND2_X1 U788 ( .A1(n693), .A2(n692), .ZN(n694) );
  NAND2_X1 U789 ( .A1(n695), .A2(n694), .ZN(n894) );
  NAND2_X1 U790 ( .A1(G1991), .A2(n894), .ZN(n697) );
  NAND2_X1 U791 ( .A1(G1996), .A2(n878), .ZN(n696) );
  NAND2_X1 U792 ( .A1(n697), .A2(n696), .ZN(n931) );
  NAND2_X1 U793 ( .A1(n824), .A2(n931), .ZN(n819) );
  NOR2_X1 U794 ( .A1(G1986), .A2(G290), .ZN(n698) );
  XOR2_X1 U795 ( .A(n698), .B(KEYINPUT102), .Z(n699) );
  OR2_X1 U796 ( .A1(n894), .A2(G1991), .ZN(n932) );
  NAND2_X1 U797 ( .A1(n699), .A2(n932), .ZN(n700) );
  NAND2_X1 U798 ( .A1(n819), .A2(n700), .ZN(n701) );
  XNOR2_X1 U799 ( .A(KEYINPUT103), .B(n701), .ZN(n702) );
  NOR2_X1 U800 ( .A1(n939), .A2(n702), .ZN(n703) );
  XNOR2_X1 U801 ( .A(n703), .B(KEYINPUT39), .ZN(n714) );
  NAND2_X1 U802 ( .A1(G104), .A2(n881), .ZN(n705) );
  NAND2_X1 U803 ( .A1(G140), .A2(n882), .ZN(n704) );
  NAND2_X1 U804 ( .A1(n705), .A2(n704), .ZN(n706) );
  XNOR2_X1 U805 ( .A(KEYINPUT34), .B(n706), .ZN(n712) );
  NAND2_X1 U806 ( .A1(n885), .A2(G116), .ZN(n707) );
  XOR2_X1 U807 ( .A(KEYINPUT85), .B(n707), .Z(n709) );
  NAND2_X1 U808 ( .A1(n886), .A2(G128), .ZN(n708) );
  NAND2_X1 U809 ( .A1(n709), .A2(n708), .ZN(n710) );
  XOR2_X1 U810 ( .A(KEYINPUT35), .B(n710), .Z(n711) );
  NOR2_X1 U811 ( .A1(n712), .A2(n711), .ZN(n713) );
  XNOR2_X1 U812 ( .A(KEYINPUT36), .B(n713), .ZN(n900) );
  INV_X1 U813 ( .A(G2067), .ZN(n842) );
  XOR2_X1 U814 ( .A(KEYINPUT37), .B(n842), .Z(n715) );
  NOR2_X1 U815 ( .A1(n900), .A2(n715), .ZN(n948) );
  NAND2_X1 U816 ( .A1(n824), .A2(n948), .ZN(n820) );
  NAND2_X1 U817 ( .A1(n714), .A2(n820), .ZN(n716) );
  NAND2_X1 U818 ( .A1(n900), .A2(n715), .ZN(n945) );
  NAND2_X1 U819 ( .A1(n716), .A2(n945), .ZN(n717) );
  NAND2_X1 U820 ( .A1(n717), .A2(n824), .ZN(n830) );
  INV_X1 U821 ( .A(n718), .ZN(n757) );
  OR2_X1 U822 ( .A1(n755), .A2(n757), .ZN(n773) );
  NAND2_X1 U823 ( .A1(n773), .A2(G1341), .ZN(n719) );
  XNOR2_X1 U824 ( .A(n719), .B(KEYINPUT92), .ZN(n720) );
  NAND2_X1 U825 ( .A1(n720), .A2(n962), .ZN(n723) );
  NAND2_X1 U826 ( .A1(G1996), .A2(n760), .ZN(n721) );
  XOR2_X1 U827 ( .A(KEYINPUT26), .B(n721), .Z(n722) );
  NOR2_X1 U828 ( .A1(n723), .A2(n722), .ZN(n725) );
  OR2_X1 U829 ( .A1(n725), .A2(n724), .ZN(n732) );
  NAND2_X1 U830 ( .A1(n725), .A2(n724), .ZN(n730) );
  NOR2_X1 U831 ( .A1(n773), .A2(n842), .ZN(n726) );
  XNOR2_X1 U832 ( .A(n726), .B(KEYINPUT93), .ZN(n728) );
  NAND2_X1 U833 ( .A1(n773), .A2(G1348), .ZN(n727) );
  NAND2_X1 U834 ( .A1(n728), .A2(n727), .ZN(n729) );
  NAND2_X1 U835 ( .A1(n730), .A2(n729), .ZN(n731) );
  NAND2_X1 U836 ( .A1(n732), .A2(n731), .ZN(n738) );
  NAND2_X1 U837 ( .A1(n748), .A2(G2072), .ZN(n734) );
  INV_X1 U838 ( .A(G1956), .ZN(n854) );
  NOR2_X1 U839 ( .A1(n748), .A2(n854), .ZN(n735) );
  NOR2_X1 U840 ( .A1(n736), .A2(n735), .ZN(n740) );
  NAND2_X1 U841 ( .A1(n739), .A2(n740), .ZN(n737) );
  NAND2_X1 U842 ( .A1(n738), .A2(n737), .ZN(n744) );
  NOR2_X1 U843 ( .A1(n740), .A2(n739), .ZN(n742) );
  XNOR2_X1 U844 ( .A(KEYINPUT91), .B(KEYINPUT28), .ZN(n741) );
  XNOR2_X1 U845 ( .A(n742), .B(n741), .ZN(n743) );
  NAND2_X1 U846 ( .A1(n744), .A2(n743), .ZN(n746) );
  XOR2_X1 U847 ( .A(KEYINPUT94), .B(KEYINPUT29), .Z(n745) );
  XNOR2_X1 U848 ( .A(n746), .B(n745), .ZN(n754) );
  XNOR2_X1 U849 ( .A(G2078), .B(KEYINPUT25), .ZN(n1007) );
  NAND2_X1 U850 ( .A1(n760), .A2(n1007), .ZN(n747) );
  XNOR2_X1 U851 ( .A(n747), .B(KEYINPUT87), .ZN(n750) );
  NOR2_X1 U852 ( .A1(n748), .A2(G1961), .ZN(n749) );
  NOR2_X1 U853 ( .A1(n750), .A2(n749), .ZN(n751) );
  XNOR2_X1 U854 ( .A(KEYINPUT88), .B(n751), .ZN(n766) );
  NOR2_X1 U855 ( .A1(G301), .A2(n766), .ZN(n752) );
  XNOR2_X1 U856 ( .A(KEYINPUT89), .B(n752), .ZN(n753) );
  NAND2_X1 U857 ( .A1(n754), .A2(n753), .ZN(n772) );
  XOR2_X1 U858 ( .A(KEYINPUT30), .B(KEYINPUT96), .Z(n765) );
  OR2_X1 U859 ( .A1(n755), .A2(G2084), .ZN(n756) );
  NOR2_X1 U860 ( .A1(n757), .A2(n756), .ZN(n787) );
  INV_X1 U861 ( .A(G8), .ZN(n758) );
  OR2_X1 U862 ( .A1(n758), .A2(G1966), .ZN(n759) );
  NOR2_X1 U863 ( .A1(n760), .A2(n759), .ZN(n784) );
  NOR2_X1 U864 ( .A1(n787), .A2(n784), .ZN(n762) );
  XNOR2_X1 U865 ( .A(n762), .B(n761), .ZN(n763) );
  NAND2_X1 U866 ( .A1(n763), .A2(G8), .ZN(n764) );
  NOR2_X1 U867 ( .A1(G168), .A2(n519), .ZN(n768) );
  AND2_X1 U868 ( .A1(G301), .A2(n766), .ZN(n767) );
  NOR2_X1 U869 ( .A1(n768), .A2(n767), .ZN(n769) );
  XNOR2_X1 U870 ( .A(KEYINPUT31), .B(n769), .ZN(n770) );
  INV_X1 U871 ( .A(n770), .ZN(n771) );
  NAND2_X1 U872 ( .A1(n772), .A2(n771), .ZN(n785) );
  NAND2_X1 U873 ( .A1(n785), .A2(G286), .ZN(n780) );
  AND2_X1 U874 ( .A1(G8), .A2(n773), .ZN(n793) );
  INV_X1 U875 ( .A(n793), .ZN(n817) );
  NOR2_X1 U876 ( .A1(G1971), .A2(n817), .ZN(n774) );
  XNOR2_X1 U877 ( .A(KEYINPUT97), .B(n774), .ZN(n777) );
  NOR2_X1 U878 ( .A1(G2090), .A2(n773), .ZN(n775) );
  NOR2_X1 U879 ( .A1(G166), .A2(n775), .ZN(n776) );
  NAND2_X1 U880 ( .A1(n777), .A2(n776), .ZN(n778) );
  OR2_X1 U881 ( .A1(n758), .A2(n778), .ZN(n779) );
  NAND2_X1 U882 ( .A1(n780), .A2(n779), .ZN(n782) );
  INV_X1 U883 ( .A(KEYINPUT32), .ZN(n781) );
  XNOR2_X1 U884 ( .A(n782), .B(n781), .ZN(n806) );
  INV_X1 U885 ( .A(KEYINPUT33), .ZN(n783) );
  AND2_X1 U886 ( .A1(n806), .A2(n783), .ZN(n791) );
  INV_X1 U887 ( .A(n785), .ZN(n786) );
  NOR2_X1 U888 ( .A1(n784), .A2(n786), .ZN(n789) );
  NAND2_X1 U889 ( .A1(G8), .A2(n787), .ZN(n788) );
  NAND2_X1 U890 ( .A1(n789), .A2(n788), .ZN(n807) );
  NAND2_X1 U891 ( .A1(G1976), .A2(G288), .ZN(n960) );
  AND2_X1 U892 ( .A1(n807), .A2(n960), .ZN(n790) );
  NAND2_X1 U893 ( .A1(n791), .A2(n790), .ZN(n803) );
  NOR2_X1 U894 ( .A1(G1976), .A2(G288), .ZN(n796) );
  NAND2_X1 U895 ( .A1(n796), .A2(n793), .ZN(n792) );
  NAND2_X1 U896 ( .A1(n792), .A2(KEYINPUT33), .ZN(n799) );
  INV_X1 U897 ( .A(n799), .ZN(n794) );
  INV_X1 U898 ( .A(n960), .ZN(n797) );
  NOR2_X1 U899 ( .A1(G1971), .A2(G303), .ZN(n795) );
  NOR2_X1 U900 ( .A1(n796), .A2(n795), .ZN(n963) );
  OR2_X1 U901 ( .A1(n797), .A2(n963), .ZN(n798) );
  OR2_X1 U902 ( .A1(KEYINPUT33), .A2(n798), .ZN(n800) );
  AND2_X1 U903 ( .A1(n800), .A2(n799), .ZN(n801) );
  OR2_X1 U904 ( .A1(n520), .A2(n801), .ZN(n802) );
  NAND2_X1 U905 ( .A1(n803), .A2(n802), .ZN(n804) );
  XNOR2_X1 U906 ( .A(n804), .B(KEYINPUT98), .ZN(n805) );
  XOR2_X1 U907 ( .A(G1981), .B(G305), .Z(n953) );
  NAND2_X1 U908 ( .A1(n805), .A2(n953), .ZN(n813) );
  NAND2_X1 U909 ( .A1(n806), .A2(n807), .ZN(n810) );
  NOR2_X1 U910 ( .A1(G2090), .A2(G303), .ZN(n808) );
  NAND2_X1 U911 ( .A1(G8), .A2(n808), .ZN(n809) );
  NAND2_X1 U912 ( .A1(n810), .A2(n809), .ZN(n811) );
  NAND2_X1 U913 ( .A1(n811), .A2(n817), .ZN(n812) );
  NAND2_X1 U914 ( .A1(n813), .A2(n812), .ZN(n814) );
  NOR2_X1 U915 ( .A1(G1981), .A2(G305), .ZN(n815) );
  XOR2_X1 U916 ( .A(n815), .B(KEYINPUT24), .Z(n816) );
  NAND2_X1 U917 ( .A1(n820), .A2(n819), .ZN(n821) );
  XNOR2_X1 U918 ( .A(n823), .B(KEYINPUT100), .ZN(n826) );
  XNOR2_X1 U919 ( .A(G1986), .B(G290), .ZN(n959) );
  NAND2_X1 U920 ( .A1(n824), .A2(n959), .ZN(n825) );
  NAND2_X1 U921 ( .A1(n826), .A2(n825), .ZN(n828) );
  NAND2_X1 U922 ( .A1(n830), .A2(n829), .ZN(n831) );
  XNOR2_X1 U923 ( .A(n831), .B(KEYINPUT40), .ZN(G329) );
  NAND2_X1 U924 ( .A1(G2106), .A2(n832), .ZN(G217) );
  INV_X1 U925 ( .A(n832), .ZN(G223) );
  NAND2_X1 U926 ( .A1(G15), .A2(G2), .ZN(n833) );
  XNOR2_X1 U927 ( .A(KEYINPUT105), .B(n833), .ZN(n834) );
  NAND2_X1 U928 ( .A1(n834), .A2(G661), .ZN(n835) );
  XNOR2_X1 U929 ( .A(KEYINPUT106), .B(n835), .ZN(G259) );
  NAND2_X1 U930 ( .A1(G3), .A2(G1), .ZN(n836) );
  NAND2_X1 U931 ( .A1(n837), .A2(n836), .ZN(G188) );
  XNOR2_X1 U932 ( .A(KEYINPUT107), .B(n838), .ZN(G319) );
  XOR2_X1 U933 ( .A(G2096), .B(KEYINPUT108), .Z(n840) );
  XNOR2_X1 U934 ( .A(G2090), .B(KEYINPUT43), .ZN(n839) );
  XNOR2_X1 U935 ( .A(n840), .B(n839), .ZN(n841) );
  XOR2_X1 U936 ( .A(n841), .B(KEYINPUT42), .Z(n844) );
  XOR2_X1 U937 ( .A(n842), .B(G2072), .Z(n843) );
  XNOR2_X1 U938 ( .A(n844), .B(n843), .ZN(n848) );
  XOR2_X1 U939 ( .A(G2678), .B(G2100), .Z(n846) );
  XNOR2_X1 U940 ( .A(G2078), .B(G2084), .ZN(n845) );
  XNOR2_X1 U941 ( .A(n846), .B(n845), .ZN(n847) );
  XNOR2_X1 U942 ( .A(n848), .B(n847), .ZN(G227) );
  XOR2_X1 U943 ( .A(G1966), .B(G1971), .Z(n850) );
  XNOR2_X1 U944 ( .A(G1981), .B(G1976), .ZN(n849) );
  XNOR2_X1 U945 ( .A(n850), .B(n849), .ZN(n851) );
  XOR2_X1 U946 ( .A(n851), .B(G2474), .Z(n853) );
  XNOR2_X1 U947 ( .A(G1996), .B(G1991), .ZN(n852) );
  XNOR2_X1 U948 ( .A(n853), .B(n852), .ZN(n858) );
  XOR2_X1 U949 ( .A(KEYINPUT41), .B(G1961), .Z(n856) );
  XOR2_X1 U950 ( .A(G1986), .B(n854), .Z(n855) );
  XNOR2_X1 U951 ( .A(n856), .B(n855), .ZN(n857) );
  XNOR2_X1 U952 ( .A(n858), .B(n857), .ZN(G229) );
  NAND2_X1 U953 ( .A1(G100), .A2(n881), .ZN(n860) );
  NAND2_X1 U954 ( .A1(G136), .A2(n882), .ZN(n859) );
  NAND2_X1 U955 ( .A1(n860), .A2(n859), .ZN(n863) );
  NAND2_X1 U956 ( .A1(n885), .A2(G112), .ZN(n861) );
  XOR2_X1 U957 ( .A(KEYINPUT110), .B(n861), .Z(n862) );
  NOR2_X1 U958 ( .A1(n863), .A2(n862), .ZN(n867) );
  XOR2_X1 U959 ( .A(KEYINPUT44), .B(KEYINPUT109), .Z(n865) );
  NAND2_X1 U960 ( .A1(G124), .A2(n886), .ZN(n864) );
  XNOR2_X1 U961 ( .A(n865), .B(n864), .ZN(n866) );
  NAND2_X1 U962 ( .A1(n867), .A2(n866), .ZN(n868) );
  XNOR2_X1 U963 ( .A(n868), .B(KEYINPUT111), .ZN(G162) );
  XNOR2_X1 U964 ( .A(KEYINPUT46), .B(KEYINPUT48), .ZN(n880) );
  NAND2_X1 U965 ( .A1(G106), .A2(n881), .ZN(n870) );
  NAND2_X1 U966 ( .A1(G142), .A2(n882), .ZN(n869) );
  NAND2_X1 U967 ( .A1(n870), .A2(n869), .ZN(n871) );
  XNOR2_X1 U968 ( .A(n871), .B(KEYINPUT45), .ZN(n873) );
  NAND2_X1 U969 ( .A1(G130), .A2(n886), .ZN(n872) );
  NAND2_X1 U970 ( .A1(n873), .A2(n872), .ZN(n876) );
  NAND2_X1 U971 ( .A1(n885), .A2(G118), .ZN(n874) );
  XOR2_X1 U972 ( .A(KEYINPUT112), .B(n874), .Z(n875) );
  NOR2_X1 U973 ( .A1(n876), .A2(n875), .ZN(n877) );
  XNOR2_X1 U974 ( .A(n878), .B(n877), .ZN(n879) );
  XNOR2_X1 U975 ( .A(n880), .B(n879), .ZN(n893) );
  NAND2_X1 U976 ( .A1(G103), .A2(n881), .ZN(n884) );
  NAND2_X1 U977 ( .A1(G139), .A2(n882), .ZN(n883) );
  NAND2_X1 U978 ( .A1(n884), .A2(n883), .ZN(n892) );
  NAND2_X1 U979 ( .A1(G115), .A2(n885), .ZN(n888) );
  NAND2_X1 U980 ( .A1(G127), .A2(n886), .ZN(n887) );
  NAND2_X1 U981 ( .A1(n888), .A2(n887), .ZN(n889) );
  XNOR2_X1 U982 ( .A(KEYINPUT113), .B(n889), .ZN(n890) );
  XNOR2_X1 U983 ( .A(KEYINPUT47), .B(n890), .ZN(n891) );
  NOR2_X1 U984 ( .A1(n892), .A2(n891), .ZN(n934) );
  XOR2_X1 U985 ( .A(n893), .B(n934), .Z(n896) );
  XOR2_X1 U986 ( .A(G164), .B(n894), .Z(n895) );
  XNOR2_X1 U987 ( .A(n896), .B(n895), .ZN(n897) );
  XNOR2_X1 U988 ( .A(n928), .B(n897), .ZN(n899) );
  XNOR2_X1 U989 ( .A(G160), .B(G162), .ZN(n898) );
  XNOR2_X1 U990 ( .A(n899), .B(n898), .ZN(n901) );
  XOR2_X1 U991 ( .A(n901), .B(n900), .Z(n902) );
  NOR2_X1 U992 ( .A1(G37), .A2(n902), .ZN(G395) );
  XOR2_X1 U993 ( .A(n903), .B(G286), .Z(n905) );
  XOR2_X1 U994 ( .A(n965), .B(G171), .Z(n904) );
  XNOR2_X1 U995 ( .A(n905), .B(n904), .ZN(n906) );
  XOR2_X1 U996 ( .A(n962), .B(n906), .Z(n907) );
  NOR2_X1 U997 ( .A1(G37), .A2(n907), .ZN(n908) );
  XNOR2_X1 U998 ( .A(KEYINPUT114), .B(n908), .ZN(G397) );
  XNOR2_X1 U999 ( .A(G1341), .B(G2454), .ZN(n909) );
  XNOR2_X1 U1000 ( .A(n909), .B(G2430), .ZN(n910) );
  XNOR2_X1 U1001 ( .A(n910), .B(G1348), .ZN(n916) );
  XOR2_X1 U1002 ( .A(G2443), .B(G2427), .Z(n912) );
  XNOR2_X1 U1003 ( .A(G2438), .B(G2446), .ZN(n911) );
  XNOR2_X1 U1004 ( .A(n912), .B(n911), .ZN(n914) );
  XOR2_X1 U1005 ( .A(G2451), .B(G2435), .Z(n913) );
  XNOR2_X1 U1006 ( .A(n914), .B(n913), .ZN(n915) );
  XNOR2_X1 U1007 ( .A(n916), .B(n915), .ZN(n917) );
  NAND2_X1 U1008 ( .A1(n917), .A2(G14), .ZN(n918) );
  XNOR2_X1 U1009 ( .A(KEYINPUT104), .B(n918), .ZN(n927) );
  NAND2_X1 U1010 ( .A1(G319), .A2(n927), .ZN(n922) );
  NOR2_X1 U1011 ( .A1(G227), .A2(G229), .ZN(n919) );
  XOR2_X1 U1012 ( .A(KEYINPUT49), .B(n919), .Z(n920) );
  XNOR2_X1 U1013 ( .A(n920), .B(KEYINPUT115), .ZN(n921) );
  NOR2_X1 U1014 ( .A1(n922), .A2(n921), .ZN(n924) );
  NOR2_X1 U1015 ( .A1(G395), .A2(G397), .ZN(n923) );
  NAND2_X1 U1016 ( .A1(n924), .A2(n923), .ZN(G225) );
  XOR2_X1 U1017 ( .A(KEYINPUT116), .B(G225), .Z(G308) );
  INV_X1 U1019 ( .A(G120), .ZN(G236) );
  INV_X1 U1020 ( .A(G96), .ZN(G221) );
  INV_X1 U1021 ( .A(G69), .ZN(G235) );
  NOR2_X1 U1022 ( .A1(n926), .A2(n925), .ZN(G325) );
  INV_X1 U1023 ( .A(G325), .ZN(G261) );
  INV_X1 U1024 ( .A(n927), .ZN(G401) );
  INV_X1 U1025 ( .A(G108), .ZN(G238) );
  INV_X1 U1026 ( .A(G29), .ZN(n1024) );
  XNOR2_X1 U1027 ( .A(KEYINPUT117), .B(KEYINPUT52), .ZN(n950) );
  XNOR2_X1 U1028 ( .A(G160), .B(G2084), .ZN(n929) );
  NAND2_X1 U1029 ( .A1(n929), .A2(n928), .ZN(n930) );
  NOR2_X1 U1030 ( .A1(n931), .A2(n930), .ZN(n933) );
  NAND2_X1 U1031 ( .A1(n933), .A2(n932), .ZN(n944) );
  XOR2_X1 U1032 ( .A(G2072), .B(n934), .Z(n936) );
  XOR2_X1 U1033 ( .A(G164), .B(G2078), .Z(n935) );
  NOR2_X1 U1034 ( .A1(n936), .A2(n935), .ZN(n937) );
  XNOR2_X1 U1035 ( .A(KEYINPUT50), .B(n937), .ZN(n942) );
  XOR2_X1 U1036 ( .A(G2090), .B(G162), .Z(n938) );
  NOR2_X1 U1037 ( .A1(n939), .A2(n938), .ZN(n940) );
  XOR2_X1 U1038 ( .A(KEYINPUT51), .B(n940), .Z(n941) );
  NAND2_X1 U1039 ( .A1(n942), .A2(n941), .ZN(n943) );
  NOR2_X1 U1040 ( .A1(n944), .A2(n943), .ZN(n946) );
  NAND2_X1 U1041 ( .A1(n946), .A2(n945), .ZN(n947) );
  NOR2_X1 U1042 ( .A1(n948), .A2(n947), .ZN(n949) );
  XNOR2_X1 U1043 ( .A(n950), .B(n949), .ZN(n951) );
  XNOR2_X1 U1044 ( .A(KEYINPUT55), .B(KEYINPUT118), .ZN(n1022) );
  NOR2_X1 U1045 ( .A1(n951), .A2(n1022), .ZN(n952) );
  NOR2_X1 U1046 ( .A1(n1024), .A2(n952), .ZN(n1033) );
  INV_X1 U1047 ( .A(G16), .ZN(n998) );
  XOR2_X1 U1048 ( .A(n998), .B(KEYINPUT56), .Z(n975) );
  XNOR2_X1 U1049 ( .A(G1966), .B(G168), .ZN(n954) );
  NAND2_X1 U1050 ( .A1(n954), .A2(n953), .ZN(n955) );
  XNOR2_X1 U1051 ( .A(n955), .B(KEYINPUT57), .ZN(n973) );
  XOR2_X1 U1052 ( .A(G1961), .B(G301), .Z(n957) );
  NAND2_X1 U1053 ( .A1(G1971), .A2(G303), .ZN(n956) );
  NAND2_X1 U1054 ( .A1(n957), .A2(n956), .ZN(n958) );
  NOR2_X1 U1055 ( .A1(n959), .A2(n958), .ZN(n961) );
  NAND2_X1 U1056 ( .A1(n961), .A2(n960), .ZN(n971) );
  XNOR2_X1 U1057 ( .A(n962), .B(G1341), .ZN(n969) );
  XOR2_X1 U1058 ( .A(G299), .B(G1956), .Z(n964) );
  NAND2_X1 U1059 ( .A1(n964), .A2(n963), .ZN(n967) );
  XNOR2_X1 U1060 ( .A(G1348), .B(n965), .ZN(n966) );
  NOR2_X1 U1061 ( .A1(n967), .A2(n966), .ZN(n968) );
  NAND2_X1 U1062 ( .A1(n969), .A2(n968), .ZN(n970) );
  NOR2_X1 U1063 ( .A1(n971), .A2(n970), .ZN(n972) );
  NAND2_X1 U1064 ( .A1(n973), .A2(n972), .ZN(n974) );
  NAND2_X1 U1065 ( .A1(n975), .A2(n974), .ZN(n1000) );
  XNOR2_X1 U1066 ( .A(G1981), .B(G6), .ZN(n977) );
  XNOR2_X1 U1067 ( .A(G1341), .B(G19), .ZN(n976) );
  NOR2_X1 U1068 ( .A1(n977), .A2(n976), .ZN(n978) );
  XNOR2_X1 U1069 ( .A(KEYINPUT126), .B(n978), .ZN(n980) );
  XOR2_X1 U1070 ( .A(G1956), .B(G20), .Z(n979) );
  NAND2_X1 U1071 ( .A1(n980), .A2(n979), .ZN(n983) );
  XOR2_X1 U1072 ( .A(KEYINPUT59), .B(G1348), .Z(n981) );
  XNOR2_X1 U1073 ( .A(G4), .B(n981), .ZN(n982) );
  NOR2_X1 U1074 ( .A1(n983), .A2(n982), .ZN(n984) );
  XNOR2_X1 U1075 ( .A(KEYINPUT60), .B(n984), .ZN(n988) );
  XNOR2_X1 U1076 ( .A(G1966), .B(G21), .ZN(n986) );
  XNOR2_X1 U1077 ( .A(G1961), .B(G5), .ZN(n985) );
  NOR2_X1 U1078 ( .A1(n986), .A2(n985), .ZN(n987) );
  NAND2_X1 U1079 ( .A1(n988), .A2(n987), .ZN(n995) );
  XNOR2_X1 U1080 ( .A(G1986), .B(G24), .ZN(n990) );
  XNOR2_X1 U1081 ( .A(G1971), .B(G22), .ZN(n989) );
  NOR2_X1 U1082 ( .A1(n990), .A2(n989), .ZN(n992) );
  XOR2_X1 U1083 ( .A(G1976), .B(G23), .Z(n991) );
  NAND2_X1 U1084 ( .A1(n992), .A2(n991), .ZN(n993) );
  XNOR2_X1 U1085 ( .A(KEYINPUT58), .B(n993), .ZN(n994) );
  NOR2_X1 U1086 ( .A1(n995), .A2(n994), .ZN(n996) );
  XNOR2_X1 U1087 ( .A(KEYINPUT61), .B(n996), .ZN(n997) );
  NAND2_X1 U1088 ( .A1(n998), .A2(n997), .ZN(n999) );
  NAND2_X1 U1089 ( .A1(n1000), .A2(n999), .ZN(n1030) );
  XOR2_X1 U1090 ( .A(G25), .B(G1991), .Z(n1006) );
  XOR2_X1 U1091 ( .A(G26), .B(G2067), .Z(n1001) );
  NAND2_X1 U1092 ( .A1(n1001), .A2(G28), .ZN(n1004) );
  XNOR2_X1 U1093 ( .A(KEYINPUT120), .B(G2072), .ZN(n1002) );
  XNOR2_X1 U1094 ( .A(G33), .B(n1002), .ZN(n1003) );
  NOR2_X1 U1095 ( .A1(n1004), .A2(n1003), .ZN(n1005) );
  NAND2_X1 U1096 ( .A1(n1006), .A2(n1005), .ZN(n1012) );
  XOR2_X1 U1097 ( .A(G1996), .B(G32), .Z(n1009) );
  XNOR2_X1 U1098 ( .A(n1007), .B(G27), .ZN(n1008) );
  NAND2_X1 U1099 ( .A1(n1009), .A2(n1008), .ZN(n1010) );
  XOR2_X1 U1100 ( .A(n1010), .B(KEYINPUT121), .Z(n1011) );
  NOR2_X1 U1101 ( .A1(n1012), .A2(n1011), .ZN(n1013) );
  XOR2_X1 U1102 ( .A(KEYINPUT122), .B(n1013), .Z(n1014) );
  XNOR2_X1 U1103 ( .A(KEYINPUT53), .B(n1014), .ZN(n1017) );
  XNOR2_X1 U1104 ( .A(G2090), .B(G35), .ZN(n1015) );
  XNOR2_X1 U1105 ( .A(n1015), .B(KEYINPUT119), .ZN(n1016) );
  NAND2_X1 U1106 ( .A1(n1017), .A2(n1016), .ZN(n1018) );
  XNOR2_X1 U1107 ( .A(n1018), .B(KEYINPUT123), .ZN(n1021) );
  XOR2_X1 U1108 ( .A(G2084), .B(G34), .Z(n1019) );
  XNOR2_X1 U1109 ( .A(KEYINPUT54), .B(n1019), .ZN(n1020) );
  NAND2_X1 U1110 ( .A1(n1021), .A2(n1020), .ZN(n1023) );
  XOR2_X1 U1111 ( .A(n1023), .B(n1022), .Z(n1026) );
  XNOR2_X1 U1112 ( .A(n1024), .B(KEYINPUT124), .ZN(n1025) );
  NAND2_X1 U1113 ( .A1(n1026), .A2(n1025), .ZN(n1027) );
  NAND2_X1 U1114 ( .A1(n1027), .A2(G11), .ZN(n1028) );
  XOR2_X1 U1115 ( .A(KEYINPUT125), .B(n1028), .Z(n1029) );
  NOR2_X1 U1116 ( .A1(n1030), .A2(n1029), .ZN(n1031) );
  XNOR2_X1 U1117 ( .A(n1031), .B(KEYINPUT127), .ZN(n1032) );
  NOR2_X1 U1118 ( .A1(n1033), .A2(n1032), .ZN(n1034) );
  XOR2_X1 U1119 ( .A(KEYINPUT62), .B(n1034), .Z(G150) );
  INV_X1 U1120 ( .A(G150), .ZN(G311) );
endmodule

