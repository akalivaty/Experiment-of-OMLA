//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 0 0 0 1 1 1 0 0 0 0 1 0 1 1 0 1 1 1 1 0 1 0 0 0 1 0 1 1 0 0 0 0 0 1 0 0 0 0 0 1 1 1 1 0 0 1 1 1 1 1 1 0 1 0 0 1 0 1 1 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:15:15 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n679, new_n680,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n709, new_n710,
    new_n711, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n728, new_n729, new_n730, new_n731, new_n733, new_n734, new_n735,
    new_n736, new_n737, new_n739, new_n740, new_n741, new_n742, new_n744,
    new_n745, new_n747, new_n748, new_n749, new_n750, new_n751, new_n752,
    new_n753, new_n754, new_n755, new_n756, new_n757, new_n758, new_n759,
    new_n760, new_n761, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n774, new_n775,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n847, new_n848,
    new_n849, new_n851, new_n852, new_n853, new_n855, new_n856, new_n857,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n901, new_n902,
    new_n903, new_n904, new_n906, new_n907, new_n908, new_n909, new_n910,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n923, new_n924, new_n925, new_n927,
    new_n928, new_n929, new_n930, new_n931, new_n932, new_n933, new_n935,
    new_n936, new_n937, new_n938, new_n939, new_n940, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n948, new_n949, new_n950,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n960, new_n961, new_n962, new_n963, new_n964, new_n965, new_n966,
    new_n967, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976;
  INV_X1    g000(.A(KEYINPUT72), .ZN(new_n202));
  NAND2_X1  g001(.A1(G227gat), .A2(G233gat), .ZN(new_n203));
  XOR2_X1   g002(.A(new_n203), .B(KEYINPUT64), .Z(new_n204));
  INV_X1    g003(.A(G120gat), .ZN(new_n205));
  NAND2_X1  g004(.A1(new_n205), .A2(G113gat), .ZN(new_n206));
  INV_X1    g005(.A(G113gat), .ZN(new_n207));
  NAND2_X1  g006(.A1(new_n207), .A2(G120gat), .ZN(new_n208));
  AOI21_X1  g007(.A(KEYINPUT1), .B1(new_n206), .B2(new_n208), .ZN(new_n209));
  XNOR2_X1  g008(.A(G127gat), .B(G134gat), .ZN(new_n210));
  NAND2_X1  g009(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  INV_X1    g010(.A(G134gat), .ZN(new_n212));
  NAND2_X1  g011(.A1(new_n212), .A2(G127gat), .ZN(new_n213));
  INV_X1    g012(.A(G127gat), .ZN(new_n214));
  NAND2_X1  g013(.A1(new_n214), .A2(G134gat), .ZN(new_n215));
  AND3_X1   g014(.A1(new_n213), .A2(new_n215), .A3(KEYINPUT67), .ZN(new_n216));
  AOI21_X1  g015(.A(KEYINPUT67), .B1(new_n213), .B2(new_n215), .ZN(new_n217));
  AND2_X1   g016(.A1(new_n206), .A2(new_n208), .ZN(new_n218));
  OAI22_X1  g017(.A1(new_n216), .A2(new_n217), .B1(new_n218), .B2(KEYINPUT1), .ZN(new_n219));
  OAI21_X1  g018(.A(new_n211), .B1(new_n219), .B2(KEYINPUT68), .ZN(new_n220));
  NAND2_X1  g019(.A1(new_n210), .A2(KEYINPUT67), .ZN(new_n221));
  INV_X1    g020(.A(KEYINPUT67), .ZN(new_n222));
  NOR2_X1   g021(.A1(new_n214), .A2(G134gat), .ZN(new_n223));
  NOR2_X1   g022(.A1(new_n212), .A2(G127gat), .ZN(new_n224));
  OAI21_X1  g023(.A(new_n222), .B1(new_n223), .B2(new_n224), .ZN(new_n225));
  AOI21_X1  g024(.A(new_n209), .B1(new_n221), .B2(new_n225), .ZN(new_n226));
  INV_X1    g025(.A(KEYINPUT68), .ZN(new_n227));
  NOR2_X1   g026(.A1(new_n226), .A2(new_n227), .ZN(new_n228));
  OAI21_X1  g027(.A(KEYINPUT69), .B1(new_n220), .B2(new_n228), .ZN(new_n229));
  AOI22_X1  g028(.A1(new_n226), .A2(new_n227), .B1(new_n209), .B2(new_n210), .ZN(new_n230));
  INV_X1    g029(.A(KEYINPUT69), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n219), .A2(KEYINPUT68), .ZN(new_n232));
  NAND3_X1  g031(.A1(new_n230), .A2(new_n231), .A3(new_n232), .ZN(new_n233));
  NAND2_X1  g032(.A1(G169gat), .A2(G176gat), .ZN(new_n234));
  INV_X1    g033(.A(new_n234), .ZN(new_n235));
  NOR2_X1   g034(.A1(G169gat), .A2(G176gat), .ZN(new_n236));
  AOI21_X1  g035(.A(new_n235), .B1(KEYINPUT23), .B2(new_n236), .ZN(new_n237));
  XNOR2_X1  g036(.A(new_n237), .B(KEYINPUT66), .ZN(new_n238));
  INV_X1    g037(.A(G183gat), .ZN(new_n239));
  INV_X1    g038(.A(G190gat), .ZN(new_n240));
  NOR3_X1   g039(.A1(new_n239), .A2(new_n240), .A3(KEYINPUT24), .ZN(new_n241));
  XOR2_X1   g040(.A(G183gat), .B(G190gat), .Z(new_n242));
  AOI21_X1  g041(.A(new_n241), .B1(new_n242), .B2(KEYINPUT24), .ZN(new_n243));
  INV_X1    g042(.A(KEYINPUT23), .ZN(new_n244));
  OAI21_X1  g043(.A(new_n244), .B1(G169gat), .B2(G176gat), .ZN(new_n245));
  NAND2_X1  g044(.A1(new_n243), .A2(new_n245), .ZN(new_n246));
  OAI21_X1  g045(.A(KEYINPUT25), .B1(new_n238), .B2(new_n246), .ZN(new_n247));
  INV_X1    g046(.A(KEYINPUT28), .ZN(new_n248));
  XNOR2_X1  g047(.A(KEYINPUT27), .B(G183gat), .ZN(new_n249));
  INV_X1    g048(.A(new_n249), .ZN(new_n250));
  OAI21_X1  g049(.A(new_n248), .B1(new_n250), .B2(G190gat), .ZN(new_n251));
  NAND3_X1  g050(.A1(new_n249), .A2(KEYINPUT28), .A3(new_n240), .ZN(new_n252));
  NAND2_X1  g051(.A1(new_n251), .A2(new_n252), .ZN(new_n253));
  INV_X1    g052(.A(new_n236), .ZN(new_n254));
  OR2_X1    g053(.A1(new_n254), .A2(KEYINPUT26), .ZN(new_n255));
  AOI21_X1  g054(.A(new_n235), .B1(new_n254), .B2(KEYINPUT26), .ZN(new_n256));
  AOI22_X1  g055(.A1(new_n255), .A2(new_n256), .B1(G183gat), .B2(G190gat), .ZN(new_n257));
  INV_X1    g056(.A(KEYINPUT25), .ZN(new_n258));
  NAND3_X1  g057(.A1(new_n245), .A2(new_n258), .A3(new_n234), .ZN(new_n259));
  XNOR2_X1  g058(.A(KEYINPUT65), .B(G169gat), .ZN(new_n260));
  NOR2_X1   g059(.A1(new_n244), .A2(G176gat), .ZN(new_n261));
  AOI21_X1  g060(.A(new_n259), .B1(new_n260), .B2(new_n261), .ZN(new_n262));
  AOI22_X1  g061(.A1(new_n253), .A2(new_n257), .B1(new_n243), .B2(new_n262), .ZN(new_n263));
  AND4_X1   g062(.A1(new_n229), .A2(new_n233), .A3(new_n247), .A4(new_n263), .ZN(new_n264));
  AOI22_X1  g063(.A1(new_n229), .A2(new_n233), .B1(new_n247), .B2(new_n263), .ZN(new_n265));
  OAI21_X1  g064(.A(new_n204), .B1(new_n264), .B2(new_n265), .ZN(new_n266));
  NAND2_X1  g065(.A1(new_n266), .A2(KEYINPUT32), .ZN(new_n267));
  XNOR2_X1  g066(.A(G15gat), .B(G43gat), .ZN(new_n268));
  XNOR2_X1  g067(.A(G71gat), .B(G99gat), .ZN(new_n269));
  XNOR2_X1  g068(.A(new_n268), .B(new_n269), .ZN(new_n270));
  INV_X1    g069(.A(KEYINPUT33), .ZN(new_n271));
  NOR2_X1   g070(.A1(new_n270), .A2(new_n271), .ZN(new_n272));
  NOR2_X1   g071(.A1(new_n267), .A2(new_n272), .ZN(new_n273));
  NOR2_X1   g072(.A1(new_n264), .A2(new_n265), .ZN(new_n274));
  INV_X1    g073(.A(KEYINPUT34), .ZN(new_n275));
  INV_X1    g074(.A(new_n204), .ZN(new_n276));
  NAND4_X1  g075(.A1(new_n274), .A2(KEYINPUT71), .A3(new_n275), .A4(new_n276), .ZN(new_n277));
  INV_X1    g076(.A(KEYINPUT71), .ZN(new_n278));
  NAND2_X1  g077(.A1(new_n247), .A2(new_n263), .ZN(new_n279));
  NOR3_X1   g078(.A1(new_n220), .A2(new_n228), .A3(KEYINPUT69), .ZN(new_n280));
  AOI21_X1  g079(.A(new_n231), .B1(new_n230), .B2(new_n232), .ZN(new_n281));
  OAI21_X1  g080(.A(new_n279), .B1(new_n280), .B2(new_n281), .ZN(new_n282));
  NAND4_X1  g081(.A1(new_n229), .A2(new_n233), .A3(new_n247), .A4(new_n263), .ZN(new_n283));
  NAND3_X1  g082(.A1(new_n282), .A2(new_n276), .A3(new_n283), .ZN(new_n284));
  OAI21_X1  g083(.A(new_n278), .B1(new_n284), .B2(KEYINPUT34), .ZN(new_n285));
  NAND2_X1  g084(.A1(new_n284), .A2(KEYINPUT34), .ZN(new_n286));
  NAND3_X1  g085(.A1(new_n277), .A2(new_n285), .A3(new_n286), .ZN(new_n287));
  INV_X1    g086(.A(new_n270), .ZN(new_n288));
  AOI21_X1  g087(.A(new_n276), .B1(new_n282), .B2(new_n283), .ZN(new_n289));
  INV_X1    g088(.A(KEYINPUT32), .ZN(new_n290));
  OAI21_X1  g089(.A(new_n288), .B1(new_n289), .B2(new_n290), .ZN(new_n291));
  NOR2_X1   g090(.A1(new_n289), .A2(KEYINPUT33), .ZN(new_n292));
  OAI21_X1  g091(.A(KEYINPUT70), .B1(new_n291), .B2(new_n292), .ZN(new_n293));
  NAND2_X1  g092(.A1(new_n266), .A2(new_n271), .ZN(new_n294));
  INV_X1    g093(.A(KEYINPUT70), .ZN(new_n295));
  NAND4_X1  g094(.A1(new_n267), .A2(new_n294), .A3(new_n295), .A4(new_n288), .ZN(new_n296));
  AOI211_X1 g095(.A(new_n273), .B(new_n287), .C1(new_n293), .C2(new_n296), .ZN(new_n297));
  INV_X1    g096(.A(new_n287), .ZN(new_n298));
  NAND2_X1  g097(.A1(new_n293), .A2(new_n296), .ZN(new_n299));
  INV_X1    g098(.A(new_n273), .ZN(new_n300));
  AOI21_X1  g099(.A(new_n298), .B1(new_n299), .B2(new_n300), .ZN(new_n301));
  OAI211_X1 g100(.A(new_n202), .B(KEYINPUT36), .C1(new_n297), .C2(new_n301), .ZN(new_n302));
  NOR3_X1   g101(.A1(new_n291), .A2(new_n292), .A3(KEYINPUT70), .ZN(new_n303));
  AOI21_X1  g102(.A(new_n270), .B1(new_n266), .B2(KEYINPUT32), .ZN(new_n304));
  AOI21_X1  g103(.A(new_n295), .B1(new_n304), .B2(new_n294), .ZN(new_n305));
  OAI21_X1  g104(.A(new_n300), .B1(new_n303), .B2(new_n305), .ZN(new_n306));
  NAND2_X1  g105(.A1(new_n306), .A2(new_n287), .ZN(new_n307));
  NAND2_X1  g106(.A1(new_n202), .A2(KEYINPUT36), .ZN(new_n308));
  NAND3_X1  g107(.A1(new_n299), .A2(new_n298), .A3(new_n300), .ZN(new_n309));
  OR2_X1    g108(.A1(new_n202), .A2(KEYINPUT36), .ZN(new_n310));
  NAND4_X1  g109(.A1(new_n307), .A2(new_n308), .A3(new_n309), .A4(new_n310), .ZN(new_n311));
  NAND2_X1  g110(.A1(new_n302), .A2(new_n311), .ZN(new_n312));
  INV_X1    g111(.A(G22gat), .ZN(new_n313));
  OR2_X1    g112(.A1(G141gat), .A2(G148gat), .ZN(new_n314));
  NAND2_X1  g113(.A1(G141gat), .A2(G148gat), .ZN(new_n315));
  NAND2_X1  g114(.A1(new_n314), .A2(new_n315), .ZN(new_n316));
  INV_X1    g115(.A(KEYINPUT75), .ZN(new_n317));
  NAND2_X1  g116(.A1(new_n316), .A2(new_n317), .ZN(new_n318));
  INV_X1    g117(.A(KEYINPUT2), .ZN(new_n319));
  NAND3_X1  g118(.A1(new_n314), .A2(KEYINPUT75), .A3(new_n315), .ZN(new_n320));
  NAND3_X1  g119(.A1(new_n318), .A2(new_n319), .A3(new_n320), .ZN(new_n321));
  INV_X1    g120(.A(G155gat), .ZN(new_n322));
  INV_X1    g121(.A(G162gat), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n322), .A2(new_n323), .ZN(new_n324));
  NAND2_X1  g123(.A1(G155gat), .A2(G162gat), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n324), .A2(new_n325), .ZN(new_n326));
  INV_X1    g125(.A(new_n326), .ZN(new_n327));
  NAND2_X1  g126(.A1(new_n321), .A2(new_n327), .ZN(new_n328));
  INV_X1    g127(.A(KEYINPUT3), .ZN(new_n329));
  AOI21_X1  g128(.A(new_n316), .B1(KEYINPUT2), .B2(new_n325), .ZN(new_n330));
  NAND3_X1  g129(.A1(new_n324), .A2(KEYINPUT76), .A3(new_n325), .ZN(new_n331));
  INV_X1    g130(.A(KEYINPUT76), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n326), .A2(new_n332), .ZN(new_n333));
  NAND3_X1  g132(.A1(new_n330), .A2(new_n331), .A3(new_n333), .ZN(new_n334));
  NAND3_X1  g133(.A1(new_n328), .A2(new_n329), .A3(new_n334), .ZN(new_n335));
  INV_X1    g134(.A(KEYINPUT29), .ZN(new_n336));
  NAND2_X1  g135(.A1(new_n335), .A2(new_n336), .ZN(new_n337));
  XNOR2_X1  g136(.A(G197gat), .B(G204gat), .ZN(new_n338));
  INV_X1    g137(.A(KEYINPUT22), .ZN(new_n339));
  INV_X1    g138(.A(G211gat), .ZN(new_n340));
  INV_X1    g139(.A(G218gat), .ZN(new_n341));
  OAI21_X1  g140(.A(new_n339), .B1(new_n340), .B2(new_n341), .ZN(new_n342));
  NAND2_X1  g141(.A1(new_n338), .A2(new_n342), .ZN(new_n343));
  XOR2_X1   g142(.A(G211gat), .B(G218gat), .Z(new_n344));
  OR2_X1    g143(.A1(new_n343), .A2(new_n344), .ZN(new_n345));
  NAND2_X1  g144(.A1(new_n343), .A2(new_n344), .ZN(new_n346));
  AND2_X1   g145(.A1(new_n345), .A2(new_n346), .ZN(new_n347));
  NAND2_X1  g146(.A1(new_n337), .A2(new_n347), .ZN(new_n348));
  NAND2_X1  g147(.A1(new_n347), .A2(KEYINPUT82), .ZN(new_n349));
  INV_X1    g148(.A(new_n346), .ZN(new_n350));
  INV_X1    g149(.A(KEYINPUT82), .ZN(new_n351));
  AOI21_X1  g150(.A(KEYINPUT29), .B1(new_n350), .B2(new_n351), .ZN(new_n352));
  AOI21_X1  g151(.A(KEYINPUT3), .B1(new_n349), .B2(new_n352), .ZN(new_n353));
  AND2_X1   g152(.A1(new_n328), .A2(new_n334), .ZN(new_n354));
  OAI21_X1  g153(.A(new_n348), .B1(new_n353), .B2(new_n354), .ZN(new_n355));
  AND2_X1   g154(.A1(G228gat), .A2(G233gat), .ZN(new_n356));
  INV_X1    g155(.A(new_n356), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n355), .A2(new_n357), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n345), .A2(new_n346), .ZN(new_n359));
  AOI21_X1  g158(.A(KEYINPUT3), .B1(new_n359), .B2(new_n336), .ZN(new_n360));
  OAI211_X1 g159(.A(new_n348), .B(new_n356), .C1(new_n354), .C2(new_n360), .ZN(new_n361));
  AOI21_X1  g160(.A(new_n313), .B1(new_n358), .B2(new_n361), .ZN(new_n362));
  OR2_X1    g161(.A1(new_n362), .A2(KEYINPUT84), .ZN(new_n363));
  AND3_X1   g162(.A1(new_n358), .A2(new_n313), .A3(new_n361), .ZN(new_n364));
  XNOR2_X1  g163(.A(G78gat), .B(G106gat), .ZN(new_n365));
  INV_X1    g164(.A(G50gat), .ZN(new_n366));
  XNOR2_X1  g165(.A(new_n365), .B(new_n366), .ZN(new_n367));
  XNOR2_X1  g166(.A(KEYINPUT81), .B(KEYINPUT31), .ZN(new_n368));
  XNOR2_X1  g167(.A(new_n367), .B(new_n368), .ZN(new_n369));
  NOR2_X1   g168(.A1(new_n364), .A2(new_n369), .ZN(new_n370));
  NAND2_X1  g169(.A1(new_n362), .A2(KEYINPUT84), .ZN(new_n371));
  NAND3_X1  g170(.A1(new_n363), .A2(new_n370), .A3(new_n371), .ZN(new_n372));
  OAI21_X1  g171(.A(new_n369), .B1(new_n364), .B2(new_n362), .ZN(new_n373));
  INV_X1    g172(.A(KEYINPUT83), .ZN(new_n374));
  NAND2_X1  g173(.A1(new_n373), .A2(new_n374), .ZN(new_n375));
  OAI211_X1 g174(.A(KEYINPUT83), .B(new_n369), .C1(new_n364), .C2(new_n362), .ZN(new_n376));
  NAND3_X1  g175(.A1(new_n372), .A2(new_n375), .A3(new_n376), .ZN(new_n377));
  INV_X1    g176(.A(KEYINPUT80), .ZN(new_n378));
  INV_X1    g177(.A(KEYINPUT5), .ZN(new_n379));
  NAND3_X1  g178(.A1(new_n354), .A2(new_n232), .A3(new_n230), .ZN(new_n380));
  NAND2_X1  g179(.A1(new_n328), .A2(new_n334), .ZN(new_n381));
  OAI21_X1  g180(.A(new_n381), .B1(new_n220), .B2(new_n228), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n380), .A2(new_n382), .ZN(new_n383));
  NAND2_X1  g182(.A1(G225gat), .A2(G233gat), .ZN(new_n384));
  INV_X1    g183(.A(new_n384), .ZN(new_n385));
  AOI21_X1  g184(.A(new_n379), .B1(new_n383), .B2(new_n385), .ZN(new_n386));
  NAND3_X1  g185(.A1(new_n229), .A2(new_n233), .A3(new_n354), .ZN(new_n387));
  XNOR2_X1  g186(.A(KEYINPUT77), .B(KEYINPUT4), .ZN(new_n388));
  INV_X1    g187(.A(new_n388), .ZN(new_n389));
  NAND2_X1  g188(.A1(new_n230), .A2(new_n232), .ZN(new_n390));
  NOR2_X1   g189(.A1(new_n390), .A2(new_n381), .ZN(new_n391));
  INV_X1    g190(.A(KEYINPUT4), .ZN(new_n392));
  AOI22_X1  g191(.A1(new_n387), .A2(new_n389), .B1(new_n391), .B2(new_n392), .ZN(new_n393));
  NAND2_X1  g192(.A1(new_n381), .A2(KEYINPUT3), .ZN(new_n394));
  NAND3_X1  g193(.A1(new_n394), .A2(new_n390), .A3(new_n335), .ZN(new_n395));
  NAND2_X1  g194(.A1(new_n395), .A2(new_n384), .ZN(new_n396));
  OAI21_X1  g195(.A(new_n386), .B1(new_n393), .B2(new_n396), .ZN(new_n397));
  NAND2_X1  g196(.A1(new_n380), .A2(KEYINPUT4), .ZN(new_n398));
  NAND4_X1  g197(.A1(new_n229), .A2(new_n233), .A3(new_n354), .A4(new_n388), .ZN(new_n399));
  NAND2_X1  g198(.A1(new_n398), .A2(new_n399), .ZN(new_n400));
  NAND4_X1  g199(.A1(new_n400), .A2(new_n379), .A3(new_n384), .A4(new_n395), .ZN(new_n401));
  NAND2_X1  g200(.A1(new_n397), .A2(new_n401), .ZN(new_n402));
  XNOR2_X1  g201(.A(G1gat), .B(G29gat), .ZN(new_n403));
  XNOR2_X1  g202(.A(new_n403), .B(KEYINPUT0), .ZN(new_n404));
  XNOR2_X1  g203(.A(G57gat), .B(G85gat), .ZN(new_n405));
  XOR2_X1   g204(.A(new_n404), .B(new_n405), .Z(new_n406));
  INV_X1    g205(.A(new_n406), .ZN(new_n407));
  XOR2_X1   g206(.A(KEYINPUT78), .B(KEYINPUT6), .Z(new_n408));
  INV_X1    g207(.A(new_n408), .ZN(new_n409));
  AND4_X1   g208(.A1(new_n378), .A2(new_n402), .A3(new_n407), .A4(new_n409), .ZN(new_n410));
  AOI21_X1  g209(.A(new_n406), .B1(new_n397), .B2(new_n401), .ZN(new_n411));
  AOI21_X1  g210(.A(new_n378), .B1(new_n411), .B2(new_n409), .ZN(new_n412));
  NOR2_X1   g211(.A1(new_n410), .A2(new_n412), .ZN(new_n413));
  AOI21_X1  g212(.A(new_n409), .B1(new_n402), .B2(new_n407), .ZN(new_n414));
  INV_X1    g213(.A(KEYINPUT79), .ZN(new_n415));
  NAND3_X1  g214(.A1(new_n397), .A2(new_n401), .A3(new_n406), .ZN(new_n416));
  AND3_X1   g215(.A1(new_n414), .A2(new_n415), .A3(new_n416), .ZN(new_n417));
  AOI21_X1  g216(.A(new_n415), .B1(new_n414), .B2(new_n416), .ZN(new_n418));
  OAI21_X1  g217(.A(new_n413), .B1(new_n417), .B2(new_n418), .ZN(new_n419));
  AND2_X1   g218(.A1(G226gat), .A2(G233gat), .ZN(new_n420));
  NAND2_X1  g219(.A1(new_n279), .A2(new_n420), .ZN(new_n421));
  AOI21_X1  g220(.A(KEYINPUT29), .B1(new_n247), .B2(new_n263), .ZN(new_n422));
  OAI21_X1  g221(.A(new_n421), .B1(new_n422), .B2(new_n420), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n423), .A2(new_n347), .ZN(new_n424));
  OAI211_X1 g223(.A(new_n421), .B(new_n359), .C1(new_n422), .C2(new_n420), .ZN(new_n425));
  XNOR2_X1  g224(.A(G8gat), .B(G36gat), .ZN(new_n426));
  XNOR2_X1  g225(.A(G64gat), .B(G92gat), .ZN(new_n427));
  XOR2_X1   g226(.A(new_n426), .B(new_n427), .Z(new_n428));
  NAND3_X1  g227(.A1(new_n424), .A2(new_n425), .A3(new_n428), .ZN(new_n429));
  XNOR2_X1  g228(.A(KEYINPUT74), .B(KEYINPUT30), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n429), .A2(new_n430), .ZN(new_n431));
  INV_X1    g230(.A(new_n428), .ZN(new_n432));
  AND2_X1   g231(.A1(new_n423), .A2(new_n347), .ZN(new_n433));
  INV_X1    g232(.A(new_n425), .ZN(new_n434));
  OAI21_X1  g233(.A(new_n432), .B1(new_n433), .B2(new_n434), .ZN(new_n435));
  INV_X1    g234(.A(KEYINPUT73), .ZN(new_n436));
  NAND4_X1  g235(.A1(new_n424), .A2(KEYINPUT30), .A3(new_n425), .A4(new_n428), .ZN(new_n437));
  NAND4_X1  g236(.A1(new_n431), .A2(new_n435), .A3(new_n436), .A4(new_n437), .ZN(new_n438));
  OR2_X1    g237(.A1(new_n437), .A2(new_n436), .ZN(new_n439));
  NAND2_X1  g238(.A1(new_n438), .A2(new_n439), .ZN(new_n440));
  AOI21_X1  g239(.A(new_n377), .B1(new_n419), .B2(new_n440), .ZN(new_n441));
  NOR2_X1   g240(.A1(new_n312), .A2(new_n441), .ZN(new_n442));
  INV_X1    g241(.A(new_n395), .ZN(new_n443));
  AOI21_X1  g242(.A(new_n443), .B1(new_n399), .B2(new_n398), .ZN(new_n444));
  OAI21_X1  g243(.A(KEYINPUT85), .B1(new_n444), .B2(new_n384), .ZN(new_n445));
  NAND2_X1  g244(.A1(new_n400), .A2(new_n395), .ZN(new_n446));
  INV_X1    g245(.A(KEYINPUT85), .ZN(new_n447));
  NAND3_X1  g246(.A1(new_n446), .A2(new_n447), .A3(new_n385), .ZN(new_n448));
  NAND2_X1  g247(.A1(new_n445), .A2(new_n448), .ZN(new_n449));
  INV_X1    g248(.A(KEYINPUT39), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n449), .A2(new_n450), .ZN(new_n451));
  NAND3_X1  g250(.A1(new_n380), .A2(new_n384), .A3(new_n382), .ZN(new_n452));
  NAND4_X1  g251(.A1(new_n445), .A2(new_n448), .A3(KEYINPUT39), .A4(new_n452), .ZN(new_n453));
  NAND3_X1  g252(.A1(new_n451), .A2(new_n453), .A3(new_n406), .ZN(new_n454));
  INV_X1    g253(.A(KEYINPUT86), .ZN(new_n455));
  NOR2_X1   g254(.A1(new_n455), .A2(KEYINPUT40), .ZN(new_n456));
  NAND2_X1  g255(.A1(new_n454), .A2(new_n456), .ZN(new_n457));
  INV_X1    g256(.A(new_n411), .ZN(new_n458));
  AND3_X1   g257(.A1(new_n438), .A2(new_n439), .A3(new_n458), .ZN(new_n459));
  INV_X1    g258(.A(new_n456), .ZN(new_n460));
  NAND4_X1  g259(.A1(new_n451), .A2(new_n460), .A3(new_n453), .A4(new_n406), .ZN(new_n461));
  AND3_X1   g260(.A1(new_n457), .A2(new_n459), .A3(new_n461), .ZN(new_n462));
  INV_X1    g261(.A(new_n412), .ZN(new_n463));
  NAND2_X1  g262(.A1(new_n414), .A2(new_n416), .ZN(new_n464));
  NAND3_X1  g263(.A1(new_n411), .A2(new_n378), .A3(new_n409), .ZN(new_n465));
  NAND3_X1  g264(.A1(new_n463), .A2(new_n464), .A3(new_n465), .ZN(new_n466));
  OAI21_X1  g265(.A(KEYINPUT37), .B1(new_n433), .B2(new_n434), .ZN(new_n467));
  INV_X1    g266(.A(KEYINPUT37), .ZN(new_n468));
  NAND3_X1  g267(.A1(new_n424), .A2(new_n468), .A3(new_n425), .ZN(new_n469));
  NAND3_X1  g268(.A1(new_n467), .A2(new_n432), .A3(new_n469), .ZN(new_n470));
  NAND2_X1  g269(.A1(new_n470), .A2(KEYINPUT38), .ZN(new_n471));
  INV_X1    g270(.A(KEYINPUT38), .ZN(new_n472));
  NAND4_X1  g271(.A1(new_n467), .A2(new_n472), .A3(new_n432), .A4(new_n469), .ZN(new_n473));
  NAND3_X1  g272(.A1(new_n471), .A2(new_n429), .A3(new_n473), .ZN(new_n474));
  OAI21_X1  g273(.A(new_n377), .B1(new_n466), .B2(new_n474), .ZN(new_n475));
  OR2_X1    g274(.A1(new_n462), .A2(new_n475), .ZN(new_n476));
  NAND2_X1  g275(.A1(new_n419), .A2(new_n440), .ZN(new_n477));
  NAND3_X1  g276(.A1(new_n377), .A2(new_n307), .A3(new_n309), .ZN(new_n478));
  OAI21_X1  g277(.A(KEYINPUT35), .B1(new_n477), .B2(new_n478), .ZN(new_n479));
  INV_X1    g278(.A(new_n478), .ZN(new_n480));
  INV_X1    g279(.A(KEYINPUT35), .ZN(new_n481));
  AND3_X1   g280(.A1(new_n466), .A2(new_n481), .A3(new_n440), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n480), .A2(new_n482), .ZN(new_n483));
  AOI22_X1  g282(.A1(new_n442), .A2(new_n476), .B1(new_n479), .B2(new_n483), .ZN(new_n484));
  XNOR2_X1  g283(.A(G113gat), .B(G141gat), .ZN(new_n485));
  XNOR2_X1  g284(.A(KEYINPUT87), .B(KEYINPUT11), .ZN(new_n486));
  XNOR2_X1  g285(.A(new_n485), .B(new_n486), .ZN(new_n487));
  XNOR2_X1  g286(.A(G169gat), .B(G197gat), .ZN(new_n488));
  XNOR2_X1  g287(.A(new_n487), .B(new_n488), .ZN(new_n489));
  XNOR2_X1  g288(.A(new_n489), .B(KEYINPUT12), .ZN(new_n490));
  INV_X1    g289(.A(new_n490), .ZN(new_n491));
  XNOR2_X1  g290(.A(G15gat), .B(G22gat), .ZN(new_n492));
  INV_X1    g291(.A(KEYINPUT16), .ZN(new_n493));
  OAI21_X1  g292(.A(new_n492), .B1(new_n493), .B2(G1gat), .ZN(new_n494));
  OAI21_X1  g293(.A(new_n494), .B1(G1gat), .B2(new_n492), .ZN(new_n495));
  XOR2_X1   g294(.A(new_n495), .B(G8gat), .Z(new_n496));
  INV_X1    g295(.A(G29gat), .ZN(new_n497));
  AND3_X1   g296(.A1(new_n497), .A2(KEYINPUT14), .A3(G36gat), .ZN(new_n498));
  XNOR2_X1  g297(.A(KEYINPUT14), .B(G29gat), .ZN(new_n499));
  INV_X1    g298(.A(G36gat), .ZN(new_n500));
  AOI21_X1  g299(.A(new_n498), .B1(new_n499), .B2(new_n500), .ZN(new_n501));
  AND2_X1   g300(.A1(G43gat), .A2(G50gat), .ZN(new_n502));
  NOR2_X1   g301(.A1(G43gat), .A2(G50gat), .ZN(new_n503));
  OAI21_X1  g302(.A(KEYINPUT15), .B1(new_n502), .B2(new_n503), .ZN(new_n504));
  INV_X1    g303(.A(G43gat), .ZN(new_n505));
  NAND2_X1  g304(.A1(new_n505), .A2(new_n366), .ZN(new_n506));
  INV_X1    g305(.A(KEYINPUT15), .ZN(new_n507));
  NAND2_X1  g306(.A1(G43gat), .A2(G50gat), .ZN(new_n508));
  NAND3_X1  g307(.A1(new_n506), .A2(new_n507), .A3(new_n508), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n504), .A2(new_n509), .ZN(new_n510));
  OAI21_X1  g309(.A(KEYINPUT88), .B1(new_n501), .B2(new_n510), .ZN(new_n511));
  INV_X1    g310(.A(new_n504), .ZN(new_n512));
  NAND2_X1  g311(.A1(new_n501), .A2(new_n512), .ZN(new_n513));
  AND2_X1   g312(.A1(KEYINPUT14), .A2(G29gat), .ZN(new_n514));
  NOR2_X1   g313(.A1(KEYINPUT14), .A2(G29gat), .ZN(new_n515));
  OAI21_X1  g314(.A(new_n500), .B1(new_n514), .B2(new_n515), .ZN(new_n516));
  NAND3_X1  g315(.A1(new_n497), .A2(KEYINPUT14), .A3(G36gat), .ZN(new_n517));
  NAND2_X1  g316(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  INV_X1    g317(.A(KEYINPUT88), .ZN(new_n519));
  NAND4_X1  g318(.A1(new_n518), .A2(new_n519), .A3(new_n504), .A4(new_n509), .ZN(new_n520));
  NAND3_X1  g319(.A1(new_n511), .A2(new_n513), .A3(new_n520), .ZN(new_n521));
  XNOR2_X1  g320(.A(new_n496), .B(new_n521), .ZN(new_n522));
  NAND2_X1  g321(.A1(G229gat), .A2(G233gat), .ZN(new_n523));
  XOR2_X1   g322(.A(new_n523), .B(KEYINPUT13), .Z(new_n524));
  INV_X1    g323(.A(new_n524), .ZN(new_n525));
  NOR2_X1   g324(.A1(new_n522), .A2(new_n525), .ZN(new_n526));
  INV_X1    g325(.A(new_n526), .ZN(new_n527));
  INV_X1    g326(.A(KEYINPUT89), .ZN(new_n528));
  AND3_X1   g327(.A1(new_n521), .A2(new_n528), .A3(KEYINPUT17), .ZN(new_n529));
  AOI21_X1  g328(.A(KEYINPUT17), .B1(new_n521), .B2(new_n528), .ZN(new_n530));
  OAI21_X1  g329(.A(new_n496), .B1(new_n529), .B2(new_n530), .ZN(new_n531));
  INV_X1    g330(.A(KEYINPUT90), .ZN(new_n532));
  XNOR2_X1  g331(.A(new_n495), .B(G8gat), .ZN(new_n533));
  AOI21_X1  g332(.A(new_n532), .B1(new_n533), .B2(new_n521), .ZN(new_n534));
  NAND2_X1  g333(.A1(new_n531), .A2(new_n534), .ZN(new_n535));
  OAI211_X1 g334(.A(new_n532), .B(new_n496), .C1(new_n529), .C2(new_n530), .ZN(new_n536));
  AOI22_X1  g335(.A1(new_n535), .A2(new_n536), .B1(G229gat), .B2(G233gat), .ZN(new_n537));
  OAI21_X1  g336(.A(new_n527), .B1(new_n537), .B2(KEYINPUT18), .ZN(new_n538));
  NAND2_X1  g337(.A1(new_n520), .A2(new_n513), .ZN(new_n539));
  AND2_X1   g338(.A1(new_n504), .A2(new_n509), .ZN(new_n540));
  AOI21_X1  g339(.A(new_n519), .B1(new_n540), .B2(new_n518), .ZN(new_n541));
  OAI21_X1  g340(.A(new_n528), .B1(new_n539), .B2(new_n541), .ZN(new_n542));
  INV_X1    g341(.A(KEYINPUT17), .ZN(new_n543));
  NAND2_X1  g342(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  NAND3_X1  g343(.A1(new_n521), .A2(new_n528), .A3(KEYINPUT17), .ZN(new_n545));
  AOI21_X1  g344(.A(new_n533), .B1(new_n544), .B2(new_n545), .ZN(new_n546));
  INV_X1    g345(.A(new_n534), .ZN(new_n547));
  OAI21_X1  g346(.A(new_n536), .B1(new_n546), .B2(new_n547), .ZN(new_n548));
  NAND2_X1  g347(.A1(new_n548), .A2(new_n523), .ZN(new_n549));
  INV_X1    g348(.A(KEYINPUT18), .ZN(new_n550));
  NOR2_X1   g349(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  OAI21_X1  g350(.A(new_n491), .B1(new_n538), .B2(new_n551), .ZN(new_n552));
  AOI21_X1  g351(.A(new_n526), .B1(new_n549), .B2(new_n550), .ZN(new_n553));
  NAND2_X1  g352(.A1(new_n537), .A2(KEYINPUT18), .ZN(new_n554));
  NAND3_X1  g353(.A1(new_n553), .A2(new_n554), .A3(new_n490), .ZN(new_n555));
  NAND2_X1  g354(.A1(new_n552), .A2(new_n555), .ZN(new_n556));
  INV_X1    g355(.A(new_n556), .ZN(new_n557));
  NOR2_X1   g356(.A1(new_n484), .A2(new_n557), .ZN(new_n558));
  OR2_X1    g357(.A1(G57gat), .A2(G64gat), .ZN(new_n559));
  NAND2_X1  g358(.A1(G57gat), .A2(G64gat), .ZN(new_n560));
  AND2_X1   g359(.A1(new_n559), .A2(new_n560), .ZN(new_n561));
  INV_X1    g360(.A(KEYINPUT9), .ZN(new_n562));
  INV_X1    g361(.A(G71gat), .ZN(new_n563));
  INV_X1    g362(.A(G78gat), .ZN(new_n564));
  OAI21_X1  g363(.A(new_n562), .B1(new_n563), .B2(new_n564), .ZN(new_n565));
  XNOR2_X1  g364(.A(G71gat), .B(G78gat), .ZN(new_n566));
  INV_X1    g365(.A(new_n566), .ZN(new_n567));
  OAI211_X1 g366(.A(new_n561), .B(new_n565), .C1(new_n567), .C2(KEYINPUT91), .ZN(new_n568));
  NAND3_X1  g367(.A1(new_n565), .A2(new_n559), .A3(new_n560), .ZN(new_n569));
  NAND3_X1  g368(.A1(new_n559), .A2(KEYINPUT91), .A3(new_n560), .ZN(new_n570));
  NAND3_X1  g369(.A1(new_n569), .A2(new_n566), .A3(new_n570), .ZN(new_n571));
  NAND2_X1  g370(.A1(new_n568), .A2(new_n571), .ZN(new_n572));
  NOR2_X1   g371(.A1(new_n572), .A2(KEYINPUT21), .ZN(new_n573));
  NAND2_X1  g372(.A1(G231gat), .A2(G233gat), .ZN(new_n574));
  XNOR2_X1  g373(.A(new_n573), .B(new_n574), .ZN(new_n575));
  XNOR2_X1  g374(.A(new_n575), .B(new_n214), .ZN(new_n576));
  AOI21_X1  g375(.A(new_n533), .B1(KEYINPUT21), .B2(new_n572), .ZN(new_n577));
  XNOR2_X1  g376(.A(new_n577), .B(KEYINPUT92), .ZN(new_n578));
  OR2_X1    g377(.A1(new_n576), .A2(new_n578), .ZN(new_n579));
  NAND2_X1  g378(.A1(new_n576), .A2(new_n578), .ZN(new_n580));
  XNOR2_X1  g379(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n581));
  XNOR2_X1  g380(.A(new_n581), .B(G155gat), .ZN(new_n582));
  XNOR2_X1  g381(.A(G183gat), .B(G211gat), .ZN(new_n583));
  XNOR2_X1  g382(.A(new_n582), .B(new_n583), .ZN(new_n584));
  AND3_X1   g383(.A1(new_n579), .A2(new_n580), .A3(new_n584), .ZN(new_n585));
  AOI21_X1  g384(.A(new_n584), .B1(new_n579), .B2(new_n580), .ZN(new_n586));
  OR2_X1    g385(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  INV_X1    g386(.A(new_n587), .ZN(new_n588));
  INV_X1    g387(.A(KEYINPUT97), .ZN(new_n589));
  NAND2_X1  g388(.A1(G232gat), .A2(G233gat), .ZN(new_n590));
  INV_X1    g389(.A(KEYINPUT41), .ZN(new_n591));
  NAND2_X1  g390(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  XNOR2_X1  g391(.A(new_n592), .B(KEYINPUT93), .ZN(new_n593));
  XNOR2_X1  g392(.A(G134gat), .B(G162gat), .ZN(new_n594));
  XNOR2_X1  g393(.A(new_n593), .B(new_n594), .ZN(new_n595));
  INV_X1    g394(.A(KEYINPUT94), .ZN(new_n596));
  OAI211_X1 g395(.A(new_n596), .B(KEYINPUT7), .C1(G85gat), .C2(G92gat), .ZN(new_n597));
  INV_X1    g396(.A(G85gat), .ZN(new_n598));
  INV_X1    g397(.A(G92gat), .ZN(new_n599));
  OAI21_X1  g398(.A(new_n597), .B1(new_n598), .B2(new_n599), .ZN(new_n600));
  INV_X1    g399(.A(G99gat), .ZN(new_n601));
  INV_X1    g400(.A(G106gat), .ZN(new_n602));
  OAI21_X1  g401(.A(KEYINPUT95), .B1(new_n601), .B2(new_n602), .ZN(new_n603));
  INV_X1    g402(.A(KEYINPUT95), .ZN(new_n604));
  NAND3_X1  g403(.A1(new_n604), .A2(G99gat), .A3(G106gat), .ZN(new_n605));
  NAND3_X1  g404(.A1(new_n603), .A2(KEYINPUT8), .A3(new_n605), .ZN(new_n606));
  NAND4_X1  g405(.A1(new_n596), .A2(KEYINPUT7), .A3(G85gat), .A4(G92gat), .ZN(new_n607));
  NAND3_X1  g406(.A1(new_n600), .A2(new_n606), .A3(new_n607), .ZN(new_n608));
  XOR2_X1   g407(.A(G99gat), .B(G106gat), .Z(new_n609));
  NAND2_X1  g408(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  INV_X1    g409(.A(new_n609), .ZN(new_n611));
  NAND4_X1  g410(.A1(new_n611), .A2(new_n606), .A3(new_n600), .A4(new_n607), .ZN(new_n612));
  NAND2_X1  g411(.A1(new_n610), .A2(new_n612), .ZN(new_n613));
  OAI21_X1  g412(.A(new_n613), .B1(new_n529), .B2(new_n530), .ZN(new_n614));
  NOR2_X1   g413(.A1(new_n590), .A2(new_n591), .ZN(new_n615));
  INV_X1    g414(.A(new_n613), .ZN(new_n616));
  AOI21_X1  g415(.A(new_n615), .B1(new_n616), .B2(new_n521), .ZN(new_n617));
  XNOR2_X1  g416(.A(G190gat), .B(G218gat), .ZN(new_n618));
  XOR2_X1   g417(.A(new_n618), .B(KEYINPUT96), .Z(new_n619));
  NAND3_X1  g418(.A1(new_n614), .A2(new_n617), .A3(new_n619), .ZN(new_n620));
  INV_X1    g419(.A(new_n620), .ZN(new_n621));
  NOR2_X1   g420(.A1(new_n618), .A2(KEYINPUT96), .ZN(new_n622));
  INV_X1    g421(.A(new_n622), .ZN(new_n623));
  AOI21_X1  g422(.A(new_n623), .B1(new_n614), .B2(new_n617), .ZN(new_n624));
  OAI211_X1 g423(.A(new_n589), .B(new_n595), .C1(new_n621), .C2(new_n624), .ZN(new_n625));
  INV_X1    g424(.A(new_n624), .ZN(new_n626));
  NAND2_X1  g425(.A1(new_n595), .A2(new_n589), .ZN(new_n627));
  OR2_X1    g426(.A1(new_n595), .A2(new_n589), .ZN(new_n628));
  NAND4_X1  g427(.A1(new_n626), .A2(new_n627), .A3(new_n620), .A4(new_n628), .ZN(new_n629));
  NAND2_X1  g428(.A1(new_n625), .A2(new_n629), .ZN(new_n630));
  NAND3_X1  g429(.A1(new_n613), .A2(new_n568), .A3(new_n571), .ZN(new_n631));
  INV_X1    g430(.A(KEYINPUT10), .ZN(new_n632));
  NAND3_X1  g431(.A1(new_n572), .A2(new_n610), .A3(new_n612), .ZN(new_n633));
  NAND3_X1  g432(.A1(new_n631), .A2(new_n632), .A3(new_n633), .ZN(new_n634));
  NAND4_X1  g433(.A1(new_n572), .A2(new_n610), .A3(KEYINPUT10), .A4(new_n612), .ZN(new_n635));
  INV_X1    g434(.A(KEYINPUT98), .ZN(new_n636));
  AND2_X1   g435(.A1(new_n635), .A2(new_n636), .ZN(new_n637));
  NAND2_X1  g436(.A1(new_n634), .A2(new_n637), .ZN(new_n638));
  NAND2_X1  g437(.A1(G230gat), .A2(G233gat), .ZN(new_n639));
  NOR2_X1   g438(.A1(new_n635), .A2(new_n636), .ZN(new_n640));
  INV_X1    g439(.A(new_n640), .ZN(new_n641));
  NAND3_X1  g440(.A1(new_n638), .A2(new_n639), .A3(new_n641), .ZN(new_n642));
  NAND2_X1  g441(.A1(new_n631), .A2(new_n633), .ZN(new_n643));
  INV_X1    g442(.A(new_n639), .ZN(new_n644));
  NAND2_X1  g443(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  AND2_X1   g444(.A1(new_n642), .A2(new_n645), .ZN(new_n646));
  XNOR2_X1  g445(.A(G120gat), .B(G148gat), .ZN(new_n647));
  XNOR2_X1  g446(.A(G176gat), .B(G204gat), .ZN(new_n648));
  XOR2_X1   g447(.A(new_n647), .B(new_n648), .Z(new_n649));
  OR2_X1    g448(.A1(new_n646), .A2(new_n649), .ZN(new_n650));
  NAND3_X1  g449(.A1(new_n642), .A2(new_n645), .A3(new_n649), .ZN(new_n651));
  AND2_X1   g450(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  NAND3_X1  g451(.A1(new_n588), .A2(new_n630), .A3(new_n652), .ZN(new_n653));
  INV_X1    g452(.A(new_n653), .ZN(new_n654));
  OR2_X1    g453(.A1(new_n419), .A2(KEYINPUT99), .ZN(new_n655));
  NAND2_X1  g454(.A1(new_n419), .A2(KEYINPUT99), .ZN(new_n656));
  NAND2_X1  g455(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  INV_X1    g456(.A(new_n657), .ZN(new_n658));
  NAND3_X1  g457(.A1(new_n558), .A2(new_n654), .A3(new_n658), .ZN(new_n659));
  XNOR2_X1  g458(.A(new_n659), .B(G1gat), .ZN(G1324gat));
  NAND2_X1  g459(.A1(new_n558), .A2(new_n654), .ZN(new_n661));
  OAI21_X1  g460(.A(G8gat), .B1(new_n661), .B2(new_n440), .ZN(new_n662));
  INV_X1    g461(.A(new_n440), .ZN(new_n663));
  XOR2_X1   g462(.A(KEYINPUT16), .B(G8gat), .Z(new_n664));
  NAND4_X1  g463(.A1(new_n558), .A2(new_n663), .A3(new_n654), .A4(new_n664), .ZN(new_n665));
  NAND2_X1  g464(.A1(new_n662), .A2(new_n665), .ZN(new_n666));
  NAND2_X1  g465(.A1(new_n666), .A2(KEYINPUT42), .ZN(new_n667));
  INV_X1    g466(.A(KEYINPUT42), .ZN(new_n668));
  NAND2_X1  g467(.A1(new_n665), .A2(new_n668), .ZN(new_n669));
  NAND2_X1  g468(.A1(new_n667), .A2(new_n669), .ZN(new_n670));
  INV_X1    g469(.A(KEYINPUT100), .ZN(new_n671));
  XNOR2_X1  g470(.A(new_n670), .B(new_n671), .ZN(G1325gat));
  INV_X1    g471(.A(new_n312), .ZN(new_n673));
  OAI21_X1  g472(.A(G15gat), .B1(new_n661), .B2(new_n673), .ZN(new_n674));
  NOR2_X1   g473(.A1(new_n297), .A2(new_n301), .ZN(new_n675));
  NOR2_X1   g474(.A1(new_n653), .A2(G15gat), .ZN(new_n676));
  NAND3_X1  g475(.A1(new_n558), .A2(new_n675), .A3(new_n676), .ZN(new_n677));
  NAND2_X1  g476(.A1(new_n674), .A2(new_n677), .ZN(G1326gat));
  NOR2_X1   g477(.A1(new_n661), .A2(new_n377), .ZN(new_n679));
  XOR2_X1   g478(.A(KEYINPUT43), .B(G22gat), .Z(new_n680));
  XNOR2_X1  g479(.A(new_n679), .B(new_n680), .ZN(G1327gat));
  NAND2_X1  g480(.A1(new_n587), .A2(new_n652), .ZN(new_n682));
  NOR4_X1   g481(.A1(new_n484), .A2(new_n557), .A3(new_n630), .A4(new_n682), .ZN(new_n683));
  NAND3_X1  g482(.A1(new_n683), .A2(new_n497), .A3(new_n658), .ZN(new_n684));
  XNOR2_X1  g483(.A(new_n684), .B(KEYINPUT45), .ZN(new_n685));
  INV_X1    g484(.A(KEYINPUT44), .ZN(new_n686));
  OAI21_X1  g485(.A(new_n686), .B1(new_n484), .B2(new_n630), .ZN(new_n687));
  AND2_X1   g486(.A1(new_n625), .A2(new_n629), .ZN(new_n688));
  NOR2_X1   g487(.A1(new_n462), .A2(new_n475), .ZN(new_n689));
  NOR3_X1   g488(.A1(new_n689), .A2(new_n312), .A3(new_n441), .ZN(new_n690));
  NAND4_X1  g489(.A1(new_n675), .A2(new_n419), .A3(new_n440), .A4(new_n377), .ZN(new_n691));
  AOI22_X1  g490(.A1(new_n691), .A2(KEYINPUT35), .B1(new_n480), .B2(new_n482), .ZN(new_n692));
  OAI211_X1 g491(.A(KEYINPUT44), .B(new_n688), .C1(new_n690), .C2(new_n692), .ZN(new_n693));
  AND2_X1   g492(.A1(new_n687), .A2(new_n693), .ZN(new_n694));
  INV_X1    g493(.A(KEYINPUT101), .ZN(new_n695));
  NAND2_X1  g494(.A1(new_n549), .A2(new_n550), .ZN(new_n696));
  AND4_X1   g495(.A1(new_n554), .A2(new_n696), .A3(new_n527), .A4(new_n490), .ZN(new_n697));
  AOI21_X1  g496(.A(new_n490), .B1(new_n553), .B2(new_n554), .ZN(new_n698));
  OAI21_X1  g497(.A(new_n695), .B1(new_n697), .B2(new_n698), .ZN(new_n699));
  NAND3_X1  g498(.A1(new_n552), .A2(new_n555), .A3(KEYINPUT101), .ZN(new_n700));
  NAND2_X1  g499(.A1(new_n699), .A2(new_n700), .ZN(new_n701));
  INV_X1    g500(.A(new_n701), .ZN(new_n702));
  NOR2_X1   g501(.A1(new_n702), .A2(new_n682), .ZN(new_n703));
  NAND2_X1  g502(.A1(new_n694), .A2(new_n703), .ZN(new_n704));
  OAI21_X1  g503(.A(KEYINPUT102), .B1(new_n704), .B2(new_n657), .ZN(new_n705));
  NAND2_X1  g504(.A1(new_n705), .A2(G29gat), .ZN(new_n706));
  NOR3_X1   g505(.A1(new_n704), .A2(KEYINPUT102), .A3(new_n657), .ZN(new_n707));
  OAI21_X1  g506(.A(new_n685), .B1(new_n706), .B2(new_n707), .ZN(G1328gat));
  NAND3_X1  g507(.A1(new_n683), .A2(new_n500), .A3(new_n663), .ZN(new_n709));
  XOR2_X1   g508(.A(new_n709), .B(KEYINPUT46), .Z(new_n710));
  OAI21_X1  g509(.A(G36gat), .B1(new_n704), .B2(new_n440), .ZN(new_n711));
  NAND2_X1  g510(.A1(new_n710), .A2(new_n711), .ZN(G1329gat));
  OAI21_X1  g511(.A(G43gat), .B1(new_n704), .B2(new_n673), .ZN(new_n713));
  AOI21_X1  g512(.A(KEYINPUT47), .B1(new_n713), .B2(KEYINPUT103), .ZN(new_n714));
  NAND3_X1  g513(.A1(new_n683), .A2(new_n505), .A3(new_n675), .ZN(new_n715));
  NAND2_X1  g514(.A1(new_n713), .A2(new_n715), .ZN(new_n716));
  NAND2_X1  g515(.A1(new_n714), .A2(new_n716), .ZN(new_n717));
  OAI211_X1 g516(.A(new_n713), .B(new_n715), .C1(KEYINPUT103), .C2(KEYINPUT47), .ZN(new_n718));
  NAND2_X1  g517(.A1(new_n717), .A2(new_n718), .ZN(G1330gat));
  OAI21_X1  g518(.A(G50gat), .B1(new_n704), .B2(new_n377), .ZN(new_n720));
  INV_X1    g519(.A(new_n377), .ZN(new_n721));
  NAND2_X1  g520(.A1(new_n721), .A2(new_n366), .ZN(new_n722));
  XNOR2_X1  g521(.A(new_n722), .B(KEYINPUT104), .ZN(new_n723));
  NAND2_X1  g522(.A1(new_n683), .A2(new_n723), .ZN(new_n724));
  NAND2_X1  g523(.A1(new_n720), .A2(new_n724), .ZN(new_n725));
  INV_X1    g524(.A(KEYINPUT48), .ZN(new_n726));
  XNOR2_X1  g525(.A(new_n725), .B(new_n726), .ZN(G1331gat));
  INV_X1    g526(.A(new_n652), .ZN(new_n728));
  NAND3_X1  g527(.A1(new_n588), .A2(new_n630), .A3(new_n728), .ZN(new_n729));
  NOR3_X1   g528(.A1(new_n484), .A2(new_n701), .A3(new_n729), .ZN(new_n730));
  NAND2_X1  g529(.A1(new_n730), .A2(new_n658), .ZN(new_n731));
  XNOR2_X1  g530(.A(new_n731), .B(G57gat), .ZN(G1332gat));
  XNOR2_X1  g531(.A(new_n440), .B(KEYINPUT105), .ZN(new_n733));
  AOI21_X1  g532(.A(new_n733), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n734));
  NAND2_X1  g533(.A1(new_n730), .A2(new_n734), .ZN(new_n735));
  XOR2_X1   g534(.A(new_n735), .B(KEYINPUT106), .Z(new_n736));
  NOR2_X1   g535(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n737));
  XNOR2_X1  g536(.A(new_n736), .B(new_n737), .ZN(G1333gat));
  NAND3_X1  g537(.A1(new_n730), .A2(new_n563), .A3(new_n675), .ZN(new_n739));
  AND2_X1   g538(.A1(new_n730), .A2(new_n312), .ZN(new_n740));
  OAI21_X1  g539(.A(new_n739), .B1(new_n740), .B2(new_n563), .ZN(new_n741));
  XOR2_X1   g540(.A(KEYINPUT107), .B(KEYINPUT50), .Z(new_n742));
  XNOR2_X1  g541(.A(new_n741), .B(new_n742), .ZN(G1334gat));
  NAND2_X1  g542(.A1(new_n730), .A2(new_n721), .ZN(new_n744));
  XNOR2_X1  g543(.A(KEYINPUT108), .B(G78gat), .ZN(new_n745));
  XNOR2_X1  g544(.A(new_n744), .B(new_n745), .ZN(G1335gat));
  NOR3_X1   g545(.A1(new_n701), .A2(new_n588), .A3(new_n652), .ZN(new_n747));
  NAND2_X1  g546(.A1(new_n694), .A2(new_n747), .ZN(new_n748));
  OAI21_X1  g547(.A(G85gat), .B1(new_n748), .B2(new_n657), .ZN(new_n749));
  NOR2_X1   g548(.A1(new_n701), .A2(new_n588), .ZN(new_n750));
  OAI211_X1 g549(.A(new_n688), .B(new_n750), .C1(new_n690), .C2(new_n692), .ZN(new_n751));
  INV_X1    g550(.A(KEYINPUT51), .ZN(new_n752));
  NAND2_X1  g551(.A1(new_n751), .A2(new_n752), .ZN(new_n753));
  NAND2_X1  g552(.A1(new_n442), .A2(new_n476), .ZN(new_n754));
  NAND2_X1  g553(.A1(new_n479), .A2(new_n483), .ZN(new_n755));
  NAND2_X1  g554(.A1(new_n754), .A2(new_n755), .ZN(new_n756));
  NAND4_X1  g555(.A1(new_n756), .A2(KEYINPUT51), .A3(new_n688), .A4(new_n750), .ZN(new_n757));
  NAND2_X1  g556(.A1(new_n753), .A2(new_n757), .ZN(new_n758));
  AOI21_X1  g557(.A(new_n652), .B1(new_n758), .B2(KEYINPUT109), .ZN(new_n759));
  OAI21_X1  g558(.A(new_n759), .B1(KEYINPUT109), .B2(new_n758), .ZN(new_n760));
  NAND2_X1  g559(.A1(new_n658), .A2(new_n598), .ZN(new_n761));
  OAI21_X1  g560(.A(new_n749), .B1(new_n760), .B2(new_n761), .ZN(G1336gat));
  INV_X1    g561(.A(new_n748), .ZN(new_n763));
  NAND2_X1  g562(.A1(new_n763), .A2(new_n663), .ZN(new_n764));
  NOR3_X1   g563(.A1(new_n733), .A2(G92gat), .A3(new_n652), .ZN(new_n765));
  AOI22_X1  g564(.A1(new_n764), .A2(G92gat), .B1(new_n758), .B2(new_n765), .ZN(new_n766));
  INV_X1    g565(.A(KEYINPUT52), .ZN(new_n767));
  INV_X1    g566(.A(new_n733), .ZN(new_n768));
  AOI21_X1  g567(.A(new_n599), .B1(new_n763), .B2(new_n768), .ZN(new_n769));
  NAND2_X1  g568(.A1(new_n758), .A2(new_n765), .ZN(new_n770));
  XNOR2_X1  g569(.A(KEYINPUT110), .B(KEYINPUT52), .ZN(new_n771));
  NAND2_X1  g570(.A1(new_n770), .A2(new_n771), .ZN(new_n772));
  OAI22_X1  g571(.A1(new_n766), .A2(new_n767), .B1(new_n769), .B2(new_n772), .ZN(G1337gat));
  OAI21_X1  g572(.A(G99gat), .B1(new_n748), .B2(new_n673), .ZN(new_n774));
  NAND2_X1  g573(.A1(new_n675), .A2(new_n601), .ZN(new_n775));
  OAI21_X1  g574(.A(new_n774), .B1(new_n760), .B2(new_n775), .ZN(G1338gat));
  INV_X1    g575(.A(KEYINPUT53), .ZN(new_n777));
  NOR2_X1   g576(.A1(new_n652), .A2(G106gat), .ZN(new_n778));
  NAND2_X1  g577(.A1(new_n721), .A2(new_n778), .ZN(new_n779));
  AOI21_X1  g578(.A(new_n779), .B1(new_n753), .B2(new_n757), .ZN(new_n780));
  NAND4_X1  g579(.A1(new_n687), .A2(new_n721), .A3(new_n693), .A4(new_n747), .ZN(new_n781));
  NAND2_X1  g580(.A1(new_n781), .A2(G106gat), .ZN(new_n782));
  INV_X1    g581(.A(KEYINPUT111), .ZN(new_n783));
  AOI21_X1  g582(.A(new_n780), .B1(new_n782), .B2(new_n783), .ZN(new_n784));
  NAND3_X1  g583(.A1(new_n781), .A2(KEYINPUT111), .A3(G106gat), .ZN(new_n785));
  AOI21_X1  g584(.A(new_n777), .B1(new_n784), .B2(new_n785), .ZN(new_n786));
  INV_X1    g585(.A(new_n780), .ZN(new_n787));
  XOR2_X1   g586(.A(KEYINPUT112), .B(KEYINPUT53), .Z(new_n788));
  NAND3_X1  g587(.A1(new_n787), .A2(new_n782), .A3(new_n788), .ZN(new_n789));
  INV_X1    g588(.A(new_n789), .ZN(new_n790));
  OAI21_X1  g589(.A(KEYINPUT113), .B1(new_n786), .B2(new_n790), .ZN(new_n791));
  INV_X1    g590(.A(KEYINPUT113), .ZN(new_n792));
  AND3_X1   g591(.A1(new_n781), .A2(KEYINPUT111), .A3(G106gat), .ZN(new_n793));
  AOI21_X1  g592(.A(KEYINPUT111), .B1(new_n781), .B2(G106gat), .ZN(new_n794));
  NOR3_X1   g593(.A1(new_n793), .A2(new_n794), .A3(new_n780), .ZN(new_n795));
  OAI211_X1 g594(.A(new_n792), .B(new_n789), .C1(new_n795), .C2(new_n777), .ZN(new_n796));
  NAND2_X1  g595(.A1(new_n791), .A2(new_n796), .ZN(G1339gat));
  NOR2_X1   g596(.A1(new_n653), .A2(new_n701), .ZN(new_n798));
  NAND2_X1  g597(.A1(new_n638), .A2(new_n641), .ZN(new_n799));
  NAND2_X1  g598(.A1(new_n799), .A2(new_n644), .ZN(new_n800));
  NAND3_X1  g599(.A1(new_n800), .A2(KEYINPUT54), .A3(new_n642), .ZN(new_n801));
  AOI211_X1 g600(.A(new_n644), .B(new_n640), .C1(new_n634), .C2(new_n637), .ZN(new_n802));
  INV_X1    g601(.A(KEYINPUT54), .ZN(new_n803));
  AOI21_X1  g602(.A(new_n649), .B1(new_n802), .B2(new_n803), .ZN(new_n804));
  NAND2_X1  g603(.A1(new_n801), .A2(new_n804), .ZN(new_n805));
  INV_X1    g604(.A(KEYINPUT55), .ZN(new_n806));
  NAND2_X1  g605(.A1(new_n805), .A2(new_n806), .ZN(new_n807));
  NAND3_X1  g606(.A1(new_n801), .A2(KEYINPUT55), .A3(new_n804), .ZN(new_n808));
  NAND3_X1  g607(.A1(new_n807), .A2(new_n651), .A3(new_n808), .ZN(new_n809));
  AOI21_X1  g608(.A(new_n809), .B1(new_n699), .B2(new_n700), .ZN(new_n810));
  NAND2_X1  g609(.A1(new_n522), .A2(new_n525), .ZN(new_n811));
  OAI21_X1  g610(.A(new_n811), .B1(new_n548), .B2(new_n523), .ZN(new_n812));
  NAND2_X1  g611(.A1(new_n812), .A2(new_n489), .ZN(new_n813));
  NAND2_X1  g612(.A1(new_n555), .A2(new_n813), .ZN(new_n814));
  NOR2_X1   g613(.A1(new_n814), .A2(new_n652), .ZN(new_n815));
  OAI21_X1  g614(.A(new_n630), .B1(new_n810), .B2(new_n815), .ZN(new_n816));
  NAND2_X1  g615(.A1(new_n808), .A2(new_n651), .ZN(new_n817));
  AOI21_X1  g616(.A(KEYINPUT55), .B1(new_n801), .B2(new_n804), .ZN(new_n818));
  NOR3_X1   g617(.A1(new_n817), .A2(new_n630), .A3(new_n818), .ZN(new_n819));
  INV_X1    g618(.A(new_n814), .ZN(new_n820));
  AOI21_X1  g619(.A(KEYINPUT114), .B1(new_n819), .B2(new_n820), .ZN(new_n821));
  NAND4_X1  g620(.A1(new_n688), .A2(new_n807), .A3(new_n651), .A4(new_n808), .ZN(new_n822));
  INV_X1    g621(.A(KEYINPUT114), .ZN(new_n823));
  NOR3_X1   g622(.A1(new_n822), .A2(new_n814), .A3(new_n823), .ZN(new_n824));
  NOR2_X1   g623(.A1(new_n821), .A2(new_n824), .ZN(new_n825));
  NAND2_X1  g624(.A1(new_n816), .A2(new_n825), .ZN(new_n826));
  AOI21_X1  g625(.A(new_n798), .B1(new_n826), .B2(new_n587), .ZN(new_n827));
  NOR2_X1   g626(.A1(new_n827), .A2(new_n657), .ZN(new_n828));
  NAND2_X1  g627(.A1(new_n828), .A2(new_n480), .ZN(new_n829));
  NOR2_X1   g628(.A1(new_n829), .A2(new_n768), .ZN(new_n830));
  NAND3_X1  g629(.A1(new_n830), .A2(new_n207), .A3(new_n701), .ZN(new_n831));
  INV_X1    g630(.A(KEYINPUT115), .ZN(new_n832));
  OAI21_X1  g631(.A(new_n832), .B1(new_n827), .B2(new_n721), .ZN(new_n833));
  AOI21_X1  g632(.A(new_n588), .B1(new_n816), .B2(new_n825), .ZN(new_n834));
  OAI211_X1 g633(.A(KEYINPUT115), .B(new_n377), .C1(new_n834), .C2(new_n798), .ZN(new_n835));
  NAND2_X1  g634(.A1(new_n833), .A2(new_n835), .ZN(new_n836));
  NOR2_X1   g635(.A1(new_n657), .A2(new_n768), .ZN(new_n837));
  NAND4_X1  g636(.A1(new_n836), .A2(new_n675), .A3(new_n556), .A4(new_n837), .ZN(new_n838));
  INV_X1    g637(.A(KEYINPUT116), .ZN(new_n839));
  AND3_X1   g638(.A1(new_n838), .A2(new_n839), .A3(G113gat), .ZN(new_n840));
  AOI21_X1  g639(.A(new_n839), .B1(new_n838), .B2(G113gat), .ZN(new_n841));
  OAI21_X1  g640(.A(new_n831), .B1(new_n840), .B2(new_n841), .ZN(new_n842));
  INV_X1    g641(.A(KEYINPUT117), .ZN(new_n843));
  NAND2_X1  g642(.A1(new_n842), .A2(new_n843), .ZN(new_n844));
  OAI211_X1 g643(.A(new_n831), .B(KEYINPUT117), .C1(new_n840), .C2(new_n841), .ZN(new_n845));
  NAND2_X1  g644(.A1(new_n844), .A2(new_n845), .ZN(G1340gat));
  NAND3_X1  g645(.A1(new_n836), .A2(new_n675), .A3(new_n837), .ZN(new_n847));
  NOR3_X1   g646(.A1(new_n847), .A2(new_n205), .A3(new_n652), .ZN(new_n848));
  AOI21_X1  g647(.A(G120gat), .B1(new_n830), .B2(new_n728), .ZN(new_n849));
  NOR2_X1   g648(.A1(new_n848), .A2(new_n849), .ZN(G1341gat));
  OAI21_X1  g649(.A(G127gat), .B1(new_n847), .B2(new_n587), .ZN(new_n851));
  NAND3_X1  g650(.A1(new_n830), .A2(new_n214), .A3(new_n588), .ZN(new_n852));
  NAND2_X1  g651(.A1(new_n851), .A2(new_n852), .ZN(new_n853));
  XNOR2_X1  g652(.A(new_n853), .B(KEYINPUT118), .ZN(G1342gat));
  NOR4_X1   g653(.A1(new_n829), .A2(G134gat), .A3(new_n663), .A4(new_n630), .ZN(new_n855));
  XNOR2_X1  g654(.A(new_n855), .B(KEYINPUT56), .ZN(new_n856));
  OAI21_X1  g655(.A(G134gat), .B1(new_n847), .B2(new_n630), .ZN(new_n857));
  NAND2_X1  g656(.A1(new_n856), .A2(new_n857), .ZN(G1343gat));
  INV_X1    g657(.A(new_n827), .ZN(new_n859));
  INV_X1    g658(.A(KEYINPUT57), .ZN(new_n860));
  NAND3_X1  g659(.A1(new_n859), .A2(new_n860), .A3(new_n721), .ZN(new_n861));
  NOR3_X1   g660(.A1(new_n657), .A2(new_n312), .A3(new_n768), .ZN(new_n862));
  NOR2_X1   g661(.A1(new_n557), .A2(new_n809), .ZN(new_n863));
  OAI21_X1  g662(.A(new_n630), .B1(new_n863), .B2(new_n815), .ZN(new_n864));
  NAND2_X1  g663(.A1(new_n825), .A2(new_n864), .ZN(new_n865));
  AOI21_X1  g664(.A(new_n798), .B1(new_n865), .B2(new_n587), .ZN(new_n866));
  OAI21_X1  g665(.A(KEYINPUT57), .B1(new_n866), .B2(new_n377), .ZN(new_n867));
  NAND3_X1  g666(.A1(new_n861), .A2(new_n862), .A3(new_n867), .ZN(new_n868));
  OAI21_X1  g667(.A(G141gat), .B1(new_n868), .B2(new_n557), .ZN(new_n869));
  NAND2_X1  g668(.A1(new_n673), .A2(new_n721), .ZN(new_n870));
  XNOR2_X1  g669(.A(new_n870), .B(KEYINPUT119), .ZN(new_n871));
  AND2_X1   g670(.A1(new_n871), .A2(new_n828), .ZN(new_n872));
  NOR2_X1   g671(.A1(new_n557), .A2(G141gat), .ZN(new_n873));
  NAND3_X1  g672(.A1(new_n872), .A2(new_n733), .A3(new_n873), .ZN(new_n874));
  XNOR2_X1  g673(.A(KEYINPUT120), .B(KEYINPUT58), .ZN(new_n875));
  NAND3_X1  g674(.A1(new_n869), .A2(new_n874), .A3(new_n875), .ZN(new_n876));
  INV_X1    g675(.A(new_n876), .ZN(new_n877));
  INV_X1    g676(.A(KEYINPUT58), .ZN(new_n878));
  OAI21_X1  g677(.A(G141gat), .B1(new_n868), .B2(new_n702), .ZN(new_n879));
  AOI21_X1  g678(.A(new_n878), .B1(new_n879), .B2(new_n874), .ZN(new_n880));
  OAI21_X1  g679(.A(KEYINPUT121), .B1(new_n877), .B2(new_n880), .ZN(new_n881));
  INV_X1    g680(.A(KEYINPUT121), .ZN(new_n882));
  AND2_X1   g681(.A1(new_n879), .A2(new_n874), .ZN(new_n883));
  OAI211_X1 g682(.A(new_n876), .B(new_n882), .C1(new_n883), .C2(new_n878), .ZN(new_n884));
  NAND2_X1  g683(.A1(new_n881), .A2(new_n884), .ZN(G1344gat));
  AND2_X1   g684(.A1(new_n872), .A2(new_n733), .ZN(new_n886));
  INV_X1    g685(.A(G148gat), .ZN(new_n887));
  NAND3_X1  g686(.A1(new_n886), .A2(new_n887), .A3(new_n728), .ZN(new_n888));
  INV_X1    g687(.A(new_n868), .ZN(new_n889));
  AOI211_X1 g688(.A(KEYINPUT59), .B(new_n887), .C1(new_n889), .C2(new_n728), .ZN(new_n890));
  INV_X1    g689(.A(KEYINPUT59), .ZN(new_n891));
  OAI21_X1  g690(.A(KEYINPUT57), .B1(new_n827), .B2(new_n377), .ZN(new_n892));
  NAND2_X1  g691(.A1(new_n819), .A2(new_n820), .ZN(new_n893));
  AOI21_X1  g692(.A(new_n588), .B1(new_n864), .B2(new_n893), .ZN(new_n894));
  NOR2_X1   g693(.A1(new_n653), .A2(new_n556), .ZN(new_n895));
  OAI211_X1 g694(.A(new_n860), .B(new_n721), .C1(new_n894), .C2(new_n895), .ZN(new_n896));
  AND2_X1   g695(.A1(new_n892), .A2(new_n896), .ZN(new_n897));
  NAND3_X1  g696(.A1(new_n897), .A2(new_n728), .A3(new_n862), .ZN(new_n898));
  AOI21_X1  g697(.A(new_n891), .B1(new_n898), .B2(G148gat), .ZN(new_n899));
  OAI21_X1  g698(.A(new_n888), .B1(new_n890), .B2(new_n899), .ZN(G1345gat));
  NAND3_X1  g699(.A1(new_n886), .A2(new_n322), .A3(new_n588), .ZN(new_n901));
  OAI21_X1  g700(.A(G155gat), .B1(new_n868), .B2(new_n587), .ZN(new_n902));
  NAND2_X1  g701(.A1(new_n901), .A2(new_n902), .ZN(new_n903));
  INV_X1    g702(.A(KEYINPUT122), .ZN(new_n904));
  XNOR2_X1  g703(.A(new_n903), .B(new_n904), .ZN(G1346gat));
  NAND4_X1  g704(.A1(new_n872), .A2(new_n323), .A3(new_n440), .A4(new_n688), .ZN(new_n906));
  INV_X1    g705(.A(KEYINPUT123), .ZN(new_n907));
  OAI21_X1  g706(.A(new_n907), .B1(new_n868), .B2(new_n630), .ZN(new_n908));
  NAND2_X1  g707(.A1(new_n908), .A2(G162gat), .ZN(new_n909));
  NOR3_X1   g708(.A1(new_n868), .A2(new_n907), .A3(new_n630), .ZN(new_n910));
  OAI21_X1  g709(.A(new_n906), .B1(new_n909), .B2(new_n910), .ZN(G1347gat));
  NOR2_X1   g710(.A1(new_n658), .A2(new_n440), .ZN(new_n912));
  NAND3_X1  g711(.A1(new_n836), .A2(new_n675), .A3(new_n912), .ZN(new_n913));
  OAI21_X1  g712(.A(G169gat), .B1(new_n913), .B2(new_n557), .ZN(new_n914));
  NAND2_X1  g713(.A1(new_n859), .A2(new_n657), .ZN(new_n915));
  OR2_X1    g714(.A1(new_n915), .A2(KEYINPUT124), .ZN(new_n916));
  AOI21_X1  g715(.A(new_n733), .B1(new_n915), .B2(KEYINPUT124), .ZN(new_n917));
  NAND2_X1  g716(.A1(new_n916), .A2(new_n917), .ZN(new_n918));
  NOR2_X1   g717(.A1(new_n918), .A2(new_n478), .ZN(new_n919));
  INV_X1    g718(.A(new_n919), .ZN(new_n920));
  NAND2_X1  g719(.A1(new_n701), .A2(new_n260), .ZN(new_n921));
  OAI21_X1  g720(.A(new_n914), .B1(new_n920), .B2(new_n921), .ZN(G1348gat));
  OAI21_X1  g721(.A(G176gat), .B1(new_n913), .B2(new_n652), .ZN(new_n923));
  INV_X1    g722(.A(G176gat), .ZN(new_n924));
  NAND2_X1  g723(.A1(new_n728), .A2(new_n924), .ZN(new_n925));
  OAI21_X1  g724(.A(new_n923), .B1(new_n920), .B2(new_n925), .ZN(G1349gat));
  INV_X1    g725(.A(KEYINPUT60), .ZN(new_n927));
  OAI21_X1  g726(.A(G183gat), .B1(new_n913), .B2(new_n587), .ZN(new_n928));
  NAND2_X1  g727(.A1(new_n588), .A2(new_n249), .ZN(new_n929));
  OAI211_X1 g728(.A(new_n927), .B(new_n928), .C1(new_n920), .C2(new_n929), .ZN(new_n930));
  NOR3_X1   g729(.A1(new_n918), .A2(new_n478), .A3(new_n929), .ZN(new_n931));
  INV_X1    g730(.A(new_n928), .ZN(new_n932));
  OAI21_X1  g731(.A(KEYINPUT60), .B1(new_n931), .B2(new_n932), .ZN(new_n933));
  NAND2_X1  g732(.A1(new_n930), .A2(new_n933), .ZN(G1350gat));
  NAND3_X1  g733(.A1(new_n919), .A2(new_n240), .A3(new_n688), .ZN(new_n935));
  INV_X1    g734(.A(KEYINPUT61), .ZN(new_n936));
  INV_X1    g735(.A(new_n913), .ZN(new_n937));
  NAND2_X1  g736(.A1(new_n937), .A2(new_n688), .ZN(new_n938));
  AOI21_X1  g737(.A(new_n936), .B1(new_n938), .B2(G190gat), .ZN(new_n939));
  AOI211_X1 g738(.A(KEYINPUT61), .B(new_n240), .C1(new_n937), .C2(new_n688), .ZN(new_n940));
  OAI21_X1  g739(.A(new_n935), .B1(new_n939), .B2(new_n940), .ZN(G1351gat));
  NOR2_X1   g740(.A1(new_n918), .A2(new_n870), .ZN(new_n942));
  AOI21_X1  g741(.A(G197gat), .B1(new_n942), .B2(new_n701), .ZN(new_n943));
  INV_X1    g742(.A(KEYINPUT125), .ZN(new_n944));
  NAND2_X1  g743(.A1(new_n897), .A2(new_n944), .ZN(new_n945));
  NOR3_X1   g744(.A1(new_n658), .A2(new_n440), .A3(new_n312), .ZN(new_n946));
  NAND2_X1  g745(.A1(new_n892), .A2(new_n896), .ZN(new_n947));
  NAND2_X1  g746(.A1(new_n947), .A2(KEYINPUT125), .ZN(new_n948));
  AND3_X1   g747(.A1(new_n945), .A2(new_n946), .A3(new_n948), .ZN(new_n949));
  AND2_X1   g748(.A1(new_n556), .A2(G197gat), .ZN(new_n950));
  AOI21_X1  g749(.A(new_n943), .B1(new_n949), .B2(new_n950), .ZN(G1352gat));
  NAND2_X1  g750(.A1(new_n949), .A2(new_n728), .ZN(new_n952));
  NAND2_X1  g751(.A1(new_n952), .A2(G204gat), .ZN(new_n953));
  NOR2_X1   g752(.A1(new_n652), .A2(G204gat), .ZN(new_n954));
  NAND2_X1  g753(.A1(new_n942), .A2(new_n954), .ZN(new_n955));
  NAND2_X1  g754(.A1(new_n955), .A2(KEYINPUT62), .ZN(new_n956));
  INV_X1    g755(.A(KEYINPUT62), .ZN(new_n957));
  NAND3_X1  g756(.A1(new_n942), .A2(new_n957), .A3(new_n954), .ZN(new_n958));
  NAND3_X1  g757(.A1(new_n953), .A2(new_n956), .A3(new_n958), .ZN(G1353gat));
  INV_X1    g758(.A(new_n870), .ZN(new_n960));
  NOR2_X1   g759(.A1(new_n587), .A2(G211gat), .ZN(new_n961));
  NAND4_X1  g760(.A1(new_n916), .A2(new_n917), .A3(new_n960), .A4(new_n961), .ZN(new_n962));
  NAND4_X1  g761(.A1(new_n892), .A2(new_n588), .A3(new_n896), .A4(new_n946), .ZN(new_n963));
  AND3_X1   g762(.A1(new_n963), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n964));
  AOI21_X1  g763(.A(KEYINPUT63), .B1(new_n963), .B2(G211gat), .ZN(new_n965));
  OAI21_X1  g764(.A(new_n962), .B1(new_n964), .B2(new_n965), .ZN(new_n966));
  INV_X1    g765(.A(KEYINPUT126), .ZN(new_n967));
  XNOR2_X1  g766(.A(new_n966), .B(new_n967), .ZN(G1354gat));
  NAND3_X1  g767(.A1(new_n916), .A2(new_n960), .A3(new_n917), .ZN(new_n969));
  OAI21_X1  g768(.A(new_n341), .B1(new_n969), .B2(new_n630), .ZN(new_n970));
  NOR2_X1   g769(.A1(new_n630), .A2(new_n341), .ZN(new_n971));
  NAND4_X1  g770(.A1(new_n945), .A2(new_n946), .A3(new_n948), .A4(new_n971), .ZN(new_n972));
  NAND2_X1  g771(.A1(new_n970), .A2(new_n972), .ZN(new_n973));
  NAND2_X1  g772(.A1(new_n973), .A2(KEYINPUT127), .ZN(new_n974));
  INV_X1    g773(.A(KEYINPUT127), .ZN(new_n975));
  NAND3_X1  g774(.A1(new_n970), .A2(new_n972), .A3(new_n975), .ZN(new_n976));
  NAND2_X1  g775(.A1(new_n974), .A2(new_n976), .ZN(G1355gat));
endmodule


