//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 1 0 0 0 1 0 0 1 0 1 0 1 1 0 1 0 1 0 1 0 1 0 1 0 1 0 1 0 0 0 1 1 0 1 0 0 1 0 0 1 0 0 1 0 1 1 0 0 0 0 1 0 1 0 0 0 1 0 1 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:31:16 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n442, new_n447, new_n451, new_n452, new_n453, new_n456, new_n457,
    new_n458, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n523, new_n524, new_n525,
    new_n526, new_n527, new_n528, new_n529, new_n530, new_n531, new_n532,
    new_n533, new_n534, new_n535, new_n536, new_n537, new_n538, new_n539,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n560, new_n561, new_n563, new_n564, new_n565, new_n566, new_n567,
    new_n568, new_n569, new_n570, new_n571, new_n572, new_n573, new_n574,
    new_n575, new_n576, new_n577, new_n578, new_n579, new_n580, new_n581,
    new_n582, new_n583, new_n584, new_n585, new_n586, new_n587, new_n589,
    new_n590, new_n591, new_n592, new_n593, new_n594, new_n596, new_n597,
    new_n598, new_n599, new_n601, new_n602, new_n603, new_n604, new_n605,
    new_n606, new_n607, new_n608, new_n609, new_n610, new_n611, new_n612,
    new_n614, new_n615, new_n616, new_n617, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n636, new_n637,
    new_n638, new_n641, new_n642, new_n644, new_n645, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n677, new_n678,
    new_n679, new_n680, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n692, new_n693,
    new_n694, new_n695, new_n696, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n713, new_n714, new_n715,
    new_n716, new_n717, new_n718, new_n719, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n851, new_n852, new_n853, new_n854, new_n855, new_n856,
    new_n857, new_n859, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1213, new_n1214;
  XNOR2_X1  g000(.A(KEYINPUT64), .B(G452), .ZN(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  XOR2_X1   g002(.A(KEYINPUT65), .B(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  XNOR2_X1  g007(.A(KEYINPUT66), .B(G2066), .ZN(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  XNOR2_X1  g015(.A(KEYINPUT67), .B(G108), .ZN(G238));
  AND2_X1   g016(.A1(G2072), .A2(G2078), .ZN(new_n442));
  NAND3_X1  g017(.A1(new_n442), .A2(G2084), .A3(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g025(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n451));
  XNOR2_X1  g026(.A(new_n451), .B(KEYINPUT2), .ZN(new_n452));
  NOR4_X1   g027(.A1(G238), .A2(G237), .A3(G235), .A4(G236), .ZN(new_n453));
  NAND2_X1  g028(.A1(new_n452), .A2(new_n453), .ZN(G261));
  INV_X1    g029(.A(G261), .ZN(G325));
  INV_X1    g030(.A(G567), .ZN(new_n456));
  NOR2_X1   g031(.A1(new_n453), .A2(new_n456), .ZN(new_n457));
  INV_X1    g032(.A(new_n452), .ZN(new_n458));
  AOI21_X1  g033(.A(new_n457), .B1(new_n458), .B2(G2106), .ZN(G319));
  INV_X1    g034(.A(G2105), .ZN(new_n460));
  NAND2_X1  g035(.A1(G113), .A2(G2104), .ZN(new_n461));
  INV_X1    g036(.A(new_n461), .ZN(new_n462));
  AND2_X1   g037(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n463));
  NOR2_X1   g038(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n464));
  OAI21_X1  g039(.A(G125), .B1(new_n463), .B2(new_n464), .ZN(new_n465));
  AOI21_X1  g040(.A(new_n462), .B1(new_n465), .B2(KEYINPUT68), .ZN(new_n466));
  INV_X1    g041(.A(KEYINPUT68), .ZN(new_n467));
  OAI211_X1 g042(.A(new_n467), .B(G125), .C1(new_n463), .C2(new_n464), .ZN(new_n468));
  AOI21_X1  g043(.A(new_n460), .B1(new_n466), .B2(new_n468), .ZN(new_n469));
  NAND2_X1  g044(.A1(G101), .A2(G2104), .ZN(new_n470));
  NOR2_X1   g045(.A1(new_n463), .A2(new_n464), .ZN(new_n471));
  INV_X1    g046(.A(G137), .ZN(new_n472));
  OAI21_X1  g047(.A(new_n470), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  AOI21_X1  g048(.A(new_n469), .B1(new_n460), .B2(new_n473), .ZN(G160));
  OAI21_X1  g049(.A(new_n460), .B1(new_n463), .B2(new_n464), .ZN(new_n475));
  INV_X1    g050(.A(new_n475), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n476), .A2(G136), .ZN(new_n477));
  INV_X1    g052(.A(KEYINPUT69), .ZN(new_n478));
  XNOR2_X1  g053(.A(new_n477), .B(new_n478), .ZN(new_n479));
  NOR2_X1   g054(.A1(new_n471), .A2(new_n460), .ZN(new_n480));
  OR2_X1    g055(.A1(G100), .A2(G2105), .ZN(new_n481));
  INV_X1    g056(.A(G2104), .ZN(new_n482));
  INV_X1    g057(.A(G112), .ZN(new_n483));
  AOI21_X1  g058(.A(new_n482), .B1(new_n483), .B2(G2105), .ZN(new_n484));
  AOI22_X1  g059(.A1(new_n480), .A2(G124), .B1(new_n481), .B2(new_n484), .ZN(new_n485));
  AND2_X1   g060(.A1(new_n479), .A2(new_n485), .ZN(G162));
  NOR2_X1   g061(.A1(KEYINPUT72), .A2(KEYINPUT4), .ZN(new_n487));
  NAND2_X1  g062(.A1(KEYINPUT72), .A2(KEYINPUT4), .ZN(new_n488));
  NAND2_X1  g063(.A1(new_n488), .A2(G138), .ZN(new_n489));
  OAI21_X1  g064(.A(new_n487), .B1(new_n475), .B2(new_n489), .ZN(new_n490));
  INV_X1    g065(.A(KEYINPUT3), .ZN(new_n491));
  NAND2_X1  g066(.A1(new_n491), .A2(new_n482), .ZN(new_n492));
  NAND2_X1  g067(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n493));
  NAND2_X1  g068(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  AND2_X1   g069(.A1(new_n488), .A2(G138), .ZN(new_n495));
  INV_X1    g070(.A(new_n487), .ZN(new_n496));
  NAND4_X1  g071(.A1(new_n494), .A2(new_n495), .A3(new_n460), .A4(new_n496), .ZN(new_n497));
  NAND2_X1  g072(.A1(new_n490), .A2(new_n497), .ZN(new_n498));
  OR2_X1    g073(.A1(G102), .A2(G2105), .ZN(new_n499));
  OAI21_X1  g074(.A(G2105), .B1(KEYINPUT70), .B2(G114), .ZN(new_n500));
  AND2_X1   g075(.A1(KEYINPUT70), .A2(G114), .ZN(new_n501));
  OAI211_X1 g076(.A(G2104), .B(new_n499), .C1(new_n500), .C2(new_n501), .ZN(new_n502));
  OAI211_X1 g077(.A(G126), .B(G2105), .C1(new_n463), .C2(new_n464), .ZN(new_n503));
  NAND2_X1  g078(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  NAND2_X1  g079(.A1(new_n504), .A2(KEYINPUT71), .ZN(new_n505));
  INV_X1    g080(.A(KEYINPUT71), .ZN(new_n506));
  NAND3_X1  g081(.A1(new_n502), .A2(new_n503), .A3(new_n506), .ZN(new_n507));
  AOI21_X1  g082(.A(new_n498), .B1(new_n505), .B2(new_n507), .ZN(G164));
  INV_X1    g083(.A(G651), .ZN(new_n509));
  AND2_X1   g084(.A1(KEYINPUT5), .A2(G543), .ZN(new_n510));
  NOR2_X1   g085(.A1(KEYINPUT5), .A2(G543), .ZN(new_n511));
  OAI21_X1  g086(.A(G62), .B1(new_n510), .B2(new_n511), .ZN(new_n512));
  NAND2_X1  g087(.A1(G75), .A2(G543), .ZN(new_n513));
  AOI21_X1  g088(.A(new_n509), .B1(new_n512), .B2(new_n513), .ZN(new_n514));
  NAND2_X1  g089(.A1(new_n509), .A2(KEYINPUT6), .ZN(new_n515));
  INV_X1    g090(.A(KEYINPUT6), .ZN(new_n516));
  NAND2_X1  g091(.A1(new_n516), .A2(G651), .ZN(new_n517));
  NAND2_X1  g092(.A1(new_n515), .A2(new_n517), .ZN(new_n518));
  OAI21_X1  g093(.A(G88), .B1(new_n510), .B2(new_n511), .ZN(new_n519));
  NAND2_X1  g094(.A1(G50), .A2(G543), .ZN(new_n520));
  AOI21_X1  g095(.A(new_n518), .B1(new_n519), .B2(new_n520), .ZN(new_n521));
  NOR2_X1   g096(.A1(new_n514), .A2(new_n521), .ZN(G166));
  INV_X1    g097(.A(G543), .ZN(new_n523));
  AOI21_X1  g098(.A(new_n523), .B1(new_n518), .B2(KEYINPUT73), .ZN(new_n524));
  XNOR2_X1  g099(.A(KEYINPUT6), .B(G651), .ZN(new_n525));
  INV_X1    g100(.A(KEYINPUT73), .ZN(new_n526));
  NAND2_X1  g101(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  AND2_X1   g102(.A1(new_n524), .A2(new_n527), .ZN(new_n528));
  NAND2_X1  g103(.A1(new_n528), .A2(G51), .ZN(new_n529));
  OR2_X1    g104(.A1(KEYINPUT5), .A2(G543), .ZN(new_n530));
  NAND2_X1  g105(.A1(KEYINPUT5), .A2(G543), .ZN(new_n531));
  NAND2_X1  g106(.A1(new_n530), .A2(new_n531), .ZN(new_n532));
  NAND2_X1  g107(.A1(new_n532), .A2(new_n525), .ZN(new_n533));
  INV_X1    g108(.A(new_n533), .ZN(new_n534));
  NAND2_X1  g109(.A1(new_n534), .A2(G89), .ZN(new_n535));
  NAND3_X1  g110(.A1(new_n532), .A2(G63), .A3(G651), .ZN(new_n536));
  NAND3_X1  g111(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n537));
  XNOR2_X1  g112(.A(new_n537), .B(KEYINPUT7), .ZN(new_n538));
  AND2_X1   g113(.A1(new_n536), .A2(new_n538), .ZN(new_n539));
  NAND3_X1  g114(.A1(new_n529), .A2(new_n535), .A3(new_n539), .ZN(G286));
  INV_X1    g115(.A(G286), .ZN(G168));
  XOR2_X1   g116(.A(KEYINPUT74), .B(G52), .Z(new_n542));
  NAND2_X1  g117(.A1(new_n528), .A2(new_n542), .ZN(new_n543));
  NAND2_X1  g118(.A1(G77), .A2(G543), .ZN(new_n544));
  NOR2_X1   g119(.A1(new_n510), .A2(new_n511), .ZN(new_n545));
  INV_X1    g120(.A(G64), .ZN(new_n546));
  OAI21_X1  g121(.A(new_n544), .B1(new_n545), .B2(new_n546), .ZN(new_n547));
  AOI22_X1  g122(.A1(new_n534), .A2(G90), .B1(new_n547), .B2(G651), .ZN(new_n548));
  NAND2_X1  g123(.A1(new_n543), .A2(new_n548), .ZN(G301));
  INV_X1    g124(.A(G301), .ZN(G171));
  NAND2_X1  g125(.A1(new_n528), .A2(G43), .ZN(new_n551));
  NAND2_X1  g126(.A1(G68), .A2(G543), .ZN(new_n552));
  INV_X1    g127(.A(G56), .ZN(new_n553));
  OAI21_X1  g128(.A(new_n552), .B1(new_n545), .B2(new_n553), .ZN(new_n554));
  AOI22_X1  g129(.A1(new_n534), .A2(G81), .B1(new_n554), .B2(G651), .ZN(new_n555));
  NAND2_X1  g130(.A1(new_n551), .A2(new_n555), .ZN(new_n556));
  INV_X1    g131(.A(new_n556), .ZN(new_n557));
  NAND2_X1  g132(.A1(new_n557), .A2(G860), .ZN(G153));
  NAND4_X1  g133(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g134(.A1(G1), .A2(G3), .ZN(new_n560));
  XNOR2_X1  g135(.A(new_n560), .B(KEYINPUT8), .ZN(new_n561));
  NAND4_X1  g136(.A1(G319), .A2(G483), .A3(G661), .A4(new_n561), .ZN(G188));
  XOR2_X1   g137(.A(KEYINPUT76), .B(G65), .Z(new_n563));
  AOI22_X1  g138(.A1(new_n563), .A2(new_n532), .B1(G78), .B2(G543), .ZN(new_n564));
  OAI21_X1  g139(.A(G651), .B1(new_n564), .B2(KEYINPUT77), .ZN(new_n565));
  NAND2_X1  g140(.A1(G78), .A2(G543), .ZN(new_n566));
  XNOR2_X1  g141(.A(KEYINPUT76), .B(G65), .ZN(new_n567));
  OAI21_X1  g142(.A(new_n566), .B1(new_n545), .B2(new_n567), .ZN(new_n568));
  INV_X1    g143(.A(KEYINPUT77), .ZN(new_n569));
  NOR2_X1   g144(.A1(new_n568), .A2(new_n569), .ZN(new_n570));
  INV_X1    g145(.A(KEYINPUT9), .ZN(new_n571));
  NAND3_X1  g146(.A1(new_n524), .A2(G53), .A3(new_n527), .ZN(new_n572));
  OAI22_X1  g147(.A1(new_n565), .A2(new_n570), .B1(new_n571), .B2(new_n572), .ZN(new_n573));
  NAND2_X1  g148(.A1(new_n572), .A2(new_n571), .ZN(new_n574));
  INV_X1    g149(.A(G91), .ZN(new_n575));
  OAI21_X1  g150(.A(KEYINPUT75), .B1(new_n533), .B2(new_n575), .ZN(new_n576));
  INV_X1    g151(.A(KEYINPUT75), .ZN(new_n577));
  NAND4_X1  g152(.A1(new_n532), .A2(new_n525), .A3(new_n577), .A4(G91), .ZN(new_n578));
  NAND2_X1  g153(.A1(new_n576), .A2(new_n578), .ZN(new_n579));
  NAND2_X1  g154(.A1(new_n574), .A2(new_n579), .ZN(new_n580));
  OAI21_X1  g155(.A(KEYINPUT78), .B1(new_n573), .B2(new_n580), .ZN(new_n581));
  AOI22_X1  g156(.A1(new_n571), .A2(new_n572), .B1(new_n576), .B2(new_n578), .ZN(new_n582));
  AOI21_X1  g157(.A(new_n509), .B1(new_n568), .B2(new_n569), .ZN(new_n583));
  OAI21_X1  g158(.A(new_n583), .B1(new_n569), .B2(new_n568), .ZN(new_n584));
  NAND3_X1  g159(.A1(new_n528), .A2(KEYINPUT9), .A3(G53), .ZN(new_n585));
  INV_X1    g160(.A(KEYINPUT78), .ZN(new_n586));
  NAND4_X1  g161(.A1(new_n582), .A2(new_n584), .A3(new_n585), .A4(new_n586), .ZN(new_n587));
  NAND2_X1  g162(.A1(new_n581), .A2(new_n587), .ZN(G299));
  INV_X1    g163(.A(new_n514), .ZN(new_n589));
  NAND2_X1  g164(.A1(new_n519), .A2(new_n520), .ZN(new_n590));
  NAND2_X1  g165(.A1(new_n590), .A2(new_n525), .ZN(new_n591));
  INV_X1    g166(.A(KEYINPUT79), .ZN(new_n592));
  NAND3_X1  g167(.A1(new_n589), .A2(new_n591), .A3(new_n592), .ZN(new_n593));
  OAI21_X1  g168(.A(KEYINPUT79), .B1(new_n514), .B2(new_n521), .ZN(new_n594));
  AND2_X1   g169(.A1(new_n593), .A2(new_n594), .ZN(G303));
  OAI21_X1  g170(.A(G651), .B1(new_n532), .B2(G74), .ZN(new_n596));
  NAND3_X1  g171(.A1(new_n532), .A2(new_n525), .A3(G87), .ZN(new_n597));
  AND2_X1   g172(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  NAND3_X1  g173(.A1(new_n524), .A2(G49), .A3(new_n527), .ZN(new_n599));
  NAND2_X1  g174(.A1(new_n598), .A2(new_n599), .ZN(G288));
  OAI21_X1  g175(.A(G86), .B1(new_n510), .B2(new_n511), .ZN(new_n601));
  NAND2_X1  g176(.A1(G48), .A2(G543), .ZN(new_n602));
  NAND2_X1  g177(.A1(new_n601), .A2(new_n602), .ZN(new_n603));
  NAND2_X1  g178(.A1(new_n603), .A2(new_n525), .ZN(new_n604));
  INV_X1    g179(.A(G61), .ZN(new_n605));
  AOI21_X1  g180(.A(new_n605), .B1(new_n530), .B2(new_n531), .ZN(new_n606));
  NAND2_X1  g181(.A1(G73), .A2(G543), .ZN(new_n607));
  INV_X1    g182(.A(KEYINPUT80), .ZN(new_n608));
  NAND2_X1  g183(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  NAND3_X1  g184(.A1(KEYINPUT80), .A2(G73), .A3(G543), .ZN(new_n610));
  NAND2_X1  g185(.A1(new_n609), .A2(new_n610), .ZN(new_n611));
  OAI21_X1  g186(.A(G651), .B1(new_n606), .B2(new_n611), .ZN(new_n612));
  NAND2_X1  g187(.A1(new_n604), .A2(new_n612), .ZN(G305));
  NAND2_X1  g188(.A1(new_n534), .A2(G85), .ZN(new_n614));
  AOI22_X1  g189(.A1(new_n532), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n615));
  NAND2_X1  g190(.A1(new_n524), .A2(new_n527), .ZN(new_n616));
  INV_X1    g191(.A(G47), .ZN(new_n617));
  OAI221_X1 g192(.A(new_n614), .B1(new_n509), .B2(new_n615), .C1(new_n616), .C2(new_n617), .ZN(G290));
  NAND2_X1  g193(.A1(G301), .A2(G868), .ZN(new_n619));
  NAND2_X1  g194(.A1(G79), .A2(G543), .ZN(new_n620));
  INV_X1    g195(.A(G66), .ZN(new_n621));
  OAI21_X1  g196(.A(new_n620), .B1(new_n545), .B2(new_n621), .ZN(new_n622));
  NAND2_X1  g197(.A1(new_n622), .A2(G651), .ZN(new_n623));
  INV_X1    g198(.A(G54), .ZN(new_n624));
  OAI21_X1  g199(.A(new_n623), .B1(new_n616), .B2(new_n624), .ZN(new_n625));
  NAND2_X1  g200(.A1(new_n625), .A2(KEYINPUT81), .ZN(new_n626));
  INV_X1    g201(.A(KEYINPUT81), .ZN(new_n627));
  OAI211_X1 g202(.A(new_n623), .B(new_n627), .C1(new_n616), .C2(new_n624), .ZN(new_n628));
  INV_X1    g203(.A(G92), .ZN(new_n629));
  NOR2_X1   g204(.A1(new_n533), .A2(new_n629), .ZN(new_n630));
  OR2_X1    g205(.A1(new_n630), .A2(KEYINPUT10), .ZN(new_n631));
  NAND2_X1  g206(.A1(new_n630), .A2(KEYINPUT10), .ZN(new_n632));
  AOI22_X1  g207(.A1(new_n626), .A2(new_n628), .B1(new_n631), .B2(new_n632), .ZN(new_n633));
  OAI21_X1  g208(.A(new_n619), .B1(new_n633), .B2(G868), .ZN(G284));
  OAI21_X1  g209(.A(new_n619), .B1(new_n633), .B2(G868), .ZN(G321));
  INV_X1    g210(.A(G868), .ZN(new_n636));
  NOR2_X1   g211(.A1(G286), .A2(new_n636), .ZN(new_n637));
  INV_X1    g212(.A(G299), .ZN(new_n638));
  AOI21_X1  g213(.A(new_n637), .B1(new_n638), .B2(new_n636), .ZN(G297));
  AOI21_X1  g214(.A(new_n637), .B1(new_n638), .B2(new_n636), .ZN(G280));
  INV_X1    g215(.A(G559), .ZN(new_n641));
  OAI21_X1  g216(.A(new_n633), .B1(new_n641), .B2(G860), .ZN(new_n642));
  XNOR2_X1  g217(.A(new_n642), .B(KEYINPUT82), .ZN(G148));
  NAND2_X1  g218(.A1(new_n633), .A2(new_n641), .ZN(new_n644));
  NAND2_X1  g219(.A1(new_n644), .A2(G868), .ZN(new_n645));
  OAI21_X1  g220(.A(new_n645), .B1(G868), .B2(new_n557), .ZN(G323));
  XNOR2_X1  g221(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND3_X1  g222(.A1(new_n460), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n648));
  XOR2_X1   g223(.A(new_n648), .B(KEYINPUT12), .Z(new_n649));
  XOR2_X1   g224(.A(new_n649), .B(KEYINPUT13), .Z(new_n650));
  INV_X1    g225(.A(G2100), .ZN(new_n651));
  OR2_X1    g226(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  OR2_X1    g227(.A1(G99), .A2(G2105), .ZN(new_n653));
  INV_X1    g228(.A(G111), .ZN(new_n654));
  AOI21_X1  g229(.A(new_n482), .B1(new_n654), .B2(G2105), .ZN(new_n655));
  AOI22_X1  g230(.A1(new_n476), .A2(G135), .B1(new_n653), .B2(new_n655), .ZN(new_n656));
  AND3_X1   g231(.A1(new_n480), .A2(KEYINPUT83), .A3(G123), .ZN(new_n657));
  AOI21_X1  g232(.A(KEYINPUT83), .B1(new_n480), .B2(G123), .ZN(new_n658));
  OAI21_X1  g233(.A(new_n656), .B1(new_n657), .B2(new_n658), .ZN(new_n659));
  INV_X1    g234(.A(G2096), .ZN(new_n660));
  XNOR2_X1  g235(.A(new_n659), .B(new_n660), .ZN(new_n661));
  NAND2_X1  g236(.A1(new_n650), .A2(new_n651), .ZN(new_n662));
  NAND3_X1  g237(.A1(new_n652), .A2(new_n661), .A3(new_n662), .ZN(G156));
  XNOR2_X1  g238(.A(G2451), .B(G2454), .ZN(new_n664));
  XNOR2_X1  g239(.A(new_n664), .B(KEYINPUT16), .ZN(new_n665));
  XOR2_X1   g240(.A(G2443), .B(G2446), .Z(new_n666));
  XNOR2_X1  g241(.A(new_n665), .B(new_n666), .ZN(new_n667));
  XOR2_X1   g242(.A(G1341), .B(G1348), .Z(new_n668));
  XNOR2_X1  g243(.A(new_n668), .B(KEYINPUT85), .ZN(new_n669));
  XNOR2_X1  g244(.A(new_n667), .B(new_n669), .ZN(new_n670));
  XNOR2_X1  g245(.A(G2427), .B(G2430), .ZN(new_n671));
  XNOR2_X1  g246(.A(KEYINPUT84), .B(G2438), .ZN(new_n672));
  XNOR2_X1  g247(.A(new_n671), .B(new_n672), .ZN(new_n673));
  XNOR2_X1  g248(.A(KEYINPUT15), .B(G2435), .ZN(new_n674));
  OR2_X1    g249(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  NAND2_X1  g250(.A1(new_n673), .A2(new_n674), .ZN(new_n676));
  AND3_X1   g251(.A1(new_n675), .A2(KEYINPUT14), .A3(new_n676), .ZN(new_n677));
  OR2_X1    g252(.A1(new_n670), .A2(new_n677), .ZN(new_n678));
  NAND2_X1  g253(.A1(new_n670), .A2(new_n677), .ZN(new_n679));
  NAND3_X1  g254(.A1(new_n678), .A2(G14), .A3(new_n679), .ZN(new_n680));
  INV_X1    g255(.A(new_n680), .ZN(G401));
  XOR2_X1   g256(.A(G2084), .B(G2090), .Z(new_n682));
  XNOR2_X1  g257(.A(G2067), .B(G2678), .ZN(new_n683));
  XNOR2_X1  g258(.A(new_n683), .B(KEYINPUT87), .ZN(new_n684));
  NOR2_X1   g259(.A1(G2072), .A2(G2078), .ZN(new_n685));
  NOR2_X1   g260(.A1(new_n442), .A2(new_n685), .ZN(new_n686));
  AOI21_X1  g261(.A(new_n682), .B1(new_n684), .B2(new_n686), .ZN(new_n687));
  XNOR2_X1  g262(.A(new_n686), .B(KEYINPUT17), .ZN(new_n688));
  OAI21_X1  g263(.A(new_n687), .B1(new_n684), .B2(new_n688), .ZN(new_n689));
  NAND3_X1  g264(.A1(new_n688), .A2(new_n684), .A3(new_n682), .ZN(new_n690));
  OAI211_X1 g265(.A(new_n682), .B(new_n683), .C1(new_n442), .C2(new_n685), .ZN(new_n691));
  XOR2_X1   g266(.A(KEYINPUT86), .B(KEYINPUT18), .Z(new_n692));
  XNOR2_X1  g267(.A(new_n691), .B(new_n692), .ZN(new_n693));
  NAND3_X1  g268(.A1(new_n689), .A2(new_n690), .A3(new_n693), .ZN(new_n694));
  XNOR2_X1  g269(.A(new_n694), .B(new_n660), .ZN(new_n695));
  XNOR2_X1  g270(.A(new_n695), .B(new_n651), .ZN(new_n696));
  INV_X1    g271(.A(new_n696), .ZN(G227));
  XNOR2_X1  g272(.A(G1971), .B(G1976), .ZN(new_n698));
  INV_X1    g273(.A(KEYINPUT19), .ZN(new_n699));
  XNOR2_X1  g274(.A(new_n698), .B(new_n699), .ZN(new_n700));
  XOR2_X1   g275(.A(G1956), .B(G2474), .Z(new_n701));
  XOR2_X1   g276(.A(G1961), .B(G1966), .Z(new_n702));
  NOR2_X1   g277(.A1(new_n701), .A2(new_n702), .ZN(new_n703));
  NAND2_X1  g278(.A1(new_n700), .A2(new_n703), .ZN(new_n704));
  AND2_X1   g279(.A1(new_n701), .A2(new_n702), .ZN(new_n705));
  NAND2_X1  g280(.A1(new_n700), .A2(new_n705), .ZN(new_n706));
  XOR2_X1   g281(.A(KEYINPUT88), .B(KEYINPUT20), .Z(new_n707));
  OR2_X1    g282(.A1(new_n705), .A2(new_n703), .ZN(new_n708));
  OAI221_X1 g283(.A(new_n704), .B1(new_n706), .B2(new_n707), .C1(new_n708), .C2(new_n700), .ZN(new_n709));
  AOI21_X1  g284(.A(new_n709), .B1(new_n706), .B2(new_n707), .ZN(new_n710));
  XNOR2_X1  g285(.A(G1981), .B(G1986), .ZN(new_n711));
  XNOR2_X1  g286(.A(new_n711), .B(KEYINPUT89), .ZN(new_n712));
  XNOR2_X1  g287(.A(new_n710), .B(new_n712), .ZN(new_n713));
  XOR2_X1   g288(.A(G1991), .B(G1996), .Z(new_n714));
  XNOR2_X1  g289(.A(new_n713), .B(new_n714), .ZN(new_n715));
  XNOR2_X1  g290(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n716));
  INV_X1    g291(.A(new_n716), .ZN(new_n717));
  OR2_X1    g292(.A1(new_n715), .A2(new_n717), .ZN(new_n718));
  NAND2_X1  g293(.A1(new_n715), .A2(new_n717), .ZN(new_n719));
  NAND2_X1  g294(.A1(new_n718), .A2(new_n719), .ZN(G229));
  INV_X1    g295(.A(G16), .ZN(new_n721));
  NAND2_X1  g296(.A1(new_n721), .A2(G20), .ZN(new_n722));
  XNOR2_X1  g297(.A(new_n722), .B(KEYINPUT23), .ZN(new_n723));
  OAI21_X1  g298(.A(new_n723), .B1(new_n638), .B2(new_n721), .ZN(new_n724));
  INV_X1    g299(.A(G1956), .ZN(new_n725));
  XNOR2_X1  g300(.A(new_n724), .B(new_n725), .ZN(new_n726));
  INV_X1    g301(.A(G29), .ZN(new_n727));
  NAND2_X1  g302(.A1(new_n727), .A2(G35), .ZN(new_n728));
  XOR2_X1   g303(.A(new_n728), .B(KEYINPUT101), .Z(new_n729));
  OAI21_X1  g304(.A(new_n729), .B1(G162), .B2(new_n727), .ZN(new_n730));
  XNOR2_X1  g305(.A(new_n730), .B(KEYINPUT29), .ZN(new_n731));
  AND2_X1   g306(.A1(new_n731), .A2(G2090), .ZN(new_n732));
  NOR2_X1   g307(.A1(new_n659), .A2(new_n727), .ZN(new_n733));
  INV_X1    g308(.A(KEYINPUT30), .ZN(new_n734));
  AND2_X1   g309(.A1(new_n734), .A2(G28), .ZN(new_n735));
  OAI21_X1  g310(.A(new_n727), .B1(new_n734), .B2(G28), .ZN(new_n736));
  AND2_X1   g311(.A1(KEYINPUT31), .A2(G11), .ZN(new_n737));
  NOR2_X1   g312(.A1(KEYINPUT31), .A2(G11), .ZN(new_n738));
  OAI22_X1  g313(.A1(new_n735), .A2(new_n736), .B1(new_n737), .B2(new_n738), .ZN(new_n739));
  NOR2_X1   g314(.A1(new_n733), .A2(new_n739), .ZN(new_n740));
  NAND2_X1  g315(.A1(new_n727), .A2(G33), .ZN(new_n741));
  NAND3_X1  g316(.A1(new_n460), .A2(G103), .A3(G2104), .ZN(new_n742));
  XOR2_X1   g317(.A(new_n742), .B(KEYINPUT25), .Z(new_n743));
  INV_X1    g318(.A(G139), .ZN(new_n744));
  OAI21_X1  g319(.A(new_n743), .B1(new_n744), .B2(new_n475), .ZN(new_n745));
  NAND2_X1  g320(.A1(new_n494), .A2(G127), .ZN(new_n746));
  NAND2_X1  g321(.A1(G115), .A2(G2104), .ZN(new_n747));
  AOI21_X1  g322(.A(new_n460), .B1(new_n746), .B2(new_n747), .ZN(new_n748));
  NOR2_X1   g323(.A1(new_n745), .A2(new_n748), .ZN(new_n749));
  OAI21_X1  g324(.A(new_n741), .B1(new_n749), .B2(new_n727), .ZN(new_n750));
  OAI21_X1  g325(.A(new_n740), .B1(G2072), .B2(new_n750), .ZN(new_n751));
  NAND2_X1  g326(.A1(new_n721), .A2(G19), .ZN(new_n752));
  OAI21_X1  g327(.A(new_n752), .B1(new_n557), .B2(new_n721), .ZN(new_n753));
  AOI21_X1  g328(.A(new_n751), .B1(G1341), .B2(new_n753), .ZN(new_n754));
  NAND2_X1  g329(.A1(new_n727), .A2(G26), .ZN(new_n755));
  XNOR2_X1  g330(.A(new_n755), .B(KEYINPUT28), .ZN(new_n756));
  NAND2_X1  g331(.A1(new_n480), .A2(G128), .ZN(new_n757));
  NAND2_X1  g332(.A1(new_n476), .A2(G140), .ZN(new_n758));
  OR2_X1    g333(.A1(G104), .A2(G2105), .ZN(new_n759));
  OAI211_X1 g334(.A(new_n759), .B(G2104), .C1(G116), .C2(new_n460), .ZN(new_n760));
  NAND3_X1  g335(.A1(new_n757), .A2(new_n758), .A3(new_n760), .ZN(new_n761));
  INV_X1    g336(.A(new_n761), .ZN(new_n762));
  OAI21_X1  g337(.A(new_n756), .B1(new_n762), .B2(new_n727), .ZN(new_n763));
  XNOR2_X1  g338(.A(new_n763), .B(G2067), .ZN(new_n764));
  INV_X1    g339(.A(G1961), .ZN(new_n765));
  AND2_X1   g340(.A1(new_n721), .A2(G5), .ZN(new_n766));
  AOI21_X1  g341(.A(new_n766), .B1(G301), .B2(G16), .ZN(new_n767));
  AOI21_X1  g342(.A(new_n764), .B1(new_n765), .B2(new_n767), .ZN(new_n768));
  NOR2_X1   g343(.A1(new_n753), .A2(G1341), .ZN(new_n769));
  NOR2_X1   g344(.A1(new_n767), .A2(new_n765), .ZN(new_n770));
  NOR2_X1   g345(.A1(new_n769), .A2(new_n770), .ZN(new_n771));
  XNOR2_X1  g346(.A(KEYINPUT27), .B(G1996), .ZN(new_n772));
  NAND2_X1  g347(.A1(new_n480), .A2(G129), .ZN(new_n773));
  NAND2_X1  g348(.A1(new_n476), .A2(G141), .ZN(new_n774));
  NAND3_X1  g349(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n775));
  XOR2_X1   g350(.A(new_n775), .B(KEYINPUT26), .Z(new_n776));
  NAND3_X1  g351(.A1(new_n460), .A2(G105), .A3(G2104), .ZN(new_n777));
  NAND4_X1  g352(.A1(new_n773), .A2(new_n774), .A3(new_n776), .A4(new_n777), .ZN(new_n778));
  NAND2_X1  g353(.A1(new_n778), .A2(G29), .ZN(new_n779));
  NAND2_X1  g354(.A1(new_n727), .A2(G32), .ZN(new_n780));
  AOI21_X1  g355(.A(new_n772), .B1(new_n779), .B2(new_n780), .ZN(new_n781));
  AND3_X1   g356(.A1(new_n779), .A2(new_n780), .A3(new_n772), .ZN(new_n782));
  AOI211_X1 g357(.A(new_n781), .B(new_n782), .C1(G2072), .C2(new_n750), .ZN(new_n783));
  NAND4_X1  g358(.A1(new_n754), .A2(new_n768), .A3(new_n771), .A4(new_n783), .ZN(new_n784));
  NOR2_X1   g359(.A1(new_n731), .A2(G2090), .ZN(new_n785));
  NOR3_X1   g360(.A1(new_n732), .A2(new_n784), .A3(new_n785), .ZN(new_n786));
  NAND2_X1  g361(.A1(new_n721), .A2(G21), .ZN(new_n787));
  OAI21_X1  g362(.A(new_n787), .B1(G168), .B2(new_n721), .ZN(new_n788));
  XNOR2_X1  g363(.A(KEYINPUT97), .B(G1966), .ZN(new_n789));
  XNOR2_X1  g364(.A(new_n788), .B(new_n789), .ZN(new_n790));
  NAND2_X1  g365(.A1(new_n727), .A2(G27), .ZN(new_n791));
  XNOR2_X1  g366(.A(new_n791), .B(KEYINPUT99), .ZN(new_n792));
  OAI21_X1  g367(.A(new_n792), .B1(G164), .B2(new_n727), .ZN(new_n793));
  INV_X1    g368(.A(new_n793), .ZN(new_n794));
  XNOR2_X1  g369(.A(KEYINPUT100), .B(G2078), .ZN(new_n795));
  AOI21_X1  g370(.A(new_n790), .B1(new_n794), .B2(new_n795), .ZN(new_n796));
  NOR2_X1   g371(.A1(G4), .A2(G16), .ZN(new_n797));
  XNOR2_X1  g372(.A(new_n797), .B(KEYINPUT95), .ZN(new_n798));
  INV_X1    g373(.A(new_n633), .ZN(new_n799));
  OAI21_X1  g374(.A(new_n798), .B1(new_n799), .B2(new_n721), .ZN(new_n800));
  XOR2_X1   g375(.A(KEYINPUT96), .B(G1348), .Z(new_n801));
  OR2_X1    g376(.A1(new_n800), .A2(new_n801), .ZN(new_n802));
  INV_X1    g377(.A(KEYINPUT24), .ZN(new_n803));
  INV_X1    g378(.A(G34), .ZN(new_n804));
  AOI21_X1  g379(.A(G29), .B1(new_n803), .B2(new_n804), .ZN(new_n805));
  OAI21_X1  g380(.A(new_n805), .B1(new_n803), .B2(new_n804), .ZN(new_n806));
  OAI21_X1  g381(.A(new_n806), .B1(G160), .B2(new_n727), .ZN(new_n807));
  INV_X1    g382(.A(new_n795), .ZN(new_n808));
  AOI22_X1  g383(.A1(new_n807), .A2(G2084), .B1(new_n793), .B2(new_n808), .ZN(new_n809));
  AND3_X1   g384(.A1(new_n796), .A2(new_n802), .A3(new_n809), .ZN(new_n810));
  OR2_X1    g385(.A1(new_n807), .A2(G2084), .ZN(new_n811));
  XNOR2_X1  g386(.A(new_n811), .B(KEYINPUT98), .ZN(new_n812));
  AOI21_X1  g387(.A(new_n812), .B1(new_n801), .B2(new_n800), .ZN(new_n813));
  AND4_X1   g388(.A1(new_n726), .A2(new_n786), .A3(new_n810), .A4(new_n813), .ZN(new_n814));
  MUX2_X1   g389(.A(G23), .B(G288), .S(G16), .Z(new_n815));
  OR2_X1    g390(.A1(new_n815), .A2(KEYINPUT33), .ZN(new_n816));
  NAND2_X1  g391(.A1(new_n815), .A2(KEYINPUT33), .ZN(new_n817));
  NAND2_X1  g392(.A1(new_n816), .A2(new_n817), .ZN(new_n818));
  INV_X1    g393(.A(G1976), .ZN(new_n819));
  NAND2_X1  g394(.A1(new_n818), .A2(new_n819), .ZN(new_n820));
  NAND3_X1  g395(.A1(new_n816), .A2(G1976), .A3(new_n817), .ZN(new_n821));
  MUX2_X1   g396(.A(G6), .B(G305), .S(G16), .Z(new_n822));
  XOR2_X1   g397(.A(KEYINPUT32), .B(G1981), .Z(new_n823));
  XNOR2_X1  g398(.A(new_n822), .B(new_n823), .ZN(new_n824));
  NAND2_X1  g399(.A1(new_n721), .A2(G22), .ZN(new_n825));
  OAI21_X1  g400(.A(new_n825), .B1(G166), .B2(new_n721), .ZN(new_n826));
  INV_X1    g401(.A(G1971), .ZN(new_n827));
  XNOR2_X1  g402(.A(new_n826), .B(new_n827), .ZN(new_n828));
  NAND4_X1  g403(.A1(new_n820), .A2(new_n821), .A3(new_n824), .A4(new_n828), .ZN(new_n829));
  OR2_X1    g404(.A1(new_n829), .A2(KEYINPUT34), .ZN(new_n830));
  NAND2_X1  g405(.A1(new_n829), .A2(KEYINPUT34), .ZN(new_n831));
  NAND2_X1  g406(.A1(new_n727), .A2(G25), .ZN(new_n832));
  XOR2_X1   g407(.A(new_n832), .B(KEYINPUT90), .Z(new_n833));
  NAND2_X1  g408(.A1(new_n480), .A2(G119), .ZN(new_n834));
  INV_X1    g409(.A(G95), .ZN(new_n835));
  AND3_X1   g410(.A1(new_n835), .A2(new_n460), .A3(KEYINPUT91), .ZN(new_n836));
  AOI21_X1  g411(.A(KEYINPUT91), .B1(new_n835), .B2(new_n460), .ZN(new_n837));
  OAI221_X1 g412(.A(G2104), .B1(G107), .B2(new_n460), .C1(new_n836), .C2(new_n837), .ZN(new_n838));
  NAND2_X1  g413(.A1(new_n476), .A2(G131), .ZN(new_n839));
  NAND3_X1  g414(.A1(new_n834), .A2(new_n838), .A3(new_n839), .ZN(new_n840));
  NAND2_X1  g415(.A1(new_n840), .A2(KEYINPUT92), .ZN(new_n841));
  INV_X1    g416(.A(KEYINPUT92), .ZN(new_n842));
  NAND4_X1  g417(.A1(new_n834), .A2(new_n838), .A3(new_n839), .A4(new_n842), .ZN(new_n843));
  NAND2_X1  g418(.A1(new_n841), .A2(new_n843), .ZN(new_n844));
  AOI21_X1  g419(.A(new_n833), .B1(new_n844), .B2(G29), .ZN(new_n845));
  XOR2_X1   g420(.A(KEYINPUT35), .B(G1991), .Z(new_n846));
  XNOR2_X1  g421(.A(new_n845), .B(new_n846), .ZN(new_n847));
  MUX2_X1   g422(.A(G24), .B(G290), .S(G16), .Z(new_n848));
  XNOR2_X1  g423(.A(new_n848), .B(G1986), .ZN(new_n849));
  AOI211_X1 g424(.A(new_n847), .B(new_n849), .C1(KEYINPUT94), .C2(KEYINPUT36), .ZN(new_n850));
  NAND3_X1  g425(.A1(new_n830), .A2(new_n831), .A3(new_n850), .ZN(new_n851));
  INV_X1    g426(.A(KEYINPUT94), .ZN(new_n852));
  INV_X1    g427(.A(KEYINPUT36), .ZN(new_n853));
  OAI21_X1  g428(.A(new_n852), .B1(new_n853), .B2(KEYINPUT93), .ZN(new_n854));
  INV_X1    g429(.A(new_n854), .ZN(new_n855));
  NAND2_X1  g430(.A1(new_n851), .A2(new_n855), .ZN(new_n856));
  NAND4_X1  g431(.A1(new_n830), .A2(new_n854), .A3(new_n831), .A4(new_n850), .ZN(new_n857));
  NAND3_X1  g432(.A1(new_n814), .A2(new_n856), .A3(new_n857), .ZN(G150));
  INV_X1    g433(.A(KEYINPUT102), .ZN(new_n859));
  XNOR2_X1  g434(.A(G150), .B(new_n859), .ZN(G311));
  NAND2_X1  g435(.A1(new_n633), .A2(G559), .ZN(new_n861));
  NAND2_X1  g436(.A1(new_n528), .A2(G55), .ZN(new_n862));
  NAND2_X1  g437(.A1(G80), .A2(G543), .ZN(new_n863));
  INV_X1    g438(.A(G67), .ZN(new_n864));
  OAI21_X1  g439(.A(new_n863), .B1(new_n545), .B2(new_n864), .ZN(new_n865));
  AOI22_X1  g440(.A1(new_n534), .A2(G93), .B1(new_n865), .B2(G651), .ZN(new_n866));
  NAND2_X1  g441(.A1(new_n862), .A2(new_n866), .ZN(new_n867));
  NAND2_X1  g442(.A1(new_n867), .A2(new_n556), .ZN(new_n868));
  NAND4_X1  g443(.A1(new_n551), .A2(new_n862), .A3(new_n555), .A4(new_n866), .ZN(new_n869));
  NAND2_X1  g444(.A1(new_n868), .A2(new_n869), .ZN(new_n870));
  XNOR2_X1  g445(.A(new_n861), .B(new_n870), .ZN(new_n871));
  XOR2_X1   g446(.A(KEYINPUT103), .B(KEYINPUT38), .Z(new_n872));
  XNOR2_X1  g447(.A(new_n871), .B(new_n872), .ZN(new_n873));
  INV_X1    g448(.A(KEYINPUT39), .ZN(new_n874));
  AOI21_X1  g449(.A(G860), .B1(new_n873), .B2(new_n874), .ZN(new_n875));
  OAI21_X1  g450(.A(new_n875), .B1(new_n874), .B2(new_n873), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n867), .A2(G860), .ZN(new_n877));
  XOR2_X1   g452(.A(new_n877), .B(KEYINPUT37), .Z(new_n878));
  NAND2_X1  g453(.A1(new_n876), .A2(new_n878), .ZN(G145));
  NAND2_X1  g454(.A1(new_n480), .A2(G130), .ZN(new_n880));
  NAND2_X1  g455(.A1(new_n476), .A2(G142), .ZN(new_n881));
  OR2_X1    g456(.A1(G106), .A2(G2105), .ZN(new_n882));
  OAI211_X1 g457(.A(new_n882), .B(G2104), .C1(G118), .C2(new_n460), .ZN(new_n883));
  NAND3_X1  g458(.A1(new_n880), .A2(new_n881), .A3(new_n883), .ZN(new_n884));
  OR2_X1    g459(.A1(new_n884), .A2(new_n649), .ZN(new_n885));
  NAND2_X1  g460(.A1(new_n884), .A2(new_n649), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n885), .A2(new_n886), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n887), .A2(new_n844), .ZN(new_n888));
  NAND4_X1  g463(.A1(new_n885), .A2(new_n841), .A3(new_n843), .A4(new_n886), .ZN(new_n889));
  NAND2_X1  g464(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  INV_X1    g465(.A(KEYINPUT104), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n890), .A2(new_n891), .ZN(new_n892));
  NAND3_X1  g467(.A1(new_n888), .A2(KEYINPUT104), .A3(new_n889), .ZN(new_n893));
  NAND2_X1  g468(.A1(new_n892), .A2(new_n893), .ZN(new_n894));
  INV_X1    g469(.A(new_n894), .ZN(new_n895));
  NAND4_X1  g470(.A1(new_n490), .A2(new_n497), .A3(new_n503), .A4(new_n502), .ZN(new_n896));
  XOR2_X1   g471(.A(new_n761), .B(new_n896), .Z(new_n897));
  INV_X1    g472(.A(new_n778), .ZN(new_n898));
  NAND2_X1  g473(.A1(new_n897), .A2(new_n898), .ZN(new_n899));
  XNOR2_X1  g474(.A(new_n761), .B(new_n896), .ZN(new_n900));
  NAND2_X1  g475(.A1(new_n900), .A2(new_n778), .ZN(new_n901));
  NAND2_X1  g476(.A1(new_n899), .A2(new_n901), .ZN(new_n902));
  INV_X1    g477(.A(new_n749), .ZN(new_n903));
  NAND2_X1  g478(.A1(new_n902), .A2(new_n903), .ZN(new_n904));
  NAND3_X1  g479(.A1(new_n899), .A2(new_n749), .A3(new_n901), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  OAI21_X1  g481(.A(KEYINPUT105), .B1(new_n895), .B2(new_n906), .ZN(new_n907));
  INV_X1    g482(.A(KEYINPUT105), .ZN(new_n908));
  NAND4_X1  g483(.A1(new_n894), .A2(new_n908), .A3(new_n905), .A4(new_n904), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n907), .A2(new_n909), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n895), .A2(new_n906), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n910), .A2(new_n911), .ZN(new_n912));
  XNOR2_X1  g487(.A(G160), .B(new_n659), .ZN(new_n913));
  XNOR2_X1  g488(.A(new_n913), .B(G162), .ZN(new_n914));
  AOI21_X1  g489(.A(G37), .B1(new_n912), .B2(new_n914), .ZN(new_n915));
  AOI21_X1  g490(.A(new_n890), .B1(new_n904), .B2(new_n905), .ZN(new_n916));
  INV_X1    g491(.A(KEYINPUT106), .ZN(new_n917));
  OR2_X1    g492(.A1(new_n916), .A2(new_n917), .ZN(new_n918));
  AOI21_X1  g493(.A(new_n914), .B1(new_n916), .B2(new_n917), .ZN(new_n919));
  AND2_X1   g494(.A1(new_n918), .A2(new_n919), .ZN(new_n920));
  AOI21_X1  g495(.A(KEYINPUT107), .B1(new_n920), .B2(new_n910), .ZN(new_n921));
  AND4_X1   g496(.A1(KEYINPUT107), .A2(new_n910), .A3(new_n918), .A4(new_n919), .ZN(new_n922));
  OAI21_X1  g497(.A(new_n915), .B1(new_n921), .B2(new_n922), .ZN(new_n923));
  XNOR2_X1  g498(.A(new_n923), .B(KEYINPUT40), .ZN(G395));
  XNOR2_X1  g499(.A(new_n644), .B(new_n870), .ZN(new_n925));
  NAND3_X1  g500(.A1(new_n581), .A2(new_n633), .A3(new_n587), .ZN(new_n926));
  INV_X1    g501(.A(new_n926), .ZN(new_n927));
  AOI21_X1  g502(.A(new_n633), .B1(new_n581), .B2(new_n587), .ZN(new_n928));
  OAI21_X1  g503(.A(new_n925), .B1(new_n927), .B2(new_n928), .ZN(new_n929));
  NAND2_X1  g504(.A1(G299), .A2(new_n799), .ZN(new_n930));
  INV_X1    g505(.A(KEYINPUT41), .ZN(new_n931));
  NAND3_X1  g506(.A1(new_n930), .A2(new_n931), .A3(new_n926), .ZN(new_n932));
  INV_X1    g507(.A(KEYINPUT108), .ZN(new_n933));
  NAND2_X1  g508(.A1(new_n932), .A2(new_n933), .ZN(new_n934));
  NAND4_X1  g509(.A1(new_n930), .A2(KEYINPUT108), .A3(new_n931), .A4(new_n926), .ZN(new_n935));
  OAI21_X1  g510(.A(KEYINPUT41), .B1(new_n927), .B2(new_n928), .ZN(new_n936));
  NAND3_X1  g511(.A1(new_n934), .A2(new_n935), .A3(new_n936), .ZN(new_n937));
  OAI21_X1  g512(.A(new_n929), .B1(new_n937), .B2(new_n925), .ZN(new_n938));
  OR2_X1    g513(.A1(new_n938), .A2(KEYINPUT42), .ZN(new_n939));
  XOR2_X1   g514(.A(G290), .B(G305), .Z(new_n940));
  XNOR2_X1  g515(.A(G288), .B(G166), .ZN(new_n941));
  XNOR2_X1  g516(.A(new_n940), .B(new_n941), .ZN(new_n942));
  INV_X1    g517(.A(new_n942), .ZN(new_n943));
  NAND2_X1  g518(.A1(new_n938), .A2(KEYINPUT42), .ZN(new_n944));
  AND3_X1   g519(.A1(new_n939), .A2(new_n943), .A3(new_n944), .ZN(new_n945));
  AOI21_X1  g520(.A(new_n943), .B1(new_n939), .B2(new_n944), .ZN(new_n946));
  OAI21_X1  g521(.A(G868), .B1(new_n945), .B2(new_n946), .ZN(new_n947));
  NAND2_X1  g522(.A1(new_n867), .A2(new_n636), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n947), .A2(new_n948), .ZN(G295));
  NAND2_X1  g524(.A1(new_n947), .A2(new_n948), .ZN(G331));
  NAND2_X1  g525(.A1(G286), .A2(G301), .ZN(new_n951));
  AND2_X1   g526(.A1(new_n539), .A2(new_n535), .ZN(new_n952));
  NAND4_X1  g527(.A1(new_n952), .A2(new_n529), .A3(new_n543), .A4(new_n548), .ZN(new_n953));
  NAND2_X1  g528(.A1(new_n951), .A2(new_n953), .ZN(new_n954));
  NAND2_X1  g529(.A1(new_n954), .A2(new_n870), .ZN(new_n955));
  NAND4_X1  g530(.A1(new_n951), .A2(new_n868), .A3(new_n953), .A4(new_n869), .ZN(new_n956));
  AND2_X1   g531(.A1(new_n955), .A2(new_n956), .ZN(new_n957));
  NOR3_X1   g532(.A1(new_n927), .A2(new_n928), .A3(KEYINPUT41), .ZN(new_n958));
  INV_X1    g533(.A(KEYINPUT110), .ZN(new_n959));
  AOI21_X1  g534(.A(new_n958), .B1(new_n959), .B2(new_n936), .ZN(new_n960));
  OR2_X1    g535(.A1(new_n936), .A2(new_n959), .ZN(new_n961));
  AOI21_X1  g536(.A(new_n957), .B1(new_n960), .B2(new_n961), .ZN(new_n962));
  INV_X1    g537(.A(KEYINPUT109), .ZN(new_n963));
  NAND3_X1  g538(.A1(new_n955), .A2(new_n963), .A3(new_n956), .ZN(new_n964));
  INV_X1    g539(.A(new_n870), .ZN(new_n965));
  NAND4_X1  g540(.A1(new_n965), .A2(KEYINPUT109), .A3(new_n951), .A4(new_n953), .ZN(new_n966));
  NAND2_X1  g541(.A1(new_n964), .A2(new_n966), .ZN(new_n967));
  NOR2_X1   g542(.A1(new_n927), .A2(new_n928), .ZN(new_n968));
  NAND2_X1  g543(.A1(new_n967), .A2(new_n968), .ZN(new_n969));
  INV_X1    g544(.A(KEYINPUT111), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n969), .A2(new_n970), .ZN(new_n971));
  NAND3_X1  g546(.A1(new_n967), .A2(KEYINPUT111), .A3(new_n968), .ZN(new_n972));
  NAND2_X1  g547(.A1(new_n971), .A2(new_n972), .ZN(new_n973));
  OAI21_X1  g548(.A(new_n943), .B1(new_n962), .B2(new_n973), .ZN(new_n974));
  AND2_X1   g549(.A1(new_n968), .A2(new_n957), .ZN(new_n975));
  INV_X1    g550(.A(new_n967), .ZN(new_n976));
  AOI21_X1  g551(.A(new_n975), .B1(new_n937), .B2(new_n976), .ZN(new_n977));
  AOI21_X1  g552(.A(G37), .B1(new_n977), .B2(new_n942), .ZN(new_n978));
  AND3_X1   g553(.A1(new_n974), .A2(new_n978), .A3(KEYINPUT43), .ZN(new_n979));
  OR2_X1    g554(.A1(new_n977), .A2(new_n942), .ZN(new_n980));
  AOI21_X1  g555(.A(KEYINPUT43), .B1(new_n980), .B2(new_n978), .ZN(new_n981));
  OAI21_X1  g556(.A(KEYINPUT44), .B1(new_n979), .B2(new_n981), .ZN(new_n982));
  INV_X1    g557(.A(KEYINPUT43), .ZN(new_n983));
  AND3_X1   g558(.A1(new_n974), .A2(new_n978), .A3(new_n983), .ZN(new_n984));
  AOI21_X1  g559(.A(new_n983), .B1(new_n980), .B2(new_n978), .ZN(new_n985));
  NOR2_X1   g560(.A1(new_n984), .A2(new_n985), .ZN(new_n986));
  OAI21_X1  g561(.A(new_n982), .B1(new_n986), .B2(KEYINPUT44), .ZN(G397));
  INV_X1    g562(.A(G2067), .ZN(new_n988));
  XNOR2_X1  g563(.A(new_n761), .B(new_n988), .ZN(new_n989));
  XNOR2_X1  g564(.A(new_n989), .B(KEYINPUT113), .ZN(new_n990));
  INV_X1    g565(.A(G1384), .ZN(new_n991));
  NAND2_X1  g566(.A1(new_n896), .A2(new_n991), .ZN(new_n992));
  INV_X1    g567(.A(KEYINPUT45), .ZN(new_n993));
  NAND2_X1  g568(.A1(new_n992), .A2(new_n993), .ZN(new_n994));
  INV_X1    g569(.A(G125), .ZN(new_n995));
  AOI21_X1  g570(.A(new_n995), .B1(new_n492), .B2(new_n493), .ZN(new_n996));
  OAI21_X1  g571(.A(new_n461), .B1(new_n996), .B2(new_n467), .ZN(new_n997));
  INV_X1    g572(.A(new_n468), .ZN(new_n998));
  OAI21_X1  g573(.A(G2105), .B1(new_n997), .B2(new_n998), .ZN(new_n999));
  INV_X1    g574(.A(KEYINPUT112), .ZN(new_n1000));
  INV_X1    g575(.A(G40), .ZN(new_n1001));
  AOI21_X1  g576(.A(new_n1001), .B1(new_n473), .B2(new_n460), .ZN(new_n1002));
  NAND3_X1  g577(.A1(new_n999), .A2(new_n1000), .A3(new_n1002), .ZN(new_n1003));
  AOI22_X1  g578(.A1(new_n494), .A2(G137), .B1(G101), .B2(G2104), .ZN(new_n1004));
  OAI21_X1  g579(.A(G40), .B1(new_n1004), .B2(G2105), .ZN(new_n1005));
  OAI21_X1  g580(.A(KEYINPUT112), .B1(new_n469), .B2(new_n1005), .ZN(new_n1006));
  AOI21_X1  g581(.A(new_n994), .B1(new_n1003), .B2(new_n1006), .ZN(new_n1007));
  NAND2_X1  g582(.A1(new_n990), .A2(new_n1007), .ZN(new_n1008));
  XOR2_X1   g583(.A(new_n1008), .B(KEYINPUT114), .Z(new_n1009));
  AOI21_X1  g584(.A(new_n846), .B1(new_n841), .B2(new_n843), .ZN(new_n1010));
  AND3_X1   g585(.A1(new_n841), .A2(new_n846), .A3(new_n843), .ZN(new_n1011));
  OAI21_X1  g586(.A(new_n1007), .B1(new_n1010), .B2(new_n1011), .ZN(new_n1012));
  XNOR2_X1  g587(.A(new_n778), .B(G1996), .ZN(new_n1013));
  NAND2_X1  g588(.A1(new_n1007), .A2(new_n1013), .ZN(new_n1014));
  AND3_X1   g589(.A1(new_n1009), .A2(new_n1012), .A3(new_n1014), .ZN(new_n1015));
  XNOR2_X1  g590(.A(G290), .B(G1986), .ZN(new_n1016));
  NAND2_X1  g591(.A1(new_n1016), .A2(new_n1007), .ZN(new_n1017));
  AND2_X1   g592(.A1(new_n1015), .A2(new_n1017), .ZN(new_n1018));
  AOI21_X1  g593(.A(new_n992), .B1(new_n1006), .B2(new_n1003), .ZN(new_n1019));
  INV_X1    g594(.A(G8), .ZN(new_n1020));
  NOR2_X1   g595(.A1(new_n1019), .A2(new_n1020), .ZN(new_n1021));
  AND2_X1   g596(.A1(new_n609), .A2(new_n610), .ZN(new_n1022));
  OAI21_X1  g597(.A(G61), .B1(new_n510), .B2(new_n511), .ZN(new_n1023));
  AOI21_X1  g598(.A(new_n509), .B1(new_n1022), .B2(new_n1023), .ZN(new_n1024));
  AOI21_X1  g599(.A(new_n518), .B1(new_n601), .B2(new_n602), .ZN(new_n1025));
  OAI21_X1  g600(.A(G1981), .B1(new_n1024), .B2(new_n1025), .ZN(new_n1026));
  INV_X1    g601(.A(G1981), .ZN(new_n1027));
  NAND3_X1  g602(.A1(new_n604), .A2(new_n612), .A3(new_n1027), .ZN(new_n1028));
  AND3_X1   g603(.A1(new_n1026), .A2(KEYINPUT49), .A3(new_n1028), .ZN(new_n1029));
  AOI21_X1  g604(.A(KEYINPUT49), .B1(new_n1026), .B2(new_n1028), .ZN(new_n1030));
  NOR2_X1   g605(.A1(new_n1029), .A2(new_n1030), .ZN(new_n1031));
  AOI211_X1 g606(.A(G1976), .B(G288), .C1(new_n1021), .C2(new_n1031), .ZN(new_n1032));
  XNOR2_X1  g607(.A(new_n1028), .B(KEYINPUT117), .ZN(new_n1033));
  OAI21_X1  g608(.A(new_n1021), .B1(new_n1032), .B2(new_n1033), .ZN(new_n1034));
  NAND2_X1  g609(.A1(new_n1006), .A2(new_n1003), .ZN(new_n1035));
  AND2_X1   g610(.A1(new_n896), .A2(new_n991), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n1035), .A2(new_n1036), .ZN(new_n1037));
  OAI21_X1  g612(.A(KEYINPUT116), .B1(G288), .B2(new_n819), .ZN(new_n1038));
  INV_X1    g613(.A(KEYINPUT116), .ZN(new_n1039));
  NAND4_X1  g614(.A1(new_n598), .A2(new_n1039), .A3(G1976), .A4(new_n599), .ZN(new_n1040));
  NAND2_X1  g615(.A1(new_n1038), .A2(new_n1040), .ZN(new_n1041));
  AOI21_X1  g616(.A(KEYINPUT52), .B1(G288), .B2(new_n819), .ZN(new_n1042));
  NAND4_X1  g617(.A1(new_n1037), .A2(new_n1041), .A3(G8), .A4(new_n1042), .ZN(new_n1043));
  NAND3_X1  g618(.A1(new_n1037), .A2(new_n1031), .A3(G8), .ZN(new_n1044));
  NAND2_X1  g619(.A1(new_n1043), .A2(new_n1044), .ZN(new_n1045));
  INV_X1    g620(.A(KEYINPUT52), .ZN(new_n1046));
  AOI21_X1  g621(.A(new_n1046), .B1(new_n1021), .B2(new_n1041), .ZN(new_n1047));
  NOR2_X1   g622(.A1(new_n1045), .A2(new_n1047), .ZN(new_n1048));
  INV_X1    g623(.A(new_n1048), .ZN(new_n1049));
  OAI21_X1  g624(.A(new_n993), .B1(G164), .B2(G1384), .ZN(new_n1050));
  NAND2_X1  g625(.A1(new_n1036), .A2(KEYINPUT45), .ZN(new_n1051));
  NAND3_X1  g626(.A1(new_n1050), .A2(new_n1035), .A3(new_n1051), .ZN(new_n1052));
  NAND2_X1  g627(.A1(new_n1052), .A2(new_n827), .ZN(new_n1053));
  OAI21_X1  g628(.A(KEYINPUT50), .B1(G164), .B2(G1384), .ZN(new_n1054));
  INV_X1    g629(.A(KEYINPUT50), .ZN(new_n1055));
  NAND2_X1  g630(.A1(new_n1036), .A2(new_n1055), .ZN(new_n1056));
  INV_X1    g631(.A(G2090), .ZN(new_n1057));
  NAND4_X1  g632(.A1(new_n1054), .A2(new_n1035), .A3(new_n1056), .A4(new_n1057), .ZN(new_n1058));
  NAND2_X1  g633(.A1(new_n1053), .A2(new_n1058), .ZN(new_n1059));
  NAND3_X1  g634(.A1(new_n593), .A2(new_n594), .A3(G8), .ZN(new_n1060));
  NAND2_X1  g635(.A1(new_n1060), .A2(KEYINPUT55), .ZN(new_n1061));
  INV_X1    g636(.A(KEYINPUT55), .ZN(new_n1062));
  NAND4_X1  g637(.A1(new_n593), .A2(new_n594), .A3(new_n1062), .A4(G8), .ZN(new_n1063));
  NAND2_X1  g638(.A1(new_n1061), .A2(new_n1063), .ZN(new_n1064));
  NAND2_X1  g639(.A1(new_n1064), .A2(KEYINPUT115), .ZN(new_n1065));
  INV_X1    g640(.A(KEYINPUT115), .ZN(new_n1066));
  NAND3_X1  g641(.A1(new_n1061), .A2(new_n1066), .A3(new_n1063), .ZN(new_n1067));
  NAND2_X1  g642(.A1(new_n1065), .A2(new_n1067), .ZN(new_n1068));
  NAND3_X1  g643(.A1(new_n1059), .A2(G8), .A3(new_n1068), .ZN(new_n1069));
  OAI21_X1  g644(.A(new_n1034), .B1(new_n1049), .B2(new_n1069), .ZN(new_n1070));
  INV_X1    g645(.A(KEYINPUT63), .ZN(new_n1071));
  INV_X1    g646(.A(new_n1064), .ZN(new_n1072));
  AOI22_X1  g647(.A1(new_n1006), .A2(new_n1003), .B1(KEYINPUT50), .B2(new_n992), .ZN(new_n1073));
  INV_X1    g648(.A(KEYINPUT118), .ZN(new_n1074));
  NAND2_X1  g649(.A1(new_n505), .A2(new_n507), .ZN(new_n1075));
  INV_X1    g650(.A(new_n498), .ZN(new_n1076));
  AOI21_X1  g651(.A(G1384), .B1(new_n1075), .B2(new_n1076), .ZN(new_n1077));
  AOI21_X1  g652(.A(new_n1074), .B1(new_n1077), .B2(new_n1055), .ZN(new_n1078));
  AND3_X1   g653(.A1(new_n502), .A2(new_n506), .A3(new_n503), .ZN(new_n1079));
  AOI21_X1  g654(.A(new_n506), .B1(new_n502), .B2(new_n503), .ZN(new_n1080));
  OAI211_X1 g655(.A(new_n490), .B(new_n497), .C1(new_n1079), .C2(new_n1080), .ZN(new_n1081));
  AND4_X1   g656(.A1(new_n1074), .A2(new_n1081), .A3(new_n1055), .A4(new_n991), .ZN(new_n1082));
  OAI211_X1 g657(.A(new_n1057), .B(new_n1073), .C1(new_n1078), .C2(new_n1082), .ZN(new_n1083));
  AOI21_X1  g658(.A(new_n1020), .B1(new_n1083), .B2(new_n1053), .ZN(new_n1084));
  OAI211_X1 g659(.A(new_n1048), .B(new_n1069), .C1(new_n1072), .C2(new_n1084), .ZN(new_n1085));
  NAND3_X1  g660(.A1(new_n1081), .A2(KEYINPUT45), .A3(new_n991), .ZN(new_n1086));
  NAND3_X1  g661(.A1(new_n1035), .A2(new_n1086), .A3(new_n994), .ZN(new_n1087));
  INV_X1    g662(.A(G1966), .ZN(new_n1088));
  NAND2_X1  g663(.A1(new_n1087), .A2(new_n1088), .ZN(new_n1089));
  INV_X1    g664(.A(G2084), .ZN(new_n1090));
  NAND4_X1  g665(.A1(new_n1054), .A2(new_n1035), .A3(new_n1056), .A4(new_n1090), .ZN(new_n1091));
  NAND2_X1  g666(.A1(new_n1089), .A2(new_n1091), .ZN(new_n1092));
  NAND3_X1  g667(.A1(new_n1092), .A2(G8), .A3(G168), .ZN(new_n1093));
  OAI21_X1  g668(.A(new_n1071), .B1(new_n1085), .B2(new_n1093), .ZN(new_n1094));
  NOR2_X1   g669(.A1(new_n1093), .A2(new_n1071), .ZN(new_n1095));
  NAND2_X1  g670(.A1(new_n1059), .A2(G8), .ZN(new_n1096));
  NAND2_X1  g671(.A1(new_n1096), .A2(new_n1064), .ZN(new_n1097));
  NAND4_X1  g672(.A1(new_n1095), .A2(new_n1069), .A3(new_n1097), .A4(new_n1048), .ZN(new_n1098));
  AOI21_X1  g673(.A(new_n1070), .B1(new_n1094), .B2(new_n1098), .ZN(new_n1099));
  NAND3_X1  g674(.A1(new_n1089), .A2(G168), .A3(new_n1091), .ZN(new_n1100));
  NAND2_X1  g675(.A1(new_n1100), .A2(G8), .ZN(new_n1101));
  NAND2_X1  g676(.A1(new_n1101), .A2(KEYINPUT51), .ZN(new_n1102));
  AOI21_X1  g677(.A(G168), .B1(new_n1089), .B2(new_n1091), .ZN(new_n1103));
  INV_X1    g678(.A(KEYINPUT51), .ZN(new_n1104));
  OAI211_X1 g679(.A(G8), .B(new_n1100), .C1(new_n1103), .C2(new_n1104), .ZN(new_n1105));
  INV_X1    g680(.A(KEYINPUT62), .ZN(new_n1106));
  AND3_X1   g681(.A1(new_n1102), .A2(new_n1105), .A3(new_n1106), .ZN(new_n1107));
  NAND2_X1  g682(.A1(new_n1083), .A2(new_n1053), .ZN(new_n1108));
  NAND2_X1  g683(.A1(new_n1108), .A2(G8), .ZN(new_n1109));
  NAND2_X1  g684(.A1(new_n1109), .A2(new_n1064), .ZN(new_n1110));
  INV_X1    g685(.A(G2078), .ZN(new_n1111));
  NAND4_X1  g686(.A1(new_n1050), .A2(new_n1035), .A3(new_n1051), .A4(new_n1111), .ZN(new_n1112));
  INV_X1    g687(.A(KEYINPUT53), .ZN(new_n1113));
  NAND3_X1  g688(.A1(new_n1054), .A2(new_n1035), .A3(new_n1056), .ZN(new_n1114));
  AOI22_X1  g689(.A1(new_n1112), .A2(new_n1113), .B1(new_n1114), .B2(new_n765), .ZN(new_n1115));
  NOR2_X1   g690(.A1(new_n1113), .A2(G2078), .ZN(new_n1116));
  INV_X1    g691(.A(new_n1116), .ZN(new_n1117));
  OR2_X1    g692(.A1(new_n1087), .A2(new_n1117), .ZN(new_n1118));
  AOI21_X1  g693(.A(G301), .B1(new_n1115), .B2(new_n1118), .ZN(new_n1119));
  NAND4_X1  g694(.A1(new_n1110), .A2(new_n1119), .A3(new_n1069), .A4(new_n1048), .ZN(new_n1120));
  NOR2_X1   g695(.A1(new_n1107), .A2(new_n1120), .ZN(new_n1121));
  AOI21_X1  g696(.A(new_n1104), .B1(new_n1092), .B2(G286), .ZN(new_n1122));
  NOR2_X1   g697(.A1(new_n1122), .A2(new_n1101), .ZN(new_n1123));
  AOI21_X1  g698(.A(new_n1104), .B1(new_n1100), .B2(G8), .ZN(new_n1124));
  OAI21_X1  g699(.A(KEYINPUT62), .B1(new_n1123), .B2(new_n1124), .ZN(new_n1125));
  AOI21_X1  g700(.A(KEYINPUT125), .B1(new_n1121), .B2(new_n1125), .ZN(new_n1126));
  INV_X1    g701(.A(new_n1119), .ZN(new_n1127));
  NOR2_X1   g702(.A1(new_n1085), .A2(new_n1127), .ZN(new_n1128));
  NAND3_X1  g703(.A1(new_n1102), .A2(new_n1105), .A3(new_n1106), .ZN(new_n1129));
  AND4_X1   g704(.A1(KEYINPUT125), .A2(new_n1128), .A3(new_n1125), .A4(new_n1129), .ZN(new_n1130));
  OAI21_X1  g705(.A(new_n1099), .B1(new_n1126), .B2(new_n1130), .ZN(new_n1131));
  NAND2_X1  g706(.A1(new_n1112), .A2(new_n1113), .ZN(new_n1132));
  NAND2_X1  g707(.A1(new_n1114), .A2(new_n765), .ZN(new_n1133));
  NOR3_X1   g708(.A1(new_n469), .A2(new_n1005), .A3(new_n1117), .ZN(new_n1134));
  NAND3_X1  g709(.A1(new_n1051), .A2(new_n994), .A3(new_n1134), .ZN(new_n1135));
  NAND3_X1  g710(.A1(new_n1132), .A2(new_n1133), .A3(new_n1135), .ZN(new_n1136));
  NAND2_X1  g711(.A1(new_n1136), .A2(G171), .ZN(new_n1137));
  NAND3_X1  g712(.A1(new_n1115), .A2(G301), .A3(new_n1118), .ZN(new_n1138));
  NAND3_X1  g713(.A1(new_n1137), .A2(KEYINPUT54), .A3(new_n1138), .ZN(new_n1139));
  NAND2_X1  g714(.A1(new_n1139), .A2(KEYINPUT124), .ZN(new_n1140));
  INV_X1    g715(.A(KEYINPUT124), .ZN(new_n1141));
  NAND4_X1  g716(.A1(new_n1137), .A2(new_n1138), .A3(new_n1141), .A4(KEYINPUT54), .ZN(new_n1142));
  NAND2_X1  g717(.A1(new_n1140), .A2(new_n1142), .ZN(new_n1143));
  AOI21_X1  g718(.A(new_n1085), .B1(new_n1102), .B2(new_n1105), .ZN(new_n1144));
  INV_X1    g719(.A(KEYINPUT54), .ZN(new_n1145));
  NOR2_X1   g720(.A1(new_n1136), .A2(G171), .ZN(new_n1146));
  OAI21_X1  g721(.A(new_n1145), .B1(new_n1146), .B2(new_n1119), .ZN(new_n1147));
  NAND3_X1  g722(.A1(new_n1143), .A2(new_n1144), .A3(new_n1147), .ZN(new_n1148));
  INV_X1    g723(.A(KEYINPUT123), .ZN(new_n1149));
  OAI21_X1  g724(.A(KEYINPUT119), .B1(new_n573), .B2(new_n580), .ZN(new_n1150));
  INV_X1    g725(.A(KEYINPUT119), .ZN(new_n1151));
  NAND4_X1  g726(.A1(new_n582), .A2(new_n584), .A3(new_n585), .A4(new_n1151), .ZN(new_n1152));
  NAND3_X1  g727(.A1(new_n1150), .A2(KEYINPUT57), .A3(new_n1152), .ZN(new_n1153));
  INV_X1    g728(.A(new_n1153), .ZN(new_n1154));
  AOI21_X1  g729(.A(KEYINPUT57), .B1(new_n1150), .B2(new_n1152), .ZN(new_n1155));
  NOR2_X1   g730(.A1(new_n1154), .A2(new_n1155), .ZN(new_n1156));
  OAI21_X1  g731(.A(new_n1073), .B1(new_n1078), .B2(new_n1082), .ZN(new_n1157));
  NAND2_X1  g732(.A1(new_n1157), .A2(new_n725), .ZN(new_n1158));
  INV_X1    g733(.A(new_n1052), .ZN(new_n1159));
  XNOR2_X1  g734(.A(KEYINPUT56), .B(G2072), .ZN(new_n1160));
  NAND2_X1  g735(.A1(new_n1159), .A2(new_n1160), .ZN(new_n1161));
  AND3_X1   g736(.A1(new_n1156), .A2(new_n1158), .A3(new_n1161), .ZN(new_n1162));
  AOI21_X1  g737(.A(new_n1156), .B1(new_n1158), .B2(new_n1161), .ZN(new_n1163));
  OAI21_X1  g738(.A(new_n1149), .B1(new_n1162), .B2(new_n1163), .ZN(new_n1164));
  NAND2_X1  g739(.A1(new_n1164), .A2(KEYINPUT61), .ZN(new_n1165));
  XNOR2_X1  g740(.A(KEYINPUT121), .B(KEYINPUT58), .ZN(new_n1166));
  XNOR2_X1  g741(.A(new_n1166), .B(G1341), .ZN(new_n1167));
  NAND2_X1  g742(.A1(new_n1037), .A2(new_n1167), .ZN(new_n1168));
  INV_X1    g743(.A(KEYINPUT122), .ZN(new_n1169));
  INV_X1    g744(.A(G1996), .ZN(new_n1170));
  NAND4_X1  g745(.A1(new_n1050), .A2(new_n1035), .A3(new_n1051), .A4(new_n1170), .ZN(new_n1171));
  AND3_X1   g746(.A1(new_n1168), .A2(new_n1169), .A3(new_n1171), .ZN(new_n1172));
  AOI21_X1  g747(.A(new_n1169), .B1(new_n1168), .B2(new_n1171), .ZN(new_n1173));
  OAI21_X1  g748(.A(new_n557), .B1(new_n1172), .B2(new_n1173), .ZN(new_n1174));
  NAND2_X1  g749(.A1(new_n1174), .A2(KEYINPUT59), .ZN(new_n1175));
  INV_X1    g750(.A(KEYINPUT59), .ZN(new_n1176));
  OAI211_X1 g751(.A(new_n1176), .B(new_n557), .C1(new_n1172), .C2(new_n1173), .ZN(new_n1177));
  INV_X1    g752(.A(G1348), .ZN(new_n1178));
  NAND2_X1  g753(.A1(new_n1114), .A2(new_n1178), .ZN(new_n1179));
  NAND2_X1  g754(.A1(new_n1019), .A2(new_n988), .ZN(new_n1180));
  NAND3_X1  g755(.A1(new_n1179), .A2(new_n1180), .A3(KEYINPUT60), .ZN(new_n1181));
  XNOR2_X1  g756(.A(new_n1181), .B(new_n633), .ZN(new_n1182));
  AND2_X1   g757(.A1(new_n1179), .A2(new_n1180), .ZN(new_n1183));
  OR2_X1    g758(.A1(new_n1183), .A2(KEYINPUT60), .ZN(new_n1184));
  AOI22_X1  g759(.A1(new_n1175), .A2(new_n1177), .B1(new_n1182), .B2(new_n1184), .ZN(new_n1185));
  INV_X1    g760(.A(KEYINPUT61), .ZN(new_n1186));
  OAI211_X1 g761(.A(new_n1149), .B(new_n1186), .C1(new_n1162), .C2(new_n1163), .ZN(new_n1187));
  NAND3_X1  g762(.A1(new_n1165), .A2(new_n1185), .A3(new_n1187), .ZN(new_n1188));
  AOI21_X1  g763(.A(new_n799), .B1(new_n1179), .B2(new_n1180), .ZN(new_n1189));
  INV_X1    g764(.A(KEYINPUT120), .ZN(new_n1190));
  AND2_X1   g765(.A1(new_n1189), .A2(new_n1190), .ZN(new_n1191));
  NOR2_X1   g766(.A1(new_n1189), .A2(new_n1190), .ZN(new_n1192));
  NOR3_X1   g767(.A1(new_n1163), .A2(new_n1191), .A3(new_n1192), .ZN(new_n1193));
  OR2_X1    g768(.A1(new_n1193), .A2(new_n1162), .ZN(new_n1194));
  AOI21_X1  g769(.A(new_n1148), .B1(new_n1188), .B2(new_n1194), .ZN(new_n1195));
  OAI21_X1  g770(.A(new_n1018), .B1(new_n1131), .B2(new_n1195), .ZN(new_n1196));
  INV_X1    g771(.A(new_n1007), .ZN(new_n1197));
  NAND3_X1  g772(.A1(new_n1009), .A2(new_n1011), .A3(new_n1014), .ZN(new_n1198));
  NAND2_X1  g773(.A1(new_n762), .A2(new_n988), .ZN(new_n1199));
  AOI21_X1  g774(.A(new_n1197), .B1(new_n1198), .B2(new_n1199), .ZN(new_n1200));
  OR2_X1    g775(.A1(new_n990), .A2(new_n778), .ZN(new_n1201));
  INV_X1    g776(.A(KEYINPUT46), .ZN(new_n1202));
  NAND2_X1  g777(.A1(new_n1007), .A2(new_n1170), .ZN(new_n1203));
  AOI22_X1  g778(.A1(new_n1201), .A2(new_n1007), .B1(new_n1202), .B2(new_n1203), .ZN(new_n1204));
  OAI21_X1  g779(.A(new_n1204), .B1(new_n1202), .B2(new_n1203), .ZN(new_n1205));
  XNOR2_X1  g780(.A(KEYINPUT126), .B(KEYINPUT47), .ZN(new_n1206));
  XNOR2_X1  g781(.A(new_n1205), .B(new_n1206), .ZN(new_n1207));
  NOR3_X1   g782(.A1(new_n1197), .A2(G1986), .A3(G290), .ZN(new_n1208));
  XOR2_X1   g783(.A(new_n1208), .B(KEYINPUT48), .Z(new_n1209));
  AOI211_X1 g784(.A(new_n1200), .B(new_n1207), .C1(new_n1015), .C2(new_n1209), .ZN(new_n1210));
  NAND2_X1  g785(.A1(new_n1196), .A2(new_n1210), .ZN(G329));
  assign    G231 = 1'b0;
  AND2_X1   g786(.A1(new_n680), .A2(G319), .ZN(new_n1213));
  AND4_X1   g787(.A1(new_n696), .A2(new_n718), .A3(new_n719), .A4(new_n1213), .ZN(new_n1214));
  OAI211_X1 g788(.A(new_n923), .B(new_n1214), .C1(new_n984), .C2(new_n985), .ZN(G225));
  INV_X1    g789(.A(G225), .ZN(G308));
endmodule


