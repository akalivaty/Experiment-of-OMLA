

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300,
         n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311,
         n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322,
         n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333,
         n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344,
         n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355,
         n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
         n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
         n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
         n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
         n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410,
         n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421,
         n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432,
         n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443,
         n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454,
         n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465,
         n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
         n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487,
         n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
         n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
         n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581;

  NOR2_X2 U322 ( .A1(n535), .A2(n496), .ZN(n423) );
  XNOR2_X2 U323 ( .A(n411), .B(n410), .ZN(n535) );
  XOR2_X1 U324 ( .A(n363), .B(n362), .Z(n571) );
  NOR2_X2 U325 ( .A1(n518), .A2(n444), .ZN(n556) );
  XOR2_X1 U326 ( .A(n422), .B(n311), .Z(n518) );
  XOR2_X1 U327 ( .A(KEYINPUT71), .B(G92GAT), .Z(n290) );
  INV_X1 U328 ( .A(KEYINPUT48), .ZN(n410) );
  NOR2_X1 U329 ( .A1(n461), .A2(n563), .ZN(n443) );
  XNOR2_X1 U330 ( .A(n441), .B(n440), .ZN(n517) );
  XNOR2_X1 U331 ( .A(n445), .B(G190GAT), .ZN(n446) );
  XNOR2_X1 U332 ( .A(n447), .B(n446), .ZN(G1351GAT) );
  XOR2_X1 U333 ( .A(KEYINPUT86), .B(G183GAT), .Z(n292) );
  XNOR2_X1 U334 ( .A(KEYINPUT85), .B(KEYINPUT19), .ZN(n291) );
  XNOR2_X1 U335 ( .A(n292), .B(n291), .ZN(n293) );
  XOR2_X1 U336 ( .A(n293), .B(KEYINPUT18), .Z(n295) );
  XNOR2_X1 U337 ( .A(KEYINPUT17), .B(KEYINPUT84), .ZN(n294) );
  XNOR2_X1 U338 ( .A(n295), .B(n294), .ZN(n422) );
  XOR2_X1 U339 ( .A(KEYINPUT83), .B(G176GAT), .Z(n297) );
  XNOR2_X1 U340 ( .A(G15GAT), .B(G190GAT), .ZN(n296) );
  XNOR2_X1 U341 ( .A(n297), .B(n296), .ZN(n298) );
  XOR2_X1 U342 ( .A(n298), .B(G99GAT), .Z(n300) );
  XOR2_X1 U343 ( .A(G120GAT), .B(G71GAT), .Z(n359) );
  XNOR2_X1 U344 ( .A(G43GAT), .B(n359), .ZN(n299) );
  XNOR2_X1 U345 ( .A(n300), .B(n299), .ZN(n304) );
  XOR2_X1 U346 ( .A(KEYINPUT20), .B(KEYINPUT82), .Z(n302) );
  NAND2_X1 U347 ( .A1(G227GAT), .A2(G233GAT), .ZN(n301) );
  XNOR2_X1 U348 ( .A(n302), .B(n301), .ZN(n303) );
  XOR2_X1 U349 ( .A(n304), .B(n303), .Z(n310) );
  XNOR2_X1 U350 ( .A(G127GAT), .B(KEYINPUT80), .ZN(n305) );
  XNOR2_X1 U351 ( .A(n305), .B(KEYINPUT0), .ZN(n306) );
  XOR2_X1 U352 ( .A(n306), .B(KEYINPUT81), .Z(n308) );
  XNOR2_X1 U353 ( .A(G113GAT), .B(G134GAT), .ZN(n307) );
  XNOR2_X1 U354 ( .A(n308), .B(n307), .ZN(n435) );
  XNOR2_X1 U355 ( .A(G169GAT), .B(n435), .ZN(n309) );
  XNOR2_X1 U356 ( .A(n310), .B(n309), .ZN(n311) );
  XOR2_X1 U357 ( .A(KEYINPUT22), .B(KEYINPUT87), .Z(n313) );
  XNOR2_X1 U358 ( .A(G204GAT), .B(KEYINPUT23), .ZN(n312) );
  XNOR2_X1 U359 ( .A(n313), .B(n312), .ZN(n314) );
  XOR2_X1 U360 ( .A(n314), .B(KEYINPUT24), .Z(n316) );
  XOR2_X1 U361 ( .A(G141GAT), .B(G22GAT), .Z(n343) );
  XNOR2_X1 U362 ( .A(G50GAT), .B(n343), .ZN(n315) );
  XNOR2_X1 U363 ( .A(n316), .B(n315), .ZN(n321) );
  XNOR2_X1 U364 ( .A(G106GAT), .B(G78GAT), .ZN(n317) );
  XNOR2_X1 U365 ( .A(n317), .B(G148GAT), .ZN(n354) );
  XOR2_X1 U366 ( .A(n354), .B(KEYINPUT92), .Z(n319) );
  NAND2_X1 U367 ( .A1(G228GAT), .A2(G233GAT), .ZN(n318) );
  XNOR2_X1 U368 ( .A(n319), .B(n318), .ZN(n320) );
  XOR2_X1 U369 ( .A(n321), .B(n320), .Z(n331) );
  XNOR2_X1 U370 ( .A(KEYINPUT2), .B(KEYINPUT90), .ZN(n322) );
  XNOR2_X1 U371 ( .A(n322), .B(KEYINPUT3), .ZN(n323) );
  XOR2_X1 U372 ( .A(n323), .B(KEYINPUT91), .Z(n325) );
  XNOR2_X1 U373 ( .A(G155GAT), .B(G162GAT), .ZN(n324) );
  XNOR2_X1 U374 ( .A(n325), .B(n324), .ZN(n434) );
  XNOR2_X1 U375 ( .A(G211GAT), .B(KEYINPUT89), .ZN(n326) );
  XNOR2_X1 U376 ( .A(n326), .B(KEYINPUT88), .ZN(n327) );
  XOR2_X1 U377 ( .A(n327), .B(KEYINPUT21), .Z(n329) );
  XNOR2_X1 U378 ( .A(G197GAT), .B(G218GAT), .ZN(n328) );
  XNOR2_X1 U379 ( .A(n329), .B(n328), .ZN(n417) );
  XNOR2_X1 U380 ( .A(n434), .B(n417), .ZN(n330) );
  XNOR2_X1 U381 ( .A(n331), .B(n330), .ZN(n461) );
  XOR2_X1 U382 ( .A(KEYINPUT8), .B(G50GAT), .Z(n333) );
  XNOR2_X1 U383 ( .A(G43GAT), .B(G29GAT), .ZN(n332) );
  XNOR2_X1 U384 ( .A(n333), .B(n332), .ZN(n334) );
  XOR2_X1 U385 ( .A(KEYINPUT7), .B(n334), .Z(n399) );
  XOR2_X1 U386 ( .A(KEYINPUT29), .B(KEYINPUT66), .Z(n336) );
  NAND2_X1 U387 ( .A1(G229GAT), .A2(G233GAT), .ZN(n335) );
  XNOR2_X1 U388 ( .A(n336), .B(n335), .ZN(n337) );
  XOR2_X1 U389 ( .A(n337), .B(KEYINPUT30), .Z(n342) );
  XNOR2_X1 U390 ( .A(G169GAT), .B(G36GAT), .ZN(n338) );
  XNOR2_X1 U391 ( .A(n338), .B(G8GAT), .ZN(n418) );
  XOR2_X1 U392 ( .A(G1GAT), .B(KEYINPUT67), .Z(n340) );
  XNOR2_X1 U393 ( .A(G15GAT), .B(KEYINPUT68), .ZN(n339) );
  XNOR2_X1 U394 ( .A(n340), .B(n339), .ZN(n371) );
  XNOR2_X1 U395 ( .A(n418), .B(n371), .ZN(n341) );
  XNOR2_X1 U396 ( .A(n342), .B(n341), .ZN(n344) );
  XOR2_X1 U397 ( .A(n344), .B(n343), .Z(n346) );
  XNOR2_X1 U398 ( .A(G113GAT), .B(G197GAT), .ZN(n345) );
  XNOR2_X1 U399 ( .A(n346), .B(n345), .ZN(n347) );
  XNOR2_X1 U400 ( .A(n399), .B(n347), .ZN(n565) );
  XOR2_X1 U401 ( .A(KEYINPUT70), .B(KEYINPUT73), .Z(n349) );
  XNOR2_X1 U402 ( .A(KEYINPUT33), .B(KEYINPUT32), .ZN(n348) );
  XNOR2_X1 U403 ( .A(n349), .B(n348), .ZN(n363) );
  XOR2_X1 U404 ( .A(KEYINPUT74), .B(KEYINPUT72), .Z(n351) );
  NAND2_X1 U405 ( .A1(G230GAT), .A2(G233GAT), .ZN(n350) );
  XNOR2_X1 U406 ( .A(n351), .B(n350), .ZN(n352) );
  XOR2_X1 U407 ( .A(n352), .B(KEYINPUT31), .Z(n356) );
  XNOR2_X1 U408 ( .A(G99GAT), .B(G85GAT), .ZN(n353) );
  XNOR2_X1 U409 ( .A(n290), .B(n353), .ZN(n391) );
  XNOR2_X1 U410 ( .A(n354), .B(n391), .ZN(n355) );
  XNOR2_X1 U411 ( .A(n356), .B(n355), .ZN(n357) );
  XOR2_X1 U412 ( .A(G57GAT), .B(KEYINPUT13), .Z(n367) );
  XOR2_X1 U413 ( .A(n357), .B(n367), .Z(n361) );
  XNOR2_X1 U414 ( .A(G176GAT), .B(G204GAT), .ZN(n358) );
  XNOR2_X1 U415 ( .A(n358), .B(G64GAT), .ZN(n415) );
  XNOR2_X1 U416 ( .A(n359), .B(n415), .ZN(n360) );
  XNOR2_X1 U417 ( .A(n361), .B(n360), .ZN(n362) );
  XNOR2_X1 U418 ( .A(n571), .B(KEYINPUT41), .ZN(n540) );
  NOR2_X1 U419 ( .A1(n565), .A2(n540), .ZN(n364) );
  XNOR2_X1 U420 ( .A(n364), .B(KEYINPUT46), .ZN(n384) );
  XOR2_X1 U421 ( .A(G155GAT), .B(G71GAT), .Z(n366) );
  XNOR2_X1 U422 ( .A(G183GAT), .B(G127GAT), .ZN(n365) );
  XNOR2_X1 U423 ( .A(n366), .B(n365), .ZN(n368) );
  XOR2_X1 U424 ( .A(n368), .B(n367), .Z(n370) );
  XNOR2_X1 U425 ( .A(G22GAT), .B(G211GAT), .ZN(n369) );
  XNOR2_X1 U426 ( .A(n370), .B(n369), .ZN(n375) );
  XOR2_X1 U427 ( .A(n371), .B(KEYINPUT12), .Z(n373) );
  NAND2_X1 U428 ( .A1(G231GAT), .A2(G233GAT), .ZN(n372) );
  XNOR2_X1 U429 ( .A(n373), .B(n372), .ZN(n374) );
  XOR2_X1 U430 ( .A(n375), .B(n374), .Z(n383) );
  XOR2_X1 U431 ( .A(KEYINPUT79), .B(G64GAT), .Z(n377) );
  XNOR2_X1 U432 ( .A(G8GAT), .B(G78GAT), .ZN(n376) );
  XNOR2_X1 U433 ( .A(n377), .B(n376), .ZN(n381) );
  XOR2_X1 U434 ( .A(KEYINPUT78), .B(KEYINPUT15), .Z(n379) );
  XNOR2_X1 U435 ( .A(KEYINPUT77), .B(KEYINPUT14), .ZN(n378) );
  XNOR2_X1 U436 ( .A(n379), .B(n378), .ZN(n380) );
  XNOR2_X1 U437 ( .A(n381), .B(n380), .ZN(n382) );
  XNOR2_X1 U438 ( .A(n383), .B(n382), .ZN(n574) );
  NOR2_X1 U439 ( .A1(n384), .A2(n574), .ZN(n385) );
  XNOR2_X1 U440 ( .A(n385), .B(KEYINPUT111), .ZN(n402) );
  XOR2_X1 U441 ( .A(KEYINPUT9), .B(KEYINPUT75), .Z(n387) );
  XNOR2_X1 U442 ( .A(G218GAT), .B(G106GAT), .ZN(n386) );
  XNOR2_X1 U443 ( .A(n387), .B(n386), .ZN(n388) );
  XOR2_X1 U444 ( .A(n388), .B(KEYINPUT65), .Z(n390) );
  XOR2_X1 U445 ( .A(G190GAT), .B(KEYINPUT76), .Z(n412) );
  XNOR2_X1 U446 ( .A(G36GAT), .B(n412), .ZN(n389) );
  XNOR2_X1 U447 ( .A(n390), .B(n389), .ZN(n395) );
  XOR2_X1 U448 ( .A(n391), .B(G134GAT), .Z(n393) );
  NAND2_X1 U449 ( .A1(G232GAT), .A2(G233GAT), .ZN(n392) );
  XNOR2_X1 U450 ( .A(n393), .B(n392), .ZN(n394) );
  XOR2_X1 U451 ( .A(n395), .B(n394), .Z(n401) );
  XOR2_X1 U452 ( .A(KEYINPUT11), .B(KEYINPUT64), .Z(n397) );
  XNOR2_X1 U453 ( .A(G162GAT), .B(KEYINPUT10), .ZN(n396) );
  XNOR2_X1 U454 ( .A(n397), .B(n396), .ZN(n398) );
  XNOR2_X1 U455 ( .A(n399), .B(n398), .ZN(n400) );
  XNOR2_X1 U456 ( .A(n401), .B(n400), .ZN(n547) );
  NOR2_X1 U457 ( .A1(n402), .A2(n547), .ZN(n403) );
  XNOR2_X1 U458 ( .A(n403), .B(KEYINPUT47), .ZN(n409) );
  XNOR2_X1 U459 ( .A(KEYINPUT45), .B(KEYINPUT112), .ZN(n405) );
  XNOR2_X1 U460 ( .A(KEYINPUT36), .B(n547), .ZN(n576) );
  NAND2_X1 U461 ( .A1(n574), .A2(n576), .ZN(n404) );
  XNOR2_X1 U462 ( .A(n405), .B(n404), .ZN(n406) );
  NOR2_X1 U463 ( .A1(n571), .A2(n406), .ZN(n407) );
  XNOR2_X1 U464 ( .A(KEYINPUT69), .B(n565), .ZN(n551) );
  INV_X1 U465 ( .A(n551), .ZN(n448) );
  NAND2_X1 U466 ( .A1(n407), .A2(n448), .ZN(n408) );
  NAND2_X1 U467 ( .A1(n409), .A2(n408), .ZN(n411) );
  XOR2_X1 U468 ( .A(n412), .B(G92GAT), .Z(n414) );
  NAND2_X1 U469 ( .A1(G226GAT), .A2(G233GAT), .ZN(n413) );
  XNOR2_X1 U470 ( .A(n414), .B(n413), .ZN(n416) );
  XOR2_X1 U471 ( .A(n416), .B(n415), .Z(n420) );
  XNOR2_X1 U472 ( .A(n418), .B(n417), .ZN(n419) );
  XNOR2_X1 U473 ( .A(n420), .B(n419), .ZN(n421) );
  XOR2_X1 U474 ( .A(n422), .B(n421), .Z(n496) );
  XNOR2_X1 U475 ( .A(KEYINPUT54), .B(n423), .ZN(n442) );
  XOR2_X1 U476 ( .A(G57GAT), .B(G148GAT), .Z(n425) );
  XNOR2_X1 U477 ( .A(G141GAT), .B(G120GAT), .ZN(n424) );
  XNOR2_X1 U478 ( .A(n425), .B(n424), .ZN(n427) );
  XOR2_X1 U479 ( .A(G29GAT), .B(G85GAT), .Z(n426) );
  XNOR2_X1 U480 ( .A(n427), .B(n426), .ZN(n439) );
  XOR2_X1 U481 ( .A(KEYINPUT94), .B(KEYINPUT95), .Z(n429) );
  XNOR2_X1 U482 ( .A(G1GAT), .B(KEYINPUT4), .ZN(n428) );
  XNOR2_X1 U483 ( .A(n429), .B(n428), .ZN(n433) );
  XOR2_X1 U484 ( .A(KEYINPUT93), .B(KEYINPUT5), .Z(n431) );
  XNOR2_X1 U485 ( .A(KEYINPUT6), .B(KEYINPUT1), .ZN(n430) );
  XNOR2_X1 U486 ( .A(n431), .B(n430), .ZN(n432) );
  XOR2_X1 U487 ( .A(n433), .B(n432), .Z(n437) );
  XNOR2_X1 U488 ( .A(n435), .B(n434), .ZN(n436) );
  XNOR2_X1 U489 ( .A(n437), .B(n436), .ZN(n438) );
  XNOR2_X1 U490 ( .A(n439), .B(n438), .ZN(n441) );
  NAND2_X1 U491 ( .A1(G225GAT), .A2(G233GAT), .ZN(n440) );
  NAND2_X1 U492 ( .A1(n442), .A2(n517), .ZN(n563) );
  XNOR2_X1 U493 ( .A(n443), .B(KEYINPUT55), .ZN(n444) );
  NAND2_X1 U494 ( .A1(n556), .A2(n547), .ZN(n447) );
  XOR2_X1 U495 ( .A(KEYINPUT58), .B(KEYINPUT123), .Z(n445) );
  NOR2_X1 U496 ( .A1(n571), .A2(n448), .ZN(n479) );
  INV_X1 U497 ( .A(n574), .ZN(n545) );
  NOR2_X1 U498 ( .A1(n547), .A2(n545), .ZN(n449) );
  XNOR2_X1 U499 ( .A(KEYINPUT16), .B(n449), .ZN(n466) );
  NOR2_X1 U500 ( .A1(n518), .A2(n496), .ZN(n450) );
  XNOR2_X1 U501 ( .A(n450), .B(KEYINPUT98), .ZN(n451) );
  NOR2_X1 U502 ( .A1(n461), .A2(n451), .ZN(n454) );
  XOR2_X1 U503 ( .A(KEYINPUT99), .B(KEYINPUT100), .Z(n452) );
  XNOR2_X1 U504 ( .A(KEYINPUT25), .B(n452), .ZN(n453) );
  XNOR2_X1 U505 ( .A(n454), .B(n453), .ZN(n455) );
  NAND2_X1 U506 ( .A1(n455), .A2(n517), .ZN(n460) );
  XOR2_X1 U507 ( .A(KEYINPUT96), .B(KEYINPUT26), .Z(n457) );
  NAND2_X1 U508 ( .A1(n461), .A2(n518), .ZN(n456) );
  XOR2_X1 U509 ( .A(n457), .B(n456), .Z(n562) );
  INV_X1 U510 ( .A(n562), .ZN(n458) );
  XOR2_X1 U511 ( .A(n496), .B(KEYINPUT27), .Z(n462) );
  NAND2_X1 U512 ( .A1(n458), .A2(n462), .ZN(n534) );
  XNOR2_X1 U513 ( .A(KEYINPUT97), .B(n534), .ZN(n459) );
  NOR2_X1 U514 ( .A1(n460), .A2(n459), .ZN(n465) );
  XOR2_X1 U515 ( .A(n461), .B(KEYINPUT28), .Z(n499) );
  NAND2_X1 U516 ( .A1(n462), .A2(n499), .ZN(n516) );
  INV_X1 U517 ( .A(n518), .ZN(n510) );
  NOR2_X1 U518 ( .A1(n516), .A2(n510), .ZN(n463) );
  NOR2_X1 U519 ( .A1(n517), .A2(n463), .ZN(n464) );
  NOR2_X1 U520 ( .A1(n465), .A2(n464), .ZN(n476) );
  NAND2_X1 U521 ( .A1(n466), .A2(n476), .ZN(n467) );
  XNOR2_X1 U522 ( .A(n467), .B(KEYINPUT101), .ZN(n492) );
  NAND2_X1 U523 ( .A1(n479), .A2(n492), .ZN(n474) );
  NOR2_X1 U524 ( .A1(n517), .A2(n474), .ZN(n469) );
  XNOR2_X1 U525 ( .A(KEYINPUT102), .B(KEYINPUT34), .ZN(n468) );
  XNOR2_X1 U526 ( .A(n469), .B(n468), .ZN(n470) );
  XOR2_X1 U527 ( .A(G1GAT), .B(n470), .Z(G1324GAT) );
  NOR2_X1 U528 ( .A1(n496), .A2(n474), .ZN(n471) );
  XOR2_X1 U529 ( .A(G8GAT), .B(n471), .Z(G1325GAT) );
  NOR2_X1 U530 ( .A1(n518), .A2(n474), .ZN(n473) );
  XNOR2_X1 U531 ( .A(G15GAT), .B(KEYINPUT35), .ZN(n472) );
  XNOR2_X1 U532 ( .A(n473), .B(n472), .ZN(G1326GAT) );
  NOR2_X1 U533 ( .A1(n499), .A2(n474), .ZN(n475) );
  XOR2_X1 U534 ( .A(G22GAT), .B(n475), .Z(G1327GAT) );
  NAND2_X1 U535 ( .A1(n476), .A2(n576), .ZN(n477) );
  NOR2_X1 U536 ( .A1(n574), .A2(n477), .ZN(n478) );
  XOR2_X1 U537 ( .A(KEYINPUT37), .B(n478), .Z(n503) );
  NAND2_X1 U538 ( .A1(n503), .A2(n479), .ZN(n480) );
  XNOR2_X1 U539 ( .A(KEYINPUT38), .B(n480), .ZN(n488) );
  NOR2_X1 U540 ( .A1(n488), .A2(n517), .ZN(n484) );
  XOR2_X1 U541 ( .A(KEYINPUT103), .B(KEYINPUT104), .Z(n482) );
  XNOR2_X1 U542 ( .A(G29GAT), .B(KEYINPUT39), .ZN(n481) );
  XNOR2_X1 U543 ( .A(n482), .B(n481), .ZN(n483) );
  XNOR2_X1 U544 ( .A(n484), .B(n483), .ZN(G1328GAT) );
  NOR2_X1 U545 ( .A1(n496), .A2(n488), .ZN(n485) );
  XOR2_X1 U546 ( .A(G36GAT), .B(n485), .Z(G1329GAT) );
  NOR2_X1 U547 ( .A1(n518), .A2(n488), .ZN(n486) );
  XOR2_X1 U548 ( .A(KEYINPUT40), .B(n486), .Z(n487) );
  XNOR2_X1 U549 ( .A(G43GAT), .B(n487), .ZN(G1330GAT) );
  XNOR2_X1 U550 ( .A(G50GAT), .B(KEYINPUT105), .ZN(n490) );
  NOR2_X1 U551 ( .A1(n499), .A2(n488), .ZN(n489) );
  XNOR2_X1 U552 ( .A(n490), .B(n489), .ZN(G1331GAT) );
  XNOR2_X1 U553 ( .A(G57GAT), .B(KEYINPUT42), .ZN(n495) );
  INV_X1 U554 ( .A(n517), .ZN(n536) );
  XOR2_X1 U555 ( .A(KEYINPUT106), .B(n540), .Z(n555) );
  NAND2_X1 U556 ( .A1(n555), .A2(n565), .ZN(n491) );
  XNOR2_X1 U557 ( .A(n491), .B(KEYINPUT107), .ZN(n504) );
  NAND2_X1 U558 ( .A1(n504), .A2(n492), .ZN(n493) );
  XOR2_X1 U559 ( .A(KEYINPUT108), .B(n493), .Z(n500) );
  NAND2_X1 U560 ( .A1(n536), .A2(n500), .ZN(n494) );
  XNOR2_X1 U561 ( .A(n495), .B(n494), .ZN(G1332GAT) );
  INV_X1 U562 ( .A(n496), .ZN(n507) );
  NAND2_X1 U563 ( .A1(n507), .A2(n500), .ZN(n497) );
  XNOR2_X1 U564 ( .A(G64GAT), .B(n497), .ZN(G1333GAT) );
  NAND2_X1 U565 ( .A1(n500), .A2(n510), .ZN(n498) );
  XNOR2_X1 U566 ( .A(n498), .B(G71GAT), .ZN(G1334GAT) );
  XOR2_X1 U567 ( .A(G78GAT), .B(KEYINPUT43), .Z(n502) );
  INV_X1 U568 ( .A(n499), .ZN(n513) );
  NAND2_X1 U569 ( .A1(n500), .A2(n513), .ZN(n501) );
  XNOR2_X1 U570 ( .A(n502), .B(n501), .ZN(G1335GAT) );
  NAND2_X1 U571 ( .A1(n504), .A2(n503), .ZN(n505) );
  XNOR2_X1 U572 ( .A(n505), .B(KEYINPUT109), .ZN(n512) );
  NAND2_X1 U573 ( .A1(n512), .A2(n536), .ZN(n506) );
  XNOR2_X1 U574 ( .A(G85GAT), .B(n506), .ZN(G1336GAT) );
  NAND2_X1 U575 ( .A1(n507), .A2(n512), .ZN(n508) );
  XNOR2_X1 U576 ( .A(n508), .B(KEYINPUT110), .ZN(n509) );
  XNOR2_X1 U577 ( .A(G92GAT), .B(n509), .ZN(G1337GAT) );
  NAND2_X1 U578 ( .A1(n510), .A2(n512), .ZN(n511) );
  XNOR2_X1 U579 ( .A(n511), .B(G99GAT), .ZN(G1338GAT) );
  NAND2_X1 U580 ( .A1(n513), .A2(n512), .ZN(n514) );
  XNOR2_X1 U581 ( .A(n514), .B(KEYINPUT44), .ZN(n515) );
  XNOR2_X1 U582 ( .A(G106GAT), .B(n515), .ZN(G1339GAT) );
  NOR2_X1 U583 ( .A1(n535), .A2(n516), .ZN(n520) );
  NOR2_X1 U584 ( .A1(n518), .A2(n517), .ZN(n519) );
  NAND2_X1 U585 ( .A1(n520), .A2(n519), .ZN(n521) );
  XNOR2_X1 U586 ( .A(KEYINPUT113), .B(n521), .ZN(n529) );
  NAND2_X1 U587 ( .A1(n529), .A2(n551), .ZN(n522) );
  XNOR2_X1 U588 ( .A(n522), .B(KEYINPUT114), .ZN(n523) );
  XNOR2_X1 U589 ( .A(G113GAT), .B(n523), .ZN(G1340GAT) );
  XOR2_X1 U590 ( .A(KEYINPUT49), .B(KEYINPUT115), .Z(n525) );
  NAND2_X1 U591 ( .A1(n529), .A2(n555), .ZN(n524) );
  XNOR2_X1 U592 ( .A(n525), .B(n524), .ZN(n526) );
  XOR2_X1 U593 ( .A(G120GAT), .B(n526), .Z(G1341GAT) );
  NAND2_X1 U594 ( .A1(n529), .A2(n574), .ZN(n527) );
  XNOR2_X1 U595 ( .A(n527), .B(KEYINPUT50), .ZN(n528) );
  XNOR2_X1 U596 ( .A(G127GAT), .B(n528), .ZN(G1342GAT) );
  XOR2_X1 U597 ( .A(KEYINPUT117), .B(KEYINPUT51), .Z(n531) );
  NAND2_X1 U598 ( .A1(n529), .A2(n547), .ZN(n530) );
  XNOR2_X1 U599 ( .A(n531), .B(n530), .ZN(n533) );
  XOR2_X1 U600 ( .A(G134GAT), .B(KEYINPUT116), .Z(n532) );
  XNOR2_X1 U601 ( .A(n533), .B(n532), .ZN(G1343GAT) );
  NOR2_X1 U602 ( .A1(n535), .A2(n534), .ZN(n537) );
  NAND2_X1 U603 ( .A1(n537), .A2(n536), .ZN(n548) );
  NOR2_X1 U604 ( .A1(n565), .A2(n548), .ZN(n538) );
  XOR2_X1 U605 ( .A(G141GAT), .B(n538), .Z(n539) );
  XNOR2_X1 U606 ( .A(KEYINPUT118), .B(n539), .ZN(G1344GAT) );
  NOR2_X1 U607 ( .A1(n548), .A2(n540), .ZN(n544) );
  XOR2_X1 U608 ( .A(KEYINPUT53), .B(KEYINPUT52), .Z(n542) );
  XNOR2_X1 U609 ( .A(G148GAT), .B(KEYINPUT119), .ZN(n541) );
  XNOR2_X1 U610 ( .A(n542), .B(n541), .ZN(n543) );
  XNOR2_X1 U611 ( .A(n544), .B(n543), .ZN(G1345GAT) );
  NOR2_X1 U612 ( .A1(n545), .A2(n548), .ZN(n546) );
  XOR2_X1 U613 ( .A(G155GAT), .B(n546), .Z(G1346GAT) );
  INV_X1 U614 ( .A(n547), .ZN(n549) );
  NOR2_X1 U615 ( .A1(n549), .A2(n548), .ZN(n550) );
  XOR2_X1 U616 ( .A(G162GAT), .B(n550), .Z(G1347GAT) );
  NAND2_X1 U617 ( .A1(n551), .A2(n556), .ZN(n552) );
  XNOR2_X1 U618 ( .A(G169GAT), .B(n552), .ZN(G1348GAT) );
  XOR2_X1 U619 ( .A(KEYINPUT122), .B(KEYINPUT121), .Z(n554) );
  XNOR2_X1 U620 ( .A(KEYINPUT56), .B(KEYINPUT57), .ZN(n553) );
  XNOR2_X1 U621 ( .A(n554), .B(n553), .ZN(n560) );
  XOR2_X1 U622 ( .A(G176GAT), .B(KEYINPUT120), .Z(n558) );
  NAND2_X1 U623 ( .A1(n556), .A2(n555), .ZN(n557) );
  XNOR2_X1 U624 ( .A(n558), .B(n557), .ZN(n559) );
  XNOR2_X1 U625 ( .A(n560), .B(n559), .ZN(G1349GAT) );
  NAND2_X1 U626 ( .A1(n556), .A2(n574), .ZN(n561) );
  XNOR2_X1 U627 ( .A(n561), .B(G183GAT), .ZN(G1350GAT) );
  NOR2_X1 U628 ( .A1(n563), .A2(n562), .ZN(n577) );
  INV_X1 U629 ( .A(n577), .ZN(n564) );
  NOR2_X1 U630 ( .A1(n565), .A2(n564), .ZN(n570) );
  XOR2_X1 U631 ( .A(KEYINPUT124), .B(KEYINPUT125), .Z(n567) );
  XNOR2_X1 U632 ( .A(G197GAT), .B(KEYINPUT59), .ZN(n566) );
  XNOR2_X1 U633 ( .A(n567), .B(n566), .ZN(n568) );
  XNOR2_X1 U634 ( .A(KEYINPUT60), .B(n568), .ZN(n569) );
  XNOR2_X1 U635 ( .A(n570), .B(n569), .ZN(G1352GAT) );
  XOR2_X1 U636 ( .A(G204GAT), .B(KEYINPUT61), .Z(n573) );
  NAND2_X1 U637 ( .A1(n577), .A2(n571), .ZN(n572) );
  XNOR2_X1 U638 ( .A(n573), .B(n572), .ZN(G1353GAT) );
  NAND2_X1 U639 ( .A1(n577), .A2(n574), .ZN(n575) );
  XNOR2_X1 U640 ( .A(n575), .B(G211GAT), .ZN(G1354GAT) );
  XNOR2_X1 U641 ( .A(G218GAT), .B(KEYINPUT62), .ZN(n581) );
  XOR2_X1 U642 ( .A(KEYINPUT126), .B(KEYINPUT127), .Z(n579) );
  NAND2_X1 U643 ( .A1(n577), .A2(n576), .ZN(n578) );
  XNOR2_X1 U644 ( .A(n579), .B(n578), .ZN(n580) );
  XNOR2_X1 U645 ( .A(n581), .B(n580), .ZN(G1355GAT) );
endmodule

