//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 0 0 1 0 1 1 1 0 0 0 0 1 1 0 1 0 0 1 0 1 0 1 0 0 1 0 1 1 1 1 0 1 0 1 1 0 0 0 0 1 0 1 0 1 1 0 0 1 1 0 1 1 1 0 0 0 0 1 1 0 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:33:19 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n447, new_n451, new_n452, new_n453, new_n454, new_n455,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n492, new_n493, new_n494, new_n495, new_n496,
    new_n497, new_n498, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n508, new_n509, new_n510, new_n511,
    new_n512, new_n513, new_n514, new_n515, new_n516, new_n518, new_n519,
    new_n520, new_n521, new_n522, new_n523, new_n524, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n547, new_n548, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n569,
    new_n570, new_n571, new_n573, new_n574, new_n575, new_n576, new_n577,
    new_n578, new_n579, new_n580, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n605, new_n608, new_n610, new_n611, new_n612,
    new_n613, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1207, new_n1208,
    new_n1209, new_n1210;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  XOR2_X1   g012(.A(KEYINPUT64), .B(G69), .Z(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  XNOR2_X1  g020(.A(KEYINPUT65), .B(KEYINPUT1), .ZN(new_n446));
  AND2_X1   g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XNOR2_X1  g022(.A(new_n446), .B(new_n447), .ZN(G223));
  NAND2_X1  g023(.A1(new_n447), .A2(G567), .ZN(G234));
  NAND2_X1  g024(.A1(new_n447), .A2(G2106), .ZN(G217));
  NOR4_X1   g025(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n451));
  XNOR2_X1  g026(.A(new_n451), .B(KEYINPUT2), .ZN(new_n452));
  INV_X1    g027(.A(new_n452), .ZN(new_n453));
  NOR4_X1   g028(.A1(G235), .A2(G237), .A3(G238), .A4(G236), .ZN(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(new_n455));
  NOR2_X1   g030(.A1(new_n453), .A2(new_n455), .ZN(G325));
  INV_X1    g031(.A(G325), .ZN(G261));
  AOI22_X1  g032(.A1(new_n453), .A2(G2106), .B1(G567), .B2(new_n455), .ZN(G319));
  INV_X1    g033(.A(G2105), .ZN(new_n459));
  INV_X1    g034(.A(KEYINPUT3), .ZN(new_n460));
  INV_X1    g035(.A(G2104), .ZN(new_n461));
  NAND2_X1  g036(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  NAND2_X1  g037(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n464), .A2(G125), .ZN(new_n465));
  NAND2_X1  g040(.A1(G113), .A2(G2104), .ZN(new_n466));
  AOI21_X1  g041(.A(new_n459), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  INV_X1    g042(.A(new_n463), .ZN(new_n468));
  NOR2_X1   g043(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n469));
  OAI211_X1 g044(.A(G137), .B(new_n459), .C1(new_n468), .C2(new_n469), .ZN(new_n470));
  NOR2_X1   g045(.A1(new_n461), .A2(G2105), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n471), .A2(G101), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n470), .A2(new_n472), .ZN(new_n473));
  NOR2_X1   g048(.A1(new_n467), .A2(new_n473), .ZN(G160));
  OR2_X1    g049(.A1(G100), .A2(G2105), .ZN(new_n475));
  OAI211_X1 g050(.A(new_n475), .B(G2104), .C1(G112), .C2(new_n459), .ZN(new_n476));
  AOI21_X1  g051(.A(new_n459), .B1(new_n462), .B2(new_n463), .ZN(new_n477));
  INV_X1    g052(.A(new_n477), .ZN(new_n478));
  INV_X1    g053(.A(G124), .ZN(new_n479));
  OAI21_X1  g054(.A(new_n476), .B1(new_n478), .B2(new_n479), .ZN(new_n480));
  AOI21_X1  g055(.A(G2105), .B1(new_n462), .B2(new_n463), .ZN(new_n481));
  AOI21_X1  g056(.A(new_n480), .B1(G136), .B2(new_n481), .ZN(G162));
  OAI211_X1 g057(.A(G126), .B(G2105), .C1(new_n468), .C2(new_n469), .ZN(new_n483));
  OR2_X1    g058(.A1(G102), .A2(G2105), .ZN(new_n484));
  OAI211_X1 g059(.A(new_n484), .B(G2104), .C1(G114), .C2(new_n459), .ZN(new_n485));
  NAND2_X1  g060(.A1(new_n483), .A2(new_n485), .ZN(new_n486));
  OAI211_X1 g061(.A(G138), .B(new_n459), .C1(new_n468), .C2(new_n469), .ZN(new_n487));
  NAND2_X1  g062(.A1(new_n487), .A2(KEYINPUT4), .ZN(new_n488));
  INV_X1    g063(.A(KEYINPUT4), .ZN(new_n489));
  NAND3_X1  g064(.A1(new_n481), .A2(new_n489), .A3(G138), .ZN(new_n490));
  AOI21_X1  g065(.A(new_n486), .B1(new_n488), .B2(new_n490), .ZN(G164));
  INV_X1    g066(.A(G543), .ZN(new_n492));
  INV_X1    g067(.A(KEYINPUT6), .ZN(new_n493));
  INV_X1    g068(.A(G651), .ZN(new_n494));
  OAI21_X1  g069(.A(new_n493), .B1(new_n494), .B2(KEYINPUT66), .ZN(new_n495));
  INV_X1    g070(.A(KEYINPUT66), .ZN(new_n496));
  NAND3_X1  g071(.A1(new_n496), .A2(KEYINPUT6), .A3(G651), .ZN(new_n497));
  AOI21_X1  g072(.A(new_n492), .B1(new_n495), .B2(new_n497), .ZN(new_n498));
  NAND2_X1  g073(.A1(new_n498), .A2(G50), .ZN(new_n499));
  INV_X1    g074(.A(G88), .ZN(new_n500));
  NAND2_X1  g075(.A1(new_n495), .A2(new_n497), .ZN(new_n501));
  XNOR2_X1  g076(.A(KEYINPUT5), .B(G543), .ZN(new_n502));
  NAND2_X1  g077(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  OAI21_X1  g078(.A(new_n499), .B1(new_n500), .B2(new_n503), .ZN(new_n504));
  AOI22_X1  g079(.A1(new_n502), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n505));
  NOR2_X1   g080(.A1(new_n505), .A2(new_n494), .ZN(new_n506));
  NOR2_X1   g081(.A1(new_n504), .A2(new_n506), .ZN(G166));
  NAND2_X1  g082(.A1(new_n498), .A2(G51), .ZN(new_n508));
  NAND3_X1  g083(.A1(new_n501), .A2(G89), .A3(new_n502), .ZN(new_n509));
  AND2_X1   g084(.A1(G63), .A2(G651), .ZN(new_n510));
  NAND3_X1  g085(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n511));
  NAND2_X1  g086(.A1(new_n511), .A2(KEYINPUT7), .ZN(new_n512));
  INV_X1    g087(.A(KEYINPUT7), .ZN(new_n513));
  NAND4_X1  g088(.A1(new_n513), .A2(G76), .A3(G543), .A4(G651), .ZN(new_n514));
  AOI22_X1  g089(.A1(new_n502), .A2(new_n510), .B1(new_n512), .B2(new_n514), .ZN(new_n515));
  NAND3_X1  g090(.A1(new_n508), .A2(new_n509), .A3(new_n515), .ZN(new_n516));
  XNOR2_X1  g091(.A(new_n516), .B(KEYINPUT67), .ZN(G168));
  AOI22_X1  g092(.A1(new_n502), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n518));
  NOR2_X1   g093(.A1(new_n518), .A2(new_n494), .ZN(new_n519));
  NAND2_X1  g094(.A1(new_n519), .A2(KEYINPUT68), .ZN(new_n520));
  INV_X1    g095(.A(new_n503), .ZN(new_n521));
  AOI22_X1  g096(.A1(new_n521), .A2(G90), .B1(G52), .B2(new_n498), .ZN(new_n522));
  NAND2_X1  g097(.A1(new_n520), .A2(new_n522), .ZN(new_n523));
  NOR2_X1   g098(.A1(new_n519), .A2(KEYINPUT68), .ZN(new_n524));
  NOR2_X1   g099(.A1(new_n523), .A2(new_n524), .ZN(G171));
  INV_X1    g100(.A(KEYINPUT69), .ZN(new_n526));
  INV_X1    g101(.A(G56), .ZN(new_n527));
  INV_X1    g102(.A(KEYINPUT5), .ZN(new_n528));
  NAND2_X1  g103(.A1(new_n528), .A2(new_n492), .ZN(new_n529));
  NAND2_X1  g104(.A1(KEYINPUT5), .A2(G543), .ZN(new_n530));
  AOI21_X1  g105(.A(new_n527), .B1(new_n529), .B2(new_n530), .ZN(new_n531));
  INV_X1    g106(.A(G68), .ZN(new_n532));
  NOR2_X1   g107(.A1(new_n532), .A2(new_n492), .ZN(new_n533));
  OAI211_X1 g108(.A(new_n526), .B(G651), .C1(new_n531), .C2(new_n533), .ZN(new_n534));
  NAND3_X1  g109(.A1(new_n501), .A2(G81), .A3(new_n502), .ZN(new_n535));
  NAND2_X1  g110(.A1(new_n498), .A2(G43), .ZN(new_n536));
  NAND3_X1  g111(.A1(new_n534), .A2(new_n535), .A3(new_n536), .ZN(new_n537));
  AND2_X1   g112(.A1(KEYINPUT5), .A2(G543), .ZN(new_n538));
  NOR2_X1   g113(.A1(KEYINPUT5), .A2(G543), .ZN(new_n539));
  NOR2_X1   g114(.A1(new_n538), .A2(new_n539), .ZN(new_n540));
  OAI22_X1  g115(.A1(new_n540), .A2(new_n527), .B1(new_n532), .B2(new_n492), .ZN(new_n541));
  AOI21_X1  g116(.A(new_n526), .B1(new_n541), .B2(G651), .ZN(new_n542));
  NOR2_X1   g117(.A1(new_n537), .A2(new_n542), .ZN(new_n543));
  NAND2_X1  g118(.A1(new_n543), .A2(G860), .ZN(new_n544));
  XNOR2_X1  g119(.A(new_n544), .B(KEYINPUT70), .ZN(G153));
  NAND4_X1  g120(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g121(.A1(G1), .A2(G3), .ZN(new_n547));
  XNOR2_X1  g122(.A(new_n547), .B(KEYINPUT8), .ZN(new_n548));
  NAND4_X1  g123(.A1(G319), .A2(G483), .A3(G661), .A4(new_n548), .ZN(G188));
  AND3_X1   g124(.A1(new_n496), .A2(KEYINPUT6), .A3(G651), .ZN(new_n550));
  AOI21_X1  g125(.A(KEYINPUT6), .B1(new_n496), .B2(G651), .ZN(new_n551));
  OAI211_X1 g126(.A(G53), .B(G543), .C1(new_n550), .C2(new_n551), .ZN(new_n552));
  NAND2_X1  g127(.A1(new_n552), .A2(KEYINPUT9), .ZN(new_n553));
  INV_X1    g128(.A(KEYINPUT9), .ZN(new_n554));
  NAND3_X1  g129(.A1(new_n498), .A2(new_n554), .A3(G53), .ZN(new_n555));
  NAND2_X1  g130(.A1(new_n553), .A2(new_n555), .ZN(new_n556));
  INV_X1    g131(.A(G65), .ZN(new_n557));
  OAI21_X1  g132(.A(KEYINPUT71), .B1(new_n538), .B2(new_n539), .ZN(new_n558));
  INV_X1    g133(.A(KEYINPUT71), .ZN(new_n559));
  NAND3_X1  g134(.A1(new_n529), .A2(new_n559), .A3(new_n530), .ZN(new_n560));
  AOI21_X1  g135(.A(new_n557), .B1(new_n558), .B2(new_n560), .ZN(new_n561));
  AND2_X1   g136(.A1(G78), .A2(G543), .ZN(new_n562));
  OAI21_X1  g137(.A(G651), .B1(new_n561), .B2(new_n562), .ZN(new_n563));
  NAND2_X1  g138(.A1(new_n521), .A2(G91), .ZN(new_n564));
  NAND3_X1  g139(.A1(new_n556), .A2(new_n563), .A3(new_n564), .ZN(G299));
  INV_X1    g140(.A(G171), .ZN(G301));
  INV_X1    g141(.A(G168), .ZN(G286));
  INV_X1    g142(.A(G166), .ZN(G303));
  NAND2_X1  g143(.A1(new_n521), .A2(G87), .ZN(new_n569));
  NAND2_X1  g144(.A1(new_n498), .A2(G49), .ZN(new_n570));
  OAI21_X1  g145(.A(G651), .B1(new_n502), .B2(G74), .ZN(new_n571));
  NAND3_X1  g146(.A1(new_n569), .A2(new_n570), .A3(new_n571), .ZN(G288));
  NAND2_X1  g147(.A1(new_n498), .A2(G48), .ZN(new_n573));
  INV_X1    g148(.A(KEYINPUT72), .ZN(new_n574));
  NAND2_X1  g149(.A1(G73), .A2(G543), .ZN(new_n575));
  INV_X1    g150(.A(G61), .ZN(new_n576));
  OAI21_X1  g151(.A(new_n575), .B1(new_n540), .B2(new_n576), .ZN(new_n577));
  AOI22_X1  g152(.A1(new_n573), .A2(new_n574), .B1(new_n577), .B2(G651), .ZN(new_n578));
  NAND2_X1  g153(.A1(new_n521), .A2(G86), .ZN(new_n579));
  NAND3_X1  g154(.A1(new_n498), .A2(KEYINPUT72), .A3(G48), .ZN(new_n580));
  NAND3_X1  g155(.A1(new_n578), .A2(new_n579), .A3(new_n580), .ZN(G305));
  NAND2_X1  g156(.A1(G72), .A2(G543), .ZN(new_n582));
  INV_X1    g157(.A(G60), .ZN(new_n583));
  OAI21_X1  g158(.A(new_n582), .B1(new_n540), .B2(new_n583), .ZN(new_n584));
  AOI22_X1  g159(.A1(new_n521), .A2(G85), .B1(new_n584), .B2(G651), .ZN(new_n585));
  NAND2_X1  g160(.A1(new_n498), .A2(G47), .ZN(new_n586));
  AND2_X1   g161(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  INV_X1    g162(.A(new_n587), .ZN(G290));
  INV_X1    g163(.A(G868), .ZN(new_n589));
  OR3_X1    g164(.A1(G171), .A2(KEYINPUT73), .A3(new_n589), .ZN(new_n590));
  OAI21_X1  g165(.A(KEYINPUT73), .B1(G171), .B2(new_n589), .ZN(new_n591));
  OAI211_X1 g166(.A(new_n502), .B(G92), .C1(new_n550), .C2(new_n551), .ZN(new_n592));
  INV_X1    g167(.A(KEYINPUT10), .ZN(new_n593));
  NAND2_X1  g168(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  NAND4_X1  g169(.A1(new_n501), .A2(KEYINPUT10), .A3(G92), .A4(new_n502), .ZN(new_n595));
  NAND2_X1  g170(.A1(new_n594), .A2(new_n595), .ZN(new_n596));
  INV_X1    g171(.A(G66), .ZN(new_n597));
  AOI21_X1  g172(.A(new_n597), .B1(new_n558), .B2(new_n560), .ZN(new_n598));
  AND2_X1   g173(.A1(G79), .A2(G543), .ZN(new_n599));
  OAI21_X1  g174(.A(G651), .B1(new_n598), .B2(new_n599), .ZN(new_n600));
  NAND2_X1  g175(.A1(new_n498), .A2(G54), .ZN(new_n601));
  AND3_X1   g176(.A1(new_n596), .A2(new_n600), .A3(new_n601), .ZN(new_n602));
  OAI211_X1 g177(.A(new_n590), .B(new_n591), .C1(G868), .C2(new_n602), .ZN(G284));
  OAI211_X1 g178(.A(new_n590), .B(new_n591), .C1(G868), .C2(new_n602), .ZN(G321));
  NOR2_X1   g179(.A1(G299), .A2(G868), .ZN(new_n605));
  AOI21_X1  g180(.A(new_n605), .B1(G868), .B2(G168), .ZN(G280));
  XOR2_X1   g181(.A(G280), .B(KEYINPUT74), .Z(G297));
  INV_X1    g182(.A(G559), .ZN(new_n608));
  OAI21_X1  g183(.A(new_n602), .B1(new_n608), .B2(G860), .ZN(G148));
  INV_X1    g184(.A(new_n543), .ZN(new_n610));
  NAND2_X1  g185(.A1(new_n610), .A2(new_n589), .ZN(new_n611));
  NAND3_X1  g186(.A1(new_n596), .A2(new_n600), .A3(new_n601), .ZN(new_n612));
  NOR2_X1   g187(.A1(new_n612), .A2(G559), .ZN(new_n613));
  OAI21_X1  g188(.A(new_n611), .B1(new_n613), .B2(new_n589), .ZN(G323));
  XNOR2_X1  g189(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g190(.A1(new_n464), .A2(new_n471), .ZN(new_n616));
  XNOR2_X1  g191(.A(new_n616), .B(KEYINPUT12), .ZN(new_n617));
  XNOR2_X1  g192(.A(new_n617), .B(KEYINPUT13), .ZN(new_n618));
  INV_X1    g193(.A(G2100), .ZN(new_n619));
  OR2_X1    g194(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  NAND2_X1  g195(.A1(new_n618), .A2(new_n619), .ZN(new_n621));
  NAND2_X1  g196(.A1(new_n481), .A2(G135), .ZN(new_n622));
  NAND2_X1  g197(.A1(new_n477), .A2(G123), .ZN(new_n623));
  NOR2_X1   g198(.A1(new_n459), .A2(G111), .ZN(new_n624));
  OAI21_X1  g199(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n625));
  OAI211_X1 g200(.A(new_n622), .B(new_n623), .C1(new_n624), .C2(new_n625), .ZN(new_n626));
  INV_X1    g201(.A(G2096), .ZN(new_n627));
  XNOR2_X1  g202(.A(new_n626), .B(new_n627), .ZN(new_n628));
  NAND3_X1  g203(.A1(new_n620), .A2(new_n621), .A3(new_n628), .ZN(G156));
  XNOR2_X1  g204(.A(KEYINPUT15), .B(G2435), .ZN(new_n630));
  XNOR2_X1  g205(.A(KEYINPUT76), .B(G2438), .ZN(new_n631));
  XNOR2_X1  g206(.A(new_n630), .B(new_n631), .ZN(new_n632));
  XOR2_X1   g207(.A(G2427), .B(G2430), .Z(new_n633));
  OR2_X1    g208(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  NAND2_X1  g209(.A1(new_n632), .A2(new_n633), .ZN(new_n635));
  NAND3_X1  g210(.A1(new_n634), .A2(KEYINPUT14), .A3(new_n635), .ZN(new_n636));
  XNOR2_X1  g211(.A(G1341), .B(G1348), .ZN(new_n637));
  XNOR2_X1  g212(.A(KEYINPUT75), .B(KEYINPUT16), .ZN(new_n638));
  XNOR2_X1  g213(.A(new_n637), .B(new_n638), .ZN(new_n639));
  XNOR2_X1  g214(.A(new_n636), .B(new_n639), .ZN(new_n640));
  XOR2_X1   g215(.A(G2451), .B(G2454), .Z(new_n641));
  XNOR2_X1  g216(.A(G2443), .B(G2446), .ZN(new_n642));
  XNOR2_X1  g217(.A(new_n641), .B(new_n642), .ZN(new_n643));
  NAND2_X1  g218(.A1(new_n640), .A2(new_n643), .ZN(new_n644));
  NAND2_X1  g219(.A1(new_n644), .A2(G14), .ZN(new_n645));
  NOR2_X1   g220(.A1(new_n640), .A2(new_n643), .ZN(new_n646));
  NOR2_X1   g221(.A1(new_n645), .A2(new_n646), .ZN(G401));
  XNOR2_X1  g222(.A(G2084), .B(G2090), .ZN(new_n648));
  XNOR2_X1  g223(.A(G2067), .B(G2678), .ZN(new_n649));
  XNOR2_X1  g224(.A(G2072), .B(G2078), .ZN(new_n650));
  OAI21_X1  g225(.A(new_n648), .B1(new_n649), .B2(new_n650), .ZN(new_n651));
  XNOR2_X1  g226(.A(new_n650), .B(KEYINPUT17), .ZN(new_n652));
  AOI21_X1  g227(.A(new_n651), .B1(new_n652), .B2(new_n649), .ZN(new_n653));
  XOR2_X1   g228(.A(new_n653), .B(KEYINPUT78), .Z(new_n654));
  NOR3_X1   g229(.A1(new_n652), .A2(new_n649), .A3(new_n648), .ZN(new_n655));
  XNOR2_X1  g230(.A(new_n655), .B(KEYINPUT79), .ZN(new_n656));
  INV_X1    g231(.A(new_n648), .ZN(new_n657));
  NAND3_X1  g232(.A1(new_n657), .A2(new_n649), .A3(new_n650), .ZN(new_n658));
  XOR2_X1   g233(.A(KEYINPUT77), .B(KEYINPUT18), .Z(new_n659));
  XNOR2_X1  g234(.A(new_n658), .B(new_n659), .ZN(new_n660));
  NAND3_X1  g235(.A1(new_n654), .A2(new_n656), .A3(new_n660), .ZN(new_n661));
  XNOR2_X1  g236(.A(new_n661), .B(new_n627), .ZN(new_n662));
  XNOR2_X1  g237(.A(KEYINPUT80), .B(G2100), .ZN(new_n663));
  XNOR2_X1  g238(.A(new_n662), .B(new_n663), .ZN(G227));
  XNOR2_X1  g239(.A(G1956), .B(G2474), .ZN(new_n665));
  XNOR2_X1  g240(.A(G1961), .B(G1966), .ZN(new_n666));
  AND2_X1   g241(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  XNOR2_X1  g242(.A(G1971), .B(G1976), .ZN(new_n668));
  XNOR2_X1  g243(.A(KEYINPUT81), .B(KEYINPUT19), .ZN(new_n669));
  XOR2_X1   g244(.A(new_n668), .B(new_n669), .Z(new_n670));
  NOR2_X1   g245(.A1(new_n665), .A2(new_n666), .ZN(new_n671));
  AOI21_X1  g246(.A(new_n667), .B1(new_n670), .B2(new_n671), .ZN(new_n672));
  NAND2_X1  g247(.A1(new_n670), .A2(KEYINPUT83), .ZN(new_n673));
  XNOR2_X1  g248(.A(new_n672), .B(new_n673), .ZN(new_n674));
  XNOR2_X1  g249(.A(new_n668), .B(new_n669), .ZN(new_n675));
  NAND2_X1  g250(.A1(new_n675), .A2(new_n671), .ZN(new_n676));
  XOR2_X1   g251(.A(KEYINPUT82), .B(KEYINPUT20), .Z(new_n677));
  XNOR2_X1  g252(.A(new_n676), .B(new_n677), .ZN(new_n678));
  NAND2_X1  g253(.A1(new_n674), .A2(new_n678), .ZN(new_n679));
  XNOR2_X1  g254(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n680));
  XNOR2_X1  g255(.A(new_n679), .B(new_n680), .ZN(new_n681));
  XOR2_X1   g256(.A(G1991), .B(G1996), .Z(new_n682));
  XNOR2_X1  g257(.A(new_n682), .B(KEYINPUT84), .ZN(new_n683));
  XNOR2_X1  g258(.A(new_n681), .B(new_n683), .ZN(new_n684));
  XNOR2_X1  g259(.A(G1981), .B(G1986), .ZN(new_n685));
  XNOR2_X1  g260(.A(new_n684), .B(new_n685), .ZN(G229));
  NOR2_X1   g261(.A1(G29), .A2(G35), .ZN(new_n687));
  AOI21_X1  g262(.A(new_n687), .B1(G162), .B2(G29), .ZN(new_n688));
  XNOR2_X1  g263(.A(KEYINPUT99), .B(KEYINPUT29), .ZN(new_n689));
  XNOR2_X1  g264(.A(new_n688), .B(new_n689), .ZN(new_n690));
  OR2_X1    g265(.A1(new_n690), .A2(G2090), .ZN(new_n691));
  NAND2_X1  g266(.A1(new_n543), .A2(G16), .ZN(new_n692));
  OAI21_X1  g267(.A(new_n692), .B1(G16), .B2(G19), .ZN(new_n693));
  XNOR2_X1  g268(.A(KEYINPUT89), .B(G1341), .ZN(new_n694));
  AOI22_X1  g269(.A1(new_n690), .A2(G2090), .B1(new_n693), .B2(new_n694), .ZN(new_n695));
  OR2_X1    g270(.A1(new_n693), .A2(new_n694), .ZN(new_n696));
  NOR2_X1   g271(.A1(G4), .A2(G16), .ZN(new_n697));
  AOI21_X1  g272(.A(new_n697), .B1(new_n602), .B2(G16), .ZN(new_n698));
  INV_X1    g273(.A(G1348), .ZN(new_n699));
  XNOR2_X1  g274(.A(new_n698), .B(new_n699), .ZN(new_n700));
  NAND4_X1  g275(.A1(new_n691), .A2(new_n695), .A3(new_n696), .A4(new_n700), .ZN(new_n701));
  INV_X1    g276(.A(G29), .ZN(new_n702));
  NAND2_X1  g277(.A1(new_n702), .A2(G26), .ZN(new_n703));
  XNOR2_X1  g278(.A(new_n703), .B(KEYINPUT92), .ZN(new_n704));
  XNOR2_X1  g279(.A(new_n704), .B(KEYINPUT28), .ZN(new_n705));
  NAND2_X1  g280(.A1(new_n477), .A2(G128), .ZN(new_n706));
  XNOR2_X1  g281(.A(new_n706), .B(KEYINPUT90), .ZN(new_n707));
  OAI21_X1  g282(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n708));
  INV_X1    g283(.A(G116), .ZN(new_n709));
  AOI21_X1  g284(.A(new_n708), .B1(new_n709), .B2(G2105), .ZN(new_n710));
  AOI21_X1  g285(.A(new_n710), .B1(G140), .B2(new_n481), .ZN(new_n711));
  NAND2_X1  g286(.A1(new_n707), .A2(new_n711), .ZN(new_n712));
  XNOR2_X1  g287(.A(new_n712), .B(KEYINPUT91), .ZN(new_n713));
  OAI21_X1  g288(.A(new_n705), .B1(new_n713), .B2(new_n702), .ZN(new_n714));
  INV_X1    g289(.A(G2067), .ZN(new_n715));
  XNOR2_X1  g290(.A(new_n714), .B(new_n715), .ZN(new_n716));
  INV_X1    g291(.A(G16), .ZN(new_n717));
  NAND2_X1  g292(.A1(new_n717), .A2(G20), .ZN(new_n718));
  XOR2_X1   g293(.A(new_n718), .B(KEYINPUT23), .Z(new_n719));
  AOI21_X1  g294(.A(new_n719), .B1(G299), .B2(G16), .ZN(new_n720));
  XNOR2_X1  g295(.A(new_n720), .B(G1956), .ZN(new_n721));
  NAND2_X1  g296(.A1(new_n716), .A2(new_n721), .ZN(new_n722));
  NAND2_X1  g297(.A1(new_n717), .A2(G21), .ZN(new_n723));
  OAI21_X1  g298(.A(new_n723), .B1(G168), .B2(new_n717), .ZN(new_n724));
  XNOR2_X1  g299(.A(new_n724), .B(G1966), .ZN(new_n725));
  OR2_X1    g300(.A1(new_n626), .A2(new_n702), .ZN(new_n726));
  AND2_X1   g301(.A1(new_n726), .A2(KEYINPUT96), .ZN(new_n727));
  NOR2_X1   g302(.A1(new_n726), .A2(KEYINPUT96), .ZN(new_n728));
  XNOR2_X1  g303(.A(KEYINPUT31), .B(G11), .ZN(new_n729));
  XOR2_X1   g304(.A(KEYINPUT30), .B(G28), .Z(new_n730));
  OAI21_X1  g305(.A(new_n729), .B1(new_n730), .B2(G29), .ZN(new_n731));
  NOR3_X1   g306(.A1(new_n727), .A2(new_n728), .A3(new_n731), .ZN(new_n732));
  INV_X1    g307(.A(KEYINPUT24), .ZN(new_n733));
  INV_X1    g308(.A(G34), .ZN(new_n734));
  AOI21_X1  g309(.A(G29), .B1(new_n733), .B2(new_n734), .ZN(new_n735));
  OAI21_X1  g310(.A(new_n735), .B1(new_n733), .B2(new_n734), .ZN(new_n736));
  OAI21_X1  g311(.A(new_n736), .B1(G160), .B2(new_n702), .ZN(new_n737));
  INV_X1    g312(.A(G2084), .ZN(new_n738));
  XNOR2_X1  g313(.A(new_n737), .B(new_n738), .ZN(new_n739));
  NOR2_X1   g314(.A1(G27), .A2(G29), .ZN(new_n740));
  AOI21_X1  g315(.A(new_n740), .B1(G164), .B2(G29), .ZN(new_n741));
  NAND2_X1  g316(.A1(new_n741), .A2(G2078), .ZN(new_n742));
  AND2_X1   g317(.A1(new_n702), .A2(G33), .ZN(new_n743));
  AND2_X1   g318(.A1(new_n464), .A2(G127), .ZN(new_n744));
  NAND2_X1  g319(.A1(G115), .A2(G2104), .ZN(new_n745));
  INV_X1    g320(.A(new_n745), .ZN(new_n746));
  OAI21_X1  g321(.A(G2105), .B1(new_n744), .B2(new_n746), .ZN(new_n747));
  NAND2_X1  g322(.A1(new_n481), .A2(G139), .ZN(new_n748));
  NAND3_X1  g323(.A1(new_n459), .A2(G103), .A3(G2104), .ZN(new_n749));
  XOR2_X1   g324(.A(new_n749), .B(KEYINPUT25), .Z(new_n750));
  NAND3_X1  g325(.A1(new_n747), .A2(new_n748), .A3(new_n750), .ZN(new_n751));
  AOI21_X1  g326(.A(new_n743), .B1(new_n751), .B2(G29), .ZN(new_n752));
  INV_X1    g327(.A(G2072), .ZN(new_n753));
  NAND2_X1  g328(.A1(new_n752), .A2(new_n753), .ZN(new_n754));
  INV_X1    g329(.A(KEYINPUT93), .ZN(new_n755));
  NAND2_X1  g330(.A1(new_n754), .A2(new_n755), .ZN(new_n756));
  NAND4_X1  g331(.A1(new_n732), .A2(new_n739), .A3(new_n742), .A4(new_n756), .ZN(new_n757));
  NOR2_X1   g332(.A1(new_n752), .A2(new_n753), .ZN(new_n758));
  NAND2_X1  g333(.A1(new_n758), .A2(KEYINPUT94), .ZN(new_n759));
  OAI21_X1  g334(.A(new_n759), .B1(G2078), .B2(new_n741), .ZN(new_n760));
  OAI22_X1  g335(.A1(new_n758), .A2(KEYINPUT94), .B1(new_n754), .B2(new_n755), .ZN(new_n761));
  NOR4_X1   g336(.A1(new_n725), .A2(new_n757), .A3(new_n760), .A4(new_n761), .ZN(new_n762));
  NOR2_X1   g337(.A1(G171), .A2(new_n717), .ZN(new_n763));
  AOI21_X1  g338(.A(new_n763), .B1(G5), .B2(new_n717), .ZN(new_n764));
  INV_X1    g339(.A(G1961), .ZN(new_n765));
  NOR2_X1   g340(.A1(new_n764), .A2(new_n765), .ZN(new_n766));
  XOR2_X1   g341(.A(new_n766), .B(KEYINPUT97), .Z(new_n767));
  NAND2_X1  g342(.A1(new_n764), .A2(new_n765), .ZN(new_n768));
  NAND2_X1  g343(.A1(new_n702), .A2(G32), .ZN(new_n769));
  NAND3_X1  g344(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n770));
  XOR2_X1   g345(.A(new_n770), .B(KEYINPUT26), .Z(new_n771));
  INV_X1    g346(.A(G129), .ZN(new_n772));
  OAI21_X1  g347(.A(new_n771), .B1(new_n478), .B2(new_n772), .ZN(new_n773));
  AOI22_X1  g348(.A1(new_n481), .A2(G141), .B1(G105), .B2(new_n471), .ZN(new_n774));
  INV_X1    g349(.A(new_n774), .ZN(new_n775));
  OR2_X1    g350(.A1(new_n773), .A2(new_n775), .ZN(new_n776));
  INV_X1    g351(.A(new_n776), .ZN(new_n777));
  OAI21_X1  g352(.A(new_n769), .B1(new_n777), .B2(new_n702), .ZN(new_n778));
  XNOR2_X1  g353(.A(new_n778), .B(KEYINPUT95), .ZN(new_n779));
  XNOR2_X1  g354(.A(KEYINPUT27), .B(G1996), .ZN(new_n780));
  XNOR2_X1  g355(.A(new_n779), .B(new_n780), .ZN(new_n781));
  AND4_X1   g356(.A1(new_n762), .A2(new_n767), .A3(new_n768), .A4(new_n781), .ZN(new_n782));
  AOI211_X1 g357(.A(new_n701), .B(new_n722), .C1(new_n782), .C2(KEYINPUT98), .ZN(new_n783));
  NAND2_X1  g358(.A1(new_n717), .A2(G23), .ZN(new_n784));
  INV_X1    g359(.A(G288), .ZN(new_n785));
  OAI21_X1  g360(.A(new_n784), .B1(new_n785), .B2(new_n717), .ZN(new_n786));
  XNOR2_X1  g361(.A(KEYINPUT33), .B(G1976), .ZN(new_n787));
  XNOR2_X1  g362(.A(new_n786), .B(new_n787), .ZN(new_n788));
  MUX2_X1   g363(.A(G6), .B(G305), .S(G16), .Z(new_n789));
  XNOR2_X1  g364(.A(KEYINPUT32), .B(G1981), .ZN(new_n790));
  OR2_X1    g365(.A1(new_n789), .A2(new_n790), .ZN(new_n791));
  NAND2_X1  g366(.A1(new_n789), .A2(new_n790), .ZN(new_n792));
  NAND2_X1  g367(.A1(new_n717), .A2(G22), .ZN(new_n793));
  OAI21_X1  g368(.A(new_n793), .B1(G166), .B2(new_n717), .ZN(new_n794));
  INV_X1    g369(.A(G1971), .ZN(new_n795));
  XNOR2_X1  g370(.A(new_n794), .B(new_n795), .ZN(new_n796));
  NAND4_X1  g371(.A1(new_n788), .A2(new_n791), .A3(new_n792), .A4(new_n796), .ZN(new_n797));
  OR2_X1    g372(.A1(new_n797), .A2(KEYINPUT34), .ZN(new_n798));
  NAND2_X1  g373(.A1(new_n797), .A2(KEYINPUT34), .ZN(new_n799));
  NAND2_X1  g374(.A1(new_n477), .A2(G119), .ZN(new_n800));
  XNOR2_X1  g375(.A(new_n800), .B(KEYINPUT85), .ZN(new_n801));
  OAI21_X1  g376(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n802));
  INV_X1    g377(.A(G107), .ZN(new_n803));
  AOI21_X1  g378(.A(new_n802), .B1(new_n803), .B2(G2105), .ZN(new_n804));
  AOI21_X1  g379(.A(new_n804), .B1(G131), .B2(new_n481), .ZN(new_n805));
  NAND2_X1  g380(.A1(new_n801), .A2(new_n805), .ZN(new_n806));
  MUX2_X1   g381(.A(G25), .B(new_n806), .S(G29), .Z(new_n807));
  XOR2_X1   g382(.A(KEYINPUT35), .B(G1991), .Z(new_n808));
  XOR2_X1   g383(.A(new_n807), .B(new_n808), .Z(new_n809));
  INV_X1    g384(.A(KEYINPUT86), .ZN(new_n810));
  NAND2_X1  g385(.A1(new_n809), .A2(new_n810), .ZN(new_n811));
  NOR2_X1   g386(.A1(new_n809), .A2(new_n810), .ZN(new_n812));
  NAND2_X1  g387(.A1(new_n717), .A2(G24), .ZN(new_n813));
  XOR2_X1   g388(.A(new_n813), .B(KEYINPUT87), .Z(new_n814));
  AOI21_X1  g389(.A(new_n814), .B1(G290), .B2(G16), .ZN(new_n815));
  INV_X1    g390(.A(G1986), .ZN(new_n816));
  XNOR2_X1  g391(.A(new_n815), .B(new_n816), .ZN(new_n817));
  NOR2_X1   g392(.A1(new_n812), .A2(new_n817), .ZN(new_n818));
  NAND4_X1  g393(.A1(new_n798), .A2(new_n799), .A3(new_n811), .A4(new_n818), .ZN(new_n819));
  INV_X1    g394(.A(KEYINPUT88), .ZN(new_n820));
  NAND2_X1  g395(.A1(new_n820), .A2(KEYINPUT36), .ZN(new_n821));
  OR2_X1    g396(.A1(new_n819), .A2(new_n821), .ZN(new_n822));
  OR2_X1    g397(.A1(new_n820), .A2(KEYINPUT36), .ZN(new_n823));
  NAND3_X1  g398(.A1(new_n819), .A2(new_n821), .A3(new_n823), .ZN(new_n824));
  OR2_X1    g399(.A1(new_n782), .A2(KEYINPUT98), .ZN(new_n825));
  NAND4_X1  g400(.A1(new_n783), .A2(new_n822), .A3(new_n824), .A4(new_n825), .ZN(G150));
  INV_X1    g401(.A(G150), .ZN(G311));
  INV_X1    g402(.A(G67), .ZN(new_n828));
  AOI21_X1  g403(.A(new_n828), .B1(new_n529), .B2(new_n530), .ZN(new_n829));
  AND2_X1   g404(.A1(G80), .A2(G543), .ZN(new_n830));
  OAI21_X1  g405(.A(G651), .B1(new_n829), .B2(new_n830), .ZN(new_n831));
  XNOR2_X1  g406(.A(KEYINPUT100), .B(G55), .ZN(new_n832));
  NAND2_X1  g407(.A1(new_n498), .A2(new_n832), .ZN(new_n833));
  NAND3_X1  g408(.A1(new_n501), .A2(G93), .A3(new_n502), .ZN(new_n834));
  NAND3_X1  g409(.A1(new_n831), .A2(new_n833), .A3(new_n834), .ZN(new_n835));
  INV_X1    g410(.A(KEYINPUT101), .ZN(new_n836));
  NAND2_X1  g411(.A1(new_n835), .A2(new_n836), .ZN(new_n837));
  INV_X1    g412(.A(new_n537), .ZN(new_n838));
  INV_X1    g413(.A(new_n542), .ZN(new_n839));
  NAND4_X1  g414(.A1(new_n831), .A2(new_n833), .A3(KEYINPUT101), .A4(new_n834), .ZN(new_n840));
  NAND4_X1  g415(.A1(new_n837), .A2(new_n838), .A3(new_n839), .A4(new_n840), .ZN(new_n841));
  OAI211_X1 g416(.A(new_n836), .B(new_n835), .C1(new_n537), .C2(new_n542), .ZN(new_n842));
  NAND2_X1  g417(.A1(new_n841), .A2(new_n842), .ZN(new_n843));
  XOR2_X1   g418(.A(new_n843), .B(KEYINPUT38), .Z(new_n844));
  NAND2_X1  g419(.A1(new_n602), .A2(G559), .ZN(new_n845));
  XNOR2_X1  g420(.A(new_n844), .B(new_n845), .ZN(new_n846));
  OR2_X1    g421(.A1(new_n846), .A2(KEYINPUT39), .ZN(new_n847));
  NAND2_X1  g422(.A1(new_n846), .A2(KEYINPUT39), .ZN(new_n848));
  XNOR2_X1  g423(.A(KEYINPUT102), .B(G860), .ZN(new_n849));
  NAND3_X1  g424(.A1(new_n847), .A2(new_n848), .A3(new_n849), .ZN(new_n850));
  INV_X1    g425(.A(new_n849), .ZN(new_n851));
  NAND2_X1  g426(.A1(new_n835), .A2(new_n851), .ZN(new_n852));
  XOR2_X1   g427(.A(new_n852), .B(KEYINPUT37), .Z(new_n853));
  NAND2_X1  g428(.A1(new_n850), .A2(new_n853), .ZN(G145));
  XOR2_X1   g429(.A(G160), .B(new_n626), .Z(new_n855));
  XOR2_X1   g430(.A(new_n855), .B(G162), .Z(new_n856));
  INV_X1    g431(.A(new_n856), .ZN(new_n857));
  NAND2_X1  g432(.A1(new_n713), .A2(G164), .ZN(new_n858));
  INV_X1    g433(.A(KEYINPUT91), .ZN(new_n859));
  XNOR2_X1  g434(.A(new_n712), .B(new_n859), .ZN(new_n860));
  NAND2_X1  g435(.A1(new_n490), .A2(new_n488), .ZN(new_n861));
  INV_X1    g436(.A(new_n486), .ZN(new_n862));
  NAND2_X1  g437(.A1(new_n861), .A2(new_n862), .ZN(new_n863));
  NAND2_X1  g438(.A1(new_n860), .A2(new_n863), .ZN(new_n864));
  AOI21_X1  g439(.A(new_n776), .B1(new_n858), .B2(new_n864), .ZN(new_n865));
  INV_X1    g440(.A(new_n865), .ZN(new_n866));
  INV_X1    g441(.A(new_n751), .ZN(new_n867));
  NAND3_X1  g442(.A1(new_n864), .A2(new_n858), .A3(new_n776), .ZN(new_n868));
  NAND3_X1  g443(.A1(new_n866), .A2(new_n867), .A3(new_n868), .ZN(new_n869));
  INV_X1    g444(.A(new_n868), .ZN(new_n870));
  OAI21_X1  g445(.A(new_n751), .B1(new_n870), .B2(new_n865), .ZN(new_n871));
  XNOR2_X1  g446(.A(new_n806), .B(new_n617), .ZN(new_n872));
  NAND2_X1  g447(.A1(new_n481), .A2(G142), .ZN(new_n873));
  NAND2_X1  g448(.A1(new_n477), .A2(G130), .ZN(new_n874));
  NOR2_X1   g449(.A1(new_n459), .A2(G118), .ZN(new_n875));
  OAI21_X1  g450(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n876));
  OAI211_X1 g451(.A(new_n873), .B(new_n874), .C1(new_n875), .C2(new_n876), .ZN(new_n877));
  XNOR2_X1  g452(.A(new_n872), .B(new_n877), .ZN(new_n878));
  NAND3_X1  g453(.A1(new_n869), .A2(new_n871), .A3(new_n878), .ZN(new_n879));
  INV_X1    g454(.A(KEYINPUT103), .ZN(new_n880));
  NAND2_X1  g455(.A1(new_n879), .A2(new_n880), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n869), .A2(new_n871), .ZN(new_n882));
  INV_X1    g457(.A(new_n878), .ZN(new_n883));
  NAND2_X1  g458(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  NAND2_X1  g459(.A1(new_n881), .A2(new_n884), .ZN(new_n885));
  NAND3_X1  g460(.A1(new_n882), .A2(new_n880), .A3(new_n883), .ZN(new_n886));
  AOI21_X1  g461(.A(new_n857), .B1(new_n885), .B2(new_n886), .ZN(new_n887));
  INV_X1    g462(.A(new_n887), .ZN(new_n888));
  AND2_X1   g463(.A1(new_n879), .A2(new_n857), .ZN(new_n889));
  AOI21_X1  g464(.A(G37), .B1(new_n889), .B2(new_n884), .ZN(new_n890));
  AOI21_X1  g465(.A(KEYINPUT40), .B1(new_n888), .B2(new_n890), .ZN(new_n891));
  INV_X1    g466(.A(new_n890), .ZN(new_n892));
  INV_X1    g467(.A(KEYINPUT40), .ZN(new_n893));
  NOR3_X1   g468(.A1(new_n892), .A2(new_n887), .A3(new_n893), .ZN(new_n894));
  NOR2_X1   g469(.A1(new_n891), .A2(new_n894), .ZN(G395));
  NAND2_X1  g470(.A1(new_n835), .A2(new_n589), .ZN(new_n896));
  AND2_X1   g471(.A1(new_n587), .A2(G305), .ZN(new_n897));
  NOR2_X1   g472(.A1(new_n587), .A2(G305), .ZN(new_n898));
  NOR2_X1   g473(.A1(new_n897), .A2(new_n898), .ZN(new_n899));
  XNOR2_X1  g474(.A(G166), .B(G288), .ZN(new_n900));
  XNOR2_X1  g475(.A(new_n899), .B(new_n900), .ZN(new_n901));
  XNOR2_X1  g476(.A(new_n901), .B(KEYINPUT42), .ZN(new_n902));
  XNOR2_X1  g477(.A(new_n843), .B(new_n613), .ZN(new_n903));
  AOI22_X1  g478(.A1(new_n594), .A2(new_n595), .B1(G54), .B2(new_n498), .ZN(new_n904));
  AOI21_X1  g479(.A(G299), .B1(new_n600), .B2(new_n904), .ZN(new_n905));
  INV_X1    g480(.A(KEYINPUT104), .ZN(new_n906));
  AND3_X1   g481(.A1(new_n556), .A2(new_n563), .A3(new_n564), .ZN(new_n907));
  OAI21_X1  g482(.A(new_n906), .B1(new_n907), .B2(new_n612), .ZN(new_n908));
  NAND3_X1  g483(.A1(new_n602), .A2(KEYINPUT104), .A3(G299), .ZN(new_n909));
  AOI21_X1  g484(.A(new_n905), .B1(new_n908), .B2(new_n909), .ZN(new_n910));
  NOR2_X1   g485(.A1(new_n903), .A2(new_n910), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n908), .A2(new_n909), .ZN(new_n912));
  OAI21_X1  g487(.A(KEYINPUT41), .B1(new_n602), .B2(G299), .ZN(new_n913));
  INV_X1    g488(.A(new_n913), .ZN(new_n914));
  NAND2_X1  g489(.A1(new_n912), .A2(new_n914), .ZN(new_n915));
  INV_X1    g490(.A(KEYINPUT105), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n915), .A2(new_n916), .ZN(new_n917));
  NOR3_X1   g492(.A1(new_n907), .A2(new_n906), .A3(new_n612), .ZN(new_n918));
  AOI21_X1  g493(.A(KEYINPUT104), .B1(new_n602), .B2(G299), .ZN(new_n919));
  OAI22_X1  g494(.A1(new_n918), .A2(new_n919), .B1(G299), .B2(new_n602), .ZN(new_n920));
  INV_X1    g495(.A(KEYINPUT41), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n920), .A2(new_n921), .ZN(new_n922));
  AOI21_X1  g497(.A(new_n913), .B1(new_n908), .B2(new_n909), .ZN(new_n923));
  NAND2_X1  g498(.A1(new_n923), .A2(KEYINPUT105), .ZN(new_n924));
  NAND3_X1  g499(.A1(new_n917), .A2(new_n922), .A3(new_n924), .ZN(new_n925));
  AOI21_X1  g500(.A(new_n911), .B1(new_n925), .B2(new_n903), .ZN(new_n926));
  XNOR2_X1  g501(.A(new_n902), .B(new_n926), .ZN(new_n927));
  OAI21_X1  g502(.A(new_n896), .B1(new_n927), .B2(new_n589), .ZN(G295));
  OAI21_X1  g503(.A(new_n896), .B1(new_n927), .B2(new_n589), .ZN(G331));
  INV_X1    g504(.A(KEYINPUT44), .ZN(new_n930));
  INV_X1    g505(.A(KEYINPUT107), .ZN(new_n931));
  INV_X1    g506(.A(KEYINPUT106), .ZN(new_n932));
  AND3_X1   g507(.A1(new_n841), .A2(G168), .A3(new_n842), .ZN(new_n933));
  AOI21_X1  g508(.A(G168), .B1(new_n841), .B2(new_n842), .ZN(new_n934));
  OAI21_X1  g509(.A(G301), .B1(new_n933), .B2(new_n934), .ZN(new_n935));
  NAND2_X1  g510(.A1(new_n843), .A2(G286), .ZN(new_n936));
  NAND3_X1  g511(.A1(new_n841), .A2(G168), .A3(new_n842), .ZN(new_n937));
  NAND3_X1  g512(.A1(new_n936), .A2(G171), .A3(new_n937), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n935), .A2(new_n938), .ZN(new_n939));
  OAI22_X1  g514(.A1(new_n923), .A2(KEYINPUT105), .B1(new_n910), .B2(KEYINPUT41), .ZN(new_n940));
  AND3_X1   g515(.A1(new_n912), .A2(new_n914), .A3(KEYINPUT105), .ZN(new_n941));
  OAI211_X1 g516(.A(new_n932), .B(new_n939), .C1(new_n940), .C2(new_n941), .ZN(new_n942));
  NAND3_X1  g517(.A1(new_n935), .A2(new_n938), .A3(new_n920), .ZN(new_n943));
  NAND2_X1  g518(.A1(new_n942), .A2(new_n943), .ZN(new_n944));
  AOI21_X1  g519(.A(new_n932), .B1(new_n925), .B2(new_n939), .ZN(new_n945));
  NOR3_X1   g520(.A1(new_n944), .A2(new_n945), .A3(new_n901), .ZN(new_n946));
  AOI22_X1  g521(.A1(new_n922), .A2(new_n915), .B1(new_n935), .B2(new_n938), .ZN(new_n947));
  INV_X1    g522(.A(new_n943), .ZN(new_n948));
  OAI21_X1  g523(.A(new_n901), .B1(new_n947), .B2(new_n948), .ZN(new_n949));
  INV_X1    g524(.A(KEYINPUT43), .ZN(new_n950));
  INV_X1    g525(.A(G37), .ZN(new_n951));
  NAND3_X1  g526(.A1(new_n949), .A2(new_n950), .A3(new_n951), .ZN(new_n952));
  OAI21_X1  g527(.A(new_n931), .B1(new_n946), .B2(new_n952), .ZN(new_n953));
  XOR2_X1   g528(.A(new_n899), .B(new_n900), .Z(new_n954));
  OAI21_X1  g529(.A(new_n915), .B1(KEYINPUT41), .B2(new_n910), .ZN(new_n955));
  NAND2_X1  g530(.A1(new_n939), .A2(new_n955), .ZN(new_n956));
  AOI21_X1  g531(.A(new_n954), .B1(new_n956), .B2(new_n943), .ZN(new_n957));
  NOR3_X1   g532(.A1(new_n957), .A2(KEYINPUT43), .A3(G37), .ZN(new_n958));
  OAI21_X1  g533(.A(new_n939), .B1(new_n940), .B2(new_n941), .ZN(new_n959));
  NAND2_X1  g534(.A1(new_n959), .A2(KEYINPUT106), .ZN(new_n960));
  NAND4_X1  g535(.A1(new_n960), .A2(new_n954), .A3(new_n943), .A4(new_n942), .ZN(new_n961));
  NAND3_X1  g536(.A1(new_n958), .A2(KEYINPUT107), .A3(new_n961), .ZN(new_n962));
  NAND2_X1  g537(.A1(new_n953), .A2(new_n962), .ZN(new_n963));
  NAND3_X1  g538(.A1(new_n960), .A2(new_n943), .A3(new_n942), .ZN(new_n964));
  AOI21_X1  g539(.A(G37), .B1(new_n964), .B2(new_n901), .ZN(new_n965));
  AOI21_X1  g540(.A(new_n950), .B1(new_n965), .B2(new_n961), .ZN(new_n966));
  OAI21_X1  g541(.A(new_n930), .B1(new_n963), .B2(new_n966), .ZN(new_n967));
  NAND2_X1  g542(.A1(new_n967), .A2(KEYINPUT108), .ZN(new_n968));
  NAND2_X1  g543(.A1(new_n949), .A2(new_n951), .ZN(new_n969));
  OAI21_X1  g544(.A(KEYINPUT43), .B1(new_n946), .B2(new_n969), .ZN(new_n970));
  OAI21_X1  g545(.A(new_n901), .B1(new_n944), .B2(new_n945), .ZN(new_n971));
  NAND4_X1  g546(.A1(new_n971), .A2(new_n961), .A3(new_n950), .A4(new_n951), .ZN(new_n972));
  NAND3_X1  g547(.A1(new_n970), .A2(new_n972), .A3(KEYINPUT44), .ZN(new_n973));
  NAND2_X1  g548(.A1(new_n973), .A2(KEYINPUT109), .ZN(new_n974));
  INV_X1    g549(.A(KEYINPUT109), .ZN(new_n975));
  NAND4_X1  g550(.A1(new_n970), .A2(new_n972), .A3(new_n975), .A4(KEYINPUT44), .ZN(new_n976));
  NAND2_X1  g551(.A1(new_n974), .A2(new_n976), .ZN(new_n977));
  INV_X1    g552(.A(KEYINPUT108), .ZN(new_n978));
  OAI211_X1 g553(.A(new_n978), .B(new_n930), .C1(new_n963), .C2(new_n966), .ZN(new_n979));
  NAND3_X1  g554(.A1(new_n968), .A2(new_n977), .A3(new_n979), .ZN(G397));
  AOI21_X1  g555(.A(G1384), .B1(new_n861), .B2(new_n862), .ZN(new_n981));
  AND2_X1   g556(.A1(new_n981), .A2(KEYINPUT110), .ZN(new_n982));
  INV_X1    g557(.A(KEYINPUT45), .ZN(new_n983));
  OAI21_X1  g558(.A(new_n983), .B1(new_n981), .B2(KEYINPUT110), .ZN(new_n984));
  NOR2_X1   g559(.A1(new_n982), .A2(new_n984), .ZN(new_n985));
  INV_X1    g560(.A(G40), .ZN(new_n986));
  NOR3_X1   g561(.A1(new_n467), .A2(new_n473), .A3(new_n986), .ZN(new_n987));
  NAND2_X1  g562(.A1(new_n985), .A2(new_n987), .ZN(new_n988));
  INV_X1    g563(.A(new_n988), .ZN(new_n989));
  INV_X1    g564(.A(G1996), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n989), .A2(new_n990), .ZN(new_n991));
  XNOR2_X1  g566(.A(new_n991), .B(KEYINPUT46), .ZN(new_n992));
  XNOR2_X1  g567(.A(new_n713), .B(G2067), .ZN(new_n993));
  NAND2_X1  g568(.A1(new_n993), .A2(new_n777), .ZN(new_n994));
  NAND2_X1  g569(.A1(new_n994), .A2(new_n989), .ZN(new_n995));
  NAND2_X1  g570(.A1(new_n992), .A2(new_n995), .ZN(new_n996));
  INV_X1    g571(.A(KEYINPUT47), .ZN(new_n997));
  NAND2_X1  g572(.A1(new_n996), .A2(new_n997), .ZN(new_n998));
  NAND3_X1  g573(.A1(new_n992), .A2(KEYINPUT47), .A3(new_n995), .ZN(new_n999));
  NAND2_X1  g574(.A1(new_n998), .A2(new_n999), .ZN(new_n1000));
  OR2_X1    g575(.A1(new_n1000), .A2(KEYINPUT127), .ZN(new_n1001));
  NAND2_X1  g576(.A1(new_n1000), .A2(KEYINPUT127), .ZN(new_n1002));
  XNOR2_X1  g577(.A(new_n776), .B(new_n990), .ZN(new_n1003));
  AND2_X1   g578(.A1(new_n993), .A2(new_n1003), .ZN(new_n1004));
  NAND4_X1  g579(.A1(new_n1004), .A2(new_n808), .A3(new_n801), .A4(new_n805), .ZN(new_n1005));
  NAND2_X1  g580(.A1(new_n713), .A2(new_n715), .ZN(new_n1006));
  AOI21_X1  g581(.A(new_n988), .B1(new_n1005), .B2(new_n1006), .ZN(new_n1007));
  XNOR2_X1  g582(.A(new_n806), .B(new_n808), .ZN(new_n1008));
  AOI21_X1  g583(.A(new_n988), .B1(new_n1004), .B2(new_n1008), .ZN(new_n1009));
  NOR3_X1   g584(.A1(new_n988), .A2(G1986), .A3(G290), .ZN(new_n1010));
  NOR2_X1   g585(.A1(new_n1010), .A2(KEYINPUT48), .ZN(new_n1011));
  NOR2_X1   g586(.A1(new_n1009), .A2(new_n1011), .ZN(new_n1012));
  NAND2_X1  g587(.A1(new_n1010), .A2(KEYINPUT48), .ZN(new_n1013));
  AOI21_X1  g588(.A(new_n1007), .B1(new_n1012), .B2(new_n1013), .ZN(new_n1014));
  AND3_X1   g589(.A1(new_n1001), .A2(new_n1002), .A3(new_n1014), .ZN(new_n1015));
  INV_X1    g590(.A(KEYINPUT61), .ZN(new_n1016));
  XNOR2_X1  g591(.A(G299), .B(KEYINPUT57), .ZN(new_n1017));
  INV_X1    g592(.A(new_n1017), .ZN(new_n1018));
  INV_X1    g593(.A(KEYINPUT50), .ZN(new_n1019));
  INV_X1    g594(.A(G1384), .ZN(new_n1020));
  NAND3_X1  g595(.A1(new_n863), .A2(new_n1019), .A3(new_n1020), .ZN(new_n1021));
  OAI21_X1  g596(.A(KEYINPUT50), .B1(G164), .B2(G1384), .ZN(new_n1022));
  NAND3_X1  g597(.A1(new_n1021), .A2(new_n1022), .A3(new_n987), .ZN(new_n1023));
  INV_X1    g598(.A(G1956), .ZN(new_n1024));
  NAND2_X1  g599(.A1(new_n1023), .A2(new_n1024), .ZN(new_n1025));
  INV_X1    g600(.A(KEYINPUT120), .ZN(new_n1026));
  NAND2_X1  g601(.A1(new_n1025), .A2(new_n1026), .ZN(new_n1027));
  NAND3_X1  g602(.A1(new_n1023), .A2(KEYINPUT120), .A3(new_n1024), .ZN(new_n1028));
  NAND2_X1  g603(.A1(new_n1027), .A2(new_n1028), .ZN(new_n1029));
  OAI21_X1  g604(.A(new_n983), .B1(G164), .B2(G1384), .ZN(new_n1030));
  NOR2_X1   g605(.A1(new_n983), .A2(G1384), .ZN(new_n1031));
  NAND2_X1  g606(.A1(new_n863), .A2(new_n1031), .ZN(new_n1032));
  NAND3_X1  g607(.A1(new_n1030), .A2(new_n987), .A3(new_n1032), .ZN(new_n1033));
  XNOR2_X1  g608(.A(KEYINPUT56), .B(G2072), .ZN(new_n1034));
  INV_X1    g609(.A(new_n1034), .ZN(new_n1035));
  NOR2_X1   g610(.A1(new_n1033), .A2(new_n1035), .ZN(new_n1036));
  INV_X1    g611(.A(new_n1036), .ZN(new_n1037));
  AOI21_X1  g612(.A(new_n1018), .B1(new_n1029), .B2(new_n1037), .ZN(new_n1038));
  AOI211_X1 g613(.A(new_n1017), .B(new_n1036), .C1(new_n1027), .C2(new_n1028), .ZN(new_n1039));
  OAI21_X1  g614(.A(new_n1016), .B1(new_n1038), .B2(new_n1039), .ZN(new_n1040));
  INV_X1    g615(.A(KEYINPUT60), .ZN(new_n1041));
  AND2_X1   g616(.A1(new_n1023), .A2(new_n699), .ZN(new_n1042));
  NAND2_X1  g617(.A1(new_n981), .A2(new_n987), .ZN(new_n1043));
  NOR2_X1   g618(.A1(new_n1043), .A2(G2067), .ZN(new_n1044));
  OAI21_X1  g619(.A(new_n602), .B1(new_n1042), .B2(new_n1044), .ZN(new_n1045));
  AOI21_X1  g620(.A(new_n1044), .B1(new_n699), .B2(new_n1023), .ZN(new_n1046));
  NAND2_X1  g621(.A1(new_n1046), .A2(new_n612), .ZN(new_n1047));
  AOI21_X1  g622(.A(new_n1041), .B1(new_n1045), .B2(new_n1047), .ZN(new_n1048));
  NAND3_X1  g623(.A1(new_n1046), .A2(new_n1041), .A3(new_n602), .ZN(new_n1049));
  INV_X1    g624(.A(KEYINPUT59), .ZN(new_n1050));
  NAND4_X1  g625(.A1(new_n1030), .A2(new_n1032), .A3(new_n990), .A4(new_n987), .ZN(new_n1051));
  XOR2_X1   g626(.A(KEYINPUT58), .B(G1341), .Z(new_n1052));
  NAND2_X1  g627(.A1(new_n1043), .A2(new_n1052), .ZN(new_n1053));
  NAND2_X1  g628(.A1(new_n1051), .A2(new_n1053), .ZN(new_n1054));
  AOI21_X1  g629(.A(new_n1050), .B1(new_n1054), .B2(new_n543), .ZN(new_n1055));
  AOI211_X1 g630(.A(KEYINPUT59), .B(new_n610), .C1(new_n1051), .C2(new_n1053), .ZN(new_n1056));
  OAI21_X1  g631(.A(new_n1049), .B1(new_n1055), .B2(new_n1056), .ZN(new_n1057));
  NOR2_X1   g632(.A1(new_n1048), .A2(new_n1057), .ZN(new_n1058));
  INV_X1    g633(.A(new_n1028), .ZN(new_n1059));
  AOI21_X1  g634(.A(KEYINPUT120), .B1(new_n1023), .B2(new_n1024), .ZN(new_n1060));
  OAI21_X1  g635(.A(new_n1037), .B1(new_n1059), .B2(new_n1060), .ZN(new_n1061));
  NAND2_X1  g636(.A1(new_n1061), .A2(new_n1017), .ZN(new_n1062));
  OAI211_X1 g637(.A(new_n1018), .B(new_n1037), .C1(new_n1059), .C2(new_n1060), .ZN(new_n1063));
  NAND3_X1  g638(.A1(new_n1062), .A2(KEYINPUT61), .A3(new_n1063), .ZN(new_n1064));
  NAND3_X1  g639(.A1(new_n1040), .A2(new_n1058), .A3(new_n1064), .ZN(new_n1065));
  INV_X1    g640(.A(new_n1045), .ZN(new_n1066));
  NAND2_X1  g641(.A1(new_n1066), .A2(new_n1063), .ZN(new_n1067));
  NAND3_X1  g642(.A1(new_n1067), .A2(KEYINPUT121), .A3(new_n1062), .ZN(new_n1068));
  NAND2_X1  g643(.A1(new_n1067), .A2(new_n1062), .ZN(new_n1069));
  INV_X1    g644(.A(KEYINPUT121), .ZN(new_n1070));
  NAND2_X1  g645(.A1(new_n1069), .A2(new_n1070), .ZN(new_n1071));
  NAND3_X1  g646(.A1(new_n1065), .A2(new_n1068), .A3(new_n1071), .ZN(new_n1072));
  INV_X1    g647(.A(KEYINPUT119), .ZN(new_n1073));
  INV_X1    g648(.A(G1966), .ZN(new_n1074));
  NOR2_X1   g649(.A1(new_n981), .A2(KEYINPUT45), .ZN(new_n1075));
  INV_X1    g650(.A(new_n1031), .ZN(new_n1076));
  OAI21_X1  g651(.A(new_n987), .B1(G164), .B2(new_n1076), .ZN(new_n1077));
  OAI211_X1 g652(.A(new_n1073), .B(new_n1074), .C1(new_n1075), .C2(new_n1077), .ZN(new_n1078));
  NAND4_X1  g653(.A1(new_n1021), .A2(new_n1022), .A3(new_n738), .A4(new_n987), .ZN(new_n1079));
  NAND2_X1  g654(.A1(new_n1078), .A2(new_n1079), .ZN(new_n1080));
  AOI21_X1  g655(.A(new_n1073), .B1(new_n1033), .B2(new_n1074), .ZN(new_n1081));
  OAI21_X1  g656(.A(KEYINPUT122), .B1(new_n1080), .B2(new_n1081), .ZN(new_n1082));
  NAND2_X1  g657(.A1(new_n1033), .A2(new_n1074), .ZN(new_n1083));
  NAND2_X1  g658(.A1(new_n1083), .A2(KEYINPUT119), .ZN(new_n1084));
  INV_X1    g659(.A(KEYINPUT122), .ZN(new_n1085));
  NAND4_X1  g660(.A1(new_n1084), .A2(new_n1085), .A3(new_n1079), .A4(new_n1078), .ZN(new_n1086));
  AOI21_X1  g661(.A(G286), .B1(new_n1082), .B2(new_n1086), .ZN(new_n1087));
  INV_X1    g662(.A(KEYINPUT51), .ZN(new_n1088));
  INV_X1    g663(.A(G8), .ZN(new_n1089));
  NOR2_X1   g664(.A1(new_n1088), .A2(new_n1089), .ZN(new_n1090));
  INV_X1    g665(.A(new_n1090), .ZN(new_n1091));
  NAND3_X1  g666(.A1(new_n1084), .A2(new_n1079), .A3(new_n1078), .ZN(new_n1092));
  AND2_X1   g667(.A1(new_n1092), .A2(G8), .ZN(new_n1093));
  OAI21_X1  g668(.A(new_n1088), .B1(G168), .B2(new_n1089), .ZN(new_n1094));
  OAI22_X1  g669(.A1(new_n1087), .A2(new_n1091), .B1(new_n1093), .B2(new_n1094), .ZN(new_n1095));
  NOR2_X1   g670(.A1(G168), .A2(new_n1089), .ZN(new_n1096));
  NAND3_X1  g671(.A1(new_n1082), .A2(new_n1086), .A3(new_n1096), .ZN(new_n1097));
  INV_X1    g672(.A(KEYINPUT123), .ZN(new_n1098));
  NAND2_X1  g673(.A1(new_n1097), .A2(new_n1098), .ZN(new_n1099));
  NAND4_X1  g674(.A1(new_n1082), .A2(new_n1086), .A3(KEYINPUT123), .A4(new_n1096), .ZN(new_n1100));
  NAND3_X1  g675(.A1(new_n1095), .A2(new_n1099), .A3(new_n1100), .ZN(new_n1101));
  INV_X1    g676(.A(KEYINPUT53), .ZN(new_n1102));
  OAI21_X1  g677(.A(new_n1102), .B1(new_n1033), .B2(G2078), .ZN(new_n1103));
  NAND2_X1  g678(.A1(new_n1023), .A2(new_n765), .ZN(new_n1104));
  NOR2_X1   g679(.A1(new_n1102), .A2(G2078), .ZN(new_n1105));
  NAND4_X1  g680(.A1(new_n1030), .A2(new_n1032), .A3(new_n987), .A4(new_n1105), .ZN(new_n1106));
  AND3_X1   g681(.A1(new_n1104), .A2(KEYINPUT124), .A3(new_n1106), .ZN(new_n1107));
  AOI21_X1  g682(.A(KEYINPUT124), .B1(new_n1104), .B2(new_n1106), .ZN(new_n1108));
  OAI211_X1 g683(.A(G301), .B(new_n1103), .C1(new_n1107), .C2(new_n1108), .ZN(new_n1109));
  INV_X1    g684(.A(KEYINPUT54), .ZN(new_n1110));
  INV_X1    g685(.A(new_n473), .ZN(new_n1111));
  AND2_X1   g686(.A1(new_n1111), .A2(KEYINPUT125), .ZN(new_n1112));
  NOR2_X1   g687(.A1(new_n1111), .A2(KEYINPUT125), .ZN(new_n1113));
  NAND2_X1  g688(.A1(new_n1105), .A2(G40), .ZN(new_n1114));
  NOR4_X1   g689(.A1(new_n1112), .A2(new_n1113), .A3(new_n467), .A4(new_n1114), .ZN(new_n1115));
  NAND2_X1  g690(.A1(new_n1115), .A2(new_n1032), .ZN(new_n1116));
  OAI211_X1 g691(.A(new_n1103), .B(new_n1104), .C1(new_n985), .C2(new_n1116), .ZN(new_n1117));
  AOI21_X1  g692(.A(new_n1110), .B1(new_n1117), .B2(G171), .ZN(new_n1118));
  NAND2_X1  g693(.A1(new_n1109), .A2(new_n1118), .ZN(new_n1119));
  INV_X1    g694(.A(KEYINPUT115), .ZN(new_n1120));
  AOI21_X1  g695(.A(new_n1120), .B1(new_n1043), .B2(G8), .ZN(new_n1121));
  AOI211_X1 g696(.A(KEYINPUT115), .B(new_n1089), .C1(new_n981), .C2(new_n987), .ZN(new_n1122));
  OR2_X1    g697(.A1(new_n1121), .A2(new_n1122), .ZN(new_n1123));
  XNOR2_X1  g698(.A(KEYINPUT116), .B(G86), .ZN(new_n1124));
  NAND2_X1  g699(.A1(new_n521), .A2(new_n1124), .ZN(new_n1125));
  NAND3_X1  g700(.A1(new_n578), .A2(new_n580), .A3(new_n1125), .ZN(new_n1126));
  NAND2_X1  g701(.A1(new_n1126), .A2(G1981), .ZN(new_n1127));
  INV_X1    g702(.A(G1981), .ZN(new_n1128));
  NAND4_X1  g703(.A1(new_n578), .A2(new_n1128), .A3(new_n579), .A4(new_n580), .ZN(new_n1129));
  NAND3_X1  g704(.A1(new_n1127), .A2(KEYINPUT117), .A3(new_n1129), .ZN(new_n1130));
  AOI21_X1  g705(.A(KEYINPUT49), .B1(new_n1130), .B2(KEYINPUT118), .ZN(new_n1131));
  NAND2_X1  g706(.A1(KEYINPUT118), .A2(KEYINPUT49), .ZN(new_n1132));
  AOI22_X1  g707(.A1(new_n1127), .A2(new_n1129), .B1(KEYINPUT117), .B2(new_n1132), .ZN(new_n1133));
  OAI21_X1  g708(.A(new_n1123), .B1(new_n1131), .B2(new_n1133), .ZN(new_n1134));
  NAND2_X1  g709(.A1(new_n785), .A2(G1976), .ZN(new_n1135));
  INV_X1    g710(.A(G1976), .ZN(new_n1136));
  AOI21_X1  g711(.A(KEYINPUT52), .B1(G288), .B2(new_n1136), .ZN(new_n1137));
  NAND3_X1  g712(.A1(new_n1123), .A2(new_n1135), .A3(new_n1137), .ZN(new_n1138));
  OAI21_X1  g713(.A(new_n1135), .B1(new_n1121), .B2(new_n1122), .ZN(new_n1139));
  NAND2_X1  g714(.A1(new_n1139), .A2(KEYINPUT52), .ZN(new_n1140));
  AND3_X1   g715(.A1(new_n1134), .A2(new_n1138), .A3(new_n1140), .ZN(new_n1141));
  NOR2_X1   g716(.A1(new_n1023), .A2(G2090), .ZN(new_n1142));
  NAND2_X1  g717(.A1(new_n1142), .A2(KEYINPUT113), .ZN(new_n1143));
  INV_X1    g718(.A(new_n1033), .ZN(new_n1144));
  OAI21_X1  g719(.A(KEYINPUT112), .B1(new_n1144), .B2(G1971), .ZN(new_n1145));
  INV_X1    g720(.A(KEYINPUT113), .ZN(new_n1146));
  OAI21_X1  g721(.A(new_n1146), .B1(new_n1023), .B2(G2090), .ZN(new_n1147));
  INV_X1    g722(.A(KEYINPUT112), .ZN(new_n1148));
  NAND3_X1  g723(.A1(new_n1033), .A2(new_n1148), .A3(new_n795), .ZN(new_n1149));
  NAND4_X1  g724(.A1(new_n1143), .A2(new_n1145), .A3(new_n1147), .A4(new_n1149), .ZN(new_n1150));
  NOR2_X1   g725(.A1(G166), .A2(new_n1089), .ZN(new_n1151));
  XNOR2_X1  g726(.A(KEYINPUT114), .B(KEYINPUT55), .ZN(new_n1152));
  NOR2_X1   g727(.A1(new_n1151), .A2(new_n1152), .ZN(new_n1153));
  INV_X1    g728(.A(KEYINPUT114), .ZN(new_n1154));
  NOR2_X1   g729(.A1(new_n1154), .A2(KEYINPUT55), .ZN(new_n1155));
  INV_X1    g730(.A(new_n1155), .ZN(new_n1156));
  AOI21_X1  g731(.A(new_n1153), .B1(new_n1151), .B2(new_n1156), .ZN(new_n1157));
  INV_X1    g732(.A(new_n1157), .ZN(new_n1158));
  NAND3_X1  g733(.A1(new_n1150), .A2(G8), .A3(new_n1158), .ZN(new_n1159));
  NOR2_X1   g734(.A1(new_n1144), .A2(G1971), .ZN(new_n1160));
  OAI21_X1  g735(.A(G8), .B1(new_n1160), .B2(new_n1142), .ZN(new_n1161));
  NAND2_X1  g736(.A1(new_n1161), .A2(new_n1157), .ZN(new_n1162));
  NAND4_X1  g737(.A1(new_n1119), .A2(new_n1141), .A3(new_n1159), .A4(new_n1162), .ZN(new_n1163));
  OAI21_X1  g738(.A(new_n1103), .B1(new_n1107), .B2(new_n1108), .ZN(new_n1164));
  NAND2_X1  g739(.A1(new_n1164), .A2(G171), .ZN(new_n1165));
  OR2_X1    g740(.A1(new_n1117), .A2(G171), .ZN(new_n1166));
  AOI21_X1  g741(.A(KEYINPUT54), .B1(new_n1165), .B2(new_n1166), .ZN(new_n1167));
  NOR2_X1   g742(.A1(new_n1163), .A2(new_n1167), .ZN(new_n1168));
  NAND3_X1  g743(.A1(new_n1072), .A2(new_n1101), .A3(new_n1168), .ZN(new_n1169));
  AOI21_X1  g744(.A(new_n1094), .B1(new_n1092), .B2(G8), .ZN(new_n1170));
  NAND2_X1  g745(.A1(new_n1082), .A2(new_n1086), .ZN(new_n1171));
  NAND2_X1  g746(.A1(new_n1171), .A2(G168), .ZN(new_n1172));
  AOI21_X1  g747(.A(new_n1170), .B1(new_n1172), .B2(new_n1090), .ZN(new_n1173));
  NAND2_X1  g748(.A1(new_n1099), .A2(new_n1100), .ZN(new_n1174));
  OAI21_X1  g749(.A(KEYINPUT62), .B1(new_n1173), .B2(new_n1174), .ZN(new_n1175));
  INV_X1    g750(.A(KEYINPUT62), .ZN(new_n1176));
  NAND4_X1  g751(.A1(new_n1095), .A2(new_n1176), .A3(new_n1099), .A4(new_n1100), .ZN(new_n1177));
  NAND2_X1  g752(.A1(new_n1159), .A2(new_n1162), .ZN(new_n1178));
  NAND3_X1  g753(.A1(new_n1134), .A2(new_n1138), .A3(new_n1140), .ZN(new_n1179));
  NOR3_X1   g754(.A1(new_n1178), .A2(new_n1179), .A3(new_n1165), .ZN(new_n1180));
  NAND3_X1  g755(.A1(new_n1175), .A2(new_n1177), .A3(new_n1180), .ZN(new_n1181));
  INV_X1    g756(.A(new_n1129), .ZN(new_n1182));
  NOR2_X1   g757(.A1(new_n1131), .A2(new_n1133), .ZN(new_n1183));
  NOR2_X1   g758(.A1(G288), .A2(G1976), .ZN(new_n1184));
  AOI21_X1  g759(.A(new_n1182), .B1(new_n1183), .B2(new_n1184), .ZN(new_n1185));
  INV_X1    g760(.A(new_n1123), .ZN(new_n1186));
  OAI22_X1  g761(.A1(new_n1159), .A2(new_n1179), .B1(new_n1185), .B2(new_n1186), .ZN(new_n1187));
  NAND2_X1  g762(.A1(new_n1150), .A2(G8), .ZN(new_n1188));
  AOI21_X1  g763(.A(new_n1179), .B1(new_n1157), .B2(new_n1188), .ZN(new_n1189));
  NAND3_X1  g764(.A1(new_n1092), .A2(G8), .A3(G168), .ZN(new_n1190));
  INV_X1    g765(.A(new_n1190), .ZN(new_n1191));
  NAND4_X1  g766(.A1(new_n1189), .A2(KEYINPUT63), .A3(new_n1159), .A4(new_n1191), .ZN(new_n1192));
  NAND4_X1  g767(.A1(new_n1141), .A2(new_n1191), .A3(new_n1159), .A4(new_n1162), .ZN(new_n1193));
  INV_X1    g768(.A(KEYINPUT63), .ZN(new_n1194));
  NAND2_X1  g769(.A1(new_n1193), .A2(new_n1194), .ZN(new_n1195));
  AOI21_X1  g770(.A(new_n1187), .B1(new_n1192), .B2(new_n1195), .ZN(new_n1196));
  NAND3_X1  g771(.A1(new_n1169), .A2(new_n1181), .A3(new_n1196), .ZN(new_n1197));
  INV_X1    g772(.A(KEYINPUT126), .ZN(new_n1198));
  NOR3_X1   g773(.A1(new_n988), .A2(new_n816), .A3(new_n587), .ZN(new_n1199));
  NOR2_X1   g774(.A1(new_n1199), .A2(new_n1010), .ZN(new_n1200));
  XNOR2_X1  g775(.A(new_n1200), .B(KEYINPUT111), .ZN(new_n1201));
  NOR2_X1   g776(.A1(new_n1201), .A2(new_n1009), .ZN(new_n1202));
  AND3_X1   g777(.A1(new_n1197), .A2(new_n1198), .A3(new_n1202), .ZN(new_n1203));
  AOI21_X1  g778(.A(new_n1198), .B1(new_n1197), .B2(new_n1202), .ZN(new_n1204));
  OAI21_X1  g779(.A(new_n1015), .B1(new_n1203), .B2(new_n1204), .ZN(G329));
  assign    G231 = 1'b0;
  OAI21_X1  g780(.A(G319), .B1(new_n645), .B2(new_n646), .ZN(new_n1207));
  NOR3_X1   g781(.A1(G229), .A2(G227), .A3(new_n1207), .ZN(new_n1208));
  OAI21_X1  g782(.A(new_n1208), .B1(new_n892), .B2(new_n887), .ZN(new_n1209));
  NOR2_X1   g783(.A1(new_n963), .A2(new_n966), .ZN(new_n1210));
  NOR2_X1   g784(.A1(new_n1209), .A2(new_n1210), .ZN(G308));
  OR2_X1    g785(.A1(new_n1209), .A2(new_n1210), .ZN(G225));
endmodule


