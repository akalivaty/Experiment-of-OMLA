//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 1 1 0 1 0 1 0 1 0 1 0 1 0 1 1 0 0 1 0 0 1 1 1 0 1 0 0 0 1 1 1 0 0 1 1 1 1 0 0 1 0 0 0 1 0 0 1 1 1 0 1 1 1 1 1 1 0 1 0 1 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:21:45 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n619, new_n620, new_n621, new_n622,
    new_n623, new_n624, new_n626, new_n627, new_n628, new_n629, new_n630,
    new_n631, new_n632, new_n633, new_n634, new_n636, new_n637, new_n638,
    new_n639, new_n640, new_n641, new_n642, new_n643, new_n644, new_n645,
    new_n646, new_n647, new_n648, new_n649, new_n650, new_n651, new_n652,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n671, new_n672, new_n673, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n689, new_n691, new_n692,
    new_n693, new_n695, new_n696, new_n697, new_n698, new_n699, new_n700,
    new_n701, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n744, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n773, new_n774, new_n775,
    new_n776, new_n777, new_n778, new_n779, new_n780, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n914, new_n915, new_n916, new_n917, new_n918, new_n920,
    new_n921, new_n922, new_n923, new_n924, new_n925, new_n926, new_n927,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n937, new_n938, new_n939, new_n940, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n963, new_n964, new_n965, new_n966,
    new_n967, new_n968, new_n969, new_n970, new_n971, new_n972, new_n973;
  XNOR2_X1  g000(.A(G110), .B(G140), .ZN(new_n187));
  INV_X1    g001(.A(G227), .ZN(new_n188));
  NOR2_X1   g002(.A1(new_n188), .A2(G953), .ZN(new_n189));
  XOR2_X1   g003(.A(new_n187), .B(new_n189), .Z(new_n190));
  INV_X1    g004(.A(new_n190), .ZN(new_n191));
  XOR2_X1   g005(.A(KEYINPUT68), .B(G131), .Z(new_n192));
  INV_X1    g006(.A(new_n192), .ZN(new_n193));
  INV_X1    g007(.A(KEYINPUT11), .ZN(new_n194));
  INV_X1    g008(.A(G134), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n195), .A2(KEYINPUT67), .ZN(new_n196));
  INV_X1    g010(.A(KEYINPUT67), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n197), .A2(G134), .ZN(new_n198));
  NAND3_X1  g012(.A1(new_n196), .A2(new_n198), .A3(G137), .ZN(new_n199));
  NOR2_X1   g013(.A1(G134), .A2(G137), .ZN(new_n200));
  INV_X1    g014(.A(new_n200), .ZN(new_n201));
  AOI21_X1  g015(.A(new_n194), .B1(new_n199), .B2(new_n201), .ZN(new_n202));
  INV_X1    g016(.A(G137), .ZN(new_n203));
  AND4_X1   g017(.A1(new_n194), .A2(new_n196), .A3(new_n198), .A4(new_n203), .ZN(new_n204));
  OAI21_X1  g018(.A(new_n193), .B1(new_n202), .B2(new_n204), .ZN(new_n205));
  XNOR2_X1  g019(.A(KEYINPUT67), .B(G134), .ZN(new_n206));
  NAND3_X1  g020(.A1(new_n206), .A2(new_n194), .A3(new_n203), .ZN(new_n207));
  AOI21_X1  g021(.A(new_n200), .B1(new_n206), .B2(G137), .ZN(new_n208));
  OAI211_X1 g022(.A(G131), .B(new_n207), .C1(new_n208), .C2(new_n194), .ZN(new_n209));
  AND2_X1   g023(.A1(new_n205), .A2(new_n209), .ZN(new_n210));
  INV_X1    g024(.A(G104), .ZN(new_n211));
  NOR2_X1   g025(.A1(new_n211), .A2(KEYINPUT3), .ZN(new_n212));
  INV_X1    g026(.A(KEYINPUT79), .ZN(new_n213));
  NOR2_X1   g027(.A1(new_n213), .A2(G107), .ZN(new_n214));
  INV_X1    g028(.A(G107), .ZN(new_n215));
  NOR2_X1   g029(.A1(new_n215), .A2(KEYINPUT79), .ZN(new_n216));
  OAI21_X1  g030(.A(new_n212), .B1(new_n214), .B2(new_n216), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n211), .A2(KEYINPUT3), .ZN(new_n218));
  OAI21_X1  g032(.A(G107), .B1(new_n211), .B2(KEYINPUT3), .ZN(new_n219));
  NAND4_X1  g033(.A1(new_n217), .A2(KEYINPUT80), .A3(new_n218), .A4(new_n219), .ZN(new_n220));
  INV_X1    g034(.A(KEYINPUT80), .ZN(new_n221));
  INV_X1    g035(.A(KEYINPUT3), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n222), .A2(G104), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n215), .A2(KEYINPUT79), .ZN(new_n224));
  NAND2_X1  g038(.A1(new_n213), .A2(G107), .ZN(new_n225));
  AOI21_X1  g039(.A(new_n223), .B1(new_n224), .B2(new_n225), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n219), .A2(new_n218), .ZN(new_n227));
  OAI21_X1  g041(.A(new_n221), .B1(new_n226), .B2(new_n227), .ZN(new_n228));
  NAND3_X1  g042(.A1(new_n220), .A2(new_n228), .A3(G101), .ZN(new_n229));
  INV_X1    g043(.A(KEYINPUT4), .ZN(new_n230));
  NOR2_X1   g044(.A1(new_n226), .A2(new_n227), .ZN(new_n231));
  INV_X1    g045(.A(G101), .ZN(new_n232));
  AOI21_X1  g046(.A(new_n230), .B1(new_n231), .B2(new_n232), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n229), .A2(new_n233), .ZN(new_n234));
  OR2_X1    g048(.A1(KEYINPUT0), .A2(G128), .ZN(new_n235));
  INV_X1    g049(.A(KEYINPUT64), .ZN(new_n236));
  NAND2_X1  g050(.A1(KEYINPUT0), .A2(G128), .ZN(new_n237));
  NAND3_X1  g051(.A1(new_n235), .A2(new_n236), .A3(new_n237), .ZN(new_n238));
  NAND3_X1  g052(.A1(KEYINPUT64), .A2(KEYINPUT0), .A3(G128), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n238), .A2(new_n239), .ZN(new_n240));
  INV_X1    g054(.A(G146), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n241), .A2(G143), .ZN(new_n242));
  INV_X1    g056(.A(G143), .ZN(new_n243));
  AND3_X1   g057(.A1(new_n243), .A2(KEYINPUT65), .A3(G146), .ZN(new_n244));
  AOI21_X1  g058(.A(KEYINPUT65), .B1(new_n243), .B2(G146), .ZN(new_n245));
  OAI21_X1  g059(.A(new_n242), .B1(new_n244), .B2(new_n245), .ZN(new_n246));
  NAND3_X1  g060(.A1(new_n240), .A2(new_n246), .A3(KEYINPUT66), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n243), .A2(G146), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n242), .A2(new_n248), .ZN(new_n249));
  NOR2_X1   g063(.A1(new_n249), .A2(new_n237), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n240), .A2(new_n246), .ZN(new_n251));
  INV_X1    g065(.A(KEYINPUT66), .ZN(new_n252));
  AOI21_X1  g066(.A(new_n250), .B1(new_n251), .B2(new_n252), .ZN(new_n253));
  NAND4_X1  g067(.A1(new_n220), .A2(new_n228), .A3(new_n230), .A4(G101), .ZN(new_n254));
  NAND4_X1  g068(.A1(new_n234), .A2(new_n247), .A3(new_n253), .A4(new_n254), .ZN(new_n255));
  INV_X1    g069(.A(KEYINPUT81), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n255), .A2(new_n256), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n251), .A2(new_n252), .ZN(new_n258));
  INV_X1    g072(.A(new_n250), .ZN(new_n259));
  NAND3_X1  g073(.A1(new_n258), .A2(new_n247), .A3(new_n259), .ZN(new_n260));
  INV_X1    g074(.A(new_n260), .ZN(new_n261));
  NAND4_X1  g075(.A1(new_n261), .A2(KEYINPUT81), .A3(new_n234), .A4(new_n254), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n257), .A2(new_n262), .ZN(new_n263));
  NOR2_X1   g077(.A1(new_n211), .A2(new_n215), .ZN(new_n264));
  INV_X1    g078(.A(new_n264), .ZN(new_n265));
  XNOR2_X1  g079(.A(KEYINPUT79), .B(G107), .ZN(new_n266));
  OAI211_X1 g080(.A(new_n265), .B(G101), .C1(new_n266), .C2(G104), .ZN(new_n267));
  OAI211_X1 g081(.A(new_n218), .B(new_n219), .C1(new_n266), .C2(new_n223), .ZN(new_n268));
  OAI21_X1  g082(.A(new_n267), .B1(new_n268), .B2(G101), .ZN(new_n269));
  INV_X1    g083(.A(KEYINPUT84), .ZN(new_n270));
  NAND2_X1  g084(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  OAI211_X1 g085(.A(new_n267), .B(KEYINPUT84), .C1(new_n268), .C2(G101), .ZN(new_n272));
  INV_X1    g086(.A(KEYINPUT71), .ZN(new_n273));
  NOR2_X1   g087(.A1(new_n243), .A2(G146), .ZN(new_n274));
  INV_X1    g088(.A(KEYINPUT1), .ZN(new_n275));
  OAI21_X1  g089(.A(G128), .B1(new_n274), .B2(new_n275), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n246), .A2(new_n276), .ZN(new_n277));
  NAND4_X1  g091(.A1(new_n242), .A2(new_n248), .A3(new_n275), .A4(G128), .ZN(new_n278));
  AOI21_X1  g092(.A(new_n273), .B1(new_n277), .B2(new_n278), .ZN(new_n279));
  INV_X1    g093(.A(KEYINPUT65), .ZN(new_n280));
  OAI21_X1  g094(.A(new_n280), .B1(new_n241), .B2(G143), .ZN(new_n281));
  NAND3_X1  g095(.A1(new_n243), .A2(KEYINPUT65), .A3(G146), .ZN(new_n282));
  AOI21_X1  g096(.A(new_n274), .B1(new_n281), .B2(new_n282), .ZN(new_n283));
  INV_X1    g097(.A(G128), .ZN(new_n284));
  AOI21_X1  g098(.A(new_n284), .B1(new_n242), .B2(KEYINPUT1), .ZN(new_n285));
  OAI211_X1 g099(.A(new_n273), .B(new_n278), .C1(new_n283), .C2(new_n285), .ZN(new_n286));
  INV_X1    g100(.A(new_n286), .ZN(new_n287));
  OAI211_X1 g101(.A(new_n271), .B(new_n272), .C1(new_n279), .C2(new_n287), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n288), .A2(KEYINPUT10), .ZN(new_n289));
  INV_X1    g103(.A(KEYINPUT82), .ZN(new_n290));
  NAND3_X1  g104(.A1(new_n276), .A2(new_n290), .A3(new_n249), .ZN(new_n291));
  XNOR2_X1  g105(.A(G143), .B(G146), .ZN(new_n292));
  OAI21_X1  g106(.A(KEYINPUT82), .B1(new_n285), .B2(new_n292), .ZN(new_n293));
  AND3_X1   g107(.A1(new_n291), .A2(new_n293), .A3(new_n278), .ZN(new_n294));
  OAI21_X1  g108(.A(KEYINPUT83), .B1(new_n294), .B2(new_n269), .ZN(new_n295));
  INV_X1    g109(.A(new_n269), .ZN(new_n296));
  INV_X1    g110(.A(KEYINPUT83), .ZN(new_n297));
  NAND3_X1  g111(.A1(new_n291), .A2(new_n293), .A3(new_n278), .ZN(new_n298));
  NAND3_X1  g112(.A1(new_n296), .A2(new_n297), .A3(new_n298), .ZN(new_n299));
  INV_X1    g113(.A(KEYINPUT10), .ZN(new_n300));
  NAND3_X1  g114(.A1(new_n295), .A2(new_n299), .A3(new_n300), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n289), .A2(new_n301), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n263), .A2(new_n302), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n303), .A2(KEYINPUT87), .ZN(new_n304));
  AOI22_X1  g118(.A1(new_n257), .A2(new_n262), .B1(new_n289), .B2(new_n301), .ZN(new_n305));
  INV_X1    g119(.A(KEYINPUT87), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n305), .A2(new_n306), .ZN(new_n307));
  AOI21_X1  g121(.A(new_n210), .B1(new_n304), .B2(new_n307), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n205), .A2(new_n209), .ZN(new_n309));
  NOR2_X1   g123(.A1(new_n303), .A2(new_n309), .ZN(new_n310));
  OAI21_X1  g124(.A(new_n191), .B1(new_n308), .B2(new_n310), .ZN(new_n311));
  INV_X1    g125(.A(KEYINPUT88), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n311), .A2(new_n312), .ZN(new_n313));
  AND3_X1   g127(.A1(new_n263), .A2(new_n306), .A3(new_n302), .ZN(new_n314));
  AOI21_X1  g128(.A(new_n306), .B1(new_n263), .B2(new_n302), .ZN(new_n315));
  OAI21_X1  g129(.A(new_n309), .B1(new_n314), .B2(new_n315), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n305), .A2(new_n210), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n316), .A2(new_n317), .ZN(new_n318));
  NAND3_X1  g132(.A1(new_n318), .A2(KEYINPUT88), .A3(new_n191), .ZN(new_n319));
  NOR2_X1   g133(.A1(new_n310), .A2(new_n191), .ZN(new_n320));
  AND2_X1   g134(.A1(new_n295), .A2(new_n299), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n277), .A2(new_n278), .ZN(new_n322));
  OAI21_X1  g136(.A(KEYINPUT85), .B1(new_n296), .B2(new_n322), .ZN(new_n323));
  AND2_X1   g137(.A1(new_n277), .A2(new_n278), .ZN(new_n324));
  INV_X1    g138(.A(KEYINPUT85), .ZN(new_n325));
  NAND3_X1  g139(.A1(new_n324), .A2(new_n325), .A3(new_n269), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n323), .A2(new_n326), .ZN(new_n327));
  OAI21_X1  g141(.A(new_n309), .B1(new_n321), .B2(new_n327), .ZN(new_n328));
  INV_X1    g142(.A(KEYINPUT12), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n328), .A2(new_n329), .ZN(new_n330));
  OAI211_X1 g144(.A(KEYINPUT12), .B(new_n309), .C1(new_n321), .C2(new_n327), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n330), .A2(new_n331), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n320), .A2(new_n332), .ZN(new_n333));
  NAND3_X1  g147(.A1(new_n313), .A2(new_n319), .A3(new_n333), .ZN(new_n334));
  INV_X1    g148(.A(G469), .ZN(new_n335));
  INV_X1    g149(.A(G902), .ZN(new_n336));
  NAND3_X1  g150(.A1(new_n334), .A2(new_n335), .A3(new_n336), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n320), .A2(new_n316), .ZN(new_n338));
  AOI22_X1  g152(.A1(new_n330), .A2(new_n331), .B1(new_n305), .B2(new_n210), .ZN(new_n339));
  OAI21_X1  g153(.A(new_n191), .B1(new_n339), .B2(KEYINPUT86), .ZN(new_n340));
  NAND3_X1  g154(.A1(new_n332), .A2(KEYINPUT86), .A3(new_n317), .ZN(new_n341));
  INV_X1    g155(.A(new_n341), .ZN(new_n342));
  OAI211_X1 g156(.A(G469), .B(new_n338), .C1(new_n340), .C2(new_n342), .ZN(new_n343));
  NAND2_X1  g157(.A1(G469), .A2(G902), .ZN(new_n344));
  NAND3_X1  g158(.A1(new_n337), .A2(new_n343), .A3(new_n344), .ZN(new_n345));
  XOR2_X1   g159(.A(KEYINPUT9), .B(G234), .Z(new_n346));
  INV_X1    g160(.A(new_n346), .ZN(new_n347));
  OAI21_X1  g161(.A(G221), .B1(new_n347), .B2(G902), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n345), .A2(new_n348), .ZN(new_n349));
  INV_X1    g163(.A(G125), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n324), .A2(new_n350), .ZN(new_n351));
  OR2_X1    g165(.A1(new_n351), .A2(KEYINPUT89), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n351), .A2(KEYINPUT89), .ZN(new_n353));
  NAND2_X1  g167(.A1(new_n260), .A2(G125), .ZN(new_n354));
  NAND3_X1  g168(.A1(new_n352), .A2(new_n353), .A3(new_n354), .ZN(new_n355));
  INV_X1    g169(.A(G224), .ZN(new_n356));
  NOR2_X1   g170(.A1(new_n356), .A2(G953), .ZN(new_n357));
  XNOR2_X1  g171(.A(new_n355), .B(new_n357), .ZN(new_n358));
  INV_X1    g172(.A(G119), .ZN(new_n359));
  NAND2_X1  g173(.A1(new_n359), .A2(G116), .ZN(new_n360));
  INV_X1    g174(.A(new_n360), .ZN(new_n361));
  XNOR2_X1  g175(.A(KEYINPUT70), .B(G116), .ZN(new_n362));
  AOI21_X1  g176(.A(new_n361), .B1(new_n362), .B2(G119), .ZN(new_n363));
  XOR2_X1   g177(.A(KEYINPUT2), .B(G113), .Z(new_n364));
  AND2_X1   g178(.A1(new_n363), .A2(new_n364), .ZN(new_n365));
  OAI21_X1  g179(.A(G113), .B1(new_n360), .B2(KEYINPUT5), .ZN(new_n366));
  INV_X1    g180(.A(new_n366), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n363), .A2(KEYINPUT5), .ZN(new_n368));
  AOI21_X1  g182(.A(new_n365), .B1(new_n367), .B2(new_n368), .ZN(new_n369));
  NAND3_X1  g183(.A1(new_n369), .A2(new_n271), .A3(new_n272), .ZN(new_n370));
  XNOR2_X1  g184(.A(new_n363), .B(new_n364), .ZN(new_n371));
  NAND3_X1  g185(.A1(new_n234), .A2(new_n371), .A3(new_n254), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n370), .A2(new_n372), .ZN(new_n373));
  XOR2_X1   g187(.A(G110), .B(G122), .Z(new_n374));
  OR2_X1    g188(.A1(new_n373), .A2(new_n374), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n373), .A2(new_n374), .ZN(new_n376));
  NAND3_X1  g190(.A1(new_n375), .A2(KEYINPUT6), .A3(new_n376), .ZN(new_n377));
  INV_X1    g191(.A(KEYINPUT6), .ZN(new_n378));
  NAND3_X1  g192(.A1(new_n373), .A2(new_n378), .A3(new_n374), .ZN(new_n379));
  NAND3_X1  g193(.A1(new_n358), .A2(new_n377), .A3(new_n379), .ZN(new_n380));
  AND2_X1   g194(.A1(new_n352), .A2(new_n354), .ZN(new_n381));
  INV_X1    g195(.A(new_n357), .ZN(new_n382));
  NAND4_X1  g196(.A1(new_n381), .A2(KEYINPUT7), .A3(new_n382), .A4(new_n353), .ZN(new_n383));
  XOR2_X1   g197(.A(new_n368), .B(KEYINPUT90), .Z(new_n384));
  NOR2_X1   g198(.A1(new_n384), .A2(new_n366), .ZN(new_n385));
  OAI21_X1  g199(.A(new_n296), .B1(new_n385), .B2(new_n365), .ZN(new_n386));
  XNOR2_X1  g200(.A(new_n374), .B(KEYINPUT8), .ZN(new_n387));
  AOI21_X1  g201(.A(new_n387), .B1(new_n369), .B2(new_n269), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n386), .A2(new_n388), .ZN(new_n389));
  INV_X1    g203(.A(KEYINPUT7), .ZN(new_n390));
  OAI21_X1  g204(.A(new_n355), .B1(new_n390), .B2(new_n357), .ZN(new_n391));
  NAND4_X1  g205(.A1(new_n383), .A2(new_n389), .A3(new_n391), .A4(new_n375), .ZN(new_n392));
  NAND3_X1  g206(.A1(new_n380), .A2(new_n336), .A3(new_n392), .ZN(new_n393));
  OAI21_X1  g207(.A(G210), .B1(G237), .B2(G902), .ZN(new_n394));
  INV_X1    g208(.A(new_n394), .ZN(new_n395));
  OAI21_X1  g209(.A(KEYINPUT92), .B1(new_n393), .B2(new_n395), .ZN(new_n396));
  INV_X1    g210(.A(KEYINPUT91), .ZN(new_n397));
  NAND3_X1  g211(.A1(new_n393), .A2(new_n397), .A3(new_n395), .ZN(new_n398));
  AOI21_X1  g212(.A(KEYINPUT92), .B1(new_n395), .B2(new_n397), .ZN(new_n399));
  NAND4_X1  g213(.A1(new_n380), .A2(new_n336), .A3(new_n392), .A4(new_n399), .ZN(new_n400));
  NAND3_X1  g214(.A1(new_n396), .A2(new_n398), .A3(new_n400), .ZN(new_n401));
  OAI21_X1  g215(.A(G214), .B1(G237), .B2(G902), .ZN(new_n402));
  INV_X1    g216(.A(G953), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n403), .A2(G952), .ZN(new_n404));
  AOI21_X1  g218(.A(new_n404), .B1(G234), .B2(G237), .ZN(new_n405));
  INV_X1    g219(.A(new_n405), .ZN(new_n406));
  AOI211_X1 g220(.A(new_n336), .B(new_n403), .C1(G234), .C2(G237), .ZN(new_n407));
  INV_X1    g221(.A(new_n407), .ZN(new_n408));
  XOR2_X1   g222(.A(KEYINPUT21), .B(G898), .Z(new_n409));
  OAI21_X1  g223(.A(new_n406), .B1(new_n408), .B2(new_n409), .ZN(new_n410));
  NAND3_X1  g224(.A1(new_n401), .A2(new_n402), .A3(new_n410), .ZN(new_n411));
  NOR2_X1   g225(.A1(new_n349), .A2(new_n411), .ZN(new_n412));
  INV_X1    g226(.A(KEYINPUT16), .ZN(new_n413));
  INV_X1    g227(.A(G140), .ZN(new_n414));
  NAND3_X1  g228(.A1(new_n413), .A2(new_n414), .A3(G125), .ZN(new_n415));
  OR2_X1    g229(.A1(new_n415), .A2(KEYINPUT76), .ZN(new_n416));
  XNOR2_X1  g230(.A(G125), .B(G140), .ZN(new_n417));
  NAND2_X1  g231(.A1(new_n417), .A2(KEYINPUT16), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n415), .A2(KEYINPUT76), .ZN(new_n419));
  NAND3_X1  g233(.A1(new_n416), .A2(new_n418), .A3(new_n419), .ZN(new_n420));
  OR2_X1    g234(.A1(new_n420), .A2(new_n241), .ZN(new_n421));
  INV_X1    g235(.A(KEYINPUT77), .ZN(new_n422));
  AOI21_X1  g236(.A(new_n422), .B1(new_n420), .B2(new_n241), .ZN(new_n423));
  OR2_X1    g237(.A1(new_n421), .A2(new_n423), .ZN(new_n424));
  XOR2_X1   g238(.A(KEYINPUT24), .B(G110), .Z(new_n425));
  XNOR2_X1  g239(.A(new_n425), .B(KEYINPUT75), .ZN(new_n426));
  XNOR2_X1  g240(.A(G119), .B(G128), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n426), .A2(new_n427), .ZN(new_n428));
  NOR3_X1   g242(.A1(new_n359), .A2(KEYINPUT23), .A3(G128), .ZN(new_n429));
  AOI21_X1  g243(.A(new_n429), .B1(new_n427), .B2(KEYINPUT23), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n430), .A2(G110), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n421), .A2(new_n423), .ZN(new_n432));
  NAND4_X1  g246(.A1(new_n424), .A2(new_n428), .A3(new_n431), .A4(new_n432), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n417), .A2(new_n241), .ZN(new_n434));
  NOR2_X1   g248(.A1(new_n426), .A2(new_n427), .ZN(new_n435));
  XOR2_X1   g249(.A(KEYINPUT78), .B(G110), .Z(new_n436));
  NOR2_X1   g250(.A1(new_n430), .A2(new_n436), .ZN(new_n437));
  OAI211_X1 g251(.A(new_n421), .B(new_n434), .C1(new_n435), .C2(new_n437), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n433), .A2(new_n438), .ZN(new_n439));
  NAND3_X1  g253(.A1(new_n403), .A2(G221), .A3(G234), .ZN(new_n440));
  XNOR2_X1  g254(.A(new_n440), .B(KEYINPUT22), .ZN(new_n441));
  XNOR2_X1  g255(.A(new_n441), .B(G137), .ZN(new_n442));
  XNOR2_X1  g256(.A(new_n439), .B(new_n442), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n443), .A2(new_n336), .ZN(new_n444));
  INV_X1    g258(.A(KEYINPUT25), .ZN(new_n445));
  XNOR2_X1  g259(.A(new_n444), .B(new_n445), .ZN(new_n446));
  INV_X1    g260(.A(G217), .ZN(new_n447));
  AOI21_X1  g261(.A(new_n447), .B1(G234), .B2(new_n336), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n446), .A2(new_n448), .ZN(new_n449));
  OR2_X1    g263(.A1(new_n444), .A2(new_n448), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n449), .A2(new_n450), .ZN(new_n451));
  INV_X1    g265(.A(KEYINPUT69), .ZN(new_n452));
  OAI21_X1  g266(.A(new_n452), .B1(new_n210), .B2(new_n260), .ZN(new_n453));
  NAND4_X1  g267(.A1(new_n309), .A2(KEYINPUT69), .A3(new_n247), .A4(new_n253), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n195), .A2(G137), .ZN(new_n455));
  INV_X1    g269(.A(new_n206), .ZN(new_n456));
  OAI21_X1  g270(.A(new_n455), .B1(new_n456), .B2(G137), .ZN(new_n457));
  NAND2_X1  g271(.A1(new_n457), .A2(G131), .ZN(new_n458));
  AND2_X1   g272(.A1(new_n205), .A2(new_n458), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n459), .A2(new_n322), .ZN(new_n460));
  NAND3_X1  g274(.A1(new_n453), .A2(new_n454), .A3(new_n460), .ZN(new_n461));
  INV_X1    g275(.A(KEYINPUT30), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n199), .A2(new_n201), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n464), .A2(KEYINPUT11), .ZN(new_n465));
  AOI21_X1  g279(.A(new_n192), .B1(new_n465), .B2(new_n207), .ZN(new_n466));
  INV_X1    g280(.A(G131), .ZN(new_n467));
  NOR3_X1   g281(.A1(new_n202), .A2(new_n467), .A3(new_n204), .ZN(new_n468));
  OAI211_X1 g282(.A(new_n247), .B(new_n253), .C1(new_n466), .C2(new_n468), .ZN(new_n469));
  OAI211_X1 g283(.A(new_n205), .B(new_n458), .C1(new_n279), .C2(new_n287), .ZN(new_n470));
  AND2_X1   g284(.A1(new_n469), .A2(new_n470), .ZN(new_n471));
  NAND2_X1  g285(.A1(new_n471), .A2(KEYINPUT30), .ZN(new_n472));
  NAND3_X1  g286(.A1(new_n463), .A2(new_n371), .A3(new_n472), .ZN(new_n473));
  INV_X1    g287(.A(new_n371), .ZN(new_n474));
  NAND3_X1  g288(.A1(new_n469), .A2(new_n470), .A3(new_n474), .ZN(new_n475));
  XNOR2_X1  g289(.A(KEYINPUT26), .B(KEYINPUT27), .ZN(new_n476));
  XNOR2_X1  g290(.A(new_n476), .B(G101), .ZN(new_n477));
  INV_X1    g291(.A(G237), .ZN(new_n478));
  NAND3_X1  g292(.A1(new_n478), .A2(new_n403), .A3(G210), .ZN(new_n479));
  XNOR2_X1  g293(.A(new_n477), .B(new_n479), .ZN(new_n480));
  NAND3_X1  g294(.A1(new_n473), .A2(new_n475), .A3(new_n480), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n481), .A2(KEYINPUT31), .ZN(new_n482));
  INV_X1    g296(.A(KEYINPUT28), .ZN(new_n483));
  AOI21_X1  g297(.A(KEYINPUT72), .B1(new_n475), .B2(new_n483), .ZN(new_n484));
  AND3_X1   g298(.A1(new_n469), .A2(new_n470), .A3(new_n474), .ZN(new_n485));
  AOI21_X1  g299(.A(new_n485), .B1(new_n461), .B2(new_n371), .ZN(new_n486));
  OAI21_X1  g300(.A(new_n484), .B1(new_n486), .B2(new_n483), .ZN(new_n487));
  INV_X1    g301(.A(new_n480), .ZN(new_n488));
  AOI22_X1  g302(.A1(new_n469), .A2(new_n452), .B1(new_n459), .B2(new_n322), .ZN(new_n489));
  AOI21_X1  g303(.A(new_n474), .B1(new_n489), .B2(new_n454), .ZN(new_n490));
  OAI211_X1 g304(.A(KEYINPUT72), .B(KEYINPUT28), .C1(new_n490), .C2(new_n485), .ZN(new_n491));
  NAND3_X1  g305(.A1(new_n487), .A2(new_n488), .A3(new_n491), .ZN(new_n492));
  INV_X1    g306(.A(KEYINPUT31), .ZN(new_n493));
  NAND4_X1  g307(.A1(new_n473), .A2(new_n493), .A3(new_n475), .A4(new_n480), .ZN(new_n494));
  NAND3_X1  g308(.A1(new_n482), .A2(new_n492), .A3(new_n494), .ZN(new_n495));
  NOR2_X1   g309(.A1(G472), .A2(G902), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  INV_X1    g311(.A(KEYINPUT32), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  INV_X1    g313(.A(KEYINPUT74), .ZN(new_n500));
  NAND3_X1  g314(.A1(new_n495), .A2(KEYINPUT32), .A3(new_n496), .ZN(new_n501));
  NAND3_X1  g315(.A1(new_n499), .A2(new_n500), .A3(new_n501), .ZN(new_n502));
  AND3_X1   g316(.A1(new_n495), .A2(KEYINPUT32), .A3(new_n496), .ZN(new_n503));
  AOI21_X1  g317(.A(KEYINPUT32), .B1(new_n495), .B2(new_n496), .ZN(new_n504));
  OAI21_X1  g318(.A(new_n503), .B1(new_n504), .B2(KEYINPUT74), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n502), .A2(new_n505), .ZN(new_n506));
  NAND3_X1  g320(.A1(new_n487), .A2(new_n480), .A3(new_n491), .ZN(new_n507));
  NAND3_X1  g321(.A1(new_n473), .A2(new_n475), .A3(new_n488), .ZN(new_n508));
  AOI21_X1  g322(.A(KEYINPUT29), .B1(new_n507), .B2(new_n508), .ZN(new_n509));
  NOR2_X1   g323(.A1(new_n485), .A2(KEYINPUT28), .ZN(new_n510));
  XNOR2_X1  g324(.A(new_n471), .B(new_n474), .ZN(new_n511));
  AOI21_X1  g325(.A(new_n510), .B1(new_n511), .B2(KEYINPUT28), .ZN(new_n512));
  INV_X1    g326(.A(KEYINPUT29), .ZN(new_n513));
  NOR2_X1   g327(.A1(new_n488), .A2(new_n513), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n512), .A2(new_n514), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n515), .A2(new_n336), .ZN(new_n516));
  OAI21_X1  g330(.A(G472), .B1(new_n509), .B2(new_n516), .ZN(new_n517));
  NAND2_X1  g331(.A1(new_n517), .A2(KEYINPUT73), .ZN(new_n518));
  INV_X1    g332(.A(KEYINPUT73), .ZN(new_n519));
  OAI211_X1 g333(.A(new_n519), .B(G472), .C1(new_n509), .C2(new_n516), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n518), .A2(new_n520), .ZN(new_n521));
  AOI21_X1  g335(.A(new_n451), .B1(new_n506), .B2(new_n521), .ZN(new_n522));
  XNOR2_X1  g336(.A(new_n417), .B(new_n241), .ZN(new_n523));
  INV_X1    g337(.A(KEYINPUT94), .ZN(new_n524));
  OR2_X1    g338(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  NAND3_X1  g339(.A1(new_n478), .A2(new_n403), .A3(G214), .ZN(new_n526));
  XNOR2_X1  g340(.A(new_n526), .B(G143), .ZN(new_n527));
  INV_X1    g341(.A(new_n527), .ZN(new_n528));
  NAND3_X1  g342(.A1(new_n528), .A2(KEYINPUT18), .A3(G131), .ZN(new_n529));
  NAND2_X1  g343(.A1(new_n523), .A2(new_n524), .ZN(new_n530));
  INV_X1    g344(.A(KEYINPUT18), .ZN(new_n531));
  OAI21_X1  g345(.A(new_n527), .B1(new_n531), .B2(new_n467), .ZN(new_n532));
  NAND4_X1  g346(.A1(new_n525), .A2(new_n529), .A3(new_n530), .A4(new_n532), .ZN(new_n533));
  XNOR2_X1  g347(.A(new_n527), .B(new_n193), .ZN(new_n534));
  XNOR2_X1  g348(.A(new_n417), .B(KEYINPUT19), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n535), .A2(new_n241), .ZN(new_n536));
  NAND3_X1  g350(.A1(new_n534), .A2(new_n421), .A3(new_n536), .ZN(new_n537));
  XOR2_X1   g351(.A(G113), .B(G122), .Z(new_n538));
  XNOR2_X1  g352(.A(new_n538), .B(KEYINPUT95), .ZN(new_n539));
  XNOR2_X1  g353(.A(new_n539), .B(new_n211), .ZN(new_n540));
  AND3_X1   g354(.A1(new_n533), .A2(new_n537), .A3(new_n540), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n424), .A2(new_n432), .ZN(new_n542));
  NAND3_X1  g356(.A1(new_n528), .A2(KEYINPUT17), .A3(new_n192), .ZN(new_n543));
  OAI211_X1 g357(.A(new_n542), .B(new_n543), .C1(KEYINPUT17), .C2(new_n534), .ZN(new_n544));
  NAND2_X1  g358(.A1(new_n544), .A2(new_n533), .ZN(new_n545));
  INV_X1    g359(.A(new_n540), .ZN(new_n546));
  AOI21_X1  g360(.A(new_n541), .B1(new_n545), .B2(new_n546), .ZN(new_n547));
  INV_X1    g361(.A(G475), .ZN(new_n548));
  NAND3_X1  g362(.A1(new_n547), .A2(new_n548), .A3(new_n336), .ZN(new_n549));
  OR2_X1    g363(.A1(new_n549), .A2(KEYINPUT20), .ZN(new_n550));
  XOR2_X1   g364(.A(KEYINPUT93), .B(KEYINPUT20), .Z(new_n551));
  NAND2_X1  g365(.A1(new_n549), .A2(new_n551), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n540), .A2(KEYINPUT96), .ZN(new_n553));
  AOI21_X1  g367(.A(G902), .B1(new_n545), .B2(new_n553), .ZN(new_n554));
  OAI21_X1  g368(.A(new_n554), .B1(new_n545), .B2(new_n553), .ZN(new_n555));
  AOI22_X1  g369(.A1(new_n550), .A2(new_n552), .B1(G475), .B2(new_n555), .ZN(new_n556));
  INV_X1    g370(.A(new_n556), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n284), .A2(G143), .ZN(new_n558));
  NOR2_X1   g372(.A1(new_n284), .A2(G143), .ZN(new_n559));
  OAI21_X1  g373(.A(new_n558), .B1(new_n559), .B2(KEYINPUT13), .ZN(new_n560));
  XNOR2_X1  g374(.A(new_n560), .B(KEYINPUT98), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n559), .A2(KEYINPUT13), .ZN(new_n562));
  AOI21_X1  g376(.A(new_n195), .B1(new_n561), .B2(new_n562), .ZN(new_n563));
  XOR2_X1   g377(.A(new_n563), .B(KEYINPUT99), .Z(new_n564));
  INV_X1    g378(.A(new_n559), .ZN(new_n565));
  NAND3_X1  g379(.A1(new_n456), .A2(new_n565), .A3(new_n558), .ZN(new_n566));
  INV_X1    g380(.A(G116), .ZN(new_n567));
  NOR2_X1   g381(.A1(new_n567), .A2(G122), .ZN(new_n568));
  XNOR2_X1  g382(.A(new_n568), .B(KEYINPUT97), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n362), .A2(G122), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n569), .A2(new_n570), .ZN(new_n571));
  NOR2_X1   g385(.A1(new_n571), .A2(new_n266), .ZN(new_n572));
  AND2_X1   g386(.A1(new_n571), .A2(new_n266), .ZN(new_n573));
  OAI211_X1 g387(.A(new_n564), .B(new_n566), .C1(new_n572), .C2(new_n573), .ZN(new_n574));
  NOR3_X1   g388(.A1(new_n347), .A2(new_n447), .A3(G953), .ZN(new_n575));
  XOR2_X1   g389(.A(new_n572), .B(KEYINPUT100), .Z(new_n576));
  NAND2_X1  g390(.A1(new_n565), .A2(new_n558), .ZN(new_n577));
  NAND2_X1  g391(.A1(new_n577), .A2(new_n206), .ZN(new_n578));
  NAND2_X1  g392(.A1(new_n566), .A2(new_n578), .ZN(new_n579));
  INV_X1    g393(.A(new_n570), .ZN(new_n580));
  INV_X1    g394(.A(KEYINPUT14), .ZN(new_n581));
  NAND2_X1  g395(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  INV_X1    g396(.A(new_n582), .ZN(new_n583));
  OAI21_X1  g397(.A(new_n569), .B1(new_n580), .B2(new_n581), .ZN(new_n584));
  OAI21_X1  g398(.A(G107), .B1(new_n583), .B2(new_n584), .ZN(new_n585));
  NAND3_X1  g399(.A1(new_n576), .A2(new_n579), .A3(new_n585), .ZN(new_n586));
  NAND3_X1  g400(.A1(new_n574), .A2(new_n575), .A3(new_n586), .ZN(new_n587));
  INV_X1    g401(.A(new_n587), .ZN(new_n588));
  AOI21_X1  g402(.A(new_n575), .B1(new_n574), .B2(new_n586), .ZN(new_n589));
  OAI21_X1  g403(.A(new_n336), .B1(new_n588), .B2(new_n589), .ZN(new_n590));
  INV_X1    g404(.A(G478), .ZN(new_n591));
  NOR2_X1   g405(.A1(new_n591), .A2(KEYINPUT15), .ZN(new_n592));
  XNOR2_X1  g406(.A(new_n590), .B(new_n592), .ZN(new_n593));
  NOR2_X1   g407(.A1(new_n557), .A2(new_n593), .ZN(new_n594));
  NAND3_X1  g408(.A1(new_n412), .A2(new_n522), .A3(new_n594), .ZN(new_n595));
  XNOR2_X1  g409(.A(new_n595), .B(G101), .ZN(G3));
  NAND2_X1  g410(.A1(new_n495), .A2(new_n336), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n597), .A2(G472), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n598), .A2(new_n497), .ZN(new_n599));
  NOR2_X1   g413(.A1(new_n349), .A2(new_n599), .ZN(new_n600));
  INV_X1    g414(.A(new_n451), .ZN(new_n601));
  XNOR2_X1  g415(.A(new_n393), .B(new_n394), .ZN(new_n602));
  INV_X1    g416(.A(new_n402), .ZN(new_n603));
  NOR2_X1   g417(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  AND2_X1   g418(.A1(new_n604), .A2(new_n410), .ZN(new_n605));
  OAI211_X1 g419(.A(new_n591), .B(new_n336), .C1(new_n588), .C2(new_n589), .ZN(new_n606));
  NAND2_X1  g420(.A1(G478), .A2(G902), .ZN(new_n607));
  OAI21_X1  g421(.A(KEYINPUT33), .B1(new_n588), .B2(new_n589), .ZN(new_n608));
  INV_X1    g422(.A(new_n589), .ZN(new_n609));
  INV_X1    g423(.A(KEYINPUT33), .ZN(new_n610));
  NAND3_X1  g424(.A1(new_n609), .A2(new_n610), .A3(new_n587), .ZN(new_n611));
  NAND2_X1  g425(.A1(new_n608), .A2(new_n611), .ZN(new_n612));
  OAI211_X1 g426(.A(new_n606), .B(new_n607), .C1(new_n612), .C2(new_n591), .ZN(new_n613));
  NOR2_X1   g427(.A1(new_n613), .A2(new_n556), .ZN(new_n614));
  AND2_X1   g428(.A1(new_n605), .A2(new_n614), .ZN(new_n615));
  NAND3_X1  g429(.A1(new_n600), .A2(new_n601), .A3(new_n615), .ZN(new_n616));
  XOR2_X1   g430(.A(KEYINPUT34), .B(G104), .Z(new_n617));
  XNOR2_X1  g431(.A(new_n616), .B(new_n617), .ZN(G6));
  NAND2_X1  g432(.A1(new_n555), .A2(G475), .ZN(new_n619));
  XNOR2_X1  g433(.A(new_n549), .B(new_n551), .ZN(new_n620));
  AND2_X1   g434(.A1(new_n593), .A2(new_n620), .ZN(new_n621));
  AND3_X1   g435(.A1(new_n605), .A2(new_n619), .A3(new_n621), .ZN(new_n622));
  NAND3_X1  g436(.A1(new_n600), .A2(new_n622), .A3(new_n601), .ZN(new_n623));
  XOR2_X1   g437(.A(KEYINPUT35), .B(G107), .Z(new_n624));
  XNOR2_X1  g438(.A(new_n623), .B(new_n624), .ZN(G9));
  INV_X1    g439(.A(new_n599), .ZN(new_n626));
  INV_X1    g440(.A(new_n442), .ZN(new_n627));
  NOR2_X1   g441(.A1(new_n627), .A2(KEYINPUT36), .ZN(new_n628));
  XNOR2_X1  g442(.A(new_n439), .B(new_n628), .ZN(new_n629));
  NOR2_X1   g443(.A1(new_n448), .A2(G902), .ZN(new_n630));
  NAND2_X1  g444(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n449), .A2(new_n631), .ZN(new_n632));
  NAND4_X1  g446(.A1(new_n412), .A2(new_n594), .A3(new_n626), .A4(new_n632), .ZN(new_n633));
  XOR2_X1   g447(.A(new_n633), .B(KEYINPUT37), .Z(new_n634));
  XNOR2_X1  g448(.A(new_n634), .B(G110), .ZN(G12));
  NOR3_X1   g449(.A1(new_n503), .A2(new_n504), .A3(KEYINPUT74), .ZN(new_n636));
  NOR3_X1   g450(.A1(new_n497), .A2(new_n500), .A3(new_n498), .ZN(new_n637));
  OAI21_X1  g451(.A(new_n521), .B1(new_n636), .B2(new_n637), .ZN(new_n638));
  NAND3_X1  g452(.A1(new_n638), .A2(new_n604), .A3(new_n632), .ZN(new_n639));
  XOR2_X1   g453(.A(KEYINPUT101), .B(G900), .Z(new_n640));
  AOI21_X1  g454(.A(new_n405), .B1(new_n407), .B2(new_n640), .ZN(new_n641));
  AOI21_X1  g455(.A(new_n641), .B1(new_n555), .B2(G475), .ZN(new_n642));
  NAND3_X1  g456(.A1(new_n593), .A2(new_n620), .A3(new_n642), .ZN(new_n643));
  INV_X1    g457(.A(new_n643), .ZN(new_n644));
  NAND3_X1  g458(.A1(new_n345), .A2(new_n644), .A3(new_n348), .ZN(new_n645));
  OAI21_X1  g459(.A(KEYINPUT102), .B1(new_n639), .B2(new_n645), .ZN(new_n646));
  AND3_X1   g460(.A1(new_n345), .A2(new_n348), .A3(new_n644), .ZN(new_n647));
  INV_X1    g461(.A(KEYINPUT102), .ZN(new_n648));
  AOI22_X1  g462(.A1(new_n446), .A2(new_n448), .B1(new_n629), .B2(new_n630), .ZN(new_n649));
  AOI21_X1  g463(.A(new_n649), .B1(new_n506), .B2(new_n521), .ZN(new_n650));
  NAND4_X1  g464(.A1(new_n647), .A2(new_n648), .A3(new_n604), .A4(new_n650), .ZN(new_n651));
  NAND2_X1  g465(.A1(new_n646), .A2(new_n651), .ZN(new_n652));
  XNOR2_X1  g466(.A(new_n652), .B(G128), .ZN(G30));
  INV_X1    g467(.A(new_n349), .ZN(new_n654));
  XOR2_X1   g468(.A(new_n641), .B(KEYINPUT39), .Z(new_n655));
  NAND2_X1  g469(.A1(new_n654), .A2(new_n655), .ZN(new_n656));
  NOR2_X1   g470(.A1(new_n656), .A2(KEYINPUT40), .ZN(new_n657));
  INV_X1    g471(.A(new_n593), .ZN(new_n658));
  NOR3_X1   g472(.A1(new_n657), .A2(new_n658), .A3(new_n556), .ZN(new_n659));
  AOI21_X1  g473(.A(new_n632), .B1(new_n656), .B2(KEYINPUT40), .ZN(new_n660));
  AOI21_X1  g474(.A(new_n488), .B1(new_n473), .B2(new_n475), .ZN(new_n661));
  OAI21_X1  g475(.A(new_n336), .B1(new_n511), .B2(new_n480), .ZN(new_n662));
  OAI21_X1  g476(.A(G472), .B1(new_n661), .B2(new_n662), .ZN(new_n663));
  NAND2_X1  g477(.A1(new_n506), .A2(new_n663), .ZN(new_n664));
  INV_X1    g478(.A(new_n664), .ZN(new_n665));
  NOR2_X1   g479(.A1(new_n665), .A2(new_n603), .ZN(new_n666));
  XOR2_X1   g480(.A(new_n401), .B(KEYINPUT103), .Z(new_n667));
  XNOR2_X1  g481(.A(new_n667), .B(KEYINPUT38), .ZN(new_n668));
  NAND4_X1  g482(.A1(new_n659), .A2(new_n660), .A3(new_n666), .A4(new_n668), .ZN(new_n669));
  XNOR2_X1  g483(.A(new_n669), .B(G143), .ZN(G45));
  NOR3_X1   g484(.A1(new_n613), .A2(new_n556), .A3(new_n641), .ZN(new_n671));
  NAND3_X1  g485(.A1(new_n345), .A2(new_n671), .A3(new_n348), .ZN(new_n672));
  NOR2_X1   g486(.A1(new_n639), .A2(new_n672), .ZN(new_n673));
  XNOR2_X1  g487(.A(new_n673), .B(new_n241), .ZN(G48));
  AOI21_X1  g488(.A(KEYINPUT88), .B1(new_n318), .B2(new_n191), .ZN(new_n675));
  AOI211_X1 g489(.A(new_n312), .B(new_n190), .C1(new_n316), .C2(new_n317), .ZN(new_n676));
  INV_X1    g490(.A(new_n333), .ZN(new_n677));
  NOR3_X1   g491(.A1(new_n675), .A2(new_n676), .A3(new_n677), .ZN(new_n678));
  OAI21_X1  g492(.A(G469), .B1(new_n678), .B2(G902), .ZN(new_n679));
  NAND3_X1  g493(.A1(new_n679), .A2(new_n348), .A3(new_n337), .ZN(new_n680));
  INV_X1    g494(.A(KEYINPUT104), .ZN(new_n681));
  NAND2_X1  g495(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  NAND4_X1  g496(.A1(new_n679), .A2(KEYINPUT104), .A3(new_n348), .A4(new_n337), .ZN(new_n683));
  AND3_X1   g497(.A1(new_n682), .A2(KEYINPUT105), .A3(new_n683), .ZN(new_n684));
  AOI21_X1  g498(.A(KEYINPUT105), .B1(new_n682), .B2(new_n683), .ZN(new_n685));
  OAI211_X1 g499(.A(new_n522), .B(new_n615), .C1(new_n684), .C2(new_n685), .ZN(new_n686));
  XNOR2_X1  g500(.A(KEYINPUT41), .B(G113), .ZN(new_n687));
  XNOR2_X1  g501(.A(new_n686), .B(new_n687), .ZN(G15));
  OAI211_X1 g502(.A(new_n522), .B(new_n622), .C1(new_n684), .C2(new_n685), .ZN(new_n689));
  XNOR2_X1  g503(.A(new_n689), .B(G116), .ZN(G18));
  NAND4_X1  g504(.A1(new_n682), .A2(new_n604), .A3(new_n650), .A4(new_n683), .ZN(new_n691));
  NAND2_X1  g505(.A1(new_n594), .A2(new_n410), .ZN(new_n692));
  NOR2_X1   g506(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  XNOR2_X1  g507(.A(new_n693), .B(new_n359), .ZN(G21));
  OAI211_X1 g508(.A(new_n482), .B(new_n494), .C1(new_n480), .C2(new_n512), .ZN(new_n695));
  XOR2_X1   g509(.A(new_n496), .B(KEYINPUT106), .Z(new_n696));
  AND2_X1   g510(.A1(new_n695), .A2(new_n696), .ZN(new_n697));
  AOI211_X1 g511(.A(new_n697), .B(new_n451), .C1(G472), .C2(new_n597), .ZN(new_n698));
  NOR2_X1   g512(.A1(new_n658), .A2(new_n556), .ZN(new_n699));
  AND3_X1   g513(.A1(new_n699), .A2(new_n410), .A3(new_n604), .ZN(new_n700));
  OAI211_X1 g514(.A(new_n698), .B(new_n700), .C1(new_n684), .C2(new_n685), .ZN(new_n701));
  XNOR2_X1  g515(.A(new_n701), .B(G122), .ZN(G24));
  AND3_X1   g516(.A1(new_n334), .A2(new_n335), .A3(new_n336), .ZN(new_n703));
  AOI21_X1  g517(.A(new_n335), .B1(new_n334), .B2(new_n336), .ZN(new_n704));
  NOR2_X1   g518(.A1(new_n703), .A2(new_n704), .ZN(new_n705));
  AOI21_X1  g519(.A(KEYINPUT104), .B1(new_n705), .B2(new_n348), .ZN(new_n706));
  INV_X1    g520(.A(new_n683), .ZN(new_n707));
  NOR2_X1   g521(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  INV_X1    g522(.A(new_n697), .ZN(new_n709));
  AND3_X1   g523(.A1(new_n632), .A2(new_n598), .A3(new_n709), .ZN(new_n710));
  NAND4_X1  g524(.A1(new_n708), .A2(new_n604), .A3(new_n671), .A4(new_n710), .ZN(new_n711));
  XNOR2_X1  g525(.A(new_n711), .B(G125), .ZN(G27));
  INV_X1    g526(.A(KEYINPUT107), .ZN(new_n713));
  NAND2_X1  g527(.A1(new_n343), .A2(new_n713), .ZN(new_n714));
  NAND2_X1  g528(.A1(new_n332), .A2(new_n317), .ZN(new_n715));
  INV_X1    g529(.A(KEYINPUT86), .ZN(new_n716));
  NAND2_X1  g530(.A1(new_n715), .A2(new_n716), .ZN(new_n717));
  NAND3_X1  g531(.A1(new_n717), .A2(new_n341), .A3(new_n191), .ZN(new_n718));
  NAND4_X1  g532(.A1(new_n718), .A2(KEYINPUT107), .A3(G469), .A4(new_n338), .ZN(new_n719));
  NAND2_X1  g533(.A1(new_n714), .A2(new_n719), .ZN(new_n720));
  NAND3_X1  g534(.A1(new_n337), .A2(new_n720), .A3(new_n344), .ZN(new_n721));
  NAND4_X1  g535(.A1(new_n396), .A2(new_n398), .A3(new_n402), .A4(new_n400), .ZN(new_n722));
  INV_X1    g536(.A(new_n348), .ZN(new_n723));
  NOR2_X1   g537(.A1(new_n722), .A2(new_n723), .ZN(new_n724));
  AND3_X1   g538(.A1(new_n721), .A2(new_n671), .A3(new_n724), .ZN(new_n725));
  AOI21_X1  g539(.A(new_n503), .B1(new_n518), .B2(new_n520), .ZN(new_n726));
  AOI211_X1 g540(.A(KEYINPUT108), .B(new_n451), .C1(new_n726), .C2(new_n499), .ZN(new_n727));
  INV_X1    g541(.A(KEYINPUT108), .ZN(new_n728));
  NAND2_X1  g542(.A1(new_n507), .A2(new_n508), .ZN(new_n729));
  NAND2_X1  g543(.A1(new_n729), .A2(new_n513), .ZN(new_n730));
  AOI21_X1  g544(.A(G902), .B1(new_n512), .B2(new_n514), .ZN(new_n731));
  NAND2_X1  g545(.A1(new_n730), .A2(new_n731), .ZN(new_n732));
  AOI21_X1  g546(.A(new_n519), .B1(new_n732), .B2(G472), .ZN(new_n733));
  INV_X1    g547(.A(new_n520), .ZN(new_n734));
  OAI211_X1 g548(.A(new_n501), .B(new_n499), .C1(new_n733), .C2(new_n734), .ZN(new_n735));
  AOI21_X1  g549(.A(new_n728), .B1(new_n735), .B2(new_n601), .ZN(new_n736));
  OAI211_X1 g550(.A(KEYINPUT42), .B(new_n725), .C1(new_n727), .C2(new_n736), .ZN(new_n737));
  INV_X1    g551(.A(KEYINPUT42), .ZN(new_n738));
  NAND4_X1  g552(.A1(new_n638), .A2(new_n601), .A3(new_n721), .A4(new_n724), .ZN(new_n739));
  INV_X1    g553(.A(new_n671), .ZN(new_n740));
  OAI21_X1  g554(.A(new_n738), .B1(new_n739), .B2(new_n740), .ZN(new_n741));
  NAND2_X1  g555(.A1(new_n737), .A2(new_n741), .ZN(new_n742));
  XNOR2_X1  g556(.A(new_n742), .B(G131), .ZN(G33));
  NAND4_X1  g557(.A1(new_n522), .A2(new_n644), .A3(new_n721), .A4(new_n724), .ZN(new_n744));
  XNOR2_X1  g558(.A(new_n744), .B(G134), .ZN(G36));
  NOR3_X1   g559(.A1(new_n557), .A2(new_n613), .A3(KEYINPUT43), .ZN(new_n746));
  XNOR2_X1  g560(.A(new_n556), .B(KEYINPUT111), .ZN(new_n747));
  OR2_X1    g561(.A1(new_n747), .A2(new_n613), .ZN(new_n748));
  AOI21_X1  g562(.A(new_n746), .B1(new_n748), .B2(KEYINPUT43), .ZN(new_n749));
  NAND4_X1  g563(.A1(new_n749), .A2(KEYINPUT44), .A3(new_n599), .A4(new_n632), .ZN(new_n750));
  INV_X1    g564(.A(KEYINPUT112), .ZN(new_n751));
  OR2_X1    g565(.A1(new_n750), .A2(new_n751), .ZN(new_n752));
  NAND3_X1  g566(.A1(new_n749), .A2(new_n599), .A3(new_n632), .ZN(new_n753));
  INV_X1    g567(.A(KEYINPUT44), .ZN(new_n754));
  AOI21_X1  g568(.A(new_n722), .B1(new_n753), .B2(new_n754), .ZN(new_n755));
  NAND2_X1  g569(.A1(new_n750), .A2(new_n751), .ZN(new_n756));
  NAND3_X1  g570(.A1(new_n752), .A2(new_n755), .A3(new_n756), .ZN(new_n757));
  OR2_X1    g571(.A1(new_n757), .A2(KEYINPUT113), .ZN(new_n758));
  NAND2_X1  g572(.A1(new_n757), .A2(KEYINPUT113), .ZN(new_n759));
  NAND2_X1  g573(.A1(new_n718), .A2(new_n338), .ZN(new_n760));
  XNOR2_X1  g574(.A(new_n760), .B(KEYINPUT45), .ZN(new_n761));
  NAND2_X1  g575(.A1(new_n761), .A2(G469), .ZN(new_n762));
  XNOR2_X1  g576(.A(new_n762), .B(KEYINPUT109), .ZN(new_n763));
  NAND2_X1  g577(.A1(new_n763), .A2(new_n344), .ZN(new_n764));
  INV_X1    g578(.A(KEYINPUT46), .ZN(new_n765));
  OR3_X1    g579(.A1(new_n764), .A2(KEYINPUT110), .A3(new_n765), .ZN(new_n766));
  AOI21_X1  g580(.A(new_n703), .B1(new_n764), .B2(new_n765), .ZN(new_n767));
  OAI21_X1  g581(.A(KEYINPUT110), .B1(new_n764), .B2(new_n765), .ZN(new_n768));
  NAND3_X1  g582(.A1(new_n766), .A2(new_n767), .A3(new_n768), .ZN(new_n769));
  AND2_X1   g583(.A1(new_n769), .A2(new_n348), .ZN(new_n770));
  NAND4_X1  g584(.A1(new_n758), .A2(new_n655), .A3(new_n759), .A4(new_n770), .ZN(new_n771));
  XNOR2_X1  g585(.A(new_n771), .B(G137), .ZN(G39));
  INV_X1    g586(.A(KEYINPUT47), .ZN(new_n773));
  AOI22_X1  g587(.A1(new_n769), .A2(new_n348), .B1(KEYINPUT114), .B2(new_n773), .ZN(new_n774));
  XOR2_X1   g588(.A(KEYINPUT114), .B(KEYINPUT47), .Z(new_n775));
  AOI21_X1  g589(.A(new_n774), .B1(new_n770), .B2(new_n775), .ZN(new_n776));
  INV_X1    g590(.A(new_n722), .ZN(new_n777));
  NOR2_X1   g591(.A1(new_n638), .A2(new_n601), .ZN(new_n778));
  NAND4_X1  g592(.A1(new_n776), .A2(new_n671), .A3(new_n777), .A4(new_n778), .ZN(new_n779));
  XNOR2_X1  g593(.A(new_n779), .B(KEYINPUT115), .ZN(new_n780));
  XNOR2_X1  g594(.A(new_n780), .B(new_n414), .ZN(G42));
  AND2_X1   g595(.A1(new_n749), .A2(new_n405), .ZN(new_n782));
  AND2_X1   g596(.A1(new_n782), .A2(new_n698), .ZN(new_n783));
  NOR3_X1   g597(.A1(new_n703), .A2(new_n704), .A3(new_n348), .ZN(new_n784));
  OAI211_X1 g598(.A(new_n777), .B(new_n783), .C1(new_n776), .C2(new_n784), .ZN(new_n785));
  INV_X1    g599(.A(KEYINPUT51), .ZN(new_n786));
  NOR3_X1   g600(.A1(new_n706), .A2(new_n707), .A3(new_n722), .ZN(new_n787));
  AND3_X1   g601(.A1(new_n782), .A2(new_n710), .A3(new_n787), .ZN(new_n788));
  NOR2_X1   g602(.A1(new_n668), .A2(new_n402), .ZN(new_n789));
  NAND3_X1  g603(.A1(new_n783), .A2(new_n708), .A3(new_n789), .ZN(new_n790));
  AOI21_X1  g604(.A(new_n788), .B1(new_n790), .B2(KEYINPUT50), .ZN(new_n791));
  INV_X1    g605(.A(KEYINPUT50), .ZN(new_n792));
  NAND4_X1  g606(.A1(new_n783), .A2(new_n792), .A3(new_n708), .A4(new_n789), .ZN(new_n793));
  AND4_X1   g607(.A1(new_n601), .A2(new_n787), .A3(new_n405), .A4(new_n665), .ZN(new_n794));
  NAND3_X1  g608(.A1(new_n794), .A2(new_n556), .A3(new_n613), .ZN(new_n795));
  NAND3_X1  g609(.A1(new_n791), .A2(new_n793), .A3(new_n795), .ZN(new_n796));
  OAI21_X1  g610(.A(new_n786), .B1(new_n796), .B2(KEYINPUT120), .ZN(new_n797));
  INV_X1    g611(.A(new_n796), .ZN(new_n798));
  AND3_X1   g612(.A1(new_n785), .A2(new_n797), .A3(new_n798), .ZN(new_n799));
  AOI21_X1  g613(.A(new_n797), .B1(new_n785), .B2(new_n798), .ZN(new_n800));
  NOR2_X1   g614(.A1(new_n799), .A2(new_n800), .ZN(new_n801));
  AOI21_X1  g615(.A(new_n673), .B1(new_n646), .B2(new_n651), .ZN(new_n802));
  NAND2_X1  g616(.A1(new_n699), .A2(new_n604), .ZN(new_n803));
  NOR2_X1   g617(.A1(new_n803), .A2(new_n641), .ZN(new_n804));
  AND2_X1   g618(.A1(new_n721), .A2(new_n649), .ZN(new_n805));
  NAND4_X1  g619(.A1(new_n804), .A2(new_n348), .A3(new_n664), .A4(new_n805), .ZN(new_n806));
  NAND3_X1  g620(.A1(new_n802), .A2(new_n711), .A3(new_n806), .ZN(new_n807));
  INV_X1    g621(.A(KEYINPUT52), .ZN(new_n808));
  NAND2_X1  g622(.A1(new_n807), .A2(new_n808), .ZN(new_n809));
  NAND4_X1  g623(.A1(new_n802), .A2(new_n711), .A3(new_n806), .A4(KEYINPUT52), .ZN(new_n810));
  NAND2_X1  g624(.A1(new_n809), .A2(new_n810), .ZN(new_n811));
  INV_X1    g625(.A(new_n693), .ZN(new_n812));
  NAND4_X1  g626(.A1(new_n686), .A2(new_n689), .A3(new_n701), .A4(new_n812), .ZN(new_n813));
  INV_X1    g627(.A(new_n411), .ZN(new_n814));
  NAND2_X1  g628(.A1(new_n556), .A2(new_n593), .ZN(new_n815));
  OAI21_X1  g629(.A(new_n815), .B1(new_n556), .B2(new_n613), .ZN(new_n816));
  NAND4_X1  g630(.A1(new_n600), .A2(new_n601), .A3(new_n814), .A4(new_n816), .ZN(new_n817));
  NAND3_X1  g631(.A1(new_n633), .A2(new_n817), .A3(new_n595), .ZN(new_n818));
  NOR2_X1   g632(.A1(new_n813), .A2(new_n818), .ZN(new_n819));
  NAND4_X1  g633(.A1(new_n710), .A2(new_n721), .A3(new_n671), .A4(new_n724), .ZN(new_n820));
  AND2_X1   g634(.A1(new_n777), .A2(new_n642), .ZN(new_n821));
  NAND3_X1  g635(.A1(new_n638), .A2(new_n620), .A3(new_n821), .ZN(new_n822));
  NOR2_X1   g636(.A1(new_n649), .A2(new_n593), .ZN(new_n823));
  NAND3_X1  g637(.A1(new_n345), .A2(new_n348), .A3(new_n823), .ZN(new_n824));
  OAI21_X1  g638(.A(new_n820), .B1(new_n822), .B2(new_n824), .ZN(new_n825));
  NAND2_X1  g639(.A1(new_n721), .A2(new_n724), .ZN(new_n826));
  AOI22_X1  g640(.A1(new_n502), .A2(new_n505), .B1(new_n520), .B2(new_n518), .ZN(new_n827));
  NOR4_X1   g641(.A1(new_n826), .A2(new_n827), .A3(new_n451), .A4(new_n643), .ZN(new_n828));
  OAI21_X1  g642(.A(KEYINPUT116), .B1(new_n825), .B2(new_n828), .ZN(new_n829));
  NAND2_X1  g643(.A1(new_n777), .A2(new_n642), .ZN(new_n830));
  AOI21_X1  g644(.A(new_n830), .B1(new_n521), .B2(new_n506), .ZN(new_n831));
  NAND4_X1  g645(.A1(new_n654), .A2(new_n831), .A3(new_n620), .A4(new_n823), .ZN(new_n832));
  INV_X1    g646(.A(KEYINPUT116), .ZN(new_n833));
  NAND4_X1  g647(.A1(new_n832), .A2(new_n833), .A3(new_n744), .A4(new_n820), .ZN(new_n834));
  AND3_X1   g648(.A1(new_n829), .A2(new_n742), .A3(new_n834), .ZN(new_n835));
  AOI21_X1  g649(.A(KEYINPUT117), .B1(new_n819), .B2(new_n835), .ZN(new_n836));
  NAND3_X1  g650(.A1(new_n829), .A2(new_n742), .A3(new_n834), .ZN(new_n837));
  INV_X1    g651(.A(KEYINPUT117), .ZN(new_n838));
  NOR4_X1   g652(.A1(new_n813), .A2(new_n837), .A3(new_n838), .A4(new_n818), .ZN(new_n839));
  OAI21_X1  g653(.A(new_n811), .B1(new_n836), .B2(new_n839), .ZN(new_n840));
  INV_X1    g654(.A(KEYINPUT53), .ZN(new_n841));
  NOR2_X1   g655(.A1(new_n840), .A2(new_n841), .ZN(new_n842));
  AND2_X1   g656(.A1(new_n686), .A2(new_n701), .ZN(new_n843));
  INV_X1    g657(.A(new_n522), .ZN(new_n844));
  INV_X1    g658(.A(KEYINPUT105), .ZN(new_n845));
  OAI21_X1  g659(.A(new_n845), .B1(new_n706), .B2(new_n707), .ZN(new_n846));
  NAND3_X1  g660(.A1(new_n682), .A2(KEYINPUT105), .A3(new_n683), .ZN(new_n847));
  AOI21_X1  g661(.A(new_n844), .B1(new_n846), .B2(new_n847), .ZN(new_n848));
  AOI21_X1  g662(.A(new_n693), .B1(new_n848), .B2(new_n622), .ZN(new_n849));
  INV_X1    g663(.A(new_n818), .ZN(new_n850));
  NAND4_X1  g664(.A1(new_n843), .A2(new_n835), .A3(new_n849), .A4(new_n850), .ZN(new_n851));
  NAND2_X1  g665(.A1(new_n851), .A2(new_n838), .ZN(new_n852));
  AND4_X1   g666(.A1(new_n686), .A2(new_n689), .A3(new_n701), .A4(new_n812), .ZN(new_n853));
  NAND4_X1  g667(.A1(new_n853), .A2(KEYINPUT117), .A3(new_n850), .A4(new_n835), .ZN(new_n854));
  NAND2_X1  g668(.A1(new_n852), .A2(new_n854), .ZN(new_n855));
  AOI21_X1  g669(.A(KEYINPUT53), .B1(new_n855), .B2(new_n811), .ZN(new_n856));
  OAI21_X1  g670(.A(KEYINPUT54), .B1(new_n842), .B2(new_n856), .ZN(new_n857));
  NAND2_X1  g671(.A1(new_n840), .A2(new_n841), .ZN(new_n858));
  NAND4_X1  g672(.A1(new_n853), .A2(KEYINPUT53), .A3(new_n850), .A4(new_n835), .ZN(new_n859));
  AND2_X1   g673(.A1(new_n809), .A2(new_n810), .ZN(new_n860));
  INV_X1    g674(.A(KEYINPUT118), .ZN(new_n861));
  NOR3_X1   g675(.A1(new_n859), .A2(new_n860), .A3(new_n861), .ZN(new_n862));
  NOR4_X1   g676(.A1(new_n813), .A2(new_n837), .A3(new_n841), .A4(new_n818), .ZN(new_n863));
  AOI21_X1  g677(.A(KEYINPUT118), .B1(new_n863), .B2(new_n811), .ZN(new_n864));
  NOR2_X1   g678(.A1(new_n862), .A2(new_n864), .ZN(new_n865));
  XNOR2_X1  g679(.A(KEYINPUT119), .B(KEYINPUT54), .ZN(new_n866));
  INV_X1    g680(.A(new_n866), .ZN(new_n867));
  NAND3_X1  g681(.A1(new_n858), .A2(new_n865), .A3(new_n867), .ZN(new_n868));
  NAND2_X1  g682(.A1(new_n782), .A2(new_n787), .ZN(new_n869));
  NOR2_X1   g683(.A1(new_n727), .A2(new_n736), .ZN(new_n870));
  NOR2_X1   g684(.A1(new_n869), .A2(new_n870), .ZN(new_n871));
  XOR2_X1   g685(.A(new_n871), .B(KEYINPUT48), .Z(new_n872));
  NAND3_X1  g686(.A1(new_n783), .A2(new_n604), .A3(new_n708), .ZN(new_n873));
  NAND2_X1  g687(.A1(new_n794), .A2(new_n614), .ZN(new_n874));
  XOR2_X1   g688(.A(new_n404), .B(KEYINPUT121), .Z(new_n875));
  NAND4_X1  g689(.A1(new_n872), .A2(new_n873), .A3(new_n874), .A4(new_n875), .ZN(new_n876));
  XNOR2_X1  g690(.A(new_n876), .B(KEYINPUT122), .ZN(new_n877));
  NAND4_X1  g691(.A1(new_n801), .A2(new_n857), .A3(new_n868), .A4(new_n877), .ZN(new_n878));
  OAI21_X1  g692(.A(new_n878), .B1(G952), .B2(G953), .ZN(new_n879));
  NOR4_X1   g693(.A1(new_n668), .A2(new_n723), .A3(new_n603), .A4(new_n664), .ZN(new_n880));
  INV_X1    g694(.A(new_n748), .ZN(new_n881));
  XNOR2_X1  g695(.A(new_n705), .B(KEYINPUT49), .ZN(new_n882));
  NAND4_X1  g696(.A1(new_n880), .A2(new_n601), .A3(new_n881), .A4(new_n882), .ZN(new_n883));
  NAND2_X1  g697(.A1(new_n879), .A2(new_n883), .ZN(G75));
  NAND2_X1  g698(.A1(new_n377), .A2(new_n379), .ZN(new_n885));
  XNOR2_X1  g699(.A(new_n885), .B(new_n358), .ZN(new_n886));
  XOR2_X1   g700(.A(new_n886), .B(KEYINPUT55), .Z(new_n887));
  OAI21_X1  g701(.A(new_n861), .B1(new_n859), .B2(new_n860), .ZN(new_n888));
  NAND3_X1  g702(.A1(new_n863), .A2(KEYINPUT118), .A3(new_n811), .ZN(new_n889));
  NAND2_X1  g703(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  OAI211_X1 g704(.A(G210), .B(G902), .C1(new_n856), .C2(new_n890), .ZN(new_n891));
  INV_X1    g705(.A(new_n891), .ZN(new_n892));
  OAI21_X1  g706(.A(new_n887), .B1(new_n892), .B2(KEYINPUT56), .ZN(new_n893));
  NOR2_X1   g707(.A1(new_n403), .A2(G952), .ZN(new_n894));
  INV_X1    g708(.A(new_n894), .ZN(new_n895));
  XNOR2_X1  g709(.A(KEYINPUT123), .B(KEYINPUT56), .ZN(new_n896));
  NOR2_X1   g710(.A1(new_n887), .A2(new_n896), .ZN(new_n897));
  NAND2_X1  g711(.A1(new_n891), .A2(new_n897), .ZN(new_n898));
  NAND3_X1  g712(.A1(new_n893), .A2(new_n895), .A3(new_n898), .ZN(new_n899));
  NAND2_X1  g713(.A1(new_n899), .A2(KEYINPUT124), .ZN(new_n900));
  INV_X1    g714(.A(KEYINPUT124), .ZN(new_n901));
  NAND4_X1  g715(.A1(new_n893), .A2(new_n901), .A3(new_n895), .A4(new_n898), .ZN(new_n902));
  NAND2_X1  g716(.A1(new_n900), .A2(new_n902), .ZN(G51));
  OAI21_X1  g717(.A(new_n866), .B1(new_n856), .B2(new_n890), .ZN(new_n904));
  NAND3_X1  g718(.A1(new_n868), .A2(new_n904), .A3(KEYINPUT125), .ZN(new_n905));
  NOR2_X1   g719(.A1(new_n856), .A2(new_n890), .ZN(new_n906));
  INV_X1    g720(.A(KEYINPUT125), .ZN(new_n907));
  NAND3_X1  g721(.A1(new_n906), .A2(new_n907), .A3(new_n867), .ZN(new_n908));
  XOR2_X1   g722(.A(new_n344), .B(KEYINPUT57), .Z(new_n909));
  NAND3_X1  g723(.A1(new_n905), .A2(new_n908), .A3(new_n909), .ZN(new_n910));
  NAND2_X1  g724(.A1(new_n910), .A2(new_n334), .ZN(new_n911));
  OR3_X1    g725(.A1(new_n906), .A2(new_n336), .A3(new_n763), .ZN(new_n912));
  AOI21_X1  g726(.A(new_n894), .B1(new_n911), .B2(new_n912), .ZN(G54));
  NAND2_X1  g727(.A1(new_n858), .A2(new_n865), .ZN(new_n914));
  NAND4_X1  g728(.A1(new_n914), .A2(KEYINPUT58), .A3(G475), .A4(G902), .ZN(new_n915));
  INV_X1    g729(.A(new_n547), .ZN(new_n916));
  AND2_X1   g730(.A1(new_n915), .A2(new_n916), .ZN(new_n917));
  NOR2_X1   g731(.A1(new_n915), .A2(new_n916), .ZN(new_n918));
  NOR3_X1   g732(.A1(new_n917), .A2(new_n918), .A3(new_n894), .ZN(G60));
  XNOR2_X1  g733(.A(new_n607), .B(KEYINPUT59), .ZN(new_n920));
  AND2_X1   g734(.A1(new_n612), .A2(new_n920), .ZN(new_n921));
  NAND3_X1  g735(.A1(new_n905), .A2(new_n908), .A3(new_n921), .ZN(new_n922));
  INV_X1    g736(.A(KEYINPUT126), .ZN(new_n923));
  AND3_X1   g737(.A1(new_n922), .A2(new_n923), .A3(new_n895), .ZN(new_n924));
  AOI21_X1  g738(.A(new_n923), .B1(new_n922), .B2(new_n895), .ZN(new_n925));
  NAND2_X1  g739(.A1(new_n857), .A2(new_n868), .ZN(new_n926));
  AOI21_X1  g740(.A(new_n612), .B1(new_n926), .B2(new_n920), .ZN(new_n927));
  NOR3_X1   g741(.A1(new_n924), .A2(new_n925), .A3(new_n927), .ZN(G63));
  NAND2_X1  g742(.A1(G217), .A2(G902), .ZN(new_n929));
  XOR2_X1   g743(.A(new_n929), .B(KEYINPUT60), .Z(new_n930));
  NAND3_X1  g744(.A1(new_n914), .A2(new_n629), .A3(new_n930), .ZN(new_n931));
  AND2_X1   g745(.A1(new_n914), .A2(new_n930), .ZN(new_n932));
  OAI211_X1 g746(.A(new_n895), .B(new_n931), .C1(new_n932), .C2(new_n443), .ZN(new_n933));
  INV_X1    g747(.A(KEYINPUT127), .ZN(new_n934));
  AOI21_X1  g748(.A(KEYINPUT61), .B1(new_n931), .B2(new_n934), .ZN(new_n935));
  XNOR2_X1  g749(.A(new_n933), .B(new_n935), .ZN(G66));
  INV_X1    g750(.A(new_n409), .ZN(new_n937));
  OAI21_X1  g751(.A(G953), .B1(new_n937), .B2(new_n356), .ZN(new_n938));
  OAI21_X1  g752(.A(new_n938), .B1(new_n819), .B2(G953), .ZN(new_n939));
  OAI21_X1  g753(.A(new_n885), .B1(G898), .B2(new_n403), .ZN(new_n940));
  XNOR2_X1  g754(.A(new_n939), .B(new_n940), .ZN(G69));
  NAND2_X1  g755(.A1(new_n522), .A2(new_n816), .ZN(new_n942));
  NOR3_X1   g756(.A1(new_n656), .A2(new_n942), .A3(new_n722), .ZN(new_n943));
  AND2_X1   g757(.A1(new_n802), .A2(new_n711), .ZN(new_n944));
  AND2_X1   g758(.A1(new_n669), .A2(new_n944), .ZN(new_n945));
  OR2_X1    g759(.A1(new_n945), .A2(KEYINPUT62), .ZN(new_n946));
  NAND2_X1  g760(.A1(new_n945), .A2(KEYINPUT62), .ZN(new_n947));
  AOI21_X1  g761(.A(new_n943), .B1(new_n946), .B2(new_n947), .ZN(new_n948));
  NAND3_X1  g762(.A1(new_n779), .A2(new_n771), .A3(new_n948), .ZN(new_n949));
  NAND2_X1  g763(.A1(new_n463), .A2(new_n472), .ZN(new_n950));
  XNOR2_X1  g764(.A(new_n950), .B(new_n535), .ZN(new_n951));
  NAND3_X1  g765(.A1(new_n949), .A2(new_n403), .A3(new_n951), .ZN(new_n952));
  INV_X1    g766(.A(G900), .ZN(new_n953));
  AOI21_X1  g767(.A(new_n953), .B1(new_n951), .B2(new_n188), .ZN(new_n954));
  NAND3_X1  g768(.A1(new_n779), .A2(new_n771), .A3(new_n944), .ZN(new_n955));
  NAND2_X1  g769(.A1(new_n770), .A2(new_n655), .ZN(new_n956));
  NOR3_X1   g770(.A1(new_n956), .A2(new_n803), .A3(new_n870), .ZN(new_n957));
  NOR3_X1   g771(.A1(new_n955), .A2(G953), .A3(new_n957), .ZN(new_n958));
  NAND2_X1  g772(.A1(new_n742), .A2(new_n744), .ZN(new_n959));
  INV_X1    g773(.A(new_n959), .ZN(new_n960));
  AOI22_X1  g774(.A1(new_n958), .A2(new_n960), .B1(G227), .B2(G953), .ZN(new_n961));
  OAI221_X1 g775(.A(new_n952), .B1(new_n403), .B2(new_n954), .C1(new_n961), .C2(new_n951), .ZN(G72));
  NAND2_X1  g776(.A1(G472), .A2(G902), .ZN(new_n963));
  XOR2_X1   g777(.A(new_n963), .B(KEYINPUT63), .Z(new_n964));
  INV_X1    g778(.A(new_n819), .ZN(new_n965));
  OAI21_X1  g779(.A(new_n964), .B1(new_n949), .B2(new_n965), .ZN(new_n966));
  AOI21_X1  g780(.A(new_n894), .B1(new_n966), .B2(new_n661), .ZN(new_n967));
  OAI211_X1 g781(.A(new_n508), .B(new_n964), .C1(new_n842), .C2(new_n856), .ZN(new_n968));
  INV_X1    g782(.A(new_n964), .ZN(new_n969));
  NOR2_X1   g783(.A1(new_n955), .A2(new_n957), .ZN(new_n970));
  NOR2_X1   g784(.A1(new_n965), .A2(new_n959), .ZN(new_n971));
  AOI21_X1  g785(.A(new_n969), .B1(new_n970), .B2(new_n971), .ZN(new_n972));
  OAI221_X1 g786(.A(new_n967), .B1(new_n661), .B2(new_n968), .C1(new_n972), .C2(new_n508), .ZN(new_n973));
  INV_X1    g787(.A(new_n973), .ZN(G57));
endmodule


