//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 1 1 1 0 1 1 0 1 0 0 0 0 0 0 1 0 1 1 0 1 1 0 0 0 1 1 1 0 1 1 0 1 1 1 1 0 1 0 0 0 0 0 1 1 1 1 0 1 0 0 1 0 0 1 0 0 1 1 1 1 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:35:43 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n203, new_n204, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n227, new_n228, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n236, new_n237, new_n238, new_n239,
    new_n240, new_n241, new_n242, new_n244, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n692, new_n693, new_n694, new_n695, new_n696,
    new_n697, new_n698, new_n699, new_n700, new_n701, new_n702, new_n703,
    new_n704, new_n705, new_n706, new_n707, new_n708, new_n709, new_n710,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n772, new_n773, new_n774, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1108, new_n1109, new_n1110, new_n1111, new_n1112,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1186, new_n1187, new_n1188, new_n1189, new_n1190, new_n1191,
    new_n1192, new_n1193, new_n1194, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1251, new_n1252,
    new_n1253, new_n1254, new_n1255, new_n1256, new_n1257, new_n1258,
    new_n1260, new_n1261, new_n1262, new_n1263, new_n1264, new_n1265,
    new_n1266, new_n1267, new_n1268, new_n1269, new_n1270, new_n1271,
    new_n1272, new_n1273, new_n1274, new_n1275, new_n1276, new_n1277,
    new_n1278, new_n1279, new_n1280, new_n1281, new_n1283, new_n1284,
    new_n1285, new_n1286, new_n1287, new_n1288, new_n1289, new_n1290,
    new_n1291, new_n1292, new_n1293, new_n1294, new_n1295, new_n1296,
    new_n1298, new_n1299, new_n1300, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1346,
    new_n1347, new_n1348, new_n1349, new_n1350, new_n1351, new_n1352,
    new_n1353, new_n1354, new_n1355, new_n1356, new_n1357, new_n1358,
    new_n1359, new_n1360, new_n1361, new_n1362, new_n1363, new_n1364,
    new_n1365, new_n1366, new_n1367, new_n1368, new_n1369, new_n1370,
    new_n1371, new_n1372, new_n1373, new_n1374, new_n1376, new_n1377,
    new_n1378, new_n1379, new_n1380, new_n1381;
  NOR4_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .A4(G77), .ZN(G353));
  OAI21_X1  g0001(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0002(.A1(G1), .A2(G20), .ZN(new_n203));
  AOI22_X1  g0003(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n204));
  XOR2_X1   g0004(.A(new_n204), .B(KEYINPUT66), .Z(new_n205));
  AOI22_X1  g0005(.A1(G58), .A2(G232), .B1(G116), .B2(G270), .ZN(new_n206));
  AOI22_X1  g0006(.A1(G50), .A2(G226), .B1(G68), .B2(G238), .ZN(new_n207));
  AOI22_X1  g0007(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n208));
  NAND3_X1  g0008(.A1(new_n206), .A2(new_n207), .A3(new_n208), .ZN(new_n209));
  OAI21_X1  g0009(.A(new_n203), .B1(new_n205), .B2(new_n209), .ZN(new_n210));
  XOR2_X1   g0010(.A(new_n210), .B(KEYINPUT67), .Z(new_n211));
  INV_X1    g0011(.A(KEYINPUT1), .ZN(new_n212));
  OR2_X1    g0012(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  NAND2_X1  g0013(.A1(new_n211), .A2(new_n212), .ZN(new_n214));
  OR3_X1    g0014(.A1(new_n203), .A2(KEYINPUT64), .A3(G13), .ZN(new_n215));
  OAI21_X1  g0015(.A(KEYINPUT64), .B1(new_n203), .B2(G13), .ZN(new_n216));
  NAND2_X1  g0016(.A1(new_n215), .A2(new_n216), .ZN(new_n217));
  OAI211_X1 g0017(.A(new_n217), .B(G250), .C1(G257), .C2(G264), .ZN(new_n218));
  XOR2_X1   g0018(.A(new_n218), .B(KEYINPUT0), .Z(new_n219));
  NAND2_X1  g0019(.A1(G1), .A2(G13), .ZN(new_n220));
  INV_X1    g0020(.A(G20), .ZN(new_n221));
  NOR2_X1   g0021(.A1(new_n220), .A2(new_n221), .ZN(new_n222));
  OAI21_X1  g0022(.A(G50), .B1(G58), .B2(G68), .ZN(new_n223));
  XOR2_X1   g0023(.A(new_n223), .B(KEYINPUT65), .Z(new_n224));
  AOI21_X1  g0024(.A(new_n219), .B1(new_n222), .B2(new_n224), .ZN(new_n225));
  AND3_X1   g0025(.A1(new_n213), .A2(new_n214), .A3(new_n225), .ZN(G361));
  XNOR2_X1  g0026(.A(G238), .B(G244), .ZN(new_n227));
  INV_X1    g0027(.A(G232), .ZN(new_n228));
  XNOR2_X1  g0028(.A(new_n227), .B(new_n228), .ZN(new_n229));
  XNOR2_X1  g0029(.A(KEYINPUT2), .B(G226), .ZN(new_n230));
  XNOR2_X1  g0030(.A(new_n229), .B(new_n230), .ZN(new_n231));
  XNOR2_X1  g0031(.A(G250), .B(G257), .ZN(new_n232));
  XNOR2_X1  g0032(.A(G264), .B(G270), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n232), .B(new_n233), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n231), .B(new_n234), .ZN(G358));
  XOR2_X1   g0035(.A(G87), .B(G97), .Z(new_n236));
  XNOR2_X1  g0036(.A(new_n236), .B(KEYINPUT68), .ZN(new_n237));
  XNOR2_X1  g0037(.A(G107), .B(G116), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XNOR2_X1  g0039(.A(G50), .B(G68), .ZN(new_n240));
  XNOR2_X1  g0040(.A(G58), .B(G77), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XOR2_X1   g0042(.A(new_n239), .B(new_n242), .Z(G351));
  NAND3_X1  g0043(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n244));
  NAND2_X1  g0044(.A1(new_n244), .A2(new_n220), .ZN(new_n245));
  XNOR2_X1  g0045(.A(KEYINPUT8), .B(G58), .ZN(new_n246));
  NAND2_X1  g0046(.A1(new_n221), .A2(G33), .ZN(new_n247));
  INV_X1    g0047(.A(G150), .ZN(new_n248));
  NOR2_X1   g0048(.A1(G20), .A2(G33), .ZN(new_n249));
  INV_X1    g0049(.A(new_n249), .ZN(new_n250));
  OAI22_X1  g0050(.A1(new_n246), .A2(new_n247), .B1(new_n248), .B2(new_n250), .ZN(new_n251));
  NOR2_X1   g0051(.A1(G58), .A2(G68), .ZN(new_n252));
  INV_X1    g0052(.A(G50), .ZN(new_n253));
  AOI21_X1  g0053(.A(new_n221), .B1(new_n252), .B2(new_n253), .ZN(new_n254));
  OAI21_X1  g0054(.A(new_n245), .B1(new_n251), .B2(new_n254), .ZN(new_n255));
  INV_X1    g0055(.A(G1), .ZN(new_n256));
  NAND3_X1  g0056(.A1(new_n256), .A2(G13), .A3(G20), .ZN(new_n257));
  INV_X1    g0057(.A(new_n257), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n258), .A2(new_n253), .ZN(new_n259));
  NAND3_X1  g0059(.A1(new_n257), .A2(new_n220), .A3(new_n244), .ZN(new_n260));
  INV_X1    g0060(.A(new_n260), .ZN(new_n261));
  INV_X1    g0061(.A(KEYINPUT69), .ZN(new_n262));
  NAND2_X1  g0062(.A1(new_n256), .A2(G20), .ZN(new_n263));
  INV_X1    g0063(.A(new_n263), .ZN(new_n264));
  OAI21_X1  g0064(.A(new_n262), .B1(new_n264), .B2(new_n253), .ZN(new_n265));
  NAND3_X1  g0065(.A1(new_n263), .A2(KEYINPUT69), .A3(G50), .ZN(new_n266));
  NAND3_X1  g0066(.A1(new_n261), .A2(new_n265), .A3(new_n266), .ZN(new_n267));
  NAND3_X1  g0067(.A1(new_n255), .A2(new_n259), .A3(new_n267), .ZN(new_n268));
  INV_X1    g0068(.A(KEYINPUT9), .ZN(new_n269));
  OR2_X1    g0069(.A1(new_n268), .A2(new_n269), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n268), .A2(new_n269), .ZN(new_n271));
  NAND2_X1  g0071(.A1(G33), .A2(G41), .ZN(new_n272));
  NAND3_X1  g0072(.A1(new_n272), .A2(G1), .A3(G13), .ZN(new_n273));
  OR2_X1    g0073(.A1(G41), .A2(G45), .ZN(new_n274));
  NAND4_X1  g0074(.A1(new_n273), .A2(new_n256), .A3(G274), .A4(new_n274), .ZN(new_n275));
  INV_X1    g0075(.A(new_n275), .ZN(new_n276));
  OAI21_X1  g0076(.A(new_n256), .B1(G41), .B2(G45), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n273), .A2(new_n277), .ZN(new_n278));
  INV_X1    g0078(.A(new_n278), .ZN(new_n279));
  AOI21_X1  g0079(.A(new_n276), .B1(G226), .B2(new_n279), .ZN(new_n280));
  XNOR2_X1  g0080(.A(KEYINPUT3), .B(G33), .ZN(new_n281));
  NOR2_X1   g0081(.A1(G222), .A2(G1698), .ZN(new_n282));
  INV_X1    g0082(.A(G1698), .ZN(new_n283));
  NOR2_X1   g0083(.A1(new_n283), .A2(G223), .ZN(new_n284));
  OAI21_X1  g0084(.A(new_n281), .B1(new_n282), .B2(new_n284), .ZN(new_n285));
  INV_X1    g0085(.A(new_n273), .ZN(new_n286));
  OAI211_X1 g0086(.A(new_n285), .B(new_n286), .C1(G77), .C2(new_n281), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n280), .A2(new_n287), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n288), .A2(G200), .ZN(new_n289));
  NAND3_X1  g0089(.A1(new_n280), .A2(G190), .A3(new_n287), .ZN(new_n290));
  NAND4_X1  g0090(.A1(new_n270), .A2(new_n271), .A3(new_n289), .A4(new_n290), .ZN(new_n291));
  XNOR2_X1  g0091(.A(new_n291), .B(KEYINPUT10), .ZN(new_n292));
  INV_X1    g0092(.A(KEYINPUT72), .ZN(new_n293));
  INV_X1    g0093(.A(G77), .ZN(new_n294));
  AOI21_X1  g0094(.A(new_n294), .B1(new_n256), .B2(G20), .ZN(new_n295));
  INV_X1    g0095(.A(new_n295), .ZN(new_n296));
  OAI21_X1  g0096(.A(KEYINPUT71), .B1(new_n260), .B2(new_n296), .ZN(new_n297));
  INV_X1    g0097(.A(new_n245), .ZN(new_n298));
  INV_X1    g0098(.A(KEYINPUT71), .ZN(new_n299));
  NAND4_X1  g0099(.A1(new_n298), .A2(new_n299), .A3(new_n257), .A4(new_n295), .ZN(new_n300));
  AOI22_X1  g0100(.A1(new_n297), .A2(new_n300), .B1(new_n294), .B2(new_n258), .ZN(new_n301));
  INV_X1    g0101(.A(G58), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n302), .A2(KEYINPUT8), .ZN(new_n303));
  INV_X1    g0103(.A(KEYINPUT8), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n304), .A2(G58), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n303), .A2(new_n305), .ZN(new_n306));
  AOI22_X1  g0106(.A1(new_n306), .A2(new_n249), .B1(G20), .B2(G77), .ZN(new_n307));
  INV_X1    g0107(.A(new_n247), .ZN(new_n308));
  INV_X1    g0108(.A(G87), .ZN(new_n309));
  AND2_X1   g0109(.A1(new_n309), .A2(KEYINPUT15), .ZN(new_n310));
  NOR2_X1   g0110(.A1(new_n309), .A2(KEYINPUT15), .ZN(new_n311));
  OAI21_X1  g0111(.A(new_n308), .B1(new_n310), .B2(new_n311), .ZN(new_n312));
  AOI211_X1 g0112(.A(KEYINPUT70), .B(new_n298), .C1(new_n307), .C2(new_n312), .ZN(new_n313));
  INV_X1    g0113(.A(KEYINPUT70), .ZN(new_n314));
  NOR2_X1   g0114(.A1(new_n304), .A2(G58), .ZN(new_n315));
  NOR2_X1   g0115(.A1(new_n302), .A2(KEYINPUT8), .ZN(new_n316));
  OAI21_X1  g0116(.A(new_n249), .B1(new_n315), .B2(new_n316), .ZN(new_n317));
  NAND2_X1  g0117(.A1(G20), .A2(G77), .ZN(new_n318));
  NAND3_X1  g0118(.A1(new_n312), .A2(new_n317), .A3(new_n318), .ZN(new_n319));
  AOI21_X1  g0119(.A(new_n314), .B1(new_n319), .B2(new_n245), .ZN(new_n320));
  OAI21_X1  g0120(.A(new_n301), .B1(new_n313), .B2(new_n320), .ZN(new_n321));
  INV_X1    g0121(.A(G200), .ZN(new_n322));
  NAND3_X1  g0122(.A1(new_n281), .A2(G232), .A3(new_n283), .ZN(new_n323));
  INV_X1    g0123(.A(G33), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n324), .A2(KEYINPUT3), .ZN(new_n325));
  INV_X1    g0125(.A(KEYINPUT3), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n326), .A2(G33), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n325), .A2(new_n327), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n328), .A2(G107), .ZN(new_n329));
  INV_X1    g0129(.A(G238), .ZN(new_n330));
  NOR2_X1   g0130(.A1(new_n330), .A2(new_n283), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n281), .A2(new_n331), .ZN(new_n332));
  NAND3_X1  g0132(.A1(new_n323), .A2(new_n329), .A3(new_n332), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n333), .A2(new_n286), .ZN(new_n334));
  INV_X1    g0134(.A(G244), .ZN(new_n335));
  OAI21_X1  g0135(.A(new_n275), .B1(new_n335), .B2(new_n278), .ZN(new_n336));
  INV_X1    g0136(.A(new_n336), .ZN(new_n337));
  AOI21_X1  g0137(.A(new_n322), .B1(new_n334), .B2(new_n337), .ZN(new_n338));
  OAI21_X1  g0138(.A(new_n293), .B1(new_n321), .B2(new_n338), .ZN(new_n339));
  AOI21_X1  g0139(.A(new_n336), .B1(new_n333), .B2(new_n286), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n340), .A2(G190), .ZN(new_n341));
  INV_X1    g0141(.A(G107), .ZN(new_n342));
  AOI21_X1  g0142(.A(new_n342), .B1(new_n325), .B2(new_n327), .ZN(new_n343));
  AOI21_X1  g0143(.A(new_n343), .B1(new_n281), .B2(new_n331), .ZN(new_n344));
  AOI21_X1  g0144(.A(new_n273), .B1(new_n344), .B2(new_n323), .ZN(new_n345));
  OAI21_X1  g0145(.A(G200), .B1(new_n345), .B2(new_n336), .ZN(new_n346));
  OAI21_X1  g0146(.A(new_n318), .B1(new_n246), .B2(new_n250), .ZN(new_n347));
  XNOR2_X1  g0147(.A(KEYINPUT15), .B(G87), .ZN(new_n348));
  NOR2_X1   g0148(.A1(new_n348), .A2(new_n247), .ZN(new_n349));
  OAI21_X1  g0149(.A(new_n245), .B1(new_n347), .B2(new_n349), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n350), .A2(KEYINPUT70), .ZN(new_n351));
  NAND3_X1  g0151(.A1(new_n319), .A2(new_n314), .A3(new_n245), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n351), .A2(new_n352), .ZN(new_n353));
  NAND4_X1  g0153(.A1(new_n346), .A2(new_n353), .A3(KEYINPUT72), .A4(new_n301), .ZN(new_n354));
  NAND3_X1  g0154(.A1(new_n339), .A2(new_n341), .A3(new_n354), .ZN(new_n355));
  INV_X1    g0155(.A(G169), .ZN(new_n356));
  OAI21_X1  g0156(.A(new_n356), .B1(new_n345), .B2(new_n336), .ZN(new_n357));
  INV_X1    g0157(.A(G179), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n340), .A2(new_n358), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n357), .A2(new_n359), .ZN(new_n360));
  INV_X1    g0160(.A(new_n321), .ZN(new_n361));
  NOR2_X1   g0161(.A1(new_n360), .A2(new_n361), .ZN(new_n362));
  INV_X1    g0162(.A(new_n362), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n288), .A2(new_n356), .ZN(new_n364));
  OAI211_X1 g0164(.A(new_n364), .B(new_n268), .C1(G179), .C2(new_n288), .ZN(new_n365));
  NAND4_X1  g0165(.A1(new_n292), .A2(new_n355), .A3(new_n363), .A4(new_n365), .ZN(new_n366));
  OR2_X1    g0166(.A1(G223), .A2(G1698), .ZN(new_n367));
  INV_X1    g0167(.A(G226), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n368), .A2(G1698), .ZN(new_n369));
  NAND4_X1  g0169(.A1(new_n325), .A2(new_n367), .A3(new_n327), .A4(new_n369), .ZN(new_n370));
  NAND2_X1  g0170(.A1(G33), .A2(G87), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n370), .A2(new_n371), .ZN(new_n372));
  AOI21_X1  g0172(.A(G190), .B1(new_n372), .B2(new_n286), .ZN(new_n373));
  NAND3_X1  g0173(.A1(new_n273), .A2(G232), .A3(new_n277), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n275), .A2(new_n374), .ZN(new_n375));
  INV_X1    g0175(.A(KEYINPUT75), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n375), .A2(new_n376), .ZN(new_n377));
  NAND3_X1  g0177(.A1(new_n275), .A2(KEYINPUT75), .A3(new_n374), .ZN(new_n378));
  NAND3_X1  g0178(.A1(new_n373), .A2(new_n377), .A3(new_n378), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n379), .A2(KEYINPUT76), .ZN(new_n380));
  AOI21_X1  g0180(.A(new_n273), .B1(new_n370), .B2(new_n371), .ZN(new_n381));
  OAI21_X1  g0181(.A(new_n322), .B1(new_n381), .B2(new_n375), .ZN(new_n382));
  INV_X1    g0182(.A(KEYINPUT76), .ZN(new_n383));
  NAND4_X1  g0183(.A1(new_n373), .A2(new_n377), .A3(new_n383), .A4(new_n378), .ZN(new_n384));
  NAND3_X1  g0184(.A1(new_n380), .A2(new_n382), .A3(new_n384), .ZN(new_n385));
  NOR2_X1   g0185(.A1(new_n246), .A2(new_n264), .ZN(new_n386));
  AOI22_X1  g0186(.A1(new_n261), .A2(new_n386), .B1(new_n258), .B2(new_n246), .ZN(new_n387));
  INV_X1    g0187(.A(new_n387), .ZN(new_n388));
  XNOR2_X1  g0188(.A(G58), .B(G68), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n389), .A2(G20), .ZN(new_n390));
  NAND2_X1  g0190(.A1(new_n249), .A2(G159), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n390), .A2(new_n391), .ZN(new_n392));
  AOI21_X1  g0192(.A(G20), .B1(new_n325), .B2(new_n327), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n221), .A2(KEYINPUT7), .ZN(new_n394));
  OAI22_X1  g0194(.A1(new_n393), .A2(KEYINPUT7), .B1(new_n281), .B2(new_n394), .ZN(new_n395));
  AOI21_X1  g0195(.A(new_n392), .B1(new_n395), .B2(G68), .ZN(new_n396));
  AOI21_X1  g0196(.A(new_n298), .B1(new_n396), .B2(KEYINPUT16), .ZN(new_n397));
  XNOR2_X1  g0197(.A(KEYINPUT73), .B(KEYINPUT16), .ZN(new_n398));
  INV_X1    g0198(.A(new_n398), .ZN(new_n399));
  INV_X1    g0199(.A(G68), .ZN(new_n400));
  NOR2_X1   g0200(.A1(new_n326), .A2(G33), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n401), .A2(KEYINPUT74), .ZN(new_n402));
  INV_X1    g0202(.A(KEYINPUT7), .ZN(new_n403));
  NOR2_X1   g0203(.A1(new_n403), .A2(G20), .ZN(new_n404));
  OAI211_X1 g0204(.A(new_n402), .B(new_n404), .C1(new_n328), .C2(KEYINPUT74), .ZN(new_n405));
  OAI21_X1  g0205(.A(new_n403), .B1(new_n281), .B2(G20), .ZN(new_n406));
  AOI21_X1  g0206(.A(new_n400), .B1(new_n405), .B2(new_n406), .ZN(new_n407));
  OAI21_X1  g0207(.A(new_n399), .B1(new_n407), .B2(new_n392), .ZN(new_n408));
  AOI21_X1  g0208(.A(new_n388), .B1(new_n397), .B2(new_n408), .ZN(new_n409));
  AND3_X1   g0209(.A1(new_n385), .A2(new_n409), .A3(KEYINPUT17), .ZN(new_n410));
  AOI21_X1  g0210(.A(KEYINPUT17), .B1(new_n385), .B2(new_n409), .ZN(new_n411));
  NOR2_X1   g0211(.A1(new_n410), .A2(new_n411), .ZN(new_n412));
  INV_X1    g0212(.A(new_n381), .ZN(new_n413));
  NAND4_X1  g0213(.A1(new_n377), .A2(new_n413), .A3(new_n378), .A4(new_n358), .ZN(new_n414));
  OAI21_X1  g0214(.A(new_n356), .B1(new_n381), .B2(new_n375), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n414), .A2(new_n415), .ZN(new_n416));
  NOR3_X1   g0216(.A1(new_n409), .A2(KEYINPUT18), .A3(new_n416), .ZN(new_n417));
  INV_X1    g0217(.A(KEYINPUT18), .ZN(new_n418));
  AOI22_X1  g0218(.A1(new_n389), .A2(G20), .B1(G159), .B2(new_n249), .ZN(new_n419));
  AOI21_X1  g0219(.A(new_n394), .B1(new_n325), .B2(new_n327), .ZN(new_n420));
  NOR2_X1   g0220(.A1(new_n324), .A2(KEYINPUT3), .ZN(new_n421));
  OAI21_X1  g0221(.A(new_n221), .B1(new_n401), .B2(new_n421), .ZN(new_n422));
  AOI21_X1  g0222(.A(new_n420), .B1(new_n422), .B2(new_n403), .ZN(new_n423));
  OAI211_X1 g0223(.A(KEYINPUT16), .B(new_n419), .C1(new_n423), .C2(new_n400), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n424), .A2(new_n245), .ZN(new_n425));
  INV_X1    g0225(.A(KEYINPUT74), .ZN(new_n426));
  AND3_X1   g0226(.A1(new_n325), .A2(new_n327), .A3(new_n426), .ZN(new_n427));
  OAI21_X1  g0227(.A(new_n404), .B1(new_n325), .B2(new_n426), .ZN(new_n428));
  OAI22_X1  g0228(.A1(new_n427), .A2(new_n428), .B1(new_n393), .B2(KEYINPUT7), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n429), .A2(G68), .ZN(new_n430));
  AOI21_X1  g0230(.A(new_n398), .B1(new_n430), .B2(new_n419), .ZN(new_n431));
  OAI21_X1  g0231(.A(new_n387), .B1(new_n425), .B2(new_n431), .ZN(new_n432));
  INV_X1    g0232(.A(new_n416), .ZN(new_n433));
  AOI21_X1  g0233(.A(new_n418), .B1(new_n432), .B2(new_n433), .ZN(new_n434));
  NOR2_X1   g0234(.A1(new_n417), .A2(new_n434), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n412), .A2(new_n435), .ZN(new_n436));
  OAI21_X1  g0236(.A(KEYINPUT12), .B1(new_n257), .B2(G68), .ZN(new_n437));
  OR3_X1    g0237(.A1(new_n257), .A2(KEYINPUT12), .A3(G68), .ZN(new_n438));
  NOR2_X1   g0238(.A1(new_n264), .A2(new_n400), .ZN(new_n439));
  AOI22_X1  g0239(.A1(new_n437), .A2(new_n438), .B1(new_n261), .B2(new_n439), .ZN(new_n440));
  AOI22_X1  g0240(.A1(new_n249), .A2(G50), .B1(G20), .B2(new_n400), .ZN(new_n441));
  OAI21_X1  g0241(.A(new_n441), .B1(new_n294), .B2(new_n247), .ZN(new_n442));
  NAND3_X1  g0242(.A1(new_n442), .A2(KEYINPUT11), .A3(new_n245), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n440), .A2(new_n443), .ZN(new_n444));
  AOI21_X1  g0244(.A(KEYINPUT11), .B1(new_n442), .B2(new_n245), .ZN(new_n445));
  NOR2_X1   g0245(.A1(new_n444), .A2(new_n445), .ZN(new_n446));
  INV_X1    g0246(.A(G190), .ZN(new_n447));
  NAND2_X1  g0247(.A1(new_n368), .A2(new_n283), .ZN(new_n448));
  NAND2_X1  g0248(.A1(new_n228), .A2(G1698), .ZN(new_n449));
  NAND4_X1  g0249(.A1(new_n325), .A2(new_n448), .A3(new_n327), .A4(new_n449), .ZN(new_n450));
  NAND2_X1  g0250(.A1(G33), .A2(G97), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n450), .A2(new_n451), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n452), .A2(new_n286), .ZN(new_n453));
  NAND3_X1  g0253(.A1(new_n273), .A2(G238), .A3(new_n277), .ZN(new_n454));
  AND2_X1   g0254(.A1(new_n275), .A2(new_n454), .ZN(new_n455));
  INV_X1    g0255(.A(KEYINPUT13), .ZN(new_n456));
  NAND3_X1  g0256(.A1(new_n453), .A2(new_n455), .A3(new_n456), .ZN(new_n457));
  AOI21_X1  g0257(.A(new_n273), .B1(new_n450), .B2(new_n451), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n275), .A2(new_n454), .ZN(new_n459));
  OAI21_X1  g0259(.A(KEYINPUT13), .B1(new_n458), .B2(new_n459), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n457), .A2(new_n460), .ZN(new_n461));
  OAI21_X1  g0261(.A(new_n446), .B1(new_n447), .B2(new_n461), .ZN(new_n462));
  AOI21_X1  g0262(.A(new_n322), .B1(new_n457), .B2(new_n460), .ZN(new_n463));
  NOR2_X1   g0263(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  INV_X1    g0264(.A(new_n464), .ZN(new_n465));
  INV_X1    g0265(.A(new_n446), .ZN(new_n466));
  INV_X1    g0266(.A(KEYINPUT14), .ZN(new_n467));
  NAND3_X1  g0267(.A1(new_n461), .A2(new_n467), .A3(G169), .ZN(new_n468));
  NAND3_X1  g0268(.A1(new_n457), .A2(G179), .A3(new_n460), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  AOI21_X1  g0270(.A(new_n467), .B1(new_n461), .B2(G169), .ZN(new_n471));
  OAI21_X1  g0271(.A(new_n466), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  NAND2_X1  g0272(.A1(new_n465), .A2(new_n472), .ZN(new_n473));
  NOR3_X1   g0273(.A1(new_n366), .A2(new_n436), .A3(new_n473), .ZN(new_n474));
  OAI21_X1  g0274(.A(KEYINPUT78), .B1(new_n324), .B2(G1), .ZN(new_n475));
  INV_X1    g0275(.A(KEYINPUT78), .ZN(new_n476));
  NAND3_X1  g0276(.A1(new_n476), .A2(new_n256), .A3(G33), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n475), .A2(new_n477), .ZN(new_n478));
  NOR3_X1   g0278(.A1(new_n478), .A2(new_n260), .A3(new_n342), .ZN(new_n479));
  NAND4_X1  g0279(.A1(new_n256), .A2(new_n342), .A3(G13), .A4(G20), .ZN(new_n480));
  XNOR2_X1  g0280(.A(new_n480), .B(KEYINPUT25), .ZN(new_n481));
  OAI21_X1  g0281(.A(KEYINPUT81), .B1(new_n479), .B2(new_n481), .ZN(new_n482));
  AND2_X1   g0282(.A1(new_n475), .A2(new_n477), .ZN(new_n483));
  NAND3_X1  g0283(.A1(new_n261), .A2(new_n483), .A3(G107), .ZN(new_n484));
  INV_X1    g0284(.A(KEYINPUT81), .ZN(new_n485));
  INV_X1    g0285(.A(KEYINPUT25), .ZN(new_n486));
  XNOR2_X1  g0286(.A(new_n480), .B(new_n486), .ZN(new_n487));
  NAND3_X1  g0287(.A1(new_n484), .A2(new_n485), .A3(new_n487), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n482), .A2(new_n488), .ZN(new_n489));
  NAND3_X1  g0289(.A1(new_n221), .A2(KEYINPUT80), .A3(G87), .ZN(new_n490));
  OAI21_X1  g0290(.A(KEYINPUT22), .B1(new_n328), .B2(new_n490), .ZN(new_n491));
  INV_X1    g0291(.A(new_n490), .ZN(new_n492));
  INV_X1    g0292(.A(KEYINPUT22), .ZN(new_n493));
  NAND3_X1  g0293(.A1(new_n281), .A2(new_n492), .A3(new_n493), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n491), .A2(new_n494), .ZN(new_n495));
  INV_X1    g0295(.A(KEYINPUT23), .ZN(new_n496));
  OAI21_X1  g0296(.A(new_n496), .B1(new_n221), .B2(G107), .ZN(new_n497));
  NAND3_X1  g0297(.A1(new_n342), .A2(KEYINPUT23), .A3(G20), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  NAND3_X1  g0299(.A1(new_n221), .A2(G33), .A3(G116), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  INV_X1    g0301(.A(new_n501), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n495), .A2(new_n502), .ZN(new_n503));
  INV_X1    g0303(.A(KEYINPUT24), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  AOI21_X1  g0305(.A(new_n501), .B1(new_n491), .B2(new_n494), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n506), .A2(KEYINPUT24), .ZN(new_n507));
  NAND3_X1  g0307(.A1(new_n505), .A2(new_n507), .A3(new_n245), .ZN(new_n508));
  INV_X1    g0308(.A(G45), .ZN(new_n509));
  NOR2_X1   g0309(.A1(new_n509), .A2(G1), .ZN(new_n510));
  AND2_X1   g0310(.A1(KEYINPUT5), .A2(G41), .ZN(new_n511));
  NOR2_X1   g0311(.A1(KEYINPUT5), .A2(G41), .ZN(new_n512));
  OAI21_X1  g0312(.A(new_n510), .B1(new_n511), .B2(new_n512), .ZN(new_n513));
  NAND3_X1  g0313(.A1(new_n513), .A2(G264), .A3(new_n273), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n514), .A2(KEYINPUT83), .ZN(new_n515));
  INV_X1    g0315(.A(KEYINPUT83), .ZN(new_n516));
  NAND4_X1  g0316(.A1(new_n513), .A2(new_n516), .A3(G264), .A4(new_n273), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n515), .A2(new_n517), .ZN(new_n518));
  INV_X1    g0318(.A(G274), .ZN(new_n519));
  AND2_X1   g0319(.A1(G1), .A2(G13), .ZN(new_n520));
  AOI21_X1  g0320(.A(new_n519), .B1(new_n520), .B2(new_n272), .ZN(new_n521));
  XNOR2_X1  g0321(.A(KEYINPUT5), .B(G41), .ZN(new_n522));
  NAND3_X1  g0322(.A1(new_n521), .A2(new_n510), .A3(new_n522), .ZN(new_n523));
  INV_X1    g0323(.A(G250), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n524), .A2(new_n283), .ZN(new_n525));
  INV_X1    g0325(.A(G257), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n526), .A2(G1698), .ZN(new_n527));
  NAND4_X1  g0327(.A1(new_n325), .A2(new_n525), .A3(new_n327), .A4(new_n527), .ZN(new_n528));
  AND2_X1   g0328(.A1(KEYINPUT82), .A2(G294), .ZN(new_n529));
  NOR2_X1   g0329(.A1(KEYINPUT82), .A2(G294), .ZN(new_n530));
  OAI21_X1  g0330(.A(G33), .B1(new_n529), .B2(new_n530), .ZN(new_n531));
  AOI21_X1  g0331(.A(new_n273), .B1(new_n528), .B2(new_n531), .ZN(new_n532));
  INV_X1    g0332(.A(new_n532), .ZN(new_n533));
  AND3_X1   g0333(.A1(new_n518), .A2(new_n523), .A3(new_n533), .ZN(new_n534));
  AOI22_X1  g0334(.A1(new_n489), .A2(new_n508), .B1(new_n534), .B2(new_n358), .ZN(new_n535));
  AOI21_X1  g0335(.A(new_n532), .B1(new_n515), .B2(new_n517), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n536), .A2(new_n523), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n537), .A2(new_n356), .ZN(new_n538));
  NAND3_X1  g0338(.A1(new_n536), .A2(new_n447), .A3(new_n523), .ZN(new_n539));
  OAI21_X1  g0339(.A(new_n539), .B1(new_n534), .B2(G200), .ZN(new_n540));
  AOI21_X1  g0340(.A(new_n298), .B1(new_n503), .B2(new_n504), .ZN(new_n541));
  AOI22_X1  g0341(.A1(new_n541), .A2(new_n507), .B1(new_n488), .B2(new_n482), .ZN(new_n542));
  AOI22_X1  g0342(.A1(new_n535), .A2(new_n538), .B1(new_n540), .B2(new_n542), .ZN(new_n543));
  NAND3_X1  g0343(.A1(KEYINPUT19), .A2(G33), .A3(G97), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n544), .A2(new_n221), .ZN(new_n545));
  NOR2_X1   g0345(.A1(G97), .A2(G107), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n546), .A2(new_n309), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n545), .A2(new_n547), .ZN(new_n548));
  NOR2_X1   g0348(.A1(new_n400), .A2(G20), .ZN(new_n549));
  NAND3_X1  g0349(.A1(new_n549), .A2(new_n325), .A3(new_n327), .ZN(new_n550));
  INV_X1    g0350(.A(KEYINPUT19), .ZN(new_n551));
  INV_X1    g0351(.A(G97), .ZN(new_n552));
  OAI21_X1  g0352(.A(new_n551), .B1(new_n247), .B2(new_n552), .ZN(new_n553));
  NAND3_X1  g0353(.A1(new_n548), .A2(new_n550), .A3(new_n553), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n554), .A2(new_n245), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n348), .A2(new_n258), .ZN(new_n556));
  INV_X1    g0356(.A(new_n348), .ZN(new_n557));
  NAND3_X1  g0357(.A1(new_n261), .A2(new_n483), .A3(new_n557), .ZN(new_n558));
  NAND3_X1  g0358(.A1(new_n555), .A2(new_n556), .A3(new_n558), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n330), .A2(new_n283), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n335), .A2(G1698), .ZN(new_n561));
  NAND4_X1  g0361(.A1(new_n325), .A2(new_n560), .A3(new_n327), .A4(new_n561), .ZN(new_n562));
  NAND2_X1  g0362(.A1(G33), .A2(G116), .ZN(new_n563));
  AOI21_X1  g0363(.A(new_n273), .B1(new_n562), .B2(new_n563), .ZN(new_n564));
  AOI21_X1  g0364(.A(new_n524), .B1(new_n256), .B2(G45), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n565), .A2(new_n273), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n273), .A2(G274), .ZN(new_n567));
  INV_X1    g0367(.A(new_n510), .ZN(new_n568));
  OAI21_X1  g0368(.A(new_n566), .B1(new_n567), .B2(new_n568), .ZN(new_n569));
  OAI21_X1  g0369(.A(new_n356), .B1(new_n564), .B2(new_n569), .ZN(new_n570));
  AOI22_X1  g0370(.A1(new_n521), .A2(new_n510), .B1(new_n273), .B2(new_n565), .ZN(new_n571));
  NOR2_X1   g0371(.A1(G238), .A2(G1698), .ZN(new_n572));
  AOI21_X1  g0372(.A(new_n572), .B1(new_n335), .B2(G1698), .ZN(new_n573));
  AOI22_X1  g0373(.A1(new_n573), .A2(new_n281), .B1(G33), .B2(G116), .ZN(new_n574));
  OAI211_X1 g0374(.A(new_n358), .B(new_n571), .C1(new_n574), .C2(new_n273), .ZN(new_n575));
  NAND3_X1  g0375(.A1(new_n559), .A2(new_n570), .A3(new_n575), .ZN(new_n576));
  OAI21_X1  g0376(.A(G200), .B1(new_n564), .B2(new_n569), .ZN(new_n577));
  OAI211_X1 g0377(.A(G190), .B(new_n571), .C1(new_n574), .C2(new_n273), .ZN(new_n578));
  AOI22_X1  g0378(.A1(new_n554), .A2(new_n245), .B1(new_n258), .B2(new_n348), .ZN(new_n579));
  NAND3_X1  g0379(.A1(new_n261), .A2(new_n483), .A3(G87), .ZN(new_n580));
  NAND4_X1  g0380(.A1(new_n577), .A2(new_n578), .A3(new_n579), .A4(new_n580), .ZN(new_n581));
  AND2_X1   g0381(.A1(new_n576), .A2(new_n581), .ZN(new_n582));
  NAND4_X1  g0382(.A1(new_n325), .A2(new_n327), .A3(G244), .A4(new_n283), .ZN(new_n583));
  INV_X1    g0383(.A(KEYINPUT4), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  NAND2_X1  g0385(.A1(G33), .A2(G283), .ZN(new_n586));
  INV_X1    g0386(.A(new_n586), .ZN(new_n587));
  NAND2_X1  g0387(.A1(G250), .A2(G1698), .ZN(new_n588));
  NAND2_X1  g0388(.A1(KEYINPUT4), .A2(G244), .ZN(new_n589));
  OAI21_X1  g0389(.A(new_n588), .B1(new_n589), .B2(G1698), .ZN(new_n590));
  AOI21_X1  g0390(.A(new_n587), .B1(new_n281), .B2(new_n590), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n585), .A2(new_n591), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n592), .A2(new_n286), .ZN(new_n593));
  NAND3_X1  g0393(.A1(new_n513), .A2(G257), .A3(new_n273), .ZN(new_n594));
  AND2_X1   g0394(.A1(new_n594), .A2(new_n523), .ZN(new_n595));
  AOI21_X1  g0395(.A(new_n356), .B1(new_n593), .B2(new_n595), .ZN(new_n596));
  AOI21_X1  g0396(.A(new_n273), .B1(new_n585), .B2(new_n591), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n594), .A2(new_n523), .ZN(new_n598));
  NOR3_X1   g0398(.A1(new_n597), .A2(new_n598), .A3(new_n358), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n429), .A2(G107), .ZN(new_n600));
  INV_X1    g0400(.A(KEYINPUT6), .ZN(new_n601));
  AND2_X1   g0401(.A1(G97), .A2(G107), .ZN(new_n602));
  OAI21_X1  g0402(.A(new_n601), .B1(new_n602), .B2(new_n546), .ZN(new_n603));
  NAND2_X1  g0403(.A1(KEYINPUT6), .A2(G97), .ZN(new_n604));
  OAI21_X1  g0404(.A(KEYINPUT77), .B1(new_n604), .B2(G107), .ZN(new_n605));
  INV_X1    g0405(.A(KEYINPUT77), .ZN(new_n606));
  NAND4_X1  g0406(.A1(new_n606), .A2(new_n342), .A3(KEYINPUT6), .A4(G97), .ZN(new_n607));
  NAND3_X1  g0407(.A1(new_n603), .A2(new_n605), .A3(new_n607), .ZN(new_n608));
  AOI22_X1  g0408(.A1(new_n608), .A2(G20), .B1(G77), .B2(new_n249), .ZN(new_n609));
  AOI21_X1  g0409(.A(new_n298), .B1(new_n600), .B2(new_n609), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n258), .A2(new_n552), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n261), .A2(new_n483), .ZN(new_n612));
  OAI21_X1  g0412(.A(new_n611), .B1(new_n612), .B2(new_n552), .ZN(new_n613));
  OAI22_X1  g0413(.A1(new_n596), .A2(new_n599), .B1(new_n610), .B2(new_n613), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n608), .A2(G20), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n249), .A2(G77), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n615), .A2(new_n616), .ZN(new_n617));
  AOI21_X1  g0417(.A(new_n342), .B1(new_n405), .B2(new_n406), .ZN(new_n618));
  OAI21_X1  g0418(.A(new_n245), .B1(new_n617), .B2(new_n618), .ZN(new_n619));
  INV_X1    g0419(.A(new_n613), .ZN(new_n620));
  AOI21_X1  g0420(.A(G200), .B1(new_n593), .B2(new_n595), .ZN(new_n621));
  NOR3_X1   g0421(.A1(new_n597), .A2(new_n598), .A3(G190), .ZN(new_n622));
  OAI211_X1 g0422(.A(new_n619), .B(new_n620), .C1(new_n621), .C2(new_n622), .ZN(new_n623));
  AND3_X1   g0423(.A1(new_n582), .A2(new_n614), .A3(new_n623), .ZN(new_n624));
  NOR2_X1   g0424(.A1(new_n283), .A2(G264), .ZN(new_n625));
  NOR2_X1   g0425(.A1(G257), .A2(G1698), .ZN(new_n626));
  OAI211_X1 g0426(.A(new_n325), .B(new_n327), .C1(new_n625), .C2(new_n626), .ZN(new_n627));
  INV_X1    g0427(.A(G303), .ZN(new_n628));
  OAI21_X1  g0428(.A(new_n628), .B1(new_n401), .B2(new_n421), .ZN(new_n629));
  NAND3_X1  g0429(.A1(new_n627), .A2(new_n629), .A3(new_n286), .ZN(new_n630));
  NAND3_X1  g0430(.A1(new_n513), .A2(G270), .A3(new_n273), .ZN(new_n631));
  NAND3_X1  g0431(.A1(new_n630), .A2(new_n523), .A3(new_n631), .ZN(new_n632));
  NAND3_X1  g0432(.A1(new_n632), .A2(KEYINPUT21), .A3(G169), .ZN(new_n633));
  NAND4_X1  g0433(.A1(new_n630), .A2(G179), .A3(new_n523), .A4(new_n631), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n633), .A2(new_n634), .ZN(new_n635));
  INV_X1    g0435(.A(G116), .ZN(new_n636));
  NAND4_X1  g0436(.A1(new_n256), .A2(new_n636), .A3(G13), .A4(G20), .ZN(new_n637));
  INV_X1    g0437(.A(KEYINPUT79), .ZN(new_n638));
  XNOR2_X1  g0438(.A(new_n637), .B(new_n638), .ZN(new_n639));
  OAI21_X1  g0439(.A(new_n639), .B1(new_n612), .B2(new_n636), .ZN(new_n640));
  AOI22_X1  g0440(.A1(new_n244), .A2(new_n220), .B1(G20), .B2(new_n636), .ZN(new_n641));
  OAI211_X1 g0441(.A(new_n586), .B(new_n221), .C1(G33), .C2(new_n552), .ZN(new_n642));
  AND3_X1   g0442(.A1(new_n641), .A2(KEYINPUT20), .A3(new_n642), .ZN(new_n643));
  AOI21_X1  g0443(.A(KEYINPUT20), .B1(new_n641), .B2(new_n642), .ZN(new_n644));
  NOR2_X1   g0444(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  NOR2_X1   g0445(.A1(new_n640), .A2(new_n645), .ZN(new_n646));
  INV_X1    g0446(.A(new_n646), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n635), .A2(new_n647), .ZN(new_n648));
  OAI211_X1 g0448(.A(G169), .B(new_n632), .C1(new_n640), .C2(new_n645), .ZN(new_n649));
  INV_X1    g0449(.A(KEYINPUT21), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n632), .A2(G200), .ZN(new_n652));
  OAI211_X1 g0452(.A(new_n646), .B(new_n652), .C1(new_n447), .C2(new_n632), .ZN(new_n653));
  AND3_X1   g0453(.A1(new_n648), .A2(new_n651), .A3(new_n653), .ZN(new_n654));
  AND4_X1   g0454(.A1(new_n474), .A2(new_n543), .A3(new_n624), .A4(new_n654), .ZN(G372));
  INV_X1    g0455(.A(new_n360), .ZN(new_n656));
  OAI211_X1 g0456(.A(new_n656), .B(new_n321), .C1(new_n462), .C2(new_n463), .ZN(new_n657));
  AND3_X1   g0457(.A1(new_n472), .A2(new_n657), .A3(KEYINPUT86), .ZN(new_n658));
  AOI21_X1  g0458(.A(KEYINPUT86), .B1(new_n472), .B2(new_n657), .ZN(new_n659));
  AOI21_X1  g0459(.A(new_n392), .B1(new_n429), .B2(G68), .ZN(new_n660));
  OAI211_X1 g0460(.A(new_n424), .B(new_n245), .C1(new_n660), .C2(new_n398), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n384), .A2(new_n382), .ZN(new_n662));
  AND3_X1   g0462(.A1(new_n275), .A2(new_n374), .A3(KEYINPUT75), .ZN(new_n663));
  AOI21_X1  g0463(.A(KEYINPUT75), .B1(new_n275), .B2(new_n374), .ZN(new_n664));
  NOR2_X1   g0464(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  AOI21_X1  g0465(.A(new_n383), .B1(new_n665), .B2(new_n373), .ZN(new_n666));
  OAI211_X1 g0466(.A(new_n661), .B(new_n387), .C1(new_n662), .C2(new_n666), .ZN(new_n667));
  INV_X1    g0467(.A(KEYINPUT17), .ZN(new_n668));
  XNOR2_X1  g0468(.A(new_n667), .B(new_n668), .ZN(new_n669));
  NOR3_X1   g0469(.A1(new_n658), .A2(new_n659), .A3(new_n669), .ZN(new_n670));
  INV_X1    g0470(.A(new_n435), .ZN(new_n671));
  OAI21_X1  g0471(.A(KEYINPUT87), .B1(new_n670), .B2(new_n671), .ZN(new_n672));
  INV_X1    g0472(.A(KEYINPUT87), .ZN(new_n673));
  AND2_X1   g0473(.A1(new_n472), .A2(new_n657), .ZN(new_n674));
  OAI21_X1  g0474(.A(new_n412), .B1(new_n674), .B2(KEYINPUT86), .ZN(new_n675));
  OAI211_X1 g0475(.A(new_n673), .B(new_n435), .C1(new_n675), .C2(new_n658), .ZN(new_n676));
  NAND3_X1  g0476(.A1(new_n672), .A2(new_n676), .A3(new_n292), .ZN(new_n677));
  AND2_X1   g0477(.A1(new_n677), .A2(new_n365), .ZN(new_n678));
  INV_X1    g0478(.A(new_n576), .ZN(new_n679));
  NAND3_X1  g0479(.A1(new_n582), .A2(new_n614), .A3(new_n623), .ZN(new_n680));
  OAI21_X1  g0480(.A(new_n245), .B1(new_n506), .B2(KEYINPUT24), .ZN(new_n681));
  AND3_X1   g0481(.A1(new_n495), .A2(KEYINPUT24), .A3(new_n502), .ZN(new_n682));
  OAI21_X1  g0482(.A(new_n489), .B1(new_n681), .B2(new_n682), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n537), .A2(new_n322), .ZN(new_n684));
  AOI21_X1  g0484(.A(new_n683), .B1(new_n539), .B2(new_n684), .ZN(new_n685));
  NOR2_X1   g0485(.A1(new_n680), .A2(new_n685), .ZN(new_n686));
  NAND3_X1  g0486(.A1(new_n536), .A2(new_n358), .A3(new_n523), .ZN(new_n687));
  NAND3_X1  g0487(.A1(new_n683), .A2(new_n538), .A3(new_n687), .ZN(new_n688));
  AOI22_X1  g0488(.A1(new_n635), .A2(new_n647), .B1(new_n649), .B2(new_n650), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  AOI21_X1  g0490(.A(new_n679), .B1(new_n686), .B2(new_n690), .ZN(new_n691));
  INV_X1    g0491(.A(KEYINPUT26), .ZN(new_n692));
  OAI21_X1  g0492(.A(KEYINPUT84), .B1(new_n596), .B2(new_n599), .ZN(new_n693));
  NAND3_X1  g0493(.A1(new_n593), .A2(G179), .A3(new_n595), .ZN(new_n694));
  INV_X1    g0494(.A(KEYINPUT84), .ZN(new_n695));
  OAI21_X1  g0495(.A(G169), .B1(new_n597), .B2(new_n598), .ZN(new_n696));
  NAND3_X1  g0496(.A1(new_n694), .A2(new_n695), .A3(new_n696), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n619), .A2(new_n620), .ZN(new_n698));
  NAND3_X1  g0498(.A1(new_n693), .A2(new_n697), .A3(new_n698), .ZN(new_n699));
  INV_X1    g0499(.A(new_n582), .ZN(new_n700));
  OAI21_X1  g0500(.A(new_n692), .B1(new_n699), .B2(new_n700), .ZN(new_n701));
  INV_X1    g0501(.A(new_n614), .ZN(new_n702));
  NAND4_X1  g0502(.A1(new_n702), .A2(KEYINPUT85), .A3(KEYINPUT26), .A4(new_n582), .ZN(new_n703));
  INV_X1    g0503(.A(KEYINPUT85), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n694), .A2(new_n696), .ZN(new_n705));
  NAND4_X1  g0505(.A1(new_n698), .A2(new_n705), .A3(new_n576), .A4(new_n581), .ZN(new_n706));
  OAI21_X1  g0506(.A(new_n704), .B1(new_n706), .B2(new_n692), .ZN(new_n707));
  NAND3_X1  g0507(.A1(new_n701), .A2(new_n703), .A3(new_n707), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n691), .A2(new_n708), .ZN(new_n709));
  NAND2_X1  g0509(.A1(new_n474), .A2(new_n709), .ZN(new_n710));
  NAND2_X1  g0510(.A1(new_n678), .A2(new_n710), .ZN(G369));
  INV_X1    g0511(.A(new_n689), .ZN(new_n712));
  NAND3_X1  g0512(.A1(new_n256), .A2(new_n221), .A3(G13), .ZN(new_n713));
  OR2_X1    g0513(.A1(new_n713), .A2(KEYINPUT27), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n713), .A2(KEYINPUT27), .ZN(new_n715));
  NAND3_X1  g0515(.A1(new_n714), .A2(new_n715), .A3(G213), .ZN(new_n716));
  INV_X1    g0516(.A(G343), .ZN(new_n717));
  NOR2_X1   g0517(.A1(new_n716), .A2(new_n717), .ZN(new_n718));
  NAND2_X1  g0518(.A1(new_n647), .A2(new_n718), .ZN(new_n719));
  MUX2_X1   g0519(.A(new_n712), .B(new_n654), .S(new_n719), .Z(new_n720));
  NAND2_X1  g0520(.A1(new_n720), .A2(G330), .ZN(new_n721));
  INV_X1    g0521(.A(new_n721), .ZN(new_n722));
  INV_X1    g0522(.A(new_n543), .ZN(new_n723));
  INV_X1    g0523(.A(new_n718), .ZN(new_n724));
  NOR2_X1   g0524(.A1(new_n542), .A2(new_n724), .ZN(new_n725));
  OAI22_X1  g0525(.A1(new_n723), .A2(new_n725), .B1(new_n688), .B2(new_n724), .ZN(new_n726));
  NAND2_X1  g0526(.A1(new_n722), .A2(new_n726), .ZN(new_n727));
  NAND3_X1  g0527(.A1(new_n535), .A2(new_n538), .A3(new_n724), .ZN(new_n728));
  NAND3_X1  g0528(.A1(new_n543), .A2(new_n712), .A3(new_n724), .ZN(new_n729));
  NAND3_X1  g0529(.A1(new_n727), .A2(new_n728), .A3(new_n729), .ZN(G399));
  NOR2_X1   g0530(.A1(new_n547), .A2(G116), .ZN(new_n731));
  NAND2_X1  g0531(.A1(new_n731), .A2(G1), .ZN(new_n732));
  INV_X1    g0532(.A(new_n217), .ZN(new_n733));
  NOR2_X1   g0533(.A1(new_n733), .A2(G41), .ZN(new_n734));
  MUX2_X1   g0534(.A(new_n732), .B(new_n223), .S(new_n734), .Z(new_n735));
  XOR2_X1   g0535(.A(new_n735), .B(KEYINPUT28), .Z(new_n736));
  INV_X1    g0536(.A(KEYINPUT29), .ZN(new_n737));
  NAND2_X1  g0537(.A1(new_n540), .A2(new_n542), .ZN(new_n738));
  NAND3_X1  g0538(.A1(new_n624), .A2(new_n690), .A3(new_n738), .ZN(new_n739));
  OAI21_X1  g0539(.A(KEYINPUT26), .B1(new_n699), .B2(new_n700), .ZN(new_n740));
  NAND3_X1  g0540(.A1(new_n702), .A2(new_n692), .A3(new_n582), .ZN(new_n741));
  NAND4_X1  g0541(.A1(new_n739), .A2(new_n576), .A3(new_n740), .A4(new_n741), .ZN(new_n742));
  AOI21_X1  g0542(.A(new_n737), .B1(new_n742), .B2(new_n724), .ZN(new_n743));
  AOI211_X1 g0543(.A(KEYINPUT29), .B(new_n718), .C1(new_n691), .C2(new_n708), .ZN(new_n744));
  INV_X1    g0544(.A(KEYINPUT88), .ZN(new_n745));
  AND3_X1   g0545(.A1(new_n630), .A2(new_n523), .A3(new_n631), .ZN(new_n746));
  OAI21_X1  g0546(.A(new_n358), .B1(new_n564), .B2(new_n569), .ZN(new_n747));
  OAI21_X1  g0547(.A(new_n745), .B1(new_n746), .B2(new_n747), .ZN(new_n748));
  NOR2_X1   g0548(.A1(new_n597), .A2(new_n598), .ZN(new_n749));
  INV_X1    g0549(.A(new_n749), .ZN(new_n750));
  OAI21_X1  g0550(.A(new_n571), .B1(new_n574), .B2(new_n273), .ZN(new_n751));
  NAND4_X1  g0551(.A1(new_n632), .A2(new_n751), .A3(KEYINPUT88), .A4(new_n358), .ZN(new_n752));
  NAND4_X1  g0552(.A1(new_n748), .A2(new_n537), .A3(new_n750), .A4(new_n752), .ZN(new_n753));
  NOR2_X1   g0553(.A1(new_n564), .A2(new_n569), .ZN(new_n754));
  AND3_X1   g0554(.A1(new_n518), .A2(new_n754), .A3(new_n533), .ZN(new_n755));
  INV_X1    g0555(.A(new_n634), .ZN(new_n756));
  NAND4_X1  g0556(.A1(new_n755), .A2(KEYINPUT30), .A3(new_n749), .A4(new_n756), .ZN(new_n757));
  NAND4_X1  g0557(.A1(new_n756), .A2(new_n749), .A3(new_n536), .A4(new_n754), .ZN(new_n758));
  INV_X1    g0558(.A(KEYINPUT30), .ZN(new_n759));
  NAND2_X1  g0559(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  NAND3_X1  g0560(.A1(new_n753), .A2(new_n757), .A3(new_n760), .ZN(new_n761));
  NAND2_X1  g0561(.A1(new_n761), .A2(new_n718), .ZN(new_n762));
  INV_X1    g0562(.A(KEYINPUT31), .ZN(new_n763));
  NAND2_X1  g0563(.A1(new_n762), .A2(new_n763), .ZN(new_n764));
  NAND4_X1  g0564(.A1(new_n543), .A2(new_n624), .A3(new_n654), .A4(new_n724), .ZN(new_n765));
  NAND2_X1  g0565(.A1(new_n753), .A2(new_n760), .ZN(new_n766));
  INV_X1    g0566(.A(KEYINPUT89), .ZN(new_n767));
  NAND2_X1  g0567(.A1(new_n766), .A2(new_n767), .ZN(new_n768));
  NAND3_X1  g0568(.A1(new_n753), .A2(new_n760), .A3(KEYINPUT89), .ZN(new_n769));
  AND3_X1   g0569(.A1(new_n768), .A2(new_n769), .A3(new_n757), .ZN(new_n770));
  NOR2_X1   g0570(.A1(new_n724), .A2(new_n763), .ZN(new_n771));
  INV_X1    g0571(.A(new_n771), .ZN(new_n772));
  OAI211_X1 g0572(.A(new_n764), .B(new_n765), .C1(new_n770), .C2(new_n772), .ZN(new_n773));
  AOI211_X1 g0573(.A(new_n743), .B(new_n744), .C1(G330), .C2(new_n773), .ZN(new_n774));
  OAI21_X1  g0574(.A(new_n736), .B1(new_n774), .B2(G1), .ZN(G364));
  INV_X1    g0575(.A(G13), .ZN(new_n776));
  NOR2_X1   g0576(.A1(new_n776), .A2(G20), .ZN(new_n777));
  AOI21_X1  g0577(.A(new_n256), .B1(new_n777), .B2(G45), .ZN(new_n778));
  INV_X1    g0578(.A(new_n778), .ZN(new_n779));
  NOR2_X1   g0579(.A1(new_n734), .A2(new_n779), .ZN(new_n780));
  NOR2_X1   g0580(.A1(new_n722), .A2(new_n780), .ZN(new_n781));
  OAI21_X1  g0581(.A(new_n781), .B1(G330), .B2(new_n720), .ZN(new_n782));
  NAND3_X1  g0582(.A1(new_n217), .A2(G355), .A3(new_n281), .ZN(new_n783));
  OAI21_X1  g0583(.A(new_n783), .B1(G116), .B2(new_n217), .ZN(new_n784));
  NOR2_X1   g0584(.A1(new_n733), .A2(new_n281), .ZN(new_n785));
  INV_X1    g0585(.A(new_n785), .ZN(new_n786));
  AOI21_X1  g0586(.A(new_n786), .B1(new_n509), .B2(new_n224), .ZN(new_n787));
  NAND2_X1  g0587(.A1(new_n242), .A2(G45), .ZN(new_n788));
  AOI21_X1  g0588(.A(new_n784), .B1(new_n787), .B2(new_n788), .ZN(new_n789));
  OAI21_X1  g0589(.A(G20), .B1(KEYINPUT90), .B2(G169), .ZN(new_n790));
  INV_X1    g0590(.A(new_n790), .ZN(new_n791));
  NAND2_X1  g0591(.A1(KEYINPUT90), .A2(G169), .ZN(new_n792));
  AOI21_X1  g0592(.A(new_n220), .B1(new_n791), .B2(new_n792), .ZN(new_n793));
  INV_X1    g0593(.A(new_n793), .ZN(new_n794));
  NOR2_X1   g0594(.A1(G13), .A2(G33), .ZN(new_n795));
  INV_X1    g0595(.A(new_n795), .ZN(new_n796));
  NOR2_X1   g0596(.A1(new_n796), .A2(G20), .ZN(new_n797));
  INV_X1    g0597(.A(new_n797), .ZN(new_n798));
  NAND2_X1  g0598(.A1(new_n794), .A2(new_n798), .ZN(new_n799));
  XNOR2_X1  g0599(.A(new_n799), .B(KEYINPUT91), .ZN(new_n800));
  OAI21_X1  g0600(.A(new_n780), .B1(new_n789), .B2(new_n800), .ZN(new_n801));
  NOR2_X1   g0601(.A1(new_n221), .A2(new_n358), .ZN(new_n802));
  NAND2_X1  g0602(.A1(new_n802), .A2(G200), .ZN(new_n803));
  NOR2_X1   g0603(.A1(new_n803), .A2(new_n447), .ZN(new_n804));
  INV_X1    g0604(.A(new_n804), .ZN(new_n805));
  XOR2_X1   g0605(.A(new_n802), .B(KEYINPUT92), .Z(new_n806));
  NOR3_X1   g0606(.A1(new_n806), .A2(new_n447), .A3(G200), .ZN(new_n807));
  INV_X1    g0607(.A(new_n807), .ZN(new_n808));
  OAI221_X1 g0608(.A(new_n281), .B1(new_n253), .B2(new_n805), .C1(new_n808), .C2(new_n302), .ZN(new_n809));
  NOR3_X1   g0609(.A1(new_n806), .A2(G190), .A3(G200), .ZN(new_n810));
  AOI21_X1  g0610(.A(new_n809), .B1(G77), .B2(new_n810), .ZN(new_n811));
  NOR2_X1   g0611(.A1(new_n221), .A2(G179), .ZN(new_n812));
  NOR2_X1   g0612(.A1(G190), .A2(G200), .ZN(new_n813));
  NAND2_X1  g0613(.A1(new_n812), .A2(new_n813), .ZN(new_n814));
  INV_X1    g0614(.A(G159), .ZN(new_n815));
  NOR2_X1   g0615(.A1(new_n814), .A2(new_n815), .ZN(new_n816));
  XNOR2_X1  g0616(.A(new_n816), .B(KEYINPUT93), .ZN(new_n817));
  NAND2_X1  g0617(.A1(new_n817), .A2(KEYINPUT32), .ZN(new_n818));
  OR2_X1    g0618(.A1(new_n817), .A2(KEYINPUT32), .ZN(new_n819));
  NAND3_X1  g0619(.A1(new_n812), .A2(G190), .A3(G200), .ZN(new_n820));
  NOR2_X1   g0620(.A1(new_n820), .A2(new_n309), .ZN(new_n821));
  NOR2_X1   g0621(.A1(new_n803), .A2(G190), .ZN(new_n822));
  INV_X1    g0622(.A(new_n822), .ZN(new_n823));
  NAND3_X1  g0623(.A1(new_n358), .A2(new_n322), .A3(G190), .ZN(new_n824));
  NAND2_X1  g0624(.A1(new_n824), .A2(G20), .ZN(new_n825));
  INV_X1    g0625(.A(new_n825), .ZN(new_n826));
  OAI22_X1  g0626(.A1(new_n823), .A2(new_n400), .B1(new_n826), .B2(new_n552), .ZN(new_n827));
  NAND3_X1  g0627(.A1(new_n812), .A2(new_n447), .A3(G200), .ZN(new_n828));
  INV_X1    g0628(.A(new_n828), .ZN(new_n829));
  AOI211_X1 g0629(.A(new_n821), .B(new_n827), .C1(G107), .C2(new_n829), .ZN(new_n830));
  NAND4_X1  g0630(.A1(new_n811), .A2(new_n818), .A3(new_n819), .A4(new_n830), .ZN(new_n831));
  INV_X1    g0631(.A(new_n814), .ZN(new_n832));
  AOI21_X1  g0632(.A(new_n281), .B1(new_n832), .B2(G329), .ZN(new_n833));
  INV_X1    g0633(.A(G283), .ZN(new_n834));
  OAI21_X1  g0634(.A(new_n833), .B1(new_n834), .B2(new_n828), .ZN(new_n835));
  AOI21_X1  g0635(.A(new_n835), .B1(new_n807), .B2(G322), .ZN(new_n836));
  NOR2_X1   g0636(.A1(new_n529), .A2(new_n530), .ZN(new_n837));
  INV_X1    g0637(.A(new_n837), .ZN(new_n838));
  AOI22_X1  g0638(.A1(new_n804), .A2(G326), .B1(new_n825), .B2(new_n838), .ZN(new_n839));
  XNOR2_X1  g0639(.A(KEYINPUT33), .B(G317), .ZN(new_n840));
  INV_X1    g0640(.A(new_n820), .ZN(new_n841));
  AOI22_X1  g0641(.A1(new_n822), .A2(new_n840), .B1(new_n841), .B2(G303), .ZN(new_n842));
  NAND2_X1  g0642(.A1(new_n810), .A2(G311), .ZN(new_n843));
  NAND4_X1  g0643(.A1(new_n836), .A2(new_n839), .A3(new_n842), .A4(new_n843), .ZN(new_n844));
  NAND2_X1  g0644(.A1(new_n831), .A2(new_n844), .ZN(new_n845));
  AOI21_X1  g0645(.A(new_n801), .B1(new_n845), .B2(new_n793), .ZN(new_n846));
  OAI21_X1  g0646(.A(new_n846), .B1(new_n720), .B2(new_n798), .ZN(new_n847));
  AND2_X1   g0647(.A1(new_n782), .A2(new_n847), .ZN(new_n848));
  INV_X1    g0648(.A(new_n848), .ZN(G396));
  AOI21_X1  g0649(.A(new_n718), .B1(new_n691), .B2(new_n708), .ZN(new_n850));
  OAI21_X1  g0650(.A(KEYINPUT96), .B1(new_n360), .B2(new_n361), .ZN(new_n851));
  INV_X1    g0651(.A(KEYINPUT96), .ZN(new_n852));
  NAND4_X1  g0652(.A1(new_n321), .A2(new_n357), .A3(new_n852), .A4(new_n359), .ZN(new_n853));
  NAND3_X1  g0653(.A1(new_n355), .A2(new_n851), .A3(new_n853), .ZN(new_n854));
  INV_X1    g0654(.A(new_n854), .ZN(new_n855));
  NAND2_X1  g0655(.A1(new_n850), .A2(new_n855), .ZN(new_n856));
  NAND2_X1  g0656(.A1(new_n321), .A2(new_n718), .ZN(new_n857));
  NAND4_X1  g0657(.A1(new_n355), .A2(new_n851), .A3(new_n857), .A4(new_n853), .ZN(new_n858));
  NAND2_X1  g0658(.A1(new_n362), .A2(new_n718), .ZN(new_n859));
  NAND2_X1  g0659(.A1(new_n858), .A2(new_n859), .ZN(new_n860));
  OAI21_X1  g0660(.A(new_n856), .B1(new_n850), .B2(new_n860), .ZN(new_n861));
  NAND2_X1  g0661(.A1(new_n773), .A2(G330), .ZN(new_n862));
  AOI21_X1  g0662(.A(new_n780), .B1(new_n861), .B2(new_n862), .ZN(new_n863));
  OAI21_X1  g0663(.A(new_n863), .B1(new_n862), .B2(new_n861), .ZN(new_n864));
  NAND2_X1  g0664(.A1(new_n794), .A2(new_n796), .ZN(new_n865));
  OAI21_X1  g0665(.A(new_n780), .B1(G77), .B2(new_n865), .ZN(new_n866));
  INV_X1    g0666(.A(new_n810), .ZN(new_n867));
  OAI221_X1 g0667(.A(new_n328), .B1(new_n552), .B2(new_n826), .C1(new_n867), .C2(new_n636), .ZN(new_n868));
  AOI21_X1  g0668(.A(new_n868), .B1(G294), .B2(new_n807), .ZN(new_n869));
  INV_X1    g0669(.A(G311), .ZN(new_n870));
  OAI22_X1  g0670(.A1(new_n828), .A2(new_n309), .B1(new_n814), .B2(new_n870), .ZN(new_n871));
  XOR2_X1   g0671(.A(new_n871), .B(KEYINPUT94), .Z(new_n872));
  OAI22_X1  g0672(.A1(new_n823), .A2(new_n834), .B1(new_n820), .B2(new_n342), .ZN(new_n873));
  AOI21_X1  g0673(.A(new_n873), .B1(G303), .B2(new_n804), .ZN(new_n874));
  NAND3_X1  g0674(.A1(new_n869), .A2(new_n872), .A3(new_n874), .ZN(new_n875));
  AOI22_X1  g0675(.A1(G137), .A2(new_n804), .B1(new_n822), .B2(G150), .ZN(new_n876));
  XNOR2_X1  g0676(.A(new_n876), .B(KEYINPUT95), .ZN(new_n877));
  INV_X1    g0677(.A(G143), .ZN(new_n878));
  OAI221_X1 g0678(.A(new_n877), .B1(new_n878), .B2(new_n808), .C1(new_n815), .C2(new_n867), .ZN(new_n879));
  XOR2_X1   g0679(.A(new_n879), .B(KEYINPUT34), .Z(new_n880));
  NAND2_X1  g0680(.A1(new_n829), .A2(G68), .ZN(new_n881));
  OAI21_X1  g0681(.A(new_n881), .B1(new_n253), .B2(new_n820), .ZN(new_n882));
  INV_X1    g0682(.A(G132), .ZN(new_n883));
  OAI221_X1 g0683(.A(new_n281), .B1(new_n814), .B2(new_n883), .C1(new_n826), .C2(new_n302), .ZN(new_n884));
  OR2_X1    g0684(.A1(new_n882), .A2(new_n884), .ZN(new_n885));
  OAI21_X1  g0685(.A(new_n875), .B1(new_n880), .B2(new_n885), .ZN(new_n886));
  AOI21_X1  g0686(.A(new_n866), .B1(new_n886), .B2(new_n793), .ZN(new_n887));
  OAI21_X1  g0687(.A(new_n887), .B1(new_n796), .B2(new_n860), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n864), .A2(new_n888), .ZN(G384));
  NOR2_X1   g0689(.A1(new_n777), .A2(new_n256), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n761), .A2(new_n771), .ZN(new_n891));
  NAND3_X1  g0691(.A1(new_n765), .A2(new_n764), .A3(new_n891), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n466), .A2(new_n718), .ZN(new_n893));
  NAND3_X1  g0693(.A1(new_n465), .A2(new_n472), .A3(new_n893), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n461), .A2(G169), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n895), .A2(KEYINPUT14), .ZN(new_n896));
  NAND3_X1  g0696(.A1(new_n896), .A2(new_n469), .A3(new_n468), .ZN(new_n897));
  OAI211_X1 g0697(.A(new_n466), .B(new_n718), .C1(new_n897), .C2(new_n464), .ZN(new_n898));
  AOI22_X1  g0698(.A1(new_n894), .A2(new_n898), .B1(new_n858), .B2(new_n859), .ZN(new_n899));
  AND3_X1   g0699(.A1(new_n892), .A2(new_n899), .A3(KEYINPUT40), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n432), .A2(new_n433), .ZN(new_n901));
  INV_X1    g0701(.A(new_n716), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n432), .A2(new_n902), .ZN(new_n903));
  NAND3_X1  g0703(.A1(new_n901), .A2(new_n903), .A3(new_n667), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n904), .A2(KEYINPUT37), .ZN(new_n905));
  INV_X1    g0705(.A(KEYINPUT98), .ZN(new_n906));
  AOI21_X1  g0706(.A(new_n416), .B1(new_n661), .B2(new_n387), .ZN(new_n907));
  AOI21_X1  g0707(.A(new_n907), .B1(new_n409), .B2(new_n385), .ZN(new_n908));
  AOI21_X1  g0708(.A(KEYINPUT37), .B1(new_n432), .B2(new_n902), .ZN(new_n909));
  AOI21_X1  g0709(.A(new_n906), .B1(new_n908), .B2(new_n909), .ZN(new_n910));
  NAND4_X1  g0710(.A1(new_n909), .A2(new_n906), .A3(new_n901), .A4(new_n667), .ZN(new_n911));
  INV_X1    g0711(.A(new_n911), .ZN(new_n912));
  OAI21_X1  g0712(.A(new_n905), .B1(new_n910), .B2(new_n912), .ZN(new_n913));
  AOI21_X1  g0713(.A(new_n903), .B1(new_n412), .B2(new_n435), .ZN(new_n914));
  INV_X1    g0714(.A(new_n914), .ZN(new_n915));
  AOI21_X1  g0715(.A(KEYINPUT38), .B1(new_n913), .B2(new_n915), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n901), .A2(new_n667), .ZN(new_n917));
  INV_X1    g0717(.A(KEYINPUT37), .ZN(new_n918));
  OAI21_X1  g0718(.A(new_n918), .B1(new_n409), .B2(new_n716), .ZN(new_n919));
  OAI21_X1  g0719(.A(KEYINPUT98), .B1(new_n917), .B2(new_n919), .ZN(new_n920));
  NOR2_X1   g0720(.A1(new_n396), .A2(new_n398), .ZN(new_n921));
  OAI21_X1  g0721(.A(new_n387), .B1(new_n425), .B2(new_n921), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n922), .A2(new_n433), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n922), .A2(new_n902), .ZN(new_n924));
  NAND3_X1  g0724(.A1(new_n923), .A2(new_n924), .A3(new_n667), .ZN(new_n925));
  AOI22_X1  g0725(.A1(new_n920), .A2(new_n911), .B1(KEYINPUT37), .B2(new_n925), .ZN(new_n926));
  AOI21_X1  g0726(.A(new_n924), .B1(new_n412), .B2(new_n435), .ZN(new_n927));
  INV_X1    g0727(.A(KEYINPUT38), .ZN(new_n928));
  NOR3_X1   g0728(.A1(new_n926), .A2(new_n927), .A3(new_n928), .ZN(new_n929));
  OAI21_X1  g0729(.A(new_n900), .B1(new_n916), .B2(new_n929), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n930), .A2(KEYINPUT100), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n925), .A2(KEYINPUT37), .ZN(new_n932));
  OAI21_X1  g0732(.A(new_n932), .B1(new_n910), .B2(new_n912), .ZN(new_n933));
  INV_X1    g0733(.A(new_n924), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n436), .A2(new_n934), .ZN(new_n935));
  NAND3_X1  g0735(.A1(new_n933), .A2(KEYINPUT38), .A3(new_n935), .ZN(new_n936));
  AOI22_X1  g0736(.A1(new_n920), .A2(new_n911), .B1(KEYINPUT37), .B2(new_n904), .ZN(new_n937));
  OAI21_X1  g0737(.A(new_n928), .B1(new_n937), .B2(new_n914), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n936), .A2(new_n938), .ZN(new_n939));
  INV_X1    g0739(.A(KEYINPUT100), .ZN(new_n940));
  NAND3_X1  g0740(.A1(new_n939), .A2(new_n940), .A3(new_n900), .ZN(new_n941));
  INV_X1    g0741(.A(KEYINPUT40), .ZN(new_n942));
  AND2_X1   g0742(.A1(new_n892), .A2(new_n899), .ZN(new_n943));
  AOI21_X1  g0743(.A(KEYINPUT38), .B1(new_n933), .B2(new_n935), .ZN(new_n944));
  OAI21_X1  g0744(.A(new_n943), .B1(new_n944), .B2(new_n929), .ZN(new_n945));
  AOI22_X1  g0745(.A1(new_n931), .A2(new_n941), .B1(new_n942), .B2(new_n945), .ZN(new_n946));
  XNOR2_X1  g0746(.A(new_n946), .B(KEYINPUT101), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n474), .A2(new_n892), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n947), .A2(new_n948), .ZN(new_n949));
  NAND2_X1  g0749(.A1(new_n949), .A2(G330), .ZN(new_n950));
  OR2_X1    g0750(.A1(new_n950), .A2(KEYINPUT102), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n950), .A2(KEYINPUT102), .ZN(new_n952));
  OAI211_X1 g0752(.A(new_n951), .B(new_n952), .C1(new_n948), .C2(new_n947), .ZN(new_n953));
  OAI21_X1  g0753(.A(new_n474), .B1(new_n744), .B2(new_n743), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n678), .A2(new_n954), .ZN(new_n955));
  XNOR2_X1  g0755(.A(new_n955), .B(KEYINPUT99), .ZN(new_n956));
  NAND2_X1  g0756(.A1(new_n894), .A2(new_n898), .ZN(new_n957));
  INV_X1    g0757(.A(new_n957), .ZN(new_n958));
  AND2_X1   g0758(.A1(new_n851), .A2(new_n853), .ZN(new_n959));
  NOR2_X1   g0759(.A1(new_n959), .A2(new_n718), .ZN(new_n960));
  INV_X1    g0760(.A(new_n960), .ZN(new_n961));
  AOI21_X1  g0761(.A(new_n958), .B1(new_n856), .B2(new_n961), .ZN(new_n962));
  OAI21_X1  g0762(.A(new_n928), .B1(new_n926), .B2(new_n927), .ZN(new_n963));
  NAND2_X1  g0763(.A1(new_n936), .A2(new_n963), .ZN(new_n964));
  AOI22_X1  g0764(.A1(new_n962), .A2(new_n964), .B1(new_n671), .B2(new_n716), .ZN(new_n965));
  INV_X1    g0765(.A(KEYINPUT39), .ZN(new_n966));
  OAI21_X1  g0766(.A(new_n966), .B1(new_n916), .B2(new_n929), .ZN(new_n967));
  NAND3_X1  g0767(.A1(new_n897), .A2(new_n466), .A3(new_n724), .ZN(new_n968));
  INV_X1    g0768(.A(new_n968), .ZN(new_n969));
  NAND3_X1  g0769(.A1(new_n936), .A2(new_n963), .A3(KEYINPUT39), .ZN(new_n970));
  NAND3_X1  g0770(.A1(new_n967), .A2(new_n969), .A3(new_n970), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n965), .A2(new_n971), .ZN(new_n972));
  XNOR2_X1  g0772(.A(new_n956), .B(new_n972), .ZN(new_n973));
  AOI21_X1  g0773(.A(new_n890), .B1(new_n953), .B2(new_n973), .ZN(new_n974));
  OAI21_X1  g0774(.A(new_n974), .B1(new_n973), .B2(new_n953), .ZN(new_n975));
  OAI21_X1  g0775(.A(G77), .B1(new_n302), .B2(new_n400), .ZN(new_n976));
  OAI22_X1  g0776(.A1(new_n976), .A2(new_n223), .B1(G50), .B2(new_n400), .ZN(new_n977));
  NAND3_X1  g0777(.A1(new_n977), .A2(G1), .A3(new_n776), .ZN(new_n978));
  XNOR2_X1  g0778(.A(new_n978), .B(KEYINPUT97), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n222), .A2(G116), .ZN(new_n980));
  AOI21_X1  g0780(.A(new_n980), .B1(new_n608), .B2(KEYINPUT35), .ZN(new_n981));
  OAI21_X1  g0781(.A(new_n981), .B1(KEYINPUT35), .B2(new_n608), .ZN(new_n982));
  INV_X1    g0782(.A(KEYINPUT36), .ZN(new_n983));
  OAI21_X1  g0783(.A(new_n979), .B1(new_n982), .B2(new_n983), .ZN(new_n984));
  AOI21_X1  g0784(.A(new_n984), .B1(new_n983), .B2(new_n982), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n975), .A2(new_n985), .ZN(G367));
  NOR2_X1   g0786(.A1(new_n699), .A2(new_n724), .ZN(new_n987));
  AND2_X1   g0787(.A1(new_n614), .A2(new_n623), .ZN(new_n988));
  NAND2_X1  g0788(.A1(new_n698), .A2(new_n718), .ZN(new_n989));
  AOI21_X1  g0789(.A(new_n987), .B1(new_n988), .B2(new_n989), .ZN(new_n990));
  OAI21_X1  g0790(.A(new_n614), .B1(new_n990), .B2(new_n688), .ZN(new_n991));
  NAND2_X1  g0791(.A1(new_n991), .A2(new_n724), .ZN(new_n992));
  OAI21_X1  g0792(.A(KEYINPUT42), .B1(new_n990), .B2(new_n729), .ZN(new_n993));
  OR3_X1    g0793(.A1(new_n990), .A2(new_n729), .A3(KEYINPUT42), .ZN(new_n994));
  NAND3_X1  g0794(.A1(new_n992), .A2(new_n993), .A3(new_n994), .ZN(new_n995));
  NAND2_X1  g0795(.A1(new_n579), .A2(new_n580), .ZN(new_n996));
  NAND2_X1  g0796(.A1(new_n996), .A2(new_n718), .ZN(new_n997));
  NAND2_X1  g0797(.A1(new_n582), .A2(new_n997), .ZN(new_n998));
  OAI21_X1  g0798(.A(new_n998), .B1(new_n576), .B2(new_n997), .ZN(new_n999));
  NAND2_X1  g0799(.A1(new_n999), .A2(KEYINPUT43), .ZN(new_n1000));
  NAND2_X1  g0800(.A1(new_n995), .A2(new_n1000), .ZN(new_n1001));
  NOR2_X1   g0801(.A1(new_n999), .A2(KEYINPUT43), .ZN(new_n1002));
  OR2_X1    g0802(.A1(new_n1001), .A2(new_n1002), .ZN(new_n1003));
  NAND2_X1  g0803(.A1(new_n1001), .A2(new_n1002), .ZN(new_n1004));
  NAND2_X1  g0804(.A1(new_n1003), .A2(new_n1004), .ZN(new_n1005));
  NOR2_X1   g0805(.A1(new_n727), .A2(new_n990), .ZN(new_n1006));
  XNOR2_X1  g0806(.A(new_n1005), .B(new_n1006), .ZN(new_n1007));
  XOR2_X1   g0807(.A(new_n734), .B(KEYINPUT41), .Z(new_n1008));
  NAND2_X1  g0808(.A1(new_n729), .A2(new_n728), .ZN(new_n1009));
  NAND2_X1  g0809(.A1(new_n1009), .A2(new_n990), .ZN(new_n1010));
  XOR2_X1   g0810(.A(new_n1010), .B(KEYINPUT44), .Z(new_n1011));
  NOR2_X1   g0811(.A1(new_n1009), .A2(new_n990), .ZN(new_n1012));
  XNOR2_X1  g0812(.A(new_n1012), .B(KEYINPUT45), .ZN(new_n1013));
  NAND2_X1  g0813(.A1(new_n1011), .A2(new_n1013), .ZN(new_n1014));
  NOR2_X1   g0814(.A1(new_n727), .A2(KEYINPUT103), .ZN(new_n1015));
  OR2_X1    g0815(.A1(new_n1014), .A2(new_n1015), .ZN(new_n1016));
  NOR2_X1   g0816(.A1(new_n689), .A2(new_n718), .ZN(new_n1017));
  OAI21_X1  g0817(.A(new_n729), .B1(new_n726), .B2(new_n1017), .ZN(new_n1018));
  XNOR2_X1  g0818(.A(new_n1018), .B(new_n721), .ZN(new_n1019));
  INV_X1    g0819(.A(new_n1019), .ZN(new_n1020));
  AND2_X1   g0820(.A1(new_n1020), .A2(new_n774), .ZN(new_n1021));
  NAND2_X1  g0821(.A1(new_n1014), .A2(new_n1015), .ZN(new_n1022));
  NAND3_X1  g0822(.A1(new_n1016), .A2(new_n1021), .A3(new_n1022), .ZN(new_n1023));
  AOI21_X1  g0823(.A(new_n1008), .B1(new_n1023), .B2(new_n774), .ZN(new_n1024));
  OAI21_X1  g0824(.A(new_n1007), .B1(new_n1024), .B2(new_n779), .ZN(new_n1025));
  INV_X1    g0825(.A(new_n800), .ZN(new_n1026));
  AOI22_X1  g0826(.A1(new_n785), .A2(new_n234), .B1(new_n733), .B2(new_n557), .ZN(new_n1027));
  AOI211_X1 g0827(.A(new_n734), .B(new_n779), .C1(new_n1026), .C2(new_n1027), .ZN(new_n1028));
  NAND2_X1  g0828(.A1(new_n825), .A2(G68), .ZN(new_n1029));
  INV_X1    g0829(.A(G137), .ZN(new_n1030));
  OAI221_X1 g0830(.A(new_n1029), .B1(new_n1030), .B2(new_n814), .C1(new_n808), .C2(new_n248), .ZN(new_n1031));
  AOI21_X1  g0831(.A(new_n1031), .B1(G50), .B2(new_n810), .ZN(new_n1032));
  AOI21_X1  g0832(.A(new_n328), .B1(new_n829), .B2(G77), .ZN(new_n1033));
  OR2_X1    g0833(.A1(new_n1033), .A2(KEYINPUT106), .ZN(new_n1034));
  NAND2_X1  g0834(.A1(new_n1033), .A2(KEYINPUT106), .ZN(new_n1035));
  OAI22_X1  g0835(.A1(new_n823), .A2(new_n815), .B1(new_n820), .B2(new_n302), .ZN(new_n1036));
  AOI21_X1  g0836(.A(new_n1036), .B1(G143), .B2(new_n804), .ZN(new_n1037));
  NAND4_X1  g0837(.A1(new_n1032), .A2(new_n1034), .A3(new_n1035), .A4(new_n1037), .ZN(new_n1038));
  NOR2_X1   g0838(.A1(new_n820), .A2(new_n636), .ZN(new_n1039));
  NOR2_X1   g0839(.A1(new_n1039), .A2(KEYINPUT46), .ZN(new_n1040));
  XNOR2_X1  g0840(.A(new_n1040), .B(KEYINPUT104), .ZN(new_n1041));
  AOI22_X1  g0841(.A1(KEYINPUT46), .A2(new_n1039), .B1(new_n822), .B2(new_n838), .ZN(new_n1042));
  AOI21_X1  g0842(.A(KEYINPUT105), .B1(new_n1041), .B2(new_n1042), .ZN(new_n1043));
  OAI22_X1  g0843(.A1(new_n834), .A2(new_n867), .B1(new_n808), .B2(new_n628), .ZN(new_n1044));
  INV_X1    g0844(.A(G317), .ZN(new_n1045));
  OAI221_X1 g0845(.A(new_n328), .B1(new_n814), .B2(new_n1045), .C1(new_n552), .C2(new_n828), .ZN(new_n1046));
  OAI22_X1  g0846(.A1(new_n805), .A2(new_n870), .B1(new_n826), .B2(new_n342), .ZN(new_n1047));
  NOR3_X1   g0847(.A1(new_n1044), .A2(new_n1046), .A3(new_n1047), .ZN(new_n1048));
  NAND3_X1  g0848(.A1(new_n1041), .A2(KEYINPUT105), .A3(new_n1042), .ZN(new_n1049));
  NAND2_X1  g0849(.A1(new_n1048), .A2(new_n1049), .ZN(new_n1050));
  OAI21_X1  g0850(.A(new_n1038), .B1(new_n1043), .B2(new_n1050), .ZN(new_n1051));
  XOR2_X1   g0851(.A(new_n1051), .B(KEYINPUT47), .Z(new_n1052));
  OAI221_X1 g0852(.A(new_n1028), .B1(new_n798), .B2(new_n999), .C1(new_n1052), .C2(new_n794), .ZN(new_n1053));
  NAND2_X1  g0853(.A1(new_n1025), .A2(new_n1053), .ZN(G387));
  INV_X1    g0854(.A(new_n734), .ZN(new_n1055));
  NOR2_X1   g0855(.A1(new_n1021), .A2(new_n1055), .ZN(new_n1056));
  OAI21_X1  g0856(.A(new_n1056), .B1(new_n774), .B2(new_n1020), .ZN(new_n1057));
  NAND3_X1  g0857(.A1(new_n231), .A2(G45), .A3(new_n328), .ZN(new_n1058));
  OAI21_X1  g0858(.A(KEYINPUT50), .B1(new_n246), .B2(G50), .ZN(new_n1059));
  OAI211_X1 g0859(.A(new_n1059), .B(new_n509), .C1(new_n400), .C2(new_n294), .ZN(new_n1060));
  NOR3_X1   g0860(.A1(new_n246), .A2(KEYINPUT50), .A3(G50), .ZN(new_n1061));
  OAI21_X1  g0861(.A(new_n328), .B1(new_n1060), .B2(new_n1061), .ZN(new_n1062));
  NAND2_X1  g0862(.A1(new_n1062), .A2(new_n731), .ZN(new_n1063));
  AOI21_X1  g0863(.A(new_n733), .B1(new_n1058), .B2(new_n1063), .ZN(new_n1064));
  OAI21_X1  g0864(.A(new_n1026), .B1(new_n342), .B2(new_n217), .ZN(new_n1065));
  OAI21_X1  g0865(.A(new_n780), .B1(new_n1064), .B2(new_n1065), .ZN(new_n1066));
  NOR2_X1   g0866(.A1(new_n826), .A2(new_n348), .ZN(new_n1067));
  OAI22_X1  g0867(.A1(new_n805), .A2(new_n815), .B1(new_n820), .B2(new_n294), .ZN(new_n1068));
  AOI211_X1 g0868(.A(new_n1067), .B(new_n1068), .C1(new_n306), .C2(new_n822), .ZN(new_n1069));
  OAI221_X1 g0869(.A(new_n281), .B1(new_n814), .B2(new_n248), .C1(new_n552), .C2(new_n828), .ZN(new_n1070));
  AOI21_X1  g0870(.A(new_n1070), .B1(new_n807), .B2(G50), .ZN(new_n1071));
  OAI211_X1 g0871(.A(new_n1069), .B(new_n1071), .C1(new_n400), .C2(new_n867), .ZN(new_n1072));
  AOI21_X1  g0872(.A(new_n281), .B1(new_n832), .B2(G326), .ZN(new_n1073));
  OAI22_X1  g0873(.A1(new_n826), .A2(new_n834), .B1(new_n837), .B2(new_n820), .ZN(new_n1074));
  AOI22_X1  g0874(.A1(G311), .A2(new_n822), .B1(new_n804), .B2(G322), .ZN(new_n1075));
  OAI221_X1 g0875(.A(new_n1075), .B1(new_n867), .B2(new_n628), .C1(new_n1045), .C2(new_n808), .ZN(new_n1076));
  INV_X1    g0876(.A(KEYINPUT48), .ZN(new_n1077));
  AOI21_X1  g0877(.A(new_n1074), .B1(new_n1076), .B2(new_n1077), .ZN(new_n1078));
  OAI21_X1  g0878(.A(new_n1078), .B1(new_n1077), .B2(new_n1076), .ZN(new_n1079));
  INV_X1    g0879(.A(KEYINPUT49), .ZN(new_n1080));
  OAI221_X1 g0880(.A(new_n1073), .B1(new_n636), .B2(new_n828), .C1(new_n1079), .C2(new_n1080), .ZN(new_n1081));
  AND2_X1   g0881(.A1(new_n1079), .A2(new_n1080), .ZN(new_n1082));
  OAI21_X1  g0882(.A(new_n1072), .B1(new_n1081), .B2(new_n1082), .ZN(new_n1083));
  AOI21_X1  g0883(.A(new_n1066), .B1(new_n1083), .B2(new_n793), .ZN(new_n1084));
  OR2_X1    g0884(.A1(new_n726), .A2(new_n798), .ZN(new_n1085));
  AOI22_X1  g0885(.A1(new_n1020), .A2(new_n779), .B1(new_n1084), .B2(new_n1085), .ZN(new_n1086));
  NAND2_X1  g0886(.A1(new_n1057), .A2(new_n1086), .ZN(G393));
  XNOR2_X1  g0887(.A(new_n1014), .B(new_n727), .ZN(new_n1088));
  OAI211_X1 g0888(.A(new_n1023), .B(new_n734), .C1(new_n1088), .C2(new_n1021), .ZN(new_n1089));
  NAND2_X1  g0889(.A1(new_n990), .A2(new_n797), .ZN(new_n1090));
  OAI21_X1  g0890(.A(new_n1026), .B1(new_n552), .B2(new_n217), .ZN(new_n1091));
  NOR2_X1   g0891(.A1(new_n239), .A2(new_n786), .ZN(new_n1092));
  OAI21_X1  g0892(.A(new_n780), .B1(new_n1091), .B2(new_n1092), .ZN(new_n1093));
  AOI22_X1  g0893(.A1(new_n807), .A2(G159), .B1(G150), .B2(new_n804), .ZN(new_n1094));
  XOR2_X1   g0894(.A(new_n1094), .B(KEYINPUT51), .Z(new_n1095));
  OAI22_X1  g0895(.A1(new_n823), .A2(new_n253), .B1(new_n826), .B2(new_n294), .ZN(new_n1096));
  AOI21_X1  g0896(.A(new_n1096), .B1(G68), .B2(new_n841), .ZN(new_n1097));
  OAI221_X1 g0897(.A(new_n281), .B1(new_n814), .B2(new_n878), .C1(new_n309), .C2(new_n828), .ZN(new_n1098));
  AOI21_X1  g0898(.A(new_n1098), .B1(new_n810), .B2(new_n306), .ZN(new_n1099));
  NAND3_X1  g0899(.A1(new_n1095), .A2(new_n1097), .A3(new_n1099), .ZN(new_n1100));
  AOI22_X1  g0900(.A1(new_n807), .A2(G311), .B1(G317), .B2(new_n804), .ZN(new_n1101));
  XNOR2_X1  g0901(.A(new_n1101), .B(KEYINPUT52), .ZN(new_n1102));
  AOI21_X1  g0902(.A(new_n281), .B1(new_n832), .B2(G322), .ZN(new_n1103));
  INV_X1    g0903(.A(G294), .ZN(new_n1104));
  OAI221_X1 g0904(.A(new_n1103), .B1(new_n342), .B2(new_n828), .C1(new_n867), .C2(new_n1104), .ZN(new_n1105));
  NOR2_X1   g0905(.A1(new_n820), .A2(new_n834), .ZN(new_n1106));
  OAI22_X1  g0906(.A1(new_n823), .A2(new_n628), .B1(new_n826), .B2(new_n636), .ZN(new_n1107));
  OR3_X1    g0907(.A1(new_n1105), .A2(new_n1106), .A3(new_n1107), .ZN(new_n1108));
  OAI21_X1  g0908(.A(new_n1100), .B1(new_n1102), .B2(new_n1108), .ZN(new_n1109));
  XOR2_X1   g0909(.A(new_n1109), .B(KEYINPUT107), .Z(new_n1110));
  AOI21_X1  g0910(.A(new_n1093), .B1(new_n1110), .B2(new_n793), .ZN(new_n1111));
  AOI22_X1  g0911(.A1(new_n1088), .A2(new_n779), .B1(new_n1090), .B2(new_n1111), .ZN(new_n1112));
  NAND2_X1  g0912(.A1(new_n1089), .A2(new_n1112), .ZN(G390));
  AOI22_X1  g0913(.A1(new_n807), .A2(G116), .B1(G77), .B2(new_n825), .ZN(new_n1114));
  XNOR2_X1  g0914(.A(new_n1114), .B(KEYINPUT114), .ZN(new_n1115));
  AOI211_X1 g0915(.A(new_n281), .B(new_n821), .C1(G294), .C2(new_n832), .ZN(new_n1116));
  OAI21_X1  g0916(.A(new_n1116), .B1(new_n867), .B2(new_n552), .ZN(new_n1117));
  OAI221_X1 g0917(.A(new_n881), .B1(new_n805), .B2(new_n834), .C1(new_n342), .C2(new_n823), .ZN(new_n1118));
  NOR3_X1   g0918(.A1(new_n1115), .A2(new_n1117), .A3(new_n1118), .ZN(new_n1119));
  INV_X1    g0919(.A(new_n1119), .ZN(new_n1120));
  OR2_X1    g0920(.A1(new_n1120), .A2(KEYINPUT115), .ZN(new_n1121));
  INV_X1    g0921(.A(G128), .ZN(new_n1122));
  OAI22_X1  g0922(.A1(new_n805), .A2(new_n1122), .B1(new_n826), .B2(new_n815), .ZN(new_n1123));
  AOI21_X1  g0923(.A(new_n1123), .B1(G137), .B2(new_n822), .ZN(new_n1124));
  AOI21_X1  g0924(.A(new_n328), .B1(new_n832), .B2(G125), .ZN(new_n1125));
  OAI21_X1  g0925(.A(new_n1125), .B1(new_n253), .B2(new_n828), .ZN(new_n1126));
  XNOR2_X1  g0926(.A(KEYINPUT54), .B(G143), .ZN(new_n1127));
  INV_X1    g0927(.A(new_n1127), .ZN(new_n1128));
  AOI21_X1  g0928(.A(new_n1126), .B1(new_n810), .B2(new_n1128), .ZN(new_n1129));
  NAND2_X1  g0929(.A1(new_n807), .A2(G132), .ZN(new_n1130));
  NOR2_X1   g0930(.A1(new_n820), .A2(new_n248), .ZN(new_n1131));
  XNOR2_X1  g0931(.A(KEYINPUT113), .B(KEYINPUT53), .ZN(new_n1132));
  XNOR2_X1  g0932(.A(new_n1131), .B(new_n1132), .ZN(new_n1133));
  NAND4_X1  g0933(.A1(new_n1124), .A2(new_n1129), .A3(new_n1130), .A4(new_n1133), .ZN(new_n1134));
  NAND2_X1  g0934(.A1(new_n1120), .A2(KEYINPUT115), .ZN(new_n1135));
  AND3_X1   g0935(.A1(new_n1121), .A2(new_n1134), .A3(new_n1135), .ZN(new_n1136));
  OAI221_X1 g0936(.A(new_n780), .B1(new_n306), .B2(new_n865), .C1(new_n1136), .C2(new_n794), .ZN(new_n1137));
  NAND2_X1  g0937(.A1(new_n967), .A2(new_n970), .ZN(new_n1138));
  AOI21_X1  g0938(.A(new_n1137), .B1(new_n1138), .B2(new_n795), .ZN(new_n1139));
  NAND3_X1  g0939(.A1(new_n892), .A2(new_n899), .A3(G330), .ZN(new_n1140));
  INV_X1    g0940(.A(KEYINPUT109), .ZN(new_n1141));
  NAND2_X1  g0941(.A1(new_n1140), .A2(new_n1141), .ZN(new_n1142));
  INV_X1    g0942(.A(G330), .ZN(new_n1143));
  AOI22_X1  g0943(.A1(new_n762), .A2(new_n763), .B1(new_n771), .B2(new_n761), .ZN(new_n1144));
  AOI21_X1  g0944(.A(new_n1143), .B1(new_n1144), .B2(new_n765), .ZN(new_n1145));
  NAND3_X1  g0945(.A1(new_n1145), .A2(KEYINPUT109), .A3(new_n899), .ZN(new_n1146));
  NAND2_X1  g0946(.A1(new_n1142), .A2(new_n1146), .ZN(new_n1147));
  AOI211_X1 g0947(.A(new_n718), .B(new_n854), .C1(new_n691), .C2(new_n708), .ZN(new_n1148));
  OAI21_X1  g0948(.A(new_n957), .B1(new_n1148), .B2(new_n960), .ZN(new_n1149));
  AOI22_X1  g0949(.A1(new_n967), .A2(new_n970), .B1(new_n1149), .B2(new_n968), .ZN(new_n1150));
  NAND3_X1  g0950(.A1(new_n742), .A2(new_n724), .A3(new_n855), .ZN(new_n1151));
  NAND2_X1  g0951(.A1(new_n1151), .A2(new_n961), .ZN(new_n1152));
  NAND2_X1  g0952(.A1(new_n1152), .A2(new_n957), .ZN(new_n1153));
  XNOR2_X1  g0953(.A(new_n968), .B(KEYINPUT108), .ZN(new_n1154));
  AND3_X1   g0954(.A1(new_n1153), .A2(new_n939), .A3(new_n1154), .ZN(new_n1155));
  OAI21_X1  g0955(.A(new_n1147), .B1(new_n1150), .B2(new_n1155), .ZN(new_n1156));
  AND3_X1   g0956(.A1(new_n936), .A2(new_n963), .A3(KEYINPUT39), .ZN(new_n1157));
  AOI21_X1  g0957(.A(KEYINPUT39), .B1(new_n936), .B2(new_n938), .ZN(new_n1158));
  OAI22_X1  g0958(.A1(new_n1157), .A2(new_n1158), .B1(new_n962), .B2(new_n969), .ZN(new_n1159));
  NAND3_X1  g0959(.A1(new_n1153), .A2(new_n939), .A3(new_n1154), .ZN(new_n1160));
  NAND2_X1  g0960(.A1(new_n765), .A2(new_n764), .ZN(new_n1161));
  INV_X1    g0961(.A(new_n757), .ZN(new_n1162));
  AOI21_X1  g0962(.A(new_n1162), .B1(new_n766), .B2(new_n767), .ZN(new_n1163));
  AOI21_X1  g0963(.A(new_n772), .B1(new_n1163), .B2(new_n769), .ZN(new_n1164));
  OAI211_X1 g0964(.A(new_n899), .B(G330), .C1(new_n1161), .C2(new_n1164), .ZN(new_n1165));
  NAND2_X1  g0965(.A1(new_n1165), .A2(KEYINPUT111), .ZN(new_n1166));
  INV_X1    g0966(.A(KEYINPUT111), .ZN(new_n1167));
  NAND4_X1  g0967(.A1(new_n773), .A2(new_n1167), .A3(G330), .A4(new_n899), .ZN(new_n1168));
  NAND2_X1  g0968(.A1(new_n1166), .A2(new_n1168), .ZN(new_n1169));
  NAND3_X1  g0969(.A1(new_n1159), .A2(new_n1160), .A3(new_n1169), .ZN(new_n1170));
  NAND3_X1  g0970(.A1(new_n1156), .A2(KEYINPUT110), .A3(new_n1170), .ZN(new_n1171));
  NAND2_X1  g0971(.A1(new_n1159), .A2(new_n1160), .ZN(new_n1172));
  INV_X1    g0972(.A(KEYINPUT110), .ZN(new_n1173));
  NAND3_X1  g0973(.A1(new_n1172), .A2(new_n1173), .A3(new_n1147), .ZN(new_n1174));
  NAND2_X1  g0974(.A1(new_n1171), .A2(new_n1174), .ZN(new_n1175));
  AOI21_X1  g0975(.A(new_n1139), .B1(new_n1175), .B2(new_n779), .ZN(new_n1176));
  OAI21_X1  g0976(.A(new_n860), .B1(new_n1145), .B2(KEYINPUT112), .ZN(new_n1177));
  AND3_X1   g0977(.A1(new_n892), .A2(KEYINPUT112), .A3(G330), .ZN(new_n1178));
  OAI21_X1  g0978(.A(new_n958), .B1(new_n1177), .B2(new_n1178), .ZN(new_n1179));
  INV_X1    g0979(.A(new_n1152), .ZN(new_n1180));
  NAND3_X1  g0980(.A1(new_n1179), .A2(new_n1169), .A3(new_n1180), .ZN(new_n1181));
  OAI211_X1 g0981(.A(G330), .B(new_n860), .C1(new_n1161), .C2(new_n1164), .ZN(new_n1182));
  NAND2_X1  g0982(.A1(new_n1182), .A2(new_n958), .ZN(new_n1183));
  NAND3_X1  g0983(.A1(new_n1183), .A2(new_n1142), .A3(new_n1146), .ZN(new_n1184));
  NAND2_X1  g0984(.A1(new_n856), .A2(new_n961), .ZN(new_n1185));
  NAND2_X1  g0985(.A1(new_n1184), .A2(new_n1185), .ZN(new_n1186));
  NAND2_X1  g0986(.A1(new_n1181), .A2(new_n1186), .ZN(new_n1187));
  NAND2_X1  g0987(.A1(new_n474), .A2(new_n1145), .ZN(new_n1188));
  NAND4_X1  g0988(.A1(new_n677), .A2(new_n954), .A3(new_n365), .A4(new_n1188), .ZN(new_n1189));
  INV_X1    g0989(.A(new_n1189), .ZN(new_n1190));
  NAND2_X1  g0990(.A1(new_n1187), .A2(new_n1190), .ZN(new_n1191));
  NAND3_X1  g0991(.A1(new_n1171), .A2(new_n1174), .A3(new_n1191), .ZN(new_n1192));
  NAND2_X1  g0992(.A1(new_n1192), .A2(new_n734), .ZN(new_n1193));
  AOI21_X1  g0993(.A(new_n1191), .B1(new_n1171), .B2(new_n1174), .ZN(new_n1194));
  OAI21_X1  g0994(.A(new_n1176), .B1(new_n1193), .B2(new_n1194), .ZN(G378));
  NAND2_X1  g0995(.A1(new_n292), .A2(new_n365), .ZN(new_n1196));
  NAND2_X1  g0996(.A1(new_n268), .A2(new_n902), .ZN(new_n1197));
  XNOR2_X1  g0997(.A(new_n1196), .B(new_n1197), .ZN(new_n1198));
  XNOR2_X1  g0998(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1199));
  XNOR2_X1  g0999(.A(new_n1198), .B(new_n1199), .ZN(new_n1200));
  AOI21_X1  g1000(.A(new_n1200), .B1(new_n946), .B2(G330), .ZN(new_n1201));
  NAND2_X1  g1001(.A1(new_n945), .A2(new_n942), .ZN(new_n1202));
  NAND3_X1  g1002(.A1(new_n892), .A2(new_n899), .A3(KEYINPUT40), .ZN(new_n1203));
  AOI211_X1 g1003(.A(KEYINPUT100), .B(new_n1203), .C1(new_n936), .C2(new_n938), .ZN(new_n1204));
  AOI21_X1  g1004(.A(new_n940), .B1(new_n939), .B2(new_n900), .ZN(new_n1205));
  OAI211_X1 g1005(.A(G330), .B(new_n1202), .C1(new_n1204), .C2(new_n1205), .ZN(new_n1206));
  INV_X1    g1006(.A(new_n1200), .ZN(new_n1207));
  NOR2_X1   g1007(.A1(new_n1206), .A2(new_n1207), .ZN(new_n1208));
  OAI21_X1  g1008(.A(new_n972), .B1(new_n1201), .B2(new_n1208), .ZN(new_n1209));
  NAND2_X1  g1009(.A1(new_n1206), .A2(new_n1207), .ZN(new_n1210));
  NAND2_X1  g1010(.A1(new_n931), .A2(new_n941), .ZN(new_n1211));
  NAND4_X1  g1011(.A1(new_n1211), .A2(G330), .A3(new_n1202), .A4(new_n1200), .ZN(new_n1212));
  INV_X1    g1012(.A(new_n972), .ZN(new_n1213));
  NAND3_X1  g1013(.A1(new_n1210), .A2(new_n1212), .A3(new_n1213), .ZN(new_n1214));
  NAND2_X1  g1014(.A1(new_n1209), .A2(new_n1214), .ZN(new_n1215));
  NAND2_X1  g1015(.A1(new_n1207), .A2(new_n795), .ZN(new_n1216));
  OAI21_X1  g1016(.A(new_n780), .B1(G50), .B2(new_n865), .ZN(new_n1217));
  OAI22_X1  g1017(.A1(new_n808), .A2(new_n1122), .B1(new_n883), .B2(new_n823), .ZN(new_n1218));
  AOI21_X1  g1018(.A(new_n1218), .B1(G137), .B2(new_n810), .ZN(new_n1219));
  AOI22_X1  g1019(.A1(new_n804), .A2(G125), .B1(new_n825), .B2(G150), .ZN(new_n1220));
  XOR2_X1   g1020(.A(new_n1220), .B(KEYINPUT117), .Z(new_n1221));
  NAND2_X1  g1021(.A1(new_n841), .A2(new_n1128), .ZN(new_n1222));
  XNOR2_X1  g1022(.A(new_n1222), .B(KEYINPUT116), .ZN(new_n1223));
  NAND3_X1  g1023(.A1(new_n1219), .A2(new_n1221), .A3(new_n1223), .ZN(new_n1224));
  OR2_X1    g1024(.A1(new_n1224), .A2(KEYINPUT59), .ZN(new_n1225));
  NAND2_X1  g1025(.A1(new_n1224), .A2(KEYINPUT59), .ZN(new_n1226));
  AOI211_X1 g1026(.A(G33), .B(G41), .C1(new_n832), .C2(G124), .ZN(new_n1227));
  OAI21_X1  g1027(.A(new_n1227), .B1(new_n815), .B2(new_n828), .ZN(new_n1228));
  XNOR2_X1  g1028(.A(new_n1228), .B(KEYINPUT118), .ZN(new_n1229));
  NAND3_X1  g1029(.A1(new_n1225), .A2(new_n1226), .A3(new_n1229), .ZN(new_n1230));
  NOR2_X1   g1030(.A1(new_n281), .A2(G41), .ZN(new_n1231));
  INV_X1    g1031(.A(new_n1231), .ZN(new_n1232));
  AOI21_X1  g1032(.A(new_n1232), .B1(G283), .B2(new_n832), .ZN(new_n1233));
  AND2_X1   g1033(.A1(new_n1233), .A2(new_n1029), .ZN(new_n1234));
  OAI221_X1 g1034(.A(new_n1234), .B1(new_n867), .B2(new_n348), .C1(new_n342), .C2(new_n808), .ZN(new_n1235));
  OAI22_X1  g1035(.A1(new_n823), .A2(new_n552), .B1(new_n820), .B2(new_n294), .ZN(new_n1236));
  OAI22_X1  g1036(.A1(new_n805), .A2(new_n636), .B1(new_n828), .B2(new_n302), .ZN(new_n1237));
  NOR3_X1   g1037(.A1(new_n1235), .A2(new_n1236), .A3(new_n1237), .ZN(new_n1238));
  NAND2_X1  g1038(.A1(new_n1238), .A2(KEYINPUT58), .ZN(new_n1239));
  OR2_X1    g1039(.A1(new_n1238), .A2(KEYINPUT58), .ZN(new_n1240));
  OAI211_X1 g1040(.A(new_n1232), .B(new_n253), .C1(G33), .C2(G41), .ZN(new_n1241));
  NAND4_X1  g1041(.A1(new_n1230), .A2(new_n1239), .A3(new_n1240), .A4(new_n1241), .ZN(new_n1242));
  AOI21_X1  g1042(.A(new_n1217), .B1(new_n1242), .B2(new_n793), .ZN(new_n1243));
  AOI22_X1  g1043(.A1(new_n1215), .A2(new_n779), .B1(new_n1216), .B2(new_n1243), .ZN(new_n1244));
  XNOR2_X1  g1044(.A(new_n1189), .B(KEYINPUT119), .ZN(new_n1245));
  INV_X1    g1045(.A(new_n1245), .ZN(new_n1246));
  INV_X1    g1046(.A(new_n1147), .ZN(new_n1247));
  AOI211_X1 g1047(.A(KEYINPUT110), .B(new_n1247), .C1(new_n1159), .C2(new_n1160), .ZN(new_n1248));
  AOI21_X1  g1048(.A(new_n1173), .B1(new_n1172), .B2(new_n1147), .ZN(new_n1249));
  AOI21_X1  g1049(.A(new_n1248), .B1(new_n1249), .B2(new_n1170), .ZN(new_n1250));
  OAI21_X1  g1050(.A(new_n1246), .B1(new_n1250), .B2(new_n1191), .ZN(new_n1251));
  AOI21_X1  g1051(.A(KEYINPUT57), .B1(new_n1251), .B2(new_n1215), .ZN(new_n1252));
  AND3_X1   g1052(.A1(new_n1210), .A2(new_n1213), .A3(new_n1212), .ZN(new_n1253));
  AOI21_X1  g1053(.A(new_n1213), .B1(new_n1210), .B2(new_n1212), .ZN(new_n1254));
  OAI21_X1  g1054(.A(KEYINPUT57), .B1(new_n1253), .B2(new_n1254), .ZN(new_n1255));
  INV_X1    g1055(.A(new_n1191), .ZN(new_n1256));
  AOI21_X1  g1056(.A(new_n1245), .B1(new_n1175), .B2(new_n1256), .ZN(new_n1257));
  OAI21_X1  g1057(.A(new_n734), .B1(new_n1255), .B2(new_n1257), .ZN(new_n1258));
  OAI21_X1  g1058(.A(new_n1244), .B1(new_n1252), .B2(new_n1258), .ZN(G375));
  NAND3_X1  g1059(.A1(new_n1181), .A2(new_n1186), .A3(new_n1189), .ZN(new_n1260));
  XNOR2_X1  g1060(.A(new_n1008), .B(KEYINPUT120), .ZN(new_n1261));
  NAND3_X1  g1061(.A1(new_n1191), .A2(new_n1260), .A3(new_n1261), .ZN(new_n1262));
  NAND2_X1  g1062(.A1(new_n958), .A2(new_n795), .ZN(new_n1263));
  OAI21_X1  g1063(.A(new_n780), .B1(G68), .B2(new_n865), .ZN(new_n1264));
  OAI22_X1  g1064(.A1(new_n823), .A2(new_n636), .B1(new_n805), .B2(new_n1104), .ZN(new_n1265));
  AOI211_X1 g1065(.A(new_n1067), .B(new_n1265), .C1(G97), .C2(new_n841), .ZN(new_n1266));
  OAI221_X1 g1066(.A(new_n328), .B1(new_n814), .B2(new_n628), .C1(new_n294), .C2(new_n828), .ZN(new_n1267));
  AOI21_X1  g1067(.A(new_n1267), .B1(new_n810), .B2(G107), .ZN(new_n1268));
  OAI211_X1 g1068(.A(new_n1266), .B(new_n1268), .C1(new_n834), .C2(new_n808), .ZN(new_n1269));
  OAI221_X1 g1069(.A(new_n281), .B1(new_n814), .B2(new_n1122), .C1(new_n302), .C2(new_n828), .ZN(new_n1270));
  AOI21_X1  g1070(.A(new_n1270), .B1(new_n810), .B2(G150), .ZN(new_n1271));
  AOI22_X1  g1071(.A1(new_n804), .A2(G132), .B1(new_n841), .B2(G159), .ZN(new_n1272));
  AOI22_X1  g1072(.A1(new_n822), .A2(new_n1128), .B1(new_n825), .B2(G50), .ZN(new_n1273));
  NAND2_X1  g1073(.A1(new_n807), .A2(G137), .ZN(new_n1274));
  NAND4_X1  g1074(.A1(new_n1271), .A2(new_n1272), .A3(new_n1273), .A4(new_n1274), .ZN(new_n1275));
  NAND2_X1  g1075(.A1(new_n1269), .A2(new_n1275), .ZN(new_n1276));
  OR2_X1    g1076(.A1(new_n1276), .A2(KEYINPUT121), .ZN(new_n1277));
  AOI21_X1  g1077(.A(new_n794), .B1(new_n1276), .B2(KEYINPUT121), .ZN(new_n1278));
  AOI21_X1  g1078(.A(new_n1264), .B1(new_n1277), .B2(new_n1278), .ZN(new_n1279));
  AOI22_X1  g1079(.A1(new_n1187), .A2(new_n779), .B1(new_n1263), .B2(new_n1279), .ZN(new_n1280));
  NAND2_X1  g1080(.A1(new_n1262), .A2(new_n1280), .ZN(new_n1281));
  XNOR2_X1  g1081(.A(new_n1281), .B(KEYINPUT122), .ZN(G381));
  INV_X1    g1082(.A(G390), .ZN(new_n1283));
  INV_X1    g1083(.A(G384), .ZN(new_n1284));
  NOR2_X1   g1084(.A1(G393), .A2(G396), .ZN(new_n1285));
  NAND3_X1  g1085(.A1(new_n1283), .A2(new_n1284), .A3(new_n1285), .ZN(new_n1286));
  NOR3_X1   g1086(.A1(new_n1286), .A2(G381), .A3(G387), .ZN(new_n1287));
  INV_X1    g1087(.A(G378), .ZN(new_n1288));
  NAND2_X1  g1088(.A1(new_n1216), .A2(new_n1243), .ZN(new_n1289));
  NOR2_X1   g1089(.A1(new_n1253), .A2(new_n1254), .ZN(new_n1290));
  OAI21_X1  g1090(.A(new_n1289), .B1(new_n1290), .B2(new_n778), .ZN(new_n1291));
  INV_X1    g1091(.A(KEYINPUT57), .ZN(new_n1292));
  AOI21_X1  g1092(.A(new_n1292), .B1(new_n1209), .B2(new_n1214), .ZN(new_n1293));
  AOI21_X1  g1093(.A(new_n1055), .B1(new_n1251), .B2(new_n1293), .ZN(new_n1294));
  OAI21_X1  g1094(.A(new_n1292), .B1(new_n1257), .B2(new_n1290), .ZN(new_n1295));
  AOI21_X1  g1095(.A(new_n1291), .B1(new_n1294), .B2(new_n1295), .ZN(new_n1296));
  NAND3_X1  g1096(.A1(new_n1287), .A2(new_n1288), .A3(new_n1296), .ZN(G407));
  NAND2_X1  g1097(.A1(new_n717), .A2(G213), .ZN(new_n1298));
  INV_X1    g1098(.A(new_n1298), .ZN(new_n1299));
  NAND3_X1  g1099(.A1(new_n1296), .A2(new_n1288), .A3(new_n1299), .ZN(new_n1300));
  NAND3_X1  g1100(.A1(G407), .A2(G213), .A3(new_n1300), .ZN(G409));
  OAI211_X1 g1101(.A(G378), .B(new_n1244), .C1(new_n1252), .C2(new_n1258), .ZN(new_n1302));
  OAI211_X1 g1102(.A(new_n1215), .B(new_n1261), .C1(new_n1194), .C2(new_n1245), .ZN(new_n1303));
  NAND2_X1  g1103(.A1(new_n1303), .A2(new_n1244), .ZN(new_n1304));
  NAND2_X1  g1104(.A1(new_n1304), .A2(new_n1288), .ZN(new_n1305));
  NAND2_X1  g1105(.A1(new_n1302), .A2(new_n1305), .ZN(new_n1306));
  NAND2_X1  g1106(.A1(new_n1306), .A2(new_n1298), .ZN(new_n1307));
  INV_X1    g1107(.A(KEYINPUT126), .ZN(new_n1308));
  INV_X1    g1108(.A(G2897), .ZN(new_n1309));
  NOR2_X1   g1109(.A1(new_n1298), .A2(new_n1309), .ZN(new_n1310));
  INV_X1    g1110(.A(new_n1310), .ZN(new_n1311));
  NAND4_X1  g1111(.A1(new_n1181), .A2(new_n1186), .A3(new_n1189), .A4(KEYINPUT60), .ZN(new_n1312));
  INV_X1    g1112(.A(KEYINPUT123), .ZN(new_n1313));
  NAND2_X1  g1113(.A1(new_n1312), .A2(new_n1313), .ZN(new_n1314));
  AOI21_X1  g1114(.A(new_n1055), .B1(new_n1187), .B2(new_n1190), .ZN(new_n1315));
  AOI21_X1  g1115(.A(new_n1152), .B1(new_n1166), .B2(new_n1168), .ZN(new_n1316));
  AOI22_X1  g1116(.A1(new_n1316), .A2(new_n1179), .B1(new_n1184), .B2(new_n1185), .ZN(new_n1317));
  NAND4_X1  g1117(.A1(new_n1317), .A2(KEYINPUT123), .A3(KEYINPUT60), .A4(new_n1189), .ZN(new_n1318));
  INV_X1    g1118(.A(KEYINPUT60), .ZN(new_n1319));
  NAND2_X1  g1119(.A1(new_n1260), .A2(new_n1319), .ZN(new_n1320));
  NAND4_X1  g1120(.A1(new_n1314), .A2(new_n1315), .A3(new_n1318), .A4(new_n1320), .ZN(new_n1321));
  AND3_X1   g1121(.A1(new_n1321), .A2(G384), .A3(new_n1280), .ZN(new_n1322));
  AOI21_X1  g1122(.A(G384), .B1(new_n1321), .B2(new_n1280), .ZN(new_n1323));
  INV_X1    g1123(.A(KEYINPUT124), .ZN(new_n1324));
  NOR3_X1   g1124(.A1(new_n1322), .A2(new_n1323), .A3(new_n1324), .ZN(new_n1325));
  NAND2_X1  g1125(.A1(new_n1321), .A2(new_n1280), .ZN(new_n1326));
  NAND2_X1  g1126(.A1(new_n1326), .A2(new_n1284), .ZN(new_n1327));
  NAND3_X1  g1127(.A1(new_n1321), .A2(G384), .A3(new_n1280), .ZN(new_n1328));
  AOI21_X1  g1128(.A(KEYINPUT124), .B1(new_n1327), .B2(new_n1328), .ZN(new_n1329));
  OAI21_X1  g1129(.A(new_n1311), .B1(new_n1325), .B2(new_n1329), .ZN(new_n1330));
  AOI21_X1  g1130(.A(new_n1311), .B1(new_n1327), .B2(new_n1328), .ZN(new_n1331));
  INV_X1    g1131(.A(new_n1331), .ZN(new_n1332));
  AOI21_X1  g1132(.A(new_n1308), .B1(new_n1330), .B2(new_n1332), .ZN(new_n1333));
  OAI21_X1  g1133(.A(new_n1324), .B1(new_n1322), .B2(new_n1323), .ZN(new_n1334));
  NAND3_X1  g1134(.A1(new_n1327), .A2(KEYINPUT124), .A3(new_n1328), .ZN(new_n1335));
  AOI21_X1  g1135(.A(new_n1310), .B1(new_n1334), .B2(new_n1335), .ZN(new_n1336));
  NOR3_X1   g1136(.A1(new_n1336), .A2(KEYINPUT126), .A3(new_n1331), .ZN(new_n1337));
  OAI21_X1  g1137(.A(new_n1307), .B1(new_n1333), .B2(new_n1337), .ZN(new_n1338));
  NAND2_X1  g1138(.A1(new_n1334), .A2(new_n1335), .ZN(new_n1339));
  NAND3_X1  g1139(.A1(new_n1306), .A2(new_n1298), .A3(new_n1339), .ZN(new_n1340));
  NAND2_X1  g1140(.A1(new_n1340), .A2(KEYINPUT62), .ZN(new_n1341));
  INV_X1    g1141(.A(KEYINPUT61), .ZN(new_n1342));
  AOI21_X1  g1142(.A(new_n1299), .B1(new_n1302), .B2(new_n1305), .ZN(new_n1343));
  INV_X1    g1143(.A(KEYINPUT62), .ZN(new_n1344));
  NAND3_X1  g1144(.A1(new_n1343), .A2(new_n1344), .A3(new_n1339), .ZN(new_n1345));
  NAND4_X1  g1145(.A1(new_n1338), .A2(new_n1341), .A3(new_n1342), .A4(new_n1345), .ZN(new_n1346));
  NAND3_X1  g1146(.A1(new_n1025), .A2(new_n1053), .A3(G390), .ZN(new_n1347));
  INV_X1    g1147(.A(new_n1347), .ZN(new_n1348));
  AOI21_X1  g1148(.A(G390), .B1(new_n1025), .B2(new_n1053), .ZN(new_n1349));
  AOI21_X1  g1149(.A(new_n848), .B1(new_n1057), .B2(new_n1086), .ZN(new_n1350));
  OAI22_X1  g1150(.A1(new_n1348), .A2(new_n1349), .B1(new_n1285), .B2(new_n1350), .ZN(new_n1351));
  INV_X1    g1151(.A(new_n1349), .ZN(new_n1352));
  NOR2_X1   g1152(.A1(new_n1285), .A2(new_n1350), .ZN(new_n1353));
  NAND3_X1  g1153(.A1(new_n1352), .A2(new_n1353), .A3(new_n1347), .ZN(new_n1354));
  NAND2_X1  g1154(.A1(new_n1351), .A2(new_n1354), .ZN(new_n1355));
  NAND2_X1  g1155(.A1(new_n1346), .A2(new_n1355), .ZN(new_n1356));
  AOI21_X1  g1156(.A(G378), .B1(new_n1244), .B2(new_n1303), .ZN(new_n1357));
  AOI21_X1  g1157(.A(new_n1357), .B1(new_n1296), .B2(G378), .ZN(new_n1358));
  OAI21_X1  g1158(.A(KEYINPUT125), .B1(new_n1358), .B2(new_n1299), .ZN(new_n1359));
  INV_X1    g1159(.A(KEYINPUT125), .ZN(new_n1360));
  NAND2_X1  g1160(.A1(new_n1343), .A2(new_n1360), .ZN(new_n1361));
  NAND2_X1  g1161(.A1(new_n1359), .A2(new_n1361), .ZN(new_n1362));
  INV_X1    g1162(.A(KEYINPUT127), .ZN(new_n1363));
  OAI21_X1  g1163(.A(new_n1363), .B1(new_n1333), .B2(new_n1337), .ZN(new_n1364));
  NAND3_X1  g1164(.A1(new_n1330), .A2(new_n1332), .A3(new_n1308), .ZN(new_n1365));
  OAI21_X1  g1165(.A(KEYINPUT126), .B1(new_n1336), .B2(new_n1331), .ZN(new_n1366));
  NAND3_X1  g1166(.A1(new_n1365), .A2(new_n1366), .A3(KEYINPUT127), .ZN(new_n1367));
  NAND3_X1  g1167(.A1(new_n1362), .A2(new_n1364), .A3(new_n1367), .ZN(new_n1368));
  NAND4_X1  g1168(.A1(new_n1306), .A2(KEYINPUT63), .A3(new_n1298), .A4(new_n1339), .ZN(new_n1369));
  AND3_X1   g1169(.A1(new_n1351), .A2(new_n1354), .A3(new_n1342), .ZN(new_n1370));
  NAND2_X1  g1170(.A1(new_n1369), .A2(new_n1370), .ZN(new_n1371));
  AOI21_X1  g1171(.A(KEYINPUT63), .B1(new_n1343), .B2(new_n1339), .ZN(new_n1372));
  NOR2_X1   g1172(.A1(new_n1371), .A2(new_n1372), .ZN(new_n1373));
  NAND2_X1  g1173(.A1(new_n1368), .A2(new_n1373), .ZN(new_n1374));
  NAND2_X1  g1174(.A1(new_n1356), .A2(new_n1374), .ZN(G405));
  NOR2_X1   g1175(.A1(new_n1296), .A2(G378), .ZN(new_n1376));
  INV_X1    g1176(.A(new_n1302), .ZN(new_n1377));
  OAI21_X1  g1177(.A(new_n1339), .B1(new_n1376), .B2(new_n1377), .ZN(new_n1378));
  NOR2_X1   g1178(.A1(new_n1322), .A2(new_n1323), .ZN(new_n1379));
  OR2_X1    g1179(.A1(new_n1376), .A2(new_n1377), .ZN(new_n1380));
  OAI21_X1  g1180(.A(new_n1378), .B1(new_n1379), .B2(new_n1380), .ZN(new_n1381));
  XNOR2_X1  g1181(.A(new_n1381), .B(new_n1355), .ZN(G402));
endmodule


