//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 1 1 0 1 1 1 1 0 1 0 1 1 0 1 1 1 0 0 0 0 1 0 0 1 0 1 0 0 0 0 1 0 0 0 1 1 1 0 1 1 0 0 1 1 1 1 1 1 0 1 0 0 1 0 1 0 0 0 1 0 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:34:19 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n442, new_n446, new_n448, new_n449, new_n453, new_n454, new_n455,
    new_n456, new_n457, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n496,
    new_n497, new_n498, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n516, new_n517, new_n518,
    new_n519, new_n520, new_n521, new_n523, new_n524, new_n525, new_n526,
    new_n527, new_n528, new_n529, new_n530, new_n531, new_n532, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n558, new_n559, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n576, new_n577, new_n578, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n589, new_n590, new_n591,
    new_n592, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n620, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n630, new_n631, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1144, new_n1145;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  XOR2_X1   g003(.A(KEYINPUT64), .B(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  AND2_X1   g016(.A1(G2072), .A2(G2078), .ZN(new_n442));
  NAND3_X1  g017(.A1(new_n442), .A2(G2084), .A3(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  NAND2_X1  g020(.A1(G94), .A2(G452), .ZN(new_n446));
  XNOR2_X1  g021(.A(new_n446), .B(KEYINPUT65), .ZN(G173));
  XNOR2_X1  g022(.A(KEYINPUT66), .B(KEYINPUT1), .ZN(new_n448));
  AND2_X1   g023(.A1(G7), .A2(G661), .ZN(new_n449));
  XNOR2_X1  g024(.A(new_n448), .B(new_n449), .ZN(G223));
  NAND2_X1  g025(.A1(new_n449), .A2(G567), .ZN(G234));
  NAND2_X1  g026(.A1(new_n449), .A2(G2106), .ZN(G217));
  NOR4_X1   g027(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n453));
  XNOR2_X1  g028(.A(new_n453), .B(KEYINPUT2), .ZN(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(new_n455));
  NOR4_X1   g030(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n456));
  INV_X1    g031(.A(new_n456), .ZN(new_n457));
  NOR2_X1   g032(.A1(new_n455), .A2(new_n457), .ZN(G325));
  INV_X1    g033(.A(G325), .ZN(G261));
  AOI22_X1  g034(.A1(new_n455), .A2(G2106), .B1(G567), .B2(new_n457), .ZN(G319));
  XNOR2_X1  g035(.A(KEYINPUT3), .B(G2104), .ZN(new_n461));
  INV_X1    g036(.A(G2105), .ZN(new_n462));
  NAND2_X1  g037(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  INV_X1    g038(.A(G137), .ZN(new_n464));
  INV_X1    g039(.A(G101), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n462), .A2(G2104), .ZN(new_n466));
  OAI22_X1  g041(.A1(new_n463), .A2(new_n464), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n461), .A2(G125), .ZN(new_n468));
  NAND2_X1  g043(.A1(G113), .A2(G2104), .ZN(new_n469));
  AOI21_X1  g044(.A(new_n462), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  NOR2_X1   g045(.A1(new_n467), .A2(new_n470), .ZN(new_n471));
  XNOR2_X1  g046(.A(new_n471), .B(KEYINPUT67), .ZN(G160));
  OR2_X1    g047(.A1(G100), .A2(G2105), .ZN(new_n473));
  OAI211_X1 g048(.A(new_n473), .B(G2104), .C1(G112), .C2(new_n462), .ZN(new_n474));
  XOR2_X1   g049(.A(new_n474), .B(KEYINPUT68), .Z(new_n475));
  AND2_X1   g050(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n476));
  NOR2_X1   g051(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n477));
  NOR2_X1   g052(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  NOR2_X1   g053(.A1(new_n478), .A2(G2105), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n479), .A2(G136), .ZN(new_n480));
  NOR2_X1   g055(.A1(new_n478), .A2(new_n462), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n481), .A2(G124), .ZN(new_n482));
  NAND3_X1  g057(.A1(new_n475), .A2(new_n480), .A3(new_n482), .ZN(new_n483));
  XOR2_X1   g058(.A(new_n483), .B(KEYINPUT69), .Z(G162));
  OAI211_X1 g059(.A(G138), .B(new_n462), .C1(new_n476), .C2(new_n477), .ZN(new_n485));
  INV_X1    g060(.A(KEYINPUT4), .ZN(new_n486));
  NAND2_X1  g061(.A1(new_n485), .A2(new_n486), .ZN(new_n487));
  OAI21_X1  g062(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n488));
  INV_X1    g063(.A(new_n488), .ZN(new_n489));
  XNOR2_X1  g064(.A(KEYINPUT70), .B(G114), .ZN(new_n490));
  OAI21_X1  g065(.A(new_n489), .B1(new_n490), .B2(new_n462), .ZN(new_n491));
  NAND4_X1  g066(.A1(new_n461), .A2(KEYINPUT4), .A3(G138), .A4(new_n462), .ZN(new_n492));
  NAND3_X1  g067(.A1(new_n461), .A2(G126), .A3(G2105), .ZN(new_n493));
  NAND4_X1  g068(.A1(new_n487), .A2(new_n491), .A3(new_n492), .A4(new_n493), .ZN(new_n494));
  INV_X1    g069(.A(new_n494), .ZN(G164));
  NAND2_X1  g070(.A1(KEYINPUT71), .A2(KEYINPUT5), .ZN(new_n496));
  INV_X1    g071(.A(G543), .ZN(new_n497));
  NAND2_X1  g072(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  NAND3_X1  g073(.A1(KEYINPUT71), .A2(KEYINPUT5), .A3(G543), .ZN(new_n499));
  NAND2_X1  g074(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  AOI22_X1  g075(.A1(new_n500), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n501));
  INV_X1    g076(.A(G651), .ZN(new_n502));
  NOR2_X1   g077(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  INV_X1    g078(.A(new_n503), .ZN(new_n504));
  OR2_X1    g079(.A1(KEYINPUT6), .A2(G651), .ZN(new_n505));
  NAND2_X1  g080(.A1(KEYINPUT6), .A2(G651), .ZN(new_n506));
  AOI22_X1  g081(.A1(new_n498), .A2(new_n499), .B1(new_n505), .B2(new_n506), .ZN(new_n507));
  NAND2_X1  g082(.A1(new_n507), .A2(G88), .ZN(new_n508));
  AOI21_X1  g083(.A(new_n497), .B1(new_n505), .B2(new_n506), .ZN(new_n509));
  NAND2_X1  g084(.A1(new_n509), .A2(G50), .ZN(new_n510));
  NAND3_X1  g085(.A1(new_n508), .A2(KEYINPUT72), .A3(new_n510), .ZN(new_n511));
  INV_X1    g086(.A(new_n511), .ZN(new_n512));
  AOI21_X1  g087(.A(KEYINPUT72), .B1(new_n508), .B2(new_n510), .ZN(new_n513));
  OAI21_X1  g088(.A(new_n504), .B1(new_n512), .B2(new_n513), .ZN(new_n514));
  INV_X1    g089(.A(new_n514), .ZN(G166));
  NAND2_X1  g090(.A1(new_n509), .A2(G51), .ZN(new_n516));
  NAND3_X1  g091(.A1(new_n500), .A2(G63), .A3(G651), .ZN(new_n517));
  NAND3_X1  g092(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n518));
  XNOR2_X1  g093(.A(new_n518), .B(KEYINPUT7), .ZN(new_n519));
  NAND3_X1  g094(.A1(new_n516), .A2(new_n517), .A3(new_n519), .ZN(new_n520));
  AND2_X1   g095(.A1(new_n507), .A2(G89), .ZN(new_n521));
  NOR2_X1   g096(.A1(new_n520), .A2(new_n521), .ZN(G168));
  AOI22_X1  g097(.A1(new_n507), .A2(G90), .B1(new_n509), .B2(G52), .ZN(new_n523));
  XNOR2_X1  g098(.A(new_n523), .B(KEYINPUT74), .ZN(new_n524));
  NAND2_X1  g099(.A1(G77), .A2(G543), .ZN(new_n525));
  AND3_X1   g100(.A1(KEYINPUT71), .A2(KEYINPUT5), .A3(G543), .ZN(new_n526));
  AOI21_X1  g101(.A(G543), .B1(KEYINPUT71), .B2(KEYINPUT5), .ZN(new_n527));
  NOR2_X1   g102(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  INV_X1    g103(.A(G64), .ZN(new_n529));
  OAI21_X1  g104(.A(new_n525), .B1(new_n528), .B2(new_n529), .ZN(new_n530));
  AOI21_X1  g105(.A(new_n502), .B1(new_n530), .B2(KEYINPUT73), .ZN(new_n531));
  OAI21_X1  g106(.A(new_n531), .B1(KEYINPUT73), .B2(new_n530), .ZN(new_n532));
  AND2_X1   g107(.A1(new_n524), .A2(new_n532), .ZN(G171));
  INV_X1    g108(.A(G56), .ZN(new_n534));
  AOI21_X1  g109(.A(new_n534), .B1(new_n498), .B2(new_n499), .ZN(new_n535));
  NAND2_X1  g110(.A1(G68), .A2(G543), .ZN(new_n536));
  INV_X1    g111(.A(new_n536), .ZN(new_n537));
  OAI21_X1  g112(.A(KEYINPUT75), .B1(new_n535), .B2(new_n537), .ZN(new_n538));
  OAI21_X1  g113(.A(G56), .B1(new_n526), .B2(new_n527), .ZN(new_n539));
  INV_X1    g114(.A(KEYINPUT75), .ZN(new_n540));
  NAND3_X1  g115(.A1(new_n539), .A2(new_n540), .A3(new_n536), .ZN(new_n541));
  NAND3_X1  g116(.A1(new_n538), .A2(G651), .A3(new_n541), .ZN(new_n542));
  INV_X1    g117(.A(KEYINPUT76), .ZN(new_n543));
  NAND2_X1  g118(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  NAND4_X1  g119(.A1(new_n538), .A2(KEYINPUT76), .A3(G651), .A4(new_n541), .ZN(new_n545));
  XNOR2_X1  g120(.A(KEYINPUT77), .B(G43), .ZN(new_n546));
  NAND2_X1  g121(.A1(new_n509), .A2(new_n546), .ZN(new_n547));
  INV_X1    g122(.A(G81), .ZN(new_n548));
  INV_X1    g123(.A(new_n506), .ZN(new_n549));
  NOR2_X1   g124(.A1(KEYINPUT6), .A2(G651), .ZN(new_n550));
  OAI22_X1  g125(.A1(new_n526), .A2(new_n527), .B1(new_n549), .B2(new_n550), .ZN(new_n551));
  OAI21_X1  g126(.A(new_n547), .B1(new_n548), .B2(new_n551), .ZN(new_n552));
  INV_X1    g127(.A(new_n552), .ZN(new_n553));
  NAND3_X1  g128(.A1(new_n544), .A2(new_n545), .A3(new_n553), .ZN(new_n554));
  INV_X1    g129(.A(new_n554), .ZN(new_n555));
  NAND2_X1  g130(.A1(new_n555), .A2(G860), .ZN(G153));
  NAND4_X1  g131(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g132(.A1(G1), .A2(G3), .ZN(new_n558));
  XNOR2_X1  g133(.A(new_n558), .B(KEYINPUT8), .ZN(new_n559));
  NAND4_X1  g134(.A1(G319), .A2(G483), .A3(G661), .A4(new_n559), .ZN(G188));
  OAI211_X1 g135(.A(G53), .B(G543), .C1(new_n549), .C2(new_n550), .ZN(new_n561));
  NAND2_X1  g136(.A1(new_n561), .A2(KEYINPUT9), .ZN(new_n562));
  NAND2_X1  g137(.A1(new_n505), .A2(new_n506), .ZN(new_n563));
  INV_X1    g138(.A(KEYINPUT9), .ZN(new_n564));
  NAND4_X1  g139(.A1(new_n563), .A2(new_n564), .A3(G53), .A4(G543), .ZN(new_n565));
  AOI22_X1  g140(.A1(new_n562), .A2(new_n565), .B1(new_n507), .B2(G91), .ZN(new_n566));
  OAI21_X1  g141(.A(G65), .B1(new_n526), .B2(new_n527), .ZN(new_n567));
  NAND2_X1  g142(.A1(G78), .A2(G543), .ZN(new_n568));
  NAND2_X1  g143(.A1(new_n567), .A2(new_n568), .ZN(new_n569));
  AOI21_X1  g144(.A(KEYINPUT78), .B1(new_n569), .B2(G651), .ZN(new_n570));
  INV_X1    g145(.A(KEYINPUT78), .ZN(new_n571));
  AOI211_X1 g146(.A(new_n571), .B(new_n502), .C1(new_n567), .C2(new_n568), .ZN(new_n572));
  OAI21_X1  g147(.A(new_n566), .B1(new_n570), .B2(new_n572), .ZN(G299));
  NAND2_X1  g148(.A1(new_n524), .A2(new_n532), .ZN(G301));
  INV_X1    g149(.A(G168), .ZN(G286));
  INV_X1    g150(.A(KEYINPUT79), .ZN(new_n576));
  NAND2_X1  g151(.A1(new_n514), .A2(new_n576), .ZN(new_n577));
  OAI211_X1 g152(.A(KEYINPUT79), .B(new_n504), .C1(new_n512), .C2(new_n513), .ZN(new_n578));
  AND2_X1   g153(.A1(new_n577), .A2(new_n578), .ZN(G303));
  NAND3_X1  g154(.A1(new_n563), .A2(G49), .A3(G543), .ZN(new_n580));
  NAND2_X1  g155(.A1(new_n580), .A2(KEYINPUT80), .ZN(new_n581));
  INV_X1    g156(.A(KEYINPUT80), .ZN(new_n582));
  NAND3_X1  g157(.A1(new_n509), .A2(new_n582), .A3(G49), .ZN(new_n583));
  NAND2_X1  g158(.A1(new_n581), .A2(new_n583), .ZN(new_n584));
  INV_X1    g159(.A(G74), .ZN(new_n585));
  NAND2_X1  g160(.A1(new_n528), .A2(new_n585), .ZN(new_n586));
  AOI22_X1  g161(.A1(new_n586), .A2(G651), .B1(new_n507), .B2(G87), .ZN(new_n587));
  NAND2_X1  g162(.A1(new_n584), .A2(new_n587), .ZN(G288));
  AOI22_X1  g163(.A1(new_n500), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n589));
  OR2_X1    g164(.A1(new_n589), .A2(new_n502), .ZN(new_n590));
  NAND2_X1  g165(.A1(new_n507), .A2(G86), .ZN(new_n591));
  NAND2_X1  g166(.A1(new_n509), .A2(G48), .ZN(new_n592));
  NAND3_X1  g167(.A1(new_n590), .A2(new_n591), .A3(new_n592), .ZN(G305));
  AOI22_X1  g168(.A1(new_n500), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n594));
  NOR2_X1   g169(.A1(new_n594), .A2(new_n502), .ZN(new_n595));
  NAND2_X1  g170(.A1(new_n509), .A2(G47), .ZN(new_n596));
  INV_X1    g171(.A(G85), .ZN(new_n597));
  OAI21_X1  g172(.A(new_n596), .B1(new_n597), .B2(new_n551), .ZN(new_n598));
  NOR2_X1   g173(.A1(new_n595), .A2(new_n598), .ZN(new_n599));
  INV_X1    g174(.A(new_n599), .ZN(G290));
  XNOR2_X1  g175(.A(KEYINPUT83), .B(G66), .ZN(new_n601));
  NOR2_X1   g176(.A1(new_n528), .A2(new_n601), .ZN(new_n602));
  NAND2_X1  g177(.A1(G79), .A2(G543), .ZN(new_n603));
  NAND2_X1  g178(.A1(new_n603), .A2(KEYINPUT82), .ZN(new_n604));
  INV_X1    g179(.A(KEYINPUT82), .ZN(new_n605));
  NAND3_X1  g180(.A1(new_n605), .A2(G79), .A3(G543), .ZN(new_n606));
  NAND2_X1  g181(.A1(new_n604), .A2(new_n606), .ZN(new_n607));
  OAI21_X1  g182(.A(G651), .B1(new_n602), .B2(new_n607), .ZN(new_n608));
  NAND2_X1  g183(.A1(new_n509), .A2(G54), .ZN(new_n609));
  XNOR2_X1  g184(.A(KEYINPUT81), .B(KEYINPUT10), .ZN(new_n610));
  INV_X1    g185(.A(new_n610), .ZN(new_n611));
  NAND3_X1  g186(.A1(new_n507), .A2(G92), .A3(new_n611), .ZN(new_n612));
  INV_X1    g187(.A(G92), .ZN(new_n613));
  OAI21_X1  g188(.A(new_n610), .B1(new_n551), .B2(new_n613), .ZN(new_n614));
  NAND4_X1  g189(.A1(new_n608), .A2(new_n609), .A3(new_n612), .A4(new_n614), .ZN(new_n615));
  INV_X1    g190(.A(G868), .ZN(new_n616));
  NAND2_X1  g191(.A1(new_n615), .A2(new_n616), .ZN(new_n617));
  OAI21_X1  g192(.A(new_n617), .B1(G171), .B2(new_n616), .ZN(G284));
  OAI21_X1  g193(.A(new_n617), .B1(G171), .B2(new_n616), .ZN(G321));
  NAND2_X1  g194(.A1(G299), .A2(new_n616), .ZN(new_n620));
  OAI21_X1  g195(.A(new_n620), .B1(new_n616), .B2(G168), .ZN(G297));
  OAI21_X1  g196(.A(new_n620), .B1(new_n616), .B2(G168), .ZN(G280));
  INV_X1    g197(.A(new_n601), .ZN(new_n623));
  AOI21_X1  g198(.A(new_n607), .B1(new_n623), .B2(new_n500), .ZN(new_n624));
  OAI21_X1  g199(.A(new_n609), .B1(new_n624), .B2(new_n502), .ZN(new_n625));
  NAND2_X1  g200(.A1(new_n614), .A2(new_n612), .ZN(new_n626));
  NOR2_X1   g201(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  INV_X1    g202(.A(G559), .ZN(new_n628));
  OAI21_X1  g203(.A(new_n627), .B1(new_n628), .B2(G860), .ZN(G148));
  NAND2_X1  g204(.A1(new_n554), .A2(new_n616), .ZN(new_n630));
  NOR2_X1   g205(.A1(new_n615), .A2(G559), .ZN(new_n631));
  OAI21_X1  g206(.A(new_n630), .B1(new_n631), .B2(new_n616), .ZN(G323));
  XNOR2_X1  g207(.A(G323), .B(KEYINPUT11), .ZN(G282));
  INV_X1    g208(.A(new_n466), .ZN(new_n634));
  NAND2_X1  g209(.A1(new_n461), .A2(new_n634), .ZN(new_n635));
  XOR2_X1   g210(.A(new_n635), .B(KEYINPUT12), .Z(new_n636));
  INV_X1    g211(.A(new_n636), .ZN(new_n637));
  INV_X1    g212(.A(KEYINPUT13), .ZN(new_n638));
  AOI22_X1  g213(.A1(new_n637), .A2(new_n638), .B1(KEYINPUT84), .B2(G2100), .ZN(new_n639));
  OAI21_X1  g214(.A(new_n639), .B1(new_n638), .B2(new_n637), .ZN(new_n640));
  NOR2_X1   g215(.A1(KEYINPUT84), .A2(G2100), .ZN(new_n641));
  XNOR2_X1  g216(.A(new_n640), .B(new_n641), .ZN(new_n642));
  NAND2_X1  g217(.A1(new_n479), .A2(G135), .ZN(new_n643));
  NAND2_X1  g218(.A1(new_n481), .A2(G123), .ZN(new_n644));
  NOR2_X1   g219(.A1(new_n462), .A2(G111), .ZN(new_n645));
  OAI21_X1  g220(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n646));
  OAI211_X1 g221(.A(new_n643), .B(new_n644), .C1(new_n645), .C2(new_n646), .ZN(new_n647));
  XNOR2_X1  g222(.A(new_n647), .B(KEYINPUT85), .ZN(new_n648));
  XNOR2_X1  g223(.A(new_n648), .B(G2096), .ZN(new_n649));
  NAND2_X1  g224(.A1(new_n642), .A2(new_n649), .ZN(G156));
  XNOR2_X1  g225(.A(G2427), .B(G2438), .ZN(new_n651));
  XNOR2_X1  g226(.A(new_n651), .B(G2430), .ZN(new_n652));
  XNOR2_X1  g227(.A(KEYINPUT15), .B(G2435), .ZN(new_n653));
  OR2_X1    g228(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  NAND2_X1  g229(.A1(new_n652), .A2(new_n653), .ZN(new_n655));
  NAND3_X1  g230(.A1(new_n654), .A2(KEYINPUT14), .A3(new_n655), .ZN(new_n656));
  XNOR2_X1  g231(.A(new_n656), .B(KEYINPUT86), .ZN(new_n657));
  XNOR2_X1  g232(.A(G2451), .B(G2454), .ZN(new_n658));
  XNOR2_X1  g233(.A(new_n658), .B(KEYINPUT16), .ZN(new_n659));
  XNOR2_X1  g234(.A(G2443), .B(G2446), .ZN(new_n660));
  XNOR2_X1  g235(.A(new_n659), .B(new_n660), .ZN(new_n661));
  XNOR2_X1  g236(.A(new_n657), .B(new_n661), .ZN(new_n662));
  XNOR2_X1  g237(.A(G1341), .B(G1348), .ZN(new_n663));
  OR2_X1    g238(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  NAND2_X1  g239(.A1(new_n662), .A2(new_n663), .ZN(new_n665));
  NAND3_X1  g240(.A1(new_n664), .A2(G14), .A3(new_n665), .ZN(new_n666));
  XNOR2_X1  g241(.A(new_n666), .B(KEYINPUT87), .ZN(G401));
  XNOR2_X1  g242(.A(G2084), .B(G2090), .ZN(new_n668));
  XNOR2_X1  g243(.A(new_n668), .B(KEYINPUT88), .ZN(new_n669));
  XNOR2_X1  g244(.A(G2067), .B(G2678), .ZN(new_n670));
  NAND2_X1  g245(.A1(new_n669), .A2(new_n670), .ZN(new_n671));
  AND2_X1   g246(.A1(new_n671), .A2(KEYINPUT17), .ZN(new_n672));
  OR2_X1    g247(.A1(new_n669), .A2(new_n670), .ZN(new_n673));
  AOI21_X1  g248(.A(KEYINPUT18), .B1(new_n672), .B2(new_n673), .ZN(new_n674));
  XNOR2_X1  g249(.A(KEYINPUT89), .B(G2100), .ZN(new_n675));
  XNOR2_X1  g250(.A(new_n674), .B(new_n675), .ZN(new_n676));
  NOR2_X1   g251(.A1(G2072), .A2(G2078), .ZN(new_n677));
  NOR2_X1   g252(.A1(new_n442), .A2(new_n677), .ZN(new_n678));
  AOI21_X1  g253(.A(new_n678), .B1(new_n671), .B2(KEYINPUT18), .ZN(new_n679));
  XOR2_X1   g254(.A(new_n679), .B(G2096), .Z(new_n680));
  XNOR2_X1  g255(.A(new_n676), .B(new_n680), .ZN(G227));
  XNOR2_X1  g256(.A(G1956), .B(G2474), .ZN(new_n682));
  XNOR2_X1  g257(.A(new_n682), .B(KEYINPUT90), .ZN(new_n683));
  XNOR2_X1  g258(.A(G1961), .B(G1966), .ZN(new_n684));
  INV_X1    g259(.A(new_n684), .ZN(new_n685));
  NAND2_X1  g260(.A1(new_n683), .A2(new_n685), .ZN(new_n686));
  XNOR2_X1  g261(.A(G1971), .B(G1976), .ZN(new_n687));
  XNOR2_X1  g262(.A(new_n687), .B(KEYINPUT19), .ZN(new_n688));
  NOR2_X1   g263(.A1(new_n686), .A2(new_n688), .ZN(new_n689));
  XOR2_X1   g264(.A(new_n689), .B(KEYINPUT20), .Z(new_n690));
  NOR2_X1   g265(.A1(new_n683), .A2(new_n685), .ZN(new_n691));
  INV_X1    g266(.A(new_n691), .ZN(new_n692));
  NAND3_X1  g267(.A1(new_n692), .A2(new_n688), .A3(new_n686), .ZN(new_n693));
  OAI211_X1 g268(.A(new_n690), .B(new_n693), .C1(new_n688), .C2(new_n692), .ZN(new_n694));
  XNOR2_X1  g269(.A(new_n694), .B(KEYINPUT92), .ZN(new_n695));
  XOR2_X1   g270(.A(G1981), .B(G1986), .Z(new_n696));
  XNOR2_X1  g271(.A(G1991), .B(G1996), .ZN(new_n697));
  XNOR2_X1  g272(.A(new_n696), .B(new_n697), .ZN(new_n698));
  XNOR2_X1  g273(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n699));
  XNOR2_X1  g274(.A(new_n699), .B(KEYINPUT91), .ZN(new_n700));
  XNOR2_X1  g275(.A(new_n698), .B(new_n700), .ZN(new_n701));
  XNOR2_X1  g276(.A(new_n695), .B(new_n701), .ZN(G229));
  INV_X1    g277(.A(G16), .ZN(new_n703));
  NAND2_X1  g278(.A1(new_n703), .A2(G23), .ZN(new_n704));
  INV_X1    g279(.A(G288), .ZN(new_n705));
  OAI21_X1  g280(.A(new_n704), .B1(new_n705), .B2(new_n703), .ZN(new_n706));
  XNOR2_X1  g281(.A(new_n706), .B(KEYINPUT33), .ZN(new_n707));
  INV_X1    g282(.A(G1976), .ZN(new_n708));
  XNOR2_X1  g283(.A(new_n707), .B(new_n708), .ZN(new_n709));
  XOR2_X1   g284(.A(KEYINPUT96), .B(G16), .Z(new_n710));
  NAND2_X1  g285(.A1(new_n710), .A2(G22), .ZN(new_n711));
  OAI21_X1  g286(.A(new_n711), .B1(G166), .B2(new_n710), .ZN(new_n712));
  XNOR2_X1  g287(.A(new_n712), .B(G1971), .ZN(new_n713));
  MUX2_X1   g288(.A(G6), .B(G305), .S(G16), .Z(new_n714));
  XOR2_X1   g289(.A(KEYINPUT32), .B(G1981), .Z(new_n715));
  XOR2_X1   g290(.A(new_n714), .B(new_n715), .Z(new_n716));
  NOR3_X1   g291(.A1(new_n709), .A2(new_n713), .A3(new_n716), .ZN(new_n717));
  INV_X1    g292(.A(KEYINPUT34), .ZN(new_n718));
  OR2_X1    g293(.A1(new_n717), .A2(new_n718), .ZN(new_n719));
  NAND2_X1  g294(.A1(new_n717), .A2(new_n718), .ZN(new_n720));
  INV_X1    g295(.A(G29), .ZN(new_n721));
  NAND2_X1  g296(.A1(new_n721), .A2(G25), .ZN(new_n722));
  NAND2_X1  g297(.A1(new_n481), .A2(G119), .ZN(new_n723));
  INV_X1    g298(.A(KEYINPUT94), .ZN(new_n724));
  XNOR2_X1  g299(.A(new_n723), .B(new_n724), .ZN(new_n725));
  INV_X1    g300(.A(G95), .ZN(new_n726));
  AND3_X1   g301(.A1(new_n726), .A2(new_n462), .A3(KEYINPUT95), .ZN(new_n727));
  AOI21_X1  g302(.A(KEYINPUT95), .B1(new_n726), .B2(new_n462), .ZN(new_n728));
  OAI221_X1 g303(.A(G2104), .B1(G107), .B2(new_n462), .C1(new_n727), .C2(new_n728), .ZN(new_n729));
  AND2_X1   g304(.A1(new_n725), .A2(new_n729), .ZN(new_n730));
  NAND2_X1  g305(.A1(new_n479), .A2(G131), .ZN(new_n731));
  XOR2_X1   g306(.A(new_n731), .B(KEYINPUT93), .Z(new_n732));
  NAND2_X1  g307(.A1(new_n730), .A2(new_n732), .ZN(new_n733));
  INV_X1    g308(.A(new_n733), .ZN(new_n734));
  OAI21_X1  g309(.A(new_n722), .B1(new_n734), .B2(new_n721), .ZN(new_n735));
  XOR2_X1   g310(.A(KEYINPUT35), .B(G1991), .Z(new_n736));
  AND2_X1   g311(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  NOR2_X1   g312(.A1(new_n735), .A2(new_n736), .ZN(new_n738));
  INV_X1    g313(.A(new_n710), .ZN(new_n739));
  NOR2_X1   g314(.A1(new_n739), .A2(G24), .ZN(new_n740));
  AOI21_X1  g315(.A(new_n740), .B1(new_n599), .B2(new_n739), .ZN(new_n741));
  XOR2_X1   g316(.A(new_n741), .B(G1986), .Z(new_n742));
  OAI22_X1  g317(.A1(new_n737), .A2(new_n738), .B1(KEYINPUT97), .B2(new_n742), .ZN(new_n743));
  AOI21_X1  g318(.A(new_n743), .B1(KEYINPUT97), .B2(new_n742), .ZN(new_n744));
  NAND3_X1  g319(.A1(new_n719), .A2(new_n720), .A3(new_n744), .ZN(new_n745));
  INV_X1    g320(.A(KEYINPUT98), .ZN(new_n746));
  NAND2_X1  g321(.A1(new_n746), .A2(KEYINPUT36), .ZN(new_n747));
  XNOR2_X1  g322(.A(new_n745), .B(new_n747), .ZN(new_n748));
  NAND2_X1  g323(.A1(new_n479), .A2(G139), .ZN(new_n749));
  XOR2_X1   g324(.A(new_n749), .B(KEYINPUT99), .Z(new_n750));
  NAND3_X1  g325(.A1(new_n462), .A2(G103), .A3(G2104), .ZN(new_n751));
  XOR2_X1   g326(.A(new_n751), .B(KEYINPUT25), .Z(new_n752));
  AOI22_X1  g327(.A1(new_n461), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n753));
  OAI211_X1 g328(.A(new_n750), .B(new_n752), .C1(new_n462), .C2(new_n753), .ZN(new_n754));
  OR2_X1    g329(.A1(new_n754), .A2(KEYINPUT100), .ZN(new_n755));
  NAND2_X1  g330(.A1(new_n754), .A2(KEYINPUT100), .ZN(new_n756));
  NAND2_X1  g331(.A1(new_n755), .A2(new_n756), .ZN(new_n757));
  MUX2_X1   g332(.A(G33), .B(new_n757), .S(G29), .Z(new_n758));
  NOR2_X1   g333(.A1(new_n758), .A2(G2072), .ZN(new_n759));
  XOR2_X1   g334(.A(new_n759), .B(KEYINPUT101), .Z(new_n760));
  NOR2_X1   g335(.A1(new_n739), .A2(G19), .ZN(new_n761));
  AOI21_X1  g336(.A(new_n761), .B1(new_n555), .B2(new_n739), .ZN(new_n762));
  XNOR2_X1  g337(.A(new_n762), .B(G1341), .ZN(new_n763));
  INV_X1    g338(.A(new_n763), .ZN(new_n764));
  NAND2_X1  g339(.A1(G162), .A2(G29), .ZN(new_n765));
  OAI21_X1  g340(.A(new_n765), .B1(G29), .B2(G35), .ZN(new_n766));
  XOR2_X1   g341(.A(KEYINPUT29), .B(G2090), .Z(new_n767));
  INV_X1    g342(.A(G1348), .ZN(new_n768));
  NAND2_X1  g343(.A1(new_n627), .A2(G16), .ZN(new_n769));
  OAI21_X1  g344(.A(new_n769), .B1(G4), .B2(G16), .ZN(new_n770));
  AOI22_X1  g345(.A1(new_n766), .A2(new_n767), .B1(new_n768), .B2(new_n770), .ZN(new_n771));
  OAI21_X1  g346(.A(new_n771), .B1(new_n766), .B2(new_n767), .ZN(new_n772));
  OR2_X1    g347(.A1(new_n770), .A2(new_n768), .ZN(new_n773));
  NAND2_X1  g348(.A1(new_n703), .A2(G21), .ZN(new_n774));
  OAI21_X1  g349(.A(new_n774), .B1(G168), .B2(new_n703), .ZN(new_n775));
  INV_X1    g350(.A(G1966), .ZN(new_n776));
  XNOR2_X1  g351(.A(new_n775), .B(new_n776), .ZN(new_n777));
  NAND2_X1  g352(.A1(new_n773), .A2(new_n777), .ZN(new_n778));
  NAND3_X1  g353(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n779));
  XNOR2_X1  g354(.A(new_n779), .B(KEYINPUT26), .ZN(new_n780));
  AOI21_X1  g355(.A(new_n780), .B1(G129), .B2(new_n481), .ZN(new_n781));
  AOI22_X1  g356(.A1(new_n479), .A2(G141), .B1(G105), .B2(new_n634), .ZN(new_n782));
  NAND2_X1  g357(.A1(new_n781), .A2(new_n782), .ZN(new_n783));
  MUX2_X1   g358(.A(G32), .B(new_n783), .S(G29), .Z(new_n784));
  XNOR2_X1  g359(.A(new_n784), .B(KEYINPUT102), .ZN(new_n785));
  XOR2_X1   g360(.A(KEYINPUT27), .B(G1996), .Z(new_n786));
  XNOR2_X1  g361(.A(new_n785), .B(new_n786), .ZN(new_n787));
  NAND2_X1  g362(.A1(new_n703), .A2(G5), .ZN(new_n788));
  OAI21_X1  g363(.A(new_n788), .B1(G171), .B2(new_n703), .ZN(new_n789));
  INV_X1    g364(.A(G1961), .ZN(new_n790));
  XNOR2_X1  g365(.A(new_n789), .B(new_n790), .ZN(new_n791));
  NAND2_X1  g366(.A1(new_n710), .A2(G20), .ZN(new_n792));
  XOR2_X1   g367(.A(new_n792), .B(KEYINPUT23), .Z(new_n793));
  AOI21_X1  g368(.A(new_n793), .B1(G299), .B2(G16), .ZN(new_n794));
  XNOR2_X1  g369(.A(new_n794), .B(G1956), .ZN(new_n795));
  NAND2_X1  g370(.A1(new_n791), .A2(new_n795), .ZN(new_n796));
  NOR4_X1   g371(.A1(new_n772), .A2(new_n778), .A3(new_n787), .A4(new_n796), .ZN(new_n797));
  INV_X1    g372(.A(G34), .ZN(new_n798));
  AND2_X1   g373(.A1(new_n798), .A2(KEYINPUT24), .ZN(new_n799));
  NOR2_X1   g374(.A1(new_n798), .A2(KEYINPUT24), .ZN(new_n800));
  OAI21_X1  g375(.A(new_n721), .B1(new_n799), .B2(new_n800), .ZN(new_n801));
  OAI21_X1  g376(.A(new_n801), .B1(G160), .B2(new_n721), .ZN(new_n802));
  XNOR2_X1  g377(.A(new_n802), .B(G2084), .ZN(new_n803));
  NAND2_X1  g378(.A1(new_n479), .A2(G140), .ZN(new_n804));
  NAND2_X1  g379(.A1(new_n481), .A2(G128), .ZN(new_n805));
  NOR2_X1   g380(.A1(new_n462), .A2(G116), .ZN(new_n806));
  OAI21_X1  g381(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n807));
  OAI211_X1 g382(.A(new_n804), .B(new_n805), .C1(new_n806), .C2(new_n807), .ZN(new_n808));
  NAND2_X1  g383(.A1(new_n808), .A2(G29), .ZN(new_n809));
  NAND2_X1  g384(.A1(new_n721), .A2(G26), .ZN(new_n810));
  XNOR2_X1  g385(.A(new_n810), .B(KEYINPUT28), .ZN(new_n811));
  NAND2_X1  g386(.A1(new_n809), .A2(new_n811), .ZN(new_n812));
  XOR2_X1   g387(.A(new_n812), .B(G2067), .Z(new_n813));
  NOR2_X1   g388(.A1(G27), .A2(G29), .ZN(new_n814));
  AOI21_X1  g389(.A(new_n814), .B1(G164), .B2(G29), .ZN(new_n815));
  INV_X1    g390(.A(G2078), .ZN(new_n816));
  XNOR2_X1  g391(.A(new_n815), .B(new_n816), .ZN(new_n817));
  XNOR2_X1  g392(.A(KEYINPUT30), .B(G28), .ZN(new_n818));
  OR2_X1    g393(.A1(KEYINPUT31), .A2(G11), .ZN(new_n819));
  NAND2_X1  g394(.A1(KEYINPUT31), .A2(G11), .ZN(new_n820));
  AOI22_X1  g395(.A1(new_n818), .A2(new_n721), .B1(new_n819), .B2(new_n820), .ZN(new_n821));
  OAI21_X1  g396(.A(new_n821), .B1(new_n647), .B2(new_n721), .ZN(new_n822));
  XNOR2_X1  g397(.A(new_n822), .B(KEYINPUT103), .ZN(new_n823));
  NAND3_X1  g398(.A1(new_n813), .A2(new_n817), .A3(new_n823), .ZN(new_n824));
  AOI211_X1 g399(.A(new_n803), .B(new_n824), .C1(new_n758), .C2(G2072), .ZN(new_n825));
  NAND4_X1  g400(.A1(new_n760), .A2(new_n764), .A3(new_n797), .A4(new_n825), .ZN(new_n826));
  NOR2_X1   g401(.A1(new_n748), .A2(new_n826), .ZN(G311));
  OR2_X1    g402(.A1(new_n748), .A2(new_n826), .ZN(G150));
  NAND2_X1  g403(.A1(new_n627), .A2(G559), .ZN(new_n829));
  XNOR2_X1  g404(.A(new_n829), .B(KEYINPUT38), .ZN(new_n830));
  AOI21_X1  g405(.A(new_n552), .B1(new_n542), .B2(new_n543), .ZN(new_n831));
  XNOR2_X1  g406(.A(KEYINPUT105), .B(G55), .ZN(new_n832));
  NAND2_X1  g407(.A1(new_n509), .A2(new_n832), .ZN(new_n833));
  INV_X1    g408(.A(G93), .ZN(new_n834));
  OAI21_X1  g409(.A(new_n833), .B1(new_n834), .B2(new_n551), .ZN(new_n835));
  OAI21_X1  g410(.A(G67), .B1(new_n526), .B2(new_n527), .ZN(new_n836));
  NAND2_X1  g411(.A1(G80), .A2(G543), .ZN(new_n837));
  NAND2_X1  g412(.A1(new_n836), .A2(new_n837), .ZN(new_n838));
  INV_X1    g413(.A(KEYINPUT104), .ZN(new_n839));
  AOI21_X1  g414(.A(new_n502), .B1(new_n838), .B2(new_n839), .ZN(new_n840));
  NAND3_X1  g415(.A1(new_n836), .A2(KEYINPUT104), .A3(new_n837), .ZN(new_n841));
  AOI21_X1  g416(.A(new_n835), .B1(new_n840), .B2(new_n841), .ZN(new_n842));
  AND3_X1   g417(.A1(new_n831), .A2(new_n545), .A3(new_n842), .ZN(new_n843));
  AOI21_X1  g418(.A(new_n842), .B1(new_n831), .B2(new_n545), .ZN(new_n844));
  NOR2_X1   g419(.A1(new_n843), .A2(new_n844), .ZN(new_n845));
  XOR2_X1   g420(.A(new_n830), .B(new_n845), .Z(new_n846));
  INV_X1    g421(.A(KEYINPUT39), .ZN(new_n847));
  AOI21_X1  g422(.A(G860), .B1(new_n846), .B2(new_n847), .ZN(new_n848));
  OAI21_X1  g423(.A(new_n848), .B1(new_n847), .B2(new_n846), .ZN(new_n849));
  XOR2_X1   g424(.A(new_n849), .B(KEYINPUT106), .Z(new_n850));
  INV_X1    g425(.A(new_n842), .ZN(new_n851));
  NAND2_X1  g426(.A1(new_n851), .A2(G860), .ZN(new_n852));
  XOR2_X1   g427(.A(new_n852), .B(KEYINPUT37), .Z(new_n853));
  NAND2_X1  g428(.A1(new_n850), .A2(new_n853), .ZN(G145));
  NAND3_X1  g429(.A1(new_n755), .A2(KEYINPUT107), .A3(new_n756), .ZN(new_n855));
  XNOR2_X1  g430(.A(new_n783), .B(new_n808), .ZN(new_n856));
  XNOR2_X1  g431(.A(new_n856), .B(new_n494), .ZN(new_n857));
  NAND2_X1  g432(.A1(new_n855), .A2(new_n857), .ZN(new_n858));
  XNOR2_X1  g433(.A(new_n733), .B(new_n636), .ZN(new_n859));
  INV_X1    g434(.A(new_n859), .ZN(new_n860));
  NAND2_X1  g435(.A1(new_n858), .A2(new_n860), .ZN(new_n861));
  NAND3_X1  g436(.A1(new_n855), .A2(new_n859), .A3(new_n857), .ZN(new_n862));
  NAND2_X1  g437(.A1(new_n861), .A2(new_n862), .ZN(new_n863));
  INV_X1    g438(.A(KEYINPUT107), .ZN(new_n864));
  NAND2_X1  g439(.A1(new_n757), .A2(new_n864), .ZN(new_n865));
  NAND2_X1  g440(.A1(new_n479), .A2(G142), .ZN(new_n866));
  NAND2_X1  g441(.A1(new_n481), .A2(G130), .ZN(new_n867));
  OR2_X1    g442(.A1(G106), .A2(G2105), .ZN(new_n868));
  OAI211_X1 g443(.A(new_n868), .B(G2104), .C1(G118), .C2(new_n462), .ZN(new_n869));
  NAND3_X1  g444(.A1(new_n866), .A2(new_n867), .A3(new_n869), .ZN(new_n870));
  INV_X1    g445(.A(new_n870), .ZN(new_n871));
  NAND2_X1  g446(.A1(new_n865), .A2(new_n871), .ZN(new_n872));
  NAND3_X1  g447(.A1(new_n757), .A2(new_n864), .A3(new_n870), .ZN(new_n873));
  NAND2_X1  g448(.A1(new_n872), .A2(new_n873), .ZN(new_n874));
  NAND2_X1  g449(.A1(new_n863), .A2(new_n874), .ZN(new_n875));
  XNOR2_X1  g450(.A(G160), .B(new_n647), .ZN(new_n876));
  XNOR2_X1  g451(.A(new_n876), .B(G162), .ZN(new_n877));
  NAND4_X1  g452(.A1(new_n861), .A2(new_n872), .A3(new_n862), .A4(new_n873), .ZN(new_n878));
  NAND3_X1  g453(.A1(new_n875), .A2(new_n877), .A3(new_n878), .ZN(new_n879));
  INV_X1    g454(.A(G37), .ZN(new_n880));
  AND2_X1   g455(.A1(new_n879), .A2(new_n880), .ZN(new_n881));
  AOI21_X1  g456(.A(new_n877), .B1(new_n875), .B2(new_n878), .ZN(new_n882));
  INV_X1    g457(.A(KEYINPUT108), .ZN(new_n883));
  NOR2_X1   g458(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  AOI211_X1 g459(.A(KEYINPUT108), .B(new_n877), .C1(new_n875), .C2(new_n878), .ZN(new_n885));
  OAI21_X1  g460(.A(new_n881), .B1(new_n884), .B2(new_n885), .ZN(new_n886));
  XNOR2_X1  g461(.A(new_n886), .B(KEYINPUT40), .ZN(G395));
  INV_X1    g462(.A(KEYINPUT111), .ZN(new_n888));
  INV_X1    g463(.A(KEYINPUT109), .ZN(new_n889));
  OAI21_X1  g464(.A(new_n889), .B1(new_n627), .B2(G299), .ZN(new_n890));
  INV_X1    g465(.A(new_n570), .ZN(new_n891));
  INV_X1    g466(.A(new_n572), .ZN(new_n892));
  NAND2_X1  g467(.A1(new_n891), .A2(new_n892), .ZN(new_n893));
  NAND4_X1  g468(.A1(new_n893), .A2(new_n615), .A3(KEYINPUT109), .A4(new_n566), .ZN(new_n894));
  INV_X1    g469(.A(KEYINPUT110), .ZN(new_n895));
  AND3_X1   g470(.A1(new_n890), .A2(new_n894), .A3(new_n895), .ZN(new_n896));
  AOI21_X1  g471(.A(new_n895), .B1(new_n890), .B2(new_n894), .ZN(new_n897));
  NAND2_X1  g472(.A1(new_n627), .A2(G299), .ZN(new_n898));
  INV_X1    g473(.A(new_n898), .ZN(new_n899));
  NOR3_X1   g474(.A1(new_n896), .A2(new_n897), .A3(new_n899), .ZN(new_n900));
  OAI21_X1  g475(.A(new_n888), .B1(new_n900), .B2(KEYINPUT41), .ZN(new_n901));
  NAND2_X1  g476(.A1(new_n890), .A2(new_n894), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n902), .A2(KEYINPUT110), .ZN(new_n903));
  NAND3_X1  g478(.A1(new_n890), .A2(new_n894), .A3(new_n895), .ZN(new_n904));
  NAND3_X1  g479(.A1(new_n903), .A2(new_n898), .A3(new_n904), .ZN(new_n905));
  INV_X1    g480(.A(KEYINPUT41), .ZN(new_n906));
  NAND3_X1  g481(.A1(new_n905), .A2(KEYINPUT111), .A3(new_n906), .ZN(new_n907));
  NAND4_X1  g482(.A1(new_n890), .A2(new_n894), .A3(KEYINPUT41), .A4(new_n898), .ZN(new_n908));
  NAND3_X1  g483(.A1(new_n901), .A2(new_n907), .A3(new_n908), .ZN(new_n909));
  XOR2_X1   g484(.A(new_n845), .B(new_n631), .Z(new_n910));
  NAND2_X1  g485(.A1(new_n909), .A2(new_n910), .ZN(new_n911));
  NOR2_X1   g486(.A1(new_n902), .A2(new_n899), .ZN(new_n912));
  NOR2_X1   g487(.A1(new_n910), .A2(new_n912), .ZN(new_n913));
  INV_X1    g488(.A(new_n913), .ZN(new_n914));
  XNOR2_X1  g489(.A(new_n514), .B(new_n599), .ZN(new_n915));
  XNOR2_X1  g490(.A(new_n705), .B(G305), .ZN(new_n916));
  OR2_X1    g491(.A1(new_n915), .A2(new_n916), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n915), .A2(new_n916), .ZN(new_n918));
  NAND2_X1  g493(.A1(new_n917), .A2(new_n918), .ZN(new_n919));
  XNOR2_X1  g494(.A(new_n919), .B(KEYINPUT42), .ZN(new_n920));
  AND3_X1   g495(.A1(new_n911), .A2(new_n914), .A3(new_n920), .ZN(new_n921));
  AOI21_X1  g496(.A(new_n920), .B1(new_n911), .B2(new_n914), .ZN(new_n922));
  OAI21_X1  g497(.A(G868), .B1(new_n921), .B2(new_n922), .ZN(new_n923));
  OAI21_X1  g498(.A(new_n923), .B1(G868), .B2(new_n842), .ZN(G295));
  OAI21_X1  g499(.A(new_n923), .B1(G868), .B2(new_n842), .ZN(G331));
  INV_X1    g500(.A(new_n919), .ZN(new_n926));
  OAI21_X1  g501(.A(G171), .B1(new_n843), .B2(new_n844), .ZN(new_n927));
  NAND2_X1  g502(.A1(new_n554), .A2(new_n851), .ZN(new_n928));
  NAND3_X1  g503(.A1(new_n831), .A2(new_n545), .A3(new_n842), .ZN(new_n929));
  NAND3_X1  g504(.A1(new_n928), .A2(G301), .A3(new_n929), .ZN(new_n930));
  AND3_X1   g505(.A1(new_n927), .A2(G168), .A3(new_n930), .ZN(new_n931));
  AOI21_X1  g506(.A(G168), .B1(new_n927), .B2(new_n930), .ZN(new_n932));
  NOR2_X1   g507(.A1(new_n931), .A2(new_n932), .ZN(new_n933));
  NAND4_X1  g508(.A1(new_n901), .A2(new_n933), .A3(new_n907), .A4(new_n908), .ZN(new_n934));
  OAI21_X1  g509(.A(new_n912), .B1(new_n931), .B2(new_n932), .ZN(new_n935));
  AOI21_X1  g510(.A(new_n926), .B1(new_n934), .B2(new_n935), .ZN(new_n936));
  INV_X1    g511(.A(new_n936), .ZN(new_n937));
  INV_X1    g512(.A(KEYINPUT43), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n937), .A2(new_n938), .ZN(new_n939));
  NAND3_X1  g514(.A1(new_n934), .A2(new_n926), .A3(new_n935), .ZN(new_n940));
  NAND2_X1  g515(.A1(new_n940), .A2(new_n880), .ZN(new_n941));
  NAND2_X1  g516(.A1(new_n933), .A2(KEYINPUT41), .ZN(new_n942));
  NAND2_X1  g517(.A1(new_n942), .A2(new_n912), .ZN(new_n943));
  NOR3_X1   g518(.A1(new_n931), .A2(new_n932), .A3(new_n906), .ZN(new_n944));
  AOI21_X1  g519(.A(new_n919), .B1(new_n944), .B2(new_n905), .ZN(new_n945));
  AOI21_X1  g520(.A(G37), .B1(new_n943), .B2(new_n945), .ZN(new_n946));
  AND2_X1   g521(.A1(new_n937), .A2(new_n946), .ZN(new_n947));
  OAI221_X1 g522(.A(KEYINPUT44), .B1(new_n939), .B2(new_n941), .C1(new_n947), .C2(new_n938), .ZN(new_n948));
  INV_X1    g523(.A(KEYINPUT112), .ZN(new_n949));
  OAI21_X1  g524(.A(KEYINPUT43), .B1(new_n941), .B2(new_n936), .ZN(new_n950));
  NAND3_X1  g525(.A1(new_n937), .A2(new_n946), .A3(new_n938), .ZN(new_n951));
  NAND2_X1  g526(.A1(new_n950), .A2(new_n951), .ZN(new_n952));
  INV_X1    g527(.A(KEYINPUT44), .ZN(new_n953));
  AOI21_X1  g528(.A(new_n949), .B1(new_n952), .B2(new_n953), .ZN(new_n954));
  AOI211_X1 g529(.A(KEYINPUT112), .B(KEYINPUT44), .C1(new_n950), .C2(new_n951), .ZN(new_n955));
  OAI21_X1  g530(.A(new_n948), .B1(new_n954), .B2(new_n955), .ZN(G397));
  INV_X1    g531(.A(G1384), .ZN(new_n957));
  NAND2_X1  g532(.A1(new_n494), .A2(new_n957), .ZN(new_n958));
  INV_X1    g533(.A(KEYINPUT45), .ZN(new_n959));
  NAND2_X1  g534(.A1(new_n958), .A2(new_n959), .ZN(new_n960));
  NAND2_X1  g535(.A1(new_n468), .A2(new_n469), .ZN(new_n961));
  NAND2_X1  g536(.A1(new_n961), .A2(G2105), .ZN(new_n962));
  AOI22_X1  g537(.A1(new_n479), .A2(G137), .B1(G101), .B2(new_n634), .ZN(new_n963));
  NAND3_X1  g538(.A1(new_n962), .A2(new_n963), .A3(G40), .ZN(new_n964));
  NOR2_X1   g539(.A1(new_n960), .A2(new_n964), .ZN(new_n965));
  INV_X1    g540(.A(new_n965), .ZN(new_n966));
  XNOR2_X1  g541(.A(new_n808), .B(G2067), .ZN(new_n967));
  NAND2_X1  g542(.A1(new_n967), .A2(new_n965), .ZN(new_n968));
  XOR2_X1   g543(.A(new_n968), .B(KEYINPUT113), .Z(new_n969));
  XNOR2_X1  g544(.A(new_n783), .B(G1996), .ZN(new_n970));
  AOI21_X1  g545(.A(new_n969), .B1(new_n965), .B2(new_n970), .ZN(new_n971));
  AND2_X1   g546(.A1(new_n734), .A2(new_n736), .ZN(new_n972));
  NAND2_X1  g547(.A1(new_n971), .A2(new_n972), .ZN(new_n973));
  OR2_X1    g548(.A1(new_n808), .A2(G2067), .ZN(new_n974));
  AOI21_X1  g549(.A(new_n966), .B1(new_n973), .B2(new_n974), .ZN(new_n975));
  NOR2_X1   g550(.A1(new_n734), .A2(new_n736), .ZN(new_n976));
  OAI21_X1  g551(.A(new_n965), .B1(new_n972), .B2(new_n976), .ZN(new_n977));
  NOR3_X1   g552(.A1(new_n966), .A2(G1986), .A3(G290), .ZN(new_n978));
  XOR2_X1   g553(.A(new_n978), .B(KEYINPUT48), .Z(new_n979));
  AND3_X1   g554(.A1(new_n971), .A2(new_n977), .A3(new_n979), .ZN(new_n980));
  OR3_X1    g555(.A1(new_n966), .A2(KEYINPUT46), .A3(G1996), .ZN(new_n981));
  OAI21_X1  g556(.A(KEYINPUT46), .B1(new_n966), .B2(G1996), .ZN(new_n982));
  OR2_X1    g557(.A1(new_n967), .A2(new_n783), .ZN(new_n983));
  AOI22_X1  g558(.A1(new_n981), .A2(new_n982), .B1(new_n965), .B2(new_n983), .ZN(new_n984));
  XNOR2_X1  g559(.A(new_n984), .B(KEYINPUT47), .ZN(new_n985));
  NOR3_X1   g560(.A1(new_n975), .A2(new_n980), .A3(new_n985), .ZN(new_n986));
  XNOR2_X1  g561(.A(KEYINPUT120), .B(KEYINPUT63), .ZN(new_n987));
  INV_X1    g562(.A(G1981), .ZN(new_n988));
  NAND4_X1  g563(.A1(new_n590), .A2(new_n988), .A3(new_n591), .A4(new_n592), .ZN(new_n989));
  OAI21_X1  g564(.A(new_n592), .B1(new_n589), .B2(new_n502), .ZN(new_n990));
  XNOR2_X1  g565(.A(KEYINPUT116), .B(G86), .ZN(new_n991));
  NOR2_X1   g566(.A1(new_n551), .A2(new_n991), .ZN(new_n992));
  OAI21_X1  g567(.A(G1981), .B1(new_n990), .B2(new_n992), .ZN(new_n993));
  AND3_X1   g568(.A1(new_n989), .A2(new_n993), .A3(KEYINPUT49), .ZN(new_n994));
  AOI21_X1  g569(.A(KEYINPUT49), .B1(new_n989), .B2(new_n993), .ZN(new_n995));
  OAI21_X1  g570(.A(G8), .B1(new_n964), .B2(new_n958), .ZN(new_n996));
  NOR3_X1   g571(.A1(new_n994), .A2(new_n995), .A3(new_n996), .ZN(new_n997));
  NAND3_X1  g572(.A1(new_n584), .A2(new_n587), .A3(G1976), .ZN(new_n998));
  INV_X1    g573(.A(new_n998), .ZN(new_n999));
  OAI21_X1  g574(.A(KEYINPUT52), .B1(new_n996), .B2(new_n999), .ZN(new_n1000));
  AOI21_X1  g575(.A(KEYINPUT52), .B1(G288), .B2(new_n708), .ZN(new_n1001));
  NAND4_X1  g576(.A1(new_n471), .A2(G40), .A3(new_n957), .A4(new_n494), .ZN(new_n1002));
  NAND4_X1  g577(.A1(new_n1001), .A2(G8), .A3(new_n1002), .A4(new_n998), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n1000), .A2(new_n1003), .ZN(new_n1004));
  NOR2_X1   g579(.A1(new_n997), .A2(new_n1004), .ZN(new_n1005));
  NAND3_X1  g580(.A1(new_n577), .A2(G8), .A3(new_n578), .ZN(new_n1006));
  NAND2_X1  g581(.A1(KEYINPUT115), .A2(KEYINPUT55), .ZN(new_n1007));
  NAND2_X1  g582(.A1(new_n1006), .A2(new_n1007), .ZN(new_n1008));
  XOR2_X1   g583(.A(KEYINPUT115), .B(KEYINPUT55), .Z(new_n1009));
  INV_X1    g584(.A(new_n1009), .ZN(new_n1010));
  NAND4_X1  g585(.A1(new_n577), .A2(G8), .A3(new_n578), .A4(new_n1010), .ZN(new_n1011));
  NAND2_X1  g586(.A1(new_n1008), .A2(new_n1011), .ZN(new_n1012));
  INV_X1    g587(.A(G8), .ZN(new_n1013));
  NAND3_X1  g588(.A1(new_n494), .A2(KEYINPUT45), .A3(new_n957), .ZN(new_n1014));
  AND3_X1   g589(.A1(new_n962), .A2(new_n963), .A3(G40), .ZN(new_n1015));
  NAND3_X1  g590(.A1(new_n960), .A2(new_n1014), .A3(new_n1015), .ZN(new_n1016));
  XNOR2_X1  g591(.A(KEYINPUT114), .B(G1971), .ZN(new_n1017));
  NAND2_X1  g592(.A1(new_n1016), .A2(new_n1017), .ZN(new_n1018));
  AOI21_X1  g593(.A(new_n964), .B1(KEYINPUT50), .B2(new_n958), .ZN(new_n1019));
  INV_X1    g594(.A(G2090), .ZN(new_n1020));
  INV_X1    g595(.A(KEYINPUT50), .ZN(new_n1021));
  NAND3_X1  g596(.A1(new_n494), .A2(new_n1021), .A3(new_n957), .ZN(new_n1022));
  NAND3_X1  g597(.A1(new_n1019), .A2(new_n1020), .A3(new_n1022), .ZN(new_n1023));
  AOI21_X1  g598(.A(new_n1013), .B1(new_n1018), .B2(new_n1023), .ZN(new_n1024));
  OAI21_X1  g599(.A(new_n1005), .B1(new_n1012), .B2(new_n1024), .ZN(new_n1025));
  NAND2_X1  g600(.A1(new_n1025), .A2(KEYINPUT121), .ZN(new_n1026));
  INV_X1    g601(.A(KEYINPUT121), .ZN(new_n1027));
  OAI211_X1 g602(.A(new_n1005), .B(new_n1027), .C1(new_n1012), .C2(new_n1024), .ZN(new_n1028));
  NAND2_X1  g603(.A1(new_n1026), .A2(new_n1028), .ZN(new_n1029));
  AND2_X1   g604(.A1(new_n1012), .A2(new_n1024), .ZN(new_n1030));
  INV_X1    g605(.A(KEYINPUT63), .ZN(new_n1031));
  NOR2_X1   g606(.A1(new_n1030), .A2(new_n1031), .ZN(new_n1032));
  NAND2_X1  g607(.A1(new_n1029), .A2(new_n1032), .ZN(new_n1033));
  INV_X1    g608(.A(KEYINPUT118), .ZN(new_n1034));
  AND3_X1   g609(.A1(new_n494), .A2(KEYINPUT45), .A3(new_n957), .ZN(new_n1035));
  AOI21_X1  g610(.A(KEYINPUT45), .B1(new_n494), .B2(new_n957), .ZN(new_n1036));
  NOR3_X1   g611(.A1(new_n1035), .A2(new_n1036), .A3(new_n964), .ZN(new_n1037));
  OAI21_X1  g612(.A(new_n1034), .B1(new_n1037), .B2(G1966), .ZN(new_n1038));
  INV_X1    g613(.A(new_n1038), .ZN(new_n1039));
  NAND3_X1  g614(.A1(new_n1016), .A2(KEYINPUT118), .A3(new_n776), .ZN(new_n1040));
  INV_X1    g615(.A(G2084), .ZN(new_n1041));
  NAND3_X1  g616(.A1(new_n1019), .A2(new_n1041), .A3(new_n1022), .ZN(new_n1042));
  NAND2_X1  g617(.A1(new_n1040), .A2(new_n1042), .ZN(new_n1043));
  OAI211_X1 g618(.A(G8), .B(G168), .C1(new_n1039), .C2(new_n1043), .ZN(new_n1044));
  OR2_X1    g619(.A1(new_n1044), .A2(KEYINPUT119), .ZN(new_n1045));
  NAND2_X1  g620(.A1(new_n1044), .A2(KEYINPUT119), .ZN(new_n1046));
  AND2_X1   g621(.A1(new_n1045), .A2(new_n1046), .ZN(new_n1047));
  OAI21_X1  g622(.A(new_n987), .B1(new_n1033), .B2(new_n1047), .ZN(new_n1048));
  OR3_X1    g623(.A1(new_n997), .A2(G1976), .A3(G288), .ZN(new_n1049));
  AOI21_X1  g624(.A(new_n996), .B1(new_n1049), .B2(new_n989), .ZN(new_n1050));
  AOI21_X1  g625(.A(new_n1050), .B1(new_n1005), .B2(new_n1030), .ZN(new_n1051));
  NAND2_X1  g626(.A1(new_n1048), .A2(new_n1051), .ZN(new_n1052));
  INV_X1    g627(.A(KEYINPUT125), .ZN(new_n1053));
  NAND4_X1  g628(.A1(new_n1038), .A2(G168), .A3(new_n1042), .A4(new_n1040), .ZN(new_n1054));
  OAI21_X1  g629(.A(G8), .B1(KEYINPUT124), .B2(KEYINPUT51), .ZN(new_n1055));
  INV_X1    g630(.A(new_n1055), .ZN(new_n1056));
  NAND2_X1  g631(.A1(KEYINPUT124), .A2(KEYINPUT51), .ZN(new_n1057));
  NAND3_X1  g632(.A1(new_n1054), .A2(new_n1056), .A3(new_n1057), .ZN(new_n1058));
  OAI211_X1 g633(.A(G8), .B(G286), .C1(new_n1039), .C2(new_n1043), .ZN(new_n1059));
  NAND2_X1  g634(.A1(new_n1058), .A2(new_n1059), .ZN(new_n1060));
  AOI21_X1  g635(.A(new_n1057), .B1(new_n1054), .B2(new_n1056), .ZN(new_n1061));
  OAI21_X1  g636(.A(new_n1053), .B1(new_n1060), .B2(new_n1061), .ZN(new_n1062));
  INV_X1    g637(.A(new_n1061), .ZN(new_n1063));
  NAND4_X1  g638(.A1(new_n1063), .A2(KEYINPUT125), .A3(new_n1059), .A4(new_n1058), .ZN(new_n1064));
  NAND2_X1  g639(.A1(new_n1062), .A2(new_n1064), .ZN(new_n1065));
  NAND2_X1  g640(.A1(new_n1065), .A2(KEYINPUT62), .ZN(new_n1066));
  INV_X1    g641(.A(KEYINPUT62), .ZN(new_n1067));
  NAND3_X1  g642(.A1(new_n1062), .A2(new_n1064), .A3(new_n1067), .ZN(new_n1068));
  NAND4_X1  g643(.A1(new_n960), .A2(new_n816), .A3(new_n1014), .A4(new_n1015), .ZN(new_n1069));
  INV_X1    g644(.A(KEYINPUT53), .ZN(new_n1070));
  NAND2_X1  g645(.A1(new_n1069), .A2(new_n1070), .ZN(new_n1071));
  NAND2_X1  g646(.A1(new_n958), .A2(KEYINPUT50), .ZN(new_n1072));
  NAND3_X1  g647(.A1(new_n1072), .A2(new_n1015), .A3(new_n1022), .ZN(new_n1073));
  NAND2_X1  g648(.A1(new_n1073), .A2(new_n790), .ZN(new_n1074));
  NOR2_X1   g649(.A1(new_n1036), .A2(new_n964), .ZN(new_n1075));
  NAND4_X1  g650(.A1(new_n1075), .A2(KEYINPUT53), .A3(new_n816), .A4(new_n1014), .ZN(new_n1076));
  NAND3_X1  g651(.A1(new_n1071), .A2(new_n1074), .A3(new_n1076), .ZN(new_n1077));
  NAND2_X1  g652(.A1(new_n1077), .A2(G171), .ZN(new_n1078));
  NAND2_X1  g653(.A1(new_n1078), .A2(KEYINPUT126), .ZN(new_n1079));
  INV_X1    g654(.A(KEYINPUT126), .ZN(new_n1080));
  NAND3_X1  g655(.A1(new_n1077), .A2(new_n1080), .A3(G171), .ZN(new_n1081));
  AND2_X1   g656(.A1(new_n1079), .A2(new_n1081), .ZN(new_n1082));
  NAND3_X1  g657(.A1(new_n1066), .A2(new_n1068), .A3(new_n1082), .ZN(new_n1083));
  AOI22_X1  g658(.A1(new_n1029), .A2(new_n1032), .B1(new_n1045), .B2(new_n1046), .ZN(new_n1084));
  INV_X1    g659(.A(KEYINPUT54), .ZN(new_n1085));
  NAND3_X1  g660(.A1(new_n1079), .A2(new_n1085), .A3(new_n1081), .ZN(new_n1086));
  NOR2_X1   g661(.A1(new_n1085), .A2(KEYINPUT127), .ZN(new_n1087));
  OR3_X1    g662(.A1(new_n1077), .A2(G171), .A3(new_n1087), .ZN(new_n1088));
  OR2_X1    g663(.A1(new_n1077), .A2(G171), .ZN(new_n1089));
  NAND3_X1  g664(.A1(new_n1089), .A2(new_n1078), .A3(new_n1087), .ZN(new_n1090));
  NAND3_X1  g665(.A1(new_n1086), .A2(new_n1088), .A3(new_n1090), .ZN(new_n1091));
  INV_X1    g666(.A(KEYINPUT117), .ZN(new_n1092));
  XNOR2_X1  g667(.A(new_n1022), .B(new_n1092), .ZN(new_n1093));
  NAND2_X1  g668(.A1(new_n1093), .A2(new_n1019), .ZN(new_n1094));
  INV_X1    g669(.A(G1956), .ZN(new_n1095));
  NAND2_X1  g670(.A1(new_n1094), .A2(new_n1095), .ZN(new_n1096));
  INV_X1    g671(.A(KEYINPUT122), .ZN(new_n1097));
  NAND2_X1  g672(.A1(G299), .A2(new_n1097), .ZN(new_n1098));
  XNOR2_X1  g673(.A(new_n1098), .B(KEYINPUT57), .ZN(new_n1099));
  XOR2_X1   g674(.A(KEYINPUT56), .B(G2072), .Z(new_n1100));
  NOR2_X1   g675(.A1(new_n1016), .A2(new_n1100), .ZN(new_n1101));
  INV_X1    g676(.A(new_n1101), .ZN(new_n1102));
  NAND3_X1  g677(.A1(new_n1096), .A2(new_n1099), .A3(new_n1102), .ZN(new_n1103));
  INV_X1    g678(.A(KEYINPUT57), .ZN(new_n1104));
  XNOR2_X1  g679(.A(new_n1098), .B(new_n1104), .ZN(new_n1105));
  AOI21_X1  g680(.A(G1956), .B1(new_n1093), .B2(new_n1019), .ZN(new_n1106));
  OAI21_X1  g681(.A(new_n1105), .B1(new_n1106), .B2(new_n1101), .ZN(new_n1107));
  NAND2_X1  g682(.A1(new_n1103), .A2(new_n1107), .ZN(new_n1108));
  INV_X1    g683(.A(KEYINPUT61), .ZN(new_n1109));
  NAND2_X1  g684(.A1(new_n1108), .A2(new_n1109), .ZN(new_n1110));
  INV_X1    g685(.A(G1996), .ZN(new_n1111));
  NAND2_X1  g686(.A1(new_n1037), .A2(new_n1111), .ZN(new_n1112));
  XOR2_X1   g687(.A(KEYINPUT58), .B(G1341), .Z(new_n1113));
  NAND2_X1  g688(.A1(new_n1002), .A2(new_n1113), .ZN(new_n1114));
  AOI21_X1  g689(.A(new_n554), .B1(new_n1112), .B2(new_n1114), .ZN(new_n1115));
  INV_X1    g690(.A(KEYINPUT59), .ZN(new_n1116));
  XNOR2_X1  g691(.A(new_n1115), .B(new_n1116), .ZN(new_n1117));
  NAND3_X1  g692(.A1(new_n1103), .A2(KEYINPUT61), .A3(new_n1107), .ZN(new_n1118));
  NAND2_X1  g693(.A1(new_n1073), .A2(new_n768), .ZN(new_n1119));
  OAI21_X1  g694(.A(new_n1119), .B1(G2067), .B2(new_n1002), .ZN(new_n1120));
  INV_X1    g695(.A(KEYINPUT60), .ZN(new_n1121));
  NAND2_X1  g696(.A1(new_n1120), .A2(new_n1121), .ZN(new_n1122));
  NOR2_X1   g697(.A1(new_n1002), .A2(G2067), .ZN(new_n1123));
  AOI21_X1  g698(.A(new_n1123), .B1(new_n768), .B2(new_n1073), .ZN(new_n1124));
  OR2_X1    g699(.A1(new_n627), .A2(KEYINPUT123), .ZN(new_n1125));
  NAND2_X1  g700(.A1(new_n627), .A2(KEYINPUT123), .ZN(new_n1126));
  NAND4_X1  g701(.A1(new_n1124), .A2(KEYINPUT60), .A3(new_n1125), .A4(new_n1126), .ZN(new_n1127));
  NOR2_X1   g702(.A1(new_n1120), .A2(new_n1121), .ZN(new_n1128));
  OAI211_X1 g703(.A(new_n1122), .B(new_n1127), .C1(new_n1128), .C2(new_n1125), .ZN(new_n1129));
  NAND4_X1  g704(.A1(new_n1110), .A2(new_n1117), .A3(new_n1118), .A4(new_n1129), .ZN(new_n1130));
  OAI21_X1  g705(.A(new_n1107), .B1(new_n615), .B2(new_n1124), .ZN(new_n1131));
  NAND2_X1  g706(.A1(new_n1131), .A2(new_n1103), .ZN(new_n1132));
  AOI21_X1  g707(.A(new_n1091), .B1(new_n1130), .B2(new_n1132), .ZN(new_n1133));
  AOI21_X1  g708(.A(new_n1084), .B1(new_n1133), .B2(new_n1065), .ZN(new_n1134));
  NAND2_X1  g709(.A1(new_n1083), .A2(new_n1134), .ZN(new_n1135));
  OAI21_X1  g710(.A(new_n1018), .B1(new_n1094), .B2(G2090), .ZN(new_n1136));
  AOI21_X1  g711(.A(new_n1012), .B1(G8), .B2(new_n1136), .ZN(new_n1137));
  NOR4_X1   g712(.A1(new_n1137), .A2(new_n1030), .A3(new_n997), .A4(new_n1004), .ZN(new_n1138));
  AOI21_X1  g713(.A(new_n1052), .B1(new_n1135), .B2(new_n1138), .ZN(new_n1139));
  XNOR2_X1  g714(.A(new_n599), .B(G1986), .ZN(new_n1140));
  OAI211_X1 g715(.A(new_n971), .B(new_n977), .C1(new_n966), .C2(new_n1140), .ZN(new_n1141));
  OAI21_X1  g716(.A(new_n986), .B1(new_n1139), .B2(new_n1141), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g717(.A(G319), .ZN(new_n1144));
  NOR4_X1   g718(.A1(G401), .A2(new_n1144), .A3(G227), .A4(G229), .ZN(new_n1145));
  NAND3_X1  g719(.A1(new_n1145), .A2(new_n886), .A3(new_n952), .ZN(G225));
  INV_X1    g720(.A(G225), .ZN(G308));
endmodule


