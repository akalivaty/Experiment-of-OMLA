//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 0 1 1 1 0 1 0 1 1 1 0 1 1 1 0 1 1 0 1 1 1 0 0 0 0 0 1 1 0 0 0 1 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 1 1 1 1 1 0 0 1 0 0 1 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:18:52 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n659, new_n660, new_n661, new_n663, new_n664, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n684, new_n685, new_n686, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n711, new_n712, new_n713, new_n714,
    new_n716, new_n717, new_n718, new_n719, new_n721, new_n723, new_n724,
    new_n725, new_n726, new_n727, new_n728, new_n729, new_n730, new_n731,
    new_n732, new_n733, new_n734, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n744, new_n745, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n825, new_n826, new_n828,
    new_n829, new_n830, new_n831, new_n833, new_n834, new_n835, new_n836,
    new_n837, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n873, new_n874,
    new_n875, new_n877, new_n878, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n894, new_n895, new_n896, new_n898, new_n899,
    new_n900, new_n901, new_n902, new_n903, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n924, new_n925, new_n926, new_n927, new_n929, new_n930, new_n931,
    new_n932, new_n934, new_n935;
  XNOR2_X1  g000(.A(KEYINPUT27), .B(G183gat), .ZN(new_n202));
  INV_X1    g001(.A(G190gat), .ZN(new_n203));
  NAND2_X1  g002(.A1(new_n202), .A2(new_n203), .ZN(new_n204));
  XOR2_X1   g003(.A(new_n204), .B(KEYINPUT28), .Z(new_n205));
  NAND2_X1  g004(.A1(G183gat), .A2(G190gat), .ZN(new_n206));
  AND2_X1   g005(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  NAND2_X1  g006(.A1(G169gat), .A2(G176gat), .ZN(new_n208));
  INV_X1    g007(.A(KEYINPUT26), .ZN(new_n209));
  NOR2_X1   g008(.A1(G169gat), .A2(G176gat), .ZN(new_n210));
  AND3_X1   g009(.A1(new_n210), .A2(KEYINPUT65), .A3(new_n209), .ZN(new_n211));
  AOI21_X1  g010(.A(KEYINPUT65), .B1(new_n210), .B2(new_n209), .ZN(new_n212));
  OAI221_X1 g011(.A(new_n208), .B1(new_n209), .B2(new_n210), .C1(new_n211), .C2(new_n212), .ZN(new_n213));
  INV_X1    g012(.A(G183gat), .ZN(new_n214));
  NAND2_X1  g013(.A1(new_n214), .A2(new_n203), .ZN(new_n215));
  AND3_X1   g014(.A1(new_n215), .A2(KEYINPUT24), .A3(new_n206), .ZN(new_n216));
  NOR2_X1   g015(.A1(new_n210), .A2(KEYINPUT23), .ZN(new_n217));
  OAI21_X1  g016(.A(new_n208), .B1(new_n206), .B2(KEYINPUT24), .ZN(new_n218));
  NOR3_X1   g017(.A1(new_n216), .A2(new_n217), .A3(new_n218), .ZN(new_n219));
  NAND2_X1  g018(.A1(new_n210), .A2(KEYINPUT23), .ZN(new_n220));
  OAI211_X1 g019(.A(new_n219), .B(new_n220), .C1(KEYINPUT64), .C2(KEYINPUT25), .ZN(new_n221));
  AOI21_X1  g020(.A(KEYINPUT25), .B1(new_n219), .B2(KEYINPUT64), .ZN(new_n222));
  NAND2_X1  g021(.A1(new_n219), .A2(new_n220), .ZN(new_n223));
  NAND2_X1  g022(.A1(new_n222), .A2(new_n223), .ZN(new_n224));
  AOI22_X1  g023(.A1(new_n207), .A2(new_n213), .B1(new_n221), .B2(new_n224), .ZN(new_n225));
  XOR2_X1   g024(.A(KEYINPUT66), .B(G120gat), .Z(new_n226));
  NAND2_X1  g025(.A1(new_n226), .A2(G113gat), .ZN(new_n227));
  XNOR2_X1  g026(.A(G127gat), .B(G134gat), .ZN(new_n228));
  INV_X1    g027(.A(G113gat), .ZN(new_n229));
  INV_X1    g028(.A(G120gat), .ZN(new_n230));
  AOI21_X1  g029(.A(KEYINPUT1), .B1(new_n229), .B2(new_n230), .ZN(new_n231));
  NAND3_X1  g030(.A1(new_n227), .A2(new_n228), .A3(new_n231), .ZN(new_n232));
  INV_X1    g031(.A(new_n232), .ZN(new_n233));
  INV_X1    g032(.A(KEYINPUT67), .ZN(new_n234));
  NAND2_X1  g033(.A1(new_n233), .A2(new_n234), .ZN(new_n235));
  NOR2_X1   g034(.A1(new_n229), .A2(new_n230), .ZN(new_n236));
  INV_X1    g035(.A(new_n236), .ZN(new_n237));
  AOI21_X1  g036(.A(new_n228), .B1(new_n237), .B2(new_n231), .ZN(new_n238));
  NAND2_X1  g037(.A1(new_n232), .A2(KEYINPUT67), .ZN(new_n239));
  OAI21_X1  g038(.A(new_n235), .B1(new_n238), .B2(new_n239), .ZN(new_n240));
  NAND2_X1  g039(.A1(new_n225), .A2(new_n240), .ZN(new_n241));
  NAND2_X1  g040(.A1(new_n224), .A2(new_n221), .ZN(new_n242));
  NAND3_X1  g041(.A1(new_n205), .A2(new_n213), .A3(new_n206), .ZN(new_n243));
  NAND2_X1  g042(.A1(new_n242), .A2(new_n243), .ZN(new_n244));
  INV_X1    g043(.A(new_n240), .ZN(new_n245));
  NAND2_X1  g044(.A1(new_n244), .A2(new_n245), .ZN(new_n246));
  AND2_X1   g045(.A1(new_n241), .A2(new_n246), .ZN(new_n247));
  INV_X1    g046(.A(G227gat), .ZN(new_n248));
  INV_X1    g047(.A(G233gat), .ZN(new_n249));
  NOR2_X1   g048(.A1(new_n248), .A2(new_n249), .ZN(new_n250));
  INV_X1    g049(.A(new_n250), .ZN(new_n251));
  OAI21_X1  g050(.A(KEYINPUT32), .B1(new_n247), .B2(new_n251), .ZN(new_n252));
  INV_X1    g051(.A(KEYINPUT33), .ZN(new_n253));
  OAI21_X1  g052(.A(new_n253), .B1(new_n247), .B2(new_n251), .ZN(new_n254));
  XOR2_X1   g053(.A(G15gat), .B(G43gat), .Z(new_n255));
  XNOR2_X1  g054(.A(G71gat), .B(G99gat), .ZN(new_n256));
  XNOR2_X1  g055(.A(new_n255), .B(new_n256), .ZN(new_n257));
  NAND3_X1  g056(.A1(new_n252), .A2(new_n254), .A3(new_n257), .ZN(new_n258));
  INV_X1    g057(.A(KEYINPUT32), .ZN(new_n259));
  NAND2_X1  g058(.A1(new_n241), .A2(new_n246), .ZN(new_n260));
  AOI221_X4 g059(.A(new_n259), .B1(KEYINPUT33), .B2(new_n257), .C1(new_n260), .C2(new_n250), .ZN(new_n261));
  INV_X1    g060(.A(new_n261), .ZN(new_n262));
  XOR2_X1   g061(.A(KEYINPUT68), .B(KEYINPUT34), .Z(new_n263));
  INV_X1    g062(.A(new_n263), .ZN(new_n264));
  OAI21_X1  g063(.A(new_n264), .B1(new_n260), .B2(new_n250), .ZN(new_n265));
  NAND2_X1  g064(.A1(KEYINPUT68), .A2(KEYINPUT34), .ZN(new_n266));
  NAND4_X1  g065(.A1(new_n241), .A2(new_n246), .A3(new_n251), .A4(new_n266), .ZN(new_n267));
  NAND2_X1  g066(.A1(new_n265), .A2(new_n267), .ZN(new_n268));
  INV_X1    g067(.A(new_n268), .ZN(new_n269));
  NAND3_X1  g068(.A1(new_n258), .A2(new_n262), .A3(new_n269), .ZN(new_n270));
  AOI21_X1  g069(.A(new_n251), .B1(new_n241), .B2(new_n246), .ZN(new_n271));
  OAI21_X1  g070(.A(new_n257), .B1(new_n271), .B2(KEYINPUT33), .ZN(new_n272));
  NOR2_X1   g071(.A1(new_n271), .A2(new_n259), .ZN(new_n273));
  NOR2_X1   g072(.A1(new_n272), .A2(new_n273), .ZN(new_n274));
  OAI21_X1  g073(.A(new_n268), .B1(new_n274), .B2(new_n261), .ZN(new_n275));
  AOI21_X1  g074(.A(KEYINPUT36), .B1(new_n270), .B2(new_n275), .ZN(new_n276));
  INV_X1    g075(.A(KEYINPUT69), .ZN(new_n277));
  OAI211_X1 g076(.A(new_n277), .B(new_n268), .C1(new_n274), .C2(new_n261), .ZN(new_n278));
  NAND2_X1  g077(.A1(new_n270), .A2(new_n275), .ZN(new_n279));
  OAI21_X1  g078(.A(new_n278), .B1(new_n279), .B2(new_n277), .ZN(new_n280));
  AOI21_X1  g079(.A(new_n276), .B1(new_n280), .B2(KEYINPUT36), .ZN(new_n281));
  XNOR2_X1  g080(.A(G155gat), .B(G162gat), .ZN(new_n282));
  XOR2_X1   g081(.A(G141gat), .B(G148gat), .Z(new_n283));
  INV_X1    g082(.A(KEYINPUT2), .ZN(new_n284));
  AOI21_X1  g083(.A(new_n282), .B1(new_n283), .B2(new_n284), .ZN(new_n285));
  INV_X1    g084(.A(KEYINPUT76), .ZN(new_n286));
  XNOR2_X1  g085(.A(new_n282), .B(KEYINPUT74), .ZN(new_n287));
  NAND2_X1  g086(.A1(new_n287), .A2(new_n283), .ZN(new_n288));
  XOR2_X1   g087(.A(KEYINPUT75), .B(G162gat), .Z(new_n289));
  INV_X1    g088(.A(G155gat), .ZN(new_n290));
  OAI21_X1  g089(.A(KEYINPUT2), .B1(new_n289), .B2(new_n290), .ZN(new_n291));
  INV_X1    g090(.A(new_n291), .ZN(new_n292));
  OAI21_X1  g091(.A(new_n286), .B1(new_n288), .B2(new_n292), .ZN(new_n293));
  NAND4_X1  g092(.A1(new_n287), .A2(KEYINPUT76), .A3(new_n291), .A4(new_n283), .ZN(new_n294));
  AOI21_X1  g093(.A(new_n285), .B1(new_n293), .B2(new_n294), .ZN(new_n295));
  NAND2_X1  g094(.A1(new_n295), .A2(new_n240), .ZN(new_n296));
  NAND2_X1  g095(.A1(new_n296), .A2(KEYINPUT4), .ZN(new_n297));
  INV_X1    g096(.A(KEYINPUT4), .ZN(new_n298));
  NAND3_X1  g097(.A1(new_n295), .A2(new_n298), .A3(new_n240), .ZN(new_n299));
  NAND3_X1  g098(.A1(new_n297), .A2(KEYINPUT81), .A3(new_n299), .ZN(new_n300));
  INV_X1    g099(.A(KEYINPUT81), .ZN(new_n301));
  NAND3_X1  g100(.A1(new_n296), .A2(new_n301), .A3(KEYINPUT4), .ZN(new_n302));
  NAND2_X1  g101(.A1(new_n300), .A2(new_n302), .ZN(new_n303));
  INV_X1    g102(.A(KEYINPUT5), .ZN(new_n304));
  NAND2_X1  g103(.A1(G225gat), .A2(G233gat), .ZN(new_n305));
  INV_X1    g104(.A(new_n295), .ZN(new_n306));
  NOR2_X1   g105(.A1(new_n306), .A2(KEYINPUT3), .ZN(new_n307));
  INV_X1    g106(.A(KEYINPUT3), .ZN(new_n308));
  OAI21_X1  g107(.A(new_n245), .B1(new_n295), .B2(new_n308), .ZN(new_n309));
  OAI211_X1 g108(.A(new_n304), .B(new_n305), .C1(new_n307), .C2(new_n309), .ZN(new_n310));
  OAI21_X1  g109(.A(KEYINPUT82), .B1(new_n303), .B2(new_n310), .ZN(new_n311));
  INV_X1    g110(.A(new_n311), .ZN(new_n312));
  NOR3_X1   g111(.A1(new_n303), .A2(new_n310), .A3(KEYINPUT82), .ZN(new_n313));
  INV_X1    g112(.A(KEYINPUT77), .ZN(new_n314));
  NAND2_X1  g113(.A1(new_n297), .A2(new_n314), .ZN(new_n315));
  INV_X1    g114(.A(KEYINPUT78), .ZN(new_n316));
  NAND2_X1  g115(.A1(new_n299), .A2(new_n316), .ZN(new_n317));
  NAND4_X1  g116(.A1(new_n295), .A2(KEYINPUT78), .A3(new_n298), .A4(new_n240), .ZN(new_n318));
  NAND3_X1  g117(.A1(new_n296), .A2(KEYINPUT77), .A3(KEYINPUT4), .ZN(new_n319));
  NAND4_X1  g118(.A1(new_n315), .A2(new_n317), .A3(new_n318), .A4(new_n319), .ZN(new_n320));
  NOR2_X1   g119(.A1(new_n307), .A2(new_n309), .ZN(new_n321));
  INV_X1    g120(.A(new_n305), .ZN(new_n322));
  NOR2_X1   g121(.A1(new_n321), .A2(new_n322), .ZN(new_n323));
  AND2_X1   g122(.A1(new_n320), .A2(new_n323), .ZN(new_n324));
  NAND2_X1  g123(.A1(new_n306), .A2(new_n245), .ZN(new_n325));
  INV_X1    g124(.A(KEYINPUT79), .ZN(new_n326));
  AOI21_X1  g125(.A(new_n326), .B1(new_n295), .B2(new_n240), .ZN(new_n327));
  XNOR2_X1  g126(.A(new_n325), .B(new_n327), .ZN(new_n328));
  OAI21_X1  g127(.A(KEYINPUT5), .B1(new_n328), .B2(new_n305), .ZN(new_n329));
  OAI22_X1  g128(.A1(new_n312), .A2(new_n313), .B1(new_n324), .B2(new_n329), .ZN(new_n330));
  XOR2_X1   g129(.A(G1gat), .B(G29gat), .Z(new_n331));
  XNOR2_X1  g130(.A(G57gat), .B(G85gat), .ZN(new_n332));
  XNOR2_X1  g131(.A(new_n331), .B(new_n332), .ZN(new_n333));
  XNOR2_X1  g132(.A(KEYINPUT80), .B(KEYINPUT0), .ZN(new_n334));
  XNOR2_X1  g133(.A(new_n333), .B(new_n334), .ZN(new_n335));
  NAND2_X1  g134(.A1(new_n330), .A2(new_n335), .ZN(new_n336));
  OR3_X1    g135(.A1(new_n303), .A2(KEYINPUT82), .A3(new_n310), .ZN(new_n337));
  NAND2_X1  g136(.A1(new_n337), .A2(new_n311), .ZN(new_n338));
  INV_X1    g137(.A(new_n335), .ZN(new_n339));
  NAND2_X1  g138(.A1(new_n320), .A2(new_n323), .ZN(new_n340));
  OAI211_X1 g139(.A(new_n340), .B(KEYINPUT5), .C1(new_n305), .C2(new_n328), .ZN(new_n341));
  NAND3_X1  g140(.A1(new_n338), .A2(new_n339), .A3(new_n341), .ZN(new_n342));
  INV_X1    g141(.A(KEYINPUT6), .ZN(new_n343));
  NAND3_X1  g142(.A1(new_n336), .A2(new_n342), .A3(new_n343), .ZN(new_n344));
  AOI21_X1  g143(.A(new_n339), .B1(new_n338), .B2(new_n341), .ZN(new_n345));
  NAND2_X1  g144(.A1(new_n345), .A2(KEYINPUT6), .ZN(new_n346));
  NAND2_X1  g145(.A1(new_n344), .A2(new_n346), .ZN(new_n347));
  INV_X1    g146(.A(KEYINPUT73), .ZN(new_n348));
  NAND2_X1  g147(.A1(G226gat), .A2(G233gat), .ZN(new_n349));
  OAI21_X1  g148(.A(new_n348), .B1(new_n225), .B2(new_n349), .ZN(new_n350));
  NAND4_X1  g149(.A1(new_n244), .A2(KEYINPUT73), .A3(G226gat), .A4(G233gat), .ZN(new_n351));
  NOR2_X1   g150(.A1(new_n225), .A2(KEYINPUT29), .ZN(new_n352));
  XNOR2_X1  g151(.A(new_n349), .B(KEYINPUT72), .ZN(new_n353));
  OAI211_X1 g152(.A(new_n350), .B(new_n351), .C1(new_n352), .C2(new_n353), .ZN(new_n354));
  XOR2_X1   g153(.A(G211gat), .B(G218gat), .Z(new_n355));
  XNOR2_X1  g154(.A(new_n355), .B(KEYINPUT70), .ZN(new_n356));
  INV_X1    g155(.A(G211gat), .ZN(new_n357));
  INV_X1    g156(.A(G218gat), .ZN(new_n358));
  NOR2_X1   g157(.A1(new_n357), .A2(new_n358), .ZN(new_n359));
  NOR2_X1   g158(.A1(G197gat), .A2(G204gat), .ZN(new_n360));
  AND2_X1   g159(.A1(G197gat), .A2(G204gat), .ZN(new_n361));
  OAI22_X1  g160(.A1(new_n359), .A2(KEYINPUT22), .B1(new_n360), .B2(new_n361), .ZN(new_n362));
  NAND2_X1  g161(.A1(new_n362), .A2(KEYINPUT71), .ZN(new_n363));
  XNOR2_X1  g162(.A(new_n356), .B(new_n363), .ZN(new_n364));
  INV_X1    g163(.A(new_n364), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n354), .A2(new_n365), .ZN(new_n366));
  OAI21_X1  g165(.A(new_n349), .B1(new_n225), .B2(KEYINPUT29), .ZN(new_n367));
  NAND2_X1  g166(.A1(new_n244), .A2(new_n353), .ZN(new_n368));
  AND2_X1   g167(.A1(new_n367), .A2(new_n368), .ZN(new_n369));
  NAND2_X1  g168(.A1(new_n369), .A2(new_n364), .ZN(new_n370));
  NAND2_X1  g169(.A1(new_n366), .A2(new_n370), .ZN(new_n371));
  XNOR2_X1  g170(.A(G8gat), .B(G36gat), .ZN(new_n372));
  XNOR2_X1  g171(.A(G64gat), .B(G92gat), .ZN(new_n373));
  XOR2_X1   g172(.A(new_n372), .B(new_n373), .Z(new_n374));
  INV_X1    g173(.A(new_n374), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n371), .A2(new_n375), .ZN(new_n376));
  NAND3_X1  g175(.A1(new_n366), .A2(new_n370), .A3(new_n374), .ZN(new_n377));
  NAND3_X1  g176(.A1(new_n376), .A2(KEYINPUT30), .A3(new_n377), .ZN(new_n378));
  OR3_X1    g177(.A1(new_n371), .A2(KEYINPUT30), .A3(new_n375), .ZN(new_n379));
  NAND2_X1  g178(.A1(new_n378), .A2(new_n379), .ZN(new_n380));
  NAND2_X1  g179(.A1(new_n347), .A2(new_n380), .ZN(new_n381));
  INV_X1    g180(.A(KEYINPUT84), .ZN(new_n382));
  XOR2_X1   g181(.A(G78gat), .B(G106gat), .Z(new_n383));
  XNOR2_X1  g182(.A(KEYINPUT31), .B(G50gat), .ZN(new_n384));
  XNOR2_X1  g183(.A(new_n383), .B(new_n384), .ZN(new_n385));
  INV_X1    g184(.A(G22gat), .ZN(new_n386));
  AOI21_X1  g185(.A(KEYINPUT29), .B1(new_n295), .B2(new_n308), .ZN(new_n387));
  OR2_X1    g186(.A1(new_n387), .A2(new_n364), .ZN(new_n388));
  NAND2_X1  g187(.A1(G228gat), .A2(G233gat), .ZN(new_n389));
  OAI21_X1  g188(.A(new_n308), .B1(new_n365), .B2(KEYINPUT29), .ZN(new_n390));
  AOI21_X1  g189(.A(new_n389), .B1(new_n390), .B2(new_n306), .ZN(new_n391));
  NAND2_X1  g190(.A1(new_n388), .A2(new_n391), .ZN(new_n392));
  OR2_X1    g191(.A1(new_n356), .A2(new_n362), .ZN(new_n393));
  AOI21_X1  g192(.A(KEYINPUT29), .B1(new_n356), .B2(new_n362), .ZN(new_n394));
  AOI21_X1  g193(.A(KEYINPUT3), .B1(new_n393), .B2(new_n394), .ZN(new_n395));
  OAI22_X1  g194(.A1(new_n387), .A2(new_n364), .B1(new_n295), .B2(new_n395), .ZN(new_n396));
  NAND2_X1  g195(.A1(new_n396), .A2(new_n389), .ZN(new_n397));
  AOI21_X1  g196(.A(new_n386), .B1(new_n392), .B2(new_n397), .ZN(new_n398));
  INV_X1    g197(.A(KEYINPUT83), .ZN(new_n399));
  OAI211_X1 g198(.A(new_n382), .B(new_n385), .C1(new_n398), .C2(new_n399), .ZN(new_n400));
  INV_X1    g199(.A(new_n400), .ZN(new_n401));
  AOI22_X1  g200(.A1(new_n388), .A2(new_n391), .B1(new_n396), .B2(new_n389), .ZN(new_n402));
  OAI21_X1  g201(.A(KEYINPUT83), .B1(new_n402), .B2(new_n386), .ZN(new_n403));
  AOI21_X1  g202(.A(new_n382), .B1(new_n403), .B2(new_n385), .ZN(new_n404));
  INV_X1    g203(.A(new_n402), .ZN(new_n405));
  NOR2_X1   g204(.A1(new_n405), .A2(G22gat), .ZN(new_n406));
  OAI22_X1  g205(.A1(new_n401), .A2(new_n404), .B1(new_n398), .B2(new_n406), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n403), .A2(new_n385), .ZN(new_n408));
  NAND2_X1  g207(.A1(new_n408), .A2(KEYINPUT84), .ZN(new_n409));
  NOR2_X1   g208(.A1(new_n406), .A2(new_n398), .ZN(new_n410));
  NAND3_X1  g209(.A1(new_n409), .A2(new_n410), .A3(new_n400), .ZN(new_n411));
  NAND2_X1  g210(.A1(new_n407), .A2(new_n411), .ZN(new_n412));
  AOI21_X1  g211(.A(new_n281), .B1(new_n381), .B2(new_n412), .ZN(new_n413));
  INV_X1    g212(.A(KEYINPUT85), .ZN(new_n414));
  AOI21_X1  g213(.A(new_n414), .B1(new_n344), .B2(new_n346), .ZN(new_n415));
  AOI21_X1  g214(.A(KEYINPUT85), .B1(new_n345), .B2(KEYINPUT6), .ZN(new_n416));
  OAI21_X1  g215(.A(new_n375), .B1(new_n371), .B2(KEYINPUT37), .ZN(new_n417));
  INV_X1    g216(.A(KEYINPUT37), .ZN(new_n418));
  AOI21_X1  g217(.A(new_n418), .B1(new_n366), .B2(new_n370), .ZN(new_n419));
  OAI21_X1  g218(.A(KEYINPUT38), .B1(new_n417), .B2(new_n419), .ZN(new_n420));
  NAND2_X1  g219(.A1(new_n369), .A2(new_n365), .ZN(new_n421));
  NAND2_X1  g220(.A1(new_n421), .A2(KEYINPUT37), .ZN(new_n422));
  AOI21_X1  g221(.A(new_n422), .B1(new_n364), .B2(new_n354), .ZN(new_n423));
  OR2_X1    g222(.A1(new_n423), .A2(KEYINPUT38), .ZN(new_n424));
  OAI211_X1 g223(.A(new_n420), .B(new_n377), .C1(new_n424), .C2(new_n417), .ZN(new_n425));
  NOR3_X1   g224(.A1(new_n415), .A2(new_n416), .A3(new_n425), .ZN(new_n426));
  INV_X1    g225(.A(new_n412), .ZN(new_n427));
  INV_X1    g226(.A(KEYINPUT39), .ZN(new_n428));
  AOI21_X1  g227(.A(new_n428), .B1(new_n328), .B2(new_n305), .ZN(new_n429));
  OAI21_X1  g228(.A(new_n322), .B1(new_n303), .B2(new_n321), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n429), .A2(new_n430), .ZN(new_n431));
  OAI211_X1 g230(.A(new_n431), .B(new_n339), .C1(KEYINPUT39), .C2(new_n430), .ZN(new_n432));
  INV_X1    g231(.A(KEYINPUT40), .ZN(new_n433));
  OAI21_X1  g232(.A(new_n336), .B1(new_n432), .B2(new_n433), .ZN(new_n434));
  INV_X1    g233(.A(new_n380), .ZN(new_n435));
  NAND2_X1  g234(.A1(new_n432), .A2(new_n433), .ZN(new_n436));
  NAND2_X1  g235(.A1(new_n435), .A2(new_n436), .ZN(new_n437));
  OAI21_X1  g236(.A(new_n427), .B1(new_n434), .B2(new_n437), .ZN(new_n438));
  OAI21_X1  g237(.A(new_n413), .B1(new_n426), .B2(new_n438), .ZN(new_n439));
  NOR3_X1   g238(.A1(new_n435), .A2(KEYINPUT35), .A3(new_n279), .ZN(new_n440));
  OAI211_X1 g239(.A(new_n427), .B(new_n440), .C1(new_n415), .C2(new_n416), .ZN(new_n441));
  INV_X1    g240(.A(KEYINPUT35), .ZN(new_n442));
  AND3_X1   g241(.A1(new_n280), .A2(new_n407), .A3(new_n411), .ZN(new_n443));
  AOI21_X1  g242(.A(new_n435), .B1(new_n344), .B2(new_n346), .ZN(new_n444));
  AOI21_X1  g243(.A(new_n442), .B1(new_n443), .B2(new_n444), .ZN(new_n445));
  OAI21_X1  g244(.A(new_n441), .B1(new_n445), .B2(KEYINPUT86), .ZN(new_n446));
  INV_X1    g245(.A(KEYINPUT86), .ZN(new_n447));
  AOI211_X1 g246(.A(new_n447), .B(new_n442), .C1(new_n443), .C2(new_n444), .ZN(new_n448));
  OAI21_X1  g247(.A(new_n439), .B1(new_n446), .B2(new_n448), .ZN(new_n449));
  NAND2_X1  g248(.A1(G71gat), .A2(G78gat), .ZN(new_n450));
  INV_X1    g249(.A(KEYINPUT9), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n450), .A2(new_n451), .ZN(new_n452));
  INV_X1    g251(.A(G57gat), .ZN(new_n453));
  NOR2_X1   g252(.A1(new_n453), .A2(G64gat), .ZN(new_n454));
  INV_X1    g253(.A(G64gat), .ZN(new_n455));
  NOR2_X1   g254(.A1(new_n455), .A2(G57gat), .ZN(new_n456));
  OAI211_X1 g255(.A(KEYINPUT93), .B(new_n452), .C1(new_n454), .C2(new_n456), .ZN(new_n457));
  XNOR2_X1  g256(.A(G71gat), .B(G78gat), .ZN(new_n458));
  INV_X1    g257(.A(new_n458), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n457), .A2(new_n459), .ZN(new_n460));
  INV_X1    g259(.A(KEYINPUT93), .ZN(new_n461));
  NAND2_X1  g260(.A1(new_n455), .A2(G57gat), .ZN(new_n462));
  NAND2_X1  g261(.A1(new_n453), .A2(G64gat), .ZN(new_n463));
  AOI21_X1  g262(.A(new_n461), .B1(new_n462), .B2(new_n463), .ZN(new_n464));
  NAND3_X1  g263(.A1(new_n464), .A2(new_n458), .A3(new_n452), .ZN(new_n465));
  NAND2_X1  g264(.A1(new_n460), .A2(new_n465), .ZN(new_n466));
  INV_X1    g265(.A(KEYINPUT21), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  NAND2_X1  g267(.A1(G231gat), .A2(G233gat), .ZN(new_n469));
  XNOR2_X1  g268(.A(new_n468), .B(new_n469), .ZN(new_n470));
  INV_X1    g269(.A(G127gat), .ZN(new_n471));
  XNOR2_X1  g270(.A(new_n470), .B(new_n471), .ZN(new_n472));
  INV_X1    g271(.A(G1gat), .ZN(new_n473));
  NAND2_X1  g272(.A1(new_n473), .A2(KEYINPUT16), .ZN(new_n474));
  INV_X1    g273(.A(G15gat), .ZN(new_n475));
  NAND2_X1  g274(.A1(new_n475), .A2(G22gat), .ZN(new_n476));
  NAND2_X1  g275(.A1(new_n386), .A2(G15gat), .ZN(new_n477));
  AND3_X1   g276(.A1(new_n474), .A2(new_n476), .A3(new_n477), .ZN(new_n478));
  AOI21_X1  g277(.A(G1gat), .B1(new_n476), .B2(new_n477), .ZN(new_n479));
  OAI21_X1  g278(.A(G8gat), .B1(new_n478), .B2(new_n479), .ZN(new_n480));
  NAND3_X1  g279(.A1(new_n474), .A2(new_n476), .A3(new_n477), .ZN(new_n481));
  INV_X1    g280(.A(G8gat), .ZN(new_n482));
  XNOR2_X1  g281(.A(G15gat), .B(G22gat), .ZN(new_n483));
  OAI211_X1 g282(.A(new_n481), .B(new_n482), .C1(G1gat), .C2(new_n483), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n480), .A2(new_n484), .ZN(new_n485));
  NOR2_X1   g284(.A1(new_n457), .A2(new_n459), .ZN(new_n486));
  AOI21_X1  g285(.A(new_n458), .B1(new_n464), .B2(new_n452), .ZN(new_n487));
  NOR2_X1   g286(.A1(new_n486), .A2(new_n487), .ZN(new_n488));
  AOI21_X1  g287(.A(new_n485), .B1(new_n488), .B2(KEYINPUT21), .ZN(new_n489));
  XNOR2_X1  g288(.A(new_n472), .B(new_n489), .ZN(new_n490));
  XNOR2_X1  g289(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n491));
  XNOR2_X1  g290(.A(new_n491), .B(new_n290), .ZN(new_n492));
  XOR2_X1   g291(.A(G183gat), .B(G211gat), .Z(new_n493));
  XNOR2_X1  g292(.A(new_n492), .B(new_n493), .ZN(new_n494));
  INV_X1    g293(.A(new_n494), .ZN(new_n495));
  XNOR2_X1  g294(.A(new_n490), .B(new_n495), .ZN(new_n496));
  XNOR2_X1  g295(.A(G134gat), .B(G162gat), .ZN(new_n497));
  AOI21_X1  g296(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n498));
  XOR2_X1   g297(.A(new_n497), .B(new_n498), .Z(new_n499));
  INV_X1    g298(.A(new_n499), .ZN(new_n500));
  XNOR2_X1  g299(.A(G43gat), .B(G50gat), .ZN(new_n501));
  AND2_X1   g300(.A1(new_n501), .A2(KEYINPUT15), .ZN(new_n502));
  INV_X1    g301(.A(G36gat), .ZN(new_n503));
  INV_X1    g302(.A(G29gat), .ZN(new_n504));
  NAND2_X1  g303(.A1(new_n504), .A2(KEYINPUT88), .ZN(new_n505));
  INV_X1    g304(.A(KEYINPUT88), .ZN(new_n506));
  NAND2_X1  g305(.A1(new_n506), .A2(G29gat), .ZN(new_n507));
  AOI21_X1  g306(.A(new_n503), .B1(new_n505), .B2(new_n507), .ZN(new_n508));
  NAND3_X1  g307(.A1(new_n504), .A2(new_n503), .A3(KEYINPUT14), .ZN(new_n509));
  INV_X1    g308(.A(KEYINPUT14), .ZN(new_n510));
  OAI21_X1  g309(.A(new_n510), .B1(G29gat), .B2(G36gat), .ZN(new_n511));
  NAND2_X1  g310(.A1(new_n509), .A2(new_n511), .ZN(new_n512));
  NOR2_X1   g311(.A1(new_n508), .A2(new_n512), .ZN(new_n513));
  INV_X1    g312(.A(G50gat), .ZN(new_n514));
  NAND2_X1  g313(.A1(new_n514), .A2(G43gat), .ZN(new_n515));
  INV_X1    g314(.A(G43gat), .ZN(new_n516));
  NAND2_X1  g315(.A1(new_n516), .A2(G50gat), .ZN(new_n517));
  INV_X1    g316(.A(KEYINPUT89), .ZN(new_n518));
  NAND3_X1  g317(.A1(new_n515), .A2(new_n517), .A3(new_n518), .ZN(new_n519));
  INV_X1    g318(.A(KEYINPUT15), .ZN(new_n520));
  NAND3_X1  g319(.A1(new_n516), .A2(KEYINPUT89), .A3(G50gat), .ZN(new_n521));
  NAND3_X1  g320(.A1(new_n519), .A2(new_n520), .A3(new_n521), .ZN(new_n522));
  AOI21_X1  g321(.A(new_n502), .B1(new_n513), .B2(new_n522), .ZN(new_n523));
  XNOR2_X1  g322(.A(KEYINPUT88), .B(G29gat), .ZN(new_n524));
  OAI211_X1 g323(.A(new_n511), .B(new_n509), .C1(new_n524), .C2(new_n503), .ZN(new_n525));
  NAND2_X1  g324(.A1(new_n501), .A2(KEYINPUT15), .ZN(new_n526));
  NOR2_X1   g325(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  OAI21_X1  g326(.A(KEYINPUT17), .B1(new_n523), .B2(new_n527), .ZN(new_n528));
  NAND2_X1  g327(.A1(new_n521), .A2(new_n520), .ZN(new_n529));
  AOI21_X1  g328(.A(new_n529), .B1(new_n518), .B2(new_n501), .ZN(new_n530));
  OAI21_X1  g329(.A(new_n526), .B1(new_n530), .B2(new_n525), .ZN(new_n531));
  INV_X1    g330(.A(KEYINPUT17), .ZN(new_n532));
  NAND2_X1  g331(.A1(new_n513), .A2(new_n502), .ZN(new_n533));
  NAND3_X1  g332(.A1(new_n531), .A2(new_n532), .A3(new_n533), .ZN(new_n534));
  INV_X1    g333(.A(G85gat), .ZN(new_n535));
  NAND2_X1  g334(.A1(new_n535), .A2(KEYINPUT94), .ZN(new_n536));
  INV_X1    g335(.A(KEYINPUT94), .ZN(new_n537));
  NAND2_X1  g336(.A1(new_n537), .A2(G85gat), .ZN(new_n538));
  INV_X1    g337(.A(G92gat), .ZN(new_n539));
  NAND3_X1  g338(.A1(new_n536), .A2(new_n538), .A3(new_n539), .ZN(new_n540));
  NAND2_X1  g339(.A1(G85gat), .A2(G92gat), .ZN(new_n541));
  NAND2_X1  g340(.A1(new_n541), .A2(KEYINPUT7), .ZN(new_n542));
  INV_X1    g341(.A(KEYINPUT7), .ZN(new_n543));
  NAND3_X1  g342(.A1(new_n543), .A2(G85gat), .A3(G92gat), .ZN(new_n544));
  NAND2_X1  g343(.A1(new_n542), .A2(new_n544), .ZN(new_n545));
  NAND2_X1  g344(.A1(G99gat), .A2(G106gat), .ZN(new_n546));
  NAND2_X1  g345(.A1(new_n546), .A2(KEYINPUT8), .ZN(new_n547));
  NAND3_X1  g346(.A1(new_n540), .A2(new_n545), .A3(new_n547), .ZN(new_n548));
  XNOR2_X1  g347(.A(G99gat), .B(G106gat), .ZN(new_n549));
  INV_X1    g348(.A(new_n549), .ZN(new_n550));
  NAND2_X1  g349(.A1(new_n548), .A2(new_n550), .ZN(new_n551));
  NAND4_X1  g350(.A1(new_n540), .A2(new_n545), .A3(new_n549), .A4(new_n547), .ZN(new_n552));
  NAND2_X1  g351(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  NAND3_X1  g352(.A1(new_n528), .A2(new_n534), .A3(new_n553), .ZN(new_n554));
  AND3_X1   g353(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n555));
  NOR2_X1   g354(.A1(new_n523), .A2(new_n527), .ZN(new_n556));
  INV_X1    g355(.A(KEYINPUT8), .ZN(new_n557));
  AOI21_X1  g356(.A(new_n557), .B1(G99gat), .B2(G106gat), .ZN(new_n558));
  XNOR2_X1  g357(.A(KEYINPUT94), .B(G85gat), .ZN(new_n559));
  AOI21_X1  g358(.A(new_n558), .B1(new_n559), .B2(new_n539), .ZN(new_n560));
  AOI21_X1  g359(.A(new_n549), .B1(new_n560), .B2(new_n545), .ZN(new_n561));
  INV_X1    g360(.A(new_n552), .ZN(new_n562));
  NOR2_X1   g361(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  AOI21_X1  g362(.A(new_n555), .B1(new_n556), .B2(new_n563), .ZN(new_n564));
  AND2_X1   g363(.A1(new_n554), .A2(new_n564), .ZN(new_n565));
  XNOR2_X1  g364(.A(G190gat), .B(G218gat), .ZN(new_n566));
  XNOR2_X1  g365(.A(new_n566), .B(KEYINPUT95), .ZN(new_n567));
  NAND2_X1  g366(.A1(new_n565), .A2(new_n567), .ZN(new_n568));
  NOR2_X1   g367(.A1(new_n565), .A2(new_n567), .ZN(new_n569));
  OAI211_X1 g368(.A(new_n500), .B(new_n568), .C1(new_n569), .C2(KEYINPUT97), .ZN(new_n570));
  AND2_X1   g369(.A1(new_n569), .A2(KEYINPUT97), .ZN(new_n571));
  NOR2_X1   g370(.A1(new_n570), .A2(new_n571), .ZN(new_n572));
  INV_X1    g371(.A(new_n569), .ZN(new_n573));
  INV_X1    g372(.A(KEYINPUT96), .ZN(new_n574));
  AOI21_X1  g373(.A(new_n568), .B1(new_n573), .B2(new_n574), .ZN(new_n575));
  NOR2_X1   g374(.A1(new_n575), .A2(new_n500), .ZN(new_n576));
  NAND3_X1  g375(.A1(new_n573), .A2(new_n574), .A3(new_n568), .ZN(new_n577));
  AOI21_X1  g376(.A(new_n572), .B1(new_n576), .B2(new_n577), .ZN(new_n578));
  XNOR2_X1  g377(.A(G120gat), .B(G148gat), .ZN(new_n579));
  INV_X1    g378(.A(KEYINPUT99), .ZN(new_n580));
  XNOR2_X1  g379(.A(new_n579), .B(new_n580), .ZN(new_n581));
  XNOR2_X1  g380(.A(new_n581), .B(KEYINPUT100), .ZN(new_n582));
  XNOR2_X1  g381(.A(G176gat), .B(G204gat), .ZN(new_n583));
  NAND2_X1  g382(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  INV_X1    g383(.A(KEYINPUT100), .ZN(new_n585));
  XNOR2_X1  g384(.A(new_n581), .B(new_n585), .ZN(new_n586));
  INV_X1    g385(.A(new_n583), .ZN(new_n587));
  NAND2_X1  g386(.A1(new_n586), .A2(new_n587), .ZN(new_n588));
  AND2_X1   g387(.A1(new_n584), .A2(new_n588), .ZN(new_n589));
  NAND2_X1  g388(.A1(new_n553), .A2(new_n488), .ZN(new_n590));
  NAND3_X1  g389(.A1(new_n466), .A2(new_n552), .A3(new_n551), .ZN(new_n591));
  NAND2_X1  g390(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  NAND2_X1  g391(.A1(G230gat), .A2(G233gat), .ZN(new_n593));
  NOR2_X1   g392(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  INV_X1    g393(.A(new_n594), .ZN(new_n595));
  INV_X1    g394(.A(KEYINPUT10), .ZN(new_n596));
  AND3_X1   g395(.A1(new_n460), .A2(KEYINPUT10), .A3(new_n465), .ZN(new_n597));
  INV_X1    g396(.A(KEYINPUT98), .ZN(new_n598));
  NAND3_X1  g397(.A1(new_n563), .A2(new_n597), .A3(new_n598), .ZN(new_n599));
  NAND3_X1  g398(.A1(new_n460), .A2(KEYINPUT10), .A3(new_n465), .ZN(new_n600));
  OAI21_X1  g399(.A(KEYINPUT98), .B1(new_n553), .B2(new_n600), .ZN(new_n601));
  AOI22_X1  g400(.A1(new_n592), .A2(new_n596), .B1(new_n599), .B2(new_n601), .ZN(new_n602));
  INV_X1    g401(.A(new_n593), .ZN(new_n603));
  OAI211_X1 g402(.A(new_n589), .B(new_n595), .C1(new_n602), .C2(new_n603), .ZN(new_n604));
  NAND2_X1  g403(.A1(new_n604), .A2(KEYINPUT101), .ZN(new_n605));
  NOR2_X1   g404(.A1(new_n553), .A2(new_n488), .ZN(new_n606));
  AOI21_X1  g405(.A(new_n466), .B1(new_n552), .B2(new_n551), .ZN(new_n607));
  OAI21_X1  g406(.A(new_n596), .B1(new_n606), .B2(new_n607), .ZN(new_n608));
  NAND2_X1  g407(.A1(new_n599), .A2(new_n601), .ZN(new_n609));
  NAND2_X1  g408(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  NAND2_X1  g409(.A1(new_n610), .A2(new_n593), .ZN(new_n611));
  INV_X1    g410(.A(KEYINPUT101), .ZN(new_n612));
  NAND4_X1  g411(.A1(new_n611), .A2(new_n612), .A3(new_n595), .A4(new_n589), .ZN(new_n613));
  AOI21_X1  g412(.A(new_n594), .B1(new_n610), .B2(new_n593), .ZN(new_n614));
  INV_X1    g413(.A(new_n614), .ZN(new_n615));
  NAND2_X1  g414(.A1(new_n584), .A2(new_n588), .ZN(new_n616));
  AOI22_X1  g415(.A1(new_n605), .A2(new_n613), .B1(new_n615), .B2(new_n616), .ZN(new_n617));
  NAND3_X1  g416(.A1(new_n496), .A2(new_n578), .A3(new_n617), .ZN(new_n618));
  XOR2_X1   g417(.A(new_n618), .B(KEYINPUT102), .Z(new_n619));
  INV_X1    g418(.A(new_n485), .ZN(new_n620));
  NAND3_X1  g419(.A1(new_n528), .A2(new_n534), .A3(new_n620), .ZN(new_n621));
  NAND2_X1  g420(.A1(G229gat), .A2(G233gat), .ZN(new_n622));
  XOR2_X1   g421(.A(new_n622), .B(KEYINPUT90), .Z(new_n623));
  AOI21_X1  g422(.A(KEYINPUT91), .B1(new_n556), .B2(new_n485), .ZN(new_n624));
  AND4_X1   g423(.A1(KEYINPUT91), .A2(new_n531), .A3(new_n485), .A4(new_n533), .ZN(new_n625));
  OAI211_X1 g424(.A(new_n621), .B(new_n623), .C1(new_n624), .C2(new_n625), .ZN(new_n626));
  NAND2_X1  g425(.A1(new_n626), .A2(KEYINPUT92), .ZN(new_n627));
  NAND2_X1  g426(.A1(new_n627), .A2(KEYINPUT18), .ZN(new_n628));
  INV_X1    g427(.A(KEYINPUT18), .ZN(new_n629));
  NAND3_X1  g428(.A1(new_n626), .A2(KEYINPUT92), .A3(new_n629), .ZN(new_n630));
  OAI22_X1  g429(.A1(new_n624), .A2(new_n625), .B1(new_n556), .B2(new_n485), .ZN(new_n631));
  XOR2_X1   g430(.A(new_n623), .B(KEYINPUT13), .Z(new_n632));
  NAND2_X1  g431(.A1(new_n631), .A2(new_n632), .ZN(new_n633));
  NAND3_X1  g432(.A1(new_n628), .A2(new_n630), .A3(new_n633), .ZN(new_n634));
  XNOR2_X1  g433(.A(G113gat), .B(G141gat), .ZN(new_n635));
  XNOR2_X1  g434(.A(KEYINPUT87), .B(KEYINPUT11), .ZN(new_n636));
  XNOR2_X1  g435(.A(new_n635), .B(new_n636), .ZN(new_n637));
  XNOR2_X1  g436(.A(G169gat), .B(G197gat), .ZN(new_n638));
  XNOR2_X1  g437(.A(new_n637), .B(new_n638), .ZN(new_n639));
  XNOR2_X1  g438(.A(new_n639), .B(KEYINPUT12), .ZN(new_n640));
  INV_X1    g439(.A(new_n640), .ZN(new_n641));
  NAND2_X1  g440(.A1(new_n634), .A2(new_n641), .ZN(new_n642));
  NAND4_X1  g441(.A1(new_n628), .A2(new_n630), .A3(new_n633), .A4(new_n640), .ZN(new_n643));
  NAND2_X1  g442(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  INV_X1    g443(.A(new_n644), .ZN(new_n645));
  NOR2_X1   g444(.A1(new_n619), .A2(new_n645), .ZN(new_n646));
  AND2_X1   g445(.A1(new_n449), .A2(new_n646), .ZN(new_n647));
  INV_X1    g446(.A(new_n347), .ZN(new_n648));
  NAND2_X1  g447(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  XNOR2_X1  g448(.A(new_n649), .B(G1gat), .ZN(G1324gat));
  OR2_X1    g449(.A1(KEYINPUT16), .A2(G8gat), .ZN(new_n651));
  NAND2_X1  g450(.A1(KEYINPUT16), .A2(G8gat), .ZN(new_n652));
  NAND4_X1  g451(.A1(new_n647), .A2(new_n435), .A3(new_n651), .A4(new_n652), .ZN(new_n653));
  NAND2_X1  g452(.A1(new_n653), .A2(KEYINPUT103), .ZN(new_n654));
  OR2_X1    g453(.A1(new_n654), .A2(KEYINPUT42), .ZN(new_n655));
  NAND2_X1  g454(.A1(new_n654), .A2(KEYINPUT42), .ZN(new_n656));
  AND2_X1   g455(.A1(new_n647), .A2(new_n435), .ZN(new_n657));
  OAI211_X1 g456(.A(new_n655), .B(new_n656), .C1(new_n482), .C2(new_n657), .ZN(G1325gat));
  NAND3_X1  g457(.A1(new_n647), .A2(new_n275), .A3(new_n270), .ZN(new_n659));
  NAND2_X1  g458(.A1(new_n281), .A2(G15gat), .ZN(new_n660));
  XOR2_X1   g459(.A(new_n660), .B(KEYINPUT104), .Z(new_n661));
  AOI22_X1  g460(.A1(new_n659), .A2(new_n475), .B1(new_n647), .B2(new_n661), .ZN(G1326gat));
  NAND2_X1  g461(.A1(new_n647), .A2(new_n412), .ZN(new_n663));
  XNOR2_X1  g462(.A(KEYINPUT43), .B(G22gat), .ZN(new_n664));
  XNOR2_X1  g463(.A(new_n663), .B(new_n664), .ZN(G1327gat));
  INV_X1    g464(.A(new_n578), .ZN(new_n666));
  AND2_X1   g465(.A1(new_n449), .A2(new_n666), .ZN(new_n667));
  AOI21_X1  g466(.A(new_n612), .B1(new_n614), .B2(new_n589), .ZN(new_n668));
  AOI21_X1  g467(.A(new_n603), .B1(new_n608), .B2(new_n609), .ZN(new_n669));
  NOR4_X1   g468(.A1(new_n669), .A2(KEYINPUT101), .A3(new_n616), .A4(new_n594), .ZN(new_n670));
  OAI22_X1  g469(.A1(new_n668), .A2(new_n670), .B1(new_n614), .B2(new_n589), .ZN(new_n671));
  NOR3_X1   g470(.A1(new_n496), .A2(new_n645), .A3(new_n671), .ZN(new_n672));
  AND2_X1   g471(.A1(new_n667), .A2(new_n672), .ZN(new_n673));
  NAND3_X1  g472(.A1(new_n673), .A2(new_n648), .A3(new_n524), .ZN(new_n674));
  XNOR2_X1  g473(.A(new_n674), .B(KEYINPUT45), .ZN(new_n675));
  INV_X1    g474(.A(KEYINPUT105), .ZN(new_n676));
  NAND3_X1  g475(.A1(new_n449), .A2(new_n676), .A3(new_n666), .ZN(new_n677));
  INV_X1    g476(.A(KEYINPUT44), .ZN(new_n678));
  NAND2_X1  g477(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  NAND4_X1  g478(.A1(new_n449), .A2(new_n676), .A3(KEYINPUT44), .A4(new_n666), .ZN(new_n680));
  NAND3_X1  g479(.A1(new_n679), .A2(new_n680), .A3(new_n672), .ZN(new_n681));
  NOR2_X1   g480(.A1(new_n681), .A2(new_n347), .ZN(new_n682));
  OAI21_X1  g481(.A(new_n675), .B1(new_n524), .B2(new_n682), .ZN(G1328gat));
  NAND3_X1  g482(.A1(new_n673), .A2(new_n503), .A3(new_n435), .ZN(new_n684));
  XOR2_X1   g483(.A(new_n684), .B(KEYINPUT46), .Z(new_n685));
  OAI21_X1  g484(.A(G36gat), .B1(new_n681), .B2(new_n380), .ZN(new_n686));
  NAND2_X1  g485(.A1(new_n685), .A2(new_n686), .ZN(G1329gat));
  INV_X1    g486(.A(new_n281), .ZN(new_n688));
  OAI21_X1  g487(.A(G43gat), .B1(new_n681), .B2(new_n688), .ZN(new_n689));
  NOR2_X1   g488(.A1(KEYINPUT106), .A2(KEYINPUT47), .ZN(new_n690));
  NOR2_X1   g489(.A1(new_n279), .A2(G43gat), .ZN(new_n691));
  AOI21_X1  g490(.A(new_n690), .B1(new_n673), .B2(new_n691), .ZN(new_n692));
  NAND2_X1  g491(.A1(new_n689), .A2(new_n692), .ZN(new_n693));
  NAND2_X1  g492(.A1(KEYINPUT106), .A2(KEYINPUT47), .ZN(new_n694));
  XNOR2_X1  g493(.A(new_n693), .B(new_n694), .ZN(G1330gat));
  NAND4_X1  g494(.A1(new_n679), .A2(new_n412), .A3(new_n680), .A4(new_n672), .ZN(new_n696));
  AND2_X1   g495(.A1(new_n696), .A2(KEYINPUT107), .ZN(new_n697));
  NOR2_X1   g496(.A1(new_n696), .A2(KEYINPUT107), .ZN(new_n698));
  NOR3_X1   g497(.A1(new_n697), .A2(new_n698), .A3(new_n514), .ZN(new_n699));
  NAND3_X1  g498(.A1(new_n673), .A2(new_n514), .A3(new_n412), .ZN(new_n700));
  NAND2_X1  g499(.A1(new_n700), .A2(KEYINPUT48), .ZN(new_n701));
  NAND2_X1  g500(.A1(new_n696), .A2(G50gat), .ZN(new_n702));
  AND2_X1   g501(.A1(new_n702), .A2(new_n700), .ZN(new_n703));
  OAI22_X1  g502(.A1(new_n699), .A2(new_n701), .B1(KEYINPUT48), .B2(new_n703), .ZN(G1331gat));
  INV_X1    g503(.A(new_n496), .ZN(new_n705));
  NOR4_X1   g504(.A1(new_n705), .A2(new_n666), .A3(new_n644), .A4(new_n617), .ZN(new_n706));
  NAND2_X1  g505(.A1(new_n449), .A2(new_n706), .ZN(new_n707));
  NOR2_X1   g506(.A1(new_n707), .A2(new_n347), .ZN(new_n708));
  XNOR2_X1  g507(.A(KEYINPUT108), .B(G57gat), .ZN(new_n709));
  XNOR2_X1  g508(.A(new_n708), .B(new_n709), .ZN(G1332gat));
  NOR2_X1   g509(.A1(new_n707), .A2(new_n380), .ZN(new_n711));
  NOR2_X1   g510(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n712));
  AND2_X1   g511(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n713));
  OAI21_X1  g512(.A(new_n711), .B1(new_n712), .B2(new_n713), .ZN(new_n714));
  OAI21_X1  g513(.A(new_n714), .B1(new_n711), .B2(new_n712), .ZN(G1333gat));
  NOR3_X1   g514(.A1(new_n707), .A2(G71gat), .A3(new_n279), .ZN(new_n716));
  INV_X1    g515(.A(new_n707), .ZN(new_n717));
  NAND2_X1  g516(.A1(new_n717), .A2(new_n281), .ZN(new_n718));
  AOI21_X1  g517(.A(new_n716), .B1(G71gat), .B2(new_n718), .ZN(new_n719));
  XNOR2_X1  g518(.A(new_n719), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g519(.A1(new_n717), .A2(new_n412), .ZN(new_n721));
  XNOR2_X1  g520(.A(new_n721), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g521(.A1(new_n496), .A2(new_n644), .ZN(new_n723));
  XNOR2_X1  g522(.A(new_n723), .B(KEYINPUT109), .ZN(new_n724));
  NAND2_X1  g523(.A1(new_n667), .A2(new_n724), .ZN(new_n725));
  INV_X1    g524(.A(KEYINPUT51), .ZN(new_n726));
  NAND2_X1  g525(.A1(new_n725), .A2(new_n726), .ZN(new_n727));
  NAND3_X1  g526(.A1(new_n667), .A2(KEYINPUT51), .A3(new_n724), .ZN(new_n728));
  NAND2_X1  g527(.A1(new_n727), .A2(new_n728), .ZN(new_n729));
  INV_X1    g528(.A(new_n729), .ZN(new_n730));
  NAND3_X1  g529(.A1(new_n648), .A2(new_n559), .A3(new_n671), .ZN(new_n731));
  AND2_X1   g530(.A1(new_n724), .A2(new_n671), .ZN(new_n732));
  NAND3_X1  g531(.A1(new_n679), .A2(new_n680), .A3(new_n732), .ZN(new_n733));
  NOR2_X1   g532(.A1(new_n733), .A2(new_n347), .ZN(new_n734));
  OAI22_X1  g533(.A1(new_n730), .A2(new_n731), .B1(new_n559), .B2(new_n734), .ZN(G1336gat));
  NOR3_X1   g534(.A1(new_n380), .A2(G92gat), .A3(new_n617), .ZN(new_n736));
  NAND2_X1  g535(.A1(new_n729), .A2(new_n736), .ZN(new_n737));
  OAI21_X1  g536(.A(G92gat), .B1(new_n733), .B2(new_n380), .ZN(new_n738));
  NAND2_X1  g537(.A1(new_n737), .A2(new_n738), .ZN(new_n739));
  NAND2_X1  g538(.A1(new_n739), .A2(KEYINPUT52), .ZN(new_n740));
  INV_X1    g539(.A(KEYINPUT52), .ZN(new_n741));
  NAND3_X1  g540(.A1(new_n737), .A2(new_n741), .A3(new_n738), .ZN(new_n742));
  NAND2_X1  g541(.A1(new_n740), .A2(new_n742), .ZN(G1337gat));
  OAI21_X1  g542(.A(G99gat), .B1(new_n733), .B2(new_n688), .ZN(new_n744));
  OR3_X1    g543(.A1(new_n279), .A2(G99gat), .A3(new_n617), .ZN(new_n745));
  OAI21_X1  g544(.A(new_n744), .B1(new_n730), .B2(new_n745), .ZN(G1338gat));
  OR3_X1    g545(.A1(new_n427), .A2(G106gat), .A3(new_n617), .ZN(new_n747));
  XOR2_X1   g546(.A(new_n747), .B(KEYINPUT111), .Z(new_n748));
  INV_X1    g547(.A(new_n748), .ZN(new_n749));
  AOI21_X1  g548(.A(KEYINPUT53), .B1(new_n729), .B2(new_n749), .ZN(new_n750));
  NAND4_X1  g549(.A1(new_n679), .A2(new_n412), .A3(new_n680), .A4(new_n732), .ZN(new_n751));
  INV_X1    g550(.A(KEYINPUT112), .ZN(new_n752));
  NAND2_X1  g551(.A1(new_n751), .A2(new_n752), .ZN(new_n753));
  NAND2_X1  g552(.A1(new_n753), .A2(G106gat), .ZN(new_n754));
  NOR2_X1   g553(.A1(new_n751), .A2(new_n752), .ZN(new_n755));
  OAI21_X1  g554(.A(new_n750), .B1(new_n754), .B2(new_n755), .ZN(new_n756));
  INV_X1    g555(.A(KEYINPUT110), .ZN(new_n757));
  AND3_X1   g556(.A1(new_n751), .A2(new_n757), .A3(G106gat), .ZN(new_n758));
  AOI21_X1  g557(.A(new_n757), .B1(new_n751), .B2(G106gat), .ZN(new_n759));
  AOI21_X1  g558(.A(new_n748), .B1(new_n727), .B2(new_n728), .ZN(new_n760));
  NOR3_X1   g559(.A1(new_n758), .A2(new_n759), .A3(new_n760), .ZN(new_n761));
  INV_X1    g560(.A(KEYINPUT53), .ZN(new_n762));
  OAI21_X1  g561(.A(new_n756), .B1(new_n761), .B2(new_n762), .ZN(G1339gat));
  INV_X1    g562(.A(KEYINPUT54), .ZN(new_n764));
  AOI21_X1  g563(.A(new_n764), .B1(new_n610), .B2(new_n593), .ZN(new_n765));
  NAND2_X1  g564(.A1(new_n602), .A2(new_n603), .ZN(new_n766));
  NAND2_X1  g565(.A1(new_n765), .A2(new_n766), .ZN(new_n767));
  AOI21_X1  g566(.A(new_n598), .B1(new_n563), .B2(new_n597), .ZN(new_n768));
  NOR3_X1   g567(.A1(new_n553), .A2(new_n600), .A3(KEYINPUT98), .ZN(new_n769));
  NOR2_X1   g568(.A1(new_n768), .A2(new_n769), .ZN(new_n770));
  AOI21_X1  g569(.A(KEYINPUT10), .B1(new_n590), .B2(new_n591), .ZN(new_n771));
  OAI211_X1 g570(.A(new_n764), .B(new_n593), .C1(new_n770), .C2(new_n771), .ZN(new_n772));
  AND3_X1   g571(.A1(new_n772), .A2(KEYINPUT114), .A3(new_n616), .ZN(new_n773));
  AOI21_X1  g572(.A(KEYINPUT114), .B1(new_n772), .B2(new_n616), .ZN(new_n774));
  OAI21_X1  g573(.A(new_n767), .B1(new_n773), .B2(new_n774), .ZN(new_n775));
  INV_X1    g574(.A(KEYINPUT55), .ZN(new_n776));
  NAND2_X1  g575(.A1(new_n775), .A2(new_n776), .ZN(new_n777));
  AOI21_X1  g576(.A(new_n776), .B1(new_n765), .B2(new_n766), .ZN(new_n778));
  OAI21_X1  g577(.A(new_n778), .B1(new_n773), .B2(new_n774), .ZN(new_n779));
  NAND2_X1  g578(.A1(new_n605), .A2(new_n613), .ZN(new_n780));
  AND3_X1   g579(.A1(new_n779), .A2(KEYINPUT115), .A3(new_n780), .ZN(new_n781));
  AOI21_X1  g580(.A(KEYINPUT115), .B1(new_n779), .B2(new_n780), .ZN(new_n782));
  OAI211_X1 g581(.A(new_n644), .B(new_n777), .C1(new_n781), .C2(new_n782), .ZN(new_n783));
  INV_X1    g582(.A(KEYINPUT116), .ZN(new_n784));
  OR2_X1    g583(.A1(new_n624), .A2(new_n625), .ZN(new_n785));
  AOI21_X1  g584(.A(new_n623), .B1(new_n785), .B2(new_n621), .ZN(new_n786));
  NOR2_X1   g585(.A1(new_n631), .A2(new_n632), .ZN(new_n787));
  OAI21_X1  g586(.A(new_n639), .B1(new_n786), .B2(new_n787), .ZN(new_n788));
  NAND2_X1  g587(.A1(new_n643), .A2(new_n788), .ZN(new_n789));
  OAI21_X1  g588(.A(new_n784), .B1(new_n789), .B2(new_n617), .ZN(new_n790));
  NAND4_X1  g589(.A1(new_n671), .A2(KEYINPUT116), .A3(new_n643), .A4(new_n788), .ZN(new_n791));
  AND2_X1   g590(.A1(new_n790), .A2(new_n791), .ZN(new_n792));
  NAND2_X1  g591(.A1(new_n783), .A2(new_n792), .ZN(new_n793));
  INV_X1    g592(.A(KEYINPUT117), .ZN(new_n794));
  NAND2_X1  g593(.A1(new_n793), .A2(new_n794), .ZN(new_n795));
  NAND3_X1  g594(.A1(new_n783), .A2(new_n792), .A3(KEYINPUT117), .ZN(new_n796));
  NAND3_X1  g595(.A1(new_n795), .A2(new_n578), .A3(new_n796), .ZN(new_n797));
  OR2_X1    g596(.A1(new_n578), .A2(new_n789), .ZN(new_n798));
  OAI21_X1  g597(.A(new_n777), .B1(new_n781), .B2(new_n782), .ZN(new_n799));
  NOR2_X1   g598(.A1(new_n798), .A2(new_n799), .ZN(new_n800));
  INV_X1    g599(.A(new_n800), .ZN(new_n801));
  AOI21_X1  g600(.A(new_n496), .B1(new_n797), .B2(new_n801), .ZN(new_n802));
  NOR2_X1   g601(.A1(new_n618), .A2(new_n644), .ZN(new_n803));
  XNOR2_X1  g602(.A(new_n803), .B(KEYINPUT113), .ZN(new_n804));
  OAI211_X1 g603(.A(KEYINPUT118), .B(new_n427), .C1(new_n802), .C2(new_n804), .ZN(new_n805));
  INV_X1    g604(.A(new_n805), .ZN(new_n806));
  INV_X1    g605(.A(KEYINPUT113), .ZN(new_n807));
  XNOR2_X1  g606(.A(new_n803), .B(new_n807), .ZN(new_n808));
  AOI21_X1  g607(.A(new_n666), .B1(new_n793), .B2(new_n794), .ZN(new_n809));
  AOI21_X1  g608(.A(new_n800), .B1(new_n809), .B2(new_n796), .ZN(new_n810));
  OAI21_X1  g609(.A(new_n808), .B1(new_n810), .B2(new_n496), .ZN(new_n811));
  AOI21_X1  g610(.A(KEYINPUT118), .B1(new_n811), .B2(new_n427), .ZN(new_n812));
  OR2_X1    g611(.A1(new_n806), .A2(new_n812), .ZN(new_n813));
  NAND2_X1  g612(.A1(new_n648), .A2(new_n380), .ZN(new_n814));
  NOR2_X1   g613(.A1(new_n814), .A2(new_n279), .ZN(new_n815));
  NAND2_X1  g614(.A1(new_n813), .A2(new_n815), .ZN(new_n816));
  NOR3_X1   g615(.A1(new_n816), .A2(new_n229), .A3(new_n645), .ZN(new_n817));
  AND2_X1   g616(.A1(new_n811), .A2(new_n648), .ZN(new_n818));
  INV_X1    g617(.A(new_n443), .ZN(new_n819));
  NOR2_X1   g618(.A1(new_n819), .A2(new_n435), .ZN(new_n820));
  NAND2_X1  g619(.A1(new_n818), .A2(new_n820), .ZN(new_n821));
  INV_X1    g620(.A(new_n821), .ZN(new_n822));
  AOI21_X1  g621(.A(G113gat), .B1(new_n822), .B2(new_n644), .ZN(new_n823));
  NOR2_X1   g622(.A1(new_n817), .A2(new_n823), .ZN(G1340gat));
  OAI21_X1  g623(.A(G120gat), .B1(new_n816), .B2(new_n617), .ZN(new_n825));
  OR2_X1    g624(.A1(new_n617), .A2(new_n226), .ZN(new_n826));
  OAI21_X1  g625(.A(new_n825), .B1(new_n821), .B2(new_n826), .ZN(G1341gat));
  NOR3_X1   g626(.A1(new_n816), .A2(new_n471), .A3(new_n705), .ZN(new_n828));
  OAI21_X1  g627(.A(KEYINPUT119), .B1(new_n821), .B2(new_n705), .ZN(new_n829));
  NOR3_X1   g628(.A1(new_n821), .A2(KEYINPUT119), .A3(new_n705), .ZN(new_n830));
  NOR2_X1   g629(.A1(new_n830), .A2(G127gat), .ZN(new_n831));
  AOI21_X1  g630(.A(new_n828), .B1(new_n829), .B2(new_n831), .ZN(G1342gat));
  AOI21_X1  g631(.A(G134gat), .B1(KEYINPUT120), .B2(KEYINPUT56), .ZN(new_n833));
  NAND3_X1  g632(.A1(new_n822), .A2(new_n666), .A3(new_n833), .ZN(new_n834));
  NOR2_X1   g633(.A1(KEYINPUT120), .A2(KEYINPUT56), .ZN(new_n835));
  XNOR2_X1  g634(.A(new_n834), .B(new_n835), .ZN(new_n836));
  OAI21_X1  g635(.A(G134gat), .B1(new_n816), .B2(new_n578), .ZN(new_n837));
  NAND2_X1  g636(.A1(new_n836), .A2(new_n837), .ZN(G1343gat));
  NOR2_X1   g637(.A1(new_n814), .A2(new_n281), .ZN(new_n839));
  AND2_X1   g638(.A1(new_n811), .A2(new_n412), .ZN(new_n840));
  NOR2_X1   g639(.A1(new_n840), .A2(KEYINPUT57), .ZN(new_n841));
  AND2_X1   g640(.A1(new_n841), .A2(KEYINPUT121), .ZN(new_n842));
  NAND2_X1  g641(.A1(new_n644), .A2(new_n777), .ZN(new_n843));
  NAND2_X1  g642(.A1(new_n779), .A2(new_n780), .ZN(new_n844));
  OAI22_X1  g643(.A1(new_n843), .A2(new_n844), .B1(new_n617), .B2(new_n789), .ZN(new_n845));
  NAND2_X1  g644(.A1(new_n845), .A2(new_n578), .ZN(new_n846));
  AOI21_X1  g645(.A(new_n496), .B1(new_n801), .B2(new_n846), .ZN(new_n847));
  OAI211_X1 g646(.A(KEYINPUT57), .B(new_n412), .C1(new_n804), .C2(new_n847), .ZN(new_n848));
  OAI21_X1  g647(.A(new_n848), .B1(new_n841), .B2(KEYINPUT121), .ZN(new_n849));
  OAI21_X1  g648(.A(new_n839), .B1(new_n842), .B2(new_n849), .ZN(new_n850));
  OAI21_X1  g649(.A(G141gat), .B1(new_n850), .B2(new_n645), .ZN(new_n851));
  OR2_X1    g650(.A1(KEYINPUT122), .A2(KEYINPUT58), .ZN(new_n852));
  NAND4_X1  g651(.A1(new_n818), .A2(new_n412), .A3(new_n380), .A4(new_n688), .ZN(new_n853));
  NOR3_X1   g652(.A1(new_n853), .A2(G141gat), .A3(new_n645), .ZN(new_n854));
  AOI21_X1  g653(.A(new_n854), .B1(KEYINPUT122), .B2(KEYINPUT58), .ZN(new_n855));
  AND3_X1   g654(.A1(new_n851), .A2(new_n852), .A3(new_n855), .ZN(new_n856));
  AOI21_X1  g655(.A(new_n852), .B1(new_n851), .B2(new_n855), .ZN(new_n857));
  NOR2_X1   g656(.A1(new_n856), .A2(new_n857), .ZN(G1344gat));
  NOR3_X1   g657(.A1(new_n853), .A2(G148gat), .A3(new_n617), .ZN(new_n859));
  XNOR2_X1  g658(.A(new_n859), .B(KEYINPUT123), .ZN(new_n860));
  INV_X1    g659(.A(KEYINPUT59), .ZN(new_n861));
  NAND2_X1  g660(.A1(new_n861), .A2(G148gat), .ZN(new_n862));
  INV_X1    g661(.A(new_n850), .ZN(new_n863));
  AOI21_X1  g662(.A(new_n862), .B1(new_n863), .B2(new_n671), .ZN(new_n864));
  NOR2_X1   g663(.A1(new_n619), .A2(new_n644), .ZN(new_n865));
  NOR2_X1   g664(.A1(new_n865), .A2(new_n847), .ZN(new_n866));
  NOR3_X1   g665(.A1(new_n866), .A2(KEYINPUT57), .A3(new_n427), .ZN(new_n867));
  NAND2_X1  g666(.A1(new_n811), .A2(new_n412), .ZN(new_n868));
  AOI21_X1  g667(.A(new_n867), .B1(KEYINPUT57), .B2(new_n868), .ZN(new_n869));
  NAND3_X1  g668(.A1(new_n869), .A2(new_n671), .A3(new_n839), .ZN(new_n870));
  AOI21_X1  g669(.A(new_n861), .B1(new_n870), .B2(G148gat), .ZN(new_n871));
  OAI21_X1  g670(.A(new_n860), .B1(new_n864), .B2(new_n871), .ZN(G1345gat));
  OAI21_X1  g671(.A(G155gat), .B1(new_n850), .B2(new_n705), .ZN(new_n873));
  INV_X1    g672(.A(new_n853), .ZN(new_n874));
  NAND3_X1  g673(.A1(new_n874), .A2(new_n290), .A3(new_n496), .ZN(new_n875));
  NAND2_X1  g674(.A1(new_n873), .A2(new_n875), .ZN(G1346gat));
  NOR2_X1   g675(.A1(new_n578), .A2(new_n289), .ZN(new_n877));
  NAND2_X1  g676(.A1(new_n874), .A2(new_n666), .ZN(new_n878));
  AOI22_X1  g677(.A1(new_n863), .A2(new_n877), .B1(new_n289), .B2(new_n878), .ZN(G1347gat));
  AND2_X1   g678(.A1(new_n811), .A2(new_n347), .ZN(new_n880));
  NOR2_X1   g679(.A1(new_n819), .A2(new_n380), .ZN(new_n881));
  NAND2_X1  g680(.A1(new_n880), .A2(new_n881), .ZN(new_n882));
  INV_X1    g681(.A(new_n882), .ZN(new_n883));
  AOI21_X1  g682(.A(G169gat), .B1(new_n883), .B2(new_n644), .ZN(new_n884));
  NAND2_X1  g683(.A1(new_n347), .A2(new_n435), .ZN(new_n885));
  NOR2_X1   g684(.A1(new_n885), .A2(new_n279), .ZN(new_n886));
  OAI21_X1  g685(.A(new_n886), .B1(new_n806), .B2(new_n812), .ZN(new_n887));
  NAND2_X1  g686(.A1(new_n887), .A2(KEYINPUT124), .ZN(new_n888));
  INV_X1    g687(.A(KEYINPUT124), .ZN(new_n889));
  OAI211_X1 g688(.A(new_n889), .B(new_n886), .C1(new_n806), .C2(new_n812), .ZN(new_n890));
  AND2_X1   g689(.A1(new_n888), .A2(new_n890), .ZN(new_n891));
  AND2_X1   g690(.A1(new_n644), .A2(G169gat), .ZN(new_n892));
  AOI21_X1  g691(.A(new_n884), .B1(new_n891), .B2(new_n892), .ZN(G1348gat));
  NAND2_X1  g692(.A1(new_n891), .A2(new_n671), .ZN(new_n894));
  NAND2_X1  g693(.A1(new_n894), .A2(G176gat), .ZN(new_n895));
  OR2_X1    g694(.A1(new_n617), .A2(G176gat), .ZN(new_n896));
  OAI21_X1  g695(.A(new_n895), .B1(new_n882), .B2(new_n896), .ZN(G1349gat));
  AOI21_X1  g696(.A(new_n214), .B1(new_n891), .B2(new_n496), .ZN(new_n898));
  INV_X1    g697(.A(KEYINPUT125), .ZN(new_n899));
  NAND2_X1  g698(.A1(new_n496), .A2(new_n202), .ZN(new_n900));
  OAI21_X1  g699(.A(new_n899), .B1(new_n882), .B2(new_n900), .ZN(new_n901));
  OR3_X1    g700(.A1(new_n898), .A2(KEYINPUT60), .A3(new_n901), .ZN(new_n902));
  OAI21_X1  g701(.A(KEYINPUT60), .B1(new_n898), .B2(new_n901), .ZN(new_n903));
  NAND2_X1  g702(.A1(new_n902), .A2(new_n903), .ZN(G1350gat));
  NAND3_X1  g703(.A1(new_n883), .A2(new_n203), .A3(new_n666), .ZN(new_n905));
  NAND3_X1  g704(.A1(new_n888), .A2(new_n666), .A3(new_n890), .ZN(new_n906));
  INV_X1    g705(.A(KEYINPUT61), .ZN(new_n907));
  AND3_X1   g706(.A1(new_n906), .A2(new_n907), .A3(G190gat), .ZN(new_n908));
  AOI21_X1  g707(.A(new_n907), .B1(new_n906), .B2(G190gat), .ZN(new_n909));
  OAI21_X1  g708(.A(new_n905), .B1(new_n908), .B2(new_n909), .ZN(new_n910));
  NAND2_X1  g709(.A1(new_n910), .A2(KEYINPUT126), .ZN(new_n911));
  INV_X1    g710(.A(KEYINPUT126), .ZN(new_n912));
  OAI211_X1 g711(.A(new_n912), .B(new_n905), .C1(new_n908), .C2(new_n909), .ZN(new_n913));
  NAND2_X1  g712(.A1(new_n911), .A2(new_n913), .ZN(G1351gat));
  NOR3_X1   g713(.A1(new_n427), .A2(new_n281), .A3(new_n380), .ZN(new_n915));
  NAND2_X1  g714(.A1(new_n880), .A2(new_n915), .ZN(new_n916));
  INV_X1    g715(.A(new_n916), .ZN(new_n917));
  AOI21_X1  g716(.A(G197gat), .B1(new_n917), .B2(new_n644), .ZN(new_n918));
  NOR2_X1   g717(.A1(new_n885), .A2(new_n281), .ZN(new_n919));
  NAND2_X1  g718(.A1(new_n869), .A2(new_n919), .ZN(new_n920));
  INV_X1    g719(.A(new_n920), .ZN(new_n921));
  AND2_X1   g720(.A1(new_n644), .A2(G197gat), .ZN(new_n922));
  AOI21_X1  g721(.A(new_n918), .B1(new_n921), .B2(new_n922), .ZN(G1352gat));
  NOR3_X1   g722(.A1(new_n916), .A2(G204gat), .A3(new_n617), .ZN(new_n924));
  XNOR2_X1  g723(.A(KEYINPUT127), .B(KEYINPUT62), .ZN(new_n925));
  XNOR2_X1  g724(.A(new_n924), .B(new_n925), .ZN(new_n926));
  OAI21_X1  g725(.A(G204gat), .B1(new_n920), .B2(new_n617), .ZN(new_n927));
  NAND2_X1  g726(.A1(new_n926), .A2(new_n927), .ZN(G1353gat));
  NAND3_X1  g727(.A1(new_n917), .A2(new_n357), .A3(new_n496), .ZN(new_n929));
  NAND2_X1  g728(.A1(new_n921), .A2(new_n496), .ZN(new_n930));
  AND3_X1   g729(.A1(new_n930), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n931));
  AOI21_X1  g730(.A(KEYINPUT63), .B1(new_n930), .B2(G211gat), .ZN(new_n932));
  OAI21_X1  g731(.A(new_n929), .B1(new_n931), .B2(new_n932), .ZN(G1354gat));
  OAI21_X1  g732(.A(G218gat), .B1(new_n920), .B2(new_n578), .ZN(new_n934));
  NAND3_X1  g733(.A1(new_n917), .A2(new_n358), .A3(new_n666), .ZN(new_n935));
  NAND2_X1  g734(.A1(new_n934), .A2(new_n935), .ZN(G1355gat));
endmodule


