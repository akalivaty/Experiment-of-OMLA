

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368,
         n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379,
         n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390,
         n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
         n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412,
         n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423,
         n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
         n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445,
         n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456,
         n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467,
         n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478,
         n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489,
         n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500,
         n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511,
         n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588,
         n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599,
         n600, n601, n602, n603, n604, n605, n606, n607, n608, n609, n610,
         n611, n612, n613, n614, n615, n616, n617, n618, n619, n620, n621,
         n622, n623, n624, n625, n626, n627, n628, n629, n630, n631, n632,
         n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, n643,
         n644, n645, n646, n647, n648, n649, n650, n651, n652, n653, n654,
         n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, n665,
         n666, n667, n668, n669, n670, n671, n672, n673, n674, n675, n676,
         n677, n678, n679, n680, n681, n682, n683, n684, n685, n686, n687,
         n688, n689, n690, n691, n692, n693, n694, n695, n696, n697, n698,
         n699, n700, n701, n702, n703, n704, n705, n706, n707, n708, n709,
         n710, n711, n712, n713, n714, n715, n716, n717, n718, n719, n720,
         n721, n722, n723, n724, n725, n726, n727, n728, n729, n730, n731,
         n732, n733, n734, n735, n736, n737, n738, n739, n740, n741, n742,
         n743, n744, n745, n746, n747, n748, n749, n750, n751, n752, n753,
         n754, n755, n756, n757, n758, n759, n760, n761, n762, n763, n764,
         n765, n766, n767, n768, n769, n770, n771, n772, n773, n774, n775,
         n776, n777, n778, n779, n780, n781, n782, n783, n784, n785, n786,
         n787, n788, n789, n790, n791, n792, n793, n794, n795, n796, n797,
         n798, n799, n800, n801, n802, n803, n804, n805, n806, n807;

  NAND2_X1 U381 ( .A1(n391), .A2(n390), .ZN(n384) );
  AND2_X1 U382 ( .A1(n413), .A2(n805), .ZN(n381) );
  BUF_X1 U383 ( .A(n386), .Z(n593) );
  AND2_X1 U384 ( .A1(n424), .A2(n427), .ZN(n372) );
  XNOR2_X2 U385 ( .A(G143), .B(G128), .ZN(n462) );
  XNOR2_X2 U386 ( .A(n388), .B(KEYINPUT31), .ZN(n724) );
  XNOR2_X1 U387 ( .A(G143), .B(G128), .ZN(n362) );
  NOR2_X1 U388 ( .A1(n603), .A2(n590), .ZN(n592) );
  BUF_X1 U389 ( .A(G128), .Z(n364) );
  XOR2_X1 U390 ( .A(n361), .B(n394), .Z(n358) );
  XNOR2_X2 U391 ( .A(n545), .B(n544), .ZN(n602) );
  INV_X4 U392 ( .A(G953), .ZN(n801) );
  XNOR2_X2 U393 ( .A(KEYINPUT64), .B(KEYINPUT79), .ZN(n461) );
  NOR2_X1 U394 ( .A1(n441), .A2(n440), .ZN(n439) );
  INV_X1 U395 ( .A(n381), .ZN(n360) );
  INV_X1 U396 ( .A(n737), .ZN(n359) );
  AND2_X2 U397 ( .A1(n454), .A2(n668), .ZN(n798) );
  XNOR2_X1 U398 ( .A(n439), .B(KEYINPUT48), .ZN(n454) );
  XNOR2_X1 U399 ( .A(n651), .B(n650), .ZN(n441) );
  NAND2_X1 U400 ( .A1(n403), .A2(n402), .ZN(n401) );
  AND2_X1 U401 ( .A1(n407), .A2(n405), .ZN(n404) );
  AND2_X1 U402 ( .A1(n387), .A2(n741), .ZN(n711) );
  XNOR2_X1 U403 ( .A(KEYINPUT41), .B(n646), .ZN(n750) );
  NAND2_X1 U404 ( .A1(n420), .A2(n428), .ZN(n417) );
  XNOR2_X1 U405 ( .A(n521), .B(n520), .ZN(n606) );
  AND2_X1 U406 ( .A1(n429), .A2(KEYINPUT19), .ZN(n420) );
  XNOR2_X1 U407 ( .A(n675), .B(KEYINPUT62), .ZN(n676) );
  XNOR2_X1 U408 ( .A(n500), .B(n516), .ZN(n793) );
  NAND2_X1 U409 ( .A1(n414), .A2(n590), .ZN(n361) );
  NAND2_X1 U410 ( .A1(n414), .A2(n590), .ZN(n583) );
  XNOR2_X1 U411 ( .A(n583), .B(n394), .ZN(n393) );
  XNOR2_X1 U412 ( .A(KEYINPUT64), .B(KEYINPUT79), .ZN(n363) );
  NAND2_X1 U413 ( .A1(n446), .A2(n448), .ZN(n365) );
  NAND2_X1 U414 ( .A1(n446), .A2(n448), .ZN(n771) );
  BUF_X1 U415 ( .A(n672), .Z(n784) );
  NAND2_X1 U416 ( .A1(n426), .A2(n371), .ZN(n425) );
  NAND2_X1 U417 ( .A1(n452), .A2(n451), .ZN(n421) );
  NAND2_X1 U418 ( .A1(n567), .A2(n669), .ZN(n451) );
  INV_X1 U419 ( .A(n563), .ZN(n669) );
  XNOR2_X1 U420 ( .A(KEYINPUT16), .B(G122), .ZN(n559) );
  OR2_X1 U421 ( .A1(n776), .A2(G902), .ZN(n400) );
  INV_X1 U422 ( .A(KEYINPUT25), .ZN(n460) );
  XNOR2_X1 U423 ( .A(n566), .B(n565), .ZN(n567) );
  XNOR2_X1 U424 ( .A(KEYINPUT92), .B(KEYINPUT15), .ZN(n480) );
  AND2_X1 U425 ( .A1(n798), .A2(n671), .ZN(n465) );
  OR2_X1 U426 ( .A1(n798), .A2(n469), .ZN(n468) );
  INV_X1 U427 ( .A(KEYINPUT111), .ZN(n459) );
  NAND2_X1 U428 ( .A1(n675), .A2(n543), .ZN(n418) );
  NAND2_X1 U429 ( .A1(n576), .A2(n367), .ZN(n578) );
  NAND2_X1 U430 ( .A1(n415), .A2(n417), .ZN(n576) );
  XNOR2_X1 U431 ( .A(n382), .B(G134), .ZN(n516) );
  XNOR2_X1 U432 ( .A(n542), .B(n433), .ZN(n701) );
  XNOR2_X1 U433 ( .A(n557), .B(n434), .ZN(n433) );
  INV_X1 U434 ( .A(n793), .ZN(n542) );
  XNOR2_X1 U435 ( .A(n541), .B(G140), .ZN(n434) );
  XNOR2_X1 U436 ( .A(n562), .B(n780), .ZN(n689) );
  XNOR2_X1 U437 ( .A(n438), .B(n648), .ZN(n665) );
  INV_X1 U438 ( .A(n634), .ZN(n437) );
  XNOR2_X1 U439 ( .A(n519), .B(G478), .ZN(n520) );
  INV_X1 U440 ( .A(KEYINPUT103), .ZN(n519) );
  NOR2_X1 U441 ( .A1(n628), .A2(n581), .ZN(n409) );
  INV_X1 U442 ( .A(KEYINPUT87), .ZN(n394) );
  XNOR2_X1 U443 ( .A(n495), .B(n532), .ZN(n776) );
  XNOR2_X1 U444 ( .A(n494), .B(n493), .ZN(n495) );
  XNOR2_X1 U445 ( .A(n399), .B(n395), .ZN(n494) );
  NAND2_X1 U446 ( .A1(n450), .A2(n563), .ZN(n449) );
  XNOR2_X1 U447 ( .A(n432), .B(n431), .ZN(n538) );
  XNOR2_X1 U448 ( .A(G104), .B(G107), .ZN(n432) );
  XNOR2_X1 U449 ( .A(G101), .B(G110), .ZN(n431) );
  XNOR2_X1 U450 ( .A(n621), .B(KEYINPUT45), .ZN(n672) );
  XNOR2_X1 U451 ( .A(G125), .B(G140), .ZN(n484) );
  XNOR2_X1 U452 ( .A(G122), .B(KEYINPUT12), .ZN(n524) );
  XOR2_X1 U453 ( .A(KEYINPUT102), .B(KEYINPUT11), .Z(n525) );
  XNOR2_X1 U454 ( .A(G131), .B(G143), .ZN(n522) );
  XOR2_X1 U455 ( .A(G104), .B(G113), .Z(n523) );
  NAND2_X1 U456 ( .A1(n467), .A2(n671), .ZN(n466) );
  XNOR2_X1 U457 ( .A(KEYINPUT18), .B(G125), .ZN(n553) );
  NAND2_X1 U458 ( .A1(n455), .A2(n374), .ZN(n440) );
  AND2_X1 U459 ( .A1(n659), .A2(n369), .ZN(n455) );
  NOR2_X1 U460 ( .A1(n633), .A2(n436), .ZN(n435) );
  NAND2_X1 U461 ( .A1(n645), .A2(KEYINPUT19), .ZN(n427) );
  XNOR2_X1 U462 ( .A(n602), .B(n546), .ZN(n589) );
  XNOR2_X1 U463 ( .A(n550), .B(n422), .ZN(n499) );
  INV_X1 U464 ( .A(G137), .ZN(n422) );
  XNOR2_X1 U465 ( .A(KEYINPUT93), .B(KEYINPUT3), .ZN(n506) );
  INV_X1 U466 ( .A(n538), .ZN(n779) );
  XNOR2_X1 U467 ( .A(n397), .B(n396), .ZN(n395) );
  XNOR2_X1 U468 ( .A(KEYINPUT23), .B(KEYINPUT24), .ZN(n396) );
  XNOR2_X1 U469 ( .A(n398), .B(G119), .ZN(n397) );
  INV_X1 U470 ( .A(G110), .ZN(n398) );
  XNOR2_X1 U471 ( .A(n486), .B(n485), .ZN(n399) );
  XNOR2_X1 U472 ( .A(n364), .B(G137), .ZN(n486) );
  XNOR2_X1 U473 ( .A(KEYINPUT76), .B(KEYINPUT72), .ZN(n485) );
  AND2_X1 U474 ( .A1(n457), .A2(n456), .ZN(n653) );
  NOR2_X1 U475 ( .A1(n741), .A2(n639), .ZN(n640) );
  OR2_X1 U476 ( .A1(n584), .A2(n406), .ZN(n405) );
  BUF_X1 U477 ( .A(n589), .Z(n743) );
  INV_X1 U478 ( .A(KEYINPUT22), .ZN(n463) );
  XNOR2_X1 U479 ( .A(n516), .B(n471), .ZN(n517) );
  XOR2_X1 U480 ( .A(G116), .B(G107), .Z(n471) );
  XNOR2_X1 U481 ( .A(n683), .B(n682), .ZN(n684) );
  XNOR2_X1 U482 ( .A(n701), .B(n700), .ZN(n702) );
  XNOR2_X1 U483 ( .A(n690), .B(n693), .ZN(n694) );
  NOR2_X1 U484 ( .A1(n665), .A2(n709), .ZN(n649) );
  INV_X1 U485 ( .A(KEYINPUT35), .ZN(n419) );
  NAND2_X1 U486 ( .A1(n598), .A2(n597), .ZN(n599) );
  NOR2_X1 U487 ( .A1(n409), .A2(n359), .ZN(n408) );
  XNOR2_X1 U488 ( .A(n777), .B(n776), .ZN(n430) );
  XNOR2_X1 U489 ( .A(n443), .B(n442), .ZN(G75) );
  XNOR2_X1 U490 ( .A(KEYINPUT53), .B(KEYINPUT117), .ZN(n442) );
  OR2_X1 U491 ( .A1(n769), .A2(n444), .ZN(n443) );
  NAND2_X1 U492 ( .A1(n368), .A2(n770), .ZN(n444) );
  AND2_X1 U493 ( .A1(n389), .A2(n379), .ZN(n366) );
  XNOR2_X1 U494 ( .A(n511), .B(KEYINPUT94), .ZN(n754) );
  OR2_X1 U495 ( .A1(n575), .A2(n574), .ZN(n367) );
  OR2_X1 U496 ( .A1(n768), .A2(n767), .ZN(n368) );
  OR2_X1 U497 ( .A1(n664), .A2(n663), .ZN(n369) );
  OR2_X1 U498 ( .A1(n634), .A2(n633), .ZN(n370) );
  AND2_X1 U499 ( .A1(n754), .A2(n570), .ZN(n371) );
  AND2_X1 U500 ( .A1(n468), .A2(n466), .ZN(n373) );
  AND2_X1 U501 ( .A1(n637), .A2(n717), .ZN(n374) );
  BUF_X1 U502 ( .A(n602), .Z(n642) );
  XOR2_X1 U503 ( .A(n472), .B(n460), .Z(n375) );
  AND2_X1 U504 ( .A1(n628), .A2(n581), .ZN(n376) );
  NOR2_X1 U505 ( .A1(n743), .A2(n586), .ZN(n377) );
  AND2_X1 U506 ( .A1(n456), .A2(n742), .ZN(n378) );
  INV_X2 U507 ( .A(G146), .ZN(n423) );
  XNOR2_X1 U508 ( .A(n518), .B(n517), .ZN(n772) );
  AND2_X1 U509 ( .A1(n600), .A2(KEYINPUT44), .ZN(n379) );
  NAND2_X1 U510 ( .A1(n670), .A2(KEYINPUT65), .ZN(n469) );
  AND2_X1 U511 ( .A1(n415), .A2(n417), .ZN(n380) );
  XNOR2_X1 U512 ( .A(n638), .B(KEYINPUT6), .ZN(n590) );
  XNOR2_X1 U513 ( .A(n793), .B(n509), .ZN(n675) );
  AND2_X1 U514 ( .A1(n738), .A2(n737), .ZN(n742) );
  XNOR2_X1 U515 ( .A(n362), .B(n363), .ZN(n382) );
  XNOR2_X1 U516 ( .A(n462), .B(n461), .ZN(n551) );
  INV_X1 U517 ( .A(n755), .ZN(n436) );
  XNOR2_X1 U518 ( .A(n383), .B(KEYINPUT101), .ZN(n608) );
  NOR2_X2 U519 ( .A1(n724), .A2(n711), .ZN(n383) );
  BUF_X1 U520 ( .A(n413), .Z(n385) );
  NAND2_X1 U521 ( .A1(n404), .A2(n401), .ZN(n413) );
  XNOR2_X1 U522 ( .A(n453), .B(KEYINPUT99), .ZN(n387) );
  NAND2_X1 U523 ( .A1(n583), .A2(n585), .ZN(n407) );
  NAND2_X1 U524 ( .A1(n360), .A2(n366), .ZN(n410) );
  XNOR2_X1 U525 ( .A(n578), .B(n577), .ZN(n386) );
  XNOR2_X1 U526 ( .A(n578), .B(n577), .ZN(n601) );
  NAND2_X1 U527 ( .A1(n593), .A2(n748), .ZN(n388) );
  NAND2_X1 U528 ( .A1(n381), .A2(n389), .ZN(n615) );
  XNOR2_X1 U529 ( .A(n389), .B(G122), .ZN(G24) );
  XNOR2_X2 U530 ( .A(n599), .B(n419), .ZN(n389) );
  NAND2_X1 U531 ( .A1(n358), .A2(n376), .ZN(n390) );
  AND2_X2 U532 ( .A1(n392), .A2(n408), .ZN(n391) );
  NAND2_X1 U533 ( .A1(n393), .A2(KEYINPUT88), .ZN(n392) );
  XNOR2_X2 U534 ( .A(n400), .B(n375), .ZN(n737) );
  AND2_X1 U535 ( .A1(n584), .A2(n406), .ZN(n402) );
  INV_X1 U536 ( .A(n361), .ZN(n403) );
  INV_X1 U537 ( .A(n585), .ZN(n406) );
  NAND2_X1 U538 ( .A1(n411), .A2(n410), .ZN(n613) );
  NAND2_X1 U539 ( .A1(n412), .A2(KEYINPUT66), .ZN(n411) );
  NAND2_X1 U540 ( .A1(n615), .A2(KEYINPUT44), .ZN(n412) );
  XNOR2_X1 U541 ( .A(n385), .B(n708), .ZN(G21) );
  NAND2_X1 U542 ( .A1(n414), .A2(n377), .ZN(n588) );
  XNOR2_X2 U543 ( .A(n580), .B(n463), .ZN(n414) );
  NAND2_X1 U544 ( .A1(n672), .A2(n669), .ZN(n623) );
  AND2_X2 U545 ( .A1(n416), .A2(n372), .ZN(n415) );
  NAND2_X1 U546 ( .A1(n421), .A2(n371), .ZN(n416) );
  XNOR2_X2 U547 ( .A(n418), .B(G472), .ZN(n638) );
  NAND2_X1 U548 ( .A1(n589), .A2(n742), .ZN(n603) );
  INV_X1 U549 ( .A(n421), .ZN(n428) );
  XNOR2_X2 U550 ( .A(n423), .B(KEYINPUT4), .ZN(n550) );
  OR2_X1 U551 ( .A1(n689), .A2(n449), .ZN(n429) );
  OR2_X1 U552 ( .A1(n689), .A2(n425), .ZN(n424) );
  INV_X1 U553 ( .A(n449), .ZN(n426) );
  NAND2_X1 U554 ( .A1(n428), .A2(n429), .ZN(n644) );
  NAND2_X1 U555 ( .A1(n601), .A2(n579), .ZN(n580) );
  NOR2_X1 U556 ( .A1(n430), .A2(n778), .ZN(G66) );
  NAND2_X1 U557 ( .A1(n464), .A2(n373), .ZN(n447) );
  NAND2_X1 U558 ( .A1(n447), .A2(n674), .ZN(n446) );
  NAND2_X1 U559 ( .A1(n384), .A2(n609), .ZN(n611) );
  NAND2_X1 U560 ( .A1(n771), .A2(G469), .ZN(n703) );
  NAND2_X1 U561 ( .A1(n539), .A2(n540), .ZN(n557) );
  NAND2_X1 U562 ( .A1(n437), .A2(n435), .ZN(n438) );
  NAND2_X1 U563 ( .A1(n445), .A2(n674), .ZN(n448) );
  NOR2_X1 U564 ( .A1(n470), .A2(n469), .ZN(n445) );
  INV_X1 U565 ( .A(n567), .ZN(n450) );
  NAND2_X1 U566 ( .A1(n689), .A2(n567), .ZN(n452) );
  NAND2_X1 U567 ( .A1(n386), .A2(n378), .ZN(n453) );
  NAND2_X1 U568 ( .A1(n750), .A2(n653), .ZN(n647) );
  INV_X1 U569 ( .A(n642), .ZN(n456) );
  XNOR2_X1 U570 ( .A(n640), .B(n458), .ZN(n457) );
  XNOR2_X1 U571 ( .A(n641), .B(n459), .ZN(n458) );
  XNOR2_X2 U572 ( .A(n623), .B(n622), .ZN(n470) );
  NAND2_X1 U573 ( .A1(n470), .A2(n465), .ZN(n464) );
  INV_X1 U574 ( .A(n670), .ZN(n467) );
  BUF_X1 U575 ( .A(n771), .Z(n775) );
  AND2_X1 U576 ( .A1(G217), .A2(n496), .ZN(n472) );
  XNOR2_X1 U577 ( .A(KEYINPUT46), .B(KEYINPUT86), .ZN(n650) );
  INV_X1 U578 ( .A(KEYINPUT84), .ZN(n622) );
  INV_X1 U579 ( .A(n736), .ZN(n674) );
  INV_X1 U580 ( .A(KEYINPUT34), .ZN(n594) );
  XNOR2_X1 U581 ( .A(n595), .B(n594), .ZN(n598) );
  XOR2_X1 U582 ( .A(KEYINPUT108), .B(KEYINPUT109), .Z(n548) );
  XOR2_X1 U583 ( .A(KEYINPUT14), .B(KEYINPUT95), .Z(n474) );
  NAND2_X1 U584 ( .A1(G234), .A2(G237), .ZN(n473) );
  XNOR2_X1 U585 ( .A(n474), .B(n473), .ZN(n476) );
  NAND2_X1 U586 ( .A1(G902), .A2(n476), .ZN(n572) );
  NOR2_X1 U587 ( .A1(G900), .A2(n572), .ZN(n475) );
  NAND2_X1 U588 ( .A1(G953), .A2(n475), .ZN(n479) );
  NAND2_X1 U589 ( .A1(G952), .A2(n476), .ZN(n767) );
  NOR2_X1 U590 ( .A1(G953), .A2(n767), .ZN(n477) );
  XNOR2_X1 U591 ( .A(n477), .B(KEYINPUT96), .ZN(n575) );
  INV_X1 U592 ( .A(n575), .ZN(n478) );
  NAND2_X1 U593 ( .A1(n479), .A2(n478), .ZN(n483) );
  XNOR2_X1 U594 ( .A(n480), .B(G902), .ZN(n563) );
  NAND2_X1 U595 ( .A1(G234), .A2(n563), .ZN(n481) );
  XNOR2_X1 U596 ( .A(n481), .B(KEYINPUT20), .ZN(n496) );
  AND2_X1 U597 ( .A1(n496), .A2(G221), .ZN(n482) );
  XNOR2_X1 U598 ( .A(n482), .B(KEYINPUT21), .ZN(n738) );
  NAND2_X1 U599 ( .A1(n483), .A2(n738), .ZN(n631) );
  XNOR2_X1 U600 ( .A(n631), .B(KEYINPUT69), .ZN(n497) );
  XNOR2_X1 U601 ( .A(n484), .B(KEYINPUT10), .ZN(n792) );
  XNOR2_X1 U602 ( .A(n792), .B(n423), .ZN(n532) );
  INV_X1 U603 ( .A(KEYINPUT8), .ZN(n487) );
  NAND2_X1 U604 ( .A1(n487), .A2(KEYINPUT82), .ZN(n490) );
  INV_X1 U605 ( .A(KEYINPUT82), .ZN(n488) );
  NAND2_X1 U606 ( .A1(n488), .A2(KEYINPUT8), .ZN(n489) );
  NAND2_X1 U607 ( .A1(n490), .A2(n489), .ZN(n492) );
  NAND2_X1 U608 ( .A1(G234), .A2(n801), .ZN(n491) );
  XNOR2_X1 U609 ( .A(n492), .B(n491), .ZN(n512) );
  NAND2_X1 U610 ( .A1(G221), .A2(n512), .ZN(n493) );
  NAND2_X1 U611 ( .A1(n497), .A2(n359), .ZN(n498) );
  XNOR2_X1 U612 ( .A(n498), .B(KEYINPUT68), .ZN(n639) );
  XNOR2_X1 U613 ( .A(n499), .B(G131), .ZN(n500) );
  XNOR2_X1 U614 ( .A(G101), .B(KEYINPUT5), .ZN(n501) );
  XNOR2_X1 U615 ( .A(n501), .B(KEYINPUT100), .ZN(n503) );
  NOR2_X1 U616 ( .A1(G953), .A2(G237), .ZN(n528) );
  NAND2_X1 U617 ( .A1(n528), .A2(G210), .ZN(n502) );
  XNOR2_X1 U618 ( .A(n503), .B(n502), .ZN(n508) );
  XNOR2_X1 U619 ( .A(G119), .B(G116), .ZN(n505) );
  XNOR2_X1 U620 ( .A(G113), .B(KEYINPUT71), .ZN(n504) );
  XNOR2_X1 U621 ( .A(n505), .B(n504), .ZN(n507) );
  XNOR2_X1 U622 ( .A(n507), .B(n506), .ZN(n561) );
  XNOR2_X1 U623 ( .A(n508), .B(n561), .ZN(n509) );
  INV_X1 U624 ( .A(G902), .ZN(n543) );
  NOR2_X1 U625 ( .A1(n639), .A2(n590), .ZN(n536) );
  NOR2_X1 U626 ( .A1(G902), .A2(G237), .ZN(n510) );
  XNOR2_X1 U627 ( .A(n510), .B(KEYINPUT75), .ZN(n564) );
  NAND2_X1 U628 ( .A1(n564), .A2(G214), .ZN(n511) );
  INV_X1 U629 ( .A(n754), .ZN(n645) );
  NAND2_X1 U630 ( .A1(G217), .A2(n512), .ZN(n514) );
  XOR2_X1 U631 ( .A(G122), .B(KEYINPUT9), .Z(n513) );
  XNOR2_X1 U632 ( .A(n514), .B(n513), .ZN(n515) );
  XOR2_X1 U633 ( .A(n515), .B(KEYINPUT7), .Z(n518) );
  NOR2_X1 U634 ( .A1(n772), .A2(G902), .ZN(n521) );
  XNOR2_X1 U635 ( .A(n523), .B(n522), .ZN(n527) );
  XNOR2_X1 U636 ( .A(n525), .B(n524), .ZN(n526) );
  XOR2_X1 U637 ( .A(n527), .B(n526), .Z(n530) );
  NAND2_X1 U638 ( .A1(G214), .A2(n528), .ZN(n529) );
  XNOR2_X1 U639 ( .A(n530), .B(n529), .ZN(n531) );
  XNOR2_X1 U640 ( .A(n532), .B(n531), .ZN(n683) );
  NAND2_X1 U641 ( .A1(n683), .A2(n543), .ZN(n534) );
  XOR2_X1 U642 ( .A(KEYINPUT13), .B(G475), .Z(n533) );
  XNOR2_X1 U643 ( .A(n534), .B(n533), .ZN(n605) );
  NAND2_X1 U644 ( .A1(n606), .A2(n605), .ZN(n709) );
  NOR2_X1 U645 ( .A1(n645), .A2(n709), .ZN(n535) );
  NAND2_X1 U646 ( .A1(n536), .A2(n535), .ZN(n625) );
  NAND2_X1 U647 ( .A1(n779), .A2(KEYINPUT73), .ZN(n540) );
  INV_X1 U648 ( .A(KEYINPUT73), .ZN(n537) );
  NAND2_X1 U649 ( .A1(n538), .A2(n537), .ZN(n539) );
  NAND2_X1 U650 ( .A1(G227), .A2(n801), .ZN(n541) );
  NAND2_X1 U651 ( .A1(n701), .A2(n543), .ZN(n545) );
  XOR2_X1 U652 ( .A(KEYINPUT70), .B(G469), .Z(n544) );
  INV_X1 U653 ( .A(KEYINPUT1), .ZN(n546) );
  OR2_X1 U654 ( .A1(n625), .A2(n743), .ZN(n547) );
  XNOR2_X1 U655 ( .A(n548), .B(n547), .ZN(n549) );
  XNOR2_X1 U656 ( .A(KEYINPUT43), .B(n549), .ZN(n568) );
  XNOR2_X1 U657 ( .A(n551), .B(n550), .ZN(n556) );
  NAND2_X1 U658 ( .A1(n801), .A2(G224), .ZN(n552) );
  XNOR2_X1 U659 ( .A(n552), .B(KEYINPUT17), .ZN(n554) );
  XNOR2_X1 U660 ( .A(n554), .B(n553), .ZN(n555) );
  XNOR2_X1 U661 ( .A(n556), .B(n555), .ZN(n558) );
  XNOR2_X1 U662 ( .A(n558), .B(n557), .ZN(n562) );
  XNOR2_X1 U663 ( .A(n559), .B(KEYINPUT74), .ZN(n560) );
  XNOR2_X1 U664 ( .A(n561), .B(n560), .ZN(n780) );
  NAND2_X1 U665 ( .A1(n564), .A2(G210), .ZN(n566) );
  INV_X1 U666 ( .A(KEYINPUT80), .ZN(n565) );
  INV_X1 U667 ( .A(n644), .ZN(n624) );
  AND2_X1 U668 ( .A1(n568), .A2(n624), .ZN(n667) );
  XOR2_X1 U669 ( .A(n667), .B(G140), .Z(G42) );
  INV_X1 U670 ( .A(n605), .ZN(n569) );
  AND2_X1 U671 ( .A1(n606), .A2(n569), .ZN(n757) );
  AND2_X1 U672 ( .A1(n757), .A2(n738), .ZN(n579) );
  INV_X1 U673 ( .A(KEYINPUT19), .ZN(n570) );
  NOR2_X1 U674 ( .A1(G898), .A2(n801), .ZN(n571) );
  XNOR2_X1 U675 ( .A(KEYINPUT97), .B(n571), .ZN(n781) );
  NOR2_X1 U676 ( .A1(n572), .A2(n781), .ZN(n573) );
  XNOR2_X1 U677 ( .A(n573), .B(KEYINPUT98), .ZN(n574) );
  INV_X1 U678 ( .A(KEYINPUT0), .ZN(n577) );
  INV_X1 U679 ( .A(n743), .ZN(n628) );
  INV_X1 U680 ( .A(KEYINPUT88), .ZN(n581) );
  XNOR2_X1 U681 ( .A(G101), .B(KEYINPUT112), .ZN(n582) );
  XNOR2_X1 U682 ( .A(n384), .B(n582), .ZN(G3) );
  AND2_X1 U683 ( .A1(n743), .A2(n359), .ZN(n584) );
  XNOR2_X1 U684 ( .A(KEYINPUT78), .B(KEYINPUT32), .ZN(n585) );
  OR2_X1 U685 ( .A1(n638), .A2(n737), .ZN(n586) );
  INV_X1 U686 ( .A(KEYINPUT107), .ZN(n587) );
  XNOR2_X1 U687 ( .A(n588), .B(n587), .ZN(n805) );
  INV_X1 U688 ( .A(KEYINPUT33), .ZN(n591) );
  XNOR2_X1 U689 ( .A(n592), .B(n591), .ZN(n730) );
  NAND2_X1 U690 ( .A1(n730), .A2(n593), .ZN(n595) );
  INV_X1 U691 ( .A(n606), .ZN(n596) );
  NAND2_X1 U692 ( .A1(n596), .A2(n605), .ZN(n635) );
  XNOR2_X1 U693 ( .A(n635), .B(KEYINPUT77), .ZN(n597) );
  INV_X1 U694 ( .A(KEYINPUT66), .ZN(n600) );
  INV_X1 U695 ( .A(n603), .ZN(n604) );
  AND2_X1 U696 ( .A1(n638), .A2(n604), .ZN(n748) );
  NOR2_X1 U697 ( .A1(n606), .A2(n605), .ZN(n607) );
  XNOR2_X1 U698 ( .A(n607), .B(KEYINPUT104), .ZN(n725) );
  XNOR2_X1 U699 ( .A(KEYINPUT105), .B(n725), .ZN(n666) );
  NAND2_X1 U700 ( .A1(n666), .A2(n709), .ZN(n753) );
  NAND2_X1 U701 ( .A1(n608), .A2(n753), .ZN(n609) );
  INV_X1 U702 ( .A(KEYINPUT106), .ZN(n610) );
  XNOR2_X1 U703 ( .A(n611), .B(n610), .ZN(n612) );
  NAND2_X1 U704 ( .A1(n612), .A2(n613), .ZN(n614) );
  XNOR2_X1 U705 ( .A(n614), .B(KEYINPUT89), .ZN(n620) );
  BUF_X1 U706 ( .A(n615), .Z(n616) );
  INV_X1 U707 ( .A(n616), .ZN(n618) );
  INV_X1 U708 ( .A(KEYINPUT44), .ZN(n617) );
  NAND2_X1 U709 ( .A1(n618), .A2(n617), .ZN(n619) );
  NAND2_X1 U710 ( .A1(n620), .A2(n619), .ZN(n621) );
  NOR2_X1 U711 ( .A1(n625), .A2(n624), .ZN(n626) );
  XOR2_X1 U712 ( .A(KEYINPUT36), .B(n626), .Z(n627) );
  NOR2_X1 U713 ( .A1(n628), .A2(n627), .ZN(n727) );
  INV_X1 U714 ( .A(KEYINPUT47), .ZN(n660) );
  AND2_X1 U715 ( .A1(n660), .A2(KEYINPUT81), .ZN(n629) );
  NOR2_X1 U716 ( .A1(n727), .A2(n629), .ZN(n637) );
  NAND2_X1 U717 ( .A1(n638), .A2(n754), .ZN(n630) );
  XNOR2_X1 U718 ( .A(n630), .B(KEYINPUT30), .ZN(n634) );
  NOR2_X1 U719 ( .A1(n642), .A2(n631), .ZN(n632) );
  NAND2_X1 U720 ( .A1(n632), .A2(n737), .ZN(n633) );
  NOR2_X1 U721 ( .A1(n370), .A2(n635), .ZN(n636) );
  NAND2_X1 U722 ( .A1(n636), .A2(n644), .ZN(n717) );
  XNOR2_X1 U723 ( .A(KEYINPUT28), .B(KEYINPUT110), .ZN(n641) );
  INV_X1 U724 ( .A(n638), .ZN(n741) );
  INV_X1 U725 ( .A(KEYINPUT38), .ZN(n643) );
  XNOR2_X1 U726 ( .A(n644), .B(n643), .ZN(n755) );
  NOR2_X1 U727 ( .A1(n436), .A2(n645), .ZN(n752) );
  NAND2_X1 U728 ( .A1(n752), .A2(n757), .ZN(n646) );
  XNOR2_X1 U729 ( .A(KEYINPUT42), .B(n647), .ZN(n806) );
  INV_X1 U730 ( .A(KEYINPUT39), .ZN(n648) );
  XOR2_X1 U731 ( .A(KEYINPUT40), .B(n649), .Z(n807) );
  NAND2_X1 U732 ( .A1(n806), .A2(n807), .ZN(n651) );
  INV_X1 U733 ( .A(n380), .ZN(n652) );
  NAND2_X1 U734 ( .A1(n653), .A2(n652), .ZN(n663) );
  INV_X1 U735 ( .A(n663), .ZN(n718) );
  NAND2_X1 U736 ( .A1(n718), .A2(KEYINPUT67), .ZN(n657) );
  INV_X1 U737 ( .A(n753), .ZN(n655) );
  NOR2_X1 U738 ( .A1(n718), .A2(KEYINPUT81), .ZN(n654) );
  NOR2_X1 U739 ( .A1(n655), .A2(n654), .ZN(n656) );
  NAND2_X1 U740 ( .A1(n657), .A2(n656), .ZN(n658) );
  NAND2_X1 U741 ( .A1(n658), .A2(KEYINPUT47), .ZN(n659) );
  NAND2_X1 U742 ( .A1(n753), .A2(n660), .ZN(n661) );
  NOR2_X1 U743 ( .A1(KEYINPUT67), .A2(n661), .ZN(n662) );
  NOR2_X1 U744 ( .A1(n662), .A2(KEYINPUT81), .ZN(n664) );
  NOR2_X1 U745 ( .A1(n666), .A2(n665), .ZN(n729) );
  NOR2_X1 U746 ( .A1(n667), .A2(n729), .ZN(n668) );
  NAND2_X1 U747 ( .A1(n669), .A2(KEYINPUT2), .ZN(n670) );
  INV_X1 U748 ( .A(KEYINPUT65), .ZN(n671) );
  AND2_X1 U749 ( .A1(n798), .A2(KEYINPUT2), .ZN(n673) );
  AND2_X1 U750 ( .A1(n784), .A2(n673), .ZN(n736) );
  NAND2_X1 U751 ( .A1(n771), .A2(G472), .ZN(n677) );
  XNOR2_X1 U752 ( .A(n677), .B(n676), .ZN(n680) );
  INV_X1 U753 ( .A(G952), .ZN(n678) );
  NAND2_X1 U754 ( .A1(n678), .A2(G953), .ZN(n679) );
  XNOR2_X1 U755 ( .A(n679), .B(KEYINPUT91), .ZN(n778) );
  INV_X1 U756 ( .A(n778), .ZN(n704) );
  NAND2_X1 U757 ( .A1(n680), .A2(n704), .ZN(n681) );
  XNOR2_X1 U758 ( .A(n681), .B(KEYINPUT63), .ZN(G57) );
  NAND2_X1 U759 ( .A1(n365), .A2(G475), .ZN(n685) );
  XNOR2_X1 U760 ( .A(KEYINPUT121), .B(KEYINPUT59), .ZN(n682) );
  XNOR2_X1 U761 ( .A(n685), .B(n684), .ZN(n686) );
  NAND2_X1 U762 ( .A1(n686), .A2(n704), .ZN(n688) );
  INV_X1 U763 ( .A(KEYINPUT60), .ZN(n687) );
  XNOR2_X1 U764 ( .A(n688), .B(n687), .ZN(G60) );
  NAND2_X1 U765 ( .A1(n365), .A2(G210), .ZN(n695) );
  BUF_X1 U766 ( .A(n689), .Z(n690) );
  XOR2_X1 U767 ( .A(KEYINPUT55), .B(KEYINPUT90), .Z(n692) );
  XNOR2_X1 U768 ( .A(KEYINPUT54), .B(KEYINPUT118), .ZN(n691) );
  XOR2_X1 U769 ( .A(n692), .B(n691), .Z(n693) );
  XNOR2_X1 U770 ( .A(n695), .B(n694), .ZN(n696) );
  NAND2_X1 U771 ( .A1(n696), .A2(n704), .ZN(n698) );
  XNOR2_X1 U772 ( .A(KEYINPUT85), .B(KEYINPUT56), .ZN(n697) );
  XNOR2_X1 U773 ( .A(n698), .B(n697), .ZN(G51) );
  XNOR2_X1 U774 ( .A(KEYINPUT119), .B(KEYINPUT57), .ZN(n699) );
  XNOR2_X1 U775 ( .A(n699), .B(KEYINPUT58), .ZN(n700) );
  XNOR2_X1 U776 ( .A(n703), .B(n702), .ZN(n705) );
  NAND2_X1 U777 ( .A1(n705), .A2(n704), .ZN(n707) );
  INV_X1 U778 ( .A(KEYINPUT120), .ZN(n706) );
  XNOR2_X1 U779 ( .A(n707), .B(n706), .ZN(G54) );
  XOR2_X1 U780 ( .A(G119), .B(KEYINPUT127), .Z(n708) );
  INV_X1 U781 ( .A(n709), .ZN(n722) );
  NAND2_X1 U782 ( .A1(n711), .A2(n722), .ZN(n710) );
  XNOR2_X1 U783 ( .A(n710), .B(G104), .ZN(G6) );
  XOR2_X1 U784 ( .A(KEYINPUT27), .B(KEYINPUT26), .Z(n713) );
  NAND2_X1 U785 ( .A1(n711), .A2(n725), .ZN(n712) );
  XNOR2_X1 U786 ( .A(n713), .B(n712), .ZN(n714) );
  XNOR2_X1 U787 ( .A(G107), .B(n714), .ZN(G9) );
  XOR2_X1 U788 ( .A(n364), .B(KEYINPUT29), .Z(n716) );
  NAND2_X1 U789 ( .A1(n718), .A2(n725), .ZN(n715) );
  XNOR2_X1 U790 ( .A(n716), .B(n715), .ZN(G30) );
  XNOR2_X1 U791 ( .A(G143), .B(n717), .ZN(G45) );
  XOR2_X1 U792 ( .A(KEYINPUT113), .B(KEYINPUT114), .Z(n720) );
  NAND2_X1 U793 ( .A1(n718), .A2(n722), .ZN(n719) );
  XNOR2_X1 U794 ( .A(n720), .B(n719), .ZN(n721) );
  XNOR2_X1 U795 ( .A(G146), .B(n721), .ZN(G48) );
  NAND2_X1 U796 ( .A1(n724), .A2(n722), .ZN(n723) );
  XNOR2_X1 U797 ( .A(n723), .B(G113), .ZN(G15) );
  NAND2_X1 U798 ( .A1(n725), .A2(n724), .ZN(n726) );
  XNOR2_X1 U799 ( .A(n726), .B(G116), .ZN(G18) );
  XNOR2_X1 U800 ( .A(G125), .B(n727), .ZN(n728) );
  XNOR2_X1 U801 ( .A(n728), .B(KEYINPUT37), .ZN(G27) );
  XOR2_X1 U802 ( .A(G134), .B(n729), .Z(G36) );
  BUF_X1 U803 ( .A(n730), .Z(n761) );
  AND2_X1 U804 ( .A1(n750), .A2(n761), .ZN(n731) );
  NOR2_X1 U805 ( .A1(G953), .A2(n731), .ZN(n770) );
  NOR2_X1 U806 ( .A1(n784), .A2(KEYINPUT2), .ZN(n732) );
  XNOR2_X1 U807 ( .A(n732), .B(KEYINPUT83), .ZN(n734) );
  OR2_X1 U808 ( .A1(KEYINPUT2), .A2(n798), .ZN(n733) );
  NAND2_X1 U809 ( .A1(n734), .A2(n733), .ZN(n735) );
  NOR2_X1 U810 ( .A1(n736), .A2(n735), .ZN(n769) );
  NOR2_X1 U811 ( .A1(n738), .A2(n737), .ZN(n739) );
  XNOR2_X1 U812 ( .A(n739), .B(KEYINPUT49), .ZN(n740) );
  NAND2_X1 U813 ( .A1(n741), .A2(n740), .ZN(n746) );
  NOR2_X1 U814 ( .A1(n743), .A2(n742), .ZN(n744) );
  XNOR2_X1 U815 ( .A(n744), .B(KEYINPUT50), .ZN(n745) );
  NOR2_X1 U816 ( .A1(n746), .A2(n745), .ZN(n747) );
  NOR2_X1 U817 ( .A1(n748), .A2(n747), .ZN(n749) );
  XNOR2_X1 U818 ( .A(n749), .B(KEYINPUT51), .ZN(n751) );
  NAND2_X1 U819 ( .A1(n751), .A2(n750), .ZN(n764) );
  NAND2_X1 U820 ( .A1(n753), .A2(n752), .ZN(n760) );
  NOR2_X1 U821 ( .A1(n755), .A2(n754), .ZN(n756) );
  XNOR2_X1 U822 ( .A(KEYINPUT115), .B(n756), .ZN(n758) );
  NAND2_X1 U823 ( .A1(n758), .A2(n757), .ZN(n759) );
  NAND2_X1 U824 ( .A1(n760), .A2(n759), .ZN(n762) );
  NAND2_X1 U825 ( .A1(n762), .A2(n761), .ZN(n763) );
  NAND2_X1 U826 ( .A1(n764), .A2(n763), .ZN(n766) );
  XOR2_X1 U827 ( .A(KEYINPUT52), .B(KEYINPUT116), .Z(n765) );
  XNOR2_X1 U828 ( .A(n766), .B(n765), .ZN(n768) );
  NAND2_X1 U829 ( .A1(n775), .A2(G478), .ZN(n773) );
  XNOR2_X1 U830 ( .A(n773), .B(n772), .ZN(n774) );
  NOR2_X1 U831 ( .A1(n774), .A2(n778), .ZN(G63) );
  NAND2_X1 U832 ( .A1(n775), .A2(G217), .ZN(n777) );
  XNOR2_X1 U833 ( .A(n780), .B(n779), .ZN(n782) );
  NAND2_X1 U834 ( .A1(n782), .A2(n781), .ZN(n783) );
  XNOR2_X1 U835 ( .A(n783), .B(KEYINPUT123), .ZN(n791) );
  NAND2_X1 U836 ( .A1(n784), .A2(n801), .ZN(n789) );
  NAND2_X1 U837 ( .A1(G224), .A2(G953), .ZN(n785) );
  XNOR2_X1 U838 ( .A(n785), .B(KEYINPUT61), .ZN(n786) );
  XNOR2_X1 U839 ( .A(KEYINPUT122), .B(n786), .ZN(n787) );
  NAND2_X1 U840 ( .A1(G898), .A2(n787), .ZN(n788) );
  NAND2_X1 U841 ( .A1(n789), .A2(n788), .ZN(n790) );
  XNOR2_X1 U842 ( .A(n791), .B(n790), .ZN(G69) );
  XNOR2_X1 U843 ( .A(n793), .B(n792), .ZN(n794) );
  XNOR2_X1 U844 ( .A(n794), .B(KEYINPUT124), .ZN(n799) );
  XNOR2_X1 U845 ( .A(G227), .B(n799), .ZN(n795) );
  XNOR2_X1 U846 ( .A(n795), .B(KEYINPUT126), .ZN(n796) );
  NAND2_X1 U847 ( .A1(G900), .A2(n796), .ZN(n797) );
  NAND2_X1 U848 ( .A1(n797), .A2(G953), .ZN(n804) );
  XNOR2_X1 U849 ( .A(n799), .B(n798), .ZN(n800) );
  XNOR2_X1 U850 ( .A(n800), .B(KEYINPUT125), .ZN(n802) );
  NAND2_X1 U851 ( .A1(n802), .A2(n801), .ZN(n803) );
  NAND2_X1 U852 ( .A1(n804), .A2(n803), .ZN(G72) );
  XNOR2_X1 U853 ( .A(G110), .B(n805), .ZN(G12) );
  XNOR2_X1 U854 ( .A(G137), .B(n806), .ZN(G39) );
  XNOR2_X1 U855 ( .A(G131), .B(n807), .ZN(G33) );
endmodule

