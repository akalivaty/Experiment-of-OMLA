//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 1 0 1 0 1 1 0 0 1 1 1 1 0 0 0 0 0 0 1 1 1 1 1 1 1 0 0 1 0 0 1 0 1 1 1 0 1 0 1 1 1 1 1 0 0 1 1 1 0 0 1 0 1 0 0 0 0 0 0 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:18:44 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n679, new_n680, new_n681, new_n682, new_n683, new_n684, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n692, new_n693, new_n694,
    new_n695, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n719, new_n720, new_n721, new_n722, new_n723, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n759, new_n760, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n768, new_n769, new_n770, new_n772,
    new_n774, new_n775, new_n776, new_n777, new_n778, new_n779, new_n780,
    new_n781, new_n782, new_n783, new_n784, new_n785, new_n787, new_n788,
    new_n789, new_n790, new_n792, new_n793, new_n794, new_n795, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n857, new_n858, new_n860, new_n861, new_n863, new_n864,
    new_n865, new_n866, new_n867, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n907, new_n908, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n919,
    new_n920, new_n921, new_n923, new_n924, new_n925, new_n926, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n939, new_n940, new_n941, new_n942,
    new_n944, new_n945, new_n946, new_n947, new_n948, new_n949, new_n950,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n966,
    new_n967, new_n968, new_n969, new_n970, new_n972, new_n973, new_n974,
    new_n975, new_n976;
  XOR2_X1   g000(.A(KEYINPUT74), .B(G197gat), .Z(new_n202));
  NAND2_X1  g001(.A1(new_n202), .A2(G204gat), .ZN(new_n203));
  XNOR2_X1  g002(.A(KEYINPUT74), .B(G197gat), .ZN(new_n204));
  INV_X1    g003(.A(G204gat), .ZN(new_n205));
  NAND2_X1  g004(.A1(new_n204), .A2(new_n205), .ZN(new_n206));
  INV_X1    g005(.A(KEYINPUT22), .ZN(new_n207));
  INV_X1    g006(.A(G218gat), .ZN(new_n208));
  AND2_X1   g007(.A1(new_n208), .A2(KEYINPUT75), .ZN(new_n209));
  NOR2_X1   g008(.A1(new_n208), .A2(KEYINPUT75), .ZN(new_n210));
  OAI21_X1  g009(.A(new_n207), .B1(new_n209), .B2(new_n210), .ZN(new_n211));
  NAND3_X1  g010(.A1(new_n203), .A2(new_n206), .A3(new_n211), .ZN(new_n212));
  NAND2_X1  g011(.A1(new_n212), .A2(G211gat), .ZN(new_n213));
  NOR2_X1   g012(.A1(new_n207), .A2(G211gat), .ZN(new_n214));
  NAND3_X1  g013(.A1(new_n203), .A2(new_n206), .A3(new_n214), .ZN(new_n215));
  NAND2_X1  g014(.A1(new_n213), .A2(new_n215), .ZN(new_n216));
  NAND2_X1  g015(.A1(new_n216), .A2(G218gat), .ZN(new_n217));
  NAND3_X1  g016(.A1(new_n213), .A2(new_n215), .A3(new_n208), .ZN(new_n218));
  NAND2_X1  g017(.A1(new_n217), .A2(new_n218), .ZN(new_n219));
  INV_X1    g018(.A(G226gat), .ZN(new_n220));
  INV_X1    g019(.A(G233gat), .ZN(new_n221));
  NOR2_X1   g020(.A1(new_n220), .A2(new_n221), .ZN(new_n222));
  INV_X1    g021(.A(KEYINPUT23), .ZN(new_n223));
  AND2_X1   g022(.A1(new_n223), .A2(KEYINPUT65), .ZN(new_n224));
  NOR2_X1   g023(.A1(new_n223), .A2(KEYINPUT65), .ZN(new_n225));
  OAI22_X1  g024(.A1(new_n224), .A2(new_n225), .B1(G169gat), .B2(G176gat), .ZN(new_n226));
  INV_X1    g025(.A(KEYINPUT24), .ZN(new_n227));
  INV_X1    g026(.A(G183gat), .ZN(new_n228));
  INV_X1    g027(.A(G190gat), .ZN(new_n229));
  OAI21_X1  g028(.A(new_n227), .B1(new_n228), .B2(new_n229), .ZN(new_n230));
  NAND2_X1  g029(.A1(new_n228), .A2(new_n229), .ZN(new_n231));
  NAND3_X1  g030(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n232));
  NAND3_X1  g031(.A1(new_n230), .A2(new_n231), .A3(new_n232), .ZN(new_n233));
  NAND2_X1  g032(.A1(G169gat), .A2(G176gat), .ZN(new_n234));
  INV_X1    g033(.A(new_n234), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n223), .A2(KEYINPUT65), .ZN(new_n236));
  NOR2_X1   g035(.A1(G169gat), .A2(G176gat), .ZN(new_n237));
  AOI21_X1  g036(.A(new_n235), .B1(new_n236), .B2(new_n237), .ZN(new_n238));
  NAND3_X1  g037(.A1(new_n226), .A2(new_n233), .A3(new_n238), .ZN(new_n239));
  INV_X1    g038(.A(KEYINPUT25), .ZN(new_n240));
  NAND2_X1  g039(.A1(new_n239), .A2(new_n240), .ZN(new_n241));
  NAND4_X1  g040(.A1(new_n226), .A2(new_n233), .A3(new_n238), .A4(KEYINPUT25), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n241), .A2(new_n242), .ZN(new_n243));
  AND2_X1   g042(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n244));
  NOR2_X1   g043(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n245));
  OAI21_X1  g044(.A(new_n229), .B1(new_n244), .B2(new_n245), .ZN(new_n246));
  AND2_X1   g045(.A1(KEYINPUT66), .A2(KEYINPUT28), .ZN(new_n247));
  NOR2_X1   g046(.A1(KEYINPUT66), .A2(KEYINPUT28), .ZN(new_n248));
  NOR2_X1   g047(.A1(new_n247), .A2(new_n248), .ZN(new_n249));
  XNOR2_X1  g048(.A(new_n246), .B(new_n249), .ZN(new_n250));
  NOR2_X1   g049(.A1(new_n228), .A2(new_n229), .ZN(new_n251));
  NOR3_X1   g050(.A1(KEYINPUT26), .A2(G169gat), .A3(G176gat), .ZN(new_n252));
  OAI21_X1  g051(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n253));
  NAND2_X1  g052(.A1(new_n253), .A2(new_n234), .ZN(new_n254));
  INV_X1    g053(.A(KEYINPUT67), .ZN(new_n255));
  AOI21_X1  g054(.A(new_n252), .B1(new_n254), .B2(new_n255), .ZN(new_n256));
  NAND3_X1  g055(.A1(new_n253), .A2(KEYINPUT67), .A3(new_n234), .ZN(new_n257));
  AOI21_X1  g056(.A(new_n251), .B1(new_n256), .B2(new_n257), .ZN(new_n258));
  INV_X1    g057(.A(KEYINPUT68), .ZN(new_n259));
  OAI21_X1  g058(.A(new_n250), .B1(new_n258), .B2(new_n259), .ZN(new_n260));
  AND3_X1   g059(.A1(new_n253), .A2(KEYINPUT67), .A3(new_n234), .ZN(new_n261));
  AOI21_X1  g060(.A(KEYINPUT67), .B1(new_n253), .B2(new_n234), .ZN(new_n262));
  NOR3_X1   g061(.A1(new_n261), .A2(new_n262), .A3(new_n252), .ZN(new_n263));
  NOR3_X1   g062(.A1(new_n263), .A2(KEYINPUT68), .A3(new_n251), .ZN(new_n264));
  OAI21_X1  g063(.A(new_n243), .B1(new_n260), .B2(new_n264), .ZN(new_n265));
  XNOR2_X1  g064(.A(KEYINPUT76), .B(KEYINPUT29), .ZN(new_n266));
  INV_X1    g065(.A(new_n266), .ZN(new_n267));
  AOI21_X1  g066(.A(new_n222), .B1(new_n265), .B2(new_n267), .ZN(new_n268));
  INV_X1    g067(.A(new_n222), .ZN(new_n269));
  OAI21_X1  g068(.A(KEYINPUT68), .B1(new_n263), .B2(new_n251), .ZN(new_n270));
  NAND2_X1  g069(.A1(new_n258), .A2(new_n259), .ZN(new_n271));
  NAND3_X1  g070(.A1(new_n270), .A2(new_n271), .A3(new_n250), .ZN(new_n272));
  AOI21_X1  g071(.A(new_n269), .B1(new_n272), .B2(new_n243), .ZN(new_n273));
  OAI21_X1  g072(.A(new_n219), .B1(new_n268), .B2(new_n273), .ZN(new_n274));
  XNOR2_X1  g073(.A(G8gat), .B(G36gat), .ZN(new_n275));
  XNOR2_X1  g074(.A(G64gat), .B(G92gat), .ZN(new_n276));
  XNOR2_X1  g075(.A(new_n275), .B(new_n276), .ZN(new_n277));
  INV_X1    g076(.A(new_n277), .ZN(new_n278));
  NAND2_X1  g077(.A1(new_n265), .A2(new_n222), .ZN(new_n279));
  AND3_X1   g078(.A1(new_n213), .A2(new_n208), .A3(new_n215), .ZN(new_n280));
  AOI21_X1  g079(.A(new_n208), .B1(new_n213), .B2(new_n215), .ZN(new_n281));
  NOR2_X1   g080(.A1(new_n280), .A2(new_n281), .ZN(new_n282));
  AOI21_X1  g081(.A(KEYINPUT29), .B1(new_n272), .B2(new_n243), .ZN(new_n283));
  OAI211_X1 g082(.A(new_n279), .B(new_n282), .C1(new_n283), .C2(new_n222), .ZN(new_n284));
  NAND3_X1  g083(.A1(new_n274), .A2(new_n278), .A3(new_n284), .ZN(new_n285));
  NAND2_X1  g084(.A1(new_n285), .A2(KEYINPUT77), .ZN(new_n286));
  INV_X1    g085(.A(KEYINPUT77), .ZN(new_n287));
  NAND4_X1  g086(.A1(new_n274), .A2(new_n287), .A3(new_n284), .A4(new_n278), .ZN(new_n288));
  NAND2_X1  g087(.A1(new_n286), .A2(new_n288), .ZN(new_n289));
  INV_X1    g088(.A(KEYINPUT30), .ZN(new_n290));
  NAND2_X1  g089(.A1(new_n289), .A2(new_n290), .ZN(new_n291));
  NAND4_X1  g090(.A1(new_n274), .A2(KEYINPUT30), .A3(new_n284), .A4(new_n278), .ZN(new_n292));
  AND2_X1   g091(.A1(new_n274), .A2(new_n284), .ZN(new_n293));
  OAI21_X1  g092(.A(new_n292), .B1(new_n293), .B2(new_n278), .ZN(new_n294));
  INV_X1    g093(.A(new_n294), .ZN(new_n295));
  XNOR2_X1  g094(.A(G1gat), .B(G29gat), .ZN(new_n296));
  XNOR2_X1  g095(.A(new_n296), .B(G85gat), .ZN(new_n297));
  XNOR2_X1  g096(.A(KEYINPUT0), .B(G57gat), .ZN(new_n298));
  XNOR2_X1  g097(.A(new_n297), .B(new_n298), .ZN(new_n299));
  INV_X1    g098(.A(new_n299), .ZN(new_n300));
  INV_X1    g099(.A(KEYINPUT5), .ZN(new_n301));
  NAND2_X1  g100(.A1(G225gat), .A2(G233gat), .ZN(new_n302));
  AND2_X1   g101(.A1(G155gat), .A2(G162gat), .ZN(new_n303));
  NOR2_X1   g102(.A1(G155gat), .A2(G162gat), .ZN(new_n304));
  NOR2_X1   g103(.A1(new_n303), .A2(new_n304), .ZN(new_n305));
  XNOR2_X1  g104(.A(G141gat), .B(G148gat), .ZN(new_n306));
  INV_X1    g105(.A(KEYINPUT2), .ZN(new_n307));
  AOI21_X1  g106(.A(new_n307), .B1(G155gat), .B2(G162gat), .ZN(new_n308));
  OAI21_X1  g107(.A(new_n305), .B1(new_n306), .B2(new_n308), .ZN(new_n309));
  INV_X1    g108(.A(G141gat), .ZN(new_n310));
  NAND2_X1  g109(.A1(new_n310), .A2(G148gat), .ZN(new_n311));
  INV_X1    g110(.A(G148gat), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n312), .A2(G141gat), .ZN(new_n313));
  NAND2_X1  g112(.A1(new_n311), .A2(new_n313), .ZN(new_n314));
  XNOR2_X1  g113(.A(G155gat), .B(G162gat), .ZN(new_n315));
  INV_X1    g114(.A(G155gat), .ZN(new_n316));
  INV_X1    g115(.A(G162gat), .ZN(new_n317));
  OAI21_X1  g116(.A(KEYINPUT2), .B1(new_n316), .B2(new_n317), .ZN(new_n318));
  NAND3_X1  g117(.A1(new_n314), .A2(new_n315), .A3(new_n318), .ZN(new_n319));
  INV_X1    g118(.A(KEYINPUT3), .ZN(new_n320));
  AND3_X1   g119(.A1(new_n309), .A2(new_n319), .A3(new_n320), .ZN(new_n321));
  AOI21_X1  g120(.A(new_n320), .B1(new_n309), .B2(new_n319), .ZN(new_n322));
  NOR2_X1   g121(.A1(new_n321), .A2(new_n322), .ZN(new_n323));
  INV_X1    g122(.A(KEYINPUT69), .ZN(new_n324));
  INV_X1    g123(.A(G134gat), .ZN(new_n325));
  NAND3_X1  g124(.A1(new_n324), .A2(new_n325), .A3(G127gat), .ZN(new_n326));
  INV_X1    g125(.A(G127gat), .ZN(new_n327));
  AOI21_X1  g126(.A(KEYINPUT69), .B1(new_n327), .B2(G134gat), .ZN(new_n328));
  NOR2_X1   g127(.A1(new_n327), .A2(G134gat), .ZN(new_n329));
  OAI21_X1  g128(.A(new_n326), .B1(new_n328), .B2(new_n329), .ZN(new_n330));
  INV_X1    g129(.A(KEYINPUT70), .ZN(new_n331));
  NAND2_X1  g130(.A1(new_n330), .A2(new_n331), .ZN(new_n332));
  OAI211_X1 g131(.A(KEYINPUT70), .B(new_n326), .C1(new_n328), .C2(new_n329), .ZN(new_n333));
  INV_X1    g132(.A(G120gat), .ZN(new_n334));
  NAND2_X1  g133(.A1(new_n334), .A2(G113gat), .ZN(new_n335));
  INV_X1    g134(.A(G113gat), .ZN(new_n336));
  NAND2_X1  g135(.A1(new_n336), .A2(G120gat), .ZN(new_n337));
  AOI21_X1  g136(.A(KEYINPUT1), .B1(new_n335), .B2(new_n337), .ZN(new_n338));
  INV_X1    g137(.A(new_n338), .ZN(new_n339));
  NAND3_X1  g138(.A1(new_n332), .A2(new_n333), .A3(new_n339), .ZN(new_n340));
  XNOR2_X1  g139(.A(G127gat), .B(G134gat), .ZN(new_n341));
  NAND2_X1  g140(.A1(new_n338), .A2(new_n341), .ZN(new_n342));
  NAND2_X1  g141(.A1(new_n340), .A2(new_n342), .ZN(new_n343));
  NAND2_X1  g142(.A1(new_n323), .A2(new_n343), .ZN(new_n344));
  AND2_X1   g143(.A1(new_n309), .A2(new_n319), .ZN(new_n345));
  NAND3_X1  g144(.A1(new_n340), .A2(new_n345), .A3(new_n342), .ZN(new_n346));
  NOR2_X1   g145(.A1(new_n346), .A2(KEYINPUT4), .ZN(new_n347));
  INV_X1    g146(.A(KEYINPUT4), .ZN(new_n348));
  AOI21_X1  g147(.A(new_n338), .B1(new_n330), .B2(new_n331), .ZN(new_n349));
  AOI22_X1  g148(.A1(new_n349), .A2(new_n333), .B1(new_n338), .B2(new_n341), .ZN(new_n350));
  AOI21_X1  g149(.A(new_n348), .B1(new_n350), .B2(new_n345), .ZN(new_n351));
  OAI211_X1 g150(.A(new_n302), .B(new_n344), .C1(new_n347), .C2(new_n351), .ZN(new_n352));
  INV_X1    g151(.A(new_n345), .ZN(new_n353));
  NAND2_X1  g152(.A1(new_n343), .A2(new_n353), .ZN(new_n354));
  AOI21_X1  g153(.A(new_n302), .B1(new_n354), .B2(new_n346), .ZN(new_n355));
  INV_X1    g154(.A(new_n355), .ZN(new_n356));
  AOI21_X1  g155(.A(new_n301), .B1(new_n352), .B2(new_n356), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n346), .A2(KEYINPUT4), .ZN(new_n358));
  NAND3_X1  g157(.A1(new_n350), .A2(new_n348), .A3(new_n345), .ZN(new_n359));
  AOI22_X1  g158(.A1(new_n358), .A2(new_n359), .B1(new_n343), .B2(new_n323), .ZN(new_n360));
  AOI21_X1  g159(.A(KEYINPUT5), .B1(new_n360), .B2(new_n302), .ZN(new_n361));
  OAI21_X1  g160(.A(new_n300), .B1(new_n357), .B2(new_n361), .ZN(new_n362));
  NAND2_X1  g161(.A1(new_n352), .A2(new_n301), .ZN(new_n363));
  AOI21_X1  g162(.A(new_n355), .B1(new_n360), .B2(new_n302), .ZN(new_n364));
  OAI211_X1 g163(.A(new_n299), .B(new_n363), .C1(new_n364), .C2(new_n301), .ZN(new_n365));
  INV_X1    g164(.A(KEYINPUT6), .ZN(new_n366));
  NAND3_X1  g165(.A1(new_n362), .A2(new_n365), .A3(new_n366), .ZN(new_n367));
  NOR2_X1   g166(.A1(new_n357), .A2(new_n361), .ZN(new_n368));
  NAND3_X1  g167(.A1(new_n368), .A2(KEYINPUT6), .A3(new_n299), .ZN(new_n369));
  NAND2_X1  g168(.A1(new_n367), .A2(new_n369), .ZN(new_n370));
  NAND3_X1  g169(.A1(new_n291), .A2(new_n295), .A3(new_n370), .ZN(new_n371));
  XNOR2_X1  g170(.A(KEYINPUT78), .B(KEYINPUT31), .ZN(new_n372));
  INV_X1    g171(.A(G50gat), .ZN(new_n373));
  XNOR2_X1  g172(.A(new_n372), .B(new_n373), .ZN(new_n374));
  XNOR2_X1  g173(.A(G78gat), .B(G106gat), .ZN(new_n375));
  INV_X1    g174(.A(G22gat), .ZN(new_n376));
  XNOR2_X1  g175(.A(new_n375), .B(new_n376), .ZN(new_n377));
  XNOR2_X1  g176(.A(new_n374), .B(new_n377), .ZN(new_n378));
  INV_X1    g177(.A(new_n378), .ZN(new_n379));
  INV_X1    g178(.A(G228gat), .ZN(new_n380));
  NOR2_X1   g179(.A1(new_n380), .A2(new_n221), .ZN(new_n381));
  INV_X1    g180(.A(new_n381), .ZN(new_n382));
  NOR3_X1   g181(.A1(new_n280), .A2(new_n281), .A3(KEYINPUT29), .ZN(new_n383));
  OAI21_X1  g182(.A(new_n353), .B1(new_n383), .B2(KEYINPUT3), .ZN(new_n384));
  NOR2_X1   g183(.A1(new_n321), .A2(new_n266), .ZN(new_n385));
  INV_X1    g184(.A(new_n385), .ZN(new_n386));
  NAND2_X1  g185(.A1(new_n219), .A2(new_n386), .ZN(new_n387));
  AOI21_X1  g186(.A(new_n382), .B1(new_n384), .B2(new_n387), .ZN(new_n388));
  NAND3_X1  g187(.A1(new_n217), .A2(new_n218), .A3(new_n267), .ZN(new_n389));
  AOI21_X1  g188(.A(new_n345), .B1(new_n389), .B2(new_n320), .ZN(new_n390));
  NOR2_X1   g189(.A1(new_n282), .A2(new_n385), .ZN(new_n391));
  NOR3_X1   g190(.A1(new_n390), .A2(new_n391), .A3(new_n381), .ZN(new_n392));
  OAI21_X1  g191(.A(new_n379), .B1(new_n388), .B2(new_n392), .ZN(new_n393));
  AOI21_X1  g192(.A(KEYINPUT3), .B1(new_n282), .B2(new_n267), .ZN(new_n394));
  OAI211_X1 g193(.A(new_n382), .B(new_n387), .C1(new_n394), .C2(new_n345), .ZN(new_n395));
  INV_X1    g194(.A(KEYINPUT29), .ZN(new_n396));
  NAND3_X1  g195(.A1(new_n217), .A2(new_n218), .A3(new_n396), .ZN(new_n397));
  AOI21_X1  g196(.A(new_n345), .B1(new_n397), .B2(new_n320), .ZN(new_n398));
  OAI21_X1  g197(.A(new_n381), .B1(new_n398), .B2(new_n391), .ZN(new_n399));
  NAND3_X1  g198(.A1(new_n395), .A2(new_n399), .A3(new_n378), .ZN(new_n400));
  NAND2_X1  g199(.A1(new_n393), .A2(new_n400), .ZN(new_n401));
  INV_X1    g200(.A(G227gat), .ZN(new_n402));
  NOR2_X1   g201(.A1(new_n402), .A2(new_n221), .ZN(new_n403));
  XNOR2_X1  g202(.A(new_n403), .B(KEYINPUT64), .ZN(new_n404));
  INV_X1    g203(.A(new_n404), .ZN(new_n405));
  OAI211_X1 g204(.A(new_n243), .B(new_n350), .C1(new_n260), .C2(new_n264), .ZN(new_n406));
  INV_X1    g205(.A(new_n406), .ZN(new_n407));
  AOI21_X1  g206(.A(new_n350), .B1(new_n272), .B2(new_n243), .ZN(new_n408));
  OAI21_X1  g207(.A(new_n405), .B1(new_n407), .B2(new_n408), .ZN(new_n409));
  NAND2_X1  g208(.A1(new_n409), .A2(KEYINPUT32), .ZN(new_n410));
  XOR2_X1   g209(.A(G15gat), .B(G43gat), .Z(new_n411));
  XNOR2_X1  g210(.A(new_n411), .B(KEYINPUT71), .ZN(new_n412));
  XOR2_X1   g211(.A(G71gat), .B(G99gat), .Z(new_n413));
  XNOR2_X1  g212(.A(new_n413), .B(KEYINPUT72), .ZN(new_n414));
  XNOR2_X1  g213(.A(new_n412), .B(new_n414), .ZN(new_n415));
  NAND2_X1  g214(.A1(new_n265), .A2(new_n343), .ZN(new_n416));
  AOI21_X1  g215(.A(new_n404), .B1(new_n416), .B2(new_n406), .ZN(new_n417));
  OAI211_X1 g216(.A(new_n410), .B(new_n415), .C1(KEYINPUT33), .C2(new_n417), .ZN(new_n418));
  INV_X1    g217(.A(KEYINPUT73), .ZN(new_n419));
  NOR2_X1   g218(.A1(new_n405), .A2(KEYINPUT34), .ZN(new_n420));
  NAND4_X1  g219(.A1(new_n416), .A2(new_n419), .A3(new_n406), .A4(new_n420), .ZN(new_n421));
  OAI21_X1  g220(.A(new_n415), .B1(new_n417), .B2(KEYINPUT33), .ZN(new_n422));
  INV_X1    g221(.A(KEYINPUT32), .ZN(new_n423));
  NOR2_X1   g222(.A1(new_n417), .A2(new_n423), .ZN(new_n424));
  NAND2_X1  g223(.A1(new_n422), .A2(new_n424), .ZN(new_n425));
  OAI211_X1 g224(.A(new_n416), .B(new_n406), .C1(new_n402), .C2(new_n221), .ZN(new_n426));
  NAND3_X1  g225(.A1(new_n416), .A2(new_n406), .A3(new_n420), .ZN(new_n427));
  AOI22_X1  g226(.A1(new_n426), .A2(KEYINPUT34), .B1(new_n427), .B2(KEYINPUT73), .ZN(new_n428));
  NAND4_X1  g227(.A1(new_n418), .A2(new_n421), .A3(new_n425), .A4(new_n428), .ZN(new_n429));
  NAND2_X1  g228(.A1(new_n426), .A2(KEYINPUT34), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n427), .A2(KEYINPUT73), .ZN(new_n431));
  NAND3_X1  g230(.A1(new_n430), .A2(new_n421), .A3(new_n431), .ZN(new_n432));
  NOR2_X1   g231(.A1(new_n422), .A2(new_n424), .ZN(new_n433));
  NAND2_X1  g232(.A1(new_n416), .A2(new_n406), .ZN(new_n434));
  AOI221_X4 g233(.A(new_n423), .B1(KEYINPUT33), .B2(new_n415), .C1(new_n434), .C2(new_n405), .ZN(new_n435));
  OAI21_X1  g234(.A(new_n432), .B1(new_n433), .B2(new_n435), .ZN(new_n436));
  NAND3_X1  g235(.A1(new_n401), .A2(new_n429), .A3(new_n436), .ZN(new_n437));
  OAI21_X1  g236(.A(KEYINPUT35), .B1(new_n371), .B2(new_n437), .ZN(new_n438));
  INV_X1    g237(.A(KEYINPUT85), .ZN(new_n439));
  NAND2_X1  g238(.A1(new_n438), .A2(new_n439), .ZN(new_n440));
  OAI211_X1 g239(.A(KEYINPUT85), .B(KEYINPUT35), .C1(new_n371), .C2(new_n437), .ZN(new_n441));
  NOR2_X1   g240(.A1(new_n365), .A2(new_n366), .ZN(new_n442));
  INV_X1    g241(.A(KEYINPUT82), .ZN(new_n443));
  OAI21_X1  g242(.A(new_n443), .B1(new_n357), .B2(new_n361), .ZN(new_n444));
  OAI211_X1 g243(.A(KEYINPUT82), .B(new_n363), .C1(new_n364), .C2(new_n301), .ZN(new_n445));
  NAND3_X1  g244(.A1(new_n444), .A2(new_n445), .A3(new_n299), .ZN(new_n446));
  OAI21_X1  g245(.A(new_n363), .B1(new_n364), .B2(new_n301), .ZN(new_n447));
  AOI21_X1  g246(.A(KEYINPUT6), .B1(new_n447), .B2(new_n300), .ZN(new_n448));
  AOI21_X1  g247(.A(new_n442), .B1(new_n446), .B2(new_n448), .ZN(new_n449));
  NOR2_X1   g248(.A1(new_n437), .A2(new_n449), .ZN(new_n450));
  INV_X1    g249(.A(KEYINPUT35), .ZN(new_n451));
  AOI21_X1  g250(.A(KEYINPUT30), .B1(new_n286), .B2(new_n288), .ZN(new_n452));
  NOR2_X1   g251(.A1(new_n452), .A2(new_n294), .ZN(new_n453));
  NAND3_X1  g252(.A1(new_n450), .A2(new_n451), .A3(new_n453), .ZN(new_n454));
  NAND3_X1  g253(.A1(new_n440), .A2(new_n441), .A3(new_n454), .ZN(new_n455));
  AND3_X1   g254(.A1(new_n393), .A2(KEYINPUT79), .A3(new_n400), .ZN(new_n456));
  AOI21_X1  g255(.A(KEYINPUT79), .B1(new_n393), .B2(new_n400), .ZN(new_n457));
  NOR2_X1   g256(.A1(new_n456), .A2(new_n457), .ZN(new_n458));
  INV_X1    g257(.A(KEYINPUT36), .ZN(new_n459));
  NOR3_X1   g258(.A1(new_n433), .A2(new_n432), .A3(new_n435), .ZN(new_n460));
  AOI22_X1  g259(.A1(new_n418), .A2(new_n425), .B1(new_n421), .B2(new_n428), .ZN(new_n461));
  OAI21_X1  g260(.A(new_n459), .B1(new_n460), .B2(new_n461), .ZN(new_n462));
  NAND3_X1  g261(.A1(new_n429), .A2(new_n436), .A3(KEYINPUT36), .ZN(new_n463));
  AOI22_X1  g262(.A1(new_n458), .A2(new_n371), .B1(new_n462), .B2(new_n463), .ZN(new_n464));
  OAI21_X1  g263(.A(new_n344), .B1(new_n347), .B2(new_n351), .ZN(new_n465));
  NAND3_X1  g264(.A1(new_n465), .A2(G225gat), .A3(G233gat), .ZN(new_n466));
  NAND3_X1  g265(.A1(new_n354), .A2(new_n302), .A3(new_n346), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n467), .A2(KEYINPUT39), .ZN(new_n468));
  INV_X1    g267(.A(KEYINPUT81), .ZN(new_n469));
  NAND2_X1  g268(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  NAND3_X1  g269(.A1(new_n467), .A2(KEYINPUT81), .A3(KEYINPUT39), .ZN(new_n471));
  NAND3_X1  g270(.A1(new_n466), .A2(new_n470), .A3(new_n471), .ZN(new_n472));
  NOR2_X1   g271(.A1(new_n360), .A2(new_n302), .ZN(new_n473));
  XNOR2_X1  g272(.A(KEYINPUT80), .B(KEYINPUT39), .ZN(new_n474));
  AOI21_X1  g273(.A(new_n299), .B1(new_n473), .B2(new_n474), .ZN(new_n475));
  NAND2_X1  g274(.A1(new_n472), .A2(new_n475), .ZN(new_n476));
  INV_X1    g275(.A(KEYINPUT40), .ZN(new_n477));
  NAND2_X1  g276(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  NAND3_X1  g277(.A1(new_n472), .A2(new_n475), .A3(KEYINPUT40), .ZN(new_n479));
  AND3_X1   g278(.A1(new_n478), .A2(new_n446), .A3(new_n479), .ZN(new_n480));
  INV_X1    g279(.A(KEYINPUT83), .ZN(new_n481));
  OAI211_X1 g280(.A(new_n480), .B(new_n481), .C1(new_n452), .C2(new_n294), .ZN(new_n482));
  NAND3_X1  g281(.A1(new_n478), .A2(new_n446), .A3(new_n479), .ZN(new_n483));
  OAI21_X1  g282(.A(KEYINPUT83), .B1(new_n453), .B2(new_n483), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n482), .A2(new_n484), .ZN(new_n485));
  INV_X1    g284(.A(KEYINPUT37), .ZN(new_n486));
  NAND3_X1  g285(.A1(new_n274), .A2(new_n486), .A3(new_n284), .ZN(new_n487));
  NAND2_X1  g286(.A1(new_n487), .A2(new_n277), .ZN(new_n488));
  AOI21_X1  g287(.A(new_n486), .B1(new_n274), .B2(new_n284), .ZN(new_n489));
  OAI21_X1  g288(.A(KEYINPUT38), .B1(new_n488), .B2(new_n489), .ZN(new_n490));
  INV_X1    g289(.A(KEYINPUT84), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  INV_X1    g291(.A(new_n488), .ZN(new_n493));
  AOI21_X1  g292(.A(new_n266), .B1(new_n272), .B2(new_n243), .ZN(new_n494));
  OAI21_X1  g293(.A(new_n279), .B1(new_n494), .B2(new_n222), .ZN(new_n495));
  AOI21_X1  g294(.A(new_n486), .B1(new_n495), .B2(new_n282), .ZN(new_n496));
  OAI211_X1 g295(.A(new_n279), .B(new_n219), .C1(new_n283), .C2(new_n222), .ZN(new_n497));
  AOI21_X1  g296(.A(KEYINPUT38), .B1(new_n496), .B2(new_n497), .ZN(new_n498));
  AOI22_X1  g297(.A1(new_n493), .A2(new_n498), .B1(new_n286), .B2(new_n288), .ZN(new_n499));
  OAI211_X1 g298(.A(KEYINPUT84), .B(KEYINPUT38), .C1(new_n488), .C2(new_n489), .ZN(new_n500));
  NAND4_X1  g299(.A1(new_n492), .A2(new_n499), .A3(new_n449), .A4(new_n500), .ZN(new_n501));
  NAND2_X1  g300(.A1(new_n501), .A2(new_n401), .ZN(new_n502));
  OAI21_X1  g301(.A(new_n464), .B1(new_n485), .B2(new_n502), .ZN(new_n503));
  AND3_X1   g302(.A1(new_n455), .A2(new_n503), .A3(KEYINPUT86), .ZN(new_n504));
  AOI21_X1  g303(.A(KEYINPUT86), .B1(new_n455), .B2(new_n503), .ZN(new_n505));
  XNOR2_X1  g304(.A(G15gat), .B(G22gat), .ZN(new_n506));
  NOR2_X1   g305(.A1(new_n506), .A2(G1gat), .ZN(new_n507));
  OAI21_X1  g306(.A(G8gat), .B1(new_n507), .B2(KEYINPUT90), .ZN(new_n508));
  INV_X1    g307(.A(KEYINPUT16), .ZN(new_n509));
  OAI21_X1  g308(.A(new_n506), .B1(new_n509), .B2(G1gat), .ZN(new_n510));
  OAI21_X1  g309(.A(new_n510), .B1(G1gat), .B2(new_n506), .ZN(new_n511));
  XNOR2_X1  g310(.A(new_n508), .B(new_n511), .ZN(new_n512));
  XNOR2_X1  g311(.A(G43gat), .B(G50gat), .ZN(new_n513));
  AND2_X1   g312(.A1(new_n513), .A2(KEYINPUT15), .ZN(new_n514));
  INV_X1    g313(.A(KEYINPUT14), .ZN(new_n515));
  INV_X1    g314(.A(G29gat), .ZN(new_n516));
  NAND2_X1  g315(.A1(new_n516), .A2(KEYINPUT87), .ZN(new_n517));
  INV_X1    g316(.A(KEYINPUT87), .ZN(new_n518));
  NAND2_X1  g317(.A1(new_n518), .A2(G29gat), .ZN(new_n519));
  NAND3_X1  g318(.A1(new_n517), .A2(new_n519), .A3(G36gat), .ZN(new_n520));
  INV_X1    g319(.A(G36gat), .ZN(new_n521));
  NAND2_X1  g320(.A1(new_n516), .A2(new_n521), .ZN(new_n522));
  AOI21_X1  g321(.A(new_n515), .B1(new_n520), .B2(new_n522), .ZN(new_n523));
  AOI21_X1  g322(.A(KEYINPUT14), .B1(new_n516), .B2(new_n521), .ZN(new_n524));
  OAI21_X1  g323(.A(new_n514), .B1(new_n523), .B2(new_n524), .ZN(new_n525));
  NAND2_X1  g324(.A1(new_n525), .A2(KEYINPUT88), .ZN(new_n526));
  INV_X1    g325(.A(KEYINPUT88), .ZN(new_n527));
  OAI211_X1 g326(.A(new_n527), .B(new_n514), .C1(new_n523), .C2(new_n524), .ZN(new_n528));
  NAND2_X1  g327(.A1(new_n526), .A2(new_n528), .ZN(new_n529));
  INV_X1    g328(.A(KEYINPUT17), .ZN(new_n530));
  INV_X1    g329(.A(KEYINPUT89), .ZN(new_n531));
  NOR2_X1   g330(.A1(new_n513), .A2(new_n531), .ZN(new_n532));
  XNOR2_X1  g331(.A(new_n532), .B(KEYINPUT15), .ZN(new_n533));
  NOR2_X1   g332(.A1(new_n523), .A2(new_n524), .ZN(new_n534));
  NAND2_X1  g333(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  AND3_X1   g334(.A1(new_n529), .A2(new_n530), .A3(new_n535), .ZN(new_n536));
  AOI21_X1  g335(.A(new_n530), .B1(new_n529), .B2(new_n535), .ZN(new_n537));
  OAI21_X1  g336(.A(new_n512), .B1(new_n536), .B2(new_n537), .ZN(new_n538));
  NAND2_X1  g337(.A1(G229gat), .A2(G233gat), .ZN(new_n539));
  NAND2_X1  g338(.A1(new_n529), .A2(new_n535), .ZN(new_n540));
  INV_X1    g339(.A(new_n512), .ZN(new_n541));
  NAND2_X1  g340(.A1(new_n540), .A2(new_n541), .ZN(new_n542));
  NAND3_X1  g341(.A1(new_n538), .A2(new_n539), .A3(new_n542), .ZN(new_n543));
  INV_X1    g342(.A(KEYINPUT18), .ZN(new_n544));
  NAND2_X1  g343(.A1(new_n543), .A2(new_n544), .ZN(new_n545));
  INV_X1    g344(.A(new_n545), .ZN(new_n546));
  NAND2_X1  g345(.A1(new_n546), .A2(KEYINPUT93), .ZN(new_n547));
  NAND4_X1  g346(.A1(new_n538), .A2(KEYINPUT18), .A3(new_n539), .A4(new_n542), .ZN(new_n548));
  XNOR2_X1  g347(.A(new_n539), .B(KEYINPUT13), .ZN(new_n549));
  INV_X1    g348(.A(new_n549), .ZN(new_n550));
  INV_X1    g349(.A(KEYINPUT91), .ZN(new_n551));
  INV_X1    g350(.A(new_n540), .ZN(new_n552));
  AOI21_X1  g351(.A(new_n551), .B1(new_n552), .B2(new_n512), .ZN(new_n553));
  NAND4_X1  g352(.A1(new_n512), .A2(new_n529), .A3(new_n551), .A4(new_n535), .ZN(new_n554));
  NAND2_X1  g353(.A1(new_n542), .A2(new_n554), .ZN(new_n555));
  OAI21_X1  g354(.A(new_n550), .B1(new_n553), .B2(new_n555), .ZN(new_n556));
  XNOR2_X1  g355(.A(G113gat), .B(G141gat), .ZN(new_n557));
  XNOR2_X1  g356(.A(new_n557), .B(G197gat), .ZN(new_n558));
  XNOR2_X1  g357(.A(KEYINPUT11), .B(G169gat), .ZN(new_n559));
  XNOR2_X1  g358(.A(new_n558), .B(new_n559), .ZN(new_n560));
  XOR2_X1   g359(.A(new_n560), .B(KEYINPUT12), .Z(new_n561));
  NAND3_X1  g360(.A1(new_n548), .A2(new_n556), .A3(new_n561), .ZN(new_n562));
  INV_X1    g361(.A(new_n562), .ZN(new_n563));
  AOI21_X1  g362(.A(KEYINPUT93), .B1(new_n543), .B2(new_n544), .ZN(new_n564));
  INV_X1    g363(.A(new_n564), .ZN(new_n565));
  NAND3_X1  g364(.A1(new_n547), .A2(new_n563), .A3(new_n565), .ZN(new_n566));
  AND3_X1   g365(.A1(new_n548), .A2(new_n556), .A3(KEYINPUT92), .ZN(new_n567));
  AOI21_X1  g366(.A(KEYINPUT92), .B1(new_n548), .B2(new_n556), .ZN(new_n568));
  NOR3_X1   g367(.A1(new_n567), .A2(new_n568), .A3(new_n546), .ZN(new_n569));
  OAI21_X1  g368(.A(new_n566), .B1(new_n569), .B2(new_n561), .ZN(new_n570));
  INV_X1    g369(.A(new_n570), .ZN(new_n571));
  NOR3_X1   g370(.A1(new_n504), .A2(new_n505), .A3(new_n571), .ZN(new_n572));
  XOR2_X1   g371(.A(G183gat), .B(G211gat), .Z(new_n573));
  XNOR2_X1  g372(.A(new_n573), .B(KEYINPUT97), .ZN(new_n574));
  XNOR2_X1  g373(.A(new_n574), .B(KEYINPUT19), .ZN(new_n575));
  XNOR2_X1  g374(.A(new_n575), .B(KEYINPUT20), .ZN(new_n576));
  INV_X1    g375(.A(new_n576), .ZN(new_n577));
  INV_X1    g376(.A(KEYINPUT21), .ZN(new_n578));
  NAND2_X1  g377(.A1(G71gat), .A2(G78gat), .ZN(new_n579));
  INV_X1    g378(.A(G71gat), .ZN(new_n580));
  INV_X1    g379(.A(G78gat), .ZN(new_n581));
  NAND2_X1  g380(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  XNOR2_X1  g381(.A(G57gat), .B(G64gat), .ZN(new_n583));
  INV_X1    g382(.A(KEYINPUT9), .ZN(new_n584));
  OAI211_X1 g383(.A(new_n579), .B(new_n582), .C1(new_n583), .C2(new_n584), .ZN(new_n585));
  INV_X1    g384(.A(KEYINPUT94), .ZN(new_n586));
  NAND2_X1  g385(.A1(new_n583), .A2(new_n586), .ZN(new_n587));
  NAND3_X1  g386(.A1(new_n580), .A2(new_n581), .A3(KEYINPUT9), .ZN(new_n588));
  NAND2_X1  g387(.A1(new_n588), .A2(new_n579), .ZN(new_n589));
  NAND2_X1  g388(.A1(new_n587), .A2(new_n589), .ZN(new_n590));
  NOR2_X1   g389(.A1(new_n583), .A2(new_n586), .ZN(new_n591));
  OAI21_X1  g390(.A(new_n585), .B1(new_n590), .B2(new_n591), .ZN(new_n592));
  OAI21_X1  g391(.A(new_n512), .B1(new_n578), .B2(new_n592), .ZN(new_n593));
  XNOR2_X1  g392(.A(new_n593), .B(KEYINPUT96), .ZN(new_n594));
  XOR2_X1   g393(.A(G127gat), .B(G155gat), .Z(new_n595));
  NAND2_X1  g394(.A1(new_n594), .A2(new_n595), .ZN(new_n596));
  INV_X1    g395(.A(new_n596), .ZN(new_n597));
  NOR2_X1   g396(.A1(new_n594), .A2(new_n595), .ZN(new_n598));
  OAI21_X1  g397(.A(new_n577), .B1(new_n597), .B2(new_n598), .ZN(new_n599));
  INV_X1    g398(.A(new_n598), .ZN(new_n600));
  NAND3_X1  g399(.A1(new_n600), .A2(new_n596), .A3(new_n576), .ZN(new_n601));
  NAND2_X1  g400(.A1(new_n592), .A2(new_n578), .ZN(new_n602));
  NAND2_X1  g401(.A1(G231gat), .A2(G233gat), .ZN(new_n603));
  XNOR2_X1  g402(.A(new_n603), .B(KEYINPUT95), .ZN(new_n604));
  XNOR2_X1  g403(.A(new_n602), .B(new_n604), .ZN(new_n605));
  AND3_X1   g404(.A1(new_n599), .A2(new_n601), .A3(new_n605), .ZN(new_n606));
  AOI21_X1  g405(.A(new_n605), .B1(new_n599), .B2(new_n601), .ZN(new_n607));
  NOR2_X1   g406(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  INV_X1    g407(.A(new_n608), .ZN(new_n609));
  NAND2_X1  g408(.A1(G99gat), .A2(G106gat), .ZN(new_n610));
  INV_X1    g409(.A(G85gat), .ZN(new_n611));
  INV_X1    g410(.A(G92gat), .ZN(new_n612));
  AOI22_X1  g411(.A1(KEYINPUT8), .A2(new_n610), .B1(new_n611), .B2(new_n612), .ZN(new_n613));
  INV_X1    g412(.A(KEYINPUT7), .ZN(new_n614));
  OAI21_X1  g413(.A(new_n614), .B1(new_n611), .B2(new_n612), .ZN(new_n615));
  NAND3_X1  g414(.A1(KEYINPUT7), .A2(G85gat), .A3(G92gat), .ZN(new_n616));
  NAND3_X1  g415(.A1(new_n613), .A2(new_n615), .A3(new_n616), .ZN(new_n617));
  XNOR2_X1  g416(.A(G99gat), .B(G106gat), .ZN(new_n618));
  INV_X1    g417(.A(new_n618), .ZN(new_n619));
  NAND2_X1  g418(.A1(new_n617), .A2(new_n619), .ZN(new_n620));
  NAND4_X1  g419(.A1(new_n613), .A2(new_n618), .A3(new_n615), .A4(new_n616), .ZN(new_n621));
  NAND2_X1  g420(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  INV_X1    g421(.A(new_n622), .ZN(new_n623));
  AND2_X1   g422(.A1(G232gat), .A2(G233gat), .ZN(new_n624));
  AOI22_X1  g423(.A1(new_n540), .A2(new_n623), .B1(KEYINPUT41), .B2(new_n624), .ZN(new_n625));
  NOR2_X1   g424(.A1(new_n536), .A2(new_n537), .ZN(new_n626));
  XOR2_X1   g425(.A(new_n622), .B(KEYINPUT98), .Z(new_n627));
  OAI21_X1  g426(.A(new_n625), .B1(new_n626), .B2(new_n627), .ZN(new_n628));
  NAND2_X1  g427(.A1(new_n628), .A2(KEYINPUT99), .ZN(new_n629));
  INV_X1    g428(.A(KEYINPUT99), .ZN(new_n630));
  OAI211_X1 g429(.A(new_n630), .B(new_n625), .C1(new_n626), .C2(new_n627), .ZN(new_n631));
  XNOR2_X1  g430(.A(G190gat), .B(G218gat), .ZN(new_n632));
  NAND3_X1  g431(.A1(new_n629), .A2(new_n631), .A3(new_n632), .ZN(new_n633));
  INV_X1    g432(.A(new_n632), .ZN(new_n634));
  NAND3_X1  g433(.A1(new_n628), .A2(KEYINPUT99), .A3(new_n634), .ZN(new_n635));
  NAND2_X1  g434(.A1(new_n633), .A2(new_n635), .ZN(new_n636));
  INV_X1    g435(.A(KEYINPUT100), .ZN(new_n637));
  NOR2_X1   g436(.A1(new_n624), .A2(KEYINPUT41), .ZN(new_n638));
  XNOR2_X1  g437(.A(G134gat), .B(G162gat), .ZN(new_n639));
  XNOR2_X1  g438(.A(new_n638), .B(new_n639), .ZN(new_n640));
  OAI21_X1  g439(.A(new_n636), .B1(new_n637), .B2(new_n640), .ZN(new_n641));
  XNOR2_X1  g440(.A(new_n640), .B(KEYINPUT100), .ZN(new_n642));
  INV_X1    g441(.A(new_n642), .ZN(new_n643));
  NAND3_X1  g442(.A1(new_n633), .A2(new_n643), .A3(new_n635), .ZN(new_n644));
  NAND2_X1  g443(.A1(new_n641), .A2(new_n644), .ZN(new_n645));
  NOR2_X1   g444(.A1(new_n609), .A2(new_n645), .ZN(new_n646));
  NAND2_X1  g445(.A1(G230gat), .A2(G233gat), .ZN(new_n647));
  INV_X1    g446(.A(new_n647), .ZN(new_n648));
  NAND2_X1  g447(.A1(new_n592), .A2(new_n622), .ZN(new_n649));
  OR2_X1    g448(.A1(new_n583), .A2(new_n586), .ZN(new_n650));
  NAND3_X1  g449(.A1(new_n650), .A2(new_n589), .A3(new_n587), .ZN(new_n651));
  NAND4_X1  g450(.A1(new_n651), .A2(new_n585), .A3(new_n621), .A4(new_n620), .ZN(new_n652));
  INV_X1    g451(.A(KEYINPUT10), .ZN(new_n653));
  NAND3_X1  g452(.A1(new_n649), .A2(new_n652), .A3(new_n653), .ZN(new_n654));
  NAND4_X1  g453(.A1(new_n623), .A2(KEYINPUT10), .A3(new_n651), .A4(new_n585), .ZN(new_n655));
  AOI21_X1  g454(.A(new_n648), .B1(new_n654), .B2(new_n655), .ZN(new_n656));
  NAND2_X1  g455(.A1(new_n649), .A2(new_n652), .ZN(new_n657));
  AOI21_X1  g456(.A(new_n656), .B1(new_n657), .B2(new_n648), .ZN(new_n658));
  XNOR2_X1  g457(.A(G176gat), .B(G204gat), .ZN(new_n659));
  XNOR2_X1  g458(.A(new_n659), .B(KEYINPUT101), .ZN(new_n660));
  XNOR2_X1  g459(.A(G120gat), .B(G148gat), .ZN(new_n661));
  XNOR2_X1  g460(.A(new_n660), .B(new_n661), .ZN(new_n662));
  OR2_X1    g461(.A1(new_n658), .A2(new_n662), .ZN(new_n663));
  NAND2_X1  g462(.A1(new_n654), .A2(new_n655), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n664), .A2(new_n647), .ZN(new_n665));
  NAND2_X1  g464(.A1(new_n657), .A2(new_n648), .ZN(new_n666));
  NAND3_X1  g465(.A1(new_n665), .A2(new_n666), .A3(new_n662), .ZN(new_n667));
  NAND2_X1  g466(.A1(new_n663), .A2(new_n667), .ZN(new_n668));
  INV_X1    g467(.A(new_n668), .ZN(new_n669));
  NAND3_X1  g468(.A1(new_n572), .A2(new_n646), .A3(new_n669), .ZN(new_n670));
  INV_X1    g469(.A(new_n670), .ZN(new_n671));
  INV_X1    g470(.A(new_n370), .ZN(new_n672));
  AND2_X1   g471(.A1(new_n672), .A2(KEYINPUT102), .ZN(new_n673));
  NOR2_X1   g472(.A1(new_n672), .A2(KEYINPUT102), .ZN(new_n674));
  NOR2_X1   g473(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  INV_X1    g474(.A(new_n675), .ZN(new_n676));
  NAND2_X1  g475(.A1(new_n671), .A2(new_n676), .ZN(new_n677));
  XNOR2_X1  g476(.A(new_n677), .B(G1gat), .ZN(G1324gat));
  NOR2_X1   g477(.A1(new_n670), .A2(new_n453), .ZN(new_n679));
  NOR2_X1   g478(.A1(KEYINPUT103), .A2(KEYINPUT42), .ZN(new_n680));
  XNOR2_X1  g479(.A(new_n680), .B(new_n509), .ZN(new_n681));
  NAND2_X1  g480(.A1(new_n679), .A2(new_n681), .ZN(new_n682));
  OR2_X1    g481(.A1(new_n682), .A2(G8gat), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n682), .A2(G8gat), .ZN(new_n684));
  OAI211_X1 g483(.A(new_n683), .B(new_n684), .C1(KEYINPUT42), .C2(new_n679), .ZN(G1325gat));
  NAND2_X1  g484(.A1(new_n462), .A2(new_n463), .ZN(new_n686));
  INV_X1    g485(.A(new_n686), .ZN(new_n687));
  AND3_X1   g486(.A1(new_n671), .A2(G15gat), .A3(new_n687), .ZN(new_n688));
  NOR2_X1   g487(.A1(new_n460), .A2(new_n461), .ZN(new_n689));
  AOI21_X1  g488(.A(G15gat), .B1(new_n671), .B2(new_n689), .ZN(new_n690));
  NOR2_X1   g489(.A1(new_n688), .A2(new_n690), .ZN(G1326gat));
  INV_X1    g490(.A(new_n458), .ZN(new_n692));
  NOR2_X1   g491(.A1(new_n670), .A2(new_n692), .ZN(new_n693));
  XNOR2_X1  g492(.A(new_n693), .B(new_n376), .ZN(new_n694));
  XNOR2_X1  g493(.A(KEYINPUT104), .B(KEYINPUT43), .ZN(new_n695));
  XNOR2_X1  g494(.A(new_n694), .B(new_n695), .ZN(G1327gat));
  NAND2_X1  g495(.A1(new_n455), .A2(new_n503), .ZN(new_n697));
  INV_X1    g496(.A(KEYINPUT86), .ZN(new_n698));
  NAND2_X1  g497(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  NAND3_X1  g498(.A1(new_n455), .A2(new_n503), .A3(KEYINPUT86), .ZN(new_n700));
  NAND2_X1  g499(.A1(new_n609), .A2(new_n669), .ZN(new_n701));
  AND2_X1   g500(.A1(new_n641), .A2(new_n644), .ZN(new_n702));
  NOR2_X1   g501(.A1(new_n701), .A2(new_n702), .ZN(new_n703));
  NAND4_X1  g502(.A1(new_n699), .A2(new_n570), .A3(new_n700), .A4(new_n703), .ZN(new_n704));
  INV_X1    g503(.A(new_n704), .ZN(new_n705));
  NAND2_X1  g504(.A1(new_n517), .A2(new_n519), .ZN(new_n706));
  NAND3_X1  g505(.A1(new_n705), .A2(new_n706), .A3(new_n676), .ZN(new_n707));
  XNOR2_X1  g506(.A(new_n707), .B(KEYINPUT45), .ZN(new_n708));
  AOI21_X1  g507(.A(new_n702), .B1(new_n455), .B2(new_n503), .ZN(new_n709));
  XOR2_X1   g508(.A(KEYINPUT105), .B(KEYINPUT44), .Z(new_n710));
  NAND2_X1  g509(.A1(new_n709), .A2(new_n710), .ZN(new_n711));
  NOR3_X1   g510(.A1(new_n504), .A2(new_n505), .A3(new_n702), .ZN(new_n712));
  INV_X1    g511(.A(KEYINPUT44), .ZN(new_n713));
  OAI21_X1  g512(.A(new_n711), .B1(new_n712), .B2(new_n713), .ZN(new_n714));
  NOR2_X1   g513(.A1(new_n701), .A2(new_n571), .ZN(new_n715));
  NAND2_X1  g514(.A1(new_n714), .A2(new_n715), .ZN(new_n716));
  NOR2_X1   g515(.A1(new_n716), .A2(new_n675), .ZN(new_n717));
  OAI21_X1  g516(.A(new_n708), .B1(new_n706), .B2(new_n717), .ZN(G1328gat));
  INV_X1    g517(.A(new_n453), .ZN(new_n719));
  NAND3_X1  g518(.A1(new_n705), .A2(new_n521), .A3(new_n719), .ZN(new_n720));
  NAND2_X1  g519(.A1(new_n720), .A2(KEYINPUT46), .ZN(new_n721));
  XNOR2_X1  g520(.A(new_n721), .B(KEYINPUT106), .ZN(new_n722));
  OAI21_X1  g521(.A(G36gat), .B1(new_n716), .B2(new_n453), .ZN(new_n723));
  OAI211_X1 g522(.A(new_n722), .B(new_n723), .C1(KEYINPUT46), .C2(new_n720), .ZN(G1329gat));
  INV_X1    g523(.A(new_n689), .ZN(new_n725));
  NOR3_X1   g524(.A1(new_n704), .A2(G43gat), .A3(new_n725), .ZN(new_n726));
  INV_X1    g525(.A(new_n715), .ZN(new_n727));
  NAND3_X1  g526(.A1(new_n699), .A2(new_n700), .A3(new_n645), .ZN(new_n728));
  NAND2_X1  g527(.A1(new_n728), .A2(KEYINPUT44), .ZN(new_n729));
  AOI21_X1  g528(.A(new_n727), .B1(new_n729), .B2(new_n711), .ZN(new_n730));
  NAND2_X1  g529(.A1(new_n730), .A2(new_n687), .ZN(new_n731));
  AOI21_X1  g530(.A(new_n726), .B1(new_n731), .B2(G43gat), .ZN(new_n732));
  XNOR2_X1  g531(.A(new_n732), .B(KEYINPUT47), .ZN(G1330gat));
  INV_X1    g532(.A(KEYINPUT48), .ZN(new_n734));
  INV_X1    g533(.A(new_n401), .ZN(new_n735));
  NAND3_X1  g534(.A1(new_n714), .A2(new_n735), .A3(new_n715), .ZN(new_n736));
  NAND2_X1  g535(.A1(new_n736), .A2(G50gat), .ZN(new_n737));
  NOR2_X1   g536(.A1(new_n692), .A2(G50gat), .ZN(new_n738));
  NAND2_X1  g537(.A1(new_n705), .A2(new_n738), .ZN(new_n739));
  AOI21_X1  g538(.A(new_n734), .B1(new_n737), .B2(new_n739), .ZN(new_n740));
  NAND4_X1  g539(.A1(new_n572), .A2(KEYINPUT107), .A3(new_n703), .A4(new_n738), .ZN(new_n741));
  INV_X1    g540(.A(KEYINPUT107), .ZN(new_n742));
  INV_X1    g541(.A(new_n738), .ZN(new_n743));
  OAI21_X1  g542(.A(new_n742), .B1(new_n704), .B2(new_n743), .ZN(new_n744));
  NAND3_X1  g543(.A1(new_n741), .A2(new_n744), .A3(new_n734), .ZN(new_n745));
  NAND2_X1  g544(.A1(new_n730), .A2(new_n458), .ZN(new_n746));
  AOI21_X1  g545(.A(new_n745), .B1(new_n746), .B2(G50gat), .ZN(new_n747));
  NOR3_X1   g546(.A1(new_n740), .A2(KEYINPUT108), .A3(new_n747), .ZN(new_n748));
  INV_X1    g547(.A(KEYINPUT108), .ZN(new_n749));
  AOI21_X1  g548(.A(new_n373), .B1(new_n730), .B2(new_n735), .ZN(new_n750));
  INV_X1    g549(.A(new_n739), .ZN(new_n751));
  OAI21_X1  g550(.A(KEYINPUT48), .B1(new_n750), .B2(new_n751), .ZN(new_n752));
  AND2_X1   g551(.A1(new_n744), .A2(new_n734), .ZN(new_n753));
  AOI22_X1  g552(.A1(new_n728), .A2(KEYINPUT44), .B1(new_n709), .B2(new_n710), .ZN(new_n754));
  NOR3_X1   g553(.A1(new_n754), .A2(new_n692), .A3(new_n727), .ZN(new_n755));
  OAI211_X1 g554(.A(new_n741), .B(new_n753), .C1(new_n755), .C2(new_n373), .ZN(new_n756));
  AOI21_X1  g555(.A(new_n749), .B1(new_n752), .B2(new_n756), .ZN(new_n757));
  NOR2_X1   g556(.A1(new_n748), .A2(new_n757), .ZN(G1331gat));
  NAND4_X1  g557(.A1(new_n697), .A2(new_n571), .A3(new_n646), .A4(new_n668), .ZN(new_n759));
  NOR2_X1   g558(.A1(new_n759), .A2(new_n675), .ZN(new_n760));
  XOR2_X1   g559(.A(new_n760), .B(G57gat), .Z(G1332gat));
  XOR2_X1   g560(.A(new_n759), .B(KEYINPUT109), .Z(new_n762));
  NOR2_X1   g561(.A1(new_n762), .A2(new_n453), .ZN(new_n763));
  NOR2_X1   g562(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n764));
  AND2_X1   g563(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n765));
  OAI21_X1  g564(.A(new_n763), .B1(new_n764), .B2(new_n765), .ZN(new_n766));
  OAI21_X1  g565(.A(new_n766), .B1(new_n763), .B2(new_n764), .ZN(G1333gat));
  NOR3_X1   g566(.A1(new_n759), .A2(G71gat), .A3(new_n725), .ZN(new_n768));
  OR2_X1    g567(.A1(new_n762), .A2(new_n686), .ZN(new_n769));
  AOI21_X1  g568(.A(new_n768), .B1(new_n769), .B2(G71gat), .ZN(new_n770));
  XNOR2_X1  g569(.A(new_n770), .B(KEYINPUT50), .ZN(G1334gat));
  NOR2_X1   g570(.A1(new_n762), .A2(new_n692), .ZN(new_n772));
  XNOR2_X1  g571(.A(new_n772), .B(new_n581), .ZN(G1335gat));
  NAND3_X1  g572(.A1(new_n609), .A2(new_n571), .A3(new_n668), .ZN(new_n774));
  NOR2_X1   g573(.A1(new_n754), .A2(new_n774), .ZN(new_n775));
  INV_X1    g574(.A(new_n775), .ZN(new_n776));
  OAI21_X1  g575(.A(G85gat), .B1(new_n776), .B2(new_n675), .ZN(new_n777));
  INV_X1    g576(.A(KEYINPUT51), .ZN(new_n778));
  AOI211_X1 g577(.A(new_n570), .B(new_n608), .C1(KEYINPUT110), .C2(new_n778), .ZN(new_n779));
  NAND2_X1  g578(.A1(new_n709), .A2(new_n779), .ZN(new_n780));
  NOR2_X1   g579(.A1(new_n778), .A2(KEYINPUT110), .ZN(new_n781));
  INV_X1    g580(.A(new_n781), .ZN(new_n782));
  XNOR2_X1  g581(.A(new_n780), .B(new_n782), .ZN(new_n783));
  AND2_X1   g582(.A1(new_n783), .A2(new_n668), .ZN(new_n784));
  NAND3_X1  g583(.A1(new_n784), .A2(new_n611), .A3(new_n676), .ZN(new_n785));
  NAND2_X1  g584(.A1(new_n777), .A2(new_n785), .ZN(G1336gat));
  NAND2_X1  g585(.A1(new_n775), .A2(new_n719), .ZN(new_n787));
  NOR2_X1   g586(.A1(new_n453), .A2(G92gat), .ZN(new_n788));
  AOI22_X1  g587(.A1(new_n787), .A2(G92gat), .B1(new_n784), .B2(new_n788), .ZN(new_n789));
  XOR2_X1   g588(.A(KEYINPUT111), .B(KEYINPUT52), .Z(new_n790));
  XNOR2_X1  g589(.A(new_n789), .B(new_n790), .ZN(G1337gat));
  OAI21_X1  g590(.A(G99gat), .B1(new_n776), .B2(new_n686), .ZN(new_n792));
  NOR3_X1   g591(.A1(new_n725), .A2(G99gat), .A3(new_n669), .ZN(new_n793));
  XNOR2_X1  g592(.A(new_n793), .B(KEYINPUT112), .ZN(new_n794));
  NAND2_X1  g593(.A1(new_n783), .A2(new_n794), .ZN(new_n795));
  NAND2_X1  g594(.A1(new_n792), .A2(new_n795), .ZN(G1338gat));
  OAI21_X1  g595(.A(G106gat), .B1(new_n776), .B2(new_n401), .ZN(new_n797));
  NOR2_X1   g596(.A1(new_n401), .A2(G106gat), .ZN(new_n798));
  AOI21_X1  g597(.A(KEYINPUT53), .B1(new_n784), .B2(new_n798), .ZN(new_n799));
  NAND2_X1  g598(.A1(new_n797), .A2(new_n799), .ZN(new_n800));
  NAND2_X1  g599(.A1(new_n775), .A2(new_n458), .ZN(new_n801));
  AOI22_X1  g600(.A1(new_n801), .A2(G106gat), .B1(new_n784), .B2(new_n798), .ZN(new_n802));
  INV_X1    g601(.A(KEYINPUT53), .ZN(new_n803));
  OAI21_X1  g602(.A(new_n800), .B1(new_n802), .B2(new_n803), .ZN(G1339gat));
  INV_X1    g603(.A(KEYINPUT113), .ZN(new_n805));
  NAND3_X1  g604(.A1(new_n654), .A2(new_n655), .A3(new_n648), .ZN(new_n806));
  NAND3_X1  g605(.A1(new_n665), .A2(KEYINPUT54), .A3(new_n806), .ZN(new_n807));
  INV_X1    g606(.A(KEYINPUT54), .ZN(new_n808));
  AOI21_X1  g607(.A(new_n662), .B1(new_n656), .B2(new_n808), .ZN(new_n809));
  NAND3_X1  g608(.A1(new_n807), .A2(KEYINPUT55), .A3(new_n809), .ZN(new_n810));
  NAND2_X1  g609(.A1(new_n810), .A2(new_n667), .ZN(new_n811));
  AOI21_X1  g610(.A(KEYINPUT55), .B1(new_n807), .B2(new_n809), .ZN(new_n812));
  OAI21_X1  g611(.A(new_n805), .B1(new_n811), .B2(new_n812), .ZN(new_n813));
  INV_X1    g612(.A(new_n812), .ZN(new_n814));
  NAND4_X1  g613(.A1(new_n814), .A2(KEYINPUT113), .A3(new_n667), .A4(new_n810), .ZN(new_n815));
  AND2_X1   g614(.A1(new_n813), .A2(new_n815), .ZN(new_n816));
  INV_X1    g615(.A(new_n561), .ZN(new_n817));
  AND2_X1   g616(.A1(new_n548), .A2(new_n556), .ZN(new_n818));
  OAI21_X1  g617(.A(new_n545), .B1(new_n818), .B2(KEYINPUT92), .ZN(new_n819));
  OAI21_X1  g618(.A(new_n817), .B1(new_n819), .B2(new_n567), .ZN(new_n820));
  AOI21_X1  g619(.A(new_n816), .B1(new_n820), .B2(new_n566), .ZN(new_n821));
  INV_X1    g620(.A(KEYINPUT93), .ZN(new_n822));
  NOR2_X1   g621(.A1(new_n545), .A2(new_n822), .ZN(new_n823));
  NOR3_X1   g622(.A1(new_n823), .A2(new_n562), .A3(new_n564), .ZN(new_n824));
  NAND2_X1  g623(.A1(new_n538), .A2(new_n542), .ZN(new_n825));
  NAND3_X1  g624(.A1(new_n825), .A2(G229gat), .A3(G233gat), .ZN(new_n826));
  OR3_X1    g625(.A1(new_n553), .A2(new_n555), .A3(new_n550), .ZN(new_n827));
  AOI21_X1  g626(.A(new_n560), .B1(new_n826), .B2(new_n827), .ZN(new_n828));
  NOR3_X1   g627(.A1(new_n824), .A2(new_n669), .A3(new_n828), .ZN(new_n829));
  OAI21_X1  g628(.A(new_n702), .B1(new_n821), .B2(new_n829), .ZN(new_n830));
  INV_X1    g629(.A(KEYINPUT114), .ZN(new_n831));
  OAI21_X1  g630(.A(new_n831), .B1(new_n824), .B2(new_n828), .ZN(new_n832));
  INV_X1    g631(.A(new_n828), .ZN(new_n833));
  NAND3_X1  g632(.A1(new_n566), .A2(new_n833), .A3(KEYINPUT114), .ZN(new_n834));
  NAND2_X1  g633(.A1(new_n813), .A2(new_n815), .ZN(new_n835));
  NAND4_X1  g634(.A1(new_n645), .A2(new_n832), .A3(new_n834), .A4(new_n835), .ZN(new_n836));
  AOI21_X1  g635(.A(new_n608), .B1(new_n830), .B2(new_n836), .ZN(new_n837));
  AND4_X1   g636(.A1(new_n571), .A2(new_n702), .A3(new_n608), .A4(new_n669), .ZN(new_n838));
  OAI21_X1  g637(.A(new_n692), .B1(new_n837), .B2(new_n838), .ZN(new_n839));
  INV_X1    g638(.A(KEYINPUT115), .ZN(new_n840));
  AOI21_X1  g639(.A(new_n725), .B1(new_n839), .B2(new_n840), .ZN(new_n841));
  NAND2_X1  g640(.A1(new_n676), .A2(new_n453), .ZN(new_n842));
  INV_X1    g641(.A(new_n842), .ZN(new_n843));
  OAI211_X1 g642(.A(KEYINPUT115), .B(new_n692), .C1(new_n837), .C2(new_n838), .ZN(new_n844));
  NAND3_X1  g643(.A1(new_n841), .A2(new_n843), .A3(new_n844), .ZN(new_n845));
  OAI21_X1  g644(.A(G113gat), .B1(new_n845), .B2(new_n571), .ZN(new_n846));
  NOR2_X1   g645(.A1(new_n823), .A2(new_n564), .ZN(new_n847));
  AOI21_X1  g646(.A(new_n828), .B1(new_n847), .B2(new_n563), .ZN(new_n848));
  AOI22_X1  g647(.A1(new_n570), .A2(new_n835), .B1(new_n848), .B2(new_n668), .ZN(new_n849));
  OAI21_X1  g648(.A(new_n836), .B1(new_n849), .B2(new_n645), .ZN(new_n850));
  AOI21_X1  g649(.A(new_n838), .B1(new_n850), .B2(new_n609), .ZN(new_n851));
  NOR2_X1   g650(.A1(new_n851), .A2(new_n437), .ZN(new_n852));
  NAND2_X1  g651(.A1(new_n852), .A2(new_n843), .ZN(new_n853));
  INV_X1    g652(.A(new_n853), .ZN(new_n854));
  NAND3_X1  g653(.A1(new_n854), .A2(new_n336), .A3(new_n570), .ZN(new_n855));
  NAND2_X1  g654(.A1(new_n846), .A2(new_n855), .ZN(G1340gat));
  OAI21_X1  g655(.A(G120gat), .B1(new_n845), .B2(new_n669), .ZN(new_n857));
  NAND3_X1  g656(.A1(new_n854), .A2(new_n334), .A3(new_n668), .ZN(new_n858));
  NAND2_X1  g657(.A1(new_n857), .A2(new_n858), .ZN(G1341gat));
  NOR3_X1   g658(.A1(new_n845), .A2(new_n327), .A3(new_n609), .ZN(new_n860));
  AOI21_X1  g659(.A(G127gat), .B1(new_n854), .B2(new_n608), .ZN(new_n861));
  NOR2_X1   g660(.A1(new_n860), .A2(new_n861), .ZN(G1342gat));
  NOR2_X1   g661(.A1(new_n702), .A2(new_n719), .ZN(new_n863));
  NAND4_X1  g662(.A1(new_n852), .A2(new_n325), .A3(new_n676), .A4(new_n863), .ZN(new_n864));
  XOR2_X1   g663(.A(KEYINPUT116), .B(KEYINPUT56), .Z(new_n865));
  XNOR2_X1  g664(.A(new_n864), .B(new_n865), .ZN(new_n866));
  OAI21_X1  g665(.A(G134gat), .B1(new_n845), .B2(new_n702), .ZN(new_n867));
  NAND2_X1  g666(.A1(new_n866), .A2(new_n867), .ZN(G1343gat));
  NOR2_X1   g667(.A1(new_n851), .A2(new_n401), .ZN(new_n869));
  NOR2_X1   g668(.A1(new_n675), .A2(new_n687), .ZN(new_n870));
  NAND2_X1  g669(.A1(new_n870), .A2(new_n453), .ZN(new_n871));
  INV_X1    g670(.A(new_n871), .ZN(new_n872));
  NAND2_X1  g671(.A1(new_n869), .A2(new_n872), .ZN(new_n873));
  NOR3_X1   g672(.A1(new_n873), .A2(G141gat), .A3(new_n571), .ZN(new_n874));
  OR2_X1    g673(.A1(new_n869), .A2(KEYINPUT57), .ZN(new_n875));
  NOR2_X1   g674(.A1(new_n811), .A2(new_n812), .ZN(new_n876));
  AOI21_X1  g675(.A(new_n829), .B1(new_n570), .B2(new_n876), .ZN(new_n877));
  OR2_X1    g676(.A1(new_n877), .A2(new_n645), .ZN(new_n878));
  AOI21_X1  g677(.A(new_n608), .B1(new_n878), .B2(new_n836), .ZN(new_n879));
  OAI211_X1 g678(.A(KEYINPUT57), .B(new_n458), .C1(new_n879), .C2(new_n838), .ZN(new_n880));
  AOI21_X1  g679(.A(new_n871), .B1(new_n875), .B2(new_n880), .ZN(new_n881));
  NAND2_X1  g680(.A1(new_n881), .A2(new_n570), .ZN(new_n882));
  AOI21_X1  g681(.A(new_n874), .B1(new_n882), .B2(G141gat), .ZN(new_n883));
  INV_X1    g682(.A(KEYINPUT58), .ZN(new_n884));
  XNOR2_X1  g683(.A(new_n883), .B(new_n884), .ZN(G1344gat));
  INV_X1    g684(.A(KEYINPUT59), .ZN(new_n886));
  OAI211_X1 g685(.A(KEYINPUT57), .B(new_n735), .C1(new_n837), .C2(new_n838), .ZN(new_n887));
  XNOR2_X1  g686(.A(new_n887), .B(KEYINPUT117), .ZN(new_n888));
  INV_X1    g687(.A(new_n838), .ZN(new_n889));
  NAND4_X1  g688(.A1(new_n645), .A2(new_n832), .A3(new_n834), .A4(new_n876), .ZN(new_n890));
  AOI21_X1  g689(.A(KEYINPUT118), .B1(new_n878), .B2(new_n890), .ZN(new_n891));
  OAI211_X1 g690(.A(KEYINPUT118), .B(new_n890), .C1(new_n877), .C2(new_n645), .ZN(new_n892));
  NAND2_X1  g691(.A1(new_n892), .A2(new_n609), .ZN(new_n893));
  OAI21_X1  g692(.A(new_n889), .B1(new_n891), .B2(new_n893), .ZN(new_n894));
  AOI21_X1  g693(.A(KEYINPUT57), .B1(new_n894), .B2(new_n458), .ZN(new_n895));
  OAI211_X1 g694(.A(new_n668), .B(new_n872), .C1(new_n888), .C2(new_n895), .ZN(new_n896));
  AOI21_X1  g695(.A(new_n886), .B1(new_n896), .B2(G148gat), .ZN(new_n897));
  AOI211_X1 g696(.A(KEYINPUT59), .B(new_n312), .C1(new_n881), .C2(new_n668), .ZN(new_n898));
  NAND2_X1  g697(.A1(new_n668), .A2(new_n312), .ZN(new_n899));
  OAI22_X1  g698(.A1(new_n897), .A2(new_n898), .B1(new_n873), .B2(new_n899), .ZN(G1345gat));
  NAND3_X1  g699(.A1(new_n881), .A2(G155gat), .A3(new_n608), .ZN(new_n901));
  NOR3_X1   g700(.A1(new_n873), .A2(KEYINPUT119), .A3(new_n609), .ZN(new_n902));
  OAI21_X1  g701(.A(KEYINPUT119), .B1(new_n873), .B2(new_n609), .ZN(new_n903));
  NAND2_X1  g702(.A1(new_n903), .A2(new_n316), .ZN(new_n904));
  OAI21_X1  g703(.A(new_n901), .B1(new_n902), .B2(new_n904), .ZN(new_n905));
  XNOR2_X1  g704(.A(new_n905), .B(KEYINPUT120), .ZN(G1346gat));
  NAND4_X1  g705(.A1(new_n869), .A2(new_n317), .A3(new_n863), .A4(new_n870), .ZN(new_n907));
  AND2_X1   g706(.A1(new_n881), .A2(new_n645), .ZN(new_n908));
  OAI21_X1  g707(.A(new_n907), .B1(new_n908), .B2(new_n317), .ZN(G1347gat));
  NAND2_X1  g708(.A1(new_n675), .A2(new_n719), .ZN(new_n910));
  NOR3_X1   g709(.A1(new_n851), .A2(new_n437), .A3(new_n910), .ZN(new_n911));
  INV_X1    g710(.A(new_n911), .ZN(new_n912));
  OR3_X1    g711(.A1(new_n912), .A2(G169gat), .A3(new_n571), .ZN(new_n913));
  OAI21_X1  g712(.A(new_n840), .B1(new_n851), .B2(new_n458), .ZN(new_n914));
  INV_X1    g713(.A(new_n910), .ZN(new_n915));
  NAND4_X1  g714(.A1(new_n914), .A2(new_n689), .A3(new_n844), .A4(new_n915), .ZN(new_n916));
  OAI21_X1  g715(.A(G169gat), .B1(new_n916), .B2(new_n571), .ZN(new_n917));
  NAND2_X1  g716(.A1(new_n913), .A2(new_n917), .ZN(G1348gat));
  INV_X1    g717(.A(G176gat), .ZN(new_n919));
  NOR3_X1   g718(.A1(new_n916), .A2(new_n919), .A3(new_n669), .ZN(new_n920));
  AOI21_X1  g719(.A(G176gat), .B1(new_n911), .B2(new_n668), .ZN(new_n921));
  NOR2_X1   g720(.A1(new_n920), .A2(new_n921), .ZN(G1349gat));
  OAI21_X1  g721(.A(G183gat), .B1(new_n916), .B2(new_n609), .ZN(new_n923));
  INV_X1    g722(.A(KEYINPUT121), .ZN(new_n924));
  OAI21_X1  g723(.A(new_n608), .B1(new_n245), .B2(new_n244), .ZN(new_n925));
  OAI211_X1 g724(.A(new_n923), .B(new_n924), .C1(new_n912), .C2(new_n925), .ZN(new_n926));
  XNOR2_X1  g725(.A(new_n926), .B(KEYINPUT60), .ZN(G1350gat));
  NAND3_X1  g726(.A1(new_n911), .A2(new_n229), .A3(new_n645), .ZN(new_n928));
  INV_X1    g727(.A(KEYINPUT123), .ZN(new_n929));
  NAND4_X1  g728(.A1(new_n841), .A2(new_n645), .A3(new_n844), .A4(new_n915), .ZN(new_n930));
  AND3_X1   g729(.A1(new_n930), .A2(KEYINPUT122), .A3(G190gat), .ZN(new_n931));
  AOI21_X1  g730(.A(KEYINPUT122), .B1(new_n930), .B2(G190gat), .ZN(new_n932));
  OAI211_X1 g731(.A(new_n929), .B(KEYINPUT61), .C1(new_n931), .C2(new_n932), .ZN(new_n933));
  OAI21_X1  g732(.A(G190gat), .B1(new_n916), .B2(new_n702), .ZN(new_n934));
  INV_X1    g733(.A(KEYINPUT122), .ZN(new_n935));
  NAND2_X1  g734(.A1(new_n934), .A2(new_n935), .ZN(new_n936));
  INV_X1    g735(.A(KEYINPUT61), .ZN(new_n937));
  NAND3_X1  g736(.A1(new_n930), .A2(KEYINPUT122), .A3(G190gat), .ZN(new_n938));
  NAND3_X1  g737(.A1(new_n936), .A2(new_n937), .A3(new_n938), .ZN(new_n939));
  NAND2_X1  g738(.A1(new_n933), .A2(new_n939), .ZN(new_n940));
  NAND2_X1  g739(.A1(new_n936), .A2(new_n938), .ZN(new_n941));
  AOI21_X1  g740(.A(new_n929), .B1(new_n941), .B2(KEYINPUT61), .ZN(new_n942));
  OAI21_X1  g741(.A(new_n928), .B1(new_n940), .B2(new_n942), .ZN(G1351gat));
  NOR2_X1   g742(.A1(new_n910), .A2(new_n687), .ZN(new_n944));
  NAND2_X1  g743(.A1(new_n869), .A2(new_n944), .ZN(new_n945));
  INV_X1    g744(.A(new_n945), .ZN(new_n946));
  INV_X1    g745(.A(G197gat), .ZN(new_n947));
  NAND3_X1  g746(.A1(new_n946), .A2(new_n947), .A3(new_n570), .ZN(new_n948));
  OAI211_X1 g747(.A(new_n570), .B(new_n944), .C1(new_n888), .C2(new_n895), .ZN(new_n949));
  INV_X1    g748(.A(new_n949), .ZN(new_n950));
  OAI21_X1  g749(.A(new_n948), .B1(new_n950), .B2(new_n947), .ZN(G1352gat));
  OAI211_X1 g750(.A(new_n668), .B(new_n944), .C1(new_n888), .C2(new_n895), .ZN(new_n952));
  NAND2_X1  g751(.A1(new_n952), .A2(G204gat), .ZN(new_n953));
  NAND2_X1  g752(.A1(new_n668), .A2(new_n205), .ZN(new_n954));
  NOR3_X1   g753(.A1(new_n945), .A2(KEYINPUT62), .A3(new_n954), .ZN(new_n955));
  OAI21_X1  g754(.A(KEYINPUT62), .B1(new_n945), .B2(new_n954), .ZN(new_n956));
  INV_X1    g755(.A(KEYINPUT124), .ZN(new_n957));
  NAND2_X1  g756(.A1(new_n956), .A2(new_n957), .ZN(new_n958));
  OAI211_X1 g757(.A(KEYINPUT124), .B(KEYINPUT62), .C1(new_n945), .C2(new_n954), .ZN(new_n959));
  AOI21_X1  g758(.A(new_n955), .B1(new_n958), .B2(new_n959), .ZN(new_n960));
  NAND2_X1  g759(.A1(new_n953), .A2(new_n960), .ZN(new_n961));
  NAND2_X1  g760(.A1(new_n961), .A2(KEYINPUT125), .ZN(new_n962));
  INV_X1    g761(.A(KEYINPUT125), .ZN(new_n963));
  NAND3_X1  g762(.A1(new_n953), .A2(new_n960), .A3(new_n963), .ZN(new_n964));
  NAND2_X1  g763(.A1(new_n962), .A2(new_n964), .ZN(G1353gat));
  NOR3_X1   g764(.A1(new_n945), .A2(G211gat), .A3(new_n609), .ZN(new_n966));
  XNOR2_X1  g765(.A(new_n966), .B(KEYINPUT126), .ZN(new_n967));
  OAI211_X1 g766(.A(new_n608), .B(new_n944), .C1(new_n888), .C2(new_n895), .ZN(new_n968));
  AND3_X1   g767(.A1(new_n968), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n969));
  AOI21_X1  g768(.A(KEYINPUT63), .B1(new_n968), .B2(G211gat), .ZN(new_n970));
  OAI21_X1  g769(.A(new_n967), .B1(new_n969), .B2(new_n970), .ZN(G1354gat));
  AOI21_X1  g770(.A(G218gat), .B1(new_n946), .B2(new_n645), .ZN(new_n972));
  NOR2_X1   g771(.A1(new_n888), .A2(new_n895), .ZN(new_n973));
  NOR3_X1   g772(.A1(new_n973), .A2(new_n687), .A3(new_n910), .ZN(new_n974));
  NOR3_X1   g773(.A1(new_n702), .A2(new_n209), .A3(new_n210), .ZN(new_n975));
  XNOR2_X1  g774(.A(new_n975), .B(KEYINPUT127), .ZN(new_n976));
  AOI21_X1  g775(.A(new_n972), .B1(new_n974), .B2(new_n976), .ZN(G1355gat));
endmodule


