//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 1 0 1 1 0 0 0 1 0 1 0 0 1 1 0 0 1 0 1 0 0 0 0 0 0 1 1 1 1 1 0 1 0 0 1 1 0 1 1 1 0 0 0 1 0 0 0 0 0 0 1 0 1 1 1 1 1 1 1 0 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:32:19 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n448, new_n449, new_n452, new_n453, new_n454, new_n457,
    new_n458, new_n459, new_n460, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n495, new_n496,
    new_n497, new_n498, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n518, new_n519,
    new_n520, new_n521, new_n522, new_n523, new_n524, new_n525, new_n528,
    new_n529, new_n530, new_n531, new_n532, new_n533, new_n534, new_n535,
    new_n536, new_n537, new_n538, new_n539, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n558, new_n559,
    new_n561, new_n562, new_n563, new_n564, new_n565, new_n566, new_n567,
    new_n568, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n578, new_n579, new_n580, new_n581, new_n582, new_n583, new_n584,
    new_n585, new_n586, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n611, new_n612, new_n613, new_n614, new_n615, new_n616,
    new_n617, new_n620, new_n622, new_n623, new_n624, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1213, new_n1214,
    new_n1215, new_n1217, new_n1218;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  XOR2_X1   g007(.A(KEYINPUT64), .B(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  XNOR2_X1  g013(.A(KEYINPUT65), .B(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  INV_X1    g022(.A(G567), .ZN(new_n448));
  NOR2_X1   g023(.A1(new_n446), .A2(new_n448), .ZN(new_n449));
  XOR2_X1   g024(.A(new_n449), .B(KEYINPUT66), .Z(G234));
  NAND3_X1  g025(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g026(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n452));
  XNOR2_X1  g027(.A(new_n452), .B(KEYINPUT2), .ZN(new_n453));
  NOR4_X1   g028(.A1(G236), .A2(G237), .A3(G235), .A4(G238), .ZN(new_n454));
  NAND2_X1  g029(.A1(new_n453), .A2(new_n454), .ZN(G261));
  INV_X1    g030(.A(G261), .ZN(G325));
  INV_X1    g031(.A(new_n453), .ZN(new_n457));
  NAND2_X1  g032(.A1(new_n457), .A2(G2106), .ZN(new_n458));
  OR2_X1    g033(.A1(new_n454), .A2(new_n448), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  INV_X1    g035(.A(new_n460), .ZN(G319));
  INV_X1    g036(.A(G2105), .ZN(new_n462));
  XNOR2_X1  g037(.A(KEYINPUT3), .B(G2104), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n463), .A2(G125), .ZN(new_n464));
  NAND2_X1  g039(.A1(G113), .A2(G2104), .ZN(new_n465));
  AOI21_X1  g040(.A(new_n462), .B1(new_n464), .B2(new_n465), .ZN(new_n466));
  NAND3_X1  g041(.A1(new_n463), .A2(G137), .A3(new_n462), .ZN(new_n467));
  INV_X1    g042(.A(G2104), .ZN(new_n468));
  NOR2_X1   g043(.A1(new_n468), .A2(G2105), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n469), .A2(G101), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n467), .A2(new_n470), .ZN(new_n471));
  NOR2_X1   g046(.A1(new_n466), .A2(new_n471), .ZN(G160));
  OR2_X1    g047(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n473));
  NAND2_X1  g048(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n474));
  AOI21_X1  g049(.A(G2105), .B1(new_n473), .B2(new_n474), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n475), .A2(G136), .ZN(new_n476));
  AOI21_X1  g051(.A(new_n462), .B1(new_n473), .B2(new_n474), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n477), .A2(G124), .ZN(new_n478));
  OR2_X1    g053(.A1(G100), .A2(G2105), .ZN(new_n479));
  OAI211_X1 g054(.A(new_n479), .B(G2104), .C1(G112), .C2(new_n462), .ZN(new_n480));
  NAND3_X1  g055(.A1(new_n476), .A2(new_n478), .A3(new_n480), .ZN(new_n481));
  INV_X1    g056(.A(new_n481), .ZN(G162));
  AND2_X1   g057(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n483));
  NOR2_X1   g058(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n484));
  OAI211_X1 g059(.A(G126), .B(G2105), .C1(new_n483), .C2(new_n484), .ZN(new_n485));
  INV_X1    g060(.A(G114), .ZN(new_n486));
  NAND2_X1  g061(.A1(new_n486), .A2(G2105), .ZN(new_n487));
  OAI211_X1 g062(.A(new_n487), .B(G2104), .C1(G102), .C2(G2105), .ZN(new_n488));
  NAND2_X1  g063(.A1(new_n485), .A2(new_n488), .ZN(new_n489));
  OAI211_X1 g064(.A(G138), .B(new_n462), .C1(new_n483), .C2(new_n484), .ZN(new_n490));
  NAND2_X1  g065(.A1(new_n490), .A2(KEYINPUT4), .ZN(new_n491));
  INV_X1    g066(.A(KEYINPUT4), .ZN(new_n492));
  NAND4_X1  g067(.A1(new_n463), .A2(new_n492), .A3(G138), .A4(new_n462), .ZN(new_n493));
  AOI21_X1  g068(.A(new_n489), .B1(new_n491), .B2(new_n493), .ZN(G164));
  INV_X1    g069(.A(KEYINPUT68), .ZN(new_n495));
  INV_X1    g070(.A(G651), .ZN(new_n496));
  OAI21_X1  g071(.A(new_n495), .B1(new_n496), .B2(KEYINPUT6), .ZN(new_n497));
  INV_X1    g072(.A(KEYINPUT6), .ZN(new_n498));
  NAND3_X1  g073(.A1(new_n498), .A2(KEYINPUT68), .A3(G651), .ZN(new_n499));
  AND2_X1   g074(.A1(new_n497), .A2(new_n499), .ZN(new_n500));
  NAND2_X1  g075(.A1(new_n496), .A2(KEYINPUT67), .ZN(new_n501));
  INV_X1    g076(.A(KEYINPUT67), .ZN(new_n502));
  NAND2_X1  g077(.A1(new_n502), .A2(G651), .ZN(new_n503));
  NAND3_X1  g078(.A1(new_n501), .A2(new_n503), .A3(KEYINPUT6), .ZN(new_n504));
  AND3_X1   g079(.A1(new_n500), .A2(G543), .A3(new_n504), .ZN(new_n505));
  NAND2_X1  g080(.A1(new_n505), .A2(G50), .ZN(new_n506));
  OR2_X1    g081(.A1(KEYINPUT5), .A2(G543), .ZN(new_n507));
  NAND2_X1  g082(.A1(KEYINPUT5), .A2(G543), .ZN(new_n508));
  NAND2_X1  g083(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  AND3_X1   g084(.A1(new_n500), .A2(new_n504), .A3(new_n509), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n510), .A2(G88), .ZN(new_n511));
  AOI22_X1  g086(.A1(new_n509), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n512));
  NAND2_X1  g087(.A1(new_n501), .A2(new_n503), .ZN(new_n513));
  INV_X1    g088(.A(new_n513), .ZN(new_n514));
  OR2_X1    g089(.A1(new_n512), .A2(new_n514), .ZN(new_n515));
  NAND3_X1  g090(.A1(new_n506), .A2(new_n511), .A3(new_n515), .ZN(G303));
  INV_X1    g091(.A(G303), .ZN(G166));
  NAND2_X1  g092(.A1(new_n505), .A2(G51), .ZN(new_n518));
  NAND2_X1  g093(.A1(new_n510), .A2(G89), .ZN(new_n519));
  NAND2_X1  g094(.A1(new_n509), .A2(G651), .ZN(new_n520));
  INV_X1    g095(.A(new_n520), .ZN(new_n521));
  NAND3_X1  g096(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n522));
  NAND2_X1  g097(.A1(new_n522), .A2(KEYINPUT7), .ZN(new_n523));
  OR2_X1    g098(.A1(new_n522), .A2(KEYINPUT7), .ZN(new_n524));
  AOI22_X1  g099(.A1(new_n521), .A2(G63), .B1(new_n523), .B2(new_n524), .ZN(new_n525));
  NAND3_X1  g100(.A1(new_n518), .A2(new_n519), .A3(new_n525), .ZN(G286));
  INV_X1    g101(.A(G286), .ZN(G168));
  NAND2_X1  g102(.A1(G77), .A2(G543), .ZN(new_n528));
  AND2_X1   g103(.A1(KEYINPUT5), .A2(G543), .ZN(new_n529));
  NOR2_X1   g104(.A1(KEYINPUT5), .A2(G543), .ZN(new_n530));
  NOR2_X1   g105(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  INV_X1    g106(.A(G64), .ZN(new_n532));
  OAI21_X1  g107(.A(new_n528), .B1(new_n531), .B2(new_n532), .ZN(new_n533));
  NAND2_X1  g108(.A1(new_n533), .A2(new_n513), .ZN(new_n534));
  NAND4_X1  g109(.A1(new_n500), .A2(G52), .A3(G543), .A4(new_n504), .ZN(new_n535));
  NAND3_X1  g110(.A1(new_n500), .A2(new_n504), .A3(new_n509), .ZN(new_n536));
  INV_X1    g111(.A(G90), .ZN(new_n537));
  OAI211_X1 g112(.A(new_n534), .B(new_n535), .C1(new_n536), .C2(new_n537), .ZN(new_n538));
  INV_X1    g113(.A(KEYINPUT69), .ZN(new_n539));
  XNOR2_X1  g114(.A(new_n538), .B(new_n539), .ZN(G171));
  NAND4_X1  g115(.A1(new_n500), .A2(G43), .A3(G543), .A4(new_n504), .ZN(new_n541));
  NAND4_X1  g116(.A1(new_n500), .A2(G81), .A3(new_n504), .A4(new_n509), .ZN(new_n542));
  NAND2_X1  g117(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  INV_X1    g118(.A(KEYINPUT71), .ZN(new_n544));
  NAND2_X1  g119(.A1(new_n543), .A2(new_n544), .ZN(new_n545));
  AND2_X1   g120(.A1(new_n509), .A2(G56), .ZN(new_n546));
  AND2_X1   g121(.A1(G68), .A2(G543), .ZN(new_n547));
  OAI211_X1 g122(.A(KEYINPUT70), .B(new_n513), .C1(new_n546), .C2(new_n547), .ZN(new_n548));
  INV_X1    g123(.A(KEYINPUT70), .ZN(new_n549));
  AOI21_X1  g124(.A(new_n547), .B1(new_n509), .B2(G56), .ZN(new_n550));
  OAI21_X1  g125(.A(new_n549), .B1(new_n550), .B2(new_n514), .ZN(new_n551));
  NAND2_X1  g126(.A1(new_n548), .A2(new_n551), .ZN(new_n552));
  NAND3_X1  g127(.A1(new_n541), .A2(new_n542), .A3(KEYINPUT71), .ZN(new_n553));
  NAND3_X1  g128(.A1(new_n545), .A2(new_n552), .A3(new_n553), .ZN(new_n554));
  INV_X1    g129(.A(new_n554), .ZN(new_n555));
  NAND2_X1  g130(.A1(new_n555), .A2(G860), .ZN(G153));
  NAND4_X1  g131(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g132(.A1(G1), .A2(G3), .ZN(new_n558));
  XNOR2_X1  g133(.A(new_n558), .B(KEYINPUT8), .ZN(new_n559));
  NAND4_X1  g134(.A1(G319), .A2(G483), .A3(G661), .A4(new_n559), .ZN(G188));
  NAND2_X1  g135(.A1(new_n509), .A2(G65), .ZN(new_n561));
  NAND2_X1  g136(.A1(G78), .A2(G543), .ZN(new_n562));
  AOI21_X1  g137(.A(new_n496), .B1(new_n561), .B2(new_n562), .ZN(new_n563));
  AOI21_X1  g138(.A(new_n563), .B1(new_n510), .B2(G91), .ZN(new_n564));
  NAND4_X1  g139(.A1(new_n500), .A2(G53), .A3(G543), .A4(new_n504), .ZN(new_n565));
  NAND2_X1  g140(.A1(new_n565), .A2(KEYINPUT9), .ZN(new_n566));
  INV_X1    g141(.A(new_n566), .ZN(new_n567));
  NOR2_X1   g142(.A1(new_n565), .A2(KEYINPUT9), .ZN(new_n568));
  OAI21_X1  g143(.A(new_n564), .B1(new_n567), .B2(new_n568), .ZN(G299));
  INV_X1    g144(.A(G171), .ZN(G301));
  NAND4_X1  g145(.A1(new_n500), .A2(G87), .A3(new_n504), .A4(new_n509), .ZN(new_n571));
  NAND4_X1  g146(.A1(new_n500), .A2(G49), .A3(G543), .A4(new_n504), .ZN(new_n572));
  NAND2_X1  g147(.A1(G74), .A2(G651), .ZN(new_n573));
  NAND3_X1  g148(.A1(new_n520), .A2(KEYINPUT72), .A3(new_n573), .ZN(new_n574));
  INV_X1    g149(.A(KEYINPUT72), .ZN(new_n575));
  OAI211_X1 g150(.A(new_n575), .B(G651), .C1(new_n509), .C2(G74), .ZN(new_n576));
  NAND4_X1  g151(.A1(new_n571), .A2(new_n572), .A3(new_n574), .A4(new_n576), .ZN(G288));
  NAND3_X1  g152(.A1(new_n509), .A2(KEYINPUT73), .A3(G61), .ZN(new_n578));
  INV_X1    g153(.A(new_n578), .ZN(new_n579));
  NAND2_X1  g154(.A1(G73), .A2(G543), .ZN(new_n580));
  INV_X1    g155(.A(G61), .ZN(new_n581));
  AOI21_X1  g156(.A(new_n581), .B1(new_n507), .B2(new_n508), .ZN(new_n582));
  OAI21_X1  g157(.A(new_n580), .B1(new_n582), .B2(KEYINPUT73), .ZN(new_n583));
  OAI21_X1  g158(.A(new_n513), .B1(new_n579), .B2(new_n583), .ZN(new_n584));
  NAND4_X1  g159(.A1(new_n500), .A2(G86), .A3(new_n504), .A4(new_n509), .ZN(new_n585));
  NAND4_X1  g160(.A1(new_n500), .A2(G48), .A3(G543), .A4(new_n504), .ZN(new_n586));
  NAND3_X1  g161(.A1(new_n584), .A2(new_n585), .A3(new_n586), .ZN(G305));
  NAND2_X1  g162(.A1(G72), .A2(G543), .ZN(new_n588));
  INV_X1    g163(.A(G60), .ZN(new_n589));
  OAI21_X1  g164(.A(new_n588), .B1(new_n531), .B2(new_n589), .ZN(new_n590));
  NAND2_X1  g165(.A1(new_n590), .A2(new_n513), .ZN(new_n591));
  NAND3_X1  g166(.A1(new_n500), .A2(G543), .A3(new_n504), .ZN(new_n592));
  INV_X1    g167(.A(G47), .ZN(new_n593));
  INV_X1    g168(.A(G85), .ZN(new_n594));
  OAI221_X1 g169(.A(new_n591), .B1(new_n592), .B2(new_n593), .C1(new_n594), .C2(new_n536), .ZN(G290));
  NAND2_X1  g170(.A1(G79), .A2(G543), .ZN(new_n596));
  INV_X1    g171(.A(G66), .ZN(new_n597));
  OAI21_X1  g172(.A(new_n596), .B1(new_n531), .B2(new_n597), .ZN(new_n598));
  NAND2_X1  g173(.A1(new_n598), .A2(G651), .ZN(new_n599));
  INV_X1    g174(.A(G54), .ZN(new_n600));
  OAI21_X1  g175(.A(new_n599), .B1(new_n592), .B2(new_n600), .ZN(new_n601));
  NAND3_X1  g176(.A1(new_n510), .A2(KEYINPUT10), .A3(G92), .ZN(new_n602));
  INV_X1    g177(.A(KEYINPUT10), .ZN(new_n603));
  INV_X1    g178(.A(G92), .ZN(new_n604));
  OAI21_X1  g179(.A(new_n603), .B1(new_n536), .B2(new_n604), .ZN(new_n605));
  AOI21_X1  g180(.A(new_n601), .B1(new_n602), .B2(new_n605), .ZN(new_n606));
  INV_X1    g181(.A(new_n606), .ZN(new_n607));
  NOR2_X1   g182(.A1(new_n607), .A2(G868), .ZN(new_n608));
  AOI21_X1  g183(.A(new_n608), .B1(G868), .B2(G171), .ZN(G284));
  AOI21_X1  g184(.A(new_n608), .B1(G868), .B2(G171), .ZN(G321));
  NAND2_X1  g185(.A1(G286), .A2(G868), .ZN(new_n611));
  INV_X1    g186(.A(G91), .ZN(new_n612));
  AOI22_X1  g187(.A1(new_n509), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n613));
  OAI22_X1  g188(.A1(new_n536), .A2(new_n612), .B1(new_n613), .B2(new_n496), .ZN(new_n614));
  INV_X1    g189(.A(KEYINPUT9), .ZN(new_n615));
  NAND3_X1  g190(.A1(new_n505), .A2(new_n615), .A3(G53), .ZN(new_n616));
  AOI21_X1  g191(.A(new_n614), .B1(new_n616), .B2(new_n566), .ZN(new_n617));
  OAI21_X1  g192(.A(new_n611), .B1(G868), .B2(new_n617), .ZN(G297));
  OAI21_X1  g193(.A(new_n611), .B1(G868), .B2(new_n617), .ZN(G280));
  INV_X1    g194(.A(G559), .ZN(new_n620));
  OAI21_X1  g195(.A(new_n606), .B1(new_n620), .B2(G860), .ZN(G148));
  NAND2_X1  g196(.A1(new_n606), .A2(new_n620), .ZN(new_n622));
  NAND2_X1  g197(.A1(new_n622), .A2(G868), .ZN(new_n623));
  OAI21_X1  g198(.A(new_n623), .B1(G868), .B2(new_n555), .ZN(new_n624));
  XOR2_X1   g199(.A(new_n624), .B(KEYINPUT74), .Z(G323));
  XNOR2_X1  g200(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NOR2_X1   g201(.A1(new_n483), .A2(new_n484), .ZN(new_n627));
  INV_X1    g202(.A(new_n469), .ZN(new_n628));
  NOR2_X1   g203(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  XNOR2_X1  g204(.A(KEYINPUT75), .B(KEYINPUT12), .ZN(new_n630));
  XOR2_X1   g205(.A(new_n629), .B(new_n630), .Z(new_n631));
  XOR2_X1   g206(.A(new_n631), .B(KEYINPUT13), .Z(new_n632));
  OR2_X1    g207(.A1(new_n632), .A2(G2100), .ZN(new_n633));
  NAND2_X1  g208(.A1(new_n632), .A2(G2100), .ZN(new_n634));
  NAND2_X1  g209(.A1(new_n475), .A2(G135), .ZN(new_n635));
  NAND2_X1  g210(.A1(new_n477), .A2(G123), .ZN(new_n636));
  NOR2_X1   g211(.A1(new_n462), .A2(G111), .ZN(new_n637));
  OAI21_X1  g212(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n638));
  OAI211_X1 g213(.A(new_n635), .B(new_n636), .C1(new_n637), .C2(new_n638), .ZN(new_n639));
  XOR2_X1   g214(.A(new_n639), .B(G2096), .Z(new_n640));
  NAND3_X1  g215(.A1(new_n633), .A2(new_n634), .A3(new_n640), .ZN(G156));
  XNOR2_X1  g216(.A(G2427), .B(G2438), .ZN(new_n642));
  XNOR2_X1  g217(.A(new_n642), .B(G2430), .ZN(new_n643));
  XNOR2_X1  g218(.A(KEYINPUT15), .B(G2435), .ZN(new_n644));
  OR2_X1    g219(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  NAND2_X1  g220(.A1(new_n643), .A2(new_n644), .ZN(new_n646));
  NAND3_X1  g221(.A1(new_n645), .A2(KEYINPUT14), .A3(new_n646), .ZN(new_n647));
  XNOR2_X1  g222(.A(G2443), .B(G2446), .ZN(new_n648));
  XNOR2_X1  g223(.A(new_n647), .B(new_n648), .ZN(new_n649));
  XOR2_X1   g224(.A(G2451), .B(G2454), .Z(new_n650));
  XNOR2_X1  g225(.A(new_n650), .B(KEYINPUT16), .ZN(new_n651));
  XNOR2_X1  g226(.A(new_n651), .B(KEYINPUT76), .ZN(new_n652));
  XNOR2_X1  g227(.A(new_n649), .B(new_n652), .ZN(new_n653));
  XOR2_X1   g228(.A(G1341), .B(G1348), .Z(new_n654));
  XNOR2_X1  g229(.A(new_n654), .B(KEYINPUT77), .ZN(new_n655));
  NAND2_X1  g230(.A1(new_n653), .A2(new_n655), .ZN(new_n656));
  XOR2_X1   g231(.A(new_n656), .B(KEYINPUT78), .Z(new_n657));
  OAI21_X1  g232(.A(G14), .B1(new_n653), .B2(new_n655), .ZN(new_n658));
  NOR2_X1   g233(.A1(new_n657), .A2(new_n658), .ZN(G401));
  XNOR2_X1  g234(.A(G2072), .B(G2078), .ZN(new_n660));
  XNOR2_X1  g235(.A(new_n660), .B(KEYINPUT17), .ZN(new_n661));
  XNOR2_X1  g236(.A(G2067), .B(G2678), .ZN(new_n662));
  XNOR2_X1  g237(.A(new_n662), .B(KEYINPUT79), .ZN(new_n663));
  XOR2_X1   g238(.A(G2084), .B(G2090), .Z(new_n664));
  INV_X1    g239(.A(new_n664), .ZN(new_n665));
  NOR3_X1   g240(.A1(new_n661), .A2(new_n663), .A3(new_n665), .ZN(new_n666));
  XNOR2_X1  g241(.A(new_n666), .B(KEYINPUT80), .ZN(new_n667));
  AOI21_X1  g242(.A(new_n664), .B1(new_n661), .B2(new_n663), .ZN(new_n668));
  OAI21_X1  g243(.A(new_n668), .B1(new_n660), .B2(new_n663), .ZN(new_n669));
  NAND3_X1  g244(.A1(new_n664), .A2(new_n660), .A3(new_n662), .ZN(new_n670));
  XOR2_X1   g245(.A(new_n670), .B(KEYINPUT18), .Z(new_n671));
  NAND3_X1  g246(.A1(new_n667), .A2(new_n669), .A3(new_n671), .ZN(new_n672));
  XOR2_X1   g247(.A(G2096), .B(G2100), .Z(new_n673));
  XNOR2_X1  g248(.A(new_n672), .B(new_n673), .ZN(G227));
  XNOR2_X1  g249(.A(G1971), .B(G1976), .ZN(new_n675));
  XNOR2_X1  g250(.A(KEYINPUT81), .B(KEYINPUT19), .ZN(new_n676));
  XNOR2_X1  g251(.A(new_n675), .B(new_n676), .ZN(new_n677));
  XNOR2_X1  g252(.A(G1956), .B(G2474), .ZN(new_n678));
  INV_X1    g253(.A(new_n678), .ZN(new_n679));
  XNOR2_X1  g254(.A(G1961), .B(G1966), .ZN(new_n680));
  INV_X1    g255(.A(new_n680), .ZN(new_n681));
  NAND3_X1  g256(.A1(new_n677), .A2(new_n679), .A3(new_n681), .ZN(new_n682));
  XOR2_X1   g257(.A(KEYINPUT82), .B(KEYINPUT20), .Z(new_n683));
  OR2_X1    g258(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  NAND2_X1  g259(.A1(new_n682), .A2(new_n683), .ZN(new_n685));
  NAND3_X1  g260(.A1(new_n677), .A2(new_n678), .A3(new_n680), .ZN(new_n686));
  XNOR2_X1  g261(.A(new_n678), .B(new_n680), .ZN(new_n687));
  OR2_X1    g262(.A1(new_n687), .A2(new_n677), .ZN(new_n688));
  NAND4_X1  g263(.A1(new_n684), .A2(new_n685), .A3(new_n686), .A4(new_n688), .ZN(new_n689));
  XOR2_X1   g264(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n690));
  XNOR2_X1  g265(.A(new_n689), .B(new_n690), .ZN(new_n691));
  XNOR2_X1  g266(.A(G1991), .B(G1996), .ZN(new_n692));
  XNOR2_X1  g267(.A(new_n691), .B(new_n692), .ZN(new_n693));
  XNOR2_X1  g268(.A(G1981), .B(G1986), .ZN(new_n694));
  XNOR2_X1  g269(.A(new_n693), .B(new_n694), .ZN(new_n695));
  INV_X1    g270(.A(new_n695), .ZN(G229));
  INV_X1    g271(.A(G29), .ZN(new_n697));
  INV_X1    g272(.A(G127), .ZN(new_n698));
  INV_X1    g273(.A(G115), .ZN(new_n699));
  OAI22_X1  g274(.A1(new_n627), .A2(new_n698), .B1(new_n699), .B2(new_n468), .ZN(new_n700));
  NAND2_X1  g275(.A1(new_n700), .A2(KEYINPUT89), .ZN(new_n701));
  INV_X1    g276(.A(KEYINPUT89), .ZN(new_n702));
  OAI221_X1 g277(.A(new_n702), .B1(new_n699), .B2(new_n468), .C1(new_n627), .C2(new_n698), .ZN(new_n703));
  NAND3_X1  g278(.A1(new_n701), .A2(G2105), .A3(new_n703), .ZN(new_n704));
  NAND3_X1  g279(.A1(new_n462), .A2(G103), .A3(G2104), .ZN(new_n705));
  XNOR2_X1  g280(.A(new_n705), .B(KEYINPUT25), .ZN(new_n706));
  AOI21_X1  g281(.A(new_n706), .B1(G139), .B2(new_n475), .ZN(new_n707));
  NAND2_X1  g282(.A1(new_n704), .A2(new_n707), .ZN(new_n708));
  INV_X1    g283(.A(KEYINPUT90), .ZN(new_n709));
  NAND2_X1  g284(.A1(new_n708), .A2(new_n709), .ZN(new_n710));
  NAND3_X1  g285(.A1(new_n704), .A2(KEYINPUT90), .A3(new_n707), .ZN(new_n711));
  NAND2_X1  g286(.A1(new_n710), .A2(new_n711), .ZN(new_n712));
  NAND2_X1  g287(.A1(new_n712), .A2(KEYINPUT91), .ZN(new_n713));
  INV_X1    g288(.A(KEYINPUT91), .ZN(new_n714));
  NAND3_X1  g289(.A1(new_n710), .A2(new_n714), .A3(new_n711), .ZN(new_n715));
  AOI21_X1  g290(.A(new_n697), .B1(new_n713), .B2(new_n715), .ZN(new_n716));
  AOI21_X1  g291(.A(new_n716), .B1(new_n697), .B2(G33), .ZN(new_n717));
  INV_X1    g292(.A(G2072), .ZN(new_n718));
  NOR2_X1   g293(.A1(new_n717), .A2(new_n718), .ZN(new_n719));
  XOR2_X1   g294(.A(new_n719), .B(KEYINPUT92), .Z(new_n720));
  NOR2_X1   g295(.A1(G29), .A2(G32), .ZN(new_n721));
  AOI22_X1  g296(.A1(G129), .A2(new_n477), .B1(new_n475), .B2(G141), .ZN(new_n722));
  XNOR2_X1  g297(.A(KEYINPUT93), .B(KEYINPUT26), .ZN(new_n723));
  AND3_X1   g298(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n724));
  XNOR2_X1  g299(.A(new_n723), .B(new_n724), .ZN(new_n725));
  NAND2_X1  g300(.A1(new_n469), .A2(G105), .ZN(new_n726));
  NAND3_X1  g301(.A1(new_n722), .A2(new_n725), .A3(new_n726), .ZN(new_n727));
  AND2_X1   g302(.A1(new_n727), .A2(KEYINPUT94), .ZN(new_n728));
  NOR2_X1   g303(.A1(new_n727), .A2(KEYINPUT94), .ZN(new_n729));
  NOR2_X1   g304(.A1(new_n728), .A2(new_n729), .ZN(new_n730));
  AOI21_X1  g305(.A(new_n721), .B1(new_n730), .B2(G29), .ZN(new_n731));
  XOR2_X1   g306(.A(KEYINPUT27), .B(G1996), .Z(new_n732));
  XNOR2_X1  g307(.A(new_n731), .B(new_n732), .ZN(new_n733));
  XNOR2_X1  g308(.A(KEYINPUT30), .B(G28), .ZN(new_n734));
  OR2_X1    g309(.A1(KEYINPUT31), .A2(G11), .ZN(new_n735));
  NAND2_X1  g310(.A1(KEYINPUT31), .A2(G11), .ZN(new_n736));
  AOI22_X1  g311(.A1(new_n734), .A2(new_n697), .B1(new_n735), .B2(new_n736), .ZN(new_n737));
  OAI21_X1  g312(.A(new_n737), .B1(new_n639), .B2(new_n697), .ZN(new_n738));
  INV_X1    g313(.A(KEYINPUT24), .ZN(new_n739));
  OAI21_X1  g314(.A(new_n697), .B1(new_n739), .B2(G34), .ZN(new_n740));
  AOI21_X1  g315(.A(new_n740), .B1(new_n739), .B2(G34), .ZN(new_n741));
  AOI21_X1  g316(.A(new_n741), .B1(G160), .B2(G29), .ZN(new_n742));
  AOI21_X1  g317(.A(new_n738), .B1(new_n742), .B2(G2084), .ZN(new_n743));
  OAI21_X1  g318(.A(new_n743), .B1(G2084), .B2(new_n742), .ZN(new_n744));
  NAND2_X1  g319(.A1(new_n697), .A2(G27), .ZN(new_n745));
  XOR2_X1   g320(.A(new_n745), .B(KEYINPUT95), .Z(new_n746));
  AND2_X1   g321(.A1(new_n485), .A2(new_n488), .ZN(new_n747));
  AOI21_X1  g322(.A(new_n492), .B1(new_n475), .B2(G138), .ZN(new_n748));
  NOR2_X1   g323(.A1(new_n490), .A2(KEYINPUT4), .ZN(new_n749));
  OAI21_X1  g324(.A(new_n747), .B1(new_n748), .B2(new_n749), .ZN(new_n750));
  AOI21_X1  g325(.A(new_n746), .B1(new_n750), .B2(G29), .ZN(new_n751));
  INV_X1    g326(.A(G2078), .ZN(new_n752));
  XNOR2_X1  g327(.A(new_n751), .B(new_n752), .ZN(new_n753));
  NOR3_X1   g328(.A1(new_n733), .A2(new_n744), .A3(new_n753), .ZN(new_n754));
  NAND2_X1  g329(.A1(new_n717), .A2(new_n718), .ZN(new_n755));
  INV_X1    g330(.A(G16), .ZN(new_n756));
  NAND2_X1  g331(.A1(new_n756), .A2(G21), .ZN(new_n757));
  OAI21_X1  g332(.A(new_n757), .B1(G168), .B2(new_n756), .ZN(new_n758));
  AND2_X1   g333(.A1(new_n758), .A2(G1966), .ZN(new_n759));
  XNOR2_X1  g334(.A(KEYINPUT88), .B(KEYINPUT28), .ZN(new_n760));
  NAND2_X1  g335(.A1(new_n697), .A2(G26), .ZN(new_n761));
  XNOR2_X1  g336(.A(new_n760), .B(new_n761), .ZN(new_n762));
  NAND2_X1  g337(.A1(new_n477), .A2(G128), .ZN(new_n763));
  INV_X1    g338(.A(KEYINPUT87), .ZN(new_n764));
  NAND2_X1  g339(.A1(new_n763), .A2(new_n764), .ZN(new_n765));
  NAND3_X1  g340(.A1(new_n477), .A2(KEYINPUT87), .A3(G128), .ZN(new_n766));
  NAND2_X1  g341(.A1(new_n765), .A2(new_n766), .ZN(new_n767));
  NOR2_X1   g342(.A1(new_n462), .A2(G116), .ZN(new_n768));
  OAI21_X1  g343(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n769));
  OR2_X1    g344(.A1(new_n768), .A2(new_n769), .ZN(new_n770));
  NAND2_X1  g345(.A1(new_n475), .A2(G140), .ZN(new_n771));
  NAND3_X1  g346(.A1(new_n767), .A2(new_n770), .A3(new_n771), .ZN(new_n772));
  AOI21_X1  g347(.A(new_n762), .B1(new_n772), .B2(G29), .ZN(new_n773));
  INV_X1    g348(.A(G2067), .ZN(new_n774));
  XNOR2_X1  g349(.A(new_n773), .B(new_n774), .ZN(new_n775));
  NOR2_X1   g350(.A1(new_n758), .A2(G1966), .ZN(new_n776));
  NOR3_X1   g351(.A1(new_n759), .A2(new_n775), .A3(new_n776), .ZN(new_n777));
  INV_X1    g352(.A(G19), .ZN(new_n778));
  OR3_X1    g353(.A1(new_n778), .A2(KEYINPUT85), .A3(G16), .ZN(new_n779));
  OAI21_X1  g354(.A(KEYINPUT85), .B1(new_n778), .B2(G16), .ZN(new_n780));
  OAI211_X1 g355(.A(new_n779), .B(new_n780), .C1(new_n555), .C2(new_n756), .ZN(new_n781));
  XNOR2_X1  g356(.A(KEYINPUT86), .B(G1341), .ZN(new_n782));
  XNOR2_X1  g357(.A(new_n781), .B(new_n782), .ZN(new_n783));
  NAND4_X1  g358(.A1(new_n754), .A2(new_n755), .A3(new_n777), .A4(new_n783), .ZN(new_n784));
  NAND2_X1  g359(.A1(new_n697), .A2(G35), .ZN(new_n785));
  OAI21_X1  g360(.A(new_n785), .B1(G162), .B2(new_n697), .ZN(new_n786));
  XOR2_X1   g361(.A(new_n786), .B(KEYINPUT29), .Z(new_n787));
  INV_X1    g362(.A(G2090), .ZN(new_n788));
  NAND2_X1  g363(.A1(new_n787), .A2(new_n788), .ZN(new_n789));
  XNOR2_X1  g364(.A(new_n789), .B(KEYINPUT96), .ZN(new_n790));
  OR2_X1    g365(.A1(new_n787), .A2(new_n788), .ZN(new_n791));
  INV_X1    g366(.A(KEYINPUT97), .ZN(new_n792));
  INV_X1    g367(.A(G1348), .ZN(new_n793));
  NOR2_X1   g368(.A1(new_n606), .A2(new_n756), .ZN(new_n794));
  AOI21_X1  g369(.A(new_n794), .B1(G4), .B2(new_n756), .ZN(new_n795));
  OAI22_X1  g370(.A1(new_n791), .A2(new_n792), .B1(new_n793), .B2(new_n795), .ZN(new_n796));
  OR2_X1    g371(.A1(new_n790), .A2(new_n796), .ZN(new_n797));
  NOR2_X1   g372(.A1(G5), .A2(G16), .ZN(new_n798));
  AOI21_X1  g373(.A(new_n798), .B1(G171), .B2(G16), .ZN(new_n799));
  XNOR2_X1  g374(.A(new_n799), .B(G1961), .ZN(new_n800));
  NAND2_X1  g375(.A1(new_n791), .A2(new_n792), .ZN(new_n801));
  NAND2_X1  g376(.A1(new_n795), .A2(new_n793), .ZN(new_n802));
  NAND2_X1  g377(.A1(new_n756), .A2(G20), .ZN(new_n803));
  XOR2_X1   g378(.A(new_n803), .B(KEYINPUT23), .Z(new_n804));
  AOI21_X1  g379(.A(new_n804), .B1(G299), .B2(G16), .ZN(new_n805));
  XNOR2_X1  g380(.A(new_n805), .B(G1956), .ZN(new_n806));
  NAND3_X1  g381(.A1(new_n801), .A2(new_n802), .A3(new_n806), .ZN(new_n807));
  NOR4_X1   g382(.A1(new_n784), .A2(new_n797), .A3(new_n800), .A4(new_n807), .ZN(new_n808));
  NAND2_X1  g383(.A1(new_n756), .A2(G22), .ZN(new_n809));
  OAI21_X1  g384(.A(new_n809), .B1(G166), .B2(new_n756), .ZN(new_n810));
  INV_X1    g385(.A(G1971), .ZN(new_n811));
  XNOR2_X1  g386(.A(new_n810), .B(new_n811), .ZN(new_n812));
  NOR2_X1   g387(.A1(G6), .A2(G16), .ZN(new_n813));
  NAND2_X1  g388(.A1(new_n585), .A2(new_n586), .ZN(new_n814));
  OAI21_X1  g389(.A(G61), .B1(new_n529), .B2(new_n530), .ZN(new_n815));
  INV_X1    g390(.A(KEYINPUT73), .ZN(new_n816));
  AOI22_X1  g391(.A1(new_n815), .A2(new_n816), .B1(G73), .B2(G543), .ZN(new_n817));
  AOI21_X1  g392(.A(new_n514), .B1(new_n817), .B2(new_n578), .ZN(new_n818));
  NOR2_X1   g393(.A1(new_n814), .A2(new_n818), .ZN(new_n819));
  AOI21_X1  g394(.A(new_n813), .B1(new_n819), .B2(G16), .ZN(new_n820));
  XOR2_X1   g395(.A(KEYINPUT32), .B(G1981), .Z(new_n821));
  XNOR2_X1  g396(.A(new_n820), .B(new_n821), .ZN(new_n822));
  NAND2_X1  g397(.A1(new_n756), .A2(G23), .ZN(new_n823));
  INV_X1    g398(.A(G288), .ZN(new_n824));
  OAI21_X1  g399(.A(new_n823), .B1(new_n824), .B2(new_n756), .ZN(new_n825));
  XNOR2_X1  g400(.A(KEYINPUT33), .B(G1976), .ZN(new_n826));
  XNOR2_X1  g401(.A(new_n825), .B(new_n826), .ZN(new_n827));
  NAND3_X1  g402(.A1(new_n812), .A2(new_n822), .A3(new_n827), .ZN(new_n828));
  XOR2_X1   g403(.A(new_n828), .B(KEYINPUT34), .Z(new_n829));
  NAND2_X1  g404(.A1(new_n697), .A2(G25), .ZN(new_n830));
  INV_X1    g405(.A(G95), .ZN(new_n831));
  AND3_X1   g406(.A1(new_n831), .A2(new_n462), .A3(KEYINPUT83), .ZN(new_n832));
  AOI21_X1  g407(.A(KEYINPUT83), .B1(new_n831), .B2(new_n462), .ZN(new_n833));
  OAI221_X1 g408(.A(G2104), .B1(G107), .B2(new_n462), .C1(new_n832), .C2(new_n833), .ZN(new_n834));
  NAND2_X1  g409(.A1(new_n475), .A2(G131), .ZN(new_n835));
  NAND2_X1  g410(.A1(new_n477), .A2(G119), .ZN(new_n836));
  NAND3_X1  g411(.A1(new_n834), .A2(new_n835), .A3(new_n836), .ZN(new_n837));
  INV_X1    g412(.A(new_n837), .ZN(new_n838));
  OAI21_X1  g413(.A(new_n830), .B1(new_n838), .B2(new_n697), .ZN(new_n839));
  XOR2_X1   g414(.A(KEYINPUT35), .B(G1991), .Z(new_n840));
  XNOR2_X1  g415(.A(new_n840), .B(KEYINPUT84), .ZN(new_n841));
  XNOR2_X1  g416(.A(new_n839), .B(new_n841), .ZN(new_n842));
  MUX2_X1   g417(.A(G24), .B(G290), .S(G16), .Z(new_n843));
  XOR2_X1   g418(.A(new_n843), .B(G1986), .Z(new_n844));
  NAND3_X1  g419(.A1(new_n829), .A2(new_n842), .A3(new_n844), .ZN(new_n845));
  AND2_X1   g420(.A1(new_n845), .A2(KEYINPUT36), .ZN(new_n846));
  NOR2_X1   g421(.A1(new_n845), .A2(KEYINPUT36), .ZN(new_n847));
  OAI211_X1 g422(.A(new_n720), .B(new_n808), .C1(new_n846), .C2(new_n847), .ZN(G150));
  INV_X1    g423(.A(G150), .ZN(G311));
  NAND2_X1  g424(.A1(new_n606), .A2(G559), .ZN(new_n850));
  XOR2_X1   g425(.A(KEYINPUT98), .B(KEYINPUT38), .Z(new_n851));
  XNOR2_X1  g426(.A(new_n850), .B(new_n851), .ZN(new_n852));
  XOR2_X1   g427(.A(KEYINPUT99), .B(G55), .Z(new_n853));
  NAND4_X1  g428(.A1(new_n500), .A2(G543), .A3(new_n504), .A4(new_n853), .ZN(new_n854));
  NAND2_X1  g429(.A1(G80), .A2(G543), .ZN(new_n855));
  INV_X1    g430(.A(G67), .ZN(new_n856));
  OAI21_X1  g431(.A(new_n855), .B1(new_n531), .B2(new_n856), .ZN(new_n857));
  NAND2_X1  g432(.A1(new_n857), .A2(new_n513), .ZN(new_n858));
  NAND4_X1  g433(.A1(new_n500), .A2(G93), .A3(new_n504), .A4(new_n509), .ZN(new_n859));
  NAND3_X1  g434(.A1(new_n854), .A2(new_n858), .A3(new_n859), .ZN(new_n860));
  NAND2_X1  g435(.A1(new_n554), .A2(new_n860), .ZN(new_n861));
  INV_X1    g436(.A(new_n860), .ZN(new_n862));
  NAND4_X1  g437(.A1(new_n862), .A2(new_n545), .A3(new_n552), .A4(new_n553), .ZN(new_n863));
  NAND2_X1  g438(.A1(new_n861), .A2(new_n863), .ZN(new_n864));
  INV_X1    g439(.A(new_n864), .ZN(new_n865));
  XNOR2_X1  g440(.A(new_n852), .B(new_n865), .ZN(new_n866));
  AND2_X1   g441(.A1(new_n866), .A2(KEYINPUT39), .ZN(new_n867));
  NOR2_X1   g442(.A1(new_n866), .A2(KEYINPUT39), .ZN(new_n868));
  NOR3_X1   g443(.A1(new_n867), .A2(new_n868), .A3(G860), .ZN(new_n869));
  NAND2_X1  g444(.A1(new_n860), .A2(G860), .ZN(new_n870));
  XNOR2_X1  g445(.A(new_n870), .B(KEYINPUT37), .ZN(new_n871));
  OR2_X1    g446(.A1(new_n869), .A2(new_n871), .ZN(G145));
  AOI22_X1  g447(.A1(G130), .A2(new_n477), .B1(new_n475), .B2(G142), .ZN(new_n873));
  OAI21_X1  g448(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n874));
  INV_X1    g449(.A(G118), .ZN(new_n875));
  AOI22_X1  g450(.A1(new_n874), .A2(KEYINPUT101), .B1(new_n875), .B2(G2105), .ZN(new_n876));
  OAI21_X1  g451(.A(new_n876), .B1(KEYINPUT101), .B2(new_n874), .ZN(new_n877));
  NAND2_X1  g452(.A1(new_n873), .A2(new_n877), .ZN(new_n878));
  XNOR2_X1  g453(.A(new_n878), .B(new_n837), .ZN(new_n879));
  INV_X1    g454(.A(new_n879), .ZN(new_n880));
  NAND2_X1  g455(.A1(new_n772), .A2(G164), .ZN(new_n881));
  NAND4_X1  g456(.A1(new_n750), .A2(new_n767), .A3(new_n770), .A4(new_n771), .ZN(new_n882));
  NAND2_X1  g457(.A1(new_n881), .A2(new_n882), .ZN(new_n883));
  NAND2_X1  g458(.A1(new_n883), .A2(new_n730), .ZN(new_n884));
  OAI211_X1 g459(.A(new_n881), .B(new_n882), .C1(new_n728), .C2(new_n729), .ZN(new_n885));
  NAND4_X1  g460(.A1(new_n713), .A2(new_n884), .A3(new_n715), .A4(new_n885), .ZN(new_n886));
  INV_X1    g461(.A(new_n631), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n883), .A2(new_n727), .ZN(new_n888));
  INV_X1    g463(.A(new_n727), .ZN(new_n889));
  NAND3_X1  g464(.A1(new_n881), .A2(new_n889), .A3(new_n882), .ZN(new_n890));
  NAND3_X1  g465(.A1(new_n888), .A2(new_n712), .A3(new_n890), .ZN(new_n891));
  NAND3_X1  g466(.A1(new_n886), .A2(new_n887), .A3(new_n891), .ZN(new_n892));
  INV_X1    g467(.A(new_n892), .ZN(new_n893));
  AOI21_X1  g468(.A(new_n887), .B1(new_n886), .B2(new_n891), .ZN(new_n894));
  OAI21_X1  g469(.A(new_n880), .B1(new_n893), .B2(new_n894), .ZN(new_n895));
  INV_X1    g470(.A(new_n894), .ZN(new_n896));
  NAND3_X1  g471(.A1(new_n896), .A2(new_n879), .A3(new_n892), .ZN(new_n897));
  XNOR2_X1  g472(.A(G160), .B(new_n481), .ZN(new_n898));
  XNOR2_X1  g473(.A(new_n898), .B(KEYINPUT100), .ZN(new_n899));
  XOR2_X1   g474(.A(new_n899), .B(new_n639), .Z(new_n900));
  NAND3_X1  g475(.A1(new_n895), .A2(new_n897), .A3(new_n900), .ZN(new_n901));
  INV_X1    g476(.A(G37), .ZN(new_n902));
  AND2_X1   g477(.A1(new_n901), .A2(new_n902), .ZN(new_n903));
  AOI21_X1  g478(.A(new_n900), .B1(new_n895), .B2(new_n897), .ZN(new_n904));
  NOR2_X1   g479(.A1(new_n904), .A2(KEYINPUT102), .ZN(new_n905));
  INV_X1    g480(.A(KEYINPUT102), .ZN(new_n906));
  AOI211_X1 g481(.A(new_n906), .B(new_n900), .C1(new_n895), .C2(new_n897), .ZN(new_n907));
  OAI21_X1  g482(.A(new_n903), .B1(new_n905), .B2(new_n907), .ZN(new_n908));
  XNOR2_X1  g483(.A(KEYINPUT103), .B(KEYINPUT40), .ZN(new_n909));
  XNOR2_X1  g484(.A(new_n908), .B(new_n909), .ZN(G395));
  NOR2_X1   g485(.A1(new_n860), .A2(G868), .ZN(new_n911));
  INV_X1    g486(.A(KEYINPUT105), .ZN(new_n912));
  XNOR2_X1  g487(.A(G290), .B(new_n912), .ZN(new_n913));
  OR2_X1    g488(.A1(new_n913), .A2(new_n824), .ZN(new_n914));
  NAND2_X1  g489(.A1(new_n913), .A2(new_n824), .ZN(new_n915));
  NAND2_X1  g490(.A1(new_n914), .A2(new_n915), .ZN(new_n916));
  XNOR2_X1  g491(.A(G303), .B(G305), .ZN(new_n917));
  INV_X1    g492(.A(new_n917), .ZN(new_n918));
  NAND2_X1  g493(.A1(new_n916), .A2(new_n918), .ZN(new_n919));
  NAND3_X1  g494(.A1(new_n914), .A2(new_n917), .A3(new_n915), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  XNOR2_X1  g496(.A(new_n921), .B(KEYINPUT42), .ZN(new_n922));
  XOR2_X1   g497(.A(new_n864), .B(new_n622), .Z(new_n923));
  INV_X1    g498(.A(KEYINPUT41), .ZN(new_n924));
  INV_X1    g499(.A(KEYINPUT104), .ZN(new_n925));
  OAI211_X1 g500(.A(new_n564), .B(new_n925), .C1(new_n567), .C2(new_n568), .ZN(new_n926));
  NAND2_X1  g501(.A1(new_n926), .A2(new_n606), .ZN(new_n927));
  NOR2_X1   g502(.A1(new_n617), .A2(new_n925), .ZN(new_n928));
  NOR2_X1   g503(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  NOR3_X1   g504(.A1(new_n606), .A2(new_n617), .A3(new_n925), .ZN(new_n930));
  OAI21_X1  g505(.A(new_n924), .B1(new_n929), .B2(new_n930), .ZN(new_n931));
  NAND2_X1  g506(.A1(new_n927), .A2(new_n928), .ZN(new_n932));
  NAND2_X1  g507(.A1(G299), .A2(KEYINPUT104), .ZN(new_n933));
  NAND3_X1  g508(.A1(new_n933), .A2(new_n606), .A3(new_n926), .ZN(new_n934));
  NAND3_X1  g509(.A1(new_n932), .A2(new_n934), .A3(KEYINPUT41), .ZN(new_n935));
  NAND2_X1  g510(.A1(new_n931), .A2(new_n935), .ZN(new_n936));
  AND2_X1   g511(.A1(new_n923), .A2(new_n936), .ZN(new_n937));
  NOR2_X1   g512(.A1(new_n929), .A2(new_n930), .ZN(new_n938));
  NOR2_X1   g513(.A1(new_n923), .A2(new_n938), .ZN(new_n939));
  OAI21_X1  g514(.A(KEYINPUT106), .B1(new_n937), .B2(new_n939), .ZN(new_n940));
  NAND2_X1  g515(.A1(new_n922), .A2(new_n940), .ZN(new_n941));
  NOR3_X1   g516(.A1(new_n937), .A2(new_n939), .A3(KEYINPUT106), .ZN(new_n942));
  XNOR2_X1  g517(.A(new_n941), .B(new_n942), .ZN(new_n943));
  AOI21_X1  g518(.A(new_n911), .B1(new_n943), .B2(G868), .ZN(G295));
  AOI21_X1  g519(.A(new_n911), .B1(new_n943), .B2(G868), .ZN(G331));
  INV_X1    g520(.A(KEYINPUT44), .ZN(new_n946));
  AND3_X1   g521(.A1(new_n861), .A2(G171), .A3(new_n863), .ZN(new_n947));
  AOI21_X1  g522(.A(G171), .B1(new_n861), .B2(new_n863), .ZN(new_n948));
  OAI21_X1  g523(.A(G286), .B1(new_n947), .B2(new_n948), .ZN(new_n949));
  NAND2_X1  g524(.A1(new_n864), .A2(G301), .ZN(new_n950));
  NAND3_X1  g525(.A1(new_n861), .A2(G171), .A3(new_n863), .ZN(new_n951));
  NAND3_X1  g526(.A1(new_n950), .A2(G168), .A3(new_n951), .ZN(new_n952));
  NAND2_X1  g527(.A1(new_n949), .A2(new_n952), .ZN(new_n953));
  NOR3_X1   g528(.A1(new_n929), .A2(new_n924), .A3(new_n930), .ZN(new_n954));
  AOI21_X1  g529(.A(KEYINPUT41), .B1(new_n932), .B2(new_n934), .ZN(new_n955));
  NOR2_X1   g530(.A1(new_n954), .A2(new_n955), .ZN(new_n956));
  INV_X1    g531(.A(KEYINPUT108), .ZN(new_n957));
  NAND3_X1  g532(.A1(new_n953), .A2(new_n956), .A3(new_n957), .ZN(new_n958));
  NAND3_X1  g533(.A1(new_n949), .A2(new_n952), .A3(new_n938), .ZN(new_n959));
  NAND2_X1  g534(.A1(new_n958), .A2(new_n959), .ZN(new_n960));
  AOI21_X1  g535(.A(new_n957), .B1(new_n953), .B2(new_n956), .ZN(new_n961));
  NOR3_X1   g536(.A1(new_n960), .A2(new_n921), .A3(new_n961), .ZN(new_n962));
  AOI21_X1  g537(.A(new_n936), .B1(new_n952), .B2(new_n949), .ZN(new_n963));
  INV_X1    g538(.A(new_n959), .ZN(new_n964));
  OAI21_X1  g539(.A(new_n921), .B1(new_n963), .B2(new_n964), .ZN(new_n965));
  NAND2_X1  g540(.A1(new_n965), .A2(new_n902), .ZN(new_n966));
  OAI21_X1  g541(.A(KEYINPUT43), .B1(new_n962), .B2(new_n966), .ZN(new_n967));
  OAI21_X1  g542(.A(new_n921), .B1(new_n960), .B2(new_n961), .ZN(new_n968));
  NAND2_X1  g543(.A1(new_n953), .A2(new_n956), .ZN(new_n969));
  NAND2_X1  g544(.A1(new_n969), .A2(KEYINPUT108), .ZN(new_n970));
  INV_X1    g545(.A(new_n921), .ZN(new_n971));
  NAND4_X1  g546(.A1(new_n970), .A2(new_n971), .A3(new_n959), .A4(new_n958), .ZN(new_n972));
  XNOR2_X1  g547(.A(KEYINPUT107), .B(KEYINPUT43), .ZN(new_n973));
  NAND4_X1  g548(.A1(new_n968), .A2(new_n972), .A3(new_n902), .A4(new_n973), .ZN(new_n974));
  AOI21_X1  g549(.A(new_n946), .B1(new_n967), .B2(new_n974), .ZN(new_n975));
  INV_X1    g550(.A(new_n966), .ZN(new_n976));
  INV_X1    g551(.A(new_n973), .ZN(new_n977));
  NOR2_X1   g552(.A1(new_n962), .A2(new_n977), .ZN(new_n978));
  NAND3_X1  g553(.A1(new_n968), .A2(new_n902), .A3(new_n972), .ZN(new_n979));
  AOI22_X1  g554(.A1(new_n976), .A2(new_n978), .B1(new_n979), .B2(new_n977), .ZN(new_n980));
  AOI21_X1  g555(.A(new_n975), .B1(new_n980), .B2(new_n946), .ZN(G397));
  OR2_X1    g556(.A1(G290), .A2(G1986), .ZN(new_n982));
  NAND2_X1  g557(.A1(G290), .A2(G1986), .ZN(new_n983));
  NAND3_X1  g558(.A1(new_n982), .A2(KEYINPUT109), .A3(new_n983), .ZN(new_n984));
  INV_X1    g559(.A(KEYINPUT45), .ZN(new_n985));
  OAI21_X1  g560(.A(new_n985), .B1(G164), .B2(G1384), .ZN(new_n986));
  NAND2_X1  g561(.A1(G160), .A2(G40), .ZN(new_n987));
  NOR2_X1   g562(.A1(new_n986), .A2(new_n987), .ZN(new_n988));
  OAI211_X1 g563(.A(new_n984), .B(new_n988), .C1(KEYINPUT109), .C2(new_n983), .ZN(new_n989));
  OR2_X1    g564(.A1(new_n989), .A2(KEYINPUT110), .ZN(new_n990));
  INV_X1    g565(.A(G1996), .ZN(new_n991));
  NAND2_X1  g566(.A1(new_n730), .A2(new_n991), .ZN(new_n992));
  XNOR2_X1  g567(.A(new_n772), .B(new_n774), .ZN(new_n993));
  OAI211_X1 g568(.A(new_n992), .B(new_n993), .C1(new_n991), .C2(new_n889), .ZN(new_n994));
  XNOR2_X1  g569(.A(new_n837), .B(new_n841), .ZN(new_n995));
  XNOR2_X1  g570(.A(new_n995), .B(KEYINPUT111), .ZN(new_n996));
  OAI21_X1  g571(.A(new_n988), .B1(new_n994), .B2(new_n996), .ZN(new_n997));
  NAND2_X1  g572(.A1(new_n989), .A2(KEYINPUT110), .ZN(new_n998));
  NAND3_X1  g573(.A1(new_n990), .A2(new_n997), .A3(new_n998), .ZN(new_n999));
  XNOR2_X1  g574(.A(new_n999), .B(KEYINPUT112), .ZN(new_n1000));
  INV_X1    g575(.A(KEYINPUT61), .ZN(new_n1001));
  OAI21_X1  g576(.A(KEYINPUT50), .B1(G164), .B2(G1384), .ZN(new_n1002));
  INV_X1    g577(.A(KEYINPUT50), .ZN(new_n1003));
  INV_X1    g578(.A(G1384), .ZN(new_n1004));
  NAND3_X1  g579(.A1(new_n750), .A2(new_n1003), .A3(new_n1004), .ZN(new_n1005));
  INV_X1    g580(.A(G40), .ZN(new_n1006));
  NOR3_X1   g581(.A1(new_n466), .A2(new_n471), .A3(new_n1006), .ZN(new_n1007));
  NAND3_X1  g582(.A1(new_n1002), .A2(new_n1005), .A3(new_n1007), .ZN(new_n1008));
  INV_X1    g583(.A(KEYINPUT120), .ZN(new_n1009));
  INV_X1    g584(.A(G1956), .ZN(new_n1010));
  AND3_X1   g585(.A1(new_n1008), .A2(new_n1009), .A3(new_n1010), .ZN(new_n1011));
  AOI21_X1  g586(.A(new_n1009), .B1(new_n1008), .B2(new_n1010), .ZN(new_n1012));
  NOR2_X1   g587(.A1(new_n1011), .A2(new_n1012), .ZN(new_n1013));
  INV_X1    g588(.A(KEYINPUT57), .ZN(new_n1014));
  OAI21_X1  g589(.A(new_n1014), .B1(new_n614), .B2(KEYINPUT121), .ZN(new_n1015));
  XNOR2_X1  g590(.A(G299), .B(new_n1015), .ZN(new_n1016));
  XNOR2_X1  g591(.A(KEYINPUT122), .B(KEYINPUT56), .ZN(new_n1017));
  XNOR2_X1  g592(.A(new_n1017), .B(G2072), .ZN(new_n1018));
  INV_X1    g593(.A(new_n1018), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n491), .A2(new_n493), .ZN(new_n1020));
  AOI21_X1  g595(.A(G1384), .B1(new_n1020), .B2(new_n747), .ZN(new_n1021));
  NAND2_X1  g596(.A1(new_n1021), .A2(KEYINPUT45), .ZN(new_n1022));
  INV_X1    g597(.A(KEYINPUT113), .ZN(new_n1023));
  NAND3_X1  g598(.A1(new_n1022), .A2(new_n986), .A3(new_n1023), .ZN(new_n1024));
  OAI211_X1 g599(.A(KEYINPUT113), .B(new_n985), .C1(G164), .C2(G1384), .ZN(new_n1025));
  AOI211_X1 g600(.A(new_n987), .B(new_n1019), .C1(new_n1024), .C2(new_n1025), .ZN(new_n1026));
  NOR3_X1   g601(.A1(new_n1013), .A2(new_n1016), .A3(new_n1026), .ZN(new_n1027));
  INV_X1    g602(.A(new_n1016), .ZN(new_n1028));
  NAND2_X1  g603(.A1(new_n1008), .A2(new_n1010), .ZN(new_n1029));
  NAND2_X1  g604(.A1(new_n1029), .A2(KEYINPUT120), .ZN(new_n1030));
  NAND3_X1  g605(.A1(new_n1008), .A2(new_n1009), .A3(new_n1010), .ZN(new_n1031));
  NAND2_X1  g606(.A1(new_n1030), .A2(new_n1031), .ZN(new_n1032));
  AOI21_X1  g607(.A(new_n987), .B1(new_n1024), .B2(new_n1025), .ZN(new_n1033));
  NAND2_X1  g608(.A1(new_n1033), .A2(new_n1018), .ZN(new_n1034));
  AOI21_X1  g609(.A(new_n1028), .B1(new_n1032), .B2(new_n1034), .ZN(new_n1035));
  OAI21_X1  g610(.A(new_n1001), .B1(new_n1027), .B2(new_n1035), .ZN(new_n1036));
  OAI21_X1  g611(.A(new_n1007), .B1(new_n1021), .B2(new_n1003), .ZN(new_n1037));
  INV_X1    g612(.A(new_n1037), .ZN(new_n1038));
  NAND4_X1  g613(.A1(new_n750), .A2(KEYINPUT114), .A3(new_n1003), .A4(new_n1004), .ZN(new_n1039));
  INV_X1    g614(.A(KEYINPUT114), .ZN(new_n1040));
  NAND2_X1  g615(.A1(new_n1003), .A2(new_n1004), .ZN(new_n1041));
  OAI21_X1  g616(.A(new_n1040), .B1(G164), .B2(new_n1041), .ZN(new_n1042));
  NAND2_X1  g617(.A1(new_n1039), .A2(new_n1042), .ZN(new_n1043));
  AOI21_X1  g618(.A(G1348), .B1(new_n1038), .B2(new_n1043), .ZN(new_n1044));
  NOR4_X1   g619(.A1(new_n987), .A2(G1384), .A3(G2067), .A4(G164), .ZN(new_n1045));
  NOR2_X1   g620(.A1(new_n1044), .A2(new_n1045), .ZN(new_n1046));
  AOI21_X1  g621(.A(new_n607), .B1(new_n1046), .B2(KEYINPUT60), .ZN(new_n1047));
  INV_X1    g622(.A(KEYINPUT60), .ZN(new_n1048));
  NOR4_X1   g623(.A1(new_n1044), .A2(new_n1048), .A3(new_n606), .A4(new_n1045), .ZN(new_n1049));
  OAI22_X1  g624(.A1(new_n1047), .A2(new_n1049), .B1(KEYINPUT60), .B2(new_n1046), .ZN(new_n1050));
  AND2_X1   g625(.A1(new_n555), .A2(KEYINPUT123), .ZN(new_n1051));
  AOI211_X1 g626(.A(G1996), .B(new_n987), .C1(new_n1024), .C2(new_n1025), .ZN(new_n1052));
  XNOR2_X1  g627(.A(KEYINPUT58), .B(G1341), .ZN(new_n1053));
  AOI21_X1  g628(.A(new_n1053), .B1(new_n1007), .B2(new_n1021), .ZN(new_n1054));
  OAI21_X1  g629(.A(new_n1051), .B1(new_n1052), .B2(new_n1054), .ZN(new_n1055));
  NAND2_X1  g630(.A1(new_n1055), .A2(KEYINPUT59), .ZN(new_n1056));
  INV_X1    g631(.A(KEYINPUT59), .ZN(new_n1057));
  OAI211_X1 g632(.A(new_n1057), .B(new_n1051), .C1(new_n1052), .C2(new_n1054), .ZN(new_n1058));
  NAND2_X1  g633(.A1(new_n1056), .A2(new_n1058), .ZN(new_n1059));
  OAI21_X1  g634(.A(new_n1016), .B1(new_n1013), .B2(new_n1026), .ZN(new_n1060));
  NAND3_X1  g635(.A1(new_n1032), .A2(new_n1028), .A3(new_n1034), .ZN(new_n1061));
  NAND3_X1  g636(.A1(new_n1060), .A2(KEYINPUT61), .A3(new_n1061), .ZN(new_n1062));
  NAND4_X1  g637(.A1(new_n1036), .A2(new_n1050), .A3(new_n1059), .A4(new_n1062), .ZN(new_n1063));
  NOR2_X1   g638(.A1(new_n1046), .A2(new_n607), .ZN(new_n1064));
  OAI21_X1  g639(.A(new_n1061), .B1(new_n1035), .B2(new_n1064), .ZN(new_n1065));
  NAND2_X1  g640(.A1(new_n1063), .A2(new_n1065), .ZN(new_n1066));
  AOI21_X1  g641(.A(KEYINPUT45), .B1(new_n750), .B2(new_n1004), .ZN(new_n1067));
  OAI21_X1  g642(.A(KEYINPUT118), .B1(new_n1067), .B2(new_n987), .ZN(new_n1068));
  INV_X1    g643(.A(KEYINPUT118), .ZN(new_n1069));
  NAND3_X1  g644(.A1(new_n986), .A2(new_n1069), .A3(new_n1007), .ZN(new_n1070));
  NAND3_X1  g645(.A1(new_n1068), .A2(new_n1070), .A3(new_n1022), .ZN(new_n1071));
  INV_X1    g646(.A(G1966), .ZN(new_n1072));
  NAND2_X1  g647(.A1(new_n1071), .A2(new_n1072), .ZN(new_n1073));
  AOI21_X1  g648(.A(new_n1037), .B1(new_n1042), .B2(new_n1039), .ZN(new_n1074));
  INV_X1    g649(.A(G2084), .ZN(new_n1075));
  NAND2_X1  g650(.A1(new_n1074), .A2(new_n1075), .ZN(new_n1076));
  NAND2_X1  g651(.A1(new_n1073), .A2(new_n1076), .ZN(new_n1077));
  OAI211_X1 g652(.A(KEYINPUT51), .B(G8), .C1(new_n1077), .C2(G286), .ZN(new_n1078));
  INV_X1    g653(.A(KEYINPUT124), .ZN(new_n1079));
  NAND2_X1  g654(.A1(new_n1078), .A2(new_n1079), .ZN(new_n1080));
  INV_X1    g655(.A(G8), .ZN(new_n1081));
  AOI21_X1  g656(.A(new_n1081), .B1(new_n1073), .B2(new_n1076), .ZN(new_n1082));
  NOR2_X1   g657(.A1(G168), .A2(new_n1081), .ZN(new_n1083));
  OAI211_X1 g658(.A(KEYINPUT124), .B(KEYINPUT51), .C1(new_n1082), .C2(new_n1083), .ZN(new_n1084));
  AOI22_X1  g659(.A1(new_n1071), .A2(new_n1072), .B1(new_n1074), .B2(new_n1075), .ZN(new_n1085));
  OAI21_X1  g660(.A(KEYINPUT125), .B1(new_n1085), .B2(new_n1081), .ZN(new_n1086));
  INV_X1    g661(.A(KEYINPUT125), .ZN(new_n1087));
  NAND2_X1  g662(.A1(new_n986), .A2(new_n1007), .ZN(new_n1088));
  AOI22_X1  g663(.A1(new_n1088), .A2(KEYINPUT118), .B1(KEYINPUT45), .B2(new_n1021), .ZN(new_n1089));
  AOI21_X1  g664(.A(G1966), .B1(new_n1089), .B2(new_n1070), .ZN(new_n1090));
  NAND2_X1  g665(.A1(new_n1038), .A2(new_n1043), .ZN(new_n1091));
  NOR2_X1   g666(.A1(new_n1091), .A2(G2084), .ZN(new_n1092));
  OAI211_X1 g667(.A(new_n1087), .B(G8), .C1(new_n1090), .C2(new_n1092), .ZN(new_n1093));
  NOR2_X1   g668(.A1(new_n1083), .A2(KEYINPUT51), .ZN(new_n1094));
  NAND3_X1  g669(.A1(new_n1086), .A2(new_n1093), .A3(new_n1094), .ZN(new_n1095));
  NAND3_X1  g670(.A1(new_n1080), .A2(new_n1084), .A3(new_n1095), .ZN(new_n1096));
  NAND2_X1  g671(.A1(new_n1077), .A2(new_n1083), .ZN(new_n1097));
  NAND2_X1  g672(.A1(new_n1096), .A2(new_n1097), .ZN(new_n1098));
  INV_X1    g673(.A(G1961), .ZN(new_n1099));
  NAND2_X1  g674(.A1(new_n1091), .A2(new_n1099), .ZN(new_n1100));
  NAND4_X1  g675(.A1(new_n1068), .A2(new_n752), .A3(new_n1070), .A4(new_n1022), .ZN(new_n1101));
  INV_X1    g676(.A(KEYINPUT126), .ZN(new_n1102));
  NAND2_X1  g677(.A1(new_n1101), .A2(new_n1102), .ZN(new_n1103));
  INV_X1    g678(.A(new_n1103), .ZN(new_n1104));
  OAI21_X1  g679(.A(KEYINPUT53), .B1(new_n1101), .B2(new_n1102), .ZN(new_n1105));
  OAI21_X1  g680(.A(new_n1100), .B1(new_n1104), .B2(new_n1105), .ZN(new_n1106));
  AOI211_X1 g681(.A(G2078), .B(new_n987), .C1(new_n1024), .C2(new_n1025), .ZN(new_n1107));
  NOR2_X1   g682(.A1(new_n1107), .A2(KEYINPUT53), .ZN(new_n1108));
  OAI21_X1  g683(.A(G171), .B1(new_n1106), .B2(new_n1108), .ZN(new_n1109));
  NAND2_X1  g684(.A1(new_n1033), .A2(new_n752), .ZN(new_n1110));
  INV_X1    g685(.A(KEYINPUT53), .ZN(new_n1111));
  AOI21_X1  g686(.A(G171), .B1(new_n1110), .B2(new_n1111), .ZN(new_n1112));
  INV_X1    g687(.A(new_n1088), .ZN(new_n1113));
  AOI211_X1 g688(.A(new_n1111), .B(G2078), .C1(new_n1021), .C2(KEYINPUT45), .ZN(new_n1114));
  AOI22_X1  g689(.A1(new_n1091), .A2(new_n1099), .B1(new_n1113), .B2(new_n1114), .ZN(new_n1115));
  NAND2_X1  g690(.A1(new_n1112), .A2(new_n1115), .ZN(new_n1116));
  NAND2_X1  g691(.A1(new_n1109), .A2(new_n1116), .ZN(new_n1117));
  INV_X1    g692(.A(KEYINPUT54), .ZN(new_n1118));
  NAND2_X1  g693(.A1(new_n1117), .A2(new_n1118), .ZN(new_n1119));
  OAI21_X1  g694(.A(new_n1115), .B1(new_n1107), .B2(KEYINPUT53), .ZN(new_n1120));
  AOI21_X1  g695(.A(new_n1118), .B1(new_n1120), .B2(G171), .ZN(new_n1121));
  NAND4_X1  g696(.A1(new_n1089), .A2(KEYINPUT126), .A3(new_n752), .A4(new_n1070), .ZN(new_n1122));
  NAND3_X1  g697(.A1(new_n1122), .A2(new_n1103), .A3(KEYINPUT53), .ZN(new_n1123));
  NAND3_X1  g698(.A1(new_n1123), .A2(new_n1112), .A3(new_n1100), .ZN(new_n1124));
  AND2_X1   g699(.A1(new_n1121), .A2(new_n1124), .ZN(new_n1125));
  INV_X1    g700(.A(G1981), .ZN(new_n1126));
  INV_X1    g701(.A(KEYINPUT116), .ZN(new_n1127));
  AOI21_X1  g702(.A(new_n1126), .B1(new_n584), .B2(new_n1127), .ZN(new_n1128));
  NAND2_X1  g703(.A1(new_n1128), .A2(G305), .ZN(new_n1129));
  OAI21_X1  g704(.A(G1981), .B1(new_n818), .B2(KEYINPUT116), .ZN(new_n1130));
  NAND2_X1  g705(.A1(new_n1130), .A2(new_n819), .ZN(new_n1131));
  NAND2_X1  g706(.A1(new_n1129), .A2(new_n1131), .ZN(new_n1132));
  INV_X1    g707(.A(KEYINPUT49), .ZN(new_n1133));
  NAND2_X1  g708(.A1(new_n1132), .A2(new_n1133), .ZN(new_n1134));
  NAND3_X1  g709(.A1(new_n1129), .A2(new_n1131), .A3(KEYINPUT49), .ZN(new_n1135));
  AOI21_X1  g710(.A(new_n1081), .B1(new_n1007), .B2(new_n1021), .ZN(new_n1136));
  NAND3_X1  g711(.A1(new_n1134), .A2(new_n1135), .A3(new_n1136), .ZN(new_n1137));
  INV_X1    g712(.A(KEYINPUT117), .ZN(new_n1138));
  NAND2_X1  g713(.A1(new_n1137), .A2(new_n1138), .ZN(new_n1139));
  INV_X1    g714(.A(new_n1136), .ZN(new_n1140));
  AOI21_X1  g715(.A(new_n1140), .B1(new_n1132), .B2(new_n1133), .ZN(new_n1141));
  NAND3_X1  g716(.A1(new_n1141), .A2(KEYINPUT117), .A3(new_n1135), .ZN(new_n1142));
  NAND2_X1  g717(.A1(new_n1139), .A2(new_n1142), .ZN(new_n1143));
  OAI22_X1  g718(.A1(new_n1033), .A2(G1971), .B1(G2090), .B2(new_n1008), .ZN(new_n1144));
  NAND2_X1  g719(.A1(new_n1144), .A2(G8), .ZN(new_n1145));
  NAND2_X1  g720(.A1(G303), .A2(G8), .ZN(new_n1146));
  XNOR2_X1  g721(.A(new_n1146), .B(KEYINPUT55), .ZN(new_n1147));
  NAND2_X1  g722(.A1(new_n1145), .A2(new_n1147), .ZN(new_n1148));
  INV_X1    g723(.A(new_n1147), .ZN(new_n1149));
  OAI22_X1  g724(.A1(new_n1033), .A2(G1971), .B1(new_n1091), .B2(G2090), .ZN(new_n1150));
  NAND3_X1  g725(.A1(new_n1149), .A2(new_n1150), .A3(G8), .ZN(new_n1151));
  INV_X1    g726(.A(KEYINPUT52), .ZN(new_n1152));
  AND2_X1   g727(.A1(new_n574), .A2(new_n576), .ZN(new_n1153));
  NAND4_X1  g728(.A1(new_n1153), .A2(G1976), .A3(new_n571), .A4(new_n572), .ZN(new_n1154));
  AOI21_X1  g729(.A(new_n1152), .B1(new_n1136), .B2(new_n1154), .ZN(new_n1155));
  INV_X1    g730(.A(new_n1155), .ZN(new_n1156));
  INV_X1    g731(.A(G1976), .ZN(new_n1157));
  NAND2_X1  g732(.A1(G288), .A2(new_n1157), .ZN(new_n1158));
  NAND4_X1  g733(.A1(new_n1136), .A2(new_n1152), .A3(new_n1154), .A4(new_n1158), .ZN(new_n1159));
  AOI21_X1  g734(.A(KEYINPUT115), .B1(new_n1156), .B2(new_n1159), .ZN(new_n1160));
  NAND2_X1  g735(.A1(new_n1159), .A2(KEYINPUT115), .ZN(new_n1161));
  INV_X1    g736(.A(new_n1161), .ZN(new_n1162));
  NOR2_X1   g737(.A1(new_n1160), .A2(new_n1162), .ZN(new_n1163));
  NAND4_X1  g738(.A1(new_n1143), .A2(new_n1148), .A3(new_n1151), .A4(new_n1163), .ZN(new_n1164));
  NOR2_X1   g739(.A1(new_n1125), .A2(new_n1164), .ZN(new_n1165));
  NAND4_X1  g740(.A1(new_n1066), .A2(new_n1098), .A3(new_n1119), .A4(new_n1165), .ZN(new_n1166));
  INV_X1    g741(.A(KEYINPUT115), .ZN(new_n1167));
  INV_X1    g742(.A(new_n1159), .ZN(new_n1168));
  OAI21_X1  g743(.A(new_n1167), .B1(new_n1168), .B2(new_n1155), .ZN(new_n1169));
  NAND2_X1  g744(.A1(new_n1169), .A2(new_n1161), .ZN(new_n1170));
  AOI21_X1  g745(.A(new_n1170), .B1(new_n1139), .B2(new_n1142), .ZN(new_n1171));
  INV_X1    g746(.A(new_n1151), .ZN(new_n1172));
  NAND2_X1  g747(.A1(new_n1171), .A2(new_n1172), .ZN(new_n1173));
  NOR2_X1   g748(.A1(G288), .A2(G1976), .ZN(new_n1174));
  AOI22_X1  g749(.A1(new_n1143), .A2(new_n1174), .B1(new_n1126), .B2(new_n819), .ZN(new_n1175));
  OAI21_X1  g750(.A(new_n1173), .B1(new_n1175), .B2(new_n1140), .ZN(new_n1176));
  AND3_X1   g751(.A1(new_n1141), .A2(KEYINPUT117), .A3(new_n1135), .ZN(new_n1177));
  AOI21_X1  g752(.A(KEYINPUT117), .B1(new_n1141), .B2(new_n1135), .ZN(new_n1178));
  OAI21_X1  g753(.A(new_n1163), .B1(new_n1177), .B2(new_n1178), .ZN(new_n1179));
  AOI21_X1  g754(.A(new_n1149), .B1(new_n1150), .B2(G8), .ZN(new_n1180));
  OAI21_X1  g755(.A(KEYINPUT119), .B1(new_n1179), .B2(new_n1180), .ZN(new_n1181));
  INV_X1    g756(.A(new_n1180), .ZN(new_n1182));
  INV_X1    g757(.A(KEYINPUT119), .ZN(new_n1183));
  NAND3_X1  g758(.A1(new_n1171), .A2(new_n1182), .A3(new_n1183), .ZN(new_n1184));
  NAND2_X1  g759(.A1(new_n1082), .A2(G168), .ZN(new_n1185));
  INV_X1    g760(.A(KEYINPUT63), .ZN(new_n1186));
  NOR3_X1   g761(.A1(new_n1172), .A2(new_n1185), .A3(new_n1186), .ZN(new_n1187));
  NAND3_X1  g762(.A1(new_n1181), .A2(new_n1184), .A3(new_n1187), .ZN(new_n1188));
  OAI21_X1  g763(.A(new_n1186), .B1(new_n1164), .B2(new_n1185), .ZN(new_n1189));
  AOI21_X1  g764(.A(new_n1176), .B1(new_n1188), .B2(new_n1189), .ZN(new_n1190));
  NAND2_X1  g765(.A1(new_n1166), .A2(new_n1190), .ZN(new_n1191));
  INV_X1    g766(.A(KEYINPUT62), .ZN(new_n1192));
  AND3_X1   g767(.A1(new_n1096), .A2(new_n1192), .A3(new_n1097), .ZN(new_n1193));
  AOI21_X1  g768(.A(new_n1192), .B1(new_n1096), .B2(new_n1097), .ZN(new_n1194));
  OR2_X1    g769(.A1(new_n1164), .A2(new_n1109), .ZN(new_n1195));
  NOR3_X1   g770(.A1(new_n1193), .A2(new_n1194), .A3(new_n1195), .ZN(new_n1196));
  OAI21_X1  g771(.A(new_n1000), .B1(new_n1191), .B2(new_n1196), .ZN(new_n1197));
  INV_X1    g772(.A(new_n988), .ZN(new_n1198));
  NOR2_X1   g773(.A1(new_n1198), .A2(new_n982), .ZN(new_n1199));
  XOR2_X1   g774(.A(new_n1199), .B(KEYINPUT48), .Z(new_n1200));
  AND2_X1   g775(.A1(new_n1200), .A2(new_n997), .ZN(new_n1201));
  AOI21_X1  g776(.A(new_n1198), .B1(new_n993), .B2(new_n889), .ZN(new_n1202));
  OR3_X1    g777(.A1(new_n1198), .A2(KEYINPUT46), .A3(G1996), .ZN(new_n1203));
  OAI21_X1  g778(.A(KEYINPUT46), .B1(new_n1198), .B2(G1996), .ZN(new_n1204));
  AOI21_X1  g779(.A(new_n1202), .B1(new_n1203), .B2(new_n1204), .ZN(new_n1205));
  XNOR2_X1  g780(.A(new_n1205), .B(KEYINPUT47), .ZN(new_n1206));
  NAND2_X1  g781(.A1(new_n838), .A2(new_n841), .ZN(new_n1207));
  OAI22_X1  g782(.A1(new_n994), .A2(new_n1207), .B1(G2067), .B2(new_n772), .ZN(new_n1208));
  AOI211_X1 g783(.A(new_n1201), .B(new_n1206), .C1(new_n988), .C2(new_n1208), .ZN(new_n1209));
  XNOR2_X1  g784(.A(new_n1209), .B(KEYINPUT127), .ZN(new_n1210));
  NAND2_X1  g785(.A1(new_n1197), .A2(new_n1210), .ZN(G329));
  assign    G231 = 1'b0;
  OR2_X1    g786(.A1(G227), .A2(new_n460), .ZN(new_n1213));
  NOR3_X1   g787(.A1(G401), .A2(G229), .A3(new_n1213), .ZN(new_n1214));
  NAND2_X1  g788(.A1(new_n1214), .A2(new_n908), .ZN(new_n1215));
  NOR2_X1   g789(.A1(new_n1215), .A2(new_n980), .ZN(G308));
  AND2_X1   g790(.A1(new_n979), .A2(new_n977), .ZN(new_n1217));
  NOR3_X1   g791(.A1(new_n962), .A2(new_n966), .A3(new_n977), .ZN(new_n1218));
  OAI211_X1 g792(.A(new_n908), .B(new_n1214), .C1(new_n1217), .C2(new_n1218), .ZN(G225));
endmodule


