//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 1 0 0 1 0 1 0 0 0 1 1 0 0 0 1 1 1 0 1 0 0 0 0 1 0 0 0 0 1 1 0 1 0 1 0 0 1 1 1 0 1 0 1 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 1 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:20:22 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n674, new_n675, new_n676, new_n677, new_n678, new_n680,
    new_n681, new_n682, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n703,
    new_n704, new_n705, new_n706, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n716, new_n717, new_n718, new_n719,
    new_n721, new_n722, new_n723, new_n724, new_n726, new_n727, new_n728,
    new_n729, new_n730, new_n731, new_n732, new_n733, new_n734, new_n735,
    new_n737, new_n738, new_n739, new_n741, new_n742, new_n744, new_n745,
    new_n746, new_n747, new_n748, new_n749, new_n750, new_n751, new_n752,
    new_n753, new_n754, new_n755, new_n756, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n772, new_n773, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n837, new_n838, new_n839, new_n841, new_n842,
    new_n844, new_n845, new_n846, new_n847, new_n848, new_n849, new_n850,
    new_n851, new_n852, new_n853, new_n854, new_n855, new_n856, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n923,
    new_n924, new_n925, new_n927, new_n928, new_n929, new_n930, new_n931,
    new_n932, new_n933, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n944, new_n945, new_n946, new_n948,
    new_n949, new_n950, new_n951, new_n952, new_n953, new_n954, new_n955,
    new_n956, new_n957, new_n958, new_n959, new_n960, new_n962, new_n963,
    new_n964, new_n966, new_n967, new_n968, new_n969, new_n970, new_n971,
    new_n972, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n982, new_n983, new_n984, new_n985, new_n987, new_n988,
    new_n989;
  INV_X1    g000(.A(KEYINPUT66), .ZN(new_n202));
  INV_X1    g001(.A(KEYINPUT27), .ZN(new_n203));
  NAND2_X1  g002(.A1(new_n203), .A2(G183gat), .ZN(new_n204));
  INV_X1    g003(.A(G183gat), .ZN(new_n205));
  NAND2_X1  g004(.A1(new_n205), .A2(KEYINPUT27), .ZN(new_n206));
  AOI21_X1  g005(.A(new_n202), .B1(new_n204), .B2(new_n206), .ZN(new_n207));
  OAI21_X1  g006(.A(new_n202), .B1(new_n205), .B2(KEYINPUT27), .ZN(new_n208));
  INV_X1    g007(.A(G190gat), .ZN(new_n209));
  NAND2_X1  g008(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  OAI21_X1  g009(.A(KEYINPUT67), .B1(new_n207), .B2(new_n210), .ZN(new_n211));
  AOI21_X1  g010(.A(G190gat), .B1(new_n204), .B2(new_n202), .ZN(new_n212));
  INV_X1    g011(.A(KEYINPUT67), .ZN(new_n213));
  XNOR2_X1  g012(.A(KEYINPUT27), .B(G183gat), .ZN(new_n214));
  OAI211_X1 g013(.A(new_n212), .B(new_n213), .C1(new_n202), .C2(new_n214), .ZN(new_n215));
  INV_X1    g014(.A(KEYINPUT28), .ZN(new_n216));
  NAND3_X1  g015(.A1(new_n211), .A2(new_n215), .A3(new_n216), .ZN(new_n217));
  NAND3_X1  g016(.A1(new_n214), .A2(KEYINPUT28), .A3(new_n209), .ZN(new_n218));
  NAND2_X1  g017(.A1(new_n217), .A2(new_n218), .ZN(new_n219));
  INV_X1    g018(.A(KEYINPUT69), .ZN(new_n220));
  NAND2_X1  g019(.A1(G183gat), .A2(G190gat), .ZN(new_n221));
  OAI21_X1  g020(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n222));
  NAND2_X1  g021(.A1(G169gat), .A2(G176gat), .ZN(new_n223));
  NAND3_X1  g022(.A1(new_n222), .A2(KEYINPUT68), .A3(new_n223), .ZN(new_n224));
  NOR2_X1   g023(.A1(G169gat), .A2(G176gat), .ZN(new_n225));
  INV_X1    g024(.A(new_n225), .ZN(new_n226));
  OAI21_X1  g025(.A(new_n224), .B1(KEYINPUT26), .B2(new_n226), .ZN(new_n227));
  AOI21_X1  g026(.A(KEYINPUT68), .B1(new_n222), .B2(new_n223), .ZN(new_n228));
  OAI211_X1 g027(.A(new_n220), .B(new_n221), .C1(new_n227), .C2(new_n228), .ZN(new_n229));
  OAI21_X1  g028(.A(new_n221), .B1(new_n227), .B2(new_n228), .ZN(new_n230));
  NAND2_X1  g029(.A1(new_n230), .A2(KEYINPUT69), .ZN(new_n231));
  NAND3_X1  g030(.A1(new_n219), .A2(new_n229), .A3(new_n231), .ZN(new_n232));
  XOR2_X1   g031(.A(new_n223), .B(KEYINPUT65), .Z(new_n233));
  OR2_X1    g032(.A1(new_n225), .A2(KEYINPUT23), .ZN(new_n234));
  NAND3_X1  g033(.A1(new_n233), .A2(KEYINPUT25), .A3(new_n234), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n205), .A2(new_n209), .ZN(new_n236));
  NAND3_X1  g035(.A1(new_n236), .A2(KEYINPUT24), .A3(new_n221), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n225), .A2(KEYINPUT23), .ZN(new_n238));
  OAI211_X1 g037(.A(new_n237), .B(new_n238), .C1(KEYINPUT24), .C2(new_n221), .ZN(new_n239));
  OR2_X1    g038(.A1(new_n235), .A2(new_n239), .ZN(new_n240));
  INV_X1    g039(.A(KEYINPUT25), .ZN(new_n241));
  NAND2_X1  g040(.A1(new_n234), .A2(new_n223), .ZN(new_n242));
  OAI21_X1  g041(.A(new_n241), .B1(new_n239), .B2(new_n242), .ZN(new_n243));
  NAND2_X1  g042(.A1(new_n240), .A2(new_n243), .ZN(new_n244));
  NAND2_X1  g043(.A1(new_n232), .A2(new_n244), .ZN(new_n245));
  INV_X1    g044(.A(G113gat), .ZN(new_n246));
  INV_X1    g045(.A(G120gat), .ZN(new_n247));
  AOI21_X1  g046(.A(KEYINPUT1), .B1(new_n246), .B2(new_n247), .ZN(new_n248));
  NAND2_X1  g047(.A1(G113gat), .A2(G120gat), .ZN(new_n249));
  AND2_X1   g048(.A1(new_n248), .A2(new_n249), .ZN(new_n250));
  XNOR2_X1  g049(.A(G127gat), .B(G134gat), .ZN(new_n251));
  INV_X1    g050(.A(KEYINPUT70), .ZN(new_n252));
  NAND2_X1  g051(.A1(new_n251), .A2(new_n252), .ZN(new_n253));
  INV_X1    g052(.A(G127gat), .ZN(new_n254));
  NOR2_X1   g053(.A1(new_n254), .A2(G134gat), .ZN(new_n255));
  INV_X1    g054(.A(G134gat), .ZN(new_n256));
  NOR2_X1   g055(.A1(new_n256), .A2(G127gat), .ZN(new_n257));
  OAI21_X1  g056(.A(KEYINPUT70), .B1(new_n255), .B2(new_n257), .ZN(new_n258));
  NAND3_X1  g057(.A1(new_n250), .A2(new_n253), .A3(new_n258), .ZN(new_n259));
  NAND2_X1  g058(.A1(new_n248), .A2(new_n249), .ZN(new_n260));
  NAND3_X1  g059(.A1(new_n260), .A2(new_n252), .A3(new_n251), .ZN(new_n261));
  NAND2_X1  g060(.A1(new_n259), .A2(new_n261), .ZN(new_n262));
  INV_X1    g061(.A(KEYINPUT71), .ZN(new_n263));
  NAND2_X1  g062(.A1(new_n262), .A2(new_n263), .ZN(new_n264));
  NAND3_X1  g063(.A1(new_n259), .A2(KEYINPUT71), .A3(new_n261), .ZN(new_n265));
  NAND2_X1  g064(.A1(new_n264), .A2(new_n265), .ZN(new_n266));
  NAND2_X1  g065(.A1(new_n245), .A2(new_n266), .ZN(new_n267));
  AND2_X1   g066(.A1(new_n264), .A2(new_n265), .ZN(new_n268));
  NAND3_X1  g067(.A1(new_n268), .A2(new_n232), .A3(new_n244), .ZN(new_n269));
  NAND2_X1  g068(.A1(new_n267), .A2(new_n269), .ZN(new_n270));
  NAND2_X1  g069(.A1(G227gat), .A2(G233gat), .ZN(new_n271));
  XNOR2_X1  g070(.A(new_n271), .B(KEYINPUT64), .ZN(new_n272));
  OAI21_X1  g071(.A(KEYINPUT34), .B1(new_n270), .B2(new_n272), .ZN(new_n273));
  INV_X1    g072(.A(KEYINPUT34), .ZN(new_n274));
  INV_X1    g073(.A(new_n272), .ZN(new_n275));
  NAND4_X1  g074(.A1(new_n267), .A2(new_n274), .A3(new_n275), .A4(new_n269), .ZN(new_n276));
  NAND2_X1  g075(.A1(new_n273), .A2(new_n276), .ZN(new_n277));
  XNOR2_X1  g076(.A(G15gat), .B(G43gat), .ZN(new_n278));
  XNOR2_X1  g077(.A(new_n278), .B(KEYINPUT72), .ZN(new_n279));
  INV_X1    g078(.A(G71gat), .ZN(new_n280));
  XNOR2_X1  g079(.A(new_n279), .B(new_n280), .ZN(new_n281));
  INV_X1    g080(.A(G99gat), .ZN(new_n282));
  XNOR2_X1  g081(.A(new_n281), .B(new_n282), .ZN(new_n283));
  AOI21_X1  g082(.A(new_n275), .B1(new_n267), .B2(new_n269), .ZN(new_n284));
  OAI21_X1  g083(.A(new_n283), .B1(new_n284), .B2(KEYINPUT33), .ZN(new_n285));
  INV_X1    g084(.A(KEYINPUT32), .ZN(new_n286));
  NOR2_X1   g085(.A1(new_n284), .A2(new_n286), .ZN(new_n287));
  NOR2_X1   g086(.A1(new_n285), .A2(new_n287), .ZN(new_n288));
  AOI221_X4 g087(.A(new_n286), .B1(KEYINPUT33), .B2(new_n283), .C1(new_n270), .C2(new_n272), .ZN(new_n289));
  OAI21_X1  g088(.A(new_n277), .B1(new_n288), .B2(new_n289), .ZN(new_n290));
  INV_X1    g089(.A(new_n269), .ZN(new_n291));
  AOI21_X1  g090(.A(new_n268), .B1(new_n244), .B2(new_n232), .ZN(new_n292));
  OAI21_X1  g091(.A(new_n272), .B1(new_n291), .B2(new_n292), .ZN(new_n293));
  NAND2_X1  g092(.A1(new_n293), .A2(KEYINPUT32), .ZN(new_n294));
  INV_X1    g093(.A(KEYINPUT33), .ZN(new_n295));
  NAND2_X1  g094(.A1(new_n293), .A2(new_n295), .ZN(new_n296));
  NAND3_X1  g095(.A1(new_n294), .A2(new_n296), .A3(new_n283), .ZN(new_n297));
  AND2_X1   g096(.A1(new_n273), .A2(new_n276), .ZN(new_n298));
  INV_X1    g097(.A(new_n283), .ZN(new_n299));
  OAI211_X1 g098(.A(new_n293), .B(KEYINPUT32), .C1(new_n295), .C2(new_n299), .ZN(new_n300));
  NAND3_X1  g099(.A1(new_n297), .A2(new_n298), .A3(new_n300), .ZN(new_n301));
  NAND2_X1  g100(.A1(new_n290), .A2(new_n301), .ZN(new_n302));
  INV_X1    g101(.A(new_n302), .ZN(new_n303));
  INV_X1    g102(.A(KEYINPUT36), .ZN(new_n304));
  NAND2_X1  g103(.A1(new_n303), .A2(new_n304), .ZN(new_n305));
  INV_X1    g104(.A(KEYINPUT73), .ZN(new_n306));
  AOI211_X1 g105(.A(new_n306), .B(new_n277), .C1(new_n297), .C2(new_n300), .ZN(new_n307));
  NAND2_X1  g106(.A1(new_n297), .A2(new_n300), .ZN(new_n308));
  NAND2_X1  g107(.A1(new_n308), .A2(KEYINPUT73), .ZN(new_n309));
  AOI21_X1  g108(.A(new_n307), .B1(new_n302), .B2(new_n309), .ZN(new_n310));
  OAI21_X1  g109(.A(new_n305), .B1(new_n310), .B2(new_n304), .ZN(new_n311));
  INV_X1    g110(.A(KEYINPUT3), .ZN(new_n312));
  INV_X1    g111(.A(G141gat), .ZN(new_n313));
  NAND2_X1  g112(.A1(new_n313), .A2(G148gat), .ZN(new_n314));
  INV_X1    g113(.A(G148gat), .ZN(new_n315));
  NAND2_X1  g114(.A1(new_n315), .A2(G141gat), .ZN(new_n316));
  NAND2_X1  g115(.A1(G155gat), .A2(G162gat), .ZN(new_n317));
  AOI22_X1  g116(.A1(new_n314), .A2(new_n316), .B1(KEYINPUT2), .B2(new_n317), .ZN(new_n318));
  OAI21_X1  g117(.A(KEYINPUT75), .B1(G155gat), .B2(G162gat), .ZN(new_n319));
  INV_X1    g118(.A(new_n319), .ZN(new_n320));
  NOR3_X1   g119(.A1(KEYINPUT75), .A2(G155gat), .A3(G162gat), .ZN(new_n321));
  OAI21_X1  g120(.A(new_n317), .B1(new_n320), .B2(new_n321), .ZN(new_n322));
  NAND2_X1  g121(.A1(new_n322), .A2(KEYINPUT76), .ZN(new_n323));
  INV_X1    g122(.A(new_n317), .ZN(new_n324));
  NOR2_X1   g123(.A1(G155gat), .A2(G162gat), .ZN(new_n325));
  INV_X1    g124(.A(KEYINPUT75), .ZN(new_n326));
  NAND2_X1  g125(.A1(new_n325), .A2(new_n326), .ZN(new_n327));
  AOI21_X1  g126(.A(new_n324), .B1(new_n327), .B2(new_n319), .ZN(new_n328));
  INV_X1    g127(.A(KEYINPUT76), .ZN(new_n329));
  NAND2_X1  g128(.A1(new_n328), .A2(new_n329), .ZN(new_n330));
  AOI21_X1  g129(.A(new_n318), .B1(new_n323), .B2(new_n330), .ZN(new_n331));
  NAND2_X1  g130(.A1(new_n314), .A2(new_n316), .ZN(new_n332));
  INV_X1    g131(.A(KEYINPUT2), .ZN(new_n333));
  OAI21_X1  g132(.A(new_n332), .B1(new_n333), .B2(new_n324), .ZN(new_n334));
  NOR3_X1   g133(.A1(new_n334), .A2(new_n324), .A3(new_n325), .ZN(new_n335));
  OAI21_X1  g134(.A(new_n312), .B1(new_n331), .B2(new_n335), .ZN(new_n336));
  INV_X1    g135(.A(KEYINPUT29), .ZN(new_n337));
  NAND2_X1  g136(.A1(new_n336), .A2(new_n337), .ZN(new_n338));
  INV_X1    g137(.A(KEYINPUT22), .ZN(new_n339));
  XNOR2_X1  g138(.A(KEYINPUT74), .B(G218gat), .ZN(new_n340));
  INV_X1    g139(.A(G211gat), .ZN(new_n341));
  OAI21_X1  g140(.A(new_n339), .B1(new_n340), .B2(new_n341), .ZN(new_n342));
  XNOR2_X1  g141(.A(G197gat), .B(G204gat), .ZN(new_n343));
  NAND2_X1  g142(.A1(new_n342), .A2(new_n343), .ZN(new_n344));
  INV_X1    g143(.A(new_n344), .ZN(new_n345));
  XNOR2_X1  g144(.A(G211gat), .B(G218gat), .ZN(new_n346));
  NAND2_X1  g145(.A1(new_n345), .A2(new_n346), .ZN(new_n347));
  INV_X1    g146(.A(new_n346), .ZN(new_n348));
  NAND2_X1  g147(.A1(new_n344), .A2(new_n348), .ZN(new_n349));
  NAND2_X1  g148(.A1(new_n347), .A2(new_n349), .ZN(new_n350));
  INV_X1    g149(.A(new_n350), .ZN(new_n351));
  NAND2_X1  g150(.A1(new_n338), .A2(new_n351), .ZN(new_n352));
  NOR2_X1   g151(.A1(new_n328), .A2(new_n329), .ZN(new_n353));
  AOI211_X1 g152(.A(KEYINPUT76), .B(new_n324), .C1(new_n327), .C2(new_n319), .ZN(new_n354));
  OAI21_X1  g153(.A(new_n334), .B1(new_n353), .B2(new_n354), .ZN(new_n355));
  OR3_X1    g154(.A1(new_n334), .A2(new_n324), .A3(new_n325), .ZN(new_n356));
  NAND2_X1  g155(.A1(new_n355), .A2(new_n356), .ZN(new_n357));
  INV_X1    g156(.A(new_n357), .ZN(new_n358));
  AOI21_X1  g157(.A(KEYINPUT29), .B1(new_n347), .B2(new_n349), .ZN(new_n359));
  OAI21_X1  g158(.A(new_n358), .B1(new_n359), .B2(KEYINPUT3), .ZN(new_n360));
  AND2_X1   g159(.A1(G228gat), .A2(G233gat), .ZN(new_n361));
  AND3_X1   g160(.A1(new_n352), .A2(new_n360), .A3(new_n361), .ZN(new_n362));
  AOI21_X1  g161(.A(new_n361), .B1(new_n352), .B2(new_n360), .ZN(new_n363));
  OAI21_X1  g162(.A(G22gat), .B1(new_n362), .B2(new_n363), .ZN(new_n364));
  INV_X1    g163(.A(KEYINPUT80), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n364), .A2(new_n365), .ZN(new_n366));
  XNOR2_X1  g165(.A(KEYINPUT79), .B(KEYINPUT31), .ZN(new_n367));
  INV_X1    g166(.A(G50gat), .ZN(new_n368));
  XNOR2_X1  g167(.A(new_n367), .B(new_n368), .ZN(new_n369));
  XOR2_X1   g168(.A(G78gat), .B(G106gat), .Z(new_n370));
  XNOR2_X1  g169(.A(new_n369), .B(new_n370), .ZN(new_n371));
  NAND2_X1  g170(.A1(new_n366), .A2(new_n371), .ZN(new_n372));
  OR3_X1    g171(.A1(new_n362), .A2(new_n363), .A3(G22gat), .ZN(new_n373));
  NAND2_X1  g172(.A1(new_n373), .A2(new_n364), .ZN(new_n374));
  NOR2_X1   g173(.A1(new_n372), .A2(new_n374), .ZN(new_n375));
  AOI22_X1  g174(.A1(new_n366), .A2(new_n371), .B1(new_n373), .B2(new_n364), .ZN(new_n376));
  NOR2_X1   g175(.A1(new_n375), .A2(new_n376), .ZN(new_n377));
  XNOR2_X1  g176(.A(G8gat), .B(G36gat), .ZN(new_n378));
  XNOR2_X1  g177(.A(G64gat), .B(G92gat), .ZN(new_n379));
  XOR2_X1   g178(.A(new_n378), .B(new_n379), .Z(new_n380));
  INV_X1    g179(.A(new_n380), .ZN(new_n381));
  INV_X1    g180(.A(G226gat), .ZN(new_n382));
  INV_X1    g181(.A(G233gat), .ZN(new_n383));
  NOR2_X1   g182(.A1(new_n382), .A2(new_n383), .ZN(new_n384));
  AOI21_X1  g183(.A(new_n384), .B1(new_n245), .B2(new_n337), .ZN(new_n385));
  INV_X1    g184(.A(new_n384), .ZN(new_n386));
  AOI21_X1  g185(.A(new_n386), .B1(new_n232), .B2(new_n244), .ZN(new_n387));
  NOR3_X1   g186(.A1(new_n385), .A2(new_n351), .A3(new_n387), .ZN(new_n388));
  AOI22_X1  g187(.A1(new_n217), .A2(new_n218), .B1(new_n230), .B2(KEYINPUT69), .ZN(new_n389));
  AOI22_X1  g188(.A1(new_n389), .A2(new_n229), .B1(new_n243), .B2(new_n240), .ZN(new_n390));
  OAI21_X1  g189(.A(new_n386), .B1(new_n390), .B2(KEYINPUT29), .ZN(new_n391));
  INV_X1    g190(.A(new_n387), .ZN(new_n392));
  AOI21_X1  g191(.A(new_n350), .B1(new_n391), .B2(new_n392), .ZN(new_n393));
  OAI21_X1  g192(.A(new_n381), .B1(new_n388), .B2(new_n393), .ZN(new_n394));
  OAI21_X1  g193(.A(new_n351), .B1(new_n385), .B2(new_n387), .ZN(new_n395));
  NAND3_X1  g194(.A1(new_n391), .A2(new_n350), .A3(new_n392), .ZN(new_n396));
  NAND3_X1  g195(.A1(new_n395), .A2(new_n396), .A3(new_n380), .ZN(new_n397));
  NAND3_X1  g196(.A1(new_n394), .A2(KEYINPUT30), .A3(new_n397), .ZN(new_n398));
  INV_X1    g197(.A(KEYINPUT30), .ZN(new_n399));
  NAND4_X1  g198(.A1(new_n395), .A2(new_n396), .A3(new_n399), .A4(new_n380), .ZN(new_n400));
  NAND2_X1  g199(.A1(new_n398), .A2(new_n400), .ZN(new_n401));
  INV_X1    g200(.A(KEYINPUT5), .ZN(new_n402));
  OAI21_X1  g201(.A(new_n262), .B1(new_n331), .B2(new_n335), .ZN(new_n403));
  AND2_X1   g202(.A1(new_n259), .A2(new_n261), .ZN(new_n404));
  NAND3_X1  g203(.A1(new_n404), .A2(new_n355), .A3(new_n356), .ZN(new_n405));
  NAND2_X1  g204(.A1(new_n403), .A2(new_n405), .ZN(new_n406));
  NAND2_X1  g205(.A1(G225gat), .A2(G233gat), .ZN(new_n407));
  INV_X1    g206(.A(new_n407), .ZN(new_n408));
  AOI21_X1  g207(.A(new_n402), .B1(new_n406), .B2(new_n408), .ZN(new_n409));
  NAND3_X1  g208(.A1(new_n357), .A2(new_n265), .A3(new_n264), .ZN(new_n410));
  XNOR2_X1  g209(.A(KEYINPUT77), .B(KEYINPUT4), .ZN(new_n411));
  INV_X1    g210(.A(new_n411), .ZN(new_n412));
  INV_X1    g211(.A(KEYINPUT4), .ZN(new_n413));
  AOI22_X1  g212(.A1(new_n355), .A2(new_n356), .B1(new_n261), .B2(new_n259), .ZN(new_n414));
  AOI22_X1  g213(.A1(new_n410), .A2(new_n412), .B1(new_n413), .B2(new_n414), .ZN(new_n415));
  NAND3_X1  g214(.A1(new_n355), .A2(new_n356), .A3(KEYINPUT3), .ZN(new_n416));
  NAND3_X1  g215(.A1(new_n336), .A2(new_n416), .A3(new_n404), .ZN(new_n417));
  NAND2_X1  g216(.A1(new_n417), .A2(new_n407), .ZN(new_n418));
  OAI21_X1  g217(.A(new_n409), .B1(new_n415), .B2(new_n418), .ZN(new_n419));
  OAI22_X1  g218(.A1(new_n410), .A2(new_n412), .B1(new_n413), .B2(new_n414), .ZN(new_n420));
  NAND4_X1  g219(.A1(new_n420), .A2(new_n402), .A3(new_n407), .A4(new_n417), .ZN(new_n421));
  NAND2_X1  g220(.A1(new_n419), .A2(new_n421), .ZN(new_n422));
  XNOR2_X1  g221(.A(G1gat), .B(G29gat), .ZN(new_n423));
  XNOR2_X1  g222(.A(new_n423), .B(KEYINPUT0), .ZN(new_n424));
  XNOR2_X1  g223(.A(G57gat), .B(G85gat), .ZN(new_n425));
  XOR2_X1   g224(.A(new_n424), .B(new_n425), .Z(new_n426));
  INV_X1    g225(.A(new_n426), .ZN(new_n427));
  NAND2_X1  g226(.A1(new_n422), .A2(new_n427), .ZN(new_n428));
  INV_X1    g227(.A(KEYINPUT6), .ZN(new_n429));
  NAND3_X1  g228(.A1(new_n419), .A2(new_n421), .A3(new_n426), .ZN(new_n430));
  NAND3_X1  g229(.A1(new_n428), .A2(new_n429), .A3(new_n430), .ZN(new_n431));
  NAND3_X1  g230(.A1(new_n422), .A2(KEYINPUT6), .A3(new_n427), .ZN(new_n432));
  NAND2_X1  g231(.A1(new_n431), .A2(new_n432), .ZN(new_n433));
  NAND2_X1  g232(.A1(new_n401), .A2(new_n433), .ZN(new_n434));
  INV_X1    g233(.A(KEYINPUT78), .ZN(new_n435));
  NAND2_X1  g234(.A1(new_n434), .A2(new_n435), .ZN(new_n436));
  NAND3_X1  g235(.A1(new_n401), .A2(new_n433), .A3(KEYINPUT78), .ZN(new_n437));
  AOI21_X1  g236(.A(new_n377), .B1(new_n436), .B2(new_n437), .ZN(new_n438));
  NOR2_X1   g237(.A1(new_n311), .A2(new_n438), .ZN(new_n439));
  INV_X1    g238(.A(KEYINPUT40), .ZN(new_n440));
  AOI21_X1  g239(.A(new_n407), .B1(new_n420), .B2(new_n417), .ZN(new_n441));
  NAND3_X1  g240(.A1(new_n403), .A2(new_n405), .A3(new_n407), .ZN(new_n442));
  INV_X1    g241(.A(KEYINPUT82), .ZN(new_n443));
  AND3_X1   g242(.A1(new_n442), .A2(new_n443), .A3(KEYINPUT39), .ZN(new_n444));
  AOI21_X1  g243(.A(new_n443), .B1(new_n442), .B2(KEYINPUT39), .ZN(new_n445));
  NOR3_X1   g244(.A1(new_n441), .A2(new_n444), .A3(new_n445), .ZN(new_n446));
  AND4_X1   g245(.A1(new_n357), .A2(new_n265), .A3(new_n264), .A4(new_n411), .ZN(new_n447));
  NOR2_X1   g246(.A1(new_n414), .A2(new_n413), .ZN(new_n448));
  OAI21_X1  g247(.A(new_n417), .B1(new_n447), .B2(new_n448), .ZN(new_n449));
  INV_X1    g248(.A(KEYINPUT39), .ZN(new_n450));
  NAND3_X1  g249(.A1(new_n449), .A2(new_n450), .A3(new_n408), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n451), .A2(new_n426), .ZN(new_n452));
  OAI21_X1  g251(.A(new_n440), .B1(new_n446), .B2(new_n452), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n453), .A2(new_n428), .ZN(new_n454));
  OR3_X1    g253(.A1(new_n441), .A2(new_n444), .A3(new_n445), .ZN(new_n455));
  AOI21_X1  g254(.A(new_n427), .B1(new_n441), .B2(new_n450), .ZN(new_n456));
  NAND3_X1  g255(.A1(new_n455), .A2(KEYINPUT40), .A3(new_n456), .ZN(new_n457));
  INV_X1    g256(.A(KEYINPUT83), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  NAND4_X1  g258(.A1(new_n455), .A2(KEYINPUT83), .A3(KEYINPUT40), .A4(new_n456), .ZN(new_n460));
  AOI21_X1  g259(.A(new_n454), .B1(new_n459), .B2(new_n460), .ZN(new_n461));
  INV_X1    g260(.A(KEYINPUT81), .ZN(new_n462));
  NOR2_X1   g261(.A1(new_n401), .A2(new_n462), .ZN(new_n463));
  AOI21_X1  g262(.A(KEYINPUT81), .B1(new_n398), .B2(new_n400), .ZN(new_n464));
  OAI21_X1  g263(.A(new_n461), .B1(new_n463), .B2(new_n464), .ZN(new_n465));
  OAI21_X1  g264(.A(KEYINPUT37), .B1(new_n388), .B2(new_n393), .ZN(new_n466));
  INV_X1    g265(.A(KEYINPUT38), .ZN(new_n467));
  INV_X1    g266(.A(KEYINPUT37), .ZN(new_n468));
  NAND3_X1  g267(.A1(new_n395), .A2(new_n468), .A3(new_n396), .ZN(new_n469));
  NAND4_X1  g268(.A1(new_n466), .A2(new_n467), .A3(new_n469), .A4(new_n381), .ZN(new_n470));
  NAND4_X1  g269(.A1(new_n470), .A2(new_n432), .A3(new_n431), .A4(new_n397), .ZN(new_n471));
  AND3_X1   g270(.A1(new_n466), .A2(new_n469), .A3(new_n381), .ZN(new_n472));
  OAI22_X1  g271(.A1(new_n471), .A2(KEYINPUT84), .B1(new_n467), .B2(new_n472), .ZN(new_n473));
  AND2_X1   g272(.A1(new_n471), .A2(KEYINPUT84), .ZN(new_n474));
  OAI211_X1 g273(.A(new_n465), .B(new_n377), .C1(new_n473), .C2(new_n474), .ZN(new_n475));
  NAND2_X1  g274(.A1(new_n436), .A2(new_n437), .ZN(new_n476));
  NOR3_X1   g275(.A1(new_n288), .A2(new_n289), .A3(new_n277), .ZN(new_n477));
  AOI21_X1  g276(.A(new_n298), .B1(new_n297), .B2(new_n300), .ZN(new_n478));
  OAI21_X1  g277(.A(new_n309), .B1(new_n477), .B2(new_n478), .ZN(new_n479));
  INV_X1    g278(.A(new_n307), .ZN(new_n480));
  NAND3_X1  g279(.A1(new_n479), .A2(new_n377), .A3(new_n480), .ZN(new_n481));
  OAI21_X1  g280(.A(KEYINPUT35), .B1(new_n476), .B2(new_n481), .ZN(new_n482));
  INV_X1    g281(.A(new_n433), .ZN(new_n483));
  NOR4_X1   g282(.A1(new_n483), .A2(new_n375), .A3(new_n376), .A4(KEYINPUT35), .ZN(new_n484));
  INV_X1    g283(.A(new_n463), .ZN(new_n485));
  INV_X1    g284(.A(new_n464), .ZN(new_n486));
  NAND4_X1  g285(.A1(new_n484), .A2(new_n485), .A3(new_n486), .A4(new_n303), .ZN(new_n487));
  AOI22_X1  g286(.A1(new_n439), .A2(new_n475), .B1(new_n482), .B2(new_n487), .ZN(new_n488));
  NAND2_X1  g287(.A1(G229gat), .A2(G233gat), .ZN(new_n489));
  XNOR2_X1  g288(.A(new_n489), .B(KEYINPUT13), .ZN(new_n490));
  XNOR2_X1  g289(.A(G15gat), .B(G22gat), .ZN(new_n491));
  NOR2_X1   g290(.A1(new_n491), .A2(G1gat), .ZN(new_n492));
  INV_X1    g291(.A(KEYINPUT86), .ZN(new_n493));
  OAI21_X1  g292(.A(G8gat), .B1(new_n492), .B2(new_n493), .ZN(new_n494));
  INV_X1    g293(.A(KEYINPUT16), .ZN(new_n495));
  OAI21_X1  g294(.A(new_n491), .B1(new_n495), .B2(G1gat), .ZN(new_n496));
  OAI21_X1  g295(.A(new_n496), .B1(G1gat), .B2(new_n491), .ZN(new_n497));
  XNOR2_X1  g296(.A(new_n494), .B(new_n497), .ZN(new_n498));
  INV_X1    g297(.A(new_n498), .ZN(new_n499));
  NOR2_X1   g298(.A1(G29gat), .A2(G36gat), .ZN(new_n500));
  XNOR2_X1  g299(.A(new_n500), .B(KEYINPUT14), .ZN(new_n501));
  INV_X1    g300(.A(new_n501), .ZN(new_n502));
  XNOR2_X1  g301(.A(G43gat), .B(G50gat), .ZN(new_n503));
  OR2_X1    g302(.A1(new_n503), .A2(KEYINPUT15), .ZN(new_n504));
  NAND2_X1  g303(.A1(G29gat), .A2(G36gat), .ZN(new_n505));
  INV_X1    g304(.A(KEYINPUT85), .ZN(new_n506));
  XNOR2_X1  g305(.A(new_n505), .B(new_n506), .ZN(new_n507));
  NAND2_X1  g306(.A1(new_n503), .A2(KEYINPUT15), .ZN(new_n508));
  NAND4_X1  g307(.A1(new_n502), .A2(new_n504), .A3(new_n507), .A4(new_n508), .ZN(new_n509));
  INV_X1    g308(.A(new_n505), .ZN(new_n510));
  OAI211_X1 g309(.A(KEYINPUT15), .B(new_n503), .C1(new_n501), .C2(new_n510), .ZN(new_n511));
  NAND2_X1  g310(.A1(new_n509), .A2(new_n511), .ZN(new_n512));
  NAND2_X1  g311(.A1(new_n499), .A2(new_n512), .ZN(new_n513));
  NAND3_X1  g312(.A1(new_n498), .A2(new_n511), .A3(new_n509), .ZN(new_n514));
  AOI21_X1  g313(.A(new_n490), .B1(new_n513), .B2(new_n514), .ZN(new_n515));
  INV_X1    g314(.A(KEYINPUT17), .ZN(new_n516));
  NAND3_X1  g315(.A1(new_n509), .A2(new_n516), .A3(new_n511), .ZN(new_n517));
  INV_X1    g316(.A(new_n517), .ZN(new_n518));
  AOI21_X1  g317(.A(new_n516), .B1(new_n509), .B2(new_n511), .ZN(new_n519));
  OAI21_X1  g318(.A(new_n498), .B1(new_n518), .B2(new_n519), .ZN(new_n520));
  NAND3_X1  g319(.A1(new_n513), .A2(new_n520), .A3(new_n489), .ZN(new_n521));
  INV_X1    g320(.A(KEYINPUT18), .ZN(new_n522));
  AOI21_X1  g321(.A(new_n515), .B1(new_n521), .B2(new_n522), .ZN(new_n523));
  NAND4_X1  g322(.A1(new_n513), .A2(new_n520), .A3(KEYINPUT18), .A4(new_n489), .ZN(new_n524));
  INV_X1    g323(.A(KEYINPUT87), .ZN(new_n525));
  AND2_X1   g324(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  NOR2_X1   g325(.A1(new_n524), .A2(new_n525), .ZN(new_n527));
  OAI21_X1  g326(.A(new_n523), .B1(new_n526), .B2(new_n527), .ZN(new_n528));
  XNOR2_X1  g327(.A(G113gat), .B(G141gat), .ZN(new_n529));
  XNOR2_X1  g328(.A(new_n529), .B(G197gat), .ZN(new_n530));
  XOR2_X1   g329(.A(KEYINPUT11), .B(G169gat), .Z(new_n531));
  XNOR2_X1  g330(.A(new_n530), .B(new_n531), .ZN(new_n532));
  XNOR2_X1  g331(.A(new_n532), .B(KEYINPUT12), .ZN(new_n533));
  INV_X1    g332(.A(new_n533), .ZN(new_n534));
  NAND2_X1  g333(.A1(new_n528), .A2(new_n534), .ZN(new_n535));
  OAI211_X1 g334(.A(new_n523), .B(new_n533), .C1(new_n526), .C2(new_n527), .ZN(new_n536));
  NAND2_X1  g335(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  INV_X1    g336(.A(new_n537), .ZN(new_n538));
  NOR2_X1   g337(.A1(new_n488), .A2(new_n538), .ZN(new_n539));
  NAND2_X1  g338(.A1(G99gat), .A2(G106gat), .ZN(new_n540));
  INV_X1    g339(.A(KEYINPUT95), .ZN(new_n541));
  NAND2_X1  g340(.A1(new_n540), .A2(new_n541), .ZN(new_n542));
  NAND3_X1  g341(.A1(KEYINPUT95), .A2(G99gat), .A3(G106gat), .ZN(new_n543));
  NAND3_X1  g342(.A1(new_n542), .A2(KEYINPUT8), .A3(new_n543), .ZN(new_n544));
  NAND2_X1  g343(.A1(G85gat), .A2(G92gat), .ZN(new_n545));
  INV_X1    g344(.A(new_n545), .ZN(new_n546));
  INV_X1    g345(.A(KEYINPUT94), .ZN(new_n547));
  NAND2_X1  g346(.A1(new_n547), .A2(KEYINPUT7), .ZN(new_n548));
  INV_X1    g347(.A(KEYINPUT7), .ZN(new_n549));
  NAND2_X1  g348(.A1(new_n549), .A2(KEYINPUT94), .ZN(new_n550));
  NAND3_X1  g349(.A1(new_n546), .A2(new_n548), .A3(new_n550), .ZN(new_n551));
  INV_X1    g350(.A(G85gat), .ZN(new_n552));
  NAND2_X1  g351(.A1(new_n552), .A2(KEYINPUT96), .ZN(new_n553));
  INV_X1    g352(.A(KEYINPUT96), .ZN(new_n554));
  NAND2_X1  g353(.A1(new_n554), .A2(G85gat), .ZN(new_n555));
  INV_X1    g354(.A(G92gat), .ZN(new_n556));
  NAND3_X1  g355(.A1(new_n553), .A2(new_n555), .A3(new_n556), .ZN(new_n557));
  NOR2_X1   g356(.A1(new_n547), .A2(KEYINPUT7), .ZN(new_n558));
  NAND2_X1  g357(.A1(new_n558), .A2(new_n545), .ZN(new_n559));
  NAND4_X1  g358(.A1(new_n544), .A2(new_n551), .A3(new_n557), .A4(new_n559), .ZN(new_n560));
  XOR2_X1   g359(.A(G99gat), .B(G106gat), .Z(new_n561));
  NAND2_X1  g360(.A1(new_n560), .A2(new_n561), .ZN(new_n562));
  XNOR2_X1  g361(.A(KEYINPUT96), .B(G85gat), .ZN(new_n563));
  AOI22_X1  g362(.A1(new_n563), .A2(new_n556), .B1(new_n545), .B2(new_n558), .ZN(new_n564));
  INV_X1    g363(.A(new_n561), .ZN(new_n565));
  NAND4_X1  g364(.A1(new_n564), .A2(new_n565), .A3(new_n544), .A4(new_n551), .ZN(new_n566));
  NAND3_X1  g365(.A1(new_n562), .A2(new_n566), .A3(KEYINPUT97), .ZN(new_n567));
  INV_X1    g366(.A(KEYINPUT97), .ZN(new_n568));
  NAND3_X1  g367(.A1(new_n560), .A2(new_n568), .A3(new_n561), .ZN(new_n569));
  AND2_X1   g368(.A1(new_n567), .A2(new_n569), .ZN(new_n570));
  OAI21_X1  g369(.A(new_n570), .B1(new_n519), .B2(new_n518), .ZN(new_n571));
  NAND3_X1  g370(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n572));
  INV_X1    g371(.A(new_n512), .ZN(new_n573));
  OAI211_X1 g372(.A(new_n571), .B(new_n572), .C1(new_n573), .C2(new_n570), .ZN(new_n574));
  XNOR2_X1  g373(.A(G190gat), .B(G218gat), .ZN(new_n575));
  XNOR2_X1  g374(.A(new_n575), .B(KEYINPUT98), .ZN(new_n576));
  OR2_X1    g375(.A1(new_n574), .A2(new_n576), .ZN(new_n577));
  AOI21_X1  g376(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n578));
  XNOR2_X1  g377(.A(new_n578), .B(KEYINPUT93), .ZN(new_n579));
  XNOR2_X1  g378(.A(G134gat), .B(G162gat), .ZN(new_n580));
  XNOR2_X1  g379(.A(new_n579), .B(new_n580), .ZN(new_n581));
  NAND2_X1  g380(.A1(new_n574), .A2(new_n576), .ZN(new_n582));
  AND3_X1   g381(.A1(new_n577), .A2(new_n581), .A3(new_n582), .ZN(new_n583));
  AOI21_X1  g382(.A(new_n581), .B1(new_n577), .B2(new_n582), .ZN(new_n584));
  NOR2_X1   g383(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  INV_X1    g384(.A(new_n585), .ZN(new_n586));
  NAND2_X1  g385(.A1(G71gat), .A2(G78gat), .ZN(new_n587));
  INV_X1    g386(.A(KEYINPUT9), .ZN(new_n588));
  NAND2_X1  g387(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  NAND2_X1  g388(.A1(new_n589), .A2(KEYINPUT88), .ZN(new_n590));
  INV_X1    g389(.A(KEYINPUT88), .ZN(new_n591));
  NAND3_X1  g390(.A1(new_n587), .A2(new_n591), .A3(new_n588), .ZN(new_n592));
  INV_X1    g391(.A(G57gat), .ZN(new_n593));
  NAND2_X1  g392(.A1(new_n593), .A2(G64gat), .ZN(new_n594));
  INV_X1    g393(.A(G64gat), .ZN(new_n595));
  NAND2_X1  g394(.A1(new_n595), .A2(G57gat), .ZN(new_n596));
  NAND2_X1  g395(.A1(new_n594), .A2(new_n596), .ZN(new_n597));
  NAND3_X1  g396(.A1(new_n590), .A2(new_n592), .A3(new_n597), .ZN(new_n598));
  XNOR2_X1  g397(.A(G71gat), .B(G78gat), .ZN(new_n599));
  INV_X1    g398(.A(new_n599), .ZN(new_n600));
  NAND2_X1  g399(.A1(new_n598), .A2(new_n600), .ZN(new_n601));
  INV_X1    g400(.A(KEYINPUT89), .ZN(new_n602));
  OAI21_X1  g401(.A(new_n602), .B1(new_n595), .B2(G57gat), .ZN(new_n603));
  NAND3_X1  g402(.A1(new_n593), .A2(KEYINPUT89), .A3(G64gat), .ZN(new_n604));
  NAND3_X1  g403(.A1(new_n603), .A2(new_n596), .A3(new_n604), .ZN(new_n605));
  NAND4_X1  g404(.A1(new_n605), .A2(new_n599), .A3(new_n592), .A4(new_n590), .ZN(new_n606));
  NAND2_X1  g405(.A1(new_n601), .A2(new_n606), .ZN(new_n607));
  NAND2_X1  g406(.A1(new_n607), .A2(KEYINPUT90), .ZN(new_n608));
  INV_X1    g407(.A(KEYINPUT90), .ZN(new_n609));
  NAND3_X1  g408(.A1(new_n601), .A2(new_n609), .A3(new_n606), .ZN(new_n610));
  NAND2_X1  g409(.A1(new_n608), .A2(new_n610), .ZN(new_n611));
  AOI21_X1  g410(.A(new_n499), .B1(new_n611), .B2(KEYINPUT21), .ZN(new_n612));
  XNOR2_X1  g411(.A(new_n612), .B(KEYINPUT92), .ZN(new_n613));
  XNOR2_X1  g412(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n614));
  XNOR2_X1  g413(.A(new_n614), .B(KEYINPUT91), .ZN(new_n615));
  XNOR2_X1  g414(.A(new_n615), .B(G155gat), .ZN(new_n616));
  XNOR2_X1  g415(.A(new_n613), .B(new_n616), .ZN(new_n617));
  INV_X1    g416(.A(new_n617), .ZN(new_n618));
  XNOR2_X1  g417(.A(G183gat), .B(G211gat), .ZN(new_n619));
  OR2_X1    g418(.A1(new_n611), .A2(KEYINPUT21), .ZN(new_n620));
  NAND2_X1  g419(.A1(G231gat), .A2(G233gat), .ZN(new_n621));
  XNOR2_X1  g420(.A(new_n620), .B(new_n621), .ZN(new_n622));
  AND2_X1   g421(.A1(new_n622), .A2(new_n254), .ZN(new_n623));
  NOR2_X1   g422(.A1(new_n622), .A2(new_n254), .ZN(new_n624));
  OAI21_X1  g423(.A(new_n619), .B1(new_n623), .B2(new_n624), .ZN(new_n625));
  INV_X1    g424(.A(new_n625), .ZN(new_n626));
  NOR3_X1   g425(.A1(new_n623), .A2(new_n624), .A3(new_n619), .ZN(new_n627));
  OAI21_X1  g426(.A(new_n618), .B1(new_n626), .B2(new_n627), .ZN(new_n628));
  INV_X1    g427(.A(new_n627), .ZN(new_n629));
  NAND3_X1  g428(.A1(new_n629), .A2(new_n625), .A3(new_n617), .ZN(new_n630));
  AOI21_X1  g429(.A(new_n586), .B1(new_n628), .B2(new_n630), .ZN(new_n631));
  INV_X1    g430(.A(new_n631), .ZN(new_n632));
  NAND2_X1  g431(.A1(G230gat), .A2(G233gat), .ZN(new_n633));
  INV_X1    g432(.A(new_n607), .ZN(new_n634));
  NAND3_X1  g433(.A1(new_n634), .A2(new_n562), .A3(new_n566), .ZN(new_n635));
  INV_X1    g434(.A(new_n635), .ZN(new_n636));
  NAND4_X1  g435(.A1(new_n608), .A2(new_n567), .A3(new_n610), .A4(new_n569), .ZN(new_n637));
  NAND2_X1  g436(.A1(new_n637), .A2(KEYINPUT99), .ZN(new_n638));
  AND3_X1   g437(.A1(new_n601), .A2(new_n609), .A3(new_n606), .ZN(new_n639));
  AOI21_X1  g438(.A(new_n609), .B1(new_n601), .B2(new_n606), .ZN(new_n640));
  NOR2_X1   g439(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  INV_X1    g440(.A(KEYINPUT99), .ZN(new_n642));
  NAND4_X1  g441(.A1(new_n641), .A2(new_n642), .A3(new_n569), .A4(new_n567), .ZN(new_n643));
  AOI211_X1 g442(.A(KEYINPUT10), .B(new_n636), .C1(new_n638), .C2(new_n643), .ZN(new_n644));
  INV_X1    g443(.A(KEYINPUT10), .ZN(new_n645));
  NOR3_X1   g444(.A1(new_n570), .A2(new_n641), .A3(new_n645), .ZN(new_n646));
  OAI21_X1  g445(.A(new_n633), .B1(new_n644), .B2(new_n646), .ZN(new_n647));
  AOI21_X1  g446(.A(new_n636), .B1(new_n638), .B2(new_n643), .ZN(new_n648));
  NOR2_X1   g447(.A1(new_n648), .A2(new_n633), .ZN(new_n649));
  INV_X1    g448(.A(KEYINPUT100), .ZN(new_n650));
  NAND2_X1  g449(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  OAI21_X1  g450(.A(KEYINPUT100), .B1(new_n648), .B2(new_n633), .ZN(new_n652));
  NAND3_X1  g451(.A1(new_n647), .A2(new_n651), .A3(new_n652), .ZN(new_n653));
  XOR2_X1   g452(.A(G120gat), .B(G148gat), .Z(new_n654));
  XNOR2_X1  g453(.A(new_n654), .B(KEYINPUT101), .ZN(new_n655));
  XNOR2_X1  g454(.A(G176gat), .B(G204gat), .ZN(new_n656));
  XOR2_X1   g455(.A(new_n655), .B(new_n656), .Z(new_n657));
  INV_X1    g456(.A(new_n657), .ZN(new_n658));
  NAND2_X1  g457(.A1(new_n653), .A2(new_n658), .ZN(new_n659));
  NAND4_X1  g458(.A1(new_n647), .A2(new_n651), .A3(new_n657), .A4(new_n652), .ZN(new_n660));
  NAND2_X1  g459(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  NOR2_X1   g460(.A1(new_n632), .A2(new_n661), .ZN(new_n662));
  NAND2_X1  g461(.A1(new_n539), .A2(new_n662), .ZN(new_n663));
  INV_X1    g462(.A(new_n663), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n664), .A2(new_n483), .ZN(new_n665));
  XNOR2_X1  g464(.A(new_n665), .B(G1gat), .ZN(G1324gat));
  NAND2_X1  g465(.A1(new_n485), .A2(new_n486), .ZN(new_n667));
  NAND2_X1  g466(.A1(new_n664), .A2(new_n667), .ZN(new_n668));
  AND2_X1   g467(.A1(new_n668), .A2(G8gat), .ZN(new_n669));
  XNOR2_X1  g468(.A(KEYINPUT16), .B(G8gat), .ZN(new_n670));
  NOR2_X1   g469(.A1(new_n668), .A2(new_n670), .ZN(new_n671));
  OAI21_X1  g470(.A(KEYINPUT42), .B1(new_n669), .B2(new_n671), .ZN(new_n672));
  OAI21_X1  g471(.A(new_n672), .B1(KEYINPUT42), .B2(new_n671), .ZN(G1325gat));
  NOR2_X1   g472(.A1(new_n302), .A2(KEYINPUT36), .ZN(new_n674));
  NAND2_X1  g473(.A1(new_n479), .A2(new_n480), .ZN(new_n675));
  AOI21_X1  g474(.A(new_n674), .B1(new_n675), .B2(KEYINPUT36), .ZN(new_n676));
  OAI21_X1  g475(.A(G15gat), .B1(new_n663), .B2(new_n676), .ZN(new_n677));
  OR2_X1    g476(.A1(new_n302), .A2(G15gat), .ZN(new_n678));
  OAI21_X1  g477(.A(new_n677), .B1(new_n663), .B2(new_n678), .ZN(G1326gat));
  NOR3_X1   g478(.A1(new_n488), .A2(new_n377), .A3(new_n538), .ZN(new_n680));
  NAND2_X1  g479(.A1(new_n680), .A2(new_n662), .ZN(new_n681));
  XNOR2_X1  g480(.A(KEYINPUT43), .B(G22gat), .ZN(new_n682));
  XNOR2_X1  g481(.A(new_n681), .B(new_n682), .ZN(G1327gat));
  NOR2_X1   g482(.A1(new_n488), .A2(new_n585), .ZN(new_n684));
  INV_X1    g483(.A(new_n684), .ZN(new_n685));
  NAND2_X1  g484(.A1(new_n628), .A2(new_n630), .ZN(new_n686));
  NOR2_X1   g485(.A1(new_n686), .A2(new_n661), .ZN(new_n687));
  NAND2_X1  g486(.A1(new_n687), .A2(new_n537), .ZN(new_n688));
  NOR4_X1   g487(.A1(new_n685), .A2(G29gat), .A3(new_n433), .A4(new_n688), .ZN(new_n689));
  XOR2_X1   g488(.A(new_n689), .B(KEYINPUT45), .Z(new_n690));
  INV_X1    g489(.A(KEYINPUT44), .ZN(new_n691));
  OAI21_X1  g490(.A(new_n691), .B1(new_n488), .B2(new_n585), .ZN(new_n692));
  INV_X1    g491(.A(new_n438), .ZN(new_n693));
  NAND3_X1  g492(.A1(new_n475), .A2(new_n693), .A3(new_n676), .ZN(new_n694));
  NAND2_X1  g493(.A1(new_n482), .A2(new_n487), .ZN(new_n695));
  NAND2_X1  g494(.A1(new_n694), .A2(new_n695), .ZN(new_n696));
  NAND3_X1  g495(.A1(new_n696), .A2(KEYINPUT44), .A3(new_n586), .ZN(new_n697));
  AND2_X1   g496(.A1(new_n692), .A2(new_n697), .ZN(new_n698));
  INV_X1    g497(.A(new_n688), .ZN(new_n699));
  NAND2_X1  g498(.A1(new_n698), .A2(new_n699), .ZN(new_n700));
  OAI21_X1  g499(.A(G29gat), .B1(new_n700), .B2(new_n433), .ZN(new_n701));
  NAND2_X1  g500(.A1(new_n690), .A2(new_n701), .ZN(G1328gat));
  INV_X1    g501(.A(new_n667), .ZN(new_n703));
  NOR4_X1   g502(.A1(new_n685), .A2(G36gat), .A3(new_n703), .A4(new_n688), .ZN(new_n704));
  XNOR2_X1  g503(.A(new_n704), .B(KEYINPUT46), .ZN(new_n705));
  OAI21_X1  g504(.A(G36gat), .B1(new_n700), .B2(new_n703), .ZN(new_n706));
  NAND2_X1  g505(.A1(new_n705), .A2(new_n706), .ZN(G1329gat));
  NAND3_X1  g506(.A1(new_n684), .A2(new_n303), .A3(new_n699), .ZN(new_n708));
  INV_X1    g507(.A(G43gat), .ZN(new_n709));
  INV_X1    g508(.A(KEYINPUT102), .ZN(new_n710));
  AOI22_X1  g509(.A1(new_n708), .A2(new_n709), .B1(new_n710), .B2(KEYINPUT47), .ZN(new_n711));
  NAND2_X1  g510(.A1(new_n311), .A2(G43gat), .ZN(new_n712));
  OAI21_X1  g511(.A(new_n711), .B1(new_n700), .B2(new_n712), .ZN(new_n713));
  NOR2_X1   g512(.A1(new_n710), .A2(KEYINPUT47), .ZN(new_n714));
  XOR2_X1   g513(.A(new_n713), .B(new_n714), .Z(G1330gat));
  OAI21_X1  g514(.A(G50gat), .B1(new_n700), .B2(new_n377), .ZN(new_n716));
  NAND4_X1  g515(.A1(new_n680), .A2(new_n368), .A3(new_n586), .A4(new_n687), .ZN(new_n717));
  NAND2_X1  g516(.A1(new_n716), .A2(new_n717), .ZN(new_n718));
  INV_X1    g517(.A(KEYINPUT48), .ZN(new_n719));
  XNOR2_X1  g518(.A(new_n718), .B(new_n719), .ZN(G1331gat));
  INV_X1    g519(.A(new_n661), .ZN(new_n721));
  NOR3_X1   g520(.A1(new_n632), .A2(new_n537), .A3(new_n721), .ZN(new_n722));
  NAND2_X1  g521(.A1(new_n696), .A2(new_n722), .ZN(new_n723));
  NOR2_X1   g522(.A1(new_n723), .A2(new_n433), .ZN(new_n724));
  XNOR2_X1  g523(.A(new_n724), .B(new_n593), .ZN(G1332gat));
  INV_X1    g524(.A(KEYINPUT103), .ZN(new_n726));
  XNOR2_X1  g525(.A(new_n723), .B(new_n726), .ZN(new_n727));
  AOI21_X1  g526(.A(new_n703), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n728));
  NAND2_X1  g527(.A1(new_n727), .A2(new_n728), .ZN(new_n729));
  NAND2_X1  g528(.A1(new_n729), .A2(KEYINPUT104), .ZN(new_n730));
  INV_X1    g529(.A(KEYINPUT104), .ZN(new_n731));
  NAND3_X1  g530(.A1(new_n727), .A2(new_n731), .A3(new_n728), .ZN(new_n732));
  NAND2_X1  g531(.A1(new_n730), .A2(new_n732), .ZN(new_n733));
  INV_X1    g532(.A(KEYINPUT49), .ZN(new_n734));
  NAND2_X1  g533(.A1(new_n734), .A2(new_n595), .ZN(new_n735));
  XNOR2_X1  g534(.A(new_n733), .B(new_n735), .ZN(G1333gat));
  NAND3_X1  g535(.A1(new_n727), .A2(G71gat), .A3(new_n311), .ZN(new_n737));
  OAI21_X1  g536(.A(new_n280), .B1(new_n723), .B2(new_n302), .ZN(new_n738));
  NAND2_X1  g537(.A1(new_n737), .A2(new_n738), .ZN(new_n739));
  XNOR2_X1  g538(.A(new_n739), .B(KEYINPUT50), .ZN(G1334gat));
  INV_X1    g539(.A(new_n377), .ZN(new_n741));
  NAND2_X1  g540(.A1(new_n727), .A2(new_n741), .ZN(new_n742));
  XNOR2_X1  g541(.A(new_n742), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g542(.A1(new_n686), .A2(new_n537), .ZN(new_n744));
  NAND3_X1  g543(.A1(new_n696), .A2(new_n586), .A3(new_n744), .ZN(new_n745));
  INV_X1    g544(.A(KEYINPUT51), .ZN(new_n746));
  NAND2_X1  g545(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  NAND4_X1  g546(.A1(new_n696), .A2(KEYINPUT51), .A3(new_n586), .A4(new_n744), .ZN(new_n748));
  AOI21_X1  g547(.A(new_n721), .B1(new_n747), .B2(new_n748), .ZN(new_n749));
  NAND3_X1  g548(.A1(new_n749), .A2(new_n483), .A3(new_n563), .ZN(new_n750));
  NOR3_X1   g549(.A1(new_n686), .A2(new_n537), .A3(new_n721), .ZN(new_n751));
  NAND3_X1  g550(.A1(new_n692), .A2(new_n697), .A3(new_n751), .ZN(new_n752));
  INV_X1    g551(.A(KEYINPUT105), .ZN(new_n753));
  NAND2_X1  g552(.A1(new_n752), .A2(new_n753), .ZN(new_n754));
  NAND4_X1  g553(.A1(new_n692), .A2(new_n697), .A3(KEYINPUT105), .A4(new_n751), .ZN(new_n755));
  AND3_X1   g554(.A1(new_n754), .A2(new_n483), .A3(new_n755), .ZN(new_n756));
  OAI21_X1  g555(.A(new_n750), .B1(new_n756), .B2(new_n563), .ZN(G1336gat));
  NAND3_X1  g556(.A1(new_n747), .A2(KEYINPUT106), .A3(new_n748), .ZN(new_n758));
  INV_X1    g557(.A(KEYINPUT106), .ZN(new_n759));
  NAND3_X1  g558(.A1(new_n745), .A2(new_n759), .A3(new_n746), .ZN(new_n760));
  AND2_X1   g559(.A1(new_n758), .A2(new_n760), .ZN(new_n761));
  NOR3_X1   g560(.A1(new_n703), .A2(G92gat), .A3(new_n721), .ZN(new_n762));
  NAND3_X1  g561(.A1(new_n754), .A2(new_n667), .A3(new_n755), .ZN(new_n763));
  AOI22_X1  g562(.A1(new_n761), .A2(new_n762), .B1(new_n763), .B2(G92gat), .ZN(new_n764));
  INV_X1    g563(.A(KEYINPUT52), .ZN(new_n765));
  NAND2_X1  g564(.A1(new_n747), .A2(new_n748), .ZN(new_n766));
  NAND2_X1  g565(.A1(new_n766), .A2(new_n762), .ZN(new_n767));
  NAND2_X1  g566(.A1(new_n767), .A2(new_n765), .ZN(new_n768));
  NOR2_X1   g567(.A1(new_n752), .A2(new_n703), .ZN(new_n769));
  NOR2_X1   g568(.A1(new_n769), .A2(new_n556), .ZN(new_n770));
  OAI22_X1  g569(.A1(new_n764), .A2(new_n765), .B1(new_n768), .B2(new_n770), .ZN(G1337gat));
  NAND3_X1  g570(.A1(new_n749), .A2(new_n282), .A3(new_n303), .ZN(new_n772));
  AND3_X1   g571(.A1(new_n754), .A2(new_n311), .A3(new_n755), .ZN(new_n773));
  OAI21_X1  g572(.A(new_n772), .B1(new_n773), .B2(new_n282), .ZN(G1338gat));
  NAND3_X1  g573(.A1(new_n754), .A2(new_n741), .A3(new_n755), .ZN(new_n775));
  XOR2_X1   g574(.A(KEYINPUT107), .B(G106gat), .Z(new_n776));
  NAND2_X1  g575(.A1(new_n775), .A2(new_n776), .ZN(new_n777));
  NOR3_X1   g576(.A1(new_n721), .A2(new_n377), .A3(G106gat), .ZN(new_n778));
  NAND4_X1  g577(.A1(new_n758), .A2(KEYINPUT108), .A3(new_n760), .A4(new_n778), .ZN(new_n779));
  NAND3_X1  g578(.A1(new_n758), .A2(new_n760), .A3(new_n778), .ZN(new_n780));
  INV_X1    g579(.A(KEYINPUT108), .ZN(new_n781));
  NAND2_X1  g580(.A1(new_n780), .A2(new_n781), .ZN(new_n782));
  NAND3_X1  g581(.A1(new_n777), .A2(new_n779), .A3(new_n782), .ZN(new_n783));
  NAND2_X1  g582(.A1(new_n783), .A2(KEYINPUT53), .ZN(new_n784));
  NOR2_X1   g583(.A1(new_n377), .A2(G106gat), .ZN(new_n785));
  AOI21_X1  g584(.A(KEYINPUT53), .B1(new_n749), .B2(new_n785), .ZN(new_n786));
  OAI21_X1  g585(.A(new_n776), .B1(new_n752), .B2(new_n377), .ZN(new_n787));
  NAND2_X1  g586(.A1(new_n786), .A2(new_n787), .ZN(new_n788));
  NAND2_X1  g587(.A1(new_n784), .A2(new_n788), .ZN(G1339gat));
  NAND3_X1  g588(.A1(new_n631), .A2(new_n538), .A3(new_n721), .ZN(new_n790));
  INV_X1    g589(.A(new_n790), .ZN(new_n791));
  AOI21_X1  g590(.A(new_n642), .B1(new_n570), .B2(new_n641), .ZN(new_n792));
  NOR2_X1   g591(.A1(new_n637), .A2(KEYINPUT99), .ZN(new_n793));
  OAI211_X1 g592(.A(new_n645), .B(new_n635), .C1(new_n792), .C2(new_n793), .ZN(new_n794));
  INV_X1    g593(.A(new_n633), .ZN(new_n795));
  INV_X1    g594(.A(new_n646), .ZN(new_n796));
  NAND3_X1  g595(.A1(new_n794), .A2(new_n795), .A3(new_n796), .ZN(new_n797));
  NAND3_X1  g596(.A1(new_n647), .A2(KEYINPUT54), .A3(new_n797), .ZN(new_n798));
  AOI21_X1  g597(.A(new_n795), .B1(new_n794), .B2(new_n796), .ZN(new_n799));
  INV_X1    g598(.A(KEYINPUT54), .ZN(new_n800));
  AOI21_X1  g599(.A(new_n657), .B1(new_n799), .B2(new_n800), .ZN(new_n801));
  NAND3_X1  g600(.A1(new_n798), .A2(new_n801), .A3(KEYINPUT55), .ZN(new_n802));
  NAND3_X1  g601(.A1(new_n802), .A2(new_n537), .A3(new_n660), .ZN(new_n803));
  INV_X1    g602(.A(KEYINPUT55), .ZN(new_n804));
  AND3_X1   g603(.A1(new_n647), .A2(KEYINPUT54), .A3(new_n797), .ZN(new_n805));
  OAI21_X1  g604(.A(new_n658), .B1(new_n647), .B2(KEYINPUT54), .ZN(new_n806));
  OAI21_X1  g605(.A(new_n804), .B1(new_n805), .B2(new_n806), .ZN(new_n807));
  INV_X1    g606(.A(KEYINPUT109), .ZN(new_n808));
  NAND2_X1  g607(.A1(new_n807), .A2(new_n808), .ZN(new_n809));
  AOI21_X1  g608(.A(KEYINPUT55), .B1(new_n798), .B2(new_n801), .ZN(new_n810));
  NAND2_X1  g609(.A1(new_n810), .A2(KEYINPUT109), .ZN(new_n811));
  AOI21_X1  g610(.A(new_n803), .B1(new_n809), .B2(new_n811), .ZN(new_n812));
  AND3_X1   g611(.A1(new_n513), .A2(new_n514), .A3(new_n490), .ZN(new_n813));
  AOI21_X1  g612(.A(new_n489), .B1(new_n513), .B2(new_n520), .ZN(new_n814));
  OAI21_X1  g613(.A(new_n532), .B1(new_n813), .B2(new_n814), .ZN(new_n815));
  NAND2_X1  g614(.A1(new_n536), .A2(new_n815), .ZN(new_n816));
  INV_X1    g615(.A(new_n816), .ZN(new_n817));
  NAND2_X1  g616(.A1(new_n661), .A2(new_n817), .ZN(new_n818));
  INV_X1    g617(.A(new_n818), .ZN(new_n819));
  OAI21_X1  g618(.A(new_n585), .B1(new_n812), .B2(new_n819), .ZN(new_n820));
  NAND2_X1  g619(.A1(new_n809), .A2(new_n811), .ZN(new_n821));
  NOR2_X1   g620(.A1(new_n585), .A2(new_n816), .ZN(new_n822));
  NAND4_X1  g621(.A1(new_n821), .A2(new_n660), .A3(new_n802), .A4(new_n822), .ZN(new_n823));
  NAND2_X1  g622(.A1(new_n820), .A2(new_n823), .ZN(new_n824));
  INV_X1    g623(.A(new_n686), .ZN(new_n825));
  AOI21_X1  g624(.A(new_n791), .B1(new_n824), .B2(new_n825), .ZN(new_n826));
  NOR2_X1   g625(.A1(new_n826), .A2(new_n741), .ZN(new_n827));
  NOR3_X1   g626(.A1(new_n667), .A2(new_n433), .A3(new_n302), .ZN(new_n828));
  NAND2_X1  g627(.A1(new_n827), .A2(new_n828), .ZN(new_n829));
  NOR3_X1   g628(.A1(new_n829), .A2(new_n246), .A3(new_n538), .ZN(new_n830));
  NOR2_X1   g629(.A1(new_n826), .A2(new_n433), .ZN(new_n831));
  INV_X1    g630(.A(new_n481), .ZN(new_n832));
  NAND2_X1  g631(.A1(new_n831), .A2(new_n832), .ZN(new_n833));
  NOR2_X1   g632(.A1(new_n833), .A2(new_n667), .ZN(new_n834));
  NAND2_X1  g633(.A1(new_n834), .A2(new_n537), .ZN(new_n835));
  AOI21_X1  g634(.A(new_n830), .B1(new_n835), .B2(new_n246), .ZN(G1340gat));
  NAND3_X1  g635(.A1(new_n834), .A2(new_n247), .A3(new_n661), .ZN(new_n837));
  OAI21_X1  g636(.A(G120gat), .B1(new_n829), .B2(new_n721), .ZN(new_n838));
  NAND2_X1  g637(.A1(new_n837), .A2(new_n838), .ZN(new_n839));
  XNOR2_X1  g638(.A(new_n839), .B(KEYINPUT110), .ZN(G1341gat));
  NAND3_X1  g639(.A1(new_n834), .A2(new_n254), .A3(new_n686), .ZN(new_n841));
  OAI21_X1  g640(.A(G127gat), .B1(new_n829), .B2(new_n825), .ZN(new_n842));
  NAND2_X1  g641(.A1(new_n841), .A2(new_n842), .ZN(G1342gat));
  NOR3_X1   g642(.A1(new_n667), .A2(G134gat), .A3(new_n585), .ZN(new_n844));
  NAND3_X1  g643(.A1(new_n831), .A2(new_n832), .A3(new_n844), .ZN(new_n845));
  INV_X1    g644(.A(KEYINPUT56), .ZN(new_n846));
  XNOR2_X1  g645(.A(new_n845), .B(new_n846), .ZN(new_n847));
  INV_X1    g646(.A(KEYINPUT111), .ZN(new_n848));
  NAND3_X1  g647(.A1(new_n827), .A2(new_n586), .A3(new_n828), .ZN(new_n849));
  AOI21_X1  g648(.A(new_n848), .B1(new_n849), .B2(G134gat), .ZN(new_n850));
  NAND3_X1  g649(.A1(new_n849), .A2(new_n848), .A3(G134gat), .ZN(new_n851));
  INV_X1    g650(.A(new_n851), .ZN(new_n852));
  OAI21_X1  g651(.A(new_n847), .B1(new_n850), .B2(new_n852), .ZN(new_n853));
  NAND2_X1  g652(.A1(new_n853), .A2(KEYINPUT112), .ZN(new_n854));
  INV_X1    g653(.A(KEYINPUT112), .ZN(new_n855));
  OAI211_X1 g654(.A(new_n847), .B(new_n855), .C1(new_n850), .C2(new_n852), .ZN(new_n856));
  NAND2_X1  g655(.A1(new_n854), .A2(new_n856), .ZN(G1343gat));
  NOR2_X1   g656(.A1(new_n667), .A2(new_n433), .ZN(new_n858));
  NAND2_X1  g657(.A1(new_n858), .A2(new_n676), .ZN(new_n859));
  INV_X1    g658(.A(KEYINPUT57), .ZN(new_n860));
  NOR2_X1   g659(.A1(new_n377), .A2(new_n860), .ZN(new_n861));
  OAI21_X1  g660(.A(new_n818), .B1(new_n803), .B2(new_n810), .ZN(new_n862));
  NAND2_X1  g661(.A1(new_n862), .A2(new_n585), .ZN(new_n863));
  AOI21_X1  g662(.A(new_n686), .B1(new_n823), .B2(new_n863), .ZN(new_n864));
  OAI21_X1  g663(.A(new_n861), .B1(new_n864), .B2(new_n791), .ZN(new_n865));
  INV_X1    g664(.A(new_n865), .ZN(new_n866));
  NAND2_X1  g665(.A1(new_n798), .A2(new_n801), .ZN(new_n867));
  AOI21_X1  g666(.A(KEYINPUT109), .B1(new_n867), .B2(new_n804), .ZN(new_n868));
  AOI211_X1 g667(.A(new_n808), .B(KEYINPUT55), .C1(new_n798), .C2(new_n801), .ZN(new_n869));
  NOR2_X1   g668(.A1(new_n868), .A2(new_n869), .ZN(new_n870));
  NAND4_X1  g669(.A1(new_n586), .A2(new_n802), .A3(new_n660), .A4(new_n817), .ZN(new_n871));
  NOR2_X1   g670(.A1(new_n870), .A2(new_n871), .ZN(new_n872));
  OAI21_X1  g671(.A(new_n818), .B1(new_n870), .B2(new_n803), .ZN(new_n873));
  AOI21_X1  g672(.A(new_n872), .B1(new_n873), .B2(new_n585), .ZN(new_n874));
  OAI21_X1  g673(.A(new_n790), .B1(new_n874), .B2(new_n686), .ZN(new_n875));
  AOI21_X1  g674(.A(KEYINPUT57), .B1(new_n875), .B2(new_n741), .ZN(new_n876));
  INV_X1    g675(.A(KEYINPUT113), .ZN(new_n877));
  AOI21_X1  g676(.A(new_n866), .B1(new_n876), .B2(new_n877), .ZN(new_n878));
  NOR2_X1   g677(.A1(new_n826), .A2(new_n377), .ZN(new_n879));
  OAI21_X1  g678(.A(KEYINPUT113), .B1(new_n879), .B2(KEYINPUT57), .ZN(new_n880));
  AOI21_X1  g679(.A(new_n859), .B1(new_n878), .B2(new_n880), .ZN(new_n881));
  AOI21_X1  g680(.A(new_n313), .B1(new_n881), .B2(new_n537), .ZN(new_n882));
  NOR2_X1   g681(.A1(new_n311), .A2(new_n377), .ZN(new_n883));
  AOI21_X1  g682(.A(new_n686), .B1(new_n820), .B2(new_n823), .ZN(new_n884));
  OAI211_X1 g683(.A(new_n483), .B(new_n883), .C1(new_n884), .C2(new_n791), .ZN(new_n885));
  NOR4_X1   g684(.A1(new_n885), .A2(G141gat), .A3(new_n667), .A4(new_n538), .ZN(new_n886));
  XNOR2_X1  g685(.A(new_n886), .B(KEYINPUT114), .ZN(new_n887));
  OAI21_X1  g686(.A(KEYINPUT58), .B1(new_n882), .B2(new_n887), .ZN(new_n888));
  INV_X1    g687(.A(KEYINPUT115), .ZN(new_n889));
  NAND2_X1  g688(.A1(new_n885), .A2(new_n889), .ZN(new_n890));
  NAND4_X1  g689(.A1(new_n875), .A2(KEYINPUT115), .A3(new_n483), .A4(new_n883), .ZN(new_n891));
  NOR2_X1   g690(.A1(new_n538), .A2(G141gat), .ZN(new_n892));
  NAND4_X1  g691(.A1(new_n890), .A2(new_n703), .A3(new_n891), .A4(new_n892), .ZN(new_n893));
  XOR2_X1   g692(.A(KEYINPUT116), .B(KEYINPUT58), .Z(new_n894));
  NAND2_X1  g693(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  INV_X1    g694(.A(new_n859), .ZN(new_n896));
  OAI211_X1 g695(.A(new_n877), .B(new_n860), .C1(new_n826), .C2(new_n377), .ZN(new_n897));
  NAND2_X1  g696(.A1(new_n897), .A2(new_n865), .ZN(new_n898));
  NAND2_X1  g697(.A1(new_n875), .A2(new_n741), .ZN(new_n899));
  AOI21_X1  g698(.A(new_n877), .B1(new_n899), .B2(new_n860), .ZN(new_n900));
  OAI211_X1 g699(.A(new_n537), .B(new_n896), .C1(new_n898), .C2(new_n900), .ZN(new_n901));
  AOI211_X1 g700(.A(KEYINPUT117), .B(new_n895), .C1(G141gat), .C2(new_n901), .ZN(new_n902));
  INV_X1    g701(.A(KEYINPUT117), .ZN(new_n903));
  NAND2_X1  g702(.A1(new_n901), .A2(G141gat), .ZN(new_n904));
  INV_X1    g703(.A(new_n895), .ZN(new_n905));
  AOI21_X1  g704(.A(new_n903), .B1(new_n904), .B2(new_n905), .ZN(new_n906));
  OAI21_X1  g705(.A(new_n888), .B1(new_n902), .B2(new_n906), .ZN(G1344gat));
  AOI211_X1 g706(.A(KEYINPUT59), .B(new_n315), .C1(new_n881), .C2(new_n661), .ZN(new_n908));
  INV_X1    g707(.A(KEYINPUT59), .ZN(new_n909));
  AOI21_X1  g708(.A(new_n721), .B1(new_n896), .B2(KEYINPUT118), .ZN(new_n910));
  OAI21_X1  g709(.A(new_n910), .B1(KEYINPUT118), .B2(new_n896), .ZN(new_n911));
  OAI21_X1  g710(.A(new_n741), .B1(new_n864), .B2(new_n791), .ZN(new_n912));
  NAND2_X1  g711(.A1(new_n912), .A2(new_n860), .ZN(new_n913));
  NAND2_X1  g712(.A1(new_n875), .A2(new_n861), .ZN(new_n914));
  AOI21_X1  g713(.A(new_n911), .B1(new_n913), .B2(new_n914), .ZN(new_n915));
  OR2_X1    g714(.A1(new_n915), .A2(KEYINPUT119), .ZN(new_n916));
  AOI21_X1  g715(.A(new_n315), .B1(new_n915), .B2(KEYINPUT119), .ZN(new_n917));
  AOI21_X1  g716(.A(new_n909), .B1(new_n916), .B2(new_n917), .ZN(new_n918));
  AND2_X1   g717(.A1(new_n890), .A2(new_n891), .ZN(new_n919));
  NAND2_X1  g718(.A1(new_n919), .A2(new_n703), .ZN(new_n920));
  NAND2_X1  g719(.A1(new_n661), .A2(new_n315), .ZN(new_n921));
  OAI22_X1  g720(.A1(new_n908), .A2(new_n918), .B1(new_n920), .B2(new_n921), .ZN(G1345gat));
  NAND2_X1  g721(.A1(new_n881), .A2(new_n686), .ZN(new_n923));
  NAND2_X1  g722(.A1(new_n923), .A2(G155gat), .ZN(new_n924));
  OR2_X1    g723(.A1(new_n825), .A2(G155gat), .ZN(new_n925));
  OAI21_X1  g724(.A(new_n924), .B1(new_n920), .B2(new_n925), .ZN(G1346gat));
  NAND2_X1  g725(.A1(new_n881), .A2(new_n586), .ZN(new_n927));
  INV_X1    g726(.A(KEYINPUT120), .ZN(new_n928));
  NAND2_X1  g727(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  NAND3_X1  g728(.A1(new_n881), .A2(KEYINPUT120), .A3(new_n586), .ZN(new_n930));
  NAND3_X1  g729(.A1(new_n929), .A2(G162gat), .A3(new_n930), .ZN(new_n931));
  NOR3_X1   g730(.A1(new_n667), .A2(G162gat), .A3(new_n585), .ZN(new_n932));
  NAND2_X1  g731(.A1(new_n919), .A2(new_n932), .ZN(new_n933));
  NAND2_X1  g732(.A1(new_n931), .A2(new_n933), .ZN(G1347gat));
  NAND3_X1  g733(.A1(new_n667), .A2(new_n433), .A3(new_n303), .ZN(new_n935));
  INV_X1    g734(.A(new_n935), .ZN(new_n936));
  NAND2_X1  g735(.A1(new_n827), .A2(new_n936), .ZN(new_n937));
  INV_X1    g736(.A(G169gat), .ZN(new_n938));
  NOR3_X1   g737(.A1(new_n937), .A2(new_n938), .A3(new_n538), .ZN(new_n939));
  NAND2_X1  g738(.A1(new_n667), .A2(new_n433), .ZN(new_n940));
  NOR3_X1   g739(.A1(new_n826), .A2(new_n481), .A3(new_n940), .ZN(new_n941));
  AOI21_X1  g740(.A(G169gat), .B1(new_n941), .B2(new_n537), .ZN(new_n942));
  NOR2_X1   g741(.A1(new_n939), .A2(new_n942), .ZN(G1348gat));
  OAI21_X1  g742(.A(G176gat), .B1(new_n937), .B2(new_n721), .ZN(new_n944));
  INV_X1    g743(.A(new_n941), .ZN(new_n945));
  OR2_X1    g744(.A1(new_n721), .A2(G176gat), .ZN(new_n946));
  OAI21_X1  g745(.A(new_n944), .B1(new_n945), .B2(new_n946), .ZN(G1349gat));
  INV_X1    g746(.A(KEYINPUT60), .ZN(new_n948));
  AND2_X1   g747(.A1(new_n686), .A2(new_n214), .ZN(new_n949));
  NAND2_X1  g748(.A1(new_n941), .A2(new_n949), .ZN(new_n950));
  NAND4_X1  g749(.A1(new_n875), .A2(new_n377), .A3(new_n686), .A4(new_n936), .ZN(new_n951));
  NAND2_X1  g750(.A1(new_n951), .A2(G183gat), .ZN(new_n952));
  NAND2_X1  g751(.A1(new_n950), .A2(new_n952), .ZN(new_n953));
  AOI21_X1  g752(.A(new_n948), .B1(new_n953), .B2(KEYINPUT121), .ZN(new_n954));
  INV_X1    g753(.A(KEYINPUT122), .ZN(new_n955));
  INV_X1    g754(.A(KEYINPUT121), .ZN(new_n956));
  NAND3_X1  g755(.A1(new_n950), .A2(new_n956), .A3(new_n952), .ZN(new_n957));
  AND3_X1   g756(.A1(new_n954), .A2(new_n955), .A3(new_n957), .ZN(new_n958));
  AOI21_X1  g757(.A(new_n955), .B1(new_n954), .B2(new_n957), .ZN(new_n959));
  XNOR2_X1  g758(.A(KEYINPUT123), .B(KEYINPUT60), .ZN(new_n960));
  OAI22_X1  g759(.A1(new_n958), .A2(new_n959), .B1(new_n953), .B2(new_n960), .ZN(G1350gat));
  OAI21_X1  g760(.A(G190gat), .B1(new_n937), .B2(new_n585), .ZN(new_n962));
  XNOR2_X1  g761(.A(new_n962), .B(KEYINPUT61), .ZN(new_n963));
  NAND3_X1  g762(.A1(new_n941), .A2(new_n209), .A3(new_n586), .ZN(new_n964));
  NAND2_X1  g763(.A1(new_n963), .A2(new_n964), .ZN(G1351gat));
  NOR2_X1   g764(.A1(new_n940), .A2(new_n311), .ZN(new_n966));
  NAND2_X1  g765(.A1(new_n879), .A2(new_n966), .ZN(new_n967));
  NOR3_X1   g766(.A1(new_n967), .A2(G197gat), .A3(new_n538), .ZN(new_n968));
  XOR2_X1   g767(.A(new_n966), .B(KEYINPUT124), .Z(new_n969));
  AOI21_X1  g768(.A(new_n969), .B1(new_n913), .B2(new_n914), .ZN(new_n970));
  NAND2_X1  g769(.A1(new_n970), .A2(new_n537), .ZN(new_n971));
  AOI21_X1  g770(.A(new_n968), .B1(new_n971), .B2(G197gat), .ZN(new_n972));
  XNOR2_X1  g771(.A(new_n972), .B(KEYINPUT125), .ZN(G1352gat));
  INV_X1    g772(.A(new_n967), .ZN(new_n974));
  AOI21_X1  g773(.A(G204gat), .B1(KEYINPUT126), .B2(KEYINPUT62), .ZN(new_n975));
  NAND3_X1  g774(.A1(new_n974), .A2(new_n661), .A3(new_n975), .ZN(new_n976));
  NOR2_X1   g775(.A1(KEYINPUT126), .A2(KEYINPUT62), .ZN(new_n977));
  XNOR2_X1  g776(.A(new_n976), .B(new_n977), .ZN(new_n978));
  NAND2_X1  g777(.A1(new_n970), .A2(new_n661), .ZN(new_n979));
  NAND2_X1  g778(.A1(new_n979), .A2(G204gat), .ZN(new_n980));
  NAND2_X1  g779(.A1(new_n978), .A2(new_n980), .ZN(G1353gat));
  NAND3_X1  g780(.A1(new_n974), .A2(new_n341), .A3(new_n686), .ZN(new_n982));
  NAND2_X1  g781(.A1(new_n970), .A2(new_n686), .ZN(new_n983));
  AND3_X1   g782(.A1(new_n983), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n984));
  AOI21_X1  g783(.A(KEYINPUT63), .B1(new_n983), .B2(G211gat), .ZN(new_n985));
  OAI21_X1  g784(.A(new_n982), .B1(new_n984), .B2(new_n985), .ZN(G1354gat));
  AOI21_X1  g785(.A(G218gat), .B1(new_n974), .B2(new_n586), .ZN(new_n987));
  NOR2_X1   g786(.A1(new_n585), .A2(new_n340), .ZN(new_n988));
  XOR2_X1   g787(.A(new_n988), .B(KEYINPUT127), .Z(new_n989));
  AOI21_X1  g788(.A(new_n987), .B1(new_n970), .B2(new_n989), .ZN(G1355gat));
endmodule


