//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 0 0 1 1 0 0 0 0 1 0 1 1 1 0 1 0 0 0 1 1 0 1 1 0 0 0 0 1 0 0 0 0 0 1 0 0 1 0 0 1 1 0 0 0 1 1 1 0 0 1 0 1 0 1 1 0 0 1 0 0 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:31:26 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n447, new_n451, new_n452, new_n453, new_n454, new_n455,
    new_n458, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n483, new_n484, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n532,
    new_n533, new_n534, new_n535, new_n536, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n545, new_n546, new_n547, new_n548, new_n549,
    new_n550, new_n552, new_n554, new_n555, new_n556, new_n558, new_n559,
    new_n560, new_n561, new_n562, new_n563, new_n564, new_n565, new_n566,
    new_n567, new_n568, new_n569, new_n570, new_n571, new_n572, new_n573,
    new_n574, new_n575, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n585, new_n586, new_n587, new_n588, new_n589, new_n590, new_n591,
    new_n592, new_n594, new_n595, new_n596, new_n597, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n609,
    new_n610, new_n613, new_n615, new_n616, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n824,
    new_n825, new_n826, new_n827, new_n828, new_n829, new_n830, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n895, new_n896, new_n897, new_n898,
    new_n899, new_n900, new_n901, new_n902, new_n903, new_n904, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1110, new_n1111, new_n1112,
    new_n1113;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  XOR2_X1   g004(.A(KEYINPUT64), .B(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XOR2_X1   g010(.A(KEYINPUT0), .B(G82), .Z(new_n436));
  INV_X1    g011(.A(new_n436), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  INV_X1    g015(.A(G57), .ZN(G237));
  INV_X1    g016(.A(G108), .ZN(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NAND4_X1  g025(.A1(new_n436), .A2(G44), .A3(G96), .A4(G132), .ZN(new_n451));
  XOR2_X1   g026(.A(new_n451), .B(KEYINPUT2), .Z(new_n452));
  INV_X1    g027(.A(new_n452), .ZN(new_n453));
  NOR4_X1   g028(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(new_n455));
  NOR2_X1   g030(.A1(new_n453), .A2(new_n455), .ZN(G325));
  INV_X1    g031(.A(G325), .ZN(G261));
  AOI22_X1  g032(.A1(new_n453), .A2(G2106), .B1(G567), .B2(new_n455), .ZN(new_n458));
  XOR2_X1   g033(.A(new_n458), .B(KEYINPUT65), .Z(G319));
  INV_X1    g034(.A(KEYINPUT3), .ZN(new_n460));
  NOR3_X1   g035(.A1(new_n460), .A2(KEYINPUT66), .A3(G2104), .ZN(new_n461));
  INV_X1    g036(.A(G2104), .ZN(new_n462));
  NAND2_X1  g037(.A1(new_n462), .A2(KEYINPUT3), .ZN(new_n463));
  INV_X1    g038(.A(KEYINPUT66), .ZN(new_n464));
  OAI21_X1  g039(.A(new_n464), .B1(new_n462), .B2(KEYINPUT3), .ZN(new_n465));
  AOI21_X1  g040(.A(new_n461), .B1(new_n463), .B2(new_n465), .ZN(new_n466));
  INV_X1    g041(.A(G2105), .ZN(new_n467));
  NAND4_X1  g042(.A1(new_n466), .A2(KEYINPUT67), .A3(G137), .A4(new_n467), .ZN(new_n468));
  INV_X1    g043(.A(KEYINPUT67), .ZN(new_n469));
  NAND3_X1  g044(.A1(new_n464), .A2(new_n462), .A3(KEYINPUT3), .ZN(new_n470));
  AOI21_X1  g045(.A(KEYINPUT66), .B1(new_n460), .B2(G2104), .ZN(new_n471));
  NOR2_X1   g046(.A1(new_n460), .A2(G2104), .ZN(new_n472));
  OAI211_X1 g047(.A(new_n467), .B(new_n470), .C1(new_n471), .C2(new_n472), .ZN(new_n473));
  INV_X1    g048(.A(G137), .ZN(new_n474));
  OAI21_X1  g049(.A(new_n469), .B1(new_n473), .B2(new_n474), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n468), .A2(new_n475), .ZN(new_n476));
  NAND2_X1  g051(.A1(G113), .A2(G2104), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n460), .A2(G2104), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n463), .A2(new_n478), .ZN(new_n479));
  INV_X1    g054(.A(G125), .ZN(new_n480));
  OAI21_X1  g055(.A(new_n477), .B1(new_n479), .B2(new_n480), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n481), .A2(G2105), .ZN(new_n482));
  NOR2_X1   g057(.A1(new_n462), .A2(G2105), .ZN(new_n483));
  NAND2_X1  g058(.A1(new_n483), .A2(G101), .ZN(new_n484));
  AND3_X1   g059(.A1(new_n476), .A2(new_n482), .A3(new_n484), .ZN(G160));
  INV_X1    g060(.A(KEYINPUT68), .ZN(new_n486));
  OR3_X1    g061(.A1(new_n486), .A2(G100), .A3(G2105), .ZN(new_n487));
  OAI21_X1  g062(.A(new_n486), .B1(G100), .B2(G2105), .ZN(new_n488));
  NAND3_X1  g063(.A1(new_n487), .A2(new_n488), .A3(G2104), .ZN(new_n489));
  NOR2_X1   g064(.A1(new_n467), .A2(G112), .ZN(new_n490));
  INV_X1    g065(.A(G136), .ZN(new_n491));
  OAI22_X1  g066(.A1(new_n489), .A2(new_n490), .B1(new_n473), .B2(new_n491), .ZN(new_n492));
  OAI211_X1 g067(.A(G2105), .B(new_n470), .C1(new_n471), .C2(new_n472), .ZN(new_n493));
  INV_X1    g068(.A(new_n493), .ZN(new_n494));
  AOI21_X1  g069(.A(new_n492), .B1(G124), .B2(new_n494), .ZN(G162));
  NAND4_X1  g070(.A1(new_n466), .A2(KEYINPUT69), .A3(G126), .A4(G2105), .ZN(new_n496));
  INV_X1    g071(.A(KEYINPUT69), .ZN(new_n497));
  INV_X1    g072(.A(G126), .ZN(new_n498));
  OAI21_X1  g073(.A(new_n497), .B1(new_n493), .B2(new_n498), .ZN(new_n499));
  NAND4_X1  g074(.A1(new_n463), .A2(new_n478), .A3(G138), .A4(new_n467), .ZN(new_n500));
  INV_X1    g075(.A(KEYINPUT4), .ZN(new_n501));
  OR2_X1    g076(.A1(G102), .A2(G2105), .ZN(new_n502));
  INV_X1    g077(.A(G114), .ZN(new_n503));
  AOI21_X1  g078(.A(new_n462), .B1(new_n503), .B2(G2105), .ZN(new_n504));
  AOI22_X1  g079(.A1(new_n500), .A2(new_n501), .B1(new_n502), .B2(new_n504), .ZN(new_n505));
  AND3_X1   g080(.A1(new_n467), .A2(KEYINPUT4), .A3(G138), .ZN(new_n506));
  NAND2_X1  g081(.A1(new_n466), .A2(new_n506), .ZN(new_n507));
  NAND4_X1  g082(.A1(new_n496), .A2(new_n499), .A3(new_n505), .A4(new_n507), .ZN(new_n508));
  INV_X1    g083(.A(new_n508), .ZN(G164));
  INV_X1    g084(.A(KEYINPUT71), .ZN(new_n510));
  OAI21_X1  g085(.A(G543), .B1(new_n510), .B2(KEYINPUT5), .ZN(new_n511));
  INV_X1    g086(.A(KEYINPUT70), .ZN(new_n512));
  NAND2_X1  g087(.A1(new_n512), .A2(KEYINPUT5), .ZN(new_n513));
  NAND2_X1  g088(.A1(new_n511), .A2(new_n513), .ZN(new_n514));
  NAND4_X1  g089(.A1(new_n512), .A2(new_n510), .A3(KEYINPUT5), .A4(G543), .ZN(new_n515));
  NAND2_X1  g090(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  AOI22_X1  g091(.A1(new_n516), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n517));
  INV_X1    g092(.A(G651), .ZN(new_n518));
  NOR2_X1   g093(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  NAND2_X1  g094(.A1(new_n518), .A2(KEYINPUT6), .ZN(new_n520));
  INV_X1    g095(.A(KEYINPUT6), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n521), .A2(G651), .ZN(new_n522));
  NAND2_X1  g097(.A1(new_n520), .A2(new_n522), .ZN(new_n523));
  INV_X1    g098(.A(G543), .ZN(new_n524));
  NOR2_X1   g099(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  NAND2_X1  g100(.A1(new_n525), .A2(G50), .ZN(new_n526));
  AOI21_X1  g101(.A(new_n523), .B1(new_n514), .B2(new_n515), .ZN(new_n527));
  INV_X1    g102(.A(new_n527), .ZN(new_n528));
  INV_X1    g103(.A(G88), .ZN(new_n529));
  OAI21_X1  g104(.A(new_n526), .B1(new_n528), .B2(new_n529), .ZN(new_n530));
  NOR2_X1   g105(.A1(new_n519), .A2(new_n530), .ZN(G166));
  NAND2_X1  g106(.A1(new_n527), .A2(G89), .ZN(new_n532));
  NAND3_X1  g107(.A1(new_n516), .A2(G63), .A3(G651), .ZN(new_n533));
  NAND3_X1  g108(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n534));
  XNOR2_X1  g109(.A(new_n534), .B(KEYINPUT7), .ZN(new_n535));
  NAND2_X1  g110(.A1(new_n525), .A2(G51), .ZN(new_n536));
  NAND4_X1  g111(.A1(new_n532), .A2(new_n533), .A3(new_n535), .A4(new_n536), .ZN(G286));
  INV_X1    g112(.A(G286), .ZN(G168));
  AOI22_X1  g113(.A1(new_n516), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n539));
  NOR2_X1   g114(.A1(new_n539), .A2(new_n518), .ZN(new_n540));
  NAND2_X1  g115(.A1(new_n525), .A2(G52), .ZN(new_n541));
  INV_X1    g116(.A(G90), .ZN(new_n542));
  OAI21_X1  g117(.A(new_n541), .B1(new_n528), .B2(new_n542), .ZN(new_n543));
  NOR2_X1   g118(.A1(new_n540), .A2(new_n543), .ZN(G171));
  AOI22_X1  g119(.A1(new_n516), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n545));
  NOR2_X1   g120(.A1(new_n545), .A2(new_n518), .ZN(new_n546));
  XNOR2_X1  g121(.A(new_n546), .B(KEYINPUT72), .ZN(new_n547));
  NAND2_X1  g122(.A1(new_n527), .A2(G81), .ZN(new_n548));
  NAND2_X1  g123(.A1(new_n525), .A2(G43), .ZN(new_n549));
  AND3_X1   g124(.A1(new_n547), .A2(new_n548), .A3(new_n549), .ZN(new_n550));
  NAND2_X1  g125(.A1(new_n550), .A2(G860), .ZN(G153));
  AND3_X1   g126(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n552));
  NAND2_X1  g127(.A1(new_n552), .A2(G36), .ZN(G176));
  XOR2_X1   g128(.A(KEYINPUT73), .B(KEYINPUT8), .Z(new_n554));
  NAND2_X1  g129(.A1(G1), .A2(G3), .ZN(new_n555));
  XNOR2_X1  g130(.A(new_n554), .B(new_n555), .ZN(new_n556));
  NAND2_X1  g131(.A1(new_n552), .A2(new_n556), .ZN(G188));
  NAND2_X1  g132(.A1(new_n525), .A2(G53), .ZN(new_n558));
  NAND2_X1  g133(.A1(KEYINPUT74), .A2(KEYINPUT9), .ZN(new_n559));
  XOR2_X1   g134(.A(new_n558), .B(new_n559), .Z(new_n560));
  INV_X1    g135(.A(KEYINPUT76), .ZN(new_n561));
  XNOR2_X1  g136(.A(KEYINPUT75), .B(G65), .ZN(new_n562));
  AOI21_X1  g137(.A(new_n562), .B1(new_n514), .B2(new_n515), .ZN(new_n563));
  NAND2_X1  g138(.A1(G78), .A2(G543), .ZN(new_n564));
  INV_X1    g139(.A(new_n564), .ZN(new_n565));
  OAI21_X1  g140(.A(new_n561), .B1(new_n563), .B2(new_n565), .ZN(new_n566));
  INV_X1    g141(.A(new_n562), .ZN(new_n567));
  INV_X1    g142(.A(KEYINPUT5), .ZN(new_n568));
  NAND2_X1  g143(.A1(new_n568), .A2(KEYINPUT71), .ZN(new_n569));
  AOI22_X1  g144(.A1(new_n569), .A2(G543), .B1(new_n512), .B2(KEYINPUT5), .ZN(new_n570));
  INV_X1    g145(.A(new_n515), .ZN(new_n571));
  OAI21_X1  g146(.A(new_n567), .B1(new_n570), .B2(new_n571), .ZN(new_n572));
  NAND3_X1  g147(.A1(new_n572), .A2(KEYINPUT76), .A3(new_n564), .ZN(new_n573));
  NAND3_X1  g148(.A1(new_n566), .A2(new_n573), .A3(G651), .ZN(new_n574));
  NAND2_X1  g149(.A1(new_n527), .A2(G91), .ZN(new_n575));
  NAND3_X1  g150(.A1(new_n560), .A2(new_n574), .A3(new_n575), .ZN(G299));
  INV_X1    g151(.A(G171), .ZN(G301));
  INV_X1    g152(.A(G166), .ZN(G303));
  NAND2_X1  g153(.A1(new_n527), .A2(G87), .ZN(new_n579));
  XNOR2_X1  g154(.A(new_n579), .B(KEYINPUT77), .ZN(new_n580));
  OAI21_X1  g155(.A(G651), .B1(new_n516), .B2(G74), .ZN(new_n581));
  NAND2_X1  g156(.A1(new_n525), .A2(G49), .ZN(new_n582));
  XNOR2_X1  g157(.A(new_n582), .B(KEYINPUT78), .ZN(new_n583));
  NAND3_X1  g158(.A1(new_n580), .A2(new_n581), .A3(new_n583), .ZN(G288));
  NAND2_X1  g159(.A1(new_n525), .A2(G48), .ZN(new_n585));
  INV_X1    g160(.A(G86), .ZN(new_n586));
  OAI21_X1  g161(.A(new_n585), .B1(new_n528), .B2(new_n586), .ZN(new_n587));
  NAND2_X1  g162(.A1(new_n516), .A2(G61), .ZN(new_n588));
  NAND2_X1  g163(.A1(G73), .A2(G543), .ZN(new_n589));
  XOR2_X1   g164(.A(new_n589), .B(KEYINPUT79), .Z(new_n590));
  AOI21_X1  g165(.A(new_n518), .B1(new_n588), .B2(new_n590), .ZN(new_n591));
  NOR2_X1   g166(.A1(new_n587), .A2(new_n591), .ZN(new_n592));
  INV_X1    g167(.A(new_n592), .ZN(G305));
  AOI22_X1  g168(.A1(new_n516), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n594));
  XOR2_X1   g169(.A(new_n594), .B(KEYINPUT80), .Z(new_n595));
  NAND2_X1  g170(.A1(new_n595), .A2(G651), .ZN(new_n596));
  AOI22_X1  g171(.A1(new_n527), .A2(G85), .B1(G47), .B2(new_n525), .ZN(new_n597));
  NAND2_X1  g172(.A1(new_n596), .A2(new_n597), .ZN(G290));
  NAND2_X1  g173(.A1(G301), .A2(G868), .ZN(new_n599));
  NAND2_X1  g174(.A1(new_n527), .A2(G92), .ZN(new_n600));
  XOR2_X1   g175(.A(new_n600), .B(KEYINPUT10), .Z(new_n601));
  NAND2_X1  g176(.A1(new_n525), .A2(G54), .ZN(new_n602));
  AOI22_X1  g177(.A1(new_n516), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n603));
  OR2_X1    g178(.A1(new_n603), .A2(new_n518), .ZN(new_n604));
  NAND3_X1  g179(.A1(new_n601), .A2(new_n602), .A3(new_n604), .ZN(new_n605));
  INV_X1    g180(.A(new_n605), .ZN(new_n606));
  OAI21_X1  g181(.A(new_n599), .B1(new_n606), .B2(G868), .ZN(G284));
  OAI21_X1  g182(.A(new_n599), .B1(new_n606), .B2(G868), .ZN(G321));
  NAND2_X1  g183(.A1(G286), .A2(G868), .ZN(new_n609));
  INV_X1    g184(.A(G299), .ZN(new_n610));
  OAI21_X1  g185(.A(new_n609), .B1(new_n610), .B2(G868), .ZN(G297));
  OAI21_X1  g186(.A(new_n609), .B1(new_n610), .B2(G868), .ZN(G280));
  INV_X1    g187(.A(G559), .ZN(new_n613));
  OAI21_X1  g188(.A(new_n606), .B1(new_n613), .B2(G860), .ZN(G148));
  NAND2_X1  g189(.A1(new_n606), .A2(new_n613), .ZN(new_n615));
  NAND2_X1  g190(.A1(new_n615), .A2(G868), .ZN(new_n616));
  OAI21_X1  g191(.A(new_n616), .B1(G868), .B2(new_n550), .ZN(G323));
  XNOR2_X1  g192(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g193(.A1(new_n494), .A2(G123), .ZN(new_n619));
  INV_X1    g194(.A(G135), .ZN(new_n620));
  NOR2_X1   g195(.A1(G99), .A2(G2105), .ZN(new_n621));
  OAI21_X1  g196(.A(G2104), .B1(new_n467), .B2(G111), .ZN(new_n622));
  OAI221_X1 g197(.A(new_n619), .B1(new_n620), .B2(new_n473), .C1(new_n621), .C2(new_n622), .ZN(new_n623));
  XOR2_X1   g198(.A(new_n623), .B(G2096), .Z(new_n624));
  NAND3_X1  g199(.A1(new_n467), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n625));
  XNOR2_X1  g200(.A(new_n625), .B(KEYINPUT12), .ZN(new_n626));
  XNOR2_X1  g201(.A(new_n626), .B(KEYINPUT13), .ZN(new_n627));
  XNOR2_X1  g202(.A(new_n627), .B(G2100), .ZN(new_n628));
  NAND2_X1  g203(.A1(new_n624), .A2(new_n628), .ZN(G156));
  XNOR2_X1  g204(.A(KEYINPUT15), .B(G2430), .ZN(new_n630));
  XNOR2_X1  g205(.A(new_n630), .B(G2435), .ZN(new_n631));
  XOR2_X1   g206(.A(G2427), .B(G2438), .Z(new_n632));
  XNOR2_X1  g207(.A(new_n631), .B(new_n632), .ZN(new_n633));
  NAND2_X1  g208(.A1(new_n633), .A2(KEYINPUT14), .ZN(new_n634));
  XOR2_X1   g209(.A(G2443), .B(G2446), .Z(new_n635));
  XNOR2_X1  g210(.A(new_n634), .B(new_n635), .ZN(new_n636));
  XNOR2_X1  g211(.A(G1341), .B(G1348), .ZN(new_n637));
  XNOR2_X1  g212(.A(KEYINPUT81), .B(KEYINPUT16), .ZN(new_n638));
  XNOR2_X1  g213(.A(new_n637), .B(new_n638), .ZN(new_n639));
  XNOR2_X1  g214(.A(new_n636), .B(new_n639), .ZN(new_n640));
  XNOR2_X1  g215(.A(G2451), .B(G2454), .ZN(new_n641));
  XOR2_X1   g216(.A(new_n640), .B(new_n641), .Z(new_n642));
  AND2_X1   g217(.A1(new_n642), .A2(G14), .ZN(G401));
  XOR2_X1   g218(.A(G2067), .B(G2678), .Z(new_n644));
  INV_X1    g219(.A(new_n644), .ZN(new_n645));
  XOR2_X1   g220(.A(G2084), .B(G2090), .Z(new_n646));
  NAND2_X1  g221(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  AND2_X1   g222(.A1(new_n647), .A2(KEYINPUT17), .ZN(new_n648));
  OR2_X1    g223(.A1(new_n645), .A2(new_n646), .ZN(new_n649));
  AOI21_X1  g224(.A(KEYINPUT18), .B1(new_n648), .B2(new_n649), .ZN(new_n650));
  XNOR2_X1  g225(.A(G2072), .B(G2078), .ZN(new_n651));
  XNOR2_X1  g226(.A(new_n651), .B(KEYINPUT82), .ZN(new_n652));
  AOI21_X1  g227(.A(new_n652), .B1(KEYINPUT18), .B2(new_n647), .ZN(new_n653));
  XNOR2_X1  g228(.A(new_n650), .B(new_n653), .ZN(new_n654));
  XOR2_X1   g229(.A(G2096), .B(G2100), .Z(new_n655));
  XNOR2_X1  g230(.A(new_n654), .B(new_n655), .ZN(G227));
  XNOR2_X1  g231(.A(G1971), .B(G1976), .ZN(new_n657));
  XNOR2_X1  g232(.A(new_n657), .B(KEYINPUT83), .ZN(new_n658));
  XOR2_X1   g233(.A(new_n658), .B(KEYINPUT19), .Z(new_n659));
  XOR2_X1   g234(.A(G1956), .B(G2474), .Z(new_n660));
  XOR2_X1   g235(.A(G1961), .B(G1966), .Z(new_n661));
  NOR2_X1   g236(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  INV_X1    g237(.A(new_n662), .ZN(new_n663));
  NOR2_X1   g238(.A1(new_n659), .A2(new_n663), .ZN(new_n664));
  NAND2_X1  g239(.A1(new_n660), .A2(new_n661), .ZN(new_n665));
  XNOR2_X1  g240(.A(new_n665), .B(KEYINPUT84), .ZN(new_n666));
  NOR2_X1   g241(.A1(new_n659), .A2(new_n666), .ZN(new_n667));
  AOI21_X1  g242(.A(new_n664), .B1(KEYINPUT20), .B2(new_n667), .ZN(new_n668));
  NAND3_X1  g243(.A1(new_n659), .A2(new_n665), .A3(new_n663), .ZN(new_n669));
  OAI211_X1 g244(.A(new_n668), .B(new_n669), .C1(KEYINPUT20), .C2(new_n667), .ZN(new_n670));
  XOR2_X1   g245(.A(G1991), .B(G1996), .Z(new_n671));
  XNOR2_X1  g246(.A(new_n670), .B(new_n671), .ZN(new_n672));
  XOR2_X1   g247(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n673));
  XNOR2_X1  g248(.A(new_n672), .B(new_n673), .ZN(new_n674));
  XNOR2_X1  g249(.A(G1981), .B(G1986), .ZN(new_n675));
  XNOR2_X1  g250(.A(new_n675), .B(KEYINPUT85), .ZN(new_n676));
  XNOR2_X1  g251(.A(new_n674), .B(new_n676), .ZN(G229));
  INV_X1    g252(.A(KEYINPUT88), .ZN(new_n678));
  INV_X1    g253(.A(G16), .ZN(new_n679));
  NAND2_X1  g254(.A1(new_n679), .A2(G24), .ZN(new_n680));
  INV_X1    g255(.A(G290), .ZN(new_n681));
  OAI21_X1  g256(.A(new_n680), .B1(new_n681), .B2(new_n679), .ZN(new_n682));
  XNOR2_X1  g257(.A(new_n682), .B(G1986), .ZN(new_n683));
  NAND2_X1  g258(.A1(new_n679), .A2(G23), .ZN(new_n684));
  INV_X1    g259(.A(G288), .ZN(new_n685));
  OAI21_X1  g260(.A(new_n684), .B1(new_n685), .B2(new_n679), .ZN(new_n686));
  XOR2_X1   g261(.A(new_n686), .B(KEYINPUT33), .Z(new_n687));
  OR2_X1    g262(.A1(new_n687), .A2(G1976), .ZN(new_n688));
  NAND2_X1  g263(.A1(new_n687), .A2(G1976), .ZN(new_n689));
  NAND2_X1  g264(.A1(new_n679), .A2(G6), .ZN(new_n690));
  OAI21_X1  g265(.A(new_n690), .B1(new_n592), .B2(new_n679), .ZN(new_n691));
  XOR2_X1   g266(.A(KEYINPUT32), .B(G1981), .Z(new_n692));
  XNOR2_X1  g267(.A(new_n691), .B(new_n692), .ZN(new_n693));
  NAND2_X1  g268(.A1(new_n679), .A2(G22), .ZN(new_n694));
  OAI21_X1  g269(.A(new_n694), .B1(G166), .B2(new_n679), .ZN(new_n695));
  INV_X1    g270(.A(G1971), .ZN(new_n696));
  XNOR2_X1  g271(.A(new_n695), .B(new_n696), .ZN(new_n697));
  NAND4_X1  g272(.A1(new_n688), .A2(new_n689), .A3(new_n693), .A4(new_n697), .ZN(new_n698));
  AOI211_X1 g273(.A(new_n678), .B(new_n683), .C1(new_n698), .C2(KEYINPUT34), .ZN(new_n699));
  AND2_X1   g274(.A1(KEYINPUT86), .A2(G29), .ZN(new_n700));
  NOR2_X1   g275(.A1(KEYINPUT86), .A2(G29), .ZN(new_n701));
  NOR2_X1   g276(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  INV_X1    g277(.A(new_n702), .ZN(new_n703));
  NAND2_X1  g278(.A1(new_n703), .A2(G25), .ZN(new_n704));
  INV_X1    g279(.A(G131), .ZN(new_n705));
  NOR2_X1   g280(.A1(G95), .A2(G2105), .ZN(new_n706));
  OAI21_X1  g281(.A(G2104), .B1(new_n467), .B2(G107), .ZN(new_n707));
  OAI22_X1  g282(.A1(new_n473), .A2(new_n705), .B1(new_n706), .B2(new_n707), .ZN(new_n708));
  AOI21_X1  g283(.A(new_n708), .B1(G119), .B2(new_n494), .ZN(new_n709));
  OAI21_X1  g284(.A(new_n704), .B1(new_n709), .B2(new_n703), .ZN(new_n710));
  XNOR2_X1  g285(.A(KEYINPUT35), .B(G1991), .ZN(new_n711));
  XOR2_X1   g286(.A(new_n711), .B(KEYINPUT87), .Z(new_n712));
  XNOR2_X1  g287(.A(new_n710), .B(new_n712), .ZN(new_n713));
  OAI211_X1 g288(.A(new_n699), .B(new_n713), .C1(KEYINPUT34), .C2(new_n698), .ZN(new_n714));
  INV_X1    g289(.A(KEYINPUT36), .ZN(new_n715));
  OR2_X1    g290(.A1(new_n714), .A2(new_n715), .ZN(new_n716));
  AOI22_X1  g291(.A1(new_n494), .A2(G129), .B1(G105), .B2(new_n483), .ZN(new_n717));
  NAND3_X1  g292(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n718));
  XOR2_X1   g293(.A(new_n718), .B(KEYINPUT26), .Z(new_n719));
  INV_X1    g294(.A(G141), .ZN(new_n720));
  OAI211_X1 g295(.A(new_n717), .B(new_n719), .C1(new_n720), .C2(new_n473), .ZN(new_n721));
  INV_X1    g296(.A(KEYINPUT94), .ZN(new_n722));
  OR2_X1    g297(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  NAND2_X1  g298(.A1(new_n721), .A2(new_n722), .ZN(new_n724));
  NAND2_X1  g299(.A1(new_n723), .A2(new_n724), .ZN(new_n725));
  INV_X1    g300(.A(new_n725), .ZN(new_n726));
  NAND2_X1  g301(.A1(new_n726), .A2(G29), .ZN(new_n727));
  NOR2_X1   g302(.A1(G29), .A2(G32), .ZN(new_n728));
  OAI21_X1  g303(.A(new_n727), .B1(KEYINPUT95), .B2(new_n728), .ZN(new_n729));
  OAI21_X1  g304(.A(new_n729), .B1(KEYINPUT95), .B2(new_n727), .ZN(new_n730));
  XNOR2_X1  g305(.A(KEYINPUT27), .B(G1996), .ZN(new_n731));
  XNOR2_X1  g306(.A(new_n731), .B(KEYINPUT96), .ZN(new_n732));
  XNOR2_X1  g307(.A(new_n730), .B(new_n732), .ZN(new_n733));
  NAND2_X1  g308(.A1(new_n714), .A2(new_n715), .ZN(new_n734));
  NAND2_X1  g309(.A1(new_n703), .A2(G26), .ZN(new_n735));
  XOR2_X1   g310(.A(KEYINPUT89), .B(KEYINPUT28), .Z(new_n736));
  XNOR2_X1  g311(.A(new_n735), .B(new_n736), .ZN(new_n737));
  INV_X1    g312(.A(G140), .ZN(new_n738));
  NOR2_X1   g313(.A1(G104), .A2(G2105), .ZN(new_n739));
  OAI21_X1  g314(.A(G2104), .B1(new_n467), .B2(G116), .ZN(new_n740));
  OAI22_X1  g315(.A1(new_n473), .A2(new_n738), .B1(new_n739), .B2(new_n740), .ZN(new_n741));
  AOI21_X1  g316(.A(new_n741), .B1(G128), .B2(new_n494), .ZN(new_n742));
  INV_X1    g317(.A(G29), .ZN(new_n743));
  OAI21_X1  g318(.A(new_n737), .B1(new_n742), .B2(new_n743), .ZN(new_n744));
  XNOR2_X1  g319(.A(new_n744), .B(G2067), .ZN(new_n745));
  NAND2_X1  g320(.A1(new_n679), .A2(G4), .ZN(new_n746));
  OAI21_X1  g321(.A(new_n746), .B1(new_n606), .B2(new_n679), .ZN(new_n747));
  XNOR2_X1  g322(.A(new_n747), .B(G1348), .ZN(new_n748));
  INV_X1    g323(.A(G2084), .ZN(new_n749));
  NAND2_X1  g324(.A1(G160), .A2(G29), .ZN(new_n750));
  INV_X1    g325(.A(G34), .ZN(new_n751));
  AOI21_X1  g326(.A(new_n702), .B1(KEYINPUT24), .B2(new_n751), .ZN(new_n752));
  XOR2_X1   g327(.A(new_n752), .B(KEYINPUT92), .Z(new_n753));
  OAI21_X1  g328(.A(new_n753), .B1(KEYINPUT24), .B2(new_n751), .ZN(new_n754));
  NAND2_X1  g329(.A1(new_n750), .A2(new_n754), .ZN(new_n755));
  AOI211_X1 g330(.A(new_n745), .B(new_n748), .C1(new_n749), .C2(new_n755), .ZN(new_n756));
  NAND2_X1  g331(.A1(new_n679), .A2(G5), .ZN(new_n757));
  OAI21_X1  g332(.A(new_n757), .B1(G171), .B2(new_n679), .ZN(new_n758));
  INV_X1    g333(.A(G1961), .ZN(new_n759));
  XNOR2_X1  g334(.A(new_n758), .B(new_n759), .ZN(new_n760));
  NOR2_X1   g335(.A1(new_n755), .A2(new_n749), .ZN(new_n761));
  XOR2_X1   g336(.A(new_n761), .B(KEYINPUT93), .Z(new_n762));
  NAND2_X1  g337(.A1(new_n679), .A2(G21), .ZN(new_n763));
  OAI21_X1  g338(.A(new_n763), .B1(G168), .B2(new_n679), .ZN(new_n764));
  INV_X1    g339(.A(G1966), .ZN(new_n765));
  XNOR2_X1  g340(.A(new_n764), .B(new_n765), .ZN(new_n766));
  XOR2_X1   g341(.A(KEYINPUT97), .B(G28), .Z(new_n767));
  INV_X1    g342(.A(KEYINPUT30), .ZN(new_n768));
  NOR2_X1   g343(.A1(new_n767), .A2(new_n768), .ZN(new_n769));
  NAND2_X1  g344(.A1(new_n767), .A2(new_n768), .ZN(new_n770));
  AOI21_X1  g345(.A(G29), .B1(new_n770), .B2(KEYINPUT98), .ZN(new_n771));
  OAI21_X1  g346(.A(new_n771), .B1(KEYINPUT98), .B2(new_n770), .ZN(new_n772));
  OAI221_X1 g347(.A(new_n766), .B1(new_n623), .B2(new_n703), .C1(new_n769), .C2(new_n772), .ZN(new_n773));
  NAND2_X1  g348(.A1(new_n703), .A2(G27), .ZN(new_n774));
  OAI21_X1  g349(.A(new_n774), .B1(G164), .B2(new_n703), .ZN(new_n775));
  XNOR2_X1  g350(.A(new_n775), .B(G2078), .ZN(new_n776));
  XOR2_X1   g351(.A(KEYINPUT31), .B(G11), .Z(new_n777));
  NOR3_X1   g352(.A1(new_n773), .A2(new_n776), .A3(new_n777), .ZN(new_n778));
  NAND4_X1  g353(.A1(new_n756), .A2(new_n760), .A3(new_n762), .A4(new_n778), .ZN(new_n779));
  NAND2_X1  g354(.A1(new_n550), .A2(G16), .ZN(new_n780));
  OAI21_X1  g355(.A(new_n780), .B1(G16), .B2(G19), .ZN(new_n781));
  INV_X1    g356(.A(G1341), .ZN(new_n782));
  NAND2_X1  g357(.A1(new_n703), .A2(G35), .ZN(new_n783));
  OAI21_X1  g358(.A(new_n783), .B1(G162), .B2(new_n703), .ZN(new_n784));
  XNOR2_X1  g359(.A(new_n784), .B(KEYINPUT29), .ZN(new_n785));
  AOI22_X1  g360(.A1(new_n781), .A2(new_n782), .B1(G2090), .B2(new_n785), .ZN(new_n786));
  NAND2_X1  g361(.A1(new_n743), .A2(G33), .ZN(new_n787));
  NAND2_X1  g362(.A1(new_n483), .A2(G103), .ZN(new_n788));
  XOR2_X1   g363(.A(new_n788), .B(KEYINPUT25), .Z(new_n789));
  INV_X1    g364(.A(G139), .ZN(new_n790));
  AND2_X1   g365(.A1(new_n463), .A2(new_n478), .ZN(new_n791));
  AOI22_X1  g366(.A1(new_n791), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n792));
  OAI221_X1 g367(.A(new_n789), .B1(new_n790), .B2(new_n473), .C1(new_n792), .C2(new_n467), .ZN(new_n793));
  XNOR2_X1  g368(.A(new_n793), .B(KEYINPUT90), .ZN(new_n794));
  OAI21_X1  g369(.A(new_n787), .B1(new_n794), .B2(new_n743), .ZN(new_n795));
  XNOR2_X1  g370(.A(KEYINPUT91), .B(G2072), .ZN(new_n796));
  XNOR2_X1  g371(.A(new_n795), .B(new_n796), .ZN(new_n797));
  OAI211_X1 g372(.A(new_n786), .B(new_n797), .C1(G2090), .C2(new_n785), .ZN(new_n798));
  NOR2_X1   g373(.A1(new_n781), .A2(new_n782), .ZN(new_n799));
  NAND2_X1  g374(.A1(new_n679), .A2(G20), .ZN(new_n800));
  OAI211_X1 g375(.A(KEYINPUT23), .B(new_n800), .C1(new_n610), .C2(new_n679), .ZN(new_n801));
  OAI21_X1  g376(.A(new_n801), .B1(KEYINPUT23), .B2(new_n800), .ZN(new_n802));
  INV_X1    g377(.A(G1956), .ZN(new_n803));
  XNOR2_X1  g378(.A(new_n802), .B(new_n803), .ZN(new_n804));
  NOR4_X1   g379(.A1(new_n779), .A2(new_n798), .A3(new_n799), .A4(new_n804), .ZN(new_n805));
  NAND4_X1  g380(.A1(new_n716), .A2(new_n733), .A3(new_n734), .A4(new_n805), .ZN(G150));
  INV_X1    g381(.A(G150), .ZN(G311));
  AOI22_X1  g382(.A1(new_n516), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n808));
  NOR2_X1   g383(.A1(new_n808), .A2(new_n518), .ZN(new_n809));
  XOR2_X1   g384(.A(new_n809), .B(KEYINPUT99), .Z(new_n810));
  NAND2_X1  g385(.A1(new_n525), .A2(G55), .ZN(new_n811));
  INV_X1    g386(.A(G93), .ZN(new_n812));
  OAI211_X1 g387(.A(new_n810), .B(new_n811), .C1(new_n812), .C2(new_n528), .ZN(new_n813));
  NAND2_X1  g388(.A1(new_n813), .A2(G860), .ZN(new_n814));
  XOR2_X1   g389(.A(new_n814), .B(KEYINPUT37), .Z(new_n815));
  OR2_X1    g390(.A1(new_n813), .A2(new_n550), .ZN(new_n816));
  NAND2_X1  g391(.A1(new_n813), .A2(new_n550), .ZN(new_n817));
  NAND2_X1  g392(.A1(new_n816), .A2(new_n817), .ZN(new_n818));
  XNOR2_X1  g393(.A(new_n818), .B(KEYINPUT39), .ZN(new_n819));
  NAND2_X1  g394(.A1(new_n606), .A2(G559), .ZN(new_n820));
  XNOR2_X1  g395(.A(new_n820), .B(KEYINPUT38), .ZN(new_n821));
  XNOR2_X1  g396(.A(new_n819), .B(new_n821), .ZN(new_n822));
  OAI21_X1  g397(.A(new_n815), .B1(new_n822), .B2(G860), .ZN(G145));
  XNOR2_X1  g398(.A(new_n623), .B(G162), .ZN(new_n824));
  XNOR2_X1  g399(.A(new_n824), .B(G160), .ZN(new_n825));
  INV_X1    g400(.A(new_n742), .ZN(new_n826));
  XNOR2_X1  g401(.A(new_n725), .B(new_n826), .ZN(new_n827));
  XNOR2_X1  g402(.A(new_n827), .B(new_n508), .ZN(new_n828));
  NOR2_X1   g403(.A1(new_n794), .A2(KEYINPUT100), .ZN(new_n829));
  OR2_X1    g404(.A1(new_n828), .A2(new_n829), .ZN(new_n830));
  AND2_X1   g405(.A1(new_n794), .A2(KEYINPUT100), .ZN(new_n831));
  OAI21_X1  g406(.A(new_n828), .B1(new_n829), .B2(new_n831), .ZN(new_n832));
  NAND2_X1  g407(.A1(new_n830), .A2(new_n832), .ZN(new_n833));
  INV_X1    g408(.A(G142), .ZN(new_n834));
  NOR2_X1   g409(.A1(G106), .A2(G2105), .ZN(new_n835));
  OAI21_X1  g410(.A(G2104), .B1(new_n467), .B2(G118), .ZN(new_n836));
  OAI22_X1  g411(.A1(new_n473), .A2(new_n834), .B1(new_n835), .B2(new_n836), .ZN(new_n837));
  AOI21_X1  g412(.A(new_n837), .B1(G130), .B2(new_n494), .ZN(new_n838));
  XNOR2_X1  g413(.A(new_n709), .B(new_n838), .ZN(new_n839));
  XNOR2_X1  g414(.A(new_n839), .B(KEYINPUT101), .ZN(new_n840));
  XNOR2_X1  g415(.A(new_n840), .B(new_n626), .ZN(new_n841));
  NAND2_X1  g416(.A1(new_n833), .A2(new_n841), .ZN(new_n842));
  INV_X1    g417(.A(new_n841), .ZN(new_n843));
  NAND3_X1  g418(.A1(new_n830), .A2(new_n843), .A3(new_n832), .ZN(new_n844));
  AOI21_X1  g419(.A(new_n825), .B1(new_n842), .B2(new_n844), .ZN(new_n845));
  AND2_X1   g420(.A1(new_n845), .A2(KEYINPUT102), .ZN(new_n846));
  INV_X1    g421(.A(G37), .ZN(new_n847));
  OAI21_X1  g422(.A(new_n847), .B1(new_n845), .B2(KEYINPUT102), .ZN(new_n848));
  NOR2_X1   g423(.A1(new_n846), .A2(new_n848), .ZN(new_n849));
  NAND3_X1  g424(.A1(new_n842), .A2(new_n844), .A3(new_n825), .ZN(new_n850));
  NAND2_X1  g425(.A1(new_n849), .A2(new_n850), .ZN(new_n851));
  XNOR2_X1  g426(.A(new_n851), .B(KEYINPUT40), .ZN(G395));
  XOR2_X1   g427(.A(new_n818), .B(new_n615), .Z(new_n853));
  XNOR2_X1  g428(.A(new_n610), .B(new_n605), .ZN(new_n854));
  NAND2_X1  g429(.A1(new_n853), .A2(new_n854), .ZN(new_n855));
  XOR2_X1   g430(.A(new_n855), .B(KEYINPUT103), .Z(new_n856));
  XNOR2_X1  g431(.A(new_n854), .B(KEYINPUT41), .ZN(new_n857));
  OAI21_X1  g432(.A(new_n856), .B1(new_n857), .B2(new_n853), .ZN(new_n858));
  XNOR2_X1  g433(.A(G288), .B(G303), .ZN(new_n859));
  XNOR2_X1  g434(.A(new_n859), .B(G290), .ZN(new_n860));
  XNOR2_X1  g435(.A(new_n592), .B(KEYINPUT104), .ZN(new_n861));
  XNOR2_X1  g436(.A(new_n860), .B(new_n861), .ZN(new_n862));
  XOR2_X1   g437(.A(new_n862), .B(KEYINPUT42), .Z(new_n863));
  AND2_X1   g438(.A1(new_n858), .A2(new_n863), .ZN(new_n864));
  NOR2_X1   g439(.A1(new_n858), .A2(new_n863), .ZN(new_n865));
  OAI21_X1  g440(.A(G868), .B1(new_n864), .B2(new_n865), .ZN(new_n866));
  INV_X1    g441(.A(G868), .ZN(new_n867));
  NAND2_X1  g442(.A1(new_n813), .A2(new_n867), .ZN(new_n868));
  NAND2_X1  g443(.A1(new_n866), .A2(new_n868), .ZN(G295));
  NAND2_X1  g444(.A1(new_n866), .A2(new_n868), .ZN(G331));
  NAND2_X1  g445(.A1(new_n818), .A2(G171), .ZN(new_n871));
  NAND3_X1  g446(.A1(new_n816), .A2(G301), .A3(new_n817), .ZN(new_n872));
  NAND2_X1  g447(.A1(new_n871), .A2(new_n872), .ZN(new_n873));
  NAND2_X1  g448(.A1(new_n873), .A2(G286), .ZN(new_n874));
  INV_X1    g449(.A(new_n874), .ZN(new_n875));
  NOR2_X1   g450(.A1(new_n873), .A2(G286), .ZN(new_n876));
  OAI21_X1  g451(.A(new_n857), .B1(new_n875), .B2(new_n876), .ZN(new_n877));
  INV_X1    g452(.A(new_n876), .ZN(new_n878));
  INV_X1    g453(.A(new_n854), .ZN(new_n879));
  NAND3_X1  g454(.A1(new_n878), .A2(new_n879), .A3(new_n874), .ZN(new_n880));
  NAND2_X1  g455(.A1(new_n877), .A2(new_n880), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n881), .A2(new_n862), .ZN(new_n882));
  INV_X1    g457(.A(new_n862), .ZN(new_n883));
  NAND3_X1  g458(.A1(new_n877), .A2(new_n880), .A3(new_n883), .ZN(new_n884));
  NAND3_X1  g459(.A1(new_n882), .A2(new_n847), .A3(new_n884), .ZN(new_n885));
  NAND2_X1  g460(.A1(new_n885), .A2(KEYINPUT43), .ZN(new_n886));
  XNOR2_X1  g461(.A(KEYINPUT105), .B(KEYINPUT43), .ZN(new_n887));
  INV_X1    g462(.A(new_n887), .ZN(new_n888));
  NAND4_X1  g463(.A1(new_n882), .A2(new_n847), .A3(new_n884), .A4(new_n888), .ZN(new_n889));
  NAND3_X1  g464(.A1(new_n886), .A2(KEYINPUT44), .A3(new_n889), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n885), .A2(new_n887), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n891), .A2(new_n889), .ZN(new_n892));
  INV_X1    g467(.A(new_n892), .ZN(new_n893));
  OAI21_X1  g468(.A(new_n890), .B1(new_n893), .B2(KEYINPUT44), .ZN(G397));
  INV_X1    g469(.A(G1384), .ZN(new_n895));
  NAND2_X1  g470(.A1(new_n508), .A2(new_n895), .ZN(new_n896));
  INV_X1    g471(.A(KEYINPUT45), .ZN(new_n897));
  NAND2_X1  g472(.A1(new_n896), .A2(new_n897), .ZN(new_n898));
  NAND4_X1  g473(.A1(new_n476), .A2(G40), .A3(new_n482), .A4(new_n484), .ZN(new_n899));
  INV_X1    g474(.A(new_n899), .ZN(new_n900));
  NAND3_X1  g475(.A1(new_n898), .A2(KEYINPUT109), .A3(new_n900), .ZN(new_n901));
  NAND3_X1  g476(.A1(new_n508), .A2(KEYINPUT45), .A3(new_n895), .ZN(new_n902));
  INV_X1    g477(.A(KEYINPUT109), .ZN(new_n903));
  AOI21_X1  g478(.A(KEYINPUT45), .B1(new_n508), .B2(new_n895), .ZN(new_n904));
  OAI21_X1  g479(.A(new_n903), .B1(new_n904), .B2(new_n899), .ZN(new_n905));
  NAND3_X1  g480(.A1(new_n901), .A2(new_n902), .A3(new_n905), .ZN(new_n906));
  NAND2_X1  g481(.A1(new_n906), .A2(new_n765), .ZN(new_n907));
  INV_X1    g482(.A(KEYINPUT50), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n896), .A2(new_n908), .ZN(new_n909));
  NAND3_X1  g484(.A1(new_n508), .A2(KEYINPUT50), .A3(new_n895), .ZN(new_n910));
  AOI21_X1  g485(.A(new_n899), .B1(new_n909), .B2(new_n910), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n911), .A2(new_n749), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n907), .A2(new_n912), .ZN(new_n913));
  INV_X1    g488(.A(KEYINPUT121), .ZN(new_n914));
  NAND2_X1  g489(.A1(new_n913), .A2(new_n914), .ZN(new_n915));
  NAND3_X1  g490(.A1(new_n907), .A2(KEYINPUT121), .A3(new_n912), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n915), .A2(new_n916), .ZN(new_n917));
  NAND2_X1  g492(.A1(G286), .A2(G8), .ZN(new_n918));
  XOR2_X1   g493(.A(new_n918), .B(KEYINPUT122), .Z(new_n919));
  INV_X1    g494(.A(new_n919), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n917), .A2(new_n920), .ZN(new_n921));
  XOR2_X1   g496(.A(new_n919), .B(KEYINPUT125), .Z(new_n922));
  AOI21_X1  g497(.A(KEYINPUT124), .B1(new_n917), .B2(G8), .ZN(new_n923));
  AOI221_X4 g498(.A(new_n914), .B1(new_n911), .B2(new_n749), .C1(new_n906), .C2(new_n765), .ZN(new_n924));
  AOI21_X1  g499(.A(KEYINPUT121), .B1(new_n907), .B2(new_n912), .ZN(new_n925));
  OAI211_X1 g500(.A(KEYINPUT124), .B(G8), .C1(new_n924), .C2(new_n925), .ZN(new_n926));
  INV_X1    g501(.A(new_n926), .ZN(new_n927));
  OAI21_X1  g502(.A(new_n922), .B1(new_n923), .B2(new_n927), .ZN(new_n928));
  XNOR2_X1  g503(.A(KEYINPUT123), .B(KEYINPUT51), .ZN(new_n929));
  AOI21_X1  g504(.A(KEYINPUT126), .B1(new_n928), .B2(new_n929), .ZN(new_n930));
  INV_X1    g505(.A(new_n922), .ZN(new_n931));
  OAI21_X1  g506(.A(G8), .B1(new_n924), .B2(new_n925), .ZN(new_n932));
  INV_X1    g507(.A(KEYINPUT124), .ZN(new_n933));
  NAND2_X1  g508(.A1(new_n932), .A2(new_n933), .ZN(new_n934));
  AOI21_X1  g509(.A(new_n931), .B1(new_n934), .B2(new_n926), .ZN(new_n935));
  INV_X1    g510(.A(KEYINPUT126), .ZN(new_n936));
  INV_X1    g511(.A(new_n929), .ZN(new_n937));
  NOR3_X1   g512(.A1(new_n935), .A2(new_n936), .A3(new_n937), .ZN(new_n938));
  OAI21_X1  g513(.A(new_n921), .B1(new_n930), .B2(new_n938), .ZN(new_n939));
  NAND2_X1  g514(.A1(new_n913), .A2(G8), .ZN(new_n940));
  INV_X1    g515(.A(new_n940), .ZN(new_n941));
  NOR3_X1   g516(.A1(new_n941), .A2(KEYINPUT51), .A3(new_n920), .ZN(new_n942));
  INV_X1    g517(.A(new_n942), .ZN(new_n943));
  INV_X1    g518(.A(KEYINPUT53), .ZN(new_n944));
  NOR2_X1   g519(.A1(new_n904), .A2(new_n899), .ZN(new_n945));
  XOR2_X1   g520(.A(KEYINPUT106), .B(G1384), .Z(new_n946));
  NAND3_X1  g521(.A1(new_n508), .A2(KEYINPUT45), .A3(new_n946), .ZN(new_n947));
  NAND2_X1  g522(.A1(new_n945), .A2(new_n947), .ZN(new_n948));
  OAI21_X1  g523(.A(new_n944), .B1(new_n948), .B2(G2078), .ZN(new_n949));
  INV_X1    g524(.A(new_n910), .ZN(new_n950));
  AOI21_X1  g525(.A(KEYINPUT50), .B1(new_n508), .B2(new_n895), .ZN(new_n951));
  OAI21_X1  g526(.A(new_n900), .B1(new_n950), .B2(new_n951), .ZN(new_n952));
  NAND2_X1  g527(.A1(new_n952), .A2(new_n759), .ZN(new_n953));
  NAND2_X1  g528(.A1(new_n949), .A2(new_n953), .ZN(new_n954));
  INV_X1    g529(.A(new_n906), .ZN(new_n955));
  NOR2_X1   g530(.A1(new_n944), .A2(G2078), .ZN(new_n956));
  AOI21_X1  g531(.A(new_n954), .B1(new_n955), .B2(new_n956), .ZN(new_n957));
  OR2_X1    g532(.A1(new_n957), .A2(G301), .ZN(new_n958));
  OR2_X1    g533(.A1(new_n958), .A2(KEYINPUT62), .ZN(new_n959));
  INV_X1    g534(.A(KEYINPUT61), .ZN(new_n960));
  INV_X1    g535(.A(KEYINPUT112), .ZN(new_n961));
  AND3_X1   g536(.A1(new_n574), .A2(new_n961), .A3(new_n575), .ZN(new_n962));
  AOI21_X1  g537(.A(new_n961), .B1(new_n574), .B2(new_n575), .ZN(new_n963));
  INV_X1    g538(.A(new_n560), .ZN(new_n964));
  NOR3_X1   g539(.A1(new_n962), .A2(new_n963), .A3(new_n964), .ZN(new_n965));
  OAI211_X1 g540(.A(KEYINPUT57), .B(G299), .C1(new_n965), .C2(KEYINPUT111), .ZN(new_n966));
  INV_X1    g541(.A(KEYINPUT113), .ZN(new_n967));
  INV_X1    g542(.A(KEYINPUT57), .ZN(new_n968));
  INV_X1    g543(.A(KEYINPUT111), .ZN(new_n969));
  OAI21_X1  g544(.A(new_n968), .B1(new_n965), .B2(new_n969), .ZN(new_n970));
  NAND3_X1  g545(.A1(new_n966), .A2(new_n967), .A3(new_n970), .ZN(new_n971));
  NAND2_X1  g546(.A1(new_n574), .A2(new_n575), .ZN(new_n972));
  NAND2_X1  g547(.A1(new_n972), .A2(KEYINPUT112), .ZN(new_n973));
  NAND3_X1  g548(.A1(new_n574), .A2(new_n961), .A3(new_n575), .ZN(new_n974));
  NAND3_X1  g549(.A1(new_n973), .A2(new_n560), .A3(new_n974), .ZN(new_n975));
  AOI21_X1  g550(.A(KEYINPUT57), .B1(new_n975), .B2(KEYINPUT111), .ZN(new_n976));
  NAND2_X1  g551(.A1(G299), .A2(KEYINPUT57), .ZN(new_n977));
  AOI21_X1  g552(.A(new_n977), .B1(new_n975), .B2(new_n969), .ZN(new_n978));
  OAI21_X1  g553(.A(KEYINPUT113), .B1(new_n976), .B2(new_n978), .ZN(new_n979));
  XNOR2_X1  g554(.A(KEYINPUT56), .B(G2072), .ZN(new_n980));
  NAND4_X1  g555(.A1(new_n898), .A2(new_n900), .A3(new_n947), .A4(new_n980), .ZN(new_n981));
  INV_X1    g556(.A(KEYINPUT114), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n981), .A2(new_n982), .ZN(new_n983));
  NAND4_X1  g558(.A1(new_n945), .A2(KEYINPUT114), .A3(new_n947), .A4(new_n980), .ZN(new_n984));
  NAND2_X1  g559(.A1(new_n983), .A2(new_n984), .ZN(new_n985));
  NOR3_X1   g560(.A1(new_n911), .A2(KEYINPUT110), .A3(G1956), .ZN(new_n986));
  INV_X1    g561(.A(KEYINPUT110), .ZN(new_n987));
  AOI21_X1  g562(.A(new_n987), .B1(new_n952), .B2(new_n803), .ZN(new_n988));
  OAI21_X1  g563(.A(new_n985), .B1(new_n986), .B2(new_n988), .ZN(new_n989));
  AND3_X1   g564(.A1(new_n971), .A2(new_n979), .A3(new_n989), .ZN(new_n990));
  AOI21_X1  g565(.A(new_n989), .B1(new_n971), .B2(new_n979), .ZN(new_n991));
  OAI21_X1  g566(.A(new_n960), .B1(new_n990), .B2(new_n991), .ZN(new_n992));
  INV_X1    g567(.A(KEYINPUT60), .ZN(new_n993));
  INV_X1    g568(.A(KEYINPUT115), .ZN(new_n994));
  NOR2_X1   g569(.A1(new_n896), .A2(new_n899), .ZN(new_n995));
  INV_X1    g570(.A(new_n995), .ZN(new_n996));
  OAI21_X1  g571(.A(new_n994), .B1(new_n996), .B2(G2067), .ZN(new_n997));
  INV_X1    g572(.A(G1348), .ZN(new_n998));
  NAND2_X1  g573(.A1(new_n952), .A2(new_n998), .ZN(new_n999));
  INV_X1    g574(.A(G2067), .ZN(new_n1000));
  NAND3_X1  g575(.A1(new_n995), .A2(KEYINPUT115), .A3(new_n1000), .ZN(new_n1001));
  NAND3_X1  g576(.A1(new_n997), .A2(new_n999), .A3(new_n1001), .ZN(new_n1002));
  NAND2_X1  g577(.A1(new_n1002), .A2(new_n606), .ZN(new_n1003));
  NAND4_X1  g578(.A1(new_n997), .A2(new_n999), .A3(new_n605), .A4(new_n1001), .ZN(new_n1004));
  AOI21_X1  g579(.A(new_n993), .B1(new_n1003), .B2(new_n1004), .ZN(new_n1005));
  NOR3_X1   g580(.A1(new_n1002), .A2(KEYINPUT60), .A3(new_n605), .ZN(new_n1006));
  INV_X1    g581(.A(G1996), .ZN(new_n1007));
  NAND4_X1  g582(.A1(new_n898), .A2(new_n900), .A3(new_n1007), .A4(new_n947), .ZN(new_n1008));
  NAND2_X1  g583(.A1(new_n1008), .A2(KEYINPUT118), .ZN(new_n1009));
  XOR2_X1   g584(.A(KEYINPUT58), .B(G1341), .Z(new_n1010));
  NAND2_X1  g585(.A1(new_n996), .A2(new_n1010), .ZN(new_n1011));
  INV_X1    g586(.A(KEYINPUT118), .ZN(new_n1012));
  NAND4_X1  g587(.A1(new_n945), .A2(new_n1012), .A3(new_n1007), .A4(new_n947), .ZN(new_n1013));
  NAND3_X1  g588(.A1(new_n1009), .A2(new_n1011), .A3(new_n1013), .ZN(new_n1014));
  AND4_X1   g589(.A1(KEYINPUT119), .A2(new_n547), .A3(new_n548), .A4(new_n549), .ZN(new_n1015));
  AND3_X1   g590(.A1(new_n1014), .A2(new_n1015), .A3(KEYINPUT59), .ZN(new_n1016));
  AOI21_X1  g591(.A(KEYINPUT59), .B1(new_n1014), .B2(new_n1015), .ZN(new_n1017));
  NOR4_X1   g592(.A1(new_n1005), .A2(new_n1006), .A3(new_n1016), .A4(new_n1017), .ZN(new_n1018));
  INV_X1    g593(.A(KEYINPUT120), .ZN(new_n1019));
  INV_X1    g594(.A(new_n989), .ZN(new_n1020));
  AOI21_X1  g595(.A(new_n967), .B1(new_n966), .B2(new_n970), .ZN(new_n1021));
  NOR3_X1   g596(.A1(new_n976), .A2(new_n978), .A3(KEYINPUT113), .ZN(new_n1022));
  OAI21_X1  g597(.A(new_n1020), .B1(new_n1021), .B2(new_n1022), .ZN(new_n1023));
  AOI21_X1  g598(.A(new_n1019), .B1(new_n1023), .B2(KEYINPUT61), .ZN(new_n1024));
  NOR3_X1   g599(.A1(new_n991), .A2(KEYINPUT120), .A3(new_n960), .ZN(new_n1025));
  OAI211_X1 g600(.A(new_n992), .B(new_n1018), .C1(new_n1024), .C2(new_n1025), .ZN(new_n1026));
  XNOR2_X1  g601(.A(new_n1003), .B(KEYINPUT116), .ZN(new_n1027));
  XNOR2_X1  g602(.A(new_n989), .B(KEYINPUT117), .ZN(new_n1028));
  NOR2_X1   g603(.A1(new_n1021), .A2(new_n1022), .ZN(new_n1029));
  AOI22_X1  g604(.A1(new_n1023), .A2(new_n1027), .B1(new_n1028), .B2(new_n1029), .ZN(new_n1030));
  NAND2_X1  g605(.A1(new_n1026), .A2(new_n1030), .ZN(new_n1031));
  NAND2_X1  g606(.A1(new_n508), .A2(new_n946), .ZN(new_n1032));
  NAND2_X1  g607(.A1(new_n1032), .A2(new_n897), .ZN(new_n1033));
  NAND4_X1  g608(.A1(new_n1033), .A2(new_n900), .A3(new_n947), .A4(new_n956), .ZN(new_n1034));
  NAND3_X1  g609(.A1(new_n949), .A2(new_n953), .A3(new_n1034), .ZN(new_n1035));
  OAI21_X1  g610(.A(new_n958), .B1(G171), .B2(new_n1035), .ZN(new_n1036));
  XNOR2_X1  g611(.A(KEYINPUT127), .B(KEYINPUT54), .ZN(new_n1037));
  INV_X1    g612(.A(KEYINPUT54), .ZN(new_n1038));
  AOI21_X1  g613(.A(new_n1038), .B1(new_n957), .B2(G301), .ZN(new_n1039));
  NAND2_X1  g614(.A1(new_n1035), .A2(G171), .ZN(new_n1040));
  AOI22_X1  g615(.A1(new_n1036), .A2(new_n1037), .B1(new_n1039), .B2(new_n1040), .ZN(new_n1041));
  NAND2_X1  g616(.A1(new_n1031), .A2(new_n1041), .ZN(new_n1042));
  NAND4_X1  g617(.A1(new_n939), .A2(new_n943), .A3(new_n959), .A4(new_n1042), .ZN(new_n1043));
  INV_X1    g618(.A(KEYINPUT62), .ZN(new_n1044));
  OR2_X1    g619(.A1(new_n958), .A2(new_n1044), .ZN(new_n1045));
  INV_X1    g620(.A(new_n921), .ZN(new_n1046));
  NAND3_X1  g621(.A1(new_n928), .A2(KEYINPUT126), .A3(new_n929), .ZN(new_n1047));
  OAI21_X1  g622(.A(new_n936), .B1(new_n935), .B2(new_n937), .ZN(new_n1048));
  AOI21_X1  g623(.A(new_n1046), .B1(new_n1047), .B2(new_n1048), .ZN(new_n1049));
  OAI21_X1  g624(.A(new_n1045), .B1(new_n1049), .B2(new_n942), .ZN(new_n1050));
  INV_X1    g625(.A(G8), .ZN(new_n1051));
  OR2_X1    g626(.A1(new_n952), .A2(G2090), .ZN(new_n1052));
  NAND2_X1  g627(.A1(new_n948), .A2(new_n696), .ZN(new_n1053));
  AOI21_X1  g628(.A(new_n1051), .B1(new_n1052), .B2(new_n1053), .ZN(new_n1054));
  NOR2_X1   g629(.A1(G166), .A2(new_n1051), .ZN(new_n1055));
  XNOR2_X1  g630(.A(new_n1055), .B(KEYINPUT55), .ZN(new_n1056));
  XNOR2_X1  g631(.A(new_n1054), .B(new_n1056), .ZN(new_n1057));
  XNOR2_X1  g632(.A(KEYINPUT108), .B(G1981), .ZN(new_n1058));
  NAND2_X1  g633(.A1(new_n592), .A2(new_n1058), .ZN(new_n1059));
  INV_X1    g634(.A(G1981), .ZN(new_n1060));
  OAI21_X1  g635(.A(new_n1059), .B1(new_n1060), .B2(new_n592), .ZN(new_n1061));
  XNOR2_X1  g636(.A(new_n1061), .B(KEYINPUT49), .ZN(new_n1062));
  NOR2_X1   g637(.A1(new_n995), .A2(new_n1051), .ZN(new_n1063));
  NAND2_X1  g638(.A1(new_n1062), .A2(new_n1063), .ZN(new_n1064));
  INV_X1    g639(.A(G1976), .ZN(new_n1065));
  OAI21_X1  g640(.A(new_n1063), .B1(G288), .B2(new_n1065), .ZN(new_n1066));
  NAND2_X1  g641(.A1(new_n1066), .A2(KEYINPUT52), .ZN(new_n1067));
  INV_X1    g642(.A(KEYINPUT52), .ZN(new_n1068));
  OAI21_X1  g643(.A(new_n1068), .B1(new_n685), .B2(G1976), .ZN(new_n1069));
  OAI211_X1 g644(.A(new_n1064), .B(new_n1067), .C1(new_n1066), .C2(new_n1069), .ZN(new_n1070));
  NOR2_X1   g645(.A1(new_n1057), .A2(new_n1070), .ZN(new_n1071));
  NAND3_X1  g646(.A1(new_n1043), .A2(new_n1050), .A3(new_n1071), .ZN(new_n1072));
  NAND2_X1  g647(.A1(new_n1054), .A2(new_n1056), .ZN(new_n1073));
  OR2_X1    g648(.A1(new_n1070), .A2(new_n1073), .ZN(new_n1074));
  NAND3_X1  g649(.A1(new_n1071), .A2(G168), .A3(new_n941), .ZN(new_n1075));
  XNOR2_X1  g650(.A(new_n1075), .B(KEYINPUT63), .ZN(new_n1076));
  NAND3_X1  g651(.A1(new_n1064), .A2(new_n1065), .A3(new_n685), .ZN(new_n1077));
  NAND2_X1  g652(.A1(new_n1077), .A2(new_n1059), .ZN(new_n1078));
  AOI21_X1  g653(.A(new_n1076), .B1(new_n1063), .B2(new_n1078), .ZN(new_n1079));
  NAND3_X1  g654(.A1(new_n1072), .A2(new_n1074), .A3(new_n1079), .ZN(new_n1080));
  INV_X1    g655(.A(G1986), .ZN(new_n1081));
  NOR2_X1   g656(.A1(new_n1033), .A2(new_n899), .ZN(new_n1082));
  NAND3_X1  g657(.A1(new_n681), .A2(new_n1081), .A3(new_n1082), .ZN(new_n1083));
  NAND3_X1  g658(.A1(G290), .A2(G1986), .A3(new_n1082), .ZN(new_n1084));
  NAND2_X1  g659(.A1(new_n1083), .A2(new_n1084), .ZN(new_n1085));
  XNOR2_X1  g660(.A(new_n1085), .B(KEYINPUT107), .ZN(new_n1086));
  NAND2_X1  g661(.A1(new_n726), .A2(new_n1007), .ZN(new_n1087));
  XNOR2_X1  g662(.A(new_n742), .B(G2067), .ZN(new_n1088));
  NAND2_X1  g663(.A1(new_n725), .A2(G1996), .ZN(new_n1089));
  NAND3_X1  g664(.A1(new_n1087), .A2(new_n1088), .A3(new_n1089), .ZN(new_n1090));
  INV_X1    g665(.A(new_n711), .ZN(new_n1091));
  XNOR2_X1  g666(.A(new_n709), .B(new_n1091), .ZN(new_n1092));
  OAI21_X1  g667(.A(new_n1082), .B1(new_n1090), .B2(new_n1092), .ZN(new_n1093));
  AND2_X1   g668(.A1(new_n1086), .A2(new_n1093), .ZN(new_n1094));
  NAND2_X1  g669(.A1(new_n1080), .A2(new_n1094), .ZN(new_n1095));
  NAND2_X1  g670(.A1(new_n709), .A2(new_n1091), .ZN(new_n1096));
  OAI22_X1  g671(.A1(new_n1090), .A2(new_n1096), .B1(G2067), .B2(new_n826), .ZN(new_n1097));
  AND2_X1   g672(.A1(new_n1097), .A2(new_n1082), .ZN(new_n1098));
  NOR3_X1   g673(.A1(new_n1033), .A2(G1996), .A3(new_n899), .ZN(new_n1099));
  OR2_X1    g674(.A1(new_n1099), .A2(KEYINPUT46), .ZN(new_n1100));
  INV_X1    g675(.A(new_n1088), .ZN(new_n1101));
  OAI21_X1  g676(.A(new_n1082), .B1(new_n725), .B2(new_n1101), .ZN(new_n1102));
  NAND2_X1  g677(.A1(new_n1099), .A2(KEYINPUT46), .ZN(new_n1103));
  NAND3_X1  g678(.A1(new_n1100), .A2(new_n1102), .A3(new_n1103), .ZN(new_n1104));
  XOR2_X1   g679(.A(new_n1104), .B(KEYINPUT47), .Z(new_n1105));
  XNOR2_X1  g680(.A(new_n1083), .B(KEYINPUT48), .ZN(new_n1106));
  AOI211_X1 g681(.A(new_n1098), .B(new_n1105), .C1(new_n1093), .C2(new_n1106), .ZN(new_n1107));
  NAND2_X1  g682(.A1(new_n1095), .A2(new_n1107), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g683(.A(new_n458), .ZN(new_n1110));
  OR2_X1    g684(.A1(G229), .A2(new_n1110), .ZN(new_n1111));
  AOI21_X1  g685(.A(new_n1111), .B1(new_n849), .B2(new_n850), .ZN(new_n1112));
  NOR2_X1   g686(.A1(G401), .A2(G227), .ZN(new_n1113));
  NAND3_X1  g687(.A1(new_n1112), .A2(new_n892), .A3(new_n1113), .ZN(G225));
  INV_X1    g688(.A(G225), .ZN(G308));
endmodule


