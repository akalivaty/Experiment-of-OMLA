

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300,
         n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311,
         n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322,
         n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333,
         n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344,
         n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355,
         n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
         n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
         n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
         n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
         n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410,
         n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421,
         n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432,
         n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443,
         n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454,
         n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465,
         n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
         n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487,
         n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
         n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
         n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579;

  XOR2_X1 U322 ( .A(n374), .B(n373), .Z(n290) );
  XOR2_X1 U323 ( .A(G197GAT), .B(G113GAT), .Z(n291) );
  XNOR2_X1 U324 ( .A(n372), .B(KEYINPUT107), .ZN(n373) );
  NOR2_X1 U325 ( .A1(n401), .A2(n400), .ZN(n402) );
  XNOR2_X1 U326 ( .A(n375), .B(n291), .ZN(n353) );
  XNOR2_X1 U327 ( .A(n354), .B(n353), .ZN(n356) );
  NOR2_X1 U328 ( .A1(n429), .A2(n514), .ZN(n561) );
  XOR2_X1 U329 ( .A(n567), .B(KEYINPUT41), .Z(n548) );
  XOR2_X1 U330 ( .A(n428), .B(n427), .Z(n514) );
  XOR2_X1 U331 ( .A(n463), .B(KEYINPUT28), .Z(n521) );
  XNOR2_X1 U332 ( .A(n456), .B(G190GAT), .ZN(n457) );
  XNOR2_X1 U333 ( .A(n458), .B(n457), .ZN(G1351GAT) );
  INV_X1 U334 ( .A(KEYINPUT119), .ZN(n448) );
  XOR2_X1 U335 ( .A(KEYINPUT64), .B(KEYINPUT85), .Z(n293) );
  XNOR2_X1 U336 ( .A(G71GAT), .B(KEYINPUT84), .ZN(n292) );
  XNOR2_X1 U337 ( .A(n293), .B(n292), .ZN(n297) );
  XOR2_X1 U338 ( .A(G176GAT), .B(KEYINPUT81), .Z(n295) );
  XNOR2_X1 U339 ( .A(KEYINPUT82), .B(KEYINPUT20), .ZN(n294) );
  XNOR2_X1 U340 ( .A(n295), .B(n294), .ZN(n296) );
  XOR2_X1 U341 ( .A(n297), .B(n296), .Z(n309) );
  XNOR2_X1 U342 ( .A(KEYINPUT19), .B(KEYINPUT18), .ZN(n298) );
  XNOR2_X1 U343 ( .A(n298), .B(KEYINPUT17), .ZN(n299) );
  XOR2_X1 U344 ( .A(n299), .B(KEYINPUT83), .Z(n301) );
  XNOR2_X1 U345 ( .A(G183GAT), .B(G190GAT), .ZN(n300) );
  XNOR2_X1 U346 ( .A(n301), .B(n300), .ZN(n317) );
  XOR2_X1 U347 ( .A(G99GAT), .B(G134GAT), .Z(n303) );
  XNOR2_X1 U348 ( .A(G43GAT), .B(G15GAT), .ZN(n302) );
  XNOR2_X1 U349 ( .A(n303), .B(n302), .ZN(n304) );
  XOR2_X1 U350 ( .A(G169GAT), .B(n304), .Z(n306) );
  NAND2_X1 U351 ( .A1(G227GAT), .A2(G233GAT), .ZN(n305) );
  XNOR2_X1 U352 ( .A(n306), .B(n305), .ZN(n307) );
  XNOR2_X1 U353 ( .A(n317), .B(n307), .ZN(n308) );
  XNOR2_X1 U354 ( .A(n309), .B(n308), .ZN(n313) );
  XOR2_X1 U355 ( .A(KEYINPUT80), .B(G127GAT), .Z(n311) );
  XNOR2_X1 U356 ( .A(KEYINPUT0), .B(G120GAT), .ZN(n310) );
  XNOR2_X1 U357 ( .A(n311), .B(n310), .ZN(n312) );
  XOR2_X1 U358 ( .A(G113GAT), .B(n312), .Z(n405) );
  XOR2_X1 U359 ( .A(n313), .B(n405), .Z(n530) );
  XOR2_X1 U360 ( .A(G92GAT), .B(G64GAT), .Z(n315) );
  XNOR2_X1 U361 ( .A(G204GAT), .B(KEYINPUT74), .ZN(n314) );
  XNOR2_X1 U362 ( .A(n315), .B(n314), .ZN(n316) );
  XOR2_X1 U363 ( .A(G176GAT), .B(n316), .Z(n365) );
  XNOR2_X1 U364 ( .A(n317), .B(n365), .ZN(n326) );
  XOR2_X1 U365 ( .A(G211GAT), .B(KEYINPUT21), .Z(n319) );
  XNOR2_X1 U366 ( .A(G197GAT), .B(G218GAT), .ZN(n318) );
  XNOR2_X1 U367 ( .A(n319), .B(n318), .ZN(n439) );
  XOR2_X1 U368 ( .A(n439), .B(KEYINPUT94), .Z(n321) );
  NAND2_X1 U369 ( .A1(G226GAT), .A2(G233GAT), .ZN(n320) );
  XNOR2_X1 U370 ( .A(n321), .B(n320), .ZN(n322) );
  XOR2_X1 U371 ( .A(n322), .B(KEYINPUT93), .Z(n324) );
  XOR2_X1 U372 ( .A(G169GAT), .B(G8GAT), .Z(n350) );
  XNOR2_X1 U373 ( .A(G36GAT), .B(n350), .ZN(n323) );
  XNOR2_X1 U374 ( .A(n324), .B(n323), .ZN(n325) );
  XOR2_X1 U375 ( .A(n326), .B(n325), .Z(n517) );
  INV_X1 U376 ( .A(n517), .ZN(n403) );
  XNOR2_X1 U377 ( .A(G36GAT), .B(KEYINPUT7), .ZN(n327) );
  XNOR2_X1 U378 ( .A(n327), .B(G29GAT), .ZN(n328) );
  XOR2_X1 U379 ( .A(n328), .B(KEYINPUT8), .Z(n330) );
  XNOR2_X1 U380 ( .A(G43GAT), .B(G50GAT), .ZN(n329) );
  XOR2_X1 U381 ( .A(n330), .B(n329), .Z(n355) );
  XOR2_X1 U382 ( .A(KEYINPUT75), .B(KEYINPUT11), .Z(n332) );
  XNOR2_X1 U383 ( .A(G162GAT), .B(G92GAT), .ZN(n331) );
  XNOR2_X1 U384 ( .A(n332), .B(n331), .ZN(n333) );
  XOR2_X1 U385 ( .A(n355), .B(n333), .Z(n346) );
  XOR2_X1 U386 ( .A(KEYINPUT67), .B(KEYINPUT10), .Z(n335) );
  XNOR2_X1 U387 ( .A(G190GAT), .B(G218GAT), .ZN(n334) );
  XNOR2_X1 U388 ( .A(n335), .B(n334), .ZN(n339) );
  XOR2_X1 U389 ( .A(KEYINPUT76), .B(KEYINPUT9), .Z(n337) );
  XNOR2_X1 U390 ( .A(G106GAT), .B(KEYINPUT68), .ZN(n336) );
  XNOR2_X1 U391 ( .A(n337), .B(n336), .ZN(n338) );
  XOR2_X1 U392 ( .A(n339), .B(n338), .Z(n344) );
  XOR2_X1 U393 ( .A(G134GAT), .B(KEYINPUT77), .Z(n420) );
  XOR2_X1 U394 ( .A(G99GAT), .B(G85GAT), .Z(n358) );
  XOR2_X1 U395 ( .A(n358), .B(KEYINPUT65), .Z(n341) );
  NAND2_X1 U396 ( .A1(G232GAT), .A2(G233GAT), .ZN(n340) );
  XNOR2_X1 U397 ( .A(n341), .B(n340), .ZN(n342) );
  XNOR2_X1 U398 ( .A(n420), .B(n342), .ZN(n343) );
  XNOR2_X1 U399 ( .A(n344), .B(n343), .ZN(n345) );
  XNOR2_X1 U400 ( .A(n346), .B(n345), .ZN(n553) );
  XOR2_X1 U401 ( .A(KEYINPUT69), .B(KEYINPUT29), .Z(n348) );
  NAND2_X1 U402 ( .A1(G229GAT), .A2(G233GAT), .ZN(n347) );
  XNOR2_X1 U403 ( .A(n348), .B(n347), .ZN(n349) );
  XOR2_X1 U404 ( .A(n349), .B(KEYINPUT30), .Z(n352) );
  XOR2_X1 U405 ( .A(G141GAT), .B(G22GAT), .Z(n435) );
  XNOR2_X1 U406 ( .A(n435), .B(n350), .ZN(n351) );
  XNOR2_X1 U407 ( .A(n352), .B(n351), .ZN(n354) );
  XOR2_X1 U408 ( .A(G15GAT), .B(G1GAT), .Z(n375) );
  XOR2_X1 U409 ( .A(n356), .B(n355), .Z(n500) );
  INV_X1 U410 ( .A(n500), .ZN(n562) );
  XNOR2_X1 U411 ( .A(G71GAT), .B(G57GAT), .ZN(n357) );
  XNOR2_X1 U412 ( .A(n357), .B(KEYINPUT13), .ZN(n376) );
  XNOR2_X1 U413 ( .A(KEYINPUT71), .B(n376), .ZN(n360) );
  XOR2_X1 U414 ( .A(G120GAT), .B(n358), .Z(n359) );
  XNOR2_X1 U415 ( .A(n360), .B(n359), .ZN(n364) );
  XOR2_X1 U416 ( .A(KEYINPUT31), .B(KEYINPUT32), .Z(n362) );
  NAND2_X1 U417 ( .A1(G230GAT), .A2(G233GAT), .ZN(n361) );
  XOR2_X1 U418 ( .A(n362), .B(n361), .Z(n363) );
  XNOR2_X1 U419 ( .A(n364), .B(n363), .ZN(n367) );
  XNOR2_X1 U420 ( .A(n365), .B(KEYINPUT33), .ZN(n366) );
  XNOR2_X1 U421 ( .A(n367), .B(n366), .ZN(n371) );
  XOR2_X1 U422 ( .A(G148GAT), .B(G106GAT), .Z(n369) );
  XNOR2_X1 U423 ( .A(KEYINPUT73), .B(G78GAT), .ZN(n368) );
  XNOR2_X1 U424 ( .A(n369), .B(n368), .ZN(n370) );
  XNOR2_X1 U425 ( .A(KEYINPUT72), .B(n370), .ZN(n430) );
  XNOR2_X1 U426 ( .A(n371), .B(n430), .ZN(n393) );
  INV_X1 U427 ( .A(n393), .ZN(n567) );
  NAND2_X1 U428 ( .A1(n562), .A2(n548), .ZN(n374) );
  XOR2_X1 U429 ( .A(KEYINPUT46), .B(KEYINPUT108), .Z(n372) );
  NOR2_X1 U430 ( .A1(n553), .A2(n290), .ZN(n391) );
  XOR2_X1 U431 ( .A(n376), .B(n375), .Z(n378) );
  NAND2_X1 U432 ( .A1(G231GAT), .A2(G233GAT), .ZN(n377) );
  XNOR2_X1 U433 ( .A(n378), .B(n377), .ZN(n382) );
  XOR2_X1 U434 ( .A(KEYINPUT12), .B(KEYINPUT14), .Z(n380) );
  XNOR2_X1 U435 ( .A(KEYINPUT15), .B(KEYINPUT78), .ZN(n379) );
  XNOR2_X1 U436 ( .A(n380), .B(n379), .ZN(n381) );
  XOR2_X1 U437 ( .A(n382), .B(n381), .Z(n390) );
  XOR2_X1 U438 ( .A(G211GAT), .B(G78GAT), .Z(n384) );
  XNOR2_X1 U439 ( .A(G22GAT), .B(G155GAT), .ZN(n383) );
  XNOR2_X1 U440 ( .A(n384), .B(n383), .ZN(n388) );
  XOR2_X1 U441 ( .A(G64GAT), .B(G183GAT), .Z(n386) );
  XNOR2_X1 U442 ( .A(G8GAT), .B(G127GAT), .ZN(n385) );
  XNOR2_X1 U443 ( .A(n386), .B(n385), .ZN(n387) );
  XNOR2_X1 U444 ( .A(n388), .B(n387), .ZN(n389) );
  XOR2_X1 U445 ( .A(n390), .B(n389), .Z(n572) );
  INV_X1 U446 ( .A(n572), .ZN(n486) );
  NAND2_X1 U447 ( .A1(n391), .A2(n486), .ZN(n392) );
  XNOR2_X1 U448 ( .A(n392), .B(KEYINPUT47), .ZN(n401) );
  XOR2_X1 U449 ( .A(n500), .B(KEYINPUT70), .Z(n557) );
  XNOR2_X1 U450 ( .A(KEYINPUT109), .B(KEYINPUT45), .ZN(n394) );
  XNOR2_X1 U451 ( .A(n394), .B(KEYINPUT66), .ZN(n397) );
  XNOR2_X1 U452 ( .A(n553), .B(KEYINPUT99), .ZN(n395) );
  XNOR2_X1 U453 ( .A(n395), .B(KEYINPUT36), .ZN(n577) );
  NOR2_X1 U454 ( .A1(n486), .A2(n577), .ZN(n396) );
  XOR2_X1 U455 ( .A(n397), .B(n396), .Z(n398) );
  NAND2_X1 U456 ( .A1(n393), .A2(n398), .ZN(n399) );
  NOR2_X1 U457 ( .A1(n557), .A2(n399), .ZN(n400) );
  XNOR2_X1 U458 ( .A(n402), .B(KEYINPUT48), .ZN(n527) );
  NOR2_X1 U459 ( .A1(n403), .A2(n527), .ZN(n404) );
  XOR2_X1 U460 ( .A(KEYINPUT54), .B(n404), .Z(n429) );
  INV_X1 U461 ( .A(n405), .ZN(n428) );
  XOR2_X1 U462 ( .A(KEYINPUT91), .B(KEYINPUT6), .Z(n407) );
  XNOR2_X1 U463 ( .A(KEYINPUT90), .B(KEYINPUT89), .ZN(n406) );
  XNOR2_X1 U464 ( .A(n407), .B(n406), .ZN(n411) );
  XOR2_X1 U465 ( .A(G57GAT), .B(G148GAT), .Z(n409) );
  XNOR2_X1 U466 ( .A(G141GAT), .B(G1GAT), .ZN(n408) );
  XNOR2_X1 U467 ( .A(n409), .B(n408), .ZN(n410) );
  XOR2_X1 U468 ( .A(n411), .B(n410), .Z(n419) );
  XOR2_X1 U469 ( .A(KEYINPUT2), .B(G162GAT), .Z(n413) );
  XNOR2_X1 U470 ( .A(KEYINPUT3), .B(G155GAT), .ZN(n412) );
  XNOR2_X1 U471 ( .A(n413), .B(n412), .ZN(n414) );
  XOR2_X1 U472 ( .A(KEYINPUT86), .B(n414), .Z(n431) );
  XOR2_X1 U473 ( .A(KEYINPUT1), .B(KEYINPUT5), .Z(n416) );
  XNOR2_X1 U474 ( .A(KEYINPUT4), .B(KEYINPUT88), .ZN(n415) );
  XNOR2_X1 U475 ( .A(n416), .B(n415), .ZN(n417) );
  XNOR2_X1 U476 ( .A(n431), .B(n417), .ZN(n418) );
  XNOR2_X1 U477 ( .A(n419), .B(n418), .ZN(n424) );
  XOR2_X1 U478 ( .A(n420), .B(KEYINPUT92), .Z(n422) );
  NAND2_X1 U479 ( .A1(G225GAT), .A2(G233GAT), .ZN(n421) );
  XNOR2_X1 U480 ( .A(n422), .B(n421), .ZN(n423) );
  XOR2_X1 U481 ( .A(n424), .B(n423), .Z(n426) );
  XNOR2_X1 U482 ( .A(G29GAT), .B(G85GAT), .ZN(n425) );
  XNOR2_X1 U483 ( .A(n426), .B(n425), .ZN(n427) );
  XOR2_X1 U484 ( .A(n431), .B(n430), .Z(n443) );
  XOR2_X1 U485 ( .A(KEYINPUT22), .B(KEYINPUT24), .Z(n433) );
  XNOR2_X1 U486 ( .A(G50GAT), .B(KEYINPUT87), .ZN(n432) );
  XNOR2_X1 U487 ( .A(n433), .B(n432), .ZN(n434) );
  XOR2_X1 U488 ( .A(n435), .B(n434), .Z(n437) );
  NAND2_X1 U489 ( .A1(G228GAT), .A2(G233GAT), .ZN(n436) );
  XNOR2_X1 U490 ( .A(n437), .B(n436), .ZN(n438) );
  XOR2_X1 U491 ( .A(n438), .B(KEYINPUT23), .Z(n441) );
  XNOR2_X1 U492 ( .A(n439), .B(G204GAT), .ZN(n440) );
  XNOR2_X1 U493 ( .A(n441), .B(n440), .ZN(n442) );
  XNOR2_X1 U494 ( .A(n443), .B(n442), .ZN(n463) );
  NAND2_X1 U495 ( .A1(n561), .A2(n463), .ZN(n445) );
  XOR2_X1 U496 ( .A(KEYINPUT55), .B(KEYINPUT118), .Z(n444) );
  XNOR2_X1 U497 ( .A(n445), .B(n444), .ZN(n446) );
  NOR2_X1 U498 ( .A1(n530), .A2(n446), .ZN(n447) );
  XNOR2_X1 U499 ( .A(n448), .B(n447), .ZN(n558) );
  NAND2_X1 U500 ( .A1(n558), .A2(n548), .ZN(n452) );
  XOR2_X1 U501 ( .A(KEYINPUT120), .B(KEYINPUT57), .Z(n450) );
  XNOR2_X1 U502 ( .A(G176GAT), .B(KEYINPUT56), .ZN(n449) );
  XNOR2_X1 U503 ( .A(n450), .B(n449), .ZN(n451) );
  XNOR2_X1 U504 ( .A(n452), .B(n451), .ZN(G1349GAT) );
  NAND2_X1 U505 ( .A1(n558), .A2(n572), .ZN(n455) );
  XOR2_X1 U506 ( .A(KEYINPUT121), .B(KEYINPUT122), .Z(n453) );
  XNOR2_X1 U507 ( .A(n453), .B(G183GAT), .ZN(n454) );
  XNOR2_X1 U508 ( .A(n455), .B(n454), .ZN(G1350GAT) );
  NAND2_X1 U509 ( .A1(n558), .A2(n553), .ZN(n458) );
  XOR2_X1 U510 ( .A(KEYINPUT58), .B(KEYINPUT123), .Z(n456) );
  XOR2_X1 U511 ( .A(KEYINPUT96), .B(KEYINPUT34), .Z(n476) );
  NAND2_X1 U512 ( .A1(n393), .A2(n557), .ZN(n489) );
  INV_X1 U513 ( .A(n521), .ZN(n528) );
  INV_X1 U514 ( .A(n530), .ZN(n519) );
  XNOR2_X1 U515 ( .A(n517), .B(KEYINPUT27), .ZN(n461) );
  NAND2_X1 U516 ( .A1(n461), .A2(n514), .ZN(n526) );
  NOR2_X1 U517 ( .A1(n519), .A2(n526), .ZN(n459) );
  NAND2_X1 U518 ( .A1(n528), .A2(n459), .ZN(n470) );
  NOR2_X1 U519 ( .A1(n519), .A2(n463), .ZN(n460) );
  XNOR2_X1 U520 ( .A(n460), .B(KEYINPUT26), .ZN(n560) );
  NAND2_X1 U521 ( .A1(n560), .A2(n461), .ZN(n466) );
  NAND2_X1 U522 ( .A1(n519), .A2(n517), .ZN(n462) );
  NAND2_X1 U523 ( .A1(n463), .A2(n462), .ZN(n464) );
  XOR2_X1 U524 ( .A(KEYINPUT25), .B(n464), .Z(n465) );
  NAND2_X1 U525 ( .A1(n466), .A2(n465), .ZN(n468) );
  INV_X1 U526 ( .A(n514), .ZN(n467) );
  NAND2_X1 U527 ( .A1(n468), .A2(n467), .ZN(n469) );
  NAND2_X1 U528 ( .A1(n470), .A2(n469), .ZN(n471) );
  XNOR2_X1 U529 ( .A(n471), .B(KEYINPUT95), .ZN(n484) );
  XNOR2_X1 U530 ( .A(KEYINPUT16), .B(KEYINPUT79), .ZN(n473) );
  NOR2_X1 U531 ( .A1(n553), .A2(n486), .ZN(n472) );
  XNOR2_X1 U532 ( .A(n473), .B(n472), .ZN(n474) );
  OR2_X1 U533 ( .A1(n484), .A2(n474), .ZN(n502) );
  NOR2_X1 U534 ( .A1(n489), .A2(n502), .ZN(n482) );
  NAND2_X1 U535 ( .A1(n482), .A2(n514), .ZN(n475) );
  XNOR2_X1 U536 ( .A(n476), .B(n475), .ZN(n477) );
  XOR2_X1 U537 ( .A(G1GAT), .B(n477), .Z(G1324GAT) );
  NAND2_X1 U538 ( .A1(n517), .A2(n482), .ZN(n478) );
  XNOR2_X1 U539 ( .A(n478), .B(G8GAT), .ZN(G1325GAT) );
  XOR2_X1 U540 ( .A(KEYINPUT97), .B(KEYINPUT35), .Z(n480) );
  NAND2_X1 U541 ( .A1(n482), .A2(n519), .ZN(n479) );
  XNOR2_X1 U542 ( .A(n480), .B(n479), .ZN(n481) );
  XOR2_X1 U543 ( .A(G15GAT), .B(n481), .Z(G1326GAT) );
  NAND2_X1 U544 ( .A1(n482), .A2(n521), .ZN(n483) );
  XNOR2_X1 U545 ( .A(n483), .B(G22GAT), .ZN(G1327GAT) );
  XOR2_X1 U546 ( .A(G29GAT), .B(KEYINPUT98), .Z(n492) );
  NOR2_X1 U547 ( .A1(n577), .A2(n484), .ZN(n485) );
  NAND2_X1 U548 ( .A1(n486), .A2(n485), .ZN(n487) );
  XNOR2_X1 U549 ( .A(KEYINPUT37), .B(n487), .ZN(n488) );
  XOR2_X1 U550 ( .A(KEYINPUT100), .B(n488), .Z(n513) );
  NOR2_X1 U551 ( .A1(n489), .A2(n513), .ZN(n490) );
  XNOR2_X1 U552 ( .A(n490), .B(KEYINPUT38), .ZN(n498) );
  NAND2_X1 U553 ( .A1(n498), .A2(n514), .ZN(n491) );
  XNOR2_X1 U554 ( .A(n492), .B(n491), .ZN(n494) );
  XOR2_X1 U555 ( .A(KEYINPUT39), .B(KEYINPUT101), .Z(n493) );
  XNOR2_X1 U556 ( .A(n494), .B(n493), .ZN(G1328GAT) );
  NAND2_X1 U557 ( .A1(n498), .A2(n517), .ZN(n495) );
  XNOR2_X1 U558 ( .A(n495), .B(G36GAT), .ZN(G1329GAT) );
  NAND2_X1 U559 ( .A1(n498), .A2(n519), .ZN(n496) );
  XNOR2_X1 U560 ( .A(n496), .B(KEYINPUT40), .ZN(n497) );
  XNOR2_X1 U561 ( .A(G43GAT), .B(n497), .ZN(G1330GAT) );
  NAND2_X1 U562 ( .A1(n521), .A2(n498), .ZN(n499) );
  XNOR2_X1 U563 ( .A(G50GAT), .B(n499), .ZN(G1331GAT) );
  XNOR2_X1 U564 ( .A(G57GAT), .B(KEYINPUT42), .ZN(n504) );
  NAND2_X1 U565 ( .A1(n548), .A2(n500), .ZN(n501) );
  XNOR2_X1 U566 ( .A(n501), .B(KEYINPUT102), .ZN(n512) );
  NOR2_X1 U567 ( .A1(n512), .A2(n502), .ZN(n509) );
  NAND2_X1 U568 ( .A1(n509), .A2(n514), .ZN(n503) );
  XNOR2_X1 U569 ( .A(n504), .B(n503), .ZN(G1332GAT) );
  XOR2_X1 U570 ( .A(G64GAT), .B(KEYINPUT103), .Z(n506) );
  NAND2_X1 U571 ( .A1(n509), .A2(n517), .ZN(n505) );
  XNOR2_X1 U572 ( .A(n506), .B(n505), .ZN(G1333GAT) );
  NAND2_X1 U573 ( .A1(n519), .A2(n509), .ZN(n507) );
  XNOR2_X1 U574 ( .A(n507), .B(KEYINPUT104), .ZN(n508) );
  XNOR2_X1 U575 ( .A(G71GAT), .B(n508), .ZN(G1334GAT) );
  XOR2_X1 U576 ( .A(G78GAT), .B(KEYINPUT43), .Z(n511) );
  NAND2_X1 U577 ( .A1(n509), .A2(n521), .ZN(n510) );
  XNOR2_X1 U578 ( .A(n511), .B(n510), .ZN(G1335GAT) );
  XOR2_X1 U579 ( .A(G85GAT), .B(KEYINPUT105), .Z(n516) );
  NOR2_X1 U580 ( .A1(n513), .A2(n512), .ZN(n522) );
  NAND2_X1 U581 ( .A1(n522), .A2(n514), .ZN(n515) );
  XNOR2_X1 U582 ( .A(n516), .B(n515), .ZN(G1336GAT) );
  NAND2_X1 U583 ( .A1(n517), .A2(n522), .ZN(n518) );
  XNOR2_X1 U584 ( .A(n518), .B(G92GAT), .ZN(G1337GAT) );
  NAND2_X1 U585 ( .A1(n519), .A2(n522), .ZN(n520) );
  XNOR2_X1 U586 ( .A(n520), .B(G99GAT), .ZN(G1338GAT) );
  XOR2_X1 U587 ( .A(KEYINPUT106), .B(KEYINPUT44), .Z(n524) );
  NAND2_X1 U588 ( .A1(n522), .A2(n521), .ZN(n523) );
  XNOR2_X1 U589 ( .A(n524), .B(n523), .ZN(n525) );
  XOR2_X1 U590 ( .A(G106GAT), .B(n525), .Z(G1339GAT) );
  NOR2_X1 U591 ( .A1(n527), .A2(n526), .ZN(n544) );
  NAND2_X1 U592 ( .A1(n544), .A2(n528), .ZN(n529) );
  NOR2_X1 U593 ( .A1(n530), .A2(n529), .ZN(n539) );
  NAND2_X1 U594 ( .A1(n557), .A2(n539), .ZN(n531) );
  XNOR2_X1 U595 ( .A(n531), .B(KEYINPUT110), .ZN(n532) );
  XNOR2_X1 U596 ( .A(G113GAT), .B(n532), .ZN(G1340GAT) );
  XOR2_X1 U597 ( .A(KEYINPUT112), .B(KEYINPUT49), .Z(n534) );
  NAND2_X1 U598 ( .A1(n539), .A2(n548), .ZN(n533) );
  XNOR2_X1 U599 ( .A(n534), .B(n533), .ZN(n536) );
  XOR2_X1 U600 ( .A(G120GAT), .B(KEYINPUT111), .Z(n535) );
  XNOR2_X1 U601 ( .A(n536), .B(n535), .ZN(G1341GAT) );
  NAND2_X1 U602 ( .A1(n572), .A2(n539), .ZN(n537) );
  XNOR2_X1 U603 ( .A(n537), .B(KEYINPUT50), .ZN(n538) );
  XNOR2_X1 U604 ( .A(G127GAT), .B(n538), .ZN(G1342GAT) );
  XOR2_X1 U605 ( .A(KEYINPUT114), .B(KEYINPUT51), .Z(n541) );
  NAND2_X1 U606 ( .A1(n539), .A2(n553), .ZN(n540) );
  XNOR2_X1 U607 ( .A(n541), .B(n540), .ZN(n543) );
  XOR2_X1 U608 ( .A(G134GAT), .B(KEYINPUT113), .Z(n542) );
  XNOR2_X1 U609 ( .A(n543), .B(n542), .ZN(G1343GAT) );
  XNOR2_X1 U610 ( .A(G141GAT), .B(KEYINPUT116), .ZN(n547) );
  NAND2_X1 U611 ( .A1(n560), .A2(n544), .ZN(n545) );
  XNOR2_X1 U612 ( .A(n545), .B(KEYINPUT115), .ZN(n554) );
  NAND2_X1 U613 ( .A1(n562), .A2(n554), .ZN(n546) );
  XNOR2_X1 U614 ( .A(n547), .B(n546), .ZN(G1344GAT) );
  XOR2_X1 U615 ( .A(KEYINPUT53), .B(KEYINPUT52), .Z(n550) );
  NAND2_X1 U616 ( .A1(n554), .A2(n548), .ZN(n549) );
  XNOR2_X1 U617 ( .A(n550), .B(n549), .ZN(n551) );
  XNOR2_X1 U618 ( .A(G148GAT), .B(n551), .ZN(G1345GAT) );
  NAND2_X1 U619 ( .A1(n572), .A2(n554), .ZN(n552) );
  XNOR2_X1 U620 ( .A(n552), .B(G155GAT), .ZN(G1346GAT) );
  XOR2_X1 U621 ( .A(G162GAT), .B(KEYINPUT117), .Z(n556) );
  NAND2_X1 U622 ( .A1(n554), .A2(n553), .ZN(n555) );
  XNOR2_X1 U623 ( .A(n556), .B(n555), .ZN(G1347GAT) );
  NAND2_X1 U624 ( .A1(n558), .A2(n557), .ZN(n559) );
  XNOR2_X1 U625 ( .A(G169GAT), .B(n559), .ZN(G1348GAT) );
  NAND2_X1 U626 ( .A1(n561), .A2(n560), .ZN(n576) );
  INV_X1 U627 ( .A(n576), .ZN(n571) );
  NAND2_X1 U628 ( .A1(n571), .A2(n562), .ZN(n566) );
  XOR2_X1 U629 ( .A(KEYINPUT124), .B(KEYINPUT59), .Z(n564) );
  XNOR2_X1 U630 ( .A(G197GAT), .B(KEYINPUT60), .ZN(n563) );
  XNOR2_X1 U631 ( .A(n564), .B(n563), .ZN(n565) );
  XNOR2_X1 U632 ( .A(n566), .B(n565), .ZN(G1352GAT) );
  XOR2_X1 U633 ( .A(KEYINPUT125), .B(KEYINPUT61), .Z(n569) );
  NAND2_X1 U634 ( .A1(n571), .A2(n567), .ZN(n568) );
  XNOR2_X1 U635 ( .A(n569), .B(n568), .ZN(n570) );
  XOR2_X1 U636 ( .A(G204GAT), .B(n570), .Z(G1353GAT) );
  NAND2_X1 U637 ( .A1(n572), .A2(n571), .ZN(n573) );
  XNOR2_X1 U638 ( .A(n573), .B(G211GAT), .ZN(G1354GAT) );
  XOR2_X1 U639 ( .A(KEYINPUT62), .B(KEYINPUT126), .Z(n575) );
  XNOR2_X1 U640 ( .A(G218GAT), .B(KEYINPUT127), .ZN(n574) );
  XNOR2_X1 U641 ( .A(n575), .B(n574), .ZN(n579) );
  NOR2_X1 U642 ( .A1(n577), .A2(n576), .ZN(n578) );
  XOR2_X1 U643 ( .A(n579), .B(n578), .Z(G1355GAT) );
endmodule

