//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 0 0 0 0 1 0 1 1 0 0 1 0 1 1 1 0 0 1 0 0 0 0 0 1 0 1 0 0 0 0 0 0 1 0 0 1 0 0 1 1 0 0 0 0 0 1 1 1 1 0 1 1 0 1 1 0 0 1 0 1 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:22:53 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n722, new_n723, new_n724,
    new_n725, new_n726, new_n727, new_n728, new_n729, new_n730, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n739, new_n741,
    new_n742, new_n743, new_n745, new_n746, new_n747, new_n748, new_n749,
    new_n750, new_n751, new_n752, new_n753, new_n754, new_n755, new_n756,
    new_n757, new_n758, new_n759, new_n760, new_n761, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n770, new_n771,
    new_n772, new_n773, new_n774, new_n775, new_n776, new_n777, new_n778,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n793, new_n794,
    new_n795, new_n796, new_n797, new_n798, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n825, new_n826, new_n827, new_n828, new_n829, new_n830, new_n831,
    new_n832, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n915, new_n916, new_n917,
    new_n918, new_n919, new_n920, new_n921, new_n922, new_n923, new_n924,
    new_n925, new_n926, new_n927, new_n928, new_n929, new_n930, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n944, new_n945, new_n946, new_n947,
    new_n949, new_n950, new_n951, new_n952, new_n954, new_n955, new_n956,
    new_n957, new_n958, new_n959, new_n960, new_n961, new_n962, new_n963,
    new_n964, new_n965, new_n966, new_n967, new_n968, new_n969, new_n970,
    new_n972, new_n973, new_n974, new_n975, new_n976, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011;
  INV_X1    g000(.A(G902), .ZN(new_n187));
  INV_X1    g001(.A(G146), .ZN(new_n188));
  AND2_X1   g002(.A1(KEYINPUT64), .A2(G143), .ZN(new_n189));
  NOR2_X1   g003(.A1(KEYINPUT64), .A2(G143), .ZN(new_n190));
  OAI21_X1  g004(.A(new_n188), .B1(new_n189), .B2(new_n190), .ZN(new_n191));
  INV_X1    g005(.A(G143), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n192), .A2(G146), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n191), .A2(new_n193), .ZN(new_n194));
  AND2_X1   g008(.A1(KEYINPUT0), .A2(G128), .ZN(new_n195));
  NOR2_X1   g009(.A1(KEYINPUT0), .A2(G128), .ZN(new_n196));
  NOR2_X1   g010(.A1(new_n195), .A2(new_n196), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n194), .A2(new_n197), .ZN(new_n198));
  INV_X1    g012(.A(KEYINPUT11), .ZN(new_n199));
  INV_X1    g013(.A(G134), .ZN(new_n200));
  OAI21_X1  g014(.A(new_n199), .B1(new_n200), .B2(G137), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n200), .A2(G137), .ZN(new_n202));
  INV_X1    g016(.A(G137), .ZN(new_n203));
  NAND3_X1  g017(.A1(new_n203), .A2(KEYINPUT11), .A3(G134), .ZN(new_n204));
  NAND3_X1  g018(.A1(new_n201), .A2(new_n202), .A3(new_n204), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n205), .A2(G131), .ZN(new_n206));
  INV_X1    g020(.A(G131), .ZN(new_n207));
  NAND4_X1  g021(.A1(new_n201), .A2(new_n204), .A3(new_n207), .A4(new_n202), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n206), .A2(new_n208), .ZN(new_n209));
  INV_X1    g023(.A(KEYINPUT65), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n188), .A2(G143), .ZN(new_n211));
  INV_X1    g025(.A(new_n211), .ZN(new_n212));
  NOR2_X1   g026(.A1(new_n189), .A2(new_n190), .ZN(new_n213));
  AOI21_X1  g027(.A(new_n212), .B1(new_n213), .B2(G146), .ZN(new_n214));
  AOI21_X1  g028(.A(new_n210), .B1(new_n214), .B2(new_n195), .ZN(new_n215));
  XNOR2_X1  g029(.A(KEYINPUT64), .B(G143), .ZN(new_n216));
  OAI211_X1 g030(.A(new_n211), .B(new_n195), .C1(new_n216), .C2(new_n188), .ZN(new_n217));
  NOR2_X1   g031(.A1(new_n217), .A2(KEYINPUT65), .ZN(new_n218));
  OAI211_X1 g032(.A(new_n198), .B(new_n209), .C1(new_n215), .C2(new_n218), .ZN(new_n219));
  OAI21_X1  g033(.A(new_n211), .B1(new_n216), .B2(new_n188), .ZN(new_n220));
  INV_X1    g034(.A(G128), .ZN(new_n221));
  NOR3_X1   g035(.A1(new_n220), .A2(KEYINPUT1), .A3(new_n221), .ZN(new_n222));
  OAI21_X1  g036(.A(KEYINPUT1), .B1(new_n192), .B2(G146), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n223), .A2(KEYINPUT66), .ZN(new_n224));
  INV_X1    g038(.A(KEYINPUT66), .ZN(new_n225));
  NAND3_X1  g039(.A1(new_n211), .A2(new_n225), .A3(KEYINPUT1), .ZN(new_n226));
  NAND3_X1  g040(.A1(new_n224), .A2(G128), .A3(new_n226), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n227), .A2(new_n194), .ZN(new_n228));
  INV_X1    g042(.A(KEYINPUT67), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n228), .A2(new_n229), .ZN(new_n230));
  NAND3_X1  g044(.A1(new_n227), .A2(KEYINPUT67), .A3(new_n194), .ZN(new_n231));
  AOI21_X1  g045(.A(new_n222), .B1(new_n230), .B2(new_n231), .ZN(new_n232));
  INV_X1    g046(.A(new_n202), .ZN(new_n233));
  NOR2_X1   g047(.A1(new_n200), .A2(G137), .ZN(new_n234));
  OAI21_X1  g048(.A(G131), .B1(new_n233), .B2(new_n234), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n235), .A2(new_n208), .ZN(new_n236));
  OAI21_X1  g050(.A(new_n219), .B1(new_n232), .B2(new_n236), .ZN(new_n237));
  INV_X1    g051(.A(G119), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n238), .A2(G116), .ZN(new_n239));
  INV_X1    g053(.A(G116), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n240), .A2(G119), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n239), .A2(new_n241), .ZN(new_n242));
  XNOR2_X1  g056(.A(KEYINPUT2), .B(G113), .ZN(new_n243));
  XNOR2_X1  g057(.A(new_n242), .B(new_n243), .ZN(new_n244));
  NOR2_X1   g058(.A1(new_n237), .A2(new_n244), .ZN(new_n245));
  INV_X1    g059(.A(new_n244), .ZN(new_n246));
  INV_X1    g060(.A(KEYINPUT1), .ZN(new_n247));
  NAND3_X1  g061(.A1(new_n214), .A2(new_n247), .A3(G128), .ZN(new_n248));
  AND3_X1   g062(.A1(new_n227), .A2(KEYINPUT67), .A3(new_n194), .ZN(new_n249));
  AOI21_X1  g063(.A(KEYINPUT67), .B1(new_n227), .B2(new_n194), .ZN(new_n250));
  OAI21_X1  g064(.A(new_n248), .B1(new_n249), .B2(new_n250), .ZN(new_n251));
  INV_X1    g065(.A(new_n236), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n251), .A2(new_n252), .ZN(new_n253));
  AOI21_X1  g067(.A(new_n246), .B1(new_n253), .B2(new_n219), .ZN(new_n254));
  OAI21_X1  g068(.A(KEYINPUT28), .B1(new_n245), .B2(new_n254), .ZN(new_n255));
  INV_X1    g069(.A(KEYINPUT72), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n255), .A2(new_n256), .ZN(new_n257));
  XNOR2_X1  g071(.A(KEYINPUT69), .B(G953), .ZN(new_n258));
  INV_X1    g072(.A(G237), .ZN(new_n259));
  NAND3_X1  g073(.A1(new_n258), .A2(G210), .A3(new_n259), .ZN(new_n260));
  XOR2_X1   g074(.A(KEYINPUT26), .B(G101), .Z(new_n261));
  XNOR2_X1  g075(.A(new_n260), .B(new_n261), .ZN(new_n262));
  XNOR2_X1  g076(.A(KEYINPUT70), .B(KEYINPUT27), .ZN(new_n263));
  XNOR2_X1  g077(.A(new_n262), .B(new_n263), .ZN(new_n264));
  INV_X1    g078(.A(KEYINPUT29), .ZN(new_n265));
  NOR2_X1   g079(.A1(new_n264), .A2(new_n265), .ZN(new_n266));
  INV_X1    g080(.A(KEYINPUT28), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n237), .A2(new_n244), .ZN(new_n268));
  NAND3_X1  g082(.A1(new_n253), .A2(new_n246), .A3(new_n219), .ZN(new_n269));
  AOI21_X1  g083(.A(new_n267), .B1(new_n268), .B2(new_n269), .ZN(new_n270));
  AND2_X1   g084(.A1(new_n269), .A2(new_n267), .ZN(new_n271));
  NOR2_X1   g085(.A1(new_n270), .A2(new_n271), .ZN(new_n272));
  OAI211_X1 g086(.A(new_n257), .B(new_n266), .C1(new_n272), .C2(new_n256), .ZN(new_n273));
  NOR3_X1   g087(.A1(new_n270), .A2(new_n271), .A3(new_n264), .ZN(new_n274));
  INV_X1    g088(.A(KEYINPUT71), .ZN(new_n275));
  OAI21_X1  g089(.A(new_n265), .B1(new_n274), .B2(new_n275), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n269), .A2(new_n267), .ZN(new_n277));
  INV_X1    g091(.A(new_n264), .ZN(new_n278));
  NAND4_X1  g092(.A1(new_n255), .A2(new_n275), .A3(new_n277), .A4(new_n278), .ZN(new_n279));
  INV_X1    g093(.A(KEYINPUT68), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n230), .A2(new_n231), .ZN(new_n281));
  AOI21_X1  g095(.A(new_n236), .B1(new_n281), .B2(new_n248), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n219), .A2(KEYINPUT30), .ZN(new_n283));
  OAI21_X1  g097(.A(new_n244), .B1(new_n282), .B2(new_n283), .ZN(new_n284));
  AOI21_X1  g098(.A(KEYINPUT30), .B1(new_n253), .B2(new_n219), .ZN(new_n285));
  OAI21_X1  g099(.A(new_n280), .B1(new_n284), .B2(new_n285), .ZN(new_n286));
  INV_X1    g100(.A(KEYINPUT30), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n237), .A2(new_n287), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n217), .A2(KEYINPUT65), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n213), .A2(G146), .ZN(new_n290));
  NAND4_X1  g104(.A1(new_n290), .A2(new_n210), .A3(new_n211), .A4(new_n195), .ZN(new_n291));
  AOI22_X1  g105(.A1(new_n289), .A2(new_n291), .B1(new_n194), .B2(new_n197), .ZN(new_n292));
  AOI21_X1  g106(.A(new_n287), .B1(new_n292), .B2(new_n209), .ZN(new_n293));
  AOI21_X1  g107(.A(new_n246), .B1(new_n253), .B2(new_n293), .ZN(new_n294));
  NAND3_X1  g108(.A1(new_n288), .A2(new_n294), .A3(KEYINPUT68), .ZN(new_n295));
  AOI21_X1  g109(.A(new_n245), .B1(new_n286), .B2(new_n295), .ZN(new_n296));
  OAI21_X1  g110(.A(new_n279), .B1(new_n296), .B2(new_n278), .ZN(new_n297));
  OAI211_X1 g111(.A(new_n187), .B(new_n273), .C1(new_n276), .C2(new_n297), .ZN(new_n298));
  NAND2_X1  g112(.A1(new_n298), .A2(G472), .ZN(new_n299));
  OAI21_X1  g113(.A(new_n264), .B1(new_n270), .B2(new_n271), .ZN(new_n300));
  NAND2_X1  g114(.A1(new_n286), .A2(new_n295), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n269), .A2(new_n278), .ZN(new_n302));
  INV_X1    g116(.A(new_n302), .ZN(new_n303));
  AOI21_X1  g117(.A(KEYINPUT31), .B1(new_n301), .B2(new_n303), .ZN(new_n304));
  INV_X1    g118(.A(KEYINPUT31), .ZN(new_n305));
  AOI211_X1 g119(.A(new_n305), .B(new_n302), .C1(new_n286), .C2(new_n295), .ZN(new_n306));
  OAI21_X1  g120(.A(new_n300), .B1(new_n304), .B2(new_n306), .ZN(new_n307));
  INV_X1    g121(.A(KEYINPUT32), .ZN(new_n308));
  NOR2_X1   g122(.A1(G472), .A2(G902), .ZN(new_n309));
  AND3_X1   g123(.A1(new_n307), .A2(new_n308), .A3(new_n309), .ZN(new_n310));
  AOI21_X1  g124(.A(new_n308), .B1(new_n307), .B2(new_n309), .ZN(new_n311));
  OAI21_X1  g125(.A(new_n299), .B1(new_n310), .B2(new_n311), .ZN(new_n312));
  INV_X1    g126(.A(G217), .ZN(new_n313));
  AOI21_X1  g127(.A(new_n313), .B1(G234), .B2(new_n187), .ZN(new_n314));
  INV_X1    g128(.A(new_n314), .ZN(new_n315));
  INV_X1    g129(.A(KEYINPUT75), .ZN(new_n316));
  INV_X1    g130(.A(KEYINPUT25), .ZN(new_n317));
  INV_X1    g131(.A(G125), .ZN(new_n318));
  NOR2_X1   g132(.A1(new_n318), .A2(G140), .ZN(new_n319));
  XNOR2_X1  g133(.A(G125), .B(G140), .ZN(new_n320));
  MUX2_X1   g134(.A(new_n319), .B(new_n320), .S(KEYINPUT16), .Z(new_n321));
  NOR2_X1   g135(.A1(new_n321), .A2(new_n188), .ZN(new_n322));
  AOI21_X1  g136(.A(new_n322), .B1(new_n188), .B2(new_n320), .ZN(new_n323));
  OAI21_X1  g137(.A(KEYINPUT23), .B1(new_n221), .B2(G119), .ZN(new_n324));
  OAI21_X1  g138(.A(KEYINPUT73), .B1(new_n238), .B2(G128), .ZN(new_n325));
  XOR2_X1   g139(.A(new_n324), .B(new_n325), .Z(new_n326));
  XNOR2_X1  g140(.A(G119), .B(G128), .ZN(new_n327));
  XNOR2_X1  g141(.A(KEYINPUT24), .B(G110), .ZN(new_n328));
  INV_X1    g142(.A(new_n328), .ZN(new_n329));
  OAI22_X1  g143(.A1(new_n326), .A2(G110), .B1(new_n327), .B2(new_n329), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n323), .A2(new_n330), .ZN(new_n331));
  AOI22_X1  g145(.A1(new_n326), .A2(G110), .B1(new_n327), .B2(new_n329), .ZN(new_n332));
  AND2_X1   g146(.A1(new_n321), .A2(new_n188), .ZN(new_n333));
  OAI21_X1  g147(.A(new_n332), .B1(new_n333), .B2(new_n322), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n331), .A2(new_n334), .ZN(new_n335));
  INV_X1    g149(.A(new_n335), .ZN(new_n336));
  NAND3_X1  g150(.A1(new_n258), .A2(G221), .A3(G234), .ZN(new_n337));
  XNOR2_X1  g151(.A(KEYINPUT22), .B(G137), .ZN(new_n338));
  XNOR2_X1  g152(.A(new_n337), .B(new_n338), .ZN(new_n339));
  XOR2_X1   g153(.A(new_n339), .B(KEYINPUT74), .Z(new_n340));
  OR2_X1    g154(.A1(new_n336), .A2(new_n340), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n336), .A2(new_n339), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n341), .A2(new_n342), .ZN(new_n343));
  OAI211_X1 g157(.A(new_n316), .B(new_n317), .C1(new_n343), .C2(G902), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n316), .A2(new_n317), .ZN(new_n345));
  NAND4_X1  g159(.A1(new_n341), .A2(new_n187), .A3(new_n342), .A4(new_n345), .ZN(new_n346));
  AOI21_X1  g160(.A(new_n315), .B1(new_n344), .B2(new_n346), .ZN(new_n347));
  NOR3_X1   g161(.A1(new_n343), .A2(G902), .A3(new_n314), .ZN(new_n348));
  NOR2_X1   g162(.A1(new_n347), .A2(new_n348), .ZN(new_n349));
  XNOR2_X1  g163(.A(KEYINPUT9), .B(G234), .ZN(new_n350));
  OAI21_X1  g164(.A(G221), .B1(new_n350), .B2(G902), .ZN(new_n351));
  INV_X1    g165(.A(new_n351), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n258), .A2(G227), .ZN(new_n353));
  XOR2_X1   g167(.A(G110), .B(G140), .Z(new_n354));
  XNOR2_X1  g168(.A(new_n353), .B(new_n354), .ZN(new_n355));
  INV_X1    g169(.A(KEYINPUT3), .ZN(new_n356));
  INV_X1    g170(.A(G104), .ZN(new_n357));
  OAI21_X1  g171(.A(new_n356), .B1(new_n357), .B2(G107), .ZN(new_n358));
  INV_X1    g172(.A(G107), .ZN(new_n359));
  NAND3_X1  g173(.A1(new_n359), .A2(KEYINPUT3), .A3(G104), .ZN(new_n360));
  AND2_X1   g174(.A1(new_n358), .A2(new_n360), .ZN(new_n361));
  INV_X1    g175(.A(KEYINPUT76), .ZN(new_n362));
  OAI21_X1  g176(.A(new_n362), .B1(new_n359), .B2(G104), .ZN(new_n363));
  NAND3_X1  g177(.A1(new_n357), .A2(KEYINPUT76), .A3(G107), .ZN(new_n364));
  NAND2_X1  g178(.A1(new_n363), .A2(new_n364), .ZN(new_n365));
  OAI21_X1  g179(.A(G101), .B1(new_n361), .B2(new_n365), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n366), .A2(KEYINPUT4), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n358), .A2(new_n360), .ZN(new_n368));
  INV_X1    g182(.A(G101), .ZN(new_n369));
  NAND4_X1  g183(.A1(new_n368), .A2(new_n369), .A3(new_n363), .A4(new_n364), .ZN(new_n370));
  INV_X1    g184(.A(KEYINPUT77), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n370), .A2(new_n371), .ZN(new_n372));
  INV_X1    g186(.A(new_n365), .ZN(new_n373));
  NAND4_X1  g187(.A1(new_n373), .A2(KEYINPUT77), .A3(new_n369), .A4(new_n368), .ZN(new_n374));
  AOI21_X1  g188(.A(new_n367), .B1(new_n372), .B2(new_n374), .ZN(new_n375));
  NAND3_X1  g189(.A1(new_n368), .A2(new_n363), .A3(new_n364), .ZN(new_n376));
  INV_X1    g190(.A(KEYINPUT4), .ZN(new_n377));
  NAND3_X1  g191(.A1(new_n376), .A2(new_n377), .A3(G101), .ZN(new_n378));
  OAI211_X1 g192(.A(new_n198), .B(new_n378), .C1(new_n215), .C2(new_n218), .ZN(new_n379));
  OAI21_X1  g193(.A(KEYINPUT78), .B1(new_n375), .B2(new_n379), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n372), .A2(new_n374), .ZN(new_n381));
  AOI21_X1  g195(.A(new_n377), .B1(new_n376), .B2(G101), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n381), .A2(new_n382), .ZN(new_n383));
  INV_X1    g197(.A(KEYINPUT78), .ZN(new_n384));
  NAND4_X1  g198(.A1(new_n383), .A2(new_n384), .A3(new_n292), .A4(new_n378), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n380), .A2(new_n385), .ZN(new_n386));
  INV_X1    g200(.A(new_n209), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n359), .A2(G104), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n357), .A2(G107), .ZN(new_n389));
  AOI21_X1  g203(.A(new_n369), .B1(new_n388), .B2(new_n389), .ZN(new_n390));
  AOI21_X1  g204(.A(new_n390), .B1(new_n372), .B2(new_n374), .ZN(new_n391));
  INV_X1    g205(.A(KEYINPUT79), .ZN(new_n392));
  AOI21_X1  g206(.A(new_n221), .B1(new_n191), .B2(KEYINPUT1), .ZN(new_n393));
  OAI21_X1  g207(.A(new_n392), .B1(new_n393), .B2(new_n214), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n394), .A2(new_n248), .ZN(new_n395));
  NOR3_X1   g209(.A1(new_n393), .A2(new_n214), .A3(new_n392), .ZN(new_n396));
  OAI21_X1  g210(.A(new_n391), .B1(new_n395), .B2(new_n396), .ZN(new_n397));
  INV_X1    g211(.A(KEYINPUT10), .ZN(new_n398));
  AOI211_X1 g212(.A(new_n398), .B(new_n390), .C1(new_n372), .C2(new_n374), .ZN(new_n399));
  AOI22_X1  g213(.A1(new_n397), .A2(new_n398), .B1(new_n399), .B2(new_n251), .ZN(new_n400));
  AND3_X1   g214(.A1(new_n386), .A2(new_n387), .A3(new_n400), .ZN(new_n401));
  AOI21_X1  g215(.A(new_n387), .B1(new_n386), .B2(new_n400), .ZN(new_n402));
  OAI21_X1  g216(.A(new_n355), .B1(new_n401), .B2(new_n402), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n403), .A2(KEYINPUT81), .ZN(new_n404));
  INV_X1    g218(.A(KEYINPUT81), .ZN(new_n405));
  OAI211_X1 g219(.A(new_n405), .B(new_n355), .C1(new_n401), .C2(new_n402), .ZN(new_n406));
  NAND3_X1  g220(.A1(new_n386), .A2(new_n387), .A3(new_n400), .ZN(new_n407));
  INV_X1    g221(.A(new_n355), .ZN(new_n408));
  AND2_X1   g222(.A1(new_n407), .A2(new_n408), .ZN(new_n409));
  INV_X1    g223(.A(new_n390), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n381), .A2(new_n410), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n232), .A2(new_n411), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n412), .A2(new_n397), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n413), .A2(new_n209), .ZN(new_n414));
  INV_X1    g228(.A(KEYINPUT12), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n414), .A2(new_n415), .ZN(new_n416));
  NAND3_X1  g230(.A1(new_n413), .A2(KEYINPUT12), .A3(new_n209), .ZN(new_n417));
  NAND3_X1  g231(.A1(new_n416), .A2(KEYINPUT80), .A3(new_n417), .ZN(new_n418));
  INV_X1    g232(.A(KEYINPUT80), .ZN(new_n419));
  AOI21_X1  g233(.A(KEYINPUT12), .B1(new_n413), .B2(new_n209), .ZN(new_n420));
  AOI211_X1 g234(.A(new_n415), .B(new_n387), .C1(new_n412), .C2(new_n397), .ZN(new_n421));
  OAI21_X1  g235(.A(new_n419), .B1(new_n420), .B2(new_n421), .ZN(new_n422));
  NAND3_X1  g236(.A1(new_n409), .A2(new_n418), .A3(new_n422), .ZN(new_n423));
  NAND3_X1  g237(.A1(new_n404), .A2(new_n406), .A3(new_n423), .ZN(new_n424));
  INV_X1    g238(.A(G469), .ZN(new_n425));
  NAND3_X1  g239(.A1(new_n424), .A2(new_n425), .A3(new_n187), .ZN(new_n426));
  NOR2_X1   g240(.A1(new_n425), .A2(new_n187), .ZN(new_n427));
  INV_X1    g241(.A(new_n402), .ZN(new_n428));
  OAI21_X1  g242(.A(new_n407), .B1(new_n420), .B2(new_n421), .ZN(new_n429));
  AOI22_X1  g243(.A1(new_n428), .A2(new_n409), .B1(new_n429), .B2(new_n355), .ZN(new_n430));
  AOI21_X1  g244(.A(new_n427), .B1(new_n430), .B2(G469), .ZN(new_n431));
  AOI21_X1  g245(.A(new_n352), .B1(new_n426), .B2(new_n431), .ZN(new_n432));
  NAND3_X1  g246(.A1(new_n312), .A2(new_n349), .A3(new_n432), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n240), .A2(G122), .ZN(new_n434));
  INV_X1    g248(.A(G122), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n435), .A2(G116), .ZN(new_n436));
  NAND2_X1  g250(.A1(new_n434), .A2(new_n436), .ZN(new_n437));
  NOR2_X1   g251(.A1(new_n437), .A2(KEYINPUT95), .ZN(new_n438));
  INV_X1    g252(.A(KEYINPUT95), .ZN(new_n439));
  AOI21_X1  g253(.A(new_n439), .B1(new_n434), .B2(new_n436), .ZN(new_n440));
  OAI21_X1  g254(.A(new_n359), .B1(new_n438), .B2(new_n440), .ZN(new_n441));
  INV_X1    g255(.A(KEYINPUT14), .ZN(new_n442));
  NOR2_X1   g256(.A1(new_n434), .A2(new_n442), .ZN(new_n443));
  NOR2_X1   g257(.A1(new_n443), .A2(new_n359), .ZN(new_n444));
  XNOR2_X1  g258(.A(G116), .B(G122), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n445), .A2(new_n442), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n444), .A2(new_n446), .ZN(new_n447));
  INV_X1    g261(.A(KEYINPUT96), .ZN(new_n448));
  OAI21_X1  g262(.A(new_n448), .B1(new_n192), .B2(G128), .ZN(new_n449));
  NAND3_X1  g263(.A1(new_n221), .A2(KEYINPUT96), .A3(G143), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n449), .A2(new_n450), .ZN(new_n451));
  OR2_X1    g265(.A1(KEYINPUT64), .A2(G143), .ZN(new_n452));
  NAND2_X1  g266(.A1(KEYINPUT64), .A2(G143), .ZN(new_n453));
  NAND3_X1  g267(.A1(new_n452), .A2(G128), .A3(new_n453), .ZN(new_n454));
  NAND3_X1  g268(.A1(new_n451), .A2(new_n454), .A3(new_n200), .ZN(new_n455));
  INV_X1    g269(.A(new_n455), .ZN(new_n456));
  AOI21_X1  g270(.A(new_n200), .B1(new_n451), .B2(new_n454), .ZN(new_n457));
  OAI211_X1 g271(.A(new_n441), .B(new_n447), .C1(new_n456), .C2(new_n457), .ZN(new_n458));
  INV_X1    g272(.A(KEYINPUT97), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  INV_X1    g274(.A(new_n440), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n445), .A2(new_n439), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  AOI22_X1  g277(.A1(new_n463), .A2(new_n359), .B1(new_n446), .B2(new_n444), .ZN(new_n464));
  INV_X1    g278(.A(new_n457), .ZN(new_n465));
  NAND2_X1  g279(.A1(new_n465), .A2(new_n455), .ZN(new_n466));
  NAND3_X1  g280(.A1(new_n464), .A2(new_n466), .A3(KEYINPUT97), .ZN(new_n467));
  NAND2_X1  g281(.A1(new_n460), .A2(new_n467), .ZN(new_n468));
  NAND3_X1  g282(.A1(new_n461), .A2(new_n462), .A3(G107), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n441), .A2(new_n469), .ZN(new_n470));
  INV_X1    g284(.A(KEYINPUT13), .ZN(new_n471));
  OAI21_X1  g285(.A(new_n451), .B1(new_n454), .B2(new_n471), .ZN(new_n472));
  AOI21_X1  g286(.A(KEYINPUT13), .B1(new_n213), .B2(G128), .ZN(new_n473));
  OAI21_X1  g287(.A(G134), .B1(new_n472), .B2(new_n473), .ZN(new_n474));
  NAND3_X1  g288(.A1(new_n470), .A2(new_n455), .A3(new_n474), .ZN(new_n475));
  NOR3_X1   g289(.A1(new_n350), .A2(new_n313), .A3(G953), .ZN(new_n476));
  AND3_X1   g290(.A1(new_n468), .A2(new_n475), .A3(new_n476), .ZN(new_n477));
  AOI21_X1  g291(.A(new_n476), .B1(new_n468), .B2(new_n475), .ZN(new_n478));
  OAI21_X1  g292(.A(new_n187), .B1(new_n477), .B2(new_n478), .ZN(new_n479));
  INV_X1    g293(.A(G478), .ZN(new_n480));
  NOR2_X1   g294(.A1(new_n480), .A2(KEYINPUT15), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n479), .A2(new_n481), .ZN(new_n482));
  OAI221_X1 g296(.A(new_n187), .B1(KEYINPUT15), .B2(new_n480), .C1(new_n477), .C2(new_n478), .ZN(new_n483));
  AOI21_X1  g297(.A(KEYINPUT98), .B1(new_n482), .B2(new_n483), .ZN(new_n484));
  INV_X1    g298(.A(new_n484), .ZN(new_n485));
  NAND3_X1  g299(.A1(new_n482), .A2(new_n483), .A3(KEYINPUT98), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n485), .A2(new_n486), .ZN(new_n487));
  INV_X1    g301(.A(KEYINPUT17), .ZN(new_n488));
  INV_X1    g302(.A(G953), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n489), .A2(KEYINPUT69), .ZN(new_n490));
  INV_X1    g304(.A(KEYINPUT69), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n491), .A2(G953), .ZN(new_n492));
  NAND4_X1  g306(.A1(new_n490), .A2(new_n492), .A3(G214), .A4(new_n259), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n493), .A2(new_n213), .ZN(new_n494));
  NAND4_X1  g308(.A1(new_n258), .A2(G143), .A3(G214), .A4(new_n259), .ZN(new_n495));
  NAND3_X1  g309(.A1(new_n494), .A2(new_n495), .A3(new_n207), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n494), .A2(new_n495), .ZN(new_n497));
  AOI21_X1  g311(.A(KEYINPUT93), .B1(new_n497), .B2(G131), .ZN(new_n498));
  INV_X1    g312(.A(KEYINPUT93), .ZN(new_n499));
  AOI211_X1 g313(.A(new_n499), .B(new_n207), .C1(new_n494), .C2(new_n495), .ZN(new_n500));
  OAI211_X1 g314(.A(new_n488), .B(new_n496), .C1(new_n498), .C2(new_n500), .ZN(new_n501));
  NAND2_X1  g315(.A1(new_n497), .A2(G131), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n502), .A2(new_n499), .ZN(new_n503));
  NAND3_X1  g317(.A1(new_n497), .A2(KEYINPUT93), .A3(G131), .ZN(new_n504));
  NAND3_X1  g318(.A1(new_n503), .A2(KEYINPUT17), .A3(new_n504), .ZN(new_n505));
  NOR2_X1   g319(.A1(new_n333), .A2(new_n322), .ZN(new_n506));
  NAND3_X1  g320(.A1(new_n501), .A2(new_n505), .A3(new_n506), .ZN(new_n507));
  XNOR2_X1  g321(.A(G113), .B(G122), .ZN(new_n508));
  XNOR2_X1  g322(.A(new_n508), .B(new_n357), .ZN(new_n509));
  INV_X1    g323(.A(KEYINPUT92), .ZN(new_n510));
  INV_X1    g324(.A(KEYINPUT18), .ZN(new_n511));
  AOI211_X1 g325(.A(new_n511), .B(new_n207), .C1(new_n494), .C2(new_n495), .ZN(new_n512));
  NAND2_X1  g326(.A1(KEYINPUT18), .A2(G131), .ZN(new_n513));
  NAND3_X1  g327(.A1(new_n494), .A2(new_n495), .A3(new_n513), .ZN(new_n514));
  XNOR2_X1  g328(.A(new_n320), .B(new_n188), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  OAI21_X1  g330(.A(new_n510), .B1(new_n512), .B2(new_n516), .ZN(new_n517));
  NAND3_X1  g331(.A1(new_n497), .A2(KEYINPUT18), .A3(G131), .ZN(new_n518));
  NAND4_X1  g332(.A1(new_n518), .A2(KEYINPUT92), .A3(new_n514), .A4(new_n515), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n517), .A2(new_n519), .ZN(new_n520));
  AND3_X1   g334(.A1(new_n507), .A2(new_n509), .A3(new_n520), .ZN(new_n521));
  AOI21_X1  g335(.A(new_n509), .B1(new_n507), .B2(new_n520), .ZN(new_n522));
  OAI21_X1  g336(.A(new_n187), .B1(new_n521), .B2(new_n522), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n523), .A2(G475), .ZN(new_n524));
  INV_X1    g338(.A(KEYINPUT20), .ZN(new_n525));
  OAI21_X1  g339(.A(new_n496), .B1(new_n498), .B2(new_n500), .ZN(new_n526));
  XNOR2_X1  g340(.A(new_n320), .B(KEYINPUT19), .ZN(new_n527));
  AOI21_X1  g341(.A(new_n322), .B1(new_n188), .B2(new_n527), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n526), .A2(new_n528), .ZN(new_n529));
  NAND2_X1  g343(.A1(new_n529), .A2(new_n520), .ZN(new_n530));
  INV_X1    g344(.A(new_n509), .ZN(new_n531));
  NAND2_X1  g345(.A1(new_n530), .A2(new_n531), .ZN(new_n532));
  NAND3_X1  g346(.A1(new_n507), .A2(new_n509), .A3(new_n520), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  NOR2_X1   g348(.A1(G475), .A2(G902), .ZN(new_n535));
  XNOR2_X1  g349(.A(new_n535), .B(KEYINPUT94), .ZN(new_n536));
  INV_X1    g350(.A(new_n536), .ZN(new_n537));
  AOI21_X1  g351(.A(new_n525), .B1(new_n534), .B2(new_n537), .ZN(new_n538));
  AOI211_X1 g352(.A(KEYINPUT20), .B(new_n536), .C1(new_n532), .C2(new_n533), .ZN(new_n539));
  OAI21_X1  g353(.A(new_n524), .B1(new_n538), .B2(new_n539), .ZN(new_n540));
  INV_X1    g354(.A(new_n540), .ZN(new_n541));
  INV_X1    g355(.A(G952), .ZN(new_n542));
  AOI211_X1 g356(.A(G953), .B(new_n542), .C1(G234), .C2(G237), .ZN(new_n543));
  AOI211_X1 g357(.A(new_n187), .B(new_n258), .C1(G234), .C2(G237), .ZN(new_n544));
  XNOR2_X1  g358(.A(KEYINPUT21), .B(G898), .ZN(new_n545));
  AOI21_X1  g359(.A(new_n543), .B1(new_n544), .B2(new_n545), .ZN(new_n546));
  INV_X1    g360(.A(new_n546), .ZN(new_n547));
  AND3_X1   g361(.A1(new_n487), .A2(new_n541), .A3(new_n547), .ZN(new_n548));
  OAI21_X1  g362(.A(new_n198), .B1(new_n215), .B2(new_n218), .ZN(new_n549));
  INV_X1    g363(.A(KEYINPUT84), .ZN(new_n550));
  NAND3_X1  g364(.A1(new_n549), .A2(new_n550), .A3(G125), .ZN(new_n551));
  NAND3_X1  g365(.A1(new_n281), .A2(new_n318), .A3(new_n248), .ZN(new_n552));
  OAI21_X1  g366(.A(KEYINPUT84), .B1(new_n292), .B2(new_n318), .ZN(new_n553));
  NAND3_X1  g367(.A1(new_n551), .A2(new_n552), .A3(new_n553), .ZN(new_n554));
  XNOR2_X1  g368(.A(KEYINPUT86), .B(G224), .ZN(new_n555));
  OAI21_X1  g369(.A(KEYINPUT7), .B1(new_n555), .B2(G953), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n554), .A2(new_n556), .ZN(new_n557));
  XNOR2_X1  g371(.A(G110), .B(G122), .ZN(new_n558));
  XNOR2_X1  g372(.A(new_n558), .B(KEYINPUT8), .ZN(new_n559));
  NOR2_X1   g373(.A1(new_n242), .A2(new_n243), .ZN(new_n560));
  OAI21_X1  g374(.A(G113), .B1(new_n239), .B2(KEYINPUT5), .ZN(new_n561));
  NAND3_X1  g375(.A1(new_n239), .A2(new_n241), .A3(KEYINPUT5), .ZN(new_n562));
  AOI21_X1  g376(.A(new_n561), .B1(KEYINPUT88), .B2(new_n562), .ZN(new_n563));
  OR2_X1    g377(.A1(new_n562), .A2(KEYINPUT88), .ZN(new_n564));
  AOI21_X1  g378(.A(new_n560), .B1(new_n563), .B2(new_n564), .ZN(new_n565));
  NAND4_X1  g379(.A1(new_n381), .A2(new_n565), .A3(KEYINPUT89), .A4(new_n410), .ZN(new_n566));
  INV_X1    g380(.A(new_n562), .ZN(new_n567));
  OAI22_X1  g381(.A1(new_n567), .A2(new_n561), .B1(new_n242), .B2(new_n243), .ZN(new_n568));
  INV_X1    g382(.A(new_n568), .ZN(new_n569));
  OAI21_X1  g383(.A(new_n566), .B1(new_n391), .B2(new_n569), .ZN(new_n570));
  AOI21_X1  g384(.A(KEYINPUT89), .B1(new_n391), .B2(new_n565), .ZN(new_n571));
  OAI21_X1  g385(.A(new_n559), .B1(new_n570), .B2(new_n571), .ZN(new_n572));
  INV_X1    g386(.A(new_n556), .ZN(new_n573));
  NAND4_X1  g387(.A1(new_n552), .A2(new_n551), .A3(new_n553), .A4(new_n573), .ZN(new_n574));
  NAND3_X1  g388(.A1(new_n557), .A2(new_n572), .A3(new_n574), .ZN(new_n575));
  INV_X1    g389(.A(KEYINPUT90), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n575), .A2(new_n576), .ZN(new_n577));
  NAND2_X1  g391(.A1(new_n391), .A2(new_n569), .ZN(new_n578));
  NAND2_X1  g392(.A1(new_n378), .A2(new_n244), .ZN(new_n579));
  OAI21_X1  g393(.A(new_n578), .B1(new_n375), .B2(new_n579), .ZN(new_n580));
  INV_X1    g394(.A(new_n558), .ZN(new_n581));
  NOR2_X1   g395(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  INV_X1    g396(.A(new_n582), .ZN(new_n583));
  NAND4_X1  g397(.A1(new_n557), .A2(new_n572), .A3(KEYINPUT90), .A4(new_n574), .ZN(new_n584));
  NAND3_X1  g398(.A1(new_n577), .A2(new_n583), .A3(new_n584), .ZN(new_n585));
  AOI21_X1  g399(.A(new_n579), .B1(new_n381), .B2(new_n382), .ZN(new_n586));
  AOI211_X1 g400(.A(new_n390), .B(new_n568), .C1(new_n372), .C2(new_n374), .ZN(new_n587));
  OAI21_X1  g401(.A(KEYINPUT82), .B1(new_n586), .B2(new_n587), .ZN(new_n588));
  INV_X1    g402(.A(KEYINPUT82), .ZN(new_n589));
  OAI211_X1 g403(.A(new_n578), .B(new_n589), .C1(new_n375), .C2(new_n579), .ZN(new_n590));
  INV_X1    g404(.A(KEYINPUT6), .ZN(new_n591));
  NAND4_X1  g405(.A1(new_n588), .A2(new_n590), .A3(new_n591), .A4(new_n581), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n592), .A2(KEYINPUT83), .ZN(new_n593));
  AOI21_X1  g407(.A(new_n558), .B1(new_n580), .B2(KEYINPUT82), .ZN(new_n594));
  INV_X1    g408(.A(KEYINPUT83), .ZN(new_n595));
  NAND4_X1  g409(.A1(new_n594), .A2(new_n595), .A3(new_n591), .A4(new_n590), .ZN(new_n596));
  NAND2_X1  g410(.A1(new_n593), .A2(new_n596), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n594), .A2(new_n590), .ZN(new_n598));
  NOR2_X1   g412(.A1(new_n582), .A2(new_n591), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  NAND2_X1  g414(.A1(new_n597), .A2(new_n600), .ZN(new_n601));
  INV_X1    g415(.A(KEYINPUT85), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n554), .A2(new_n602), .ZN(new_n603));
  NAND4_X1  g417(.A1(new_n552), .A2(new_n551), .A3(new_n553), .A4(KEYINPUT85), .ZN(new_n604));
  NOR2_X1   g418(.A1(new_n555), .A2(G953), .ZN(new_n605));
  XNOR2_X1  g419(.A(new_n605), .B(KEYINPUT87), .ZN(new_n606));
  NAND3_X1  g420(.A1(new_n603), .A2(new_n604), .A3(new_n606), .ZN(new_n607));
  INV_X1    g421(.A(new_n607), .ZN(new_n608));
  AOI21_X1  g422(.A(new_n606), .B1(new_n603), .B2(new_n604), .ZN(new_n609));
  NOR2_X1   g423(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  OAI211_X1 g424(.A(new_n585), .B(new_n187), .C1(new_n601), .C2(new_n610), .ZN(new_n611));
  OAI21_X1  g425(.A(G210), .B1(G237), .B2(G902), .ZN(new_n612));
  INV_X1    g426(.A(new_n612), .ZN(new_n613));
  NAND2_X1  g427(.A1(new_n613), .A2(KEYINPUT91), .ZN(new_n614));
  INV_X1    g428(.A(new_n614), .ZN(new_n615));
  NAND2_X1  g429(.A1(new_n611), .A2(new_n615), .ZN(new_n616));
  AOI22_X1  g430(.A1(new_n593), .A2(new_n596), .B1(new_n598), .B2(new_n599), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n603), .A2(new_n604), .ZN(new_n618));
  INV_X1    g432(.A(new_n606), .ZN(new_n619));
  NAND2_X1  g433(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  NAND2_X1  g434(.A1(new_n620), .A2(new_n607), .ZN(new_n621));
  AOI21_X1  g435(.A(G902), .B1(new_n617), .B2(new_n621), .ZN(new_n622));
  NAND3_X1  g436(.A1(new_n622), .A2(new_n614), .A3(new_n585), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n616), .A2(new_n623), .ZN(new_n624));
  OAI21_X1  g438(.A(G214), .B1(G237), .B2(G902), .ZN(new_n625));
  NAND3_X1  g439(.A1(new_n548), .A2(new_n624), .A3(new_n625), .ZN(new_n626));
  NOR2_X1   g440(.A1(new_n433), .A2(new_n626), .ZN(new_n627));
  XNOR2_X1  g441(.A(new_n627), .B(new_n369), .ZN(G3));
  INV_X1    g442(.A(new_n625), .ZN(new_n629));
  INV_X1    g443(.A(KEYINPUT99), .ZN(new_n630));
  NAND2_X1  g444(.A1(new_n612), .A2(new_n630), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n611), .A2(new_n631), .ZN(new_n632));
  XNOR2_X1  g446(.A(new_n612), .B(KEYINPUT99), .ZN(new_n633));
  INV_X1    g447(.A(new_n633), .ZN(new_n634));
  NAND3_X1  g448(.A1(new_n622), .A2(new_n585), .A3(new_n634), .ZN(new_n635));
  AOI21_X1  g449(.A(new_n629), .B1(new_n632), .B2(new_n635), .ZN(new_n636));
  OAI211_X1 g450(.A(new_n480), .B(new_n187), .C1(new_n477), .C2(new_n478), .ZN(new_n637));
  NOR2_X1   g451(.A1(new_n480), .A2(new_n187), .ZN(new_n638));
  INV_X1    g452(.A(new_n638), .ZN(new_n639));
  NAND2_X1  g453(.A1(new_n637), .A2(new_n639), .ZN(new_n640));
  NOR3_X1   g454(.A1(new_n477), .A2(new_n478), .A3(KEYINPUT33), .ZN(new_n641));
  INV_X1    g455(.A(KEYINPUT33), .ZN(new_n642));
  NOR2_X1   g456(.A1(new_n458), .A2(new_n459), .ZN(new_n643));
  AOI21_X1  g457(.A(KEYINPUT97), .B1(new_n464), .B2(new_n466), .ZN(new_n644));
  OAI21_X1  g458(.A(new_n475), .B1(new_n643), .B2(new_n644), .ZN(new_n645));
  INV_X1    g459(.A(new_n476), .ZN(new_n646));
  NAND2_X1  g460(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  NAND3_X1  g461(.A1(new_n468), .A2(new_n475), .A3(new_n476), .ZN(new_n648));
  AOI21_X1  g462(.A(new_n642), .B1(new_n647), .B2(new_n648), .ZN(new_n649));
  NOR2_X1   g463(.A1(new_n641), .A2(new_n649), .ZN(new_n650));
  AOI21_X1  g464(.A(new_n640), .B1(new_n650), .B2(G478), .ZN(new_n651));
  NAND2_X1  g465(.A1(new_n540), .A2(new_n651), .ZN(new_n652));
  INV_X1    g466(.A(new_n652), .ZN(new_n653));
  NAND3_X1  g467(.A1(new_n636), .A2(new_n547), .A3(new_n653), .ZN(new_n654));
  NAND2_X1  g468(.A1(new_n307), .A2(new_n187), .ZN(new_n655));
  AOI22_X1  g469(.A1(new_n655), .A2(G472), .B1(new_n307), .B2(new_n309), .ZN(new_n656));
  NAND3_X1  g470(.A1(new_n432), .A2(new_n656), .A3(new_n349), .ZN(new_n657));
  NOR2_X1   g471(.A1(new_n654), .A2(new_n657), .ZN(new_n658));
  XNOR2_X1  g472(.A(new_n658), .B(KEYINPUT100), .ZN(new_n659));
  XOR2_X1   g473(.A(KEYINPUT34), .B(G104), .Z(new_n660));
  XNOR2_X1  g474(.A(new_n659), .B(new_n660), .ZN(G6));
  INV_X1    g475(.A(new_n538), .ZN(new_n662));
  INV_X1    g476(.A(KEYINPUT101), .ZN(new_n663));
  NAND3_X1  g477(.A1(new_n534), .A2(new_n525), .A3(new_n537), .ZN(new_n664));
  NAND3_X1  g478(.A1(new_n662), .A2(new_n663), .A3(new_n664), .ZN(new_n665));
  OAI21_X1  g479(.A(KEYINPUT101), .B1(new_n538), .B2(new_n539), .ZN(new_n666));
  NAND2_X1  g480(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  NAND2_X1  g481(.A1(new_n667), .A2(new_n524), .ZN(new_n668));
  NOR2_X1   g482(.A1(new_n668), .A2(new_n487), .ZN(new_n669));
  NAND3_X1  g483(.A1(new_n669), .A2(new_n636), .A3(new_n547), .ZN(new_n670));
  NOR2_X1   g484(.A1(new_n670), .A2(new_n657), .ZN(new_n671));
  XNOR2_X1  g485(.A(KEYINPUT35), .B(G107), .ZN(new_n672));
  XNOR2_X1  g486(.A(new_n671), .B(new_n672), .ZN(G9));
  INV_X1    g487(.A(KEYINPUT36), .ZN(new_n674));
  NAND3_X1  g488(.A1(new_n336), .A2(new_n674), .A3(new_n340), .ZN(new_n675));
  NAND2_X1  g489(.A1(new_n340), .A2(new_n674), .ZN(new_n676));
  NAND2_X1  g490(.A1(new_n676), .A2(new_n335), .ZN(new_n677));
  NAND4_X1  g491(.A1(new_n675), .A2(new_n677), .A3(new_n187), .A4(new_n315), .ZN(new_n678));
  XNOR2_X1  g492(.A(new_n678), .B(KEYINPUT102), .ZN(new_n679));
  NOR2_X1   g493(.A1(new_n347), .A2(new_n679), .ZN(new_n680));
  INV_X1    g494(.A(new_n680), .ZN(new_n681));
  NAND4_X1  g495(.A1(new_n681), .A2(new_n548), .A3(new_n625), .A4(new_n624), .ZN(new_n682));
  NAND2_X1  g496(.A1(new_n432), .A2(new_n656), .ZN(new_n683));
  NOR2_X1   g497(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  XNOR2_X1  g498(.A(KEYINPUT37), .B(G110), .ZN(new_n685));
  XNOR2_X1  g499(.A(new_n684), .B(new_n685), .ZN(G12));
  INV_X1    g500(.A(G900), .ZN(new_n687));
  AOI21_X1  g501(.A(new_n543), .B1(new_n544), .B2(new_n687), .ZN(new_n688));
  INV_X1    g502(.A(new_n688), .ZN(new_n689));
  NAND4_X1  g503(.A1(new_n312), .A2(new_n432), .A3(new_n681), .A4(new_n689), .ZN(new_n690));
  INV_X1    g504(.A(new_n636), .ZN(new_n691));
  INV_X1    g505(.A(new_n669), .ZN(new_n692));
  NOR3_X1   g506(.A1(new_n690), .A2(new_n691), .A3(new_n692), .ZN(new_n693));
  XNOR2_X1  g507(.A(new_n693), .B(new_n221), .ZN(G30));
  XOR2_X1   g508(.A(new_n688), .B(KEYINPUT39), .Z(new_n695));
  NAND2_X1  g509(.A1(new_n432), .A2(new_n695), .ZN(new_n696));
  XOR2_X1   g510(.A(new_n696), .B(KEYINPUT40), .Z(new_n697));
  INV_X1    g511(.A(new_n300), .ZN(new_n698));
  NOR3_X1   g512(.A1(new_n284), .A2(new_n285), .A3(new_n280), .ZN(new_n699));
  AOI21_X1  g513(.A(KEYINPUT68), .B1(new_n288), .B2(new_n294), .ZN(new_n700));
  OAI21_X1  g514(.A(new_n303), .B1(new_n699), .B2(new_n700), .ZN(new_n701));
  NAND2_X1  g515(.A1(new_n701), .A2(new_n305), .ZN(new_n702));
  NAND3_X1  g516(.A1(new_n301), .A2(KEYINPUT31), .A3(new_n303), .ZN(new_n703));
  AOI21_X1  g517(.A(new_n698), .B1(new_n702), .B2(new_n703), .ZN(new_n704));
  INV_X1    g518(.A(new_n309), .ZN(new_n705));
  OAI21_X1  g519(.A(KEYINPUT32), .B1(new_n704), .B2(new_n705), .ZN(new_n706));
  NAND3_X1  g520(.A1(new_n307), .A2(new_n308), .A3(new_n309), .ZN(new_n707));
  NAND2_X1  g521(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  INV_X1    g522(.A(G472), .ZN(new_n709));
  NAND2_X1  g523(.A1(new_n268), .A2(new_n269), .ZN(new_n710));
  AOI21_X1  g524(.A(new_n709), .B1(new_n710), .B2(new_n264), .ZN(new_n711));
  NAND2_X1  g525(.A1(new_n701), .A2(new_n711), .ZN(new_n712));
  NAND2_X1  g526(.A1(G472), .A2(G902), .ZN(new_n713));
  NAND2_X1  g527(.A1(new_n712), .A2(new_n713), .ZN(new_n714));
  XNOR2_X1  g528(.A(new_n714), .B(KEYINPUT103), .ZN(new_n715));
  AOI21_X1  g529(.A(new_n681), .B1(new_n708), .B2(new_n715), .ZN(new_n716));
  NAND4_X1  g530(.A1(new_n485), .A2(new_n540), .A3(new_n625), .A4(new_n486), .ZN(new_n717));
  INV_X1    g531(.A(new_n717), .ZN(new_n718));
  XNOR2_X1  g532(.A(new_n624), .B(KEYINPUT38), .ZN(new_n719));
  NAND4_X1  g533(.A1(new_n697), .A2(new_n716), .A3(new_n718), .A4(new_n719), .ZN(new_n720));
  XNOR2_X1  g534(.A(new_n720), .B(new_n216), .ZN(G45));
  NAND2_X1  g535(.A1(new_n632), .A2(new_n635), .ZN(new_n722));
  NAND3_X1  g536(.A1(new_n540), .A2(new_n651), .A3(new_n689), .ZN(new_n723));
  INV_X1    g537(.A(new_n723), .ZN(new_n724));
  NAND3_X1  g538(.A1(new_n722), .A2(new_n625), .A3(new_n724), .ZN(new_n725));
  NAND2_X1  g539(.A1(new_n725), .A2(KEYINPUT104), .ZN(new_n726));
  AOI21_X1  g540(.A(new_n680), .B1(new_n708), .B2(new_n299), .ZN(new_n727));
  INV_X1    g541(.A(KEYINPUT104), .ZN(new_n728));
  NAND3_X1  g542(.A1(new_n636), .A2(new_n728), .A3(new_n724), .ZN(new_n729));
  NAND4_X1  g543(.A1(new_n726), .A2(new_n727), .A3(new_n729), .A4(new_n432), .ZN(new_n730));
  XNOR2_X1  g544(.A(new_n730), .B(G146), .ZN(G48));
  AND3_X1   g545(.A1(new_n424), .A2(new_n425), .A3(new_n187), .ZN(new_n732));
  AOI21_X1  g546(.A(new_n425), .B1(new_n424), .B2(new_n187), .ZN(new_n733));
  NOR2_X1   g547(.A1(new_n732), .A2(new_n733), .ZN(new_n734));
  NAND4_X1  g548(.A1(new_n312), .A2(new_n734), .A3(new_n349), .A4(new_n351), .ZN(new_n735));
  NOR2_X1   g549(.A1(new_n735), .A2(new_n654), .ZN(new_n736));
  XOR2_X1   g550(.A(KEYINPUT41), .B(G113), .Z(new_n737));
  XNOR2_X1  g551(.A(new_n736), .B(new_n737), .ZN(G15));
  NOR2_X1   g552(.A1(new_n735), .A2(new_n670), .ZN(new_n739));
  XNOR2_X1  g553(.A(new_n739), .B(new_n240), .ZN(G18));
  NAND3_X1  g554(.A1(new_n312), .A2(new_n548), .A3(new_n681), .ZN(new_n741));
  NAND3_X1  g555(.A1(new_n734), .A2(new_n351), .A3(new_n636), .ZN(new_n742));
  NOR2_X1   g556(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  XNOR2_X1  g557(.A(new_n743), .B(new_n238), .ZN(G21));
  AOI21_X1  g558(.A(new_n717), .B1(new_n632), .B2(new_n635), .ZN(new_n745));
  INV_X1    g559(.A(new_n745), .ZN(new_n746));
  NAND2_X1  g560(.A1(new_n424), .A2(new_n187), .ZN(new_n747));
  NAND2_X1  g561(.A1(new_n747), .A2(G469), .ZN(new_n748));
  NAND3_X1  g562(.A1(new_n748), .A2(new_n351), .A3(new_n426), .ZN(new_n749));
  NOR3_X1   g563(.A1(new_n746), .A2(new_n749), .A3(new_n546), .ZN(new_n750));
  INV_X1    g564(.A(KEYINPUT106), .ZN(new_n751));
  NAND2_X1  g565(.A1(new_n702), .A2(new_n703), .ZN(new_n752));
  OAI21_X1  g566(.A(new_n257), .B1(new_n272), .B2(new_n256), .ZN(new_n753));
  NAND2_X1  g567(.A1(new_n753), .A2(new_n264), .ZN(new_n754));
  AOI21_X1  g568(.A(new_n705), .B1(new_n752), .B2(new_n754), .ZN(new_n755));
  OAI21_X1  g569(.A(G472), .B1(new_n704), .B2(G902), .ZN(new_n756));
  NAND2_X1  g570(.A1(new_n756), .A2(KEYINPUT105), .ZN(new_n757));
  INV_X1    g571(.A(KEYINPUT105), .ZN(new_n758));
  NAND3_X1  g572(.A1(new_n655), .A2(new_n758), .A3(G472), .ZN(new_n759));
  AOI21_X1  g573(.A(new_n755), .B1(new_n757), .B2(new_n759), .ZN(new_n760));
  AOI21_X1  g574(.A(new_n751), .B1(new_n760), .B2(new_n349), .ZN(new_n761));
  INV_X1    g575(.A(new_n755), .ZN(new_n762));
  AOI21_X1  g576(.A(new_n758), .B1(new_n655), .B2(G472), .ZN(new_n763));
  AOI211_X1 g577(.A(KEYINPUT105), .B(new_n709), .C1(new_n307), .C2(new_n187), .ZN(new_n764));
  OAI211_X1 g578(.A(new_n349), .B(new_n762), .C1(new_n763), .C2(new_n764), .ZN(new_n765));
  NOR2_X1   g579(.A1(new_n765), .A2(KEYINPUT106), .ZN(new_n766));
  OAI21_X1  g580(.A(new_n750), .B1(new_n761), .B2(new_n766), .ZN(new_n767));
  XOR2_X1   g581(.A(KEYINPUT107), .B(G122), .Z(new_n768));
  XNOR2_X1  g582(.A(new_n767), .B(new_n768), .ZN(G24));
  INV_X1    g583(.A(KEYINPUT109), .ZN(new_n770));
  NAND2_X1  g584(.A1(new_n757), .A2(new_n759), .ZN(new_n771));
  XNOR2_X1  g585(.A(new_n723), .B(KEYINPUT108), .ZN(new_n772));
  NAND4_X1  g586(.A1(new_n771), .A2(new_n772), .A3(new_n681), .A4(new_n762), .ZN(new_n773));
  OAI21_X1  g587(.A(new_n770), .B1(new_n773), .B2(new_n742), .ZN(new_n774));
  AOI211_X1 g588(.A(new_n755), .B(new_n680), .C1(new_n757), .C2(new_n759), .ZN(new_n775));
  NOR2_X1   g589(.A1(new_n691), .A2(new_n749), .ZN(new_n776));
  NAND4_X1  g590(.A1(new_n775), .A2(new_n776), .A3(KEYINPUT109), .A4(new_n772), .ZN(new_n777));
  NAND2_X1  g591(.A1(new_n774), .A2(new_n777), .ZN(new_n778));
  XNOR2_X1  g592(.A(new_n778), .B(G125), .ZN(G27));
  AND3_X1   g593(.A1(new_n616), .A2(new_n625), .A3(new_n623), .ZN(new_n780));
  NAND2_X1  g594(.A1(new_n780), .A2(new_n432), .ZN(new_n781));
  INV_X1    g595(.A(new_n781), .ZN(new_n782));
  INV_X1    g596(.A(new_n349), .ZN(new_n783));
  AOI21_X1  g597(.A(new_n783), .B1(new_n708), .B2(new_n299), .ZN(new_n784));
  NAND4_X1  g598(.A1(new_n782), .A2(KEYINPUT42), .A3(new_n784), .A4(new_n772), .ZN(new_n785));
  INV_X1    g599(.A(KEYINPUT42), .ZN(new_n786));
  NAND4_X1  g600(.A1(new_n312), .A2(new_n780), .A3(new_n349), .A4(new_n432), .ZN(new_n787));
  INV_X1    g601(.A(new_n772), .ZN(new_n788));
  OAI21_X1  g602(.A(new_n786), .B1(new_n787), .B2(new_n788), .ZN(new_n789));
  NAND2_X1  g603(.A1(new_n785), .A2(new_n789), .ZN(new_n790));
  XOR2_X1   g604(.A(KEYINPUT110), .B(G131), .Z(new_n791));
  XNOR2_X1  g605(.A(new_n790), .B(new_n791), .ZN(G33));
  INV_X1    g606(.A(KEYINPUT111), .ZN(new_n793));
  NOR3_X1   g607(.A1(new_n668), .A2(new_n487), .A3(new_n688), .ZN(new_n794));
  NAND4_X1  g608(.A1(new_n782), .A2(new_n793), .A3(new_n784), .A4(new_n794), .ZN(new_n795));
  INV_X1    g609(.A(new_n794), .ZN(new_n796));
  OAI21_X1  g610(.A(KEYINPUT111), .B1(new_n787), .B2(new_n796), .ZN(new_n797));
  NAND2_X1  g611(.A1(new_n795), .A2(new_n797), .ZN(new_n798));
  XNOR2_X1  g612(.A(new_n798), .B(G134), .ZN(G36));
  OR2_X1    g613(.A1(new_n430), .A2(KEYINPUT45), .ZN(new_n800));
  NAND2_X1  g614(.A1(new_n430), .A2(KEYINPUT45), .ZN(new_n801));
  NAND3_X1  g615(.A1(new_n800), .A2(G469), .A3(new_n801), .ZN(new_n802));
  OAI21_X1  g616(.A(new_n802), .B1(new_n425), .B2(new_n187), .ZN(new_n803));
  INV_X1    g617(.A(KEYINPUT46), .ZN(new_n804));
  NAND2_X1  g618(.A1(new_n803), .A2(new_n804), .ZN(new_n805));
  NAND2_X1  g619(.A1(new_n805), .A2(new_n426), .ZN(new_n806));
  NOR2_X1   g620(.A1(new_n803), .A2(new_n804), .ZN(new_n807));
  NOR2_X1   g621(.A1(new_n806), .A2(new_n807), .ZN(new_n808));
  INV_X1    g622(.A(new_n695), .ZN(new_n809));
  NOR3_X1   g623(.A1(new_n808), .A2(new_n352), .A3(new_n809), .ZN(new_n810));
  NAND3_X1  g624(.A1(new_n616), .A2(new_n625), .A3(new_n623), .ZN(new_n811));
  OR2_X1    g625(.A1(new_n641), .A2(new_n649), .ZN(new_n812));
  OAI211_X1 g626(.A(new_n637), .B(new_n639), .C1(new_n812), .C2(new_n480), .ZN(new_n813));
  NOR3_X1   g627(.A1(new_n813), .A2(KEYINPUT43), .A3(new_n540), .ZN(new_n814));
  AOI21_X1  g628(.A(new_n813), .B1(KEYINPUT112), .B2(new_n540), .ZN(new_n815));
  OAI21_X1  g629(.A(new_n815), .B1(KEYINPUT112), .B2(new_n540), .ZN(new_n816));
  AOI21_X1  g630(.A(new_n814), .B1(new_n816), .B2(KEYINPUT43), .ZN(new_n817));
  NOR2_X1   g631(.A1(new_n656), .A2(new_n680), .ZN(new_n818));
  NAND2_X1  g632(.A1(new_n817), .A2(new_n818), .ZN(new_n819));
  INV_X1    g633(.A(new_n819), .ZN(new_n820));
  AOI21_X1  g634(.A(new_n811), .B1(new_n820), .B2(KEYINPUT44), .ZN(new_n821));
  OAI211_X1 g635(.A(new_n810), .B(new_n821), .C1(KEYINPUT44), .C2(new_n820), .ZN(new_n822));
  XNOR2_X1  g636(.A(KEYINPUT113), .B(G137), .ZN(new_n823));
  XNOR2_X1  g637(.A(new_n822), .B(new_n823), .ZN(G39));
  INV_X1    g638(.A(KEYINPUT114), .ZN(new_n825));
  INV_X1    g639(.A(KEYINPUT47), .ZN(new_n826));
  NOR2_X1   g640(.A1(new_n825), .A2(new_n826), .ZN(new_n827));
  OR3_X1    g641(.A1(new_n808), .A2(new_n352), .A3(new_n827), .ZN(new_n828));
  NOR2_X1   g642(.A1(KEYINPUT114), .A2(KEYINPUT47), .ZN(new_n829));
  OAI22_X1  g643(.A1(new_n808), .A2(new_n352), .B1(new_n829), .B2(new_n827), .ZN(new_n830));
  NOR4_X1   g644(.A1(new_n312), .A2(new_n811), .A3(new_n349), .A4(new_n723), .ZN(new_n831));
  NAND3_X1  g645(.A1(new_n828), .A2(new_n830), .A3(new_n831), .ZN(new_n832));
  XNOR2_X1  g646(.A(new_n832), .B(G140), .ZN(G42));
  AOI22_X1  g647(.A1(new_n828), .A2(new_n830), .B1(new_n352), .B2(new_n734), .ZN(new_n834));
  NOR2_X1   g648(.A1(new_n761), .A2(new_n766), .ZN(new_n835));
  NAND2_X1  g649(.A1(new_n817), .A2(new_n543), .ZN(new_n836));
  NOR2_X1   g650(.A1(new_n835), .A2(new_n836), .ZN(new_n837));
  NAND2_X1  g651(.A1(new_n837), .A2(new_n780), .ZN(new_n838));
  NOR2_X1   g652(.A1(new_n834), .A2(new_n838), .ZN(new_n839));
  NOR3_X1   g653(.A1(new_n836), .A2(new_n749), .A3(new_n811), .ZN(new_n840));
  NAND2_X1  g654(.A1(new_n708), .A2(new_n715), .ZN(new_n841));
  NAND2_X1  g655(.A1(new_n349), .A2(new_n543), .ZN(new_n842));
  NOR4_X1   g656(.A1(new_n841), .A2(new_n749), .A3(new_n842), .A4(new_n811), .ZN(new_n843));
  NOR2_X1   g657(.A1(new_n540), .A2(new_n651), .ZN(new_n844));
  AOI22_X1  g658(.A1(new_n840), .A2(new_n775), .B1(new_n843), .B2(new_n844), .ZN(new_n845));
  NOR3_X1   g659(.A1(new_n719), .A2(new_n625), .A3(new_n749), .ZN(new_n846));
  AND3_X1   g660(.A1(new_n837), .A2(KEYINPUT50), .A3(new_n846), .ZN(new_n847));
  AOI21_X1  g661(.A(KEYINPUT50), .B1(new_n837), .B2(new_n846), .ZN(new_n848));
  OAI21_X1  g662(.A(new_n845), .B1(new_n847), .B2(new_n848), .ZN(new_n849));
  AOI21_X1  g663(.A(new_n839), .B1(KEYINPUT117), .B2(new_n849), .ZN(new_n850));
  OAI21_X1  g664(.A(new_n850), .B1(KEYINPUT117), .B2(new_n849), .ZN(new_n851));
  INV_X1    g665(.A(KEYINPUT51), .ZN(new_n852));
  AND2_X1   g666(.A1(new_n851), .A2(new_n852), .ZN(new_n853));
  NAND2_X1  g667(.A1(new_n482), .A2(new_n483), .ZN(new_n854));
  INV_X1    g668(.A(new_n854), .ZN(new_n855));
  NAND4_X1  g669(.A1(new_n780), .A2(new_n524), .A3(new_n855), .A4(new_n667), .ZN(new_n856));
  OAI22_X1  g670(.A1(new_n773), .A2(new_n781), .B1(new_n690), .B2(new_n856), .ZN(new_n857));
  AOI21_X1  g671(.A(new_n857), .B1(new_n789), .B2(new_n785), .ZN(new_n858));
  AOI21_X1  g672(.A(new_n735), .B1(new_n654), .B2(new_n670), .ZN(new_n859));
  OAI22_X1  g673(.A1(new_n433), .A2(new_n626), .B1(new_n682), .B2(new_n683), .ZN(new_n860));
  OAI21_X1  g674(.A(new_n652), .B1(new_n855), .B2(new_n540), .ZN(new_n861));
  NAND4_X1  g675(.A1(new_n624), .A2(new_n861), .A3(new_n625), .A4(new_n547), .ZN(new_n862));
  OAI22_X1  g676(.A1(new_n741), .A2(new_n742), .B1(new_n657), .B2(new_n862), .ZN(new_n863));
  NOR3_X1   g677(.A1(new_n859), .A2(new_n860), .A3(new_n863), .ZN(new_n864));
  NAND4_X1  g678(.A1(new_n858), .A2(new_n864), .A3(new_n767), .A4(new_n798), .ZN(new_n865));
  AOI21_X1  g679(.A(new_n693), .B1(new_n774), .B2(new_n777), .ZN(new_n866));
  NAND2_X1  g680(.A1(new_n841), .A2(new_n680), .ZN(new_n867));
  NAND3_X1  g681(.A1(new_n745), .A2(new_n432), .A3(new_n689), .ZN(new_n868));
  OAI21_X1  g682(.A(KEYINPUT115), .B1(new_n867), .B2(new_n868), .ZN(new_n869));
  AND2_X1   g683(.A1(new_n432), .A2(new_n689), .ZN(new_n870));
  INV_X1    g684(.A(KEYINPUT115), .ZN(new_n871));
  NAND4_X1  g685(.A1(new_n716), .A2(new_n870), .A3(new_n871), .A4(new_n745), .ZN(new_n872));
  AND3_X1   g686(.A1(new_n869), .A2(new_n730), .A3(new_n872), .ZN(new_n873));
  NAND2_X1  g687(.A1(new_n866), .A2(new_n873), .ZN(new_n874));
  INV_X1    g688(.A(KEYINPUT52), .ZN(new_n875));
  NAND2_X1  g689(.A1(new_n874), .A2(new_n875), .ZN(new_n876));
  NAND3_X1  g690(.A1(new_n866), .A2(KEYINPUT52), .A3(new_n873), .ZN(new_n877));
  AOI21_X1  g691(.A(new_n865), .B1(new_n876), .B2(new_n877), .ZN(new_n878));
  XOR2_X1   g692(.A(KEYINPUT116), .B(KEYINPUT53), .Z(new_n879));
  INV_X1    g693(.A(new_n879), .ZN(new_n880));
  NAND2_X1  g694(.A1(new_n878), .A2(new_n880), .ZN(new_n881));
  OAI21_X1  g695(.A(new_n881), .B1(KEYINPUT53), .B2(new_n878), .ZN(new_n882));
  NAND2_X1  g696(.A1(new_n882), .A2(KEYINPUT54), .ZN(new_n883));
  INV_X1    g697(.A(new_n857), .ZN(new_n884));
  NAND3_X1  g698(.A1(new_n884), .A2(new_n790), .A3(new_n798), .ZN(new_n885));
  INV_X1    g699(.A(new_n863), .ZN(new_n886));
  INV_X1    g700(.A(new_n860), .ZN(new_n887));
  INV_X1    g701(.A(new_n735), .ZN(new_n888));
  INV_X1    g702(.A(new_n670), .ZN(new_n889));
  INV_X1    g703(.A(new_n654), .ZN(new_n890));
  OAI21_X1  g704(.A(new_n888), .B1(new_n889), .B2(new_n890), .ZN(new_n891));
  NAND4_X1  g705(.A1(new_n767), .A2(new_n886), .A3(new_n887), .A4(new_n891), .ZN(new_n892));
  NOR2_X1   g706(.A1(new_n885), .A2(new_n892), .ZN(new_n893));
  AND3_X1   g707(.A1(new_n866), .A2(KEYINPUT52), .A3(new_n873), .ZN(new_n894));
  AOI21_X1  g708(.A(KEYINPUT52), .B1(new_n866), .B2(new_n873), .ZN(new_n895));
  OAI21_X1  g709(.A(new_n893), .B1(new_n894), .B2(new_n895), .ZN(new_n896));
  NAND2_X1  g710(.A1(new_n896), .A2(new_n879), .ZN(new_n897));
  INV_X1    g711(.A(KEYINPUT54), .ZN(new_n898));
  OAI211_X1 g712(.A(new_n893), .B(KEYINPUT53), .C1(new_n894), .C2(new_n895), .ZN(new_n899));
  NAND3_X1  g713(.A1(new_n897), .A2(new_n898), .A3(new_n899), .ZN(new_n900));
  NAND2_X1  g714(.A1(new_n883), .A2(new_n900), .ZN(new_n901));
  AOI21_X1  g715(.A(KEYINPUT48), .B1(new_n840), .B2(new_n784), .ZN(new_n902));
  NAND3_X1  g716(.A1(new_n840), .A2(KEYINPUT48), .A3(new_n784), .ZN(new_n903));
  AOI211_X1 g717(.A(new_n542), .B(G953), .C1(new_n843), .C2(new_n653), .ZN(new_n904));
  NAND2_X1  g718(.A1(new_n903), .A2(new_n904), .ZN(new_n905));
  AOI211_X1 g719(.A(new_n902), .B(new_n905), .C1(new_n776), .C2(new_n837), .ZN(new_n906));
  OAI21_X1  g720(.A(KEYINPUT51), .B1(new_n834), .B2(new_n838), .ZN(new_n907));
  OAI21_X1  g721(.A(new_n906), .B1(new_n907), .B2(new_n849), .ZN(new_n908));
  NOR3_X1   g722(.A1(new_n853), .A2(new_n901), .A3(new_n908), .ZN(new_n909));
  NOR2_X1   g723(.A1(G952), .A2(G953), .ZN(new_n910));
  XOR2_X1   g724(.A(new_n734), .B(KEYINPUT49), .Z(new_n911));
  NAND3_X1  g725(.A1(new_n349), .A2(new_n625), .A3(new_n351), .ZN(new_n912));
  OR4_X1    g726(.A1(new_n841), .A2(new_n911), .A3(new_n816), .A4(new_n912), .ZN(new_n913));
  OAI22_X1  g727(.A1(new_n909), .A2(new_n910), .B1(new_n719), .B2(new_n913), .ZN(G75));
  NOR2_X1   g728(.A1(new_n258), .A2(G952), .ZN(new_n915));
  INV_X1    g729(.A(new_n915), .ZN(new_n916));
  AOI21_X1  g730(.A(new_n187), .B1(new_n897), .B2(new_n899), .ZN(new_n917));
  AOI21_X1  g731(.A(KEYINPUT56), .B1(new_n917), .B2(G210), .ZN(new_n918));
  XNOR2_X1  g732(.A(new_n610), .B(new_n617), .ZN(new_n919));
  XNOR2_X1  g733(.A(new_n919), .B(KEYINPUT55), .ZN(new_n920));
  OAI21_X1  g734(.A(new_n916), .B1(new_n918), .B2(new_n920), .ZN(new_n921));
  OAI21_X1  g735(.A(new_n899), .B1(new_n878), .B2(new_n880), .ZN(new_n922));
  NAND2_X1  g736(.A1(new_n922), .A2(G902), .ZN(new_n923));
  INV_X1    g737(.A(KEYINPUT118), .ZN(new_n924));
  NAND2_X1  g738(.A1(new_n923), .A2(new_n924), .ZN(new_n925));
  NAND2_X1  g739(.A1(new_n917), .A2(KEYINPUT118), .ZN(new_n926));
  AND2_X1   g740(.A1(new_n925), .A2(new_n926), .ZN(new_n927));
  NAND2_X1  g741(.A1(new_n927), .A2(new_n613), .ZN(new_n928));
  INV_X1    g742(.A(KEYINPUT56), .ZN(new_n929));
  AND2_X1   g743(.A1(new_n920), .A2(new_n929), .ZN(new_n930));
  AOI21_X1  g744(.A(new_n921), .B1(new_n928), .B2(new_n930), .ZN(G51));
  XNOR2_X1  g745(.A(KEYINPUT119), .B(KEYINPUT57), .ZN(new_n932));
  XNOR2_X1  g746(.A(new_n932), .B(new_n427), .ZN(new_n933));
  INV_X1    g747(.A(new_n900), .ZN(new_n934));
  AOI21_X1  g748(.A(new_n898), .B1(new_n897), .B2(new_n899), .ZN(new_n935));
  OAI21_X1  g749(.A(new_n933), .B1(new_n934), .B2(new_n935), .ZN(new_n936));
  INV_X1    g750(.A(KEYINPUT120), .ZN(new_n937));
  NAND2_X1  g751(.A1(new_n936), .A2(new_n937), .ZN(new_n938));
  OAI211_X1 g752(.A(KEYINPUT120), .B(new_n933), .C1(new_n934), .C2(new_n935), .ZN(new_n939));
  NAND3_X1  g753(.A1(new_n938), .A2(new_n424), .A3(new_n939), .ZN(new_n940));
  XNOR2_X1  g754(.A(new_n802), .B(KEYINPUT121), .ZN(new_n941));
  NAND2_X1  g755(.A1(new_n927), .A2(new_n941), .ZN(new_n942));
  AOI21_X1  g756(.A(new_n915), .B1(new_n940), .B2(new_n942), .ZN(G54));
  AND2_X1   g757(.A1(KEYINPUT58), .A2(G475), .ZN(new_n944));
  NAND3_X1  g758(.A1(new_n925), .A2(new_n926), .A3(new_n944), .ZN(new_n945));
  NAND3_X1  g759(.A1(new_n945), .A2(new_n533), .A3(new_n532), .ZN(new_n946));
  NAND4_X1  g760(.A1(new_n925), .A2(new_n926), .A3(new_n534), .A4(new_n944), .ZN(new_n947));
  AND3_X1   g761(.A1(new_n946), .A2(new_n916), .A3(new_n947), .ZN(G60));
  XOR2_X1   g762(.A(new_n638), .B(KEYINPUT59), .Z(new_n949));
  AOI21_X1  g763(.A(new_n812), .B1(new_n901), .B2(new_n949), .ZN(new_n950));
  OAI211_X1 g764(.A(new_n812), .B(new_n949), .C1(new_n934), .C2(new_n935), .ZN(new_n951));
  NAND2_X1  g765(.A1(new_n951), .A2(new_n916), .ZN(new_n952));
  NOR2_X1   g766(.A1(new_n950), .A2(new_n952), .ZN(G63));
  NAND2_X1  g767(.A1(G217), .A2(G902), .ZN(new_n954));
  XNOR2_X1  g768(.A(new_n954), .B(KEYINPUT60), .ZN(new_n955));
  INV_X1    g769(.A(new_n955), .ZN(new_n956));
  NAND2_X1  g770(.A1(new_n922), .A2(new_n956), .ZN(new_n957));
  NAND2_X1  g771(.A1(new_n957), .A2(KEYINPUT122), .ZN(new_n958));
  INV_X1    g772(.A(KEYINPUT122), .ZN(new_n959));
  NAND3_X1  g773(.A1(new_n922), .A2(new_n959), .A3(new_n956), .ZN(new_n960));
  XNOR2_X1  g774(.A(new_n343), .B(KEYINPUT123), .ZN(new_n961));
  NAND3_X1  g775(.A1(new_n958), .A2(new_n960), .A3(new_n961), .ZN(new_n962));
  AND2_X1   g776(.A1(new_n675), .A2(new_n677), .ZN(new_n963));
  AOI211_X1 g777(.A(KEYINPUT122), .B(new_n955), .C1(new_n897), .C2(new_n899), .ZN(new_n964));
  AOI21_X1  g778(.A(new_n959), .B1(new_n922), .B2(new_n956), .ZN(new_n965));
  OAI21_X1  g779(.A(new_n963), .B1(new_n964), .B2(new_n965), .ZN(new_n966));
  NAND3_X1  g780(.A1(new_n962), .A2(new_n966), .A3(new_n916), .ZN(new_n967));
  INV_X1    g781(.A(KEYINPUT61), .ZN(new_n968));
  NAND2_X1  g782(.A1(new_n967), .A2(new_n968), .ZN(new_n969));
  NAND4_X1  g783(.A1(new_n962), .A2(new_n966), .A3(KEYINPUT61), .A4(new_n916), .ZN(new_n970));
  NAND2_X1  g784(.A1(new_n969), .A2(new_n970), .ZN(G66));
  OAI21_X1  g785(.A(G953), .B1(new_n555), .B2(new_n545), .ZN(new_n972));
  INV_X1    g786(.A(new_n892), .ZN(new_n973));
  INV_X1    g787(.A(new_n258), .ZN(new_n974));
  OAI21_X1  g788(.A(new_n972), .B1(new_n973), .B2(new_n974), .ZN(new_n975));
  OAI21_X1  g789(.A(new_n601), .B1(G898), .B2(new_n258), .ZN(new_n976));
  XNOR2_X1  g790(.A(new_n975), .B(new_n976), .ZN(G69));
  OAI21_X1  g791(.A(new_n288), .B1(new_n282), .B2(new_n283), .ZN(new_n978));
  XNOR2_X1  g792(.A(new_n978), .B(new_n527), .ZN(new_n979));
  AOI21_X1  g793(.A(new_n979), .B1(G900), .B2(new_n974), .ZN(new_n980));
  AND3_X1   g794(.A1(new_n832), .A2(new_n822), .A3(new_n798), .ZN(new_n981));
  AND2_X1   g795(.A1(new_n866), .A2(new_n730), .ZN(new_n982));
  NAND3_X1  g796(.A1(new_n810), .A2(new_n784), .A3(new_n745), .ZN(new_n983));
  NAND4_X1  g797(.A1(new_n981), .A2(new_n790), .A3(new_n982), .A4(new_n983), .ZN(new_n984));
  OAI21_X1  g798(.A(new_n980), .B1(new_n984), .B2(new_n974), .ZN(new_n985));
  NAND4_X1  g799(.A1(new_n782), .A2(new_n784), .A3(new_n695), .A4(new_n861), .ZN(new_n986));
  XOR2_X1   g800(.A(new_n986), .B(KEYINPUT124), .Z(new_n987));
  AND3_X1   g801(.A1(new_n832), .A2(new_n822), .A3(new_n987), .ZN(new_n988));
  NAND2_X1  g802(.A1(new_n982), .A2(new_n720), .ZN(new_n989));
  NAND2_X1  g803(.A1(new_n989), .A2(KEYINPUT62), .ZN(new_n990));
  AND2_X1   g804(.A1(new_n988), .A2(new_n990), .ZN(new_n991));
  OR2_X1    g805(.A1(new_n989), .A2(KEYINPUT62), .ZN(new_n992));
  AOI21_X1  g806(.A(new_n974), .B1(new_n991), .B2(new_n992), .ZN(new_n993));
  INV_X1    g807(.A(new_n979), .ZN(new_n994));
  OAI21_X1  g808(.A(new_n985), .B1(new_n993), .B2(new_n994), .ZN(new_n995));
  AOI21_X1  g809(.A(new_n258), .B1(G227), .B2(G900), .ZN(new_n996));
  INV_X1    g810(.A(KEYINPUT125), .ZN(new_n997));
  AOI21_X1  g811(.A(new_n996), .B1(new_n985), .B2(new_n997), .ZN(new_n998));
  XOR2_X1   g812(.A(new_n995), .B(new_n998), .Z(G72));
  XNOR2_X1  g813(.A(new_n296), .B(KEYINPUT126), .ZN(new_n1000));
  NAND2_X1  g814(.A1(new_n1000), .A2(new_n278), .ZN(new_n1001));
  NAND4_X1  g815(.A1(new_n992), .A2(new_n973), .A3(new_n990), .A4(new_n988), .ZN(new_n1002));
  XOR2_X1   g816(.A(new_n713), .B(KEYINPUT63), .Z(new_n1003));
  AOI21_X1  g817(.A(new_n1001), .B1(new_n1002), .B2(new_n1003), .ZN(new_n1004));
  XOR2_X1   g818(.A(new_n1004), .B(KEYINPUT127), .Z(new_n1005));
  OAI21_X1  g819(.A(new_n1003), .B1(new_n984), .B2(new_n892), .ZN(new_n1006));
  INV_X1    g820(.A(new_n1000), .ZN(new_n1007));
  NAND3_X1  g821(.A1(new_n1006), .A2(new_n264), .A3(new_n1007), .ZN(new_n1008));
  OAI21_X1  g822(.A(new_n701), .B1(new_n296), .B2(new_n278), .ZN(new_n1009));
  NAND3_X1  g823(.A1(new_n882), .A2(new_n1003), .A3(new_n1009), .ZN(new_n1010));
  NAND3_X1  g824(.A1(new_n1008), .A2(new_n916), .A3(new_n1010), .ZN(new_n1011));
  NOR2_X1   g825(.A1(new_n1005), .A2(new_n1011), .ZN(G57));
endmodule


