//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 1 1 1 1 0 0 1 1 1 0 1 0 0 0 1 1 1 1 1 0 1 1 0 1 0 0 0 1 0 1 0 0 0 0 1 1 1 0 0 1 0 1 1 0 1 0 1 0 0 0 0 1 0 0 0 0 0 1 1 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:16:32 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n606, new_n607, new_n608,
    new_n609, new_n610, new_n611, new_n612, new_n613, new_n614, new_n615,
    new_n617, new_n618, new_n619, new_n620, new_n621, new_n622, new_n623,
    new_n624, new_n625, new_n626, new_n628, new_n629, new_n630, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n650, new_n651, new_n652, new_n653, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n677, new_n679,
    new_n680, new_n681, new_n682, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n691, new_n693, new_n694, new_n695, new_n696,
    new_n697, new_n698, new_n699, new_n700, new_n701, new_n702, new_n703,
    new_n704, new_n705, new_n706, new_n707, new_n708, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n725, new_n726,
    new_n727, new_n728, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n741, new_n742,
    new_n743, new_n744, new_n745, new_n746, new_n747, new_n748, new_n749,
    new_n750, new_n751, new_n752, new_n753, new_n754, new_n755, new_n756,
    new_n757, new_n758, new_n759, new_n760, new_n761, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n771,
    new_n772, new_n773, new_n775, new_n776, new_n778, new_n779, new_n780,
    new_n781, new_n782, new_n783, new_n784, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n799, new_n800, new_n801, new_n802, new_n803,
    new_n804, new_n805, new_n806, new_n807, new_n808, new_n809, new_n810,
    new_n811, new_n813, new_n814, new_n816, new_n817, new_n819, new_n820,
    new_n821, new_n822, new_n823, new_n824, new_n825, new_n826, new_n827,
    new_n828, new_n830, new_n831, new_n833, new_n834, new_n835, new_n836,
    new_n837, new_n839, new_n840, new_n841, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n869, new_n870, new_n871, new_n872, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880;
  INV_X1    g000(.A(KEYINPUT35), .ZN(new_n202));
  INV_X1    g001(.A(KEYINPUT34), .ZN(new_n203));
  INV_X1    g002(.A(G227gat), .ZN(new_n204));
  INV_X1    g003(.A(G233gat), .ZN(new_n205));
  NOR2_X1   g004(.A1(new_n204), .A2(new_n205), .ZN(new_n206));
  INV_X1    g005(.A(new_n206), .ZN(new_n207));
  AOI21_X1  g006(.A(new_n203), .B1(new_n207), .B2(KEYINPUT71), .ZN(new_n208));
  INV_X1    g007(.A(new_n208), .ZN(new_n209));
  INV_X1    g008(.A(KEYINPUT64), .ZN(new_n210));
  NAND2_X1  g009(.A1(G183gat), .A2(G190gat), .ZN(new_n211));
  INV_X1    g010(.A(KEYINPUT24), .ZN(new_n212));
  NOR2_X1   g011(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  AOI21_X1  g012(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n214));
  OAI21_X1  g013(.A(new_n210), .B1(new_n213), .B2(new_n214), .ZN(new_n215));
  NAND2_X1  g014(.A1(new_n211), .A2(new_n212), .ZN(new_n216));
  INV_X1    g015(.A(G183gat), .ZN(new_n217));
  INV_X1    g016(.A(G190gat), .ZN(new_n218));
  AOI22_X1  g017(.A1(new_n216), .A2(KEYINPUT64), .B1(new_n217), .B2(new_n218), .ZN(new_n219));
  INV_X1    g018(.A(KEYINPUT65), .ZN(new_n220));
  AND3_X1   g019(.A1(new_n215), .A2(new_n219), .A3(new_n220), .ZN(new_n221));
  AOI21_X1  g020(.A(new_n220), .B1(new_n215), .B2(new_n219), .ZN(new_n222));
  NOR2_X1   g021(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  AND2_X1   g022(.A1(G169gat), .A2(G176gat), .ZN(new_n224));
  NOR2_X1   g023(.A1(G169gat), .A2(G176gat), .ZN(new_n225));
  INV_X1    g024(.A(KEYINPUT23), .ZN(new_n226));
  NAND2_X1  g025(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  OAI21_X1  g026(.A(KEYINPUT23), .B1(G169gat), .B2(G176gat), .ZN(new_n228));
  AOI21_X1  g027(.A(new_n224), .B1(new_n227), .B2(new_n228), .ZN(new_n229));
  INV_X1    g028(.A(KEYINPUT66), .ZN(new_n230));
  NOR2_X1   g029(.A1(new_n229), .A2(new_n230), .ZN(new_n231));
  AOI211_X1 g030(.A(KEYINPUT66), .B(new_n224), .C1(new_n227), .C2(new_n228), .ZN(new_n232));
  NOR3_X1   g031(.A1(new_n231), .A2(new_n232), .A3(KEYINPUT25), .ZN(new_n233));
  INV_X1    g032(.A(new_n213), .ZN(new_n234));
  OAI211_X1 g033(.A(new_n234), .B(new_n216), .C1(G183gat), .C2(G190gat), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n235), .A2(new_n229), .ZN(new_n236));
  AOI22_X1  g035(.A1(new_n223), .A2(new_n233), .B1(KEYINPUT25), .B2(new_n236), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n225), .A2(KEYINPUT26), .ZN(new_n238));
  NAND2_X1  g037(.A1(new_n217), .A2(KEYINPUT27), .ZN(new_n239));
  INV_X1    g038(.A(KEYINPUT67), .ZN(new_n240));
  AOI21_X1  g039(.A(KEYINPUT28), .B1(new_n239), .B2(new_n240), .ZN(new_n241));
  XNOR2_X1  g040(.A(KEYINPUT27), .B(G183gat), .ZN(new_n242));
  OAI211_X1 g041(.A(new_n241), .B(new_n218), .C1(new_n240), .C2(new_n242), .ZN(new_n243));
  INV_X1    g042(.A(KEYINPUT27), .ZN(new_n244));
  NAND2_X1  g043(.A1(new_n244), .A2(G183gat), .ZN(new_n245));
  NAND3_X1  g044(.A1(new_n239), .A2(new_n245), .A3(new_n218), .ZN(new_n246));
  NAND2_X1  g045(.A1(new_n246), .A2(KEYINPUT28), .ZN(new_n247));
  AND3_X1   g046(.A1(new_n243), .A2(KEYINPUT68), .A3(new_n247), .ZN(new_n248));
  AOI21_X1  g047(.A(KEYINPUT68), .B1(new_n243), .B2(new_n247), .ZN(new_n249));
  OAI211_X1 g048(.A(new_n238), .B(new_n211), .C1(new_n248), .C2(new_n249), .ZN(new_n250));
  NOR3_X1   g049(.A1(new_n224), .A2(new_n225), .A3(KEYINPUT26), .ZN(new_n251));
  OAI21_X1  g050(.A(new_n237), .B1(new_n250), .B2(new_n251), .ZN(new_n252));
  INV_X1    g051(.A(G134gat), .ZN(new_n253));
  INV_X1    g052(.A(G113gat), .ZN(new_n254));
  INV_X1    g053(.A(G120gat), .ZN(new_n255));
  NAND2_X1  g054(.A1(new_n254), .A2(new_n255), .ZN(new_n256));
  INV_X1    g055(.A(KEYINPUT1), .ZN(new_n257));
  NAND2_X1  g056(.A1(G113gat), .A2(G120gat), .ZN(new_n258));
  NAND3_X1  g057(.A1(new_n256), .A2(new_n257), .A3(new_n258), .ZN(new_n259));
  INV_X1    g058(.A(G127gat), .ZN(new_n260));
  NAND3_X1  g059(.A1(new_n259), .A2(KEYINPUT69), .A3(new_n260), .ZN(new_n261));
  INV_X1    g060(.A(new_n261), .ZN(new_n262));
  AOI21_X1  g061(.A(new_n260), .B1(new_n259), .B2(KEYINPUT69), .ZN(new_n263));
  OAI21_X1  g062(.A(new_n253), .B1(new_n262), .B2(new_n263), .ZN(new_n264));
  NAND2_X1  g063(.A1(new_n259), .A2(KEYINPUT69), .ZN(new_n265));
  NAND2_X1  g064(.A1(new_n265), .A2(G127gat), .ZN(new_n266));
  NAND3_X1  g065(.A1(new_n266), .A2(G134gat), .A3(new_n261), .ZN(new_n267));
  NAND2_X1  g066(.A1(new_n264), .A2(new_n267), .ZN(new_n268));
  NAND2_X1  g067(.A1(new_n252), .A2(new_n268), .ZN(new_n269));
  NAND2_X1  g068(.A1(new_n243), .A2(new_n247), .ZN(new_n270));
  INV_X1    g069(.A(KEYINPUT68), .ZN(new_n271));
  NAND2_X1  g070(.A1(new_n270), .A2(new_n271), .ZN(new_n272));
  NAND3_X1  g071(.A1(new_n243), .A2(KEYINPUT68), .A3(new_n247), .ZN(new_n273));
  NAND2_X1  g072(.A1(new_n272), .A2(new_n273), .ZN(new_n274));
  INV_X1    g073(.A(new_n251), .ZN(new_n275));
  NAND4_X1  g074(.A1(new_n274), .A2(new_n275), .A3(new_n238), .A4(new_n211), .ZN(new_n276));
  INV_X1    g075(.A(new_n268), .ZN(new_n277));
  NAND3_X1  g076(.A1(new_n276), .A2(new_n277), .A3(new_n237), .ZN(new_n278));
  NAND3_X1  g077(.A1(new_n269), .A2(new_n206), .A3(new_n278), .ZN(new_n279));
  XNOR2_X1  g078(.A(G15gat), .B(G43gat), .ZN(new_n280));
  XNOR2_X1  g079(.A(new_n280), .B(G71gat), .ZN(new_n281));
  INV_X1    g080(.A(G99gat), .ZN(new_n282));
  XNOR2_X1  g081(.A(new_n281), .B(new_n282), .ZN(new_n283));
  NAND2_X1  g082(.A1(new_n283), .A2(KEYINPUT33), .ZN(new_n284));
  NAND3_X1  g083(.A1(new_n279), .A2(KEYINPUT32), .A3(new_n284), .ZN(new_n285));
  INV_X1    g084(.A(KEYINPUT70), .ZN(new_n286));
  NAND2_X1  g085(.A1(new_n285), .A2(new_n286), .ZN(new_n287));
  NAND4_X1  g086(.A1(new_n279), .A2(KEYINPUT70), .A3(KEYINPUT32), .A4(new_n284), .ZN(new_n288));
  NAND2_X1  g087(.A1(new_n287), .A2(new_n288), .ZN(new_n289));
  NAND2_X1  g088(.A1(new_n269), .A2(new_n278), .ZN(new_n290));
  NAND2_X1  g089(.A1(new_n290), .A2(new_n207), .ZN(new_n291));
  INV_X1    g090(.A(KEYINPUT33), .ZN(new_n292));
  OAI21_X1  g091(.A(new_n279), .B1(KEYINPUT32), .B2(new_n292), .ZN(new_n293));
  NAND2_X1  g092(.A1(new_n293), .A2(new_n283), .ZN(new_n294));
  AND3_X1   g093(.A1(new_n289), .A2(new_n291), .A3(new_n294), .ZN(new_n295));
  AOI21_X1  g094(.A(new_n291), .B1(new_n289), .B2(new_n294), .ZN(new_n296));
  OAI21_X1  g095(.A(new_n209), .B1(new_n295), .B2(new_n296), .ZN(new_n297));
  NAND2_X1  g096(.A1(new_n289), .A2(new_n294), .ZN(new_n298));
  INV_X1    g097(.A(new_n291), .ZN(new_n299));
  NAND2_X1  g098(.A1(new_n298), .A2(new_n299), .ZN(new_n300));
  NAND3_X1  g099(.A1(new_n289), .A2(new_n291), .A3(new_n294), .ZN(new_n301));
  NAND3_X1  g100(.A1(new_n300), .A2(new_n208), .A3(new_n301), .ZN(new_n302));
  XOR2_X1   g101(.A(G78gat), .B(G106gat), .Z(new_n303));
  XNOR2_X1  g102(.A(new_n303), .B(KEYINPUT31), .ZN(new_n304));
  INV_X1    g103(.A(G50gat), .ZN(new_n305));
  XNOR2_X1  g104(.A(new_n304), .B(new_n305), .ZN(new_n306));
  INV_X1    g105(.A(new_n306), .ZN(new_n307));
  INV_X1    g106(.A(KEYINPUT80), .ZN(new_n308));
  XOR2_X1   g107(.A(G155gat), .B(G162gat), .Z(new_n309));
  INV_X1    g108(.A(new_n309), .ZN(new_n310));
  INV_X1    g109(.A(G155gat), .ZN(new_n311));
  INV_X1    g110(.A(G162gat), .ZN(new_n312));
  OAI21_X1  g111(.A(KEYINPUT2), .B1(new_n311), .B2(new_n312), .ZN(new_n313));
  XOR2_X1   g112(.A(G141gat), .B(G148gat), .Z(new_n314));
  NAND3_X1  g113(.A1(new_n310), .A2(new_n313), .A3(new_n314), .ZN(new_n315));
  NAND2_X1  g114(.A1(new_n314), .A2(new_n313), .ZN(new_n316));
  NAND2_X1  g115(.A1(new_n316), .A2(new_n309), .ZN(new_n317));
  INV_X1    g116(.A(KEYINPUT3), .ZN(new_n318));
  NAND3_X1  g117(.A1(new_n315), .A2(new_n317), .A3(new_n318), .ZN(new_n319));
  INV_X1    g118(.A(KEYINPUT29), .ZN(new_n320));
  NAND2_X1  g119(.A1(new_n319), .A2(new_n320), .ZN(new_n321));
  XNOR2_X1  g120(.A(G197gat), .B(G204gat), .ZN(new_n322));
  INV_X1    g121(.A(G211gat), .ZN(new_n323));
  INV_X1    g122(.A(G218gat), .ZN(new_n324));
  NOR2_X1   g123(.A1(new_n323), .A2(new_n324), .ZN(new_n325));
  OAI21_X1  g124(.A(new_n322), .B1(KEYINPUT22), .B2(new_n325), .ZN(new_n326));
  XOR2_X1   g125(.A(G211gat), .B(G218gat), .Z(new_n327));
  XNOR2_X1  g126(.A(new_n326), .B(new_n327), .ZN(new_n328));
  INV_X1    g127(.A(new_n328), .ZN(new_n329));
  NAND2_X1  g128(.A1(new_n321), .A2(new_n329), .ZN(new_n330));
  INV_X1    g129(.A(G228gat), .ZN(new_n331));
  OAI21_X1  g130(.A(KEYINPUT78), .B1(new_n331), .B2(new_n205), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n315), .A2(new_n317), .ZN(new_n333));
  INV_X1    g132(.A(new_n333), .ZN(new_n334));
  AOI21_X1  g133(.A(KEYINPUT3), .B1(new_n328), .B2(new_n320), .ZN(new_n335));
  OAI211_X1 g134(.A(new_n330), .B(new_n332), .C1(new_n334), .C2(new_n335), .ZN(new_n336));
  NOR3_X1   g135(.A1(new_n331), .A2(new_n205), .A3(KEYINPUT78), .ZN(new_n337));
  OR2_X1    g136(.A1(new_n336), .A2(new_n337), .ZN(new_n338));
  NAND2_X1  g137(.A1(new_n336), .A2(new_n337), .ZN(new_n339));
  NAND2_X1  g138(.A1(new_n338), .A2(new_n339), .ZN(new_n340));
  XOR2_X1   g139(.A(KEYINPUT79), .B(G22gat), .Z(new_n341));
  INV_X1    g140(.A(new_n341), .ZN(new_n342));
  OAI21_X1  g141(.A(new_n308), .B1(new_n340), .B2(new_n342), .ZN(new_n343));
  NAND2_X1  g142(.A1(new_n340), .A2(new_n342), .ZN(new_n344));
  NAND2_X1  g143(.A1(new_n343), .A2(new_n344), .ZN(new_n345));
  NOR3_X1   g144(.A1(new_n340), .A2(new_n308), .A3(new_n342), .ZN(new_n346));
  OAI21_X1  g145(.A(new_n307), .B1(new_n345), .B2(new_n346), .ZN(new_n347));
  INV_X1    g146(.A(G22gat), .ZN(new_n348));
  OAI211_X1 g147(.A(new_n344), .B(new_n306), .C1(new_n348), .C2(new_n340), .ZN(new_n349));
  NAND2_X1  g148(.A1(new_n347), .A2(new_n349), .ZN(new_n350));
  NAND3_X1  g149(.A1(new_n297), .A2(new_n302), .A3(new_n350), .ZN(new_n351));
  INV_X1    g150(.A(KEYINPUT84), .ZN(new_n352));
  NAND2_X1  g151(.A1(new_n351), .A2(new_n352), .ZN(new_n353));
  NAND4_X1  g152(.A1(new_n297), .A2(new_n302), .A3(KEYINPUT84), .A4(new_n350), .ZN(new_n354));
  NAND2_X1  g153(.A1(new_n353), .A2(new_n354), .ZN(new_n355));
  NOR3_X1   g154(.A1(new_n262), .A2(new_n253), .A3(new_n263), .ZN(new_n356));
  AOI21_X1  g155(.A(G134gat), .B1(new_n266), .B2(new_n261), .ZN(new_n357));
  OAI21_X1  g156(.A(new_n334), .B1(new_n356), .B2(new_n357), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n358), .A2(KEYINPUT4), .ZN(new_n359));
  INV_X1    g158(.A(KEYINPUT4), .ZN(new_n360));
  NAND3_X1  g159(.A1(new_n268), .A2(new_n360), .A3(new_n334), .ZN(new_n361));
  NAND2_X1  g160(.A1(new_n359), .A2(new_n361), .ZN(new_n362));
  NAND2_X1  g161(.A1(new_n333), .A2(KEYINPUT3), .ZN(new_n363));
  AND3_X1   g162(.A1(new_n264), .A2(KEYINPUT74), .A3(new_n267), .ZN(new_n364));
  AOI21_X1  g163(.A(KEYINPUT74), .B1(new_n264), .B2(new_n267), .ZN(new_n365));
  OAI211_X1 g164(.A(new_n363), .B(new_n319), .C1(new_n364), .C2(new_n365), .ZN(new_n366));
  NAND2_X1  g165(.A1(G225gat), .A2(G233gat), .ZN(new_n367));
  INV_X1    g166(.A(new_n367), .ZN(new_n368));
  NOR2_X1   g167(.A1(new_n368), .A2(KEYINPUT5), .ZN(new_n369));
  AND3_X1   g168(.A1(new_n362), .A2(new_n366), .A3(new_n369), .ZN(new_n370));
  INV_X1    g169(.A(KEYINPUT5), .ZN(new_n371));
  OAI21_X1  g170(.A(new_n333), .B1(new_n364), .B2(new_n365), .ZN(new_n372));
  NAND2_X1  g171(.A1(new_n372), .A2(new_n358), .ZN(new_n373));
  AOI21_X1  g172(.A(new_n371), .B1(new_n373), .B2(new_n368), .ZN(new_n374));
  INV_X1    g173(.A(KEYINPUT75), .ZN(new_n375));
  NAND3_X1  g174(.A1(new_n359), .A2(new_n375), .A3(new_n361), .ZN(new_n376));
  OR2_X1    g175(.A1(new_n361), .A2(new_n375), .ZN(new_n377));
  NAND4_X1  g176(.A1(new_n376), .A2(new_n377), .A3(new_n366), .A4(new_n367), .ZN(new_n378));
  AOI21_X1  g177(.A(new_n370), .B1(new_n374), .B2(new_n378), .ZN(new_n379));
  XOR2_X1   g178(.A(G1gat), .B(G29gat), .Z(new_n380));
  XNOR2_X1  g179(.A(KEYINPUT76), .B(KEYINPUT0), .ZN(new_n381));
  XNOR2_X1  g180(.A(new_n380), .B(new_n381), .ZN(new_n382));
  XNOR2_X1  g181(.A(G57gat), .B(G85gat), .ZN(new_n383));
  XOR2_X1   g182(.A(new_n382), .B(new_n383), .Z(new_n384));
  INV_X1    g183(.A(new_n384), .ZN(new_n385));
  NOR2_X1   g184(.A1(new_n379), .A2(new_n385), .ZN(new_n386));
  INV_X1    g185(.A(new_n386), .ZN(new_n387));
  AOI21_X1  g186(.A(KEYINPUT6), .B1(new_n379), .B2(new_n385), .ZN(new_n388));
  NAND2_X1  g187(.A1(new_n387), .A2(new_n388), .ZN(new_n389));
  INV_X1    g188(.A(new_n379), .ZN(new_n390));
  NAND3_X1  g189(.A1(new_n390), .A2(KEYINPUT6), .A3(new_n384), .ZN(new_n391));
  NAND2_X1  g190(.A1(new_n389), .A2(new_n391), .ZN(new_n392));
  NAND2_X1  g191(.A1(new_n252), .A2(new_n320), .ZN(new_n393));
  NAND2_X1  g192(.A1(G226gat), .A2(G233gat), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n393), .A2(new_n394), .ZN(new_n395));
  INV_X1    g194(.A(new_n394), .ZN(new_n396));
  NAND2_X1  g195(.A1(new_n252), .A2(new_n396), .ZN(new_n397));
  INV_X1    g196(.A(KEYINPUT72), .ZN(new_n398));
  NAND2_X1  g197(.A1(new_n397), .A2(new_n398), .ZN(new_n399));
  NAND3_X1  g198(.A1(new_n252), .A2(KEYINPUT72), .A3(new_n396), .ZN(new_n400));
  NAND3_X1  g199(.A1(new_n395), .A2(new_n399), .A3(new_n400), .ZN(new_n401));
  INV_X1    g200(.A(KEYINPUT73), .ZN(new_n402));
  NAND3_X1  g201(.A1(new_n401), .A2(new_n402), .A3(new_n329), .ZN(new_n403));
  XOR2_X1   g202(.A(G8gat), .B(G36gat), .Z(new_n404));
  XNOR2_X1  g203(.A(new_n404), .B(G64gat), .ZN(new_n405));
  INV_X1    g204(.A(G92gat), .ZN(new_n406));
  XNOR2_X1  g205(.A(new_n405), .B(new_n406), .ZN(new_n407));
  AOI211_X1 g206(.A(new_n398), .B(new_n394), .C1(new_n276), .C2(new_n237), .ZN(new_n408));
  AOI21_X1  g207(.A(KEYINPUT72), .B1(new_n252), .B2(new_n396), .ZN(new_n409));
  NOR2_X1   g208(.A1(new_n408), .A2(new_n409), .ZN(new_n410));
  AOI21_X1  g209(.A(new_n328), .B1(new_n410), .B2(new_n395), .ZN(new_n411));
  AOI21_X1  g210(.A(KEYINPUT29), .B1(new_n276), .B2(new_n237), .ZN(new_n412));
  OAI211_X1 g211(.A(new_n397), .B(new_n328), .C1(new_n412), .C2(new_n396), .ZN(new_n413));
  NAND2_X1  g212(.A1(new_n413), .A2(KEYINPUT73), .ZN(new_n414));
  OAI211_X1 g213(.A(new_n403), .B(new_n407), .C1(new_n411), .C2(new_n414), .ZN(new_n415));
  NAND2_X1  g214(.A1(new_n415), .A2(KEYINPUT30), .ZN(new_n416));
  NAND2_X1  g215(.A1(new_n401), .A2(new_n329), .ZN(new_n417));
  NAND3_X1  g216(.A1(new_n417), .A2(KEYINPUT73), .A3(new_n413), .ZN(new_n418));
  AOI21_X1  g217(.A(new_n407), .B1(new_n418), .B2(new_n403), .ZN(new_n419));
  NOR2_X1   g218(.A1(new_n416), .A2(new_n419), .ZN(new_n420));
  AOI21_X1  g219(.A(new_n414), .B1(new_n329), .B2(new_n401), .ZN(new_n421));
  AND3_X1   g220(.A1(new_n401), .A2(new_n402), .A3(new_n329), .ZN(new_n422));
  NOR2_X1   g221(.A1(new_n421), .A2(new_n422), .ZN(new_n423));
  NOR3_X1   g222(.A1(new_n423), .A2(KEYINPUT30), .A3(new_n407), .ZN(new_n424));
  OAI21_X1  g223(.A(new_n392), .B1(new_n420), .B2(new_n424), .ZN(new_n425));
  NAND2_X1  g224(.A1(new_n425), .A2(KEYINPUT77), .ZN(new_n426));
  INV_X1    g225(.A(new_n407), .ZN(new_n427));
  OAI21_X1  g226(.A(new_n427), .B1(new_n421), .B2(new_n422), .ZN(new_n428));
  NAND3_X1  g227(.A1(new_n428), .A2(KEYINPUT30), .A3(new_n415), .ZN(new_n429));
  NAND2_X1  g228(.A1(new_n418), .A2(new_n403), .ZN(new_n430));
  INV_X1    g229(.A(KEYINPUT30), .ZN(new_n431));
  NAND3_X1  g230(.A1(new_n430), .A2(new_n431), .A3(new_n427), .ZN(new_n432));
  NAND2_X1  g231(.A1(new_n429), .A2(new_n432), .ZN(new_n433));
  INV_X1    g232(.A(KEYINPUT77), .ZN(new_n434));
  NAND3_X1  g233(.A1(new_n433), .A2(new_n434), .A3(new_n392), .ZN(new_n435));
  NAND2_X1  g234(.A1(new_n426), .A2(new_n435), .ZN(new_n436));
  AOI21_X1  g235(.A(new_n202), .B1(new_n355), .B2(new_n436), .ZN(new_n437));
  NOR3_X1   g236(.A1(new_n351), .A2(new_n425), .A3(KEYINPUT35), .ZN(new_n438));
  INV_X1    g237(.A(new_n350), .ZN(new_n439));
  NAND3_X1  g238(.A1(new_n426), .A2(new_n439), .A3(new_n435), .ZN(new_n440));
  INV_X1    g239(.A(KEYINPUT36), .ZN(new_n441));
  INV_X1    g240(.A(new_n302), .ZN(new_n442));
  AOI21_X1  g241(.A(new_n208), .B1(new_n300), .B2(new_n301), .ZN(new_n443));
  OAI21_X1  g242(.A(new_n441), .B1(new_n442), .B2(new_n443), .ZN(new_n444));
  NAND3_X1  g243(.A1(new_n297), .A2(new_n302), .A3(KEYINPUT36), .ZN(new_n445));
  NAND2_X1  g244(.A1(new_n444), .A2(new_n445), .ZN(new_n446));
  NAND2_X1  g245(.A1(new_n440), .A2(new_n446), .ZN(new_n447));
  XNOR2_X1  g246(.A(new_n388), .B(new_n386), .ZN(new_n448));
  INV_X1    g247(.A(KEYINPUT37), .ZN(new_n449));
  OAI21_X1  g248(.A(new_n449), .B1(new_n421), .B2(new_n422), .ZN(new_n450));
  INV_X1    g249(.A(KEYINPUT38), .ZN(new_n451));
  NAND3_X1  g250(.A1(new_n450), .A2(new_n451), .A3(new_n407), .ZN(new_n452));
  AOI21_X1  g251(.A(new_n449), .B1(new_n401), .B2(new_n328), .ZN(new_n453));
  NAND3_X1  g252(.A1(new_n395), .A2(new_n329), .A3(new_n397), .ZN(new_n454));
  NAND2_X1  g253(.A1(new_n453), .A2(new_n454), .ZN(new_n455));
  INV_X1    g254(.A(KEYINPUT83), .ZN(new_n456));
  NAND2_X1  g255(.A1(new_n455), .A2(new_n456), .ZN(new_n457));
  NAND3_X1  g256(.A1(new_n453), .A2(KEYINPUT83), .A3(new_n454), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  OAI211_X1 g258(.A(new_n448), .B(new_n428), .C1(new_n452), .C2(new_n459), .ZN(new_n460));
  AOI21_X1  g259(.A(new_n427), .B1(new_n430), .B2(new_n449), .ZN(new_n461));
  NAND2_X1  g260(.A1(new_n423), .A2(KEYINPUT37), .ZN(new_n462));
  AOI21_X1  g261(.A(new_n451), .B1(new_n461), .B2(new_n462), .ZN(new_n463));
  OAI21_X1  g262(.A(new_n350), .B1(new_n460), .B2(new_n463), .ZN(new_n464));
  NOR2_X1   g263(.A1(new_n373), .A2(new_n368), .ZN(new_n465));
  AOI21_X1  g264(.A(new_n367), .B1(new_n362), .B2(new_n366), .ZN(new_n466));
  INV_X1    g265(.A(KEYINPUT39), .ZN(new_n467));
  OR3_X1    g266(.A1(new_n465), .A2(new_n466), .A3(new_n467), .ZN(new_n468));
  AOI21_X1  g267(.A(new_n384), .B1(new_n466), .B2(new_n467), .ZN(new_n469));
  NAND2_X1  g268(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  INV_X1    g269(.A(KEYINPUT40), .ZN(new_n471));
  NAND2_X1  g270(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  XNOR2_X1  g271(.A(new_n472), .B(KEYINPUT81), .ZN(new_n473));
  INV_X1    g272(.A(new_n473), .ZN(new_n474));
  NAND3_X1  g273(.A1(new_n468), .A2(KEYINPUT40), .A3(new_n469), .ZN(new_n475));
  NAND4_X1  g274(.A1(new_n429), .A2(new_n387), .A3(new_n432), .A4(new_n475), .ZN(new_n476));
  OAI21_X1  g275(.A(KEYINPUT82), .B1(new_n474), .B2(new_n476), .ZN(new_n477));
  AND3_X1   g276(.A1(new_n429), .A2(new_n475), .A3(new_n432), .ZN(new_n478));
  INV_X1    g277(.A(KEYINPUT82), .ZN(new_n479));
  NAND4_X1  g278(.A1(new_n478), .A2(new_n479), .A3(new_n387), .A4(new_n473), .ZN(new_n480));
  AOI21_X1  g279(.A(new_n464), .B1(new_n477), .B2(new_n480), .ZN(new_n481));
  OAI22_X1  g280(.A1(new_n437), .A2(new_n438), .B1(new_n447), .B2(new_n481), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n482), .A2(KEYINPUT85), .ZN(new_n483));
  NAND2_X1  g282(.A1(new_n480), .A2(new_n477), .ZN(new_n484));
  INV_X1    g283(.A(new_n464), .ZN(new_n485));
  NAND2_X1  g284(.A1(new_n484), .A2(new_n485), .ZN(new_n486));
  NAND3_X1  g285(.A1(new_n486), .A2(new_n440), .A3(new_n446), .ZN(new_n487));
  INV_X1    g286(.A(new_n438), .ZN(new_n488));
  AOI22_X1  g287(.A1(new_n353), .A2(new_n354), .B1(new_n426), .B2(new_n435), .ZN(new_n489));
  OAI21_X1  g288(.A(new_n488), .B1(new_n489), .B2(new_n202), .ZN(new_n490));
  INV_X1    g289(.A(KEYINPUT85), .ZN(new_n491));
  NAND3_X1  g290(.A1(new_n487), .A2(new_n490), .A3(new_n491), .ZN(new_n492));
  XNOR2_X1  g291(.A(G43gat), .B(G50gat), .ZN(new_n493));
  NOR2_X1   g292(.A1(new_n493), .A2(KEYINPUT15), .ZN(new_n494));
  XOR2_X1   g293(.A(KEYINPUT88), .B(G36gat), .Z(new_n495));
  NAND2_X1  g294(.A1(new_n495), .A2(G29gat), .ZN(new_n496));
  INV_X1    g295(.A(KEYINPUT90), .ZN(new_n497));
  XNOR2_X1  g296(.A(new_n496), .B(new_n497), .ZN(new_n498));
  NOR2_X1   g297(.A1(G29gat), .A2(G36gat), .ZN(new_n499));
  INV_X1    g298(.A(KEYINPUT14), .ZN(new_n500));
  XNOR2_X1  g299(.A(new_n499), .B(new_n500), .ZN(new_n501));
  XNOR2_X1  g300(.A(new_n501), .B(KEYINPUT89), .ZN(new_n502));
  NAND2_X1  g301(.A1(new_n498), .A2(new_n502), .ZN(new_n503));
  NAND2_X1  g302(.A1(new_n493), .A2(KEYINPUT15), .ZN(new_n504));
  AOI21_X1  g303(.A(new_n494), .B1(new_n503), .B2(new_n504), .ZN(new_n505));
  NAND4_X1  g304(.A1(new_n496), .A2(new_n501), .A3(KEYINPUT15), .A4(new_n493), .ZN(new_n506));
  NAND2_X1  g305(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  INV_X1    g306(.A(G8gat), .ZN(new_n508));
  XNOR2_X1  g307(.A(G15gat), .B(G22gat), .ZN(new_n509));
  INV_X1    g308(.A(KEYINPUT16), .ZN(new_n510));
  OAI21_X1  g309(.A(new_n509), .B1(new_n510), .B2(G1gat), .ZN(new_n511));
  AOI21_X1  g310(.A(new_n508), .B1(new_n511), .B2(KEYINPUT91), .ZN(new_n512));
  OAI21_X1  g311(.A(new_n511), .B1(G1gat), .B2(new_n509), .ZN(new_n513));
  XNOR2_X1  g312(.A(new_n512), .B(new_n513), .ZN(new_n514));
  INV_X1    g313(.A(new_n514), .ZN(new_n515));
  NOR2_X1   g314(.A1(new_n507), .A2(new_n515), .ZN(new_n516));
  XOR2_X1   g315(.A(new_n507), .B(KEYINPUT17), .Z(new_n517));
  AOI21_X1  g316(.A(new_n516), .B1(new_n517), .B2(new_n515), .ZN(new_n518));
  NAND2_X1  g317(.A1(G229gat), .A2(G233gat), .ZN(new_n519));
  NAND2_X1  g318(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  XNOR2_X1  g319(.A(new_n520), .B(KEYINPUT18), .ZN(new_n521));
  XNOR2_X1  g320(.A(new_n507), .B(new_n515), .ZN(new_n522));
  XOR2_X1   g321(.A(new_n519), .B(KEYINPUT13), .Z(new_n523));
  NAND2_X1  g322(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  NAND2_X1  g323(.A1(new_n521), .A2(new_n524), .ZN(new_n525));
  NAND2_X1  g324(.A1(new_n525), .A2(KEYINPUT87), .ZN(new_n526));
  XNOR2_X1  g325(.A(G113gat), .B(G141gat), .ZN(new_n527));
  XNOR2_X1  g326(.A(KEYINPUT86), .B(KEYINPUT11), .ZN(new_n528));
  XNOR2_X1  g327(.A(new_n527), .B(new_n528), .ZN(new_n529));
  XOR2_X1   g328(.A(G169gat), .B(G197gat), .Z(new_n530));
  XNOR2_X1  g329(.A(new_n529), .B(new_n530), .ZN(new_n531));
  XNOR2_X1  g330(.A(new_n531), .B(KEYINPUT12), .ZN(new_n532));
  XNOR2_X1  g331(.A(new_n526), .B(new_n532), .ZN(new_n533));
  AND3_X1   g332(.A1(new_n483), .A2(new_n492), .A3(new_n533), .ZN(new_n534));
  NAND2_X1  g333(.A1(G99gat), .A2(G106gat), .ZN(new_n535));
  INV_X1    g334(.A(G85gat), .ZN(new_n536));
  AOI22_X1  g335(.A1(KEYINPUT8), .A2(new_n535), .B1(new_n536), .B2(new_n406), .ZN(new_n537));
  XNOR2_X1  g336(.A(new_n537), .B(KEYINPUT95), .ZN(new_n538));
  NAND2_X1  g337(.A1(G85gat), .A2(G92gat), .ZN(new_n539));
  XNOR2_X1  g338(.A(new_n539), .B(KEYINPUT7), .ZN(new_n540));
  NAND2_X1  g339(.A1(new_n538), .A2(new_n540), .ZN(new_n541));
  XOR2_X1   g340(.A(G99gat), .B(G106gat), .Z(new_n542));
  XNOR2_X1  g341(.A(new_n541), .B(new_n542), .ZN(new_n543));
  AND2_X1   g342(.A1(G232gat), .A2(G233gat), .ZN(new_n544));
  AOI22_X1  g343(.A1(new_n517), .A2(new_n543), .B1(KEYINPUT41), .B2(new_n544), .ZN(new_n545));
  OAI21_X1  g344(.A(new_n545), .B1(new_n507), .B2(new_n543), .ZN(new_n546));
  XOR2_X1   g345(.A(G190gat), .B(G218gat), .Z(new_n547));
  XNOR2_X1  g346(.A(new_n547), .B(KEYINPUT96), .ZN(new_n548));
  XNOR2_X1  g347(.A(new_n546), .B(new_n548), .ZN(new_n549));
  XOR2_X1   g348(.A(G134gat), .B(G162gat), .Z(new_n550));
  XNOR2_X1  g349(.A(new_n550), .B(KEYINPUT94), .ZN(new_n551));
  NOR2_X1   g350(.A1(new_n544), .A2(KEYINPUT41), .ZN(new_n552));
  XNOR2_X1  g351(.A(new_n551), .B(new_n552), .ZN(new_n553));
  OR3_X1    g352(.A1(new_n549), .A2(KEYINPUT97), .A3(new_n553), .ZN(new_n554));
  NAND2_X1  g353(.A1(new_n549), .A2(new_n553), .ZN(new_n555));
  NOR2_X1   g354(.A1(new_n546), .A2(new_n548), .ZN(new_n556));
  NAND2_X1  g355(.A1(new_n556), .A2(KEYINPUT97), .ZN(new_n557));
  NAND3_X1  g356(.A1(new_n554), .A2(new_n555), .A3(new_n557), .ZN(new_n558));
  XNOR2_X1  g357(.A(G57gat), .B(G64gat), .ZN(new_n559));
  AOI21_X1  g358(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n560));
  OR3_X1    g359(.A1(new_n559), .A2(KEYINPUT92), .A3(new_n560), .ZN(new_n561));
  XNOR2_X1  g360(.A(G71gat), .B(G78gat), .ZN(new_n562));
  XOR2_X1   g361(.A(new_n561), .B(new_n562), .Z(new_n563));
  INV_X1    g362(.A(new_n563), .ZN(new_n564));
  AOI21_X1  g363(.A(new_n514), .B1(new_n564), .B2(KEYINPUT21), .ZN(new_n565));
  XNOR2_X1  g364(.A(new_n565), .B(G183gat), .ZN(new_n566));
  XNOR2_X1  g365(.A(KEYINPUT93), .B(KEYINPUT21), .ZN(new_n567));
  NOR2_X1   g366(.A1(new_n564), .A2(new_n567), .ZN(new_n568));
  XNOR2_X1  g367(.A(new_n566), .B(new_n568), .ZN(new_n569));
  XNOR2_X1  g368(.A(G127gat), .B(G155gat), .ZN(new_n570));
  XNOR2_X1  g369(.A(new_n570), .B(G211gat), .ZN(new_n571));
  XNOR2_X1  g370(.A(new_n569), .B(new_n571), .ZN(new_n572));
  XOR2_X1   g371(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n573));
  NAND2_X1  g372(.A1(G231gat), .A2(G233gat), .ZN(new_n574));
  XNOR2_X1  g373(.A(new_n573), .B(new_n574), .ZN(new_n575));
  XNOR2_X1  g374(.A(new_n572), .B(new_n575), .ZN(new_n576));
  NAND2_X1  g375(.A1(new_n558), .A2(new_n576), .ZN(new_n577));
  XNOR2_X1  g376(.A(G120gat), .B(G148gat), .ZN(new_n578));
  INV_X1    g377(.A(G176gat), .ZN(new_n579));
  XNOR2_X1  g378(.A(new_n578), .B(new_n579), .ZN(new_n580));
  INV_X1    g379(.A(G204gat), .ZN(new_n581));
  XNOR2_X1  g380(.A(new_n580), .B(new_n581), .ZN(new_n582));
  OR2_X1    g381(.A1(new_n541), .A2(new_n542), .ZN(new_n583));
  AOI21_X1  g382(.A(new_n563), .B1(new_n583), .B2(KEYINPUT98), .ZN(new_n584));
  XNOR2_X1  g383(.A(new_n584), .B(new_n543), .ZN(new_n585));
  NAND2_X1  g384(.A1(G230gat), .A2(G233gat), .ZN(new_n586));
  XNOR2_X1  g385(.A(new_n586), .B(KEYINPUT99), .ZN(new_n587));
  INV_X1    g386(.A(new_n587), .ZN(new_n588));
  NOR2_X1   g387(.A1(new_n585), .A2(new_n588), .ZN(new_n589));
  INV_X1    g388(.A(new_n585), .ZN(new_n590));
  NAND2_X1  g389(.A1(new_n564), .A2(KEYINPUT10), .ZN(new_n591));
  OAI22_X1  g390(.A1(new_n590), .A2(KEYINPUT10), .B1(new_n543), .B2(new_n591), .ZN(new_n592));
  AOI211_X1 g391(.A(new_n582), .B(new_n589), .C1(new_n592), .C2(new_n588), .ZN(new_n593));
  XOR2_X1   g392(.A(new_n593), .B(KEYINPUT100), .Z(new_n594));
  XOR2_X1   g393(.A(new_n587), .B(KEYINPUT101), .Z(new_n595));
  NAND2_X1  g394(.A1(new_n592), .A2(new_n595), .ZN(new_n596));
  INV_X1    g395(.A(new_n596), .ZN(new_n597));
  OAI21_X1  g396(.A(new_n582), .B1(new_n597), .B2(new_n589), .ZN(new_n598));
  AND2_X1   g397(.A1(new_n594), .A2(new_n598), .ZN(new_n599));
  INV_X1    g398(.A(new_n599), .ZN(new_n600));
  NOR2_X1   g399(.A1(new_n577), .A2(new_n600), .ZN(new_n601));
  NAND2_X1  g400(.A1(new_n534), .A2(new_n601), .ZN(new_n602));
  NOR2_X1   g401(.A1(new_n602), .A2(new_n392), .ZN(new_n603));
  XOR2_X1   g402(.A(KEYINPUT102), .B(G1gat), .Z(new_n604));
  XNOR2_X1  g403(.A(new_n603), .B(new_n604), .ZN(G1324gat));
  XNOR2_X1  g404(.A(KEYINPUT16), .B(G8gat), .ZN(new_n606));
  INV_X1    g405(.A(KEYINPUT103), .ZN(new_n607));
  INV_X1    g406(.A(KEYINPUT42), .ZN(new_n608));
  AOI21_X1  g407(.A(new_n606), .B1(new_n607), .B2(new_n608), .ZN(new_n609));
  INV_X1    g408(.A(new_n602), .ZN(new_n610));
  INV_X1    g409(.A(new_n433), .ZN(new_n611));
  NAND2_X1  g410(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  AOI211_X1 g411(.A(new_n609), .B(new_n612), .C1(new_n607), .C2(new_n606), .ZN(new_n613));
  OR2_X1    g412(.A1(new_n612), .A2(new_n606), .ZN(new_n614));
  AOI21_X1  g413(.A(new_n608), .B1(new_n612), .B2(G8gat), .ZN(new_n615));
  AOI21_X1  g414(.A(new_n613), .B1(new_n614), .B2(new_n615), .ZN(G1325gat));
  INV_X1    g415(.A(G15gat), .ZN(new_n617));
  INV_X1    g416(.A(KEYINPUT104), .ZN(new_n618));
  INV_X1    g417(.A(new_n445), .ZN(new_n619));
  AOI21_X1  g418(.A(KEYINPUT36), .B1(new_n297), .B2(new_n302), .ZN(new_n620));
  OAI21_X1  g419(.A(new_n618), .B1(new_n619), .B2(new_n620), .ZN(new_n621));
  NAND3_X1  g420(.A1(new_n444), .A2(KEYINPUT104), .A3(new_n445), .ZN(new_n622));
  NAND2_X1  g421(.A1(new_n621), .A2(new_n622), .ZN(new_n623));
  NOR3_X1   g422(.A1(new_n602), .A2(new_n617), .A3(new_n623), .ZN(new_n624));
  NOR2_X1   g423(.A1(new_n442), .A2(new_n443), .ZN(new_n625));
  NAND2_X1  g424(.A1(new_n610), .A2(new_n625), .ZN(new_n626));
  AOI21_X1  g425(.A(new_n624), .B1(new_n617), .B2(new_n626), .ZN(G1326gat));
  NOR2_X1   g426(.A1(new_n602), .A2(new_n350), .ZN(new_n628));
  XOR2_X1   g427(.A(KEYINPUT43), .B(G22gat), .Z(new_n629));
  XNOR2_X1  g428(.A(new_n629), .B(KEYINPUT105), .ZN(new_n630));
  XNOR2_X1  g429(.A(new_n628), .B(new_n630), .ZN(G1327gat));
  INV_X1    g430(.A(new_n558), .ZN(new_n632));
  NOR2_X1   g431(.A1(new_n600), .A2(new_n576), .ZN(new_n633));
  AND3_X1   g432(.A1(new_n534), .A2(new_n632), .A3(new_n633), .ZN(new_n634));
  INV_X1    g433(.A(G29gat), .ZN(new_n635));
  NAND3_X1  g434(.A1(new_n634), .A2(new_n635), .A3(new_n448), .ZN(new_n636));
  XNOR2_X1  g435(.A(new_n636), .B(KEYINPUT45), .ZN(new_n637));
  INV_X1    g436(.A(KEYINPUT44), .ZN(new_n638));
  AOI22_X1  g437(.A1(new_n484), .A2(new_n485), .B1(new_n621), .B2(new_n622), .ZN(new_n639));
  NAND2_X1  g438(.A1(new_n355), .A2(new_n436), .ZN(new_n640));
  NAND2_X1  g439(.A1(new_n640), .A2(KEYINPUT35), .ZN(new_n641));
  AOI22_X1  g440(.A1(new_n639), .A2(new_n440), .B1(new_n641), .B2(new_n488), .ZN(new_n642));
  OAI21_X1  g441(.A(new_n638), .B1(new_n642), .B2(new_n558), .ZN(new_n643));
  NOR2_X1   g442(.A1(new_n558), .A2(new_n638), .ZN(new_n644));
  NAND3_X1  g443(.A1(new_n483), .A2(new_n492), .A3(new_n644), .ZN(new_n645));
  AND2_X1   g444(.A1(new_n643), .A2(new_n645), .ZN(new_n646));
  NAND3_X1  g445(.A1(new_n646), .A2(new_n533), .A3(new_n633), .ZN(new_n647));
  OAI21_X1  g446(.A(G29gat), .B1(new_n647), .B2(new_n392), .ZN(new_n648));
  NAND2_X1  g447(.A1(new_n637), .A2(new_n648), .ZN(G1328gat));
  INV_X1    g448(.A(new_n495), .ZN(new_n650));
  NAND3_X1  g449(.A1(new_n634), .A2(new_n611), .A3(new_n650), .ZN(new_n651));
  XOR2_X1   g450(.A(new_n651), .B(KEYINPUT46), .Z(new_n652));
  OAI21_X1  g451(.A(new_n495), .B1(new_n647), .B2(new_n433), .ZN(new_n653));
  NAND2_X1  g452(.A1(new_n652), .A2(new_n653), .ZN(G1329gat));
  AOI21_X1  g453(.A(G43gat), .B1(new_n634), .B2(new_n625), .ZN(new_n655));
  INV_X1    g454(.A(new_n623), .ZN(new_n656));
  INV_X1    g455(.A(G43gat), .ZN(new_n657));
  NOR2_X1   g456(.A1(new_n647), .A2(new_n657), .ZN(new_n658));
  AOI21_X1  g457(.A(new_n655), .B1(new_n656), .B2(new_n658), .ZN(new_n659));
  XOR2_X1   g458(.A(new_n659), .B(KEYINPUT47), .Z(G1330gat));
  OAI21_X1  g459(.A(G50gat), .B1(new_n647), .B2(new_n350), .ZN(new_n661));
  NAND3_X1  g460(.A1(new_n634), .A2(new_n305), .A3(new_n439), .ZN(new_n662));
  NAND3_X1  g461(.A1(new_n661), .A2(KEYINPUT48), .A3(new_n662), .ZN(new_n663));
  XNOR2_X1  g462(.A(new_n663), .B(KEYINPUT107), .ZN(new_n664));
  OR2_X1    g463(.A1(new_n662), .A2(KEYINPUT106), .ZN(new_n665));
  NAND2_X1  g464(.A1(new_n662), .A2(KEYINPUT106), .ZN(new_n666));
  AND3_X1   g465(.A1(new_n665), .A2(new_n661), .A3(new_n666), .ZN(new_n667));
  OAI21_X1  g466(.A(new_n664), .B1(KEYINPUT48), .B2(new_n667), .ZN(G1331gat));
  NAND3_X1  g467(.A1(new_n486), .A2(new_n623), .A3(new_n440), .ZN(new_n669));
  NAND2_X1  g468(.A1(new_n669), .A2(new_n490), .ZN(new_n670));
  NOR2_X1   g469(.A1(new_n577), .A2(new_n533), .ZN(new_n671));
  NAND3_X1  g470(.A1(new_n670), .A2(new_n600), .A3(new_n671), .ZN(new_n672));
  OR2_X1    g471(.A1(new_n672), .A2(KEYINPUT108), .ZN(new_n673));
  NAND2_X1  g472(.A1(new_n672), .A2(KEYINPUT108), .ZN(new_n674));
  NAND2_X1  g473(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  INV_X1    g474(.A(new_n675), .ZN(new_n676));
  NAND2_X1  g475(.A1(new_n676), .A2(new_n448), .ZN(new_n677));
  XNOR2_X1  g476(.A(new_n677), .B(G57gat), .ZN(G1332gat));
  NOR2_X1   g477(.A1(new_n675), .A2(new_n433), .ZN(new_n679));
  NOR2_X1   g478(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n680));
  AND2_X1   g479(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n681));
  OAI21_X1  g480(.A(new_n679), .B1(new_n680), .B2(new_n681), .ZN(new_n682));
  OAI21_X1  g481(.A(new_n682), .B1(new_n679), .B2(new_n680), .ZN(G1333gat));
  INV_X1    g482(.A(G71gat), .ZN(new_n684));
  NOR3_X1   g483(.A1(new_n675), .A2(new_n684), .A3(new_n623), .ZN(new_n685));
  XNOR2_X1  g484(.A(new_n685), .B(KEYINPUT109), .ZN(new_n686));
  INV_X1    g485(.A(new_n625), .ZN(new_n687));
  OAI21_X1  g486(.A(new_n684), .B1(new_n675), .B2(new_n687), .ZN(new_n688));
  NAND2_X1  g487(.A1(new_n686), .A2(new_n688), .ZN(new_n689));
  XNOR2_X1  g488(.A(new_n689), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g489(.A1(new_n676), .A2(new_n439), .ZN(new_n691));
  XNOR2_X1  g490(.A(new_n691), .B(G78gat), .ZN(G1335gat));
  INV_X1    g491(.A(KEYINPUT111), .ZN(new_n693));
  OAI21_X1  g492(.A(new_n693), .B1(new_n642), .B2(new_n558), .ZN(new_n694));
  NAND3_X1  g493(.A1(new_n670), .A2(KEYINPUT111), .A3(new_n632), .ZN(new_n695));
  NOR2_X1   g494(.A1(new_n533), .A2(new_n576), .ZN(new_n696));
  NAND3_X1  g495(.A1(new_n694), .A2(new_n695), .A3(new_n696), .ZN(new_n697));
  NAND2_X1  g496(.A1(new_n697), .A2(KEYINPUT51), .ZN(new_n698));
  INV_X1    g497(.A(KEYINPUT51), .ZN(new_n699));
  NAND4_X1  g498(.A1(new_n694), .A2(new_n699), .A3(new_n695), .A4(new_n696), .ZN(new_n700));
  NAND3_X1  g499(.A1(new_n698), .A2(new_n600), .A3(new_n700), .ZN(new_n701));
  OR2_X1    g500(.A1(new_n701), .A2(new_n392), .ZN(new_n702));
  NOR3_X1   g501(.A1(new_n533), .A2(new_n576), .A3(new_n599), .ZN(new_n703));
  NAND3_X1  g502(.A1(new_n643), .A2(new_n645), .A3(new_n703), .ZN(new_n704));
  INV_X1    g503(.A(KEYINPUT110), .ZN(new_n705));
  NAND2_X1  g504(.A1(new_n704), .A2(new_n705), .ZN(new_n706));
  NAND4_X1  g505(.A1(new_n643), .A2(new_n645), .A3(new_n703), .A4(KEYINPUT110), .ZN(new_n707));
  AOI21_X1  g506(.A(new_n536), .B1(new_n706), .B2(new_n707), .ZN(new_n708));
  AOI22_X1  g507(.A1(new_n702), .A2(new_n536), .B1(new_n448), .B2(new_n708), .ZN(G1336gat));
  NOR2_X1   g508(.A1(new_n433), .A2(G92gat), .ZN(new_n710));
  NAND4_X1  g509(.A1(new_n698), .A2(new_n700), .A3(new_n600), .A4(new_n710), .ZN(new_n711));
  INV_X1    g510(.A(KEYINPUT52), .ZN(new_n712));
  OAI21_X1  g511(.A(G92gat), .B1(new_n704), .B2(new_n433), .ZN(new_n713));
  NAND3_X1  g512(.A1(new_n711), .A2(new_n712), .A3(new_n713), .ZN(new_n714));
  AOI21_X1  g513(.A(new_n433), .B1(new_n706), .B2(new_n707), .ZN(new_n715));
  OAI21_X1  g514(.A(new_n711), .B1(new_n715), .B2(new_n406), .ZN(new_n716));
  INV_X1    g515(.A(KEYINPUT112), .ZN(new_n717));
  AND3_X1   g516(.A1(new_n716), .A2(new_n717), .A3(KEYINPUT52), .ZN(new_n718));
  AOI21_X1  g517(.A(new_n717), .B1(new_n716), .B2(KEYINPUT52), .ZN(new_n719));
  OAI21_X1  g518(.A(new_n714), .B1(new_n718), .B2(new_n719), .ZN(new_n720));
  INV_X1    g519(.A(KEYINPUT113), .ZN(new_n721));
  NAND2_X1  g520(.A1(new_n720), .A2(new_n721), .ZN(new_n722));
  OAI211_X1 g521(.A(KEYINPUT113), .B(new_n714), .C1(new_n718), .C2(new_n719), .ZN(new_n723));
  NAND2_X1  g522(.A1(new_n722), .A2(new_n723), .ZN(G1337gat));
  OAI21_X1  g523(.A(new_n282), .B1(new_n701), .B2(new_n687), .ZN(new_n725));
  NAND2_X1  g524(.A1(new_n706), .A2(new_n707), .ZN(new_n726));
  NAND3_X1  g525(.A1(new_n726), .A2(G99gat), .A3(new_n656), .ZN(new_n727));
  NAND2_X1  g526(.A1(new_n725), .A2(new_n727), .ZN(new_n728));
  XNOR2_X1  g527(.A(new_n728), .B(KEYINPUT114), .ZN(G1338gat));
  NAND3_X1  g528(.A1(new_n646), .A2(new_n439), .A3(new_n703), .ZN(new_n730));
  AOI21_X1  g529(.A(KEYINPUT53), .B1(new_n730), .B2(G106gat), .ZN(new_n731));
  NAND4_X1  g530(.A1(new_n698), .A2(new_n700), .A3(new_n439), .A4(new_n600), .ZN(new_n732));
  OAI21_X1  g531(.A(new_n731), .B1(G106gat), .B2(new_n732), .ZN(new_n733));
  INV_X1    g532(.A(new_n726), .ZN(new_n734));
  OAI21_X1  g533(.A(G106gat), .B1(new_n734), .B2(new_n350), .ZN(new_n735));
  OAI21_X1  g534(.A(new_n735), .B1(G106gat), .B2(new_n732), .ZN(new_n736));
  NAND3_X1  g535(.A1(new_n736), .A2(KEYINPUT115), .A3(KEYINPUT53), .ZN(new_n737));
  INV_X1    g536(.A(new_n737), .ZN(new_n738));
  AOI21_X1  g537(.A(KEYINPUT115), .B1(new_n736), .B2(KEYINPUT53), .ZN(new_n739));
  OAI21_X1  g538(.A(new_n733), .B1(new_n738), .B2(new_n739), .ZN(G1339gat));
  NOR3_X1   g539(.A1(new_n577), .A2(new_n533), .A3(new_n600), .ZN(new_n741));
  NAND2_X1  g540(.A1(new_n592), .A2(new_n588), .ZN(new_n742));
  OAI211_X1 g541(.A(new_n742), .B(KEYINPUT54), .C1(new_n592), .C2(new_n595), .ZN(new_n743));
  OAI211_X1 g542(.A(new_n743), .B(new_n582), .C1(KEYINPUT54), .C2(new_n596), .ZN(new_n744));
  XNOR2_X1  g543(.A(new_n744), .B(KEYINPUT55), .ZN(new_n745));
  NAND2_X1  g544(.A1(new_n745), .A2(new_n594), .ZN(new_n746));
  NOR2_X1   g545(.A1(new_n518), .A2(new_n519), .ZN(new_n747));
  NOR2_X1   g546(.A1(new_n522), .A2(new_n523), .ZN(new_n748));
  OAI21_X1  g547(.A(new_n531), .B1(new_n747), .B2(new_n748), .ZN(new_n749));
  INV_X1    g548(.A(new_n532), .ZN(new_n750));
  OAI21_X1  g549(.A(new_n749), .B1(new_n525), .B2(new_n750), .ZN(new_n751));
  NOR3_X1   g550(.A1(new_n746), .A2(new_n558), .A3(new_n751), .ZN(new_n752));
  XNOR2_X1  g551(.A(new_n752), .B(KEYINPUT116), .ZN(new_n753));
  AND2_X1   g552(.A1(new_n745), .A2(new_n594), .ZN(new_n754));
  NAND2_X1  g553(.A1(new_n754), .A2(new_n533), .ZN(new_n755));
  OR2_X1    g554(.A1(new_n599), .A2(new_n751), .ZN(new_n756));
  NAND2_X1  g555(.A1(new_n755), .A2(new_n756), .ZN(new_n757));
  NAND2_X1  g556(.A1(new_n757), .A2(new_n558), .ZN(new_n758));
  NAND2_X1  g557(.A1(new_n753), .A2(new_n758), .ZN(new_n759));
  INV_X1    g558(.A(new_n576), .ZN(new_n760));
  AOI21_X1  g559(.A(new_n741), .B1(new_n759), .B2(new_n760), .ZN(new_n761));
  NOR2_X1   g560(.A1(new_n611), .A2(new_n392), .ZN(new_n762));
  INV_X1    g561(.A(new_n762), .ZN(new_n763));
  NOR3_X1   g562(.A1(new_n761), .A2(new_n351), .A3(new_n763), .ZN(new_n764));
  AOI21_X1  g563(.A(new_n254), .B1(new_n764), .B2(new_n533), .ZN(new_n765));
  XOR2_X1   g564(.A(new_n765), .B(KEYINPUT117), .Z(new_n766));
  INV_X1    g565(.A(new_n355), .ZN(new_n767));
  NOR3_X1   g566(.A1(new_n761), .A2(new_n767), .A3(new_n763), .ZN(new_n768));
  NAND3_X1  g567(.A1(new_n768), .A2(new_n254), .A3(new_n533), .ZN(new_n769));
  NAND2_X1  g568(.A1(new_n766), .A2(new_n769), .ZN(G1340gat));
  AOI21_X1  g569(.A(new_n255), .B1(new_n764), .B2(new_n600), .ZN(new_n771));
  XNOR2_X1  g570(.A(new_n771), .B(KEYINPUT118), .ZN(new_n772));
  NAND3_X1  g571(.A1(new_n768), .A2(new_n255), .A3(new_n600), .ZN(new_n773));
  NAND2_X1  g572(.A1(new_n772), .A2(new_n773), .ZN(G1341gat));
  AOI21_X1  g573(.A(G127gat), .B1(new_n768), .B2(new_n576), .ZN(new_n775));
  NOR2_X1   g574(.A1(new_n760), .A2(new_n260), .ZN(new_n776));
  AOI21_X1  g575(.A(new_n775), .B1(new_n764), .B2(new_n776), .ZN(G1342gat));
  NAND3_X1  g576(.A1(new_n768), .A2(new_n253), .A3(new_n632), .ZN(new_n778));
  OR2_X1    g577(.A1(new_n778), .A2(KEYINPUT56), .ZN(new_n779));
  INV_X1    g578(.A(new_n764), .ZN(new_n780));
  OAI21_X1  g579(.A(G134gat), .B1(new_n780), .B2(new_n558), .ZN(new_n781));
  NAND2_X1  g580(.A1(new_n778), .A2(KEYINPUT56), .ZN(new_n782));
  NAND3_X1  g581(.A1(new_n779), .A2(new_n781), .A3(new_n782), .ZN(new_n783));
  INV_X1    g582(.A(KEYINPUT119), .ZN(new_n784));
  XNOR2_X1  g583(.A(new_n783), .B(new_n784), .ZN(G1343gat));
  AOI21_X1  g584(.A(new_n576), .B1(new_n753), .B2(new_n758), .ZN(new_n786));
  OAI21_X1  g585(.A(new_n439), .B1(new_n786), .B2(new_n741), .ZN(new_n787));
  OR2_X1    g586(.A1(new_n787), .A2(KEYINPUT57), .ZN(new_n788));
  NAND2_X1  g587(.A1(new_n787), .A2(KEYINPUT57), .ZN(new_n789));
  NOR2_X1   g588(.A1(new_n656), .A2(new_n763), .ZN(new_n790));
  NAND3_X1  g589(.A1(new_n788), .A2(new_n789), .A3(new_n790), .ZN(new_n791));
  INV_X1    g590(.A(new_n533), .ZN(new_n792));
  OAI21_X1  g591(.A(G141gat), .B1(new_n791), .B2(new_n792), .ZN(new_n793));
  NOR3_X1   g592(.A1(new_n787), .A2(new_n656), .A3(new_n763), .ZN(new_n794));
  INV_X1    g593(.A(G141gat), .ZN(new_n795));
  NAND3_X1  g594(.A1(new_n794), .A2(new_n795), .A3(new_n533), .ZN(new_n796));
  NAND2_X1  g595(.A1(new_n793), .A2(new_n796), .ZN(new_n797));
  XNOR2_X1  g596(.A(new_n797), .B(KEYINPUT58), .ZN(G1344gat));
  INV_X1    g597(.A(G148gat), .ZN(new_n799));
  NAND3_X1  g598(.A1(new_n794), .A2(new_n799), .A3(new_n600), .ZN(new_n800));
  INV_X1    g599(.A(KEYINPUT59), .ZN(new_n801));
  OAI21_X1  g600(.A(new_n801), .B1(new_n791), .B2(new_n599), .ZN(new_n802));
  NOR2_X1   g601(.A1(new_n802), .A2(new_n799), .ZN(new_n803));
  INV_X1    g602(.A(KEYINPUT57), .ZN(new_n804));
  INV_X1    g603(.A(new_n752), .ZN(new_n805));
  AOI21_X1  g604(.A(new_n576), .B1(new_n758), .B2(new_n805), .ZN(new_n806));
  OAI211_X1 g605(.A(new_n804), .B(new_n439), .C1(new_n806), .C2(new_n741), .ZN(new_n807));
  INV_X1    g606(.A(new_n807), .ZN(new_n808));
  AOI21_X1  g607(.A(new_n808), .B1(KEYINPUT57), .B2(new_n787), .ZN(new_n809));
  NAND3_X1  g608(.A1(new_n809), .A2(new_n600), .A3(new_n790), .ZN(new_n810));
  AOI21_X1  g609(.A(new_n801), .B1(new_n810), .B2(G148gat), .ZN(new_n811));
  OAI21_X1  g610(.A(new_n800), .B1(new_n803), .B2(new_n811), .ZN(G1345gat));
  AOI21_X1  g611(.A(G155gat), .B1(new_n794), .B2(new_n576), .ZN(new_n813));
  NOR2_X1   g612(.A1(new_n791), .A2(new_n311), .ZN(new_n814));
  AOI21_X1  g613(.A(new_n813), .B1(new_n814), .B2(new_n576), .ZN(G1346gat));
  AOI21_X1  g614(.A(G162gat), .B1(new_n794), .B2(new_n632), .ZN(new_n816));
  NOR2_X1   g615(.A1(new_n791), .A2(new_n312), .ZN(new_n817));
  AOI21_X1  g616(.A(new_n816), .B1(new_n817), .B2(new_n632), .ZN(G1347gat));
  NOR2_X1   g617(.A1(new_n433), .A2(new_n448), .ZN(new_n819));
  XNOR2_X1  g618(.A(new_n819), .B(KEYINPUT121), .ZN(new_n820));
  OR3_X1    g619(.A1(new_n761), .A2(new_n351), .A3(new_n820), .ZN(new_n821));
  OAI21_X1  g620(.A(G169gat), .B1(new_n821), .B2(new_n792), .ZN(new_n822));
  NOR2_X1   g621(.A1(new_n767), .A2(new_n433), .ZN(new_n823));
  NOR2_X1   g622(.A1(new_n823), .A2(KEYINPUT120), .ZN(new_n824));
  AND2_X1   g623(.A1(new_n823), .A2(KEYINPUT120), .ZN(new_n825));
  NOR4_X1   g624(.A1(new_n761), .A2(new_n448), .A3(new_n824), .A4(new_n825), .ZN(new_n826));
  INV_X1    g625(.A(G169gat), .ZN(new_n827));
  NAND3_X1  g626(.A1(new_n826), .A2(new_n827), .A3(new_n533), .ZN(new_n828));
  NAND2_X1  g627(.A1(new_n822), .A2(new_n828), .ZN(G1348gat));
  NOR3_X1   g628(.A1(new_n821), .A2(new_n579), .A3(new_n599), .ZN(new_n830));
  AOI21_X1  g629(.A(G176gat), .B1(new_n826), .B2(new_n600), .ZN(new_n831));
  NOR2_X1   g630(.A1(new_n830), .A2(new_n831), .ZN(G1349gat));
  OAI21_X1  g631(.A(G183gat), .B1(new_n821), .B2(new_n760), .ZN(new_n833));
  NAND3_X1  g632(.A1(new_n826), .A2(new_n242), .A3(new_n576), .ZN(new_n834));
  NAND2_X1  g633(.A1(new_n833), .A2(new_n834), .ZN(new_n835));
  INV_X1    g634(.A(KEYINPUT60), .ZN(new_n836));
  NOR2_X1   g635(.A1(new_n836), .A2(KEYINPUT122), .ZN(new_n837));
  XNOR2_X1  g636(.A(new_n835), .B(new_n837), .ZN(G1350gat));
  OAI21_X1  g637(.A(G190gat), .B1(new_n821), .B2(new_n558), .ZN(new_n839));
  XNOR2_X1  g638(.A(new_n839), .B(KEYINPUT61), .ZN(new_n840));
  NAND3_X1  g639(.A1(new_n826), .A2(new_n218), .A3(new_n632), .ZN(new_n841));
  NAND2_X1  g640(.A1(new_n840), .A2(new_n841), .ZN(G1351gat));
  NOR2_X1   g641(.A1(new_n656), .A2(new_n820), .ZN(new_n843));
  NAND4_X1  g642(.A1(new_n789), .A2(new_n533), .A3(new_n807), .A4(new_n843), .ZN(new_n844));
  INV_X1    g643(.A(KEYINPUT123), .ZN(new_n845));
  NAND2_X1  g644(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  NAND4_X1  g645(.A1(new_n809), .A2(KEYINPUT123), .A3(new_n533), .A4(new_n843), .ZN(new_n847));
  NAND3_X1  g646(.A1(new_n846), .A2(new_n847), .A3(G197gat), .ZN(new_n848));
  NOR2_X1   g647(.A1(new_n787), .A2(new_n656), .ZN(new_n849));
  AND2_X1   g648(.A1(new_n849), .A2(new_n819), .ZN(new_n850));
  INV_X1    g649(.A(G197gat), .ZN(new_n851));
  NAND3_X1  g650(.A1(new_n850), .A2(new_n851), .A3(new_n533), .ZN(new_n852));
  NAND2_X1  g651(.A1(new_n848), .A2(new_n852), .ZN(new_n853));
  NAND2_X1  g652(.A1(new_n853), .A2(KEYINPUT124), .ZN(new_n854));
  INV_X1    g653(.A(KEYINPUT124), .ZN(new_n855));
  NAND3_X1  g654(.A1(new_n848), .A2(new_n855), .A3(new_n852), .ZN(new_n856));
  NAND2_X1  g655(.A1(new_n854), .A2(new_n856), .ZN(G1352gat));
  NAND3_X1  g656(.A1(new_n849), .A2(new_n581), .A3(new_n819), .ZN(new_n858));
  XNOR2_X1  g657(.A(KEYINPUT125), .B(KEYINPUT62), .ZN(new_n859));
  OR3_X1    g658(.A1(new_n858), .A2(new_n599), .A3(new_n859), .ZN(new_n860));
  NAND3_X1  g659(.A1(new_n809), .A2(new_n600), .A3(new_n843), .ZN(new_n861));
  NAND2_X1  g660(.A1(new_n861), .A2(G204gat), .ZN(new_n862));
  OAI21_X1  g661(.A(new_n859), .B1(new_n858), .B2(new_n599), .ZN(new_n863));
  NAND3_X1  g662(.A1(new_n860), .A2(new_n862), .A3(new_n863), .ZN(new_n864));
  NAND2_X1  g663(.A1(new_n864), .A2(KEYINPUT126), .ZN(new_n865));
  INV_X1    g664(.A(KEYINPUT126), .ZN(new_n866));
  NAND4_X1  g665(.A1(new_n860), .A2(new_n862), .A3(new_n866), .A4(new_n863), .ZN(new_n867));
  NAND2_X1  g666(.A1(new_n865), .A2(new_n867), .ZN(G1353gat));
  NAND3_X1  g667(.A1(new_n850), .A2(new_n323), .A3(new_n576), .ZN(new_n869));
  NAND3_X1  g668(.A1(new_n809), .A2(new_n576), .A3(new_n843), .ZN(new_n870));
  AND3_X1   g669(.A1(new_n870), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n871));
  AOI21_X1  g670(.A(KEYINPUT63), .B1(new_n870), .B2(G211gat), .ZN(new_n872));
  OAI21_X1  g671(.A(new_n869), .B1(new_n871), .B2(new_n872), .ZN(G1354gat));
  NAND3_X1  g672(.A1(new_n850), .A2(new_n324), .A3(new_n632), .ZN(new_n874));
  NAND2_X1  g673(.A1(new_n789), .A2(new_n807), .ZN(new_n875));
  INV_X1    g674(.A(new_n843), .ZN(new_n876));
  NOR3_X1   g675(.A1(new_n875), .A2(KEYINPUT127), .A3(new_n876), .ZN(new_n877));
  INV_X1    g676(.A(KEYINPUT127), .ZN(new_n878));
  AOI21_X1  g677(.A(new_n878), .B1(new_n809), .B2(new_n843), .ZN(new_n879));
  NOR3_X1   g678(.A1(new_n877), .A2(new_n879), .A3(new_n558), .ZN(new_n880));
  OAI21_X1  g679(.A(new_n874), .B1(new_n880), .B2(new_n324), .ZN(G1355gat));
endmodule


