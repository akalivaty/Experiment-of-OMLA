//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 1 1 1 1 0 0 1 0 1 1 1 1 1 0 1 1 1 1 0 1 1 1 0 1 1 1 1 0 0 1 1 1 0 0 0 0 1 0 0 0 1 1 1 0 1 1 1 1 1 1 0 0 1 0 0 0 1 0 1 0 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:21:39 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n718, new_n719, new_n720, new_n721, new_n722, new_n723, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n744, new_n745, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n780, new_n781, new_n782, new_n783, new_n784, new_n785,
    new_n786, new_n787, new_n788, new_n789, new_n790, new_n791, new_n792,
    new_n793, new_n794, new_n795, new_n796, new_n797, new_n798, new_n799,
    new_n800, new_n801, new_n802, new_n803, new_n804, new_n805, new_n806,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n829,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n994,
    new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1027, new_n1028,
    new_n1029, new_n1030, new_n1031, new_n1032, new_n1034, new_n1035,
    new_n1036, new_n1037, new_n1038, new_n1039, new_n1040, new_n1041,
    new_n1042, new_n1043, new_n1044, new_n1045, new_n1046, new_n1048,
    new_n1049, new_n1050, new_n1051, new_n1052, new_n1053, new_n1055,
    new_n1056, new_n1057, new_n1058, new_n1059, new_n1060, new_n1061,
    new_n1062, new_n1063, new_n1064, new_n1065, new_n1066, new_n1067,
    new_n1068, new_n1069, new_n1070, new_n1071, new_n1072, new_n1073,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084;
  OAI21_X1  g000(.A(G214), .B1(G237), .B2(G902), .ZN(new_n187));
  INV_X1    g001(.A(G119), .ZN(new_n188));
  NAND2_X1  g002(.A1(new_n188), .A2(G116), .ZN(new_n189));
  INV_X1    g003(.A(G116), .ZN(new_n190));
  NAND2_X1  g004(.A1(new_n190), .A2(G119), .ZN(new_n191));
  INV_X1    g005(.A(G113), .ZN(new_n192));
  AND2_X1   g006(.A1(new_n192), .A2(KEYINPUT2), .ZN(new_n193));
  NOR2_X1   g007(.A1(new_n192), .A2(KEYINPUT2), .ZN(new_n194));
  OAI211_X1 g008(.A(new_n189), .B(new_n191), .C1(new_n193), .C2(new_n194), .ZN(new_n195));
  AND3_X1   g009(.A1(new_n189), .A2(new_n191), .A3(KEYINPUT5), .ZN(new_n196));
  OAI21_X1  g010(.A(G113), .B1(new_n189), .B2(KEYINPUT5), .ZN(new_n197));
  OAI21_X1  g011(.A(new_n195), .B1(new_n196), .B2(new_n197), .ZN(new_n198));
  INV_X1    g012(.A(G104), .ZN(new_n199));
  OAI21_X1  g013(.A(KEYINPUT3), .B1(new_n199), .B2(G107), .ZN(new_n200));
  INV_X1    g014(.A(KEYINPUT3), .ZN(new_n201));
  INV_X1    g015(.A(G107), .ZN(new_n202));
  NAND3_X1  g016(.A1(new_n201), .A2(new_n202), .A3(G104), .ZN(new_n203));
  INV_X1    g017(.A(G101), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n199), .A2(G107), .ZN(new_n205));
  NAND4_X1  g019(.A1(new_n200), .A2(new_n203), .A3(new_n204), .A4(new_n205), .ZN(new_n206));
  NOR2_X1   g020(.A1(new_n199), .A2(G107), .ZN(new_n207));
  NOR2_X1   g021(.A1(new_n202), .A2(G104), .ZN(new_n208));
  OAI21_X1  g022(.A(G101), .B1(new_n207), .B2(new_n208), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n206), .A2(new_n209), .ZN(new_n210));
  OR2_X1    g024(.A1(new_n198), .A2(new_n210), .ZN(new_n211));
  NAND3_X1  g025(.A1(new_n200), .A2(new_n203), .A3(new_n205), .ZN(new_n212));
  INV_X1    g026(.A(KEYINPUT79), .ZN(new_n213));
  AND3_X1   g027(.A1(new_n212), .A2(new_n213), .A3(G101), .ZN(new_n214));
  AOI21_X1  g028(.A(new_n213), .B1(new_n212), .B2(G101), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n206), .A2(KEYINPUT4), .ZN(new_n216));
  NOR3_X1   g030(.A1(new_n214), .A2(new_n215), .A3(new_n216), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n189), .A2(new_n191), .ZN(new_n218));
  XNOR2_X1  g032(.A(KEYINPUT2), .B(G113), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n218), .A2(new_n219), .ZN(new_n220));
  NAND3_X1  g034(.A1(new_n195), .A2(new_n220), .A3(KEYINPUT67), .ZN(new_n221));
  INV_X1    g035(.A(KEYINPUT67), .ZN(new_n222));
  NAND3_X1  g036(.A1(new_n218), .A2(new_n219), .A3(new_n222), .ZN(new_n223));
  INV_X1    g037(.A(KEYINPUT4), .ZN(new_n224));
  NAND3_X1  g038(.A1(new_n212), .A2(new_n224), .A3(G101), .ZN(new_n225));
  NAND3_X1  g039(.A1(new_n221), .A2(new_n223), .A3(new_n225), .ZN(new_n226));
  OAI21_X1  g040(.A(new_n211), .B1(new_n217), .B2(new_n226), .ZN(new_n227));
  XNOR2_X1  g041(.A(G110), .B(G122), .ZN(new_n228));
  INV_X1    g042(.A(new_n228), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n227), .A2(new_n229), .ZN(new_n230));
  OAI211_X1 g044(.A(new_n211), .B(new_n228), .C1(new_n217), .C2(new_n226), .ZN(new_n231));
  NAND3_X1  g045(.A1(new_n230), .A2(KEYINPUT6), .A3(new_n231), .ZN(new_n232));
  INV_X1    g046(.A(G146), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n233), .A2(G143), .ZN(new_n234));
  INV_X1    g048(.A(G143), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n235), .A2(G146), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n234), .A2(new_n236), .ZN(new_n237));
  AND2_X1   g051(.A1(KEYINPUT0), .A2(G128), .ZN(new_n238));
  INV_X1    g052(.A(new_n238), .ZN(new_n239));
  INV_X1    g053(.A(KEYINPUT64), .ZN(new_n240));
  OAI21_X1  g054(.A(new_n240), .B1(KEYINPUT0), .B2(G128), .ZN(new_n241));
  NOR2_X1   g055(.A1(KEYINPUT0), .A2(G128), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n242), .A2(KEYINPUT64), .ZN(new_n243));
  NAND4_X1  g057(.A1(new_n237), .A2(new_n239), .A3(new_n241), .A4(new_n243), .ZN(new_n244));
  XNOR2_X1  g058(.A(G143), .B(G146), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n245), .A2(new_n238), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n244), .A2(new_n246), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n247), .A2(G125), .ZN(new_n248));
  OAI21_X1  g062(.A(KEYINPUT1), .B1(new_n235), .B2(G146), .ZN(new_n249));
  NOR2_X1   g063(.A1(new_n235), .A2(G146), .ZN(new_n250));
  NOR2_X1   g064(.A1(new_n233), .A2(G143), .ZN(new_n251));
  OAI211_X1 g065(.A(G128), .B(new_n249), .C1(new_n250), .C2(new_n251), .ZN(new_n252));
  INV_X1    g066(.A(G128), .ZN(new_n253));
  OAI211_X1 g067(.A(new_n234), .B(new_n236), .C1(KEYINPUT1), .C2(new_n253), .ZN(new_n254));
  AOI21_X1  g068(.A(G125), .B1(new_n252), .B2(new_n254), .ZN(new_n255));
  INV_X1    g069(.A(new_n255), .ZN(new_n256));
  INV_X1    g070(.A(G953), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n257), .A2(G224), .ZN(new_n258));
  NAND3_X1  g072(.A1(new_n248), .A2(new_n256), .A3(new_n258), .ZN(new_n259));
  INV_X1    g073(.A(G125), .ZN(new_n260));
  AOI21_X1  g074(.A(new_n260), .B1(new_n244), .B2(new_n246), .ZN(new_n261));
  OAI211_X1 g075(.A(G224), .B(new_n257), .C1(new_n261), .C2(new_n255), .ZN(new_n262));
  AND3_X1   g076(.A1(new_n259), .A2(new_n262), .A3(KEYINPUT82), .ZN(new_n263));
  AOI21_X1  g077(.A(KEYINPUT82), .B1(new_n259), .B2(new_n262), .ZN(new_n264));
  NOR2_X1   g078(.A1(new_n263), .A2(new_n264), .ZN(new_n265));
  INV_X1    g079(.A(KEYINPUT6), .ZN(new_n266));
  NAND3_X1  g080(.A1(new_n227), .A2(new_n266), .A3(new_n229), .ZN(new_n267));
  NAND3_X1  g081(.A1(new_n232), .A2(new_n265), .A3(new_n267), .ZN(new_n268));
  INV_X1    g082(.A(KEYINPUT7), .ZN(new_n269));
  AND2_X1   g083(.A1(new_n269), .A2(KEYINPUT84), .ZN(new_n270));
  NOR2_X1   g084(.A1(new_n269), .A2(KEYINPUT84), .ZN(new_n271));
  OAI21_X1  g085(.A(new_n258), .B1(new_n270), .B2(new_n271), .ZN(new_n272));
  AOI22_X1  g086(.A1(new_n234), .A2(new_n236), .B1(new_n242), .B2(KEYINPUT64), .ZN(new_n273));
  OR2_X1    g087(.A1(KEYINPUT0), .A2(G128), .ZN(new_n274));
  AOI21_X1  g088(.A(new_n238), .B1(new_n274), .B2(new_n240), .ZN(new_n275));
  AOI22_X1  g089(.A1(new_n273), .A2(new_n275), .B1(new_n238), .B2(new_n245), .ZN(new_n276));
  OAI22_X1  g090(.A1(new_n255), .A2(KEYINPUT83), .B1(new_n276), .B2(new_n260), .ZN(new_n277));
  AND2_X1   g091(.A1(new_n255), .A2(KEYINPUT83), .ZN(new_n278));
  OAI21_X1  g092(.A(new_n272), .B1(new_n277), .B2(new_n278), .ZN(new_n279));
  NAND4_X1  g093(.A1(new_n248), .A2(new_n256), .A3(KEYINPUT7), .A4(new_n258), .ZN(new_n280));
  XNOR2_X1  g094(.A(new_n228), .B(KEYINPUT8), .ZN(new_n281));
  AND2_X1   g095(.A1(new_n198), .A2(new_n210), .ZN(new_n282));
  NOR2_X1   g096(.A1(new_n198), .A2(new_n210), .ZN(new_n283));
  OAI21_X1  g097(.A(new_n281), .B1(new_n282), .B2(new_n283), .ZN(new_n284));
  NAND4_X1  g098(.A1(new_n231), .A2(new_n279), .A3(new_n280), .A4(new_n284), .ZN(new_n285));
  INV_X1    g099(.A(G902), .ZN(new_n286));
  AND2_X1   g100(.A1(new_n285), .A2(new_n286), .ZN(new_n287));
  OAI21_X1  g101(.A(G210), .B1(G237), .B2(G902), .ZN(new_n288));
  AND3_X1   g102(.A1(new_n268), .A2(new_n287), .A3(new_n288), .ZN(new_n289));
  AOI21_X1  g103(.A(new_n288), .B1(new_n268), .B2(new_n287), .ZN(new_n290));
  OAI21_X1  g104(.A(new_n187), .B1(new_n289), .B2(new_n290), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n291), .A2(KEYINPUT85), .ZN(new_n292));
  INV_X1    g106(.A(KEYINPUT85), .ZN(new_n293));
  OAI211_X1 g107(.A(new_n293), .B(new_n187), .C1(new_n289), .C2(new_n290), .ZN(new_n294));
  AND2_X1   g108(.A1(new_n292), .A2(new_n294), .ZN(new_n295));
  INV_X1    g109(.A(KEYINPUT89), .ZN(new_n296));
  NOR2_X1   g110(.A1(G475), .A2(G902), .ZN(new_n297));
  INV_X1    g111(.A(new_n297), .ZN(new_n298));
  NOR2_X1   g112(.A1(G237), .A2(G953), .ZN(new_n299));
  AND3_X1   g113(.A1(new_n299), .A2(G143), .A3(G214), .ZN(new_n300));
  AOI21_X1  g114(.A(G143), .B1(new_n299), .B2(G214), .ZN(new_n301));
  OAI211_X1 g115(.A(KEYINPUT18), .B(G131), .C1(new_n300), .C2(new_n301), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n299), .A2(G214), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n303), .A2(new_n235), .ZN(new_n304));
  NAND3_X1  g118(.A1(new_n299), .A2(G143), .A3(G214), .ZN(new_n305));
  NAND2_X1  g119(.A1(KEYINPUT18), .A2(G131), .ZN(new_n306));
  NAND3_X1  g120(.A1(new_n304), .A2(new_n305), .A3(new_n306), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n302), .A2(new_n307), .ZN(new_n308));
  INV_X1    g122(.A(G140), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n309), .A2(G125), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n260), .A2(G140), .ZN(new_n311));
  AOI21_X1  g125(.A(new_n233), .B1(new_n310), .B2(new_n311), .ZN(new_n312));
  NAND3_X1  g126(.A1(new_n310), .A2(new_n311), .A3(new_n233), .ZN(new_n313));
  NAND2_X1  g127(.A1(new_n313), .A2(KEYINPUT75), .ZN(new_n314));
  XNOR2_X1  g128(.A(G125), .B(G140), .ZN(new_n315));
  INV_X1    g129(.A(KEYINPUT75), .ZN(new_n316));
  NAND3_X1  g130(.A1(new_n315), .A2(new_n316), .A3(new_n233), .ZN(new_n317));
  AOI21_X1  g131(.A(new_n312), .B1(new_n314), .B2(new_n317), .ZN(new_n318));
  OAI21_X1  g132(.A(KEYINPUT86), .B1(new_n308), .B2(new_n318), .ZN(new_n319));
  INV_X1    g133(.A(new_n312), .ZN(new_n320));
  AOI21_X1  g134(.A(new_n316), .B1(new_n315), .B2(new_n233), .ZN(new_n321));
  AND4_X1   g135(.A1(new_n316), .A2(new_n310), .A3(new_n311), .A4(new_n233), .ZN(new_n322));
  OAI21_X1  g136(.A(new_n320), .B1(new_n321), .B2(new_n322), .ZN(new_n323));
  INV_X1    g137(.A(KEYINPUT86), .ZN(new_n324));
  NAND4_X1  g138(.A1(new_n323), .A2(new_n324), .A3(new_n307), .A4(new_n302), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n319), .A2(new_n325), .ZN(new_n326));
  NAND3_X1  g140(.A1(new_n310), .A2(new_n311), .A3(KEYINPUT16), .ZN(new_n327));
  OR3_X1    g141(.A1(new_n260), .A2(KEYINPUT16), .A3(G140), .ZN(new_n328));
  NAND3_X1  g142(.A1(new_n327), .A2(new_n328), .A3(G146), .ZN(new_n329));
  INV_X1    g143(.A(new_n329), .ZN(new_n330));
  OAI21_X1  g144(.A(G131), .B1(new_n300), .B2(new_n301), .ZN(new_n331));
  INV_X1    g145(.A(G131), .ZN(new_n332));
  NAND3_X1  g146(.A1(new_n304), .A2(new_n332), .A3(new_n305), .ZN(new_n333));
  AOI21_X1  g147(.A(new_n330), .B1(new_n331), .B2(new_n333), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n310), .A2(new_n311), .ZN(new_n335));
  INV_X1    g149(.A(KEYINPUT19), .ZN(new_n336));
  NOR2_X1   g150(.A1(new_n335), .A2(new_n336), .ZN(new_n337));
  AOI21_X1  g151(.A(KEYINPUT19), .B1(new_n310), .B2(new_n311), .ZN(new_n338));
  OAI21_X1  g152(.A(new_n233), .B1(new_n337), .B2(new_n338), .ZN(new_n339));
  NOR2_X1   g153(.A1(new_n339), .A2(KEYINPUT87), .ZN(new_n340));
  INV_X1    g154(.A(KEYINPUT87), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n335), .A2(new_n336), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n315), .A2(KEYINPUT19), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n342), .A2(new_n343), .ZN(new_n344));
  AOI21_X1  g158(.A(new_n341), .B1(new_n344), .B2(new_n233), .ZN(new_n345));
  OAI21_X1  g159(.A(new_n334), .B1(new_n340), .B2(new_n345), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n326), .A2(new_n346), .ZN(new_n347));
  XNOR2_X1  g161(.A(G113), .B(G122), .ZN(new_n348));
  XNOR2_X1  g162(.A(new_n348), .B(new_n199), .ZN(new_n349));
  INV_X1    g163(.A(new_n349), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n347), .A2(new_n350), .ZN(new_n351));
  INV_X1    g165(.A(KEYINPUT88), .ZN(new_n352));
  AOI21_X1  g166(.A(G146), .B1(new_n327), .B2(new_n328), .ZN(new_n353));
  OAI21_X1  g167(.A(new_n352), .B1(new_n330), .B2(new_n353), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n327), .A2(new_n328), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n355), .A2(new_n233), .ZN(new_n356));
  NAND3_X1  g170(.A1(new_n356), .A2(KEYINPUT88), .A3(new_n329), .ZN(new_n357));
  AOI21_X1  g171(.A(KEYINPUT17), .B1(new_n331), .B2(new_n333), .ZN(new_n358));
  AND2_X1   g172(.A1(new_n331), .A2(KEYINPUT17), .ZN(new_n359));
  OAI211_X1 g173(.A(new_n354), .B(new_n357), .C1(new_n358), .C2(new_n359), .ZN(new_n360));
  NAND3_X1  g174(.A1(new_n326), .A2(new_n360), .A3(new_n349), .ZN(new_n361));
  AOI21_X1  g175(.A(new_n298), .B1(new_n351), .B2(new_n361), .ZN(new_n362));
  INV_X1    g176(.A(KEYINPUT20), .ZN(new_n363));
  OAI21_X1  g177(.A(new_n296), .B1(new_n362), .B2(new_n363), .ZN(new_n364));
  AND3_X1   g178(.A1(new_n326), .A2(new_n360), .A3(new_n349), .ZN(new_n365));
  AOI21_X1  g179(.A(new_n349), .B1(new_n326), .B2(new_n346), .ZN(new_n366));
  OAI21_X1  g180(.A(new_n297), .B1(new_n365), .B2(new_n366), .ZN(new_n367));
  NAND3_X1  g181(.A1(new_n367), .A2(KEYINPUT89), .A3(KEYINPUT20), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n339), .A2(KEYINPUT87), .ZN(new_n369));
  NAND3_X1  g183(.A1(new_n344), .A2(new_n341), .A3(new_n233), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n369), .A2(new_n370), .ZN(new_n371));
  AOI22_X1  g185(.A1(new_n371), .A2(new_n334), .B1(new_n319), .B2(new_n325), .ZN(new_n372));
  OAI21_X1  g186(.A(new_n361), .B1(new_n372), .B2(new_n349), .ZN(new_n373));
  AOI21_X1  g187(.A(KEYINPUT20), .B1(new_n298), .B2(KEYINPUT90), .ZN(new_n374));
  OAI211_X1 g188(.A(new_n373), .B(new_n374), .C1(KEYINPUT90), .C2(new_n298), .ZN(new_n375));
  NAND3_X1  g189(.A1(new_n364), .A2(new_n368), .A3(new_n375), .ZN(new_n376));
  INV_X1    g190(.A(G475), .ZN(new_n377));
  AOI21_X1  g191(.A(new_n349), .B1(new_n326), .B2(new_n360), .ZN(new_n378));
  OR2_X1    g192(.A1(new_n365), .A2(new_n378), .ZN(new_n379));
  AOI21_X1  g193(.A(new_n377), .B1(new_n379), .B2(new_n286), .ZN(new_n380));
  INV_X1    g194(.A(new_n380), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n376), .A2(new_n381), .ZN(new_n382));
  INV_X1    g196(.A(G478), .ZN(new_n383));
  INV_X1    g197(.A(KEYINPUT15), .ZN(new_n384));
  AOI21_X1  g198(.A(new_n383), .B1(KEYINPUT94), .B2(new_n384), .ZN(new_n385));
  OAI21_X1  g199(.A(new_n385), .B1(KEYINPUT94), .B2(new_n384), .ZN(new_n386));
  INV_X1    g200(.A(new_n386), .ZN(new_n387));
  XNOR2_X1  g201(.A(KEYINPUT9), .B(G234), .ZN(new_n388));
  INV_X1    g202(.A(G217), .ZN(new_n389));
  NOR3_X1   g203(.A1(new_n388), .A2(new_n389), .A3(G953), .ZN(new_n390));
  INV_X1    g204(.A(new_n390), .ZN(new_n391));
  OAI21_X1  g205(.A(KEYINPUT91), .B1(new_n253), .B2(G143), .ZN(new_n392));
  INV_X1    g206(.A(KEYINPUT91), .ZN(new_n393));
  NAND3_X1  g207(.A1(new_n393), .A2(new_n235), .A3(G128), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n392), .A2(new_n394), .ZN(new_n395));
  INV_X1    g209(.A(KEYINPUT93), .ZN(new_n396));
  OAI21_X1  g210(.A(new_n396), .B1(new_n235), .B2(G128), .ZN(new_n397));
  NAND3_X1  g211(.A1(new_n253), .A2(KEYINPUT93), .A3(G143), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n397), .A2(new_n398), .ZN(new_n399));
  INV_X1    g213(.A(G134), .ZN(new_n400));
  NAND3_X1  g214(.A1(new_n395), .A2(new_n399), .A3(new_n400), .ZN(new_n401));
  INV_X1    g215(.A(G122), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n402), .A2(G116), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n190), .A2(G122), .ZN(new_n404));
  AND2_X1   g218(.A1(new_n403), .A2(new_n404), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n405), .A2(G107), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n403), .A2(new_n404), .ZN(new_n407));
  NAND2_X1  g221(.A1(new_n407), .A2(new_n202), .ZN(new_n408));
  NAND3_X1  g222(.A1(new_n401), .A2(new_n406), .A3(new_n408), .ZN(new_n409));
  XOR2_X1   g223(.A(KEYINPUT92), .B(KEYINPUT13), .Z(new_n410));
  NAND2_X1  g224(.A1(new_n410), .A2(new_n395), .ZN(new_n411));
  XNOR2_X1  g225(.A(KEYINPUT92), .B(KEYINPUT13), .ZN(new_n412));
  NAND3_X1  g226(.A1(new_n412), .A2(new_n394), .A3(new_n392), .ZN(new_n413));
  NAND3_X1  g227(.A1(new_n411), .A2(new_n413), .A3(new_n399), .ZN(new_n414));
  AOI21_X1  g228(.A(new_n409), .B1(G134), .B2(new_n414), .ZN(new_n415));
  AOI21_X1  g229(.A(new_n202), .B1(new_n403), .B2(KEYINPUT14), .ZN(new_n416));
  XNOR2_X1  g230(.A(new_n416), .B(new_n407), .ZN(new_n417));
  NAND2_X1  g231(.A1(new_n395), .A2(new_n399), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n418), .A2(G134), .ZN(new_n419));
  AOI21_X1  g233(.A(new_n417), .B1(new_n401), .B2(new_n419), .ZN(new_n420));
  OAI21_X1  g234(.A(new_n391), .B1(new_n415), .B2(new_n420), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n414), .A2(G134), .ZN(new_n422));
  AND3_X1   g236(.A1(new_n401), .A2(new_n406), .A3(new_n408), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n422), .A2(new_n423), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n419), .A2(new_n401), .ZN(new_n425));
  XNOR2_X1  g239(.A(new_n405), .B(new_n416), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n425), .A2(new_n426), .ZN(new_n427));
  NAND3_X1  g241(.A1(new_n424), .A2(new_n427), .A3(new_n390), .ZN(new_n428));
  AOI21_X1  g242(.A(G902), .B1(new_n421), .B2(new_n428), .ZN(new_n429));
  INV_X1    g243(.A(KEYINPUT95), .ZN(new_n430));
  NOR2_X1   g244(.A1(new_n429), .A2(new_n430), .ZN(new_n431));
  AOI211_X1 g245(.A(KEYINPUT95), .B(G902), .C1(new_n421), .C2(new_n428), .ZN(new_n432));
  OAI21_X1  g246(.A(new_n387), .B1(new_n431), .B2(new_n432), .ZN(new_n433));
  AND3_X1   g247(.A1(new_n424), .A2(new_n427), .A3(new_n390), .ZN(new_n434));
  AOI21_X1  g248(.A(new_n390), .B1(new_n424), .B2(new_n427), .ZN(new_n435));
  OAI21_X1  g249(.A(new_n286), .B1(new_n434), .B2(new_n435), .ZN(new_n436));
  AOI21_X1  g250(.A(new_n387), .B1(new_n436), .B2(KEYINPUT95), .ZN(new_n437));
  INV_X1    g251(.A(new_n437), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n433), .A2(new_n438), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n257), .A2(G952), .ZN(new_n440));
  AOI21_X1  g254(.A(new_n440), .B1(G234), .B2(G237), .ZN(new_n441));
  NAND2_X1  g255(.A1(G234), .A2(G237), .ZN(new_n442));
  NAND3_X1  g256(.A1(new_n442), .A2(G902), .A3(G953), .ZN(new_n443));
  XOR2_X1   g257(.A(new_n443), .B(KEYINPUT96), .Z(new_n444));
  XNOR2_X1  g258(.A(KEYINPUT21), .B(G898), .ZN(new_n445));
  AOI21_X1  g259(.A(new_n441), .B1(new_n444), .B2(new_n445), .ZN(new_n446));
  NOR3_X1   g260(.A1(new_n382), .A2(new_n439), .A3(new_n446), .ZN(new_n447));
  INV_X1    g261(.A(KEYINPUT12), .ZN(new_n448));
  OAI21_X1  g262(.A(KEYINPUT11), .B1(new_n400), .B2(G137), .ZN(new_n449));
  INV_X1    g263(.A(KEYINPUT11), .ZN(new_n450));
  INV_X1    g264(.A(G137), .ZN(new_n451));
  NAND3_X1  g265(.A1(new_n450), .A2(new_n451), .A3(G134), .ZN(new_n452));
  AND2_X1   g266(.A1(new_n449), .A2(new_n452), .ZN(new_n453));
  INV_X1    g267(.A(KEYINPUT65), .ZN(new_n454));
  OAI21_X1  g268(.A(new_n454), .B1(new_n451), .B2(G134), .ZN(new_n455));
  NAND3_X1  g269(.A1(new_n400), .A2(KEYINPUT65), .A3(G137), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n455), .A2(new_n456), .ZN(new_n457));
  OAI21_X1  g271(.A(G131), .B1(new_n453), .B2(new_n457), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n449), .A2(new_n452), .ZN(new_n459));
  NAND4_X1  g273(.A1(new_n459), .A2(new_n332), .A3(new_n455), .A4(new_n456), .ZN(new_n460));
  NAND3_X1  g274(.A1(new_n458), .A2(KEYINPUT66), .A3(new_n460), .ZN(new_n461));
  INV_X1    g275(.A(KEYINPUT66), .ZN(new_n462));
  OAI211_X1 g276(.A(new_n462), .B(G131), .C1(new_n453), .C2(new_n457), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n461), .A2(new_n463), .ZN(new_n464));
  NAND4_X1  g278(.A1(new_n252), .A2(new_n206), .A3(new_n209), .A4(new_n254), .ZN(new_n465));
  INV_X1    g279(.A(new_n465), .ZN(new_n466));
  AOI22_X1  g280(.A1(new_n254), .A2(new_n252), .B1(new_n206), .B2(new_n209), .ZN(new_n467));
  NOR2_X1   g281(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  OAI21_X1  g282(.A(new_n448), .B1(new_n464), .B2(new_n468), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n252), .A2(new_n254), .ZN(new_n470));
  NAND2_X1  g284(.A1(new_n470), .A2(new_n210), .ZN(new_n471));
  NAND2_X1  g285(.A1(new_n471), .A2(new_n465), .ZN(new_n472));
  NAND4_X1  g286(.A1(new_n472), .A2(KEYINPUT12), .A3(new_n463), .A4(new_n461), .ZN(new_n473));
  NAND3_X1  g287(.A1(new_n469), .A2(KEYINPUT81), .A3(new_n473), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n212), .A2(G101), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n475), .A2(KEYINPUT79), .ZN(new_n476));
  NAND3_X1  g290(.A1(new_n212), .A2(new_n213), .A3(G101), .ZN(new_n477));
  NAND4_X1  g291(.A1(new_n476), .A2(KEYINPUT4), .A3(new_n477), .A4(new_n206), .ZN(new_n478));
  AND2_X1   g292(.A1(new_n276), .A2(new_n225), .ZN(new_n479));
  AND2_X1   g293(.A1(new_n252), .A2(new_n254), .ZN(new_n480));
  AND2_X1   g294(.A1(new_n206), .A2(new_n209), .ZN(new_n481));
  INV_X1    g295(.A(KEYINPUT10), .ZN(new_n482));
  NAND3_X1  g296(.A1(new_n480), .A2(new_n481), .A3(new_n482), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n465), .A2(KEYINPUT10), .ZN(new_n484));
  AOI22_X1  g298(.A1(new_n478), .A2(new_n479), .B1(new_n483), .B2(new_n484), .ZN(new_n485));
  INV_X1    g299(.A(KEYINPUT80), .ZN(new_n486));
  AOI21_X1  g300(.A(new_n486), .B1(new_n461), .B2(new_n463), .ZN(new_n487));
  AND3_X1   g301(.A1(new_n461), .A2(new_n486), .A3(new_n463), .ZN(new_n488));
  OAI21_X1  g302(.A(new_n485), .B1(new_n487), .B2(new_n488), .ZN(new_n489));
  XNOR2_X1  g303(.A(G110), .B(G140), .ZN(new_n490));
  INV_X1    g304(.A(G227), .ZN(new_n491));
  NOR2_X1   g305(.A1(new_n491), .A2(G953), .ZN(new_n492));
  XNOR2_X1  g306(.A(new_n490), .B(new_n492), .ZN(new_n493));
  INV_X1    g307(.A(new_n493), .ZN(new_n494));
  NAND3_X1  g308(.A1(new_n474), .A2(new_n489), .A3(new_n494), .ZN(new_n495));
  AOI21_X1  g309(.A(KEYINPUT81), .B1(new_n469), .B2(new_n473), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n478), .A2(new_n479), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n483), .A2(new_n484), .ZN(new_n498));
  AOI21_X1  g312(.A(new_n464), .B1(new_n497), .B2(new_n498), .ZN(new_n499));
  NAND2_X1  g313(.A1(new_n460), .A2(KEYINPUT66), .ZN(new_n500));
  INV_X1    g314(.A(new_n457), .ZN(new_n501));
  AOI21_X1  g315(.A(new_n332), .B1(new_n501), .B2(new_n459), .ZN(new_n502));
  NOR2_X1   g316(.A1(new_n500), .A2(new_n502), .ZN(new_n503));
  INV_X1    g317(.A(new_n463), .ZN(new_n504));
  OAI21_X1  g318(.A(KEYINPUT80), .B1(new_n503), .B2(new_n504), .ZN(new_n505));
  NAND3_X1  g319(.A1(new_n461), .A2(new_n486), .A3(new_n463), .ZN(new_n506));
  NAND2_X1  g320(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  AOI21_X1  g321(.A(new_n499), .B1(new_n485), .B2(new_n507), .ZN(new_n508));
  OAI22_X1  g322(.A1(new_n495), .A2(new_n496), .B1(new_n508), .B2(new_n494), .ZN(new_n509));
  INV_X1    g323(.A(G469), .ZN(new_n510));
  NAND3_X1  g324(.A1(new_n509), .A2(new_n510), .A3(new_n286), .ZN(new_n511));
  NAND2_X1  g325(.A1(G469), .A2(G902), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n497), .A2(new_n498), .ZN(new_n513));
  AND2_X1   g327(.A1(new_n461), .A2(new_n463), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  AND3_X1   g329(.A1(new_n489), .A2(new_n515), .A3(new_n494), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n469), .A2(new_n473), .ZN(new_n517));
  AOI21_X1  g331(.A(new_n494), .B1(new_n517), .B2(new_n489), .ZN(new_n518));
  NOR2_X1   g332(.A1(new_n516), .A2(new_n518), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n519), .A2(G469), .ZN(new_n520));
  NAND3_X1  g334(.A1(new_n511), .A2(new_n512), .A3(new_n520), .ZN(new_n521));
  OAI21_X1  g335(.A(G221), .B1(new_n388), .B2(G902), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  INV_X1    g337(.A(new_n523), .ZN(new_n524));
  AND3_X1   g338(.A1(new_n295), .A2(new_n447), .A3(new_n524), .ZN(new_n525));
  INV_X1    g339(.A(KEYINPUT78), .ZN(new_n526));
  XNOR2_X1  g340(.A(KEYINPUT22), .B(G137), .ZN(new_n527));
  AND3_X1   g341(.A1(new_n257), .A2(G221), .A3(G234), .ZN(new_n528));
  XNOR2_X1  g342(.A(new_n527), .B(new_n528), .ZN(new_n529));
  OAI21_X1  g343(.A(KEYINPUT23), .B1(new_n253), .B2(G119), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n530), .A2(KEYINPUT71), .ZN(new_n531));
  NAND2_X1  g345(.A1(new_n188), .A2(G128), .ZN(new_n532));
  INV_X1    g346(.A(KEYINPUT71), .ZN(new_n533));
  NAND3_X1  g347(.A1(new_n532), .A2(new_n533), .A3(KEYINPUT23), .ZN(new_n534));
  NAND2_X1  g348(.A1(new_n253), .A2(G119), .ZN(new_n535));
  INV_X1    g349(.A(KEYINPUT72), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  NAND3_X1  g351(.A1(new_n253), .A2(KEYINPUT72), .A3(G119), .ZN(new_n538));
  NAND4_X1  g352(.A1(new_n531), .A2(new_n534), .A3(new_n537), .A4(new_n538), .ZN(new_n539));
  NAND3_X1  g353(.A1(new_n253), .A2(KEYINPUT23), .A3(G119), .ZN(new_n540));
  XNOR2_X1  g354(.A(KEYINPUT73), .B(G110), .ZN(new_n541));
  NAND3_X1  g355(.A1(new_n539), .A2(new_n540), .A3(new_n541), .ZN(new_n542));
  NAND2_X1  g356(.A1(new_n535), .A2(new_n532), .ZN(new_n543));
  XNOR2_X1  g357(.A(KEYINPUT24), .B(G110), .ZN(new_n544));
  AND3_X1   g358(.A1(new_n543), .A2(new_n544), .A3(KEYINPUT74), .ZN(new_n545));
  AOI21_X1  g359(.A(KEYINPUT74), .B1(new_n543), .B2(new_n544), .ZN(new_n546));
  NOR2_X1   g360(.A1(new_n545), .A2(new_n546), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n542), .A2(new_n547), .ZN(new_n548));
  OAI21_X1  g362(.A(new_n329), .B1(new_n321), .B2(new_n322), .ZN(new_n549));
  INV_X1    g363(.A(new_n549), .ZN(new_n550));
  NAND2_X1  g364(.A1(new_n548), .A2(new_n550), .ZN(new_n551));
  INV_X1    g365(.A(G110), .ZN(new_n552));
  AOI21_X1  g366(.A(new_n552), .B1(new_n539), .B2(new_n540), .ZN(new_n553));
  INV_X1    g367(.A(new_n553), .ZN(new_n554));
  NOR2_X1   g368(.A1(new_n543), .A2(new_n544), .ZN(new_n555));
  AOI21_X1  g369(.A(new_n555), .B1(new_n356), .B2(new_n329), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n554), .A2(new_n556), .ZN(new_n557));
  AOI21_X1  g371(.A(new_n529), .B1(new_n551), .B2(new_n557), .ZN(new_n558));
  INV_X1    g372(.A(KEYINPUT76), .ZN(new_n559));
  OAI22_X1  g373(.A1(new_n330), .A2(new_n353), .B1(new_n543), .B2(new_n544), .ZN(new_n560));
  NOR2_X1   g374(.A1(new_n560), .A2(new_n553), .ZN(new_n561));
  AOI21_X1  g375(.A(new_n549), .B1(new_n542), .B2(new_n547), .ZN(new_n562));
  OAI21_X1  g376(.A(new_n559), .B1(new_n561), .B2(new_n562), .ZN(new_n563));
  NAND3_X1  g377(.A1(new_n551), .A2(new_n557), .A3(KEYINPUT76), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n563), .A2(new_n564), .ZN(new_n565));
  AOI21_X1  g379(.A(new_n558), .B1(new_n565), .B2(new_n529), .ZN(new_n566));
  AOI21_X1  g380(.A(new_n389), .B1(G234), .B2(new_n286), .ZN(new_n567));
  NOR2_X1   g381(.A1(new_n567), .A2(G902), .ZN(new_n568));
  XNOR2_X1  g382(.A(new_n568), .B(KEYINPUT77), .ZN(new_n569));
  INV_X1    g383(.A(new_n569), .ZN(new_n570));
  NOR2_X1   g384(.A1(new_n566), .A2(new_n570), .ZN(new_n571));
  INV_X1    g385(.A(KEYINPUT25), .ZN(new_n572));
  OAI21_X1  g386(.A(new_n572), .B1(new_n566), .B2(G902), .ZN(new_n573));
  INV_X1    g387(.A(new_n529), .ZN(new_n574));
  AOI21_X1  g388(.A(new_n574), .B1(new_n563), .B2(new_n564), .ZN(new_n575));
  OAI211_X1 g389(.A(KEYINPUT25), .B(new_n286), .C1(new_n575), .C2(new_n558), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n573), .A2(new_n576), .ZN(new_n577));
  AOI21_X1  g391(.A(new_n571), .B1(new_n577), .B2(new_n567), .ZN(new_n578));
  INV_X1    g392(.A(new_n578), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n299), .A2(G210), .ZN(new_n580));
  XNOR2_X1  g394(.A(new_n580), .B(KEYINPUT27), .ZN(new_n581));
  XNOR2_X1  g395(.A(KEYINPUT26), .B(G101), .ZN(new_n582));
  XNOR2_X1  g396(.A(new_n581), .B(new_n582), .ZN(new_n583));
  INV_X1    g397(.A(new_n583), .ZN(new_n584));
  XNOR2_X1  g398(.A(KEYINPUT68), .B(KEYINPUT28), .ZN(new_n585));
  INV_X1    g399(.A(new_n585), .ZN(new_n586));
  NAND3_X1  g400(.A1(new_n461), .A2(new_n276), .A3(new_n463), .ZN(new_n587));
  NOR2_X1   g401(.A1(new_n400), .A2(G137), .ZN(new_n588));
  NOR2_X1   g402(.A1(new_n451), .A2(G134), .ZN(new_n589));
  OAI21_X1  g403(.A(G131), .B1(new_n588), .B2(new_n589), .ZN(new_n590));
  NAND3_X1  g404(.A1(new_n480), .A2(new_n460), .A3(new_n590), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n587), .A2(new_n591), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n221), .A2(new_n223), .ZN(new_n593));
  INV_X1    g407(.A(new_n593), .ZN(new_n594));
  NAND2_X1  g408(.A1(new_n592), .A2(new_n594), .ZN(new_n595));
  NAND3_X1  g409(.A1(new_n587), .A2(new_n593), .A3(new_n591), .ZN(new_n596));
  AOI21_X1  g410(.A(new_n586), .B1(new_n595), .B2(new_n596), .ZN(new_n597));
  INV_X1    g411(.A(KEYINPUT28), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n596), .A2(new_n598), .ZN(new_n599));
  INV_X1    g413(.A(new_n599), .ZN(new_n600));
  OAI21_X1  g414(.A(new_n584), .B1(new_n597), .B2(new_n600), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n592), .A2(KEYINPUT30), .ZN(new_n602));
  INV_X1    g416(.A(KEYINPUT30), .ZN(new_n603));
  NAND3_X1  g417(.A1(new_n587), .A2(new_n603), .A3(new_n591), .ZN(new_n604));
  AOI21_X1  g418(.A(new_n593), .B1(new_n602), .B2(new_n604), .ZN(new_n605));
  NAND2_X1  g419(.A1(new_n596), .A2(new_n583), .ZN(new_n606));
  OAI21_X1  g420(.A(KEYINPUT31), .B1(new_n605), .B2(new_n606), .ZN(new_n607));
  AND3_X1   g421(.A1(new_n587), .A2(new_n603), .A3(new_n591), .ZN(new_n608));
  AOI21_X1  g422(.A(new_n603), .B1(new_n587), .B2(new_n591), .ZN(new_n609));
  OAI21_X1  g423(.A(new_n594), .B1(new_n608), .B2(new_n609), .ZN(new_n610));
  INV_X1    g424(.A(KEYINPUT31), .ZN(new_n611));
  INV_X1    g425(.A(new_n606), .ZN(new_n612));
  NAND3_X1  g426(.A1(new_n610), .A2(new_n611), .A3(new_n612), .ZN(new_n613));
  NAND3_X1  g427(.A1(new_n601), .A2(new_n607), .A3(new_n613), .ZN(new_n614));
  NOR2_X1   g428(.A1(G472), .A2(G902), .ZN(new_n615));
  XNOR2_X1  g429(.A(new_n615), .B(KEYINPUT69), .ZN(new_n616));
  AND3_X1   g430(.A1(new_n614), .A2(KEYINPUT32), .A3(new_n616), .ZN(new_n617));
  AOI21_X1  g431(.A(KEYINPUT32), .B1(new_n614), .B2(new_n616), .ZN(new_n618));
  NOR2_X1   g432(.A1(new_n617), .A2(new_n618), .ZN(new_n619));
  INV_X1    g433(.A(KEYINPUT29), .ZN(new_n620));
  AND3_X1   g434(.A1(new_n587), .A2(new_n593), .A3(new_n591), .ZN(new_n621));
  NOR3_X1   g435(.A1(new_n605), .A2(new_n583), .A3(new_n621), .ZN(new_n622));
  AOI21_X1  g436(.A(new_n593), .B1(new_n587), .B2(new_n591), .ZN(new_n623));
  OAI21_X1  g437(.A(new_n585), .B1(new_n621), .B2(new_n623), .ZN(new_n624));
  AOI21_X1  g438(.A(new_n584), .B1(new_n624), .B2(new_n599), .ZN(new_n625));
  OAI21_X1  g439(.A(new_n620), .B1(new_n622), .B2(new_n625), .ZN(new_n626));
  NAND2_X1  g440(.A1(new_n595), .A2(new_n596), .ZN(new_n627));
  NAND2_X1  g441(.A1(new_n627), .A2(KEYINPUT28), .ZN(new_n628));
  NAND2_X1  g442(.A1(new_n628), .A2(KEYINPUT70), .ZN(new_n629));
  AOI21_X1  g443(.A(new_n598), .B1(new_n595), .B2(new_n596), .ZN(new_n630));
  INV_X1    g444(.A(KEYINPUT70), .ZN(new_n631));
  AOI21_X1  g445(.A(new_n600), .B1(new_n630), .B2(new_n631), .ZN(new_n632));
  NOR2_X1   g446(.A1(new_n584), .A2(new_n620), .ZN(new_n633));
  NAND3_X1  g447(.A1(new_n629), .A2(new_n632), .A3(new_n633), .ZN(new_n634));
  NAND3_X1  g448(.A1(new_n626), .A2(new_n286), .A3(new_n634), .ZN(new_n635));
  NAND2_X1  g449(.A1(new_n635), .A2(G472), .ZN(new_n636));
  AOI211_X1 g450(.A(new_n526), .B(new_n579), .C1(new_n619), .C2(new_n636), .ZN(new_n637));
  INV_X1    g451(.A(new_n618), .ZN(new_n638));
  NAND3_X1  g452(.A1(new_n614), .A2(KEYINPUT32), .A3(new_n616), .ZN(new_n639));
  NAND3_X1  g453(.A1(new_n636), .A2(new_n638), .A3(new_n639), .ZN(new_n640));
  AOI21_X1  g454(.A(KEYINPUT78), .B1(new_n640), .B2(new_n578), .ZN(new_n641));
  OAI21_X1  g455(.A(new_n525), .B1(new_n637), .B2(new_n641), .ZN(new_n642));
  XNOR2_X1  g456(.A(new_n642), .B(G101), .ZN(G3));
  NAND2_X1  g457(.A1(new_n614), .A2(new_n286), .ZN(new_n644));
  NAND2_X1  g458(.A1(new_n644), .A2(G472), .ZN(new_n645));
  NAND2_X1  g459(.A1(new_n614), .A2(new_n616), .ZN(new_n646));
  NAND2_X1  g460(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  NOR3_X1   g461(.A1(new_n647), .A2(new_n523), .A3(new_n579), .ZN(new_n648));
  NAND2_X1  g462(.A1(new_n421), .A2(new_n428), .ZN(new_n649));
  OR2_X1    g463(.A1(new_n649), .A2(KEYINPUT33), .ZN(new_n650));
  NAND2_X1  g464(.A1(new_n649), .A2(KEYINPUT33), .ZN(new_n651));
  NAND3_X1  g465(.A1(new_n650), .A2(G478), .A3(new_n651), .ZN(new_n652));
  NOR2_X1   g466(.A1(new_n383), .A2(new_n286), .ZN(new_n653));
  AOI21_X1  g467(.A(new_n653), .B1(new_n429), .B2(new_n383), .ZN(new_n654));
  NAND2_X1  g468(.A1(new_n652), .A2(new_n654), .ZN(new_n655));
  AOI21_X1  g469(.A(new_n655), .B1(new_n376), .B2(new_n381), .ZN(new_n656));
  INV_X1    g470(.A(new_n656), .ZN(new_n657));
  NOR3_X1   g471(.A1(new_n657), .A2(new_n291), .A3(new_n446), .ZN(new_n658));
  NAND2_X1  g472(.A1(new_n648), .A2(new_n658), .ZN(new_n659));
  XOR2_X1   g473(.A(KEYINPUT34), .B(G104), .Z(new_n660));
  XNOR2_X1  g474(.A(new_n659), .B(new_n660), .ZN(G6));
  INV_X1    g475(.A(new_n187), .ZN(new_n662));
  NAND2_X1  g476(.A1(new_n268), .A2(new_n287), .ZN(new_n663));
  INV_X1    g477(.A(new_n288), .ZN(new_n664));
  NAND2_X1  g478(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  NAND3_X1  g479(.A1(new_n268), .A2(new_n287), .A3(new_n288), .ZN(new_n666));
  AOI21_X1  g480(.A(new_n662), .B1(new_n665), .B2(new_n666), .ZN(new_n667));
  AOI211_X1 g481(.A(new_n296), .B(new_n363), .C1(new_n373), .C2(new_n297), .ZN(new_n668));
  AOI21_X1  g482(.A(KEYINPUT89), .B1(new_n367), .B2(KEYINPUT20), .ZN(new_n669));
  NOR2_X1   g483(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  NAND2_X1  g484(.A1(new_n362), .A2(new_n363), .ZN(new_n671));
  AOI21_X1  g485(.A(new_n380), .B1(new_n670), .B2(new_n671), .ZN(new_n672));
  INV_X1    g486(.A(new_n446), .ZN(new_n673));
  AND4_X1   g487(.A1(new_n667), .A2(new_n672), .A3(new_n439), .A4(new_n673), .ZN(new_n674));
  NAND2_X1  g488(.A1(new_n648), .A2(new_n674), .ZN(new_n675));
  XOR2_X1   g489(.A(KEYINPUT35), .B(G107), .Z(new_n676));
  XNOR2_X1  g490(.A(new_n675), .B(new_n676), .ZN(G9));
  NOR2_X1   g491(.A1(new_n529), .A2(KEYINPUT36), .ZN(new_n678));
  AND2_X1   g492(.A1(new_n565), .A2(new_n678), .ZN(new_n679));
  NOR2_X1   g493(.A1(new_n565), .A2(new_n678), .ZN(new_n680));
  NOR3_X1   g494(.A1(new_n679), .A2(new_n680), .A3(new_n570), .ZN(new_n681));
  AOI21_X1  g495(.A(new_n681), .B1(new_n577), .B2(new_n567), .ZN(new_n682));
  NOR3_X1   g496(.A1(new_n647), .A2(new_n523), .A3(new_n682), .ZN(new_n683));
  AOI21_X1  g497(.A(new_n380), .B1(new_n670), .B2(new_n375), .ZN(new_n684));
  NOR2_X1   g498(.A1(new_n439), .A2(new_n446), .ZN(new_n685));
  AND4_X1   g499(.A1(new_n292), .A2(new_n294), .A3(new_n684), .A4(new_n685), .ZN(new_n686));
  NAND2_X1  g500(.A1(new_n683), .A2(new_n686), .ZN(new_n687));
  XOR2_X1   g501(.A(KEYINPUT37), .B(G110), .Z(new_n688));
  XNOR2_X1  g502(.A(new_n687), .B(new_n688), .ZN(G12));
  NOR2_X1   g503(.A1(new_n523), .A2(new_n682), .ZN(new_n690));
  NAND3_X1  g504(.A1(new_n364), .A2(new_n368), .A3(new_n671), .ZN(new_n691));
  INV_X1    g505(.A(G900), .ZN(new_n692));
  AOI21_X1  g506(.A(new_n441), .B1(new_n444), .B2(new_n692), .ZN(new_n693));
  INV_X1    g507(.A(new_n693), .ZN(new_n694));
  NAND4_X1  g508(.A1(new_n691), .A2(new_n439), .A3(new_n381), .A4(new_n694), .ZN(new_n695));
  INV_X1    g509(.A(new_n695), .ZN(new_n696));
  NAND4_X1  g510(.A1(new_n690), .A2(new_n640), .A3(new_n667), .A4(new_n696), .ZN(new_n697));
  XNOR2_X1  g511(.A(new_n697), .B(G128), .ZN(G30));
  XOR2_X1   g512(.A(new_n693), .B(KEYINPUT39), .Z(new_n699));
  NAND2_X1  g513(.A1(new_n524), .A2(new_n699), .ZN(new_n700));
  XNOR2_X1  g514(.A(new_n700), .B(KEYINPUT40), .ZN(new_n701));
  AOI21_X1  g515(.A(new_n584), .B1(new_n610), .B2(new_n596), .ZN(new_n702));
  OAI21_X1  g516(.A(new_n286), .B1(new_n627), .B2(new_n583), .ZN(new_n703));
  OAI21_X1  g517(.A(G472), .B1(new_n702), .B2(new_n703), .ZN(new_n704));
  NAND3_X1  g518(.A1(new_n638), .A2(new_n639), .A3(new_n704), .ZN(new_n705));
  INV_X1    g519(.A(new_n705), .ZN(new_n706));
  NAND2_X1  g520(.A1(new_n665), .A2(new_n666), .ZN(new_n707));
  XOR2_X1   g521(.A(KEYINPUT97), .B(KEYINPUT38), .Z(new_n708));
  XNOR2_X1  g522(.A(new_n707), .B(new_n708), .ZN(new_n709));
  NAND2_X1  g523(.A1(new_n436), .A2(KEYINPUT95), .ZN(new_n710));
  NAND2_X1  g524(.A1(new_n429), .A2(new_n430), .ZN(new_n711));
  NAND2_X1  g525(.A1(new_n710), .A2(new_n711), .ZN(new_n712));
  AOI21_X1  g526(.A(new_n437), .B1(new_n712), .B2(new_n387), .ZN(new_n713));
  AOI21_X1  g527(.A(new_n713), .B1(new_n376), .B2(new_n381), .ZN(new_n714));
  NAND3_X1  g528(.A1(new_n714), .A2(new_n187), .A3(new_n682), .ZN(new_n715));
  OR4_X1    g529(.A1(new_n701), .A2(new_n706), .A3(new_n709), .A4(new_n715), .ZN(new_n716));
  XNOR2_X1  g530(.A(new_n716), .B(G143), .ZN(G45));
  INV_X1    g531(.A(new_n655), .ZN(new_n718));
  NAND4_X1  g532(.A1(new_n382), .A2(new_n667), .A3(new_n718), .A4(new_n694), .ZN(new_n719));
  INV_X1    g533(.A(KEYINPUT98), .ZN(new_n720));
  NAND2_X1  g534(.A1(new_n719), .A2(new_n720), .ZN(new_n721));
  NAND4_X1  g535(.A1(new_n656), .A2(KEYINPUT98), .A3(new_n667), .A4(new_n694), .ZN(new_n722));
  NAND4_X1  g536(.A1(new_n721), .A2(new_n690), .A3(new_n640), .A4(new_n722), .ZN(new_n723));
  XNOR2_X1  g537(.A(new_n723), .B(G146), .ZN(G48));
  AOI21_X1  g538(.A(new_n579), .B1(new_n619), .B2(new_n636), .ZN(new_n725));
  NAND2_X1  g539(.A1(new_n511), .A2(new_n522), .ZN(new_n726));
  INV_X1    g540(.A(KEYINPUT99), .ZN(new_n727));
  INV_X1    g541(.A(KEYINPUT81), .ZN(new_n728));
  AOI21_X1  g542(.A(KEYINPUT12), .B1(new_n514), .B2(new_n472), .ZN(new_n729));
  INV_X1    g543(.A(new_n473), .ZN(new_n730));
  OAI21_X1  g544(.A(new_n728), .B1(new_n729), .B2(new_n730), .ZN(new_n731));
  AOI21_X1  g545(.A(new_n493), .B1(new_n507), .B2(new_n485), .ZN(new_n732));
  NAND3_X1  g546(.A1(new_n731), .A2(new_n732), .A3(new_n474), .ZN(new_n733));
  NAND2_X1  g547(.A1(new_n489), .A2(new_n515), .ZN(new_n734));
  NAND2_X1  g548(.A1(new_n734), .A2(new_n493), .ZN(new_n735));
  AOI21_X1  g549(.A(G902), .B1(new_n733), .B2(new_n735), .ZN(new_n736));
  OAI21_X1  g550(.A(new_n727), .B1(new_n736), .B2(new_n510), .ZN(new_n737));
  NAND2_X1  g551(.A1(new_n509), .A2(new_n286), .ZN(new_n738));
  NAND3_X1  g552(.A1(new_n738), .A2(KEYINPUT99), .A3(G469), .ZN(new_n739));
  AOI21_X1  g553(.A(new_n726), .B1(new_n737), .B2(new_n739), .ZN(new_n740));
  NAND3_X1  g554(.A1(new_n725), .A2(new_n658), .A3(new_n740), .ZN(new_n741));
  XNOR2_X1  g555(.A(KEYINPUT41), .B(G113), .ZN(new_n742));
  XNOR2_X1  g556(.A(new_n741), .B(new_n742), .ZN(G15));
  NAND3_X1  g557(.A1(new_n725), .A2(new_n674), .A3(new_n740), .ZN(new_n744));
  XOR2_X1   g558(.A(KEYINPUT100), .B(G116), .Z(new_n745));
  XNOR2_X1  g559(.A(new_n744), .B(new_n745), .ZN(G18));
  INV_X1    g560(.A(new_n522), .ZN(new_n747));
  AOI21_X1  g561(.A(new_n747), .B1(new_n736), .B2(new_n510), .ZN(new_n748));
  AOI21_X1  g562(.A(KEYINPUT99), .B1(new_n738), .B2(G469), .ZN(new_n749));
  NOR3_X1   g563(.A1(new_n736), .A2(new_n727), .A3(new_n510), .ZN(new_n750));
  OAI211_X1 g564(.A(new_n667), .B(new_n748), .C1(new_n749), .C2(new_n750), .ZN(new_n751));
  INV_X1    g565(.A(new_n751), .ZN(new_n752));
  NOR3_X1   g566(.A1(new_n561), .A2(new_n562), .A3(new_n559), .ZN(new_n753));
  AOI21_X1  g567(.A(KEYINPUT76), .B1(new_n551), .B2(new_n557), .ZN(new_n754));
  OAI21_X1  g568(.A(new_n529), .B1(new_n753), .B2(new_n754), .ZN(new_n755));
  INV_X1    g569(.A(new_n558), .ZN(new_n756));
  NAND2_X1  g570(.A1(new_n755), .A2(new_n756), .ZN(new_n757));
  AOI21_X1  g571(.A(KEYINPUT25), .B1(new_n757), .B2(new_n286), .ZN(new_n758));
  INV_X1    g572(.A(new_n576), .ZN(new_n759));
  OAI21_X1  g573(.A(new_n567), .B1(new_n758), .B2(new_n759), .ZN(new_n760));
  INV_X1    g574(.A(new_n681), .ZN(new_n761));
  NAND2_X1  g575(.A1(new_n760), .A2(new_n761), .ZN(new_n762));
  NAND4_X1  g576(.A1(new_n752), .A2(new_n640), .A3(new_n447), .A4(new_n762), .ZN(new_n763));
  XNOR2_X1  g577(.A(new_n763), .B(G119), .ZN(G21));
  NAND3_X1  g578(.A1(new_n382), .A2(new_n667), .A3(new_n439), .ZN(new_n765));
  INV_X1    g579(.A(KEYINPUT102), .ZN(new_n766));
  NAND2_X1  g580(.A1(new_n765), .A2(new_n766), .ZN(new_n767));
  NAND3_X1  g581(.A1(new_n714), .A2(KEYINPUT102), .A3(new_n667), .ZN(new_n768));
  NAND2_X1  g582(.A1(new_n767), .A2(new_n768), .ZN(new_n769));
  OAI211_X1 g583(.A(new_n673), .B(new_n748), .C1(new_n749), .C2(new_n750), .ZN(new_n770));
  XOR2_X1   g584(.A(new_n616), .B(KEYINPUT101), .Z(new_n771));
  AOI21_X1  g585(.A(new_n583), .B1(new_n629), .B2(new_n632), .ZN(new_n772));
  NAND2_X1  g586(.A1(new_n607), .A2(new_n613), .ZN(new_n773));
  OAI21_X1  g587(.A(new_n771), .B1(new_n772), .B2(new_n773), .ZN(new_n774));
  NAND3_X1  g588(.A1(new_n645), .A2(new_n578), .A3(new_n774), .ZN(new_n775));
  NOR2_X1   g589(.A1(new_n770), .A2(new_n775), .ZN(new_n776));
  NAND2_X1  g590(.A1(new_n769), .A2(new_n776), .ZN(new_n777));
  XOR2_X1   g591(.A(KEYINPUT103), .B(G122), .Z(new_n778));
  XNOR2_X1  g592(.A(new_n777), .B(new_n778), .ZN(G24));
  INV_X1    g593(.A(KEYINPUT105), .ZN(new_n780));
  NAND3_X1  g594(.A1(new_n382), .A2(new_n718), .A3(new_n694), .ZN(new_n781));
  INV_X1    g595(.A(KEYINPUT104), .ZN(new_n782));
  NAND2_X1  g596(.A1(new_n781), .A2(new_n782), .ZN(new_n783));
  NAND3_X1  g597(.A1(new_n656), .A2(KEYINPUT104), .A3(new_n694), .ZN(new_n784));
  NAND2_X1  g598(.A1(new_n783), .A2(new_n784), .ZN(new_n785));
  INV_X1    g599(.A(G472), .ZN(new_n786));
  AOI21_X1  g600(.A(new_n786), .B1(new_n614), .B2(new_n286), .ZN(new_n787));
  INV_X1    g601(.A(new_n771), .ZN(new_n788));
  NOR3_X1   g602(.A1(new_n605), .A2(KEYINPUT31), .A3(new_n606), .ZN(new_n789));
  AOI21_X1  g603(.A(new_n611), .B1(new_n610), .B2(new_n612), .ZN(new_n790));
  NOR2_X1   g604(.A1(new_n789), .A2(new_n790), .ZN(new_n791));
  OAI211_X1 g605(.A(new_n631), .B(KEYINPUT28), .C1(new_n621), .C2(new_n623), .ZN(new_n792));
  NAND2_X1  g606(.A1(new_n792), .A2(new_n599), .ZN(new_n793));
  AOI21_X1  g607(.A(new_n631), .B1(new_n627), .B2(KEYINPUT28), .ZN(new_n794));
  OAI21_X1  g608(.A(new_n584), .B1(new_n793), .B2(new_n794), .ZN(new_n795));
  AOI21_X1  g609(.A(new_n788), .B1(new_n791), .B2(new_n795), .ZN(new_n796));
  NOR2_X1   g610(.A1(new_n787), .A2(new_n796), .ZN(new_n797));
  NAND4_X1  g611(.A1(new_n740), .A2(new_n797), .A3(new_n667), .A4(new_n762), .ZN(new_n798));
  OAI21_X1  g612(.A(new_n780), .B1(new_n785), .B2(new_n798), .ZN(new_n799));
  AND4_X1   g613(.A1(KEYINPUT104), .A2(new_n382), .A3(new_n718), .A4(new_n694), .ZN(new_n800));
  AOI21_X1  g614(.A(KEYINPUT104), .B1(new_n656), .B2(new_n694), .ZN(new_n801));
  NOR2_X1   g615(.A1(new_n800), .A2(new_n801), .ZN(new_n802));
  NAND3_X1  g616(.A1(new_n762), .A2(new_n645), .A3(new_n774), .ZN(new_n803));
  NOR2_X1   g617(.A1(new_n803), .A2(new_n751), .ZN(new_n804));
  NAND3_X1  g618(.A1(new_n802), .A2(new_n804), .A3(KEYINPUT105), .ZN(new_n805));
  NAND2_X1  g619(.A1(new_n799), .A2(new_n805), .ZN(new_n806));
  XNOR2_X1  g620(.A(new_n806), .B(G125), .ZN(G27));
  OAI21_X1  g621(.A(KEYINPUT106), .B1(new_n516), .B2(new_n518), .ZN(new_n808));
  INV_X1    g622(.A(KEYINPUT106), .ZN(new_n809));
  AND2_X1   g623(.A1(new_n517), .A2(new_n489), .ZN(new_n810));
  OAI21_X1  g624(.A(new_n809), .B1(new_n810), .B2(new_n494), .ZN(new_n811));
  NAND3_X1  g625(.A1(new_n808), .A2(G469), .A3(new_n811), .ZN(new_n812));
  NAND3_X1  g626(.A1(new_n812), .A2(new_n511), .A3(new_n512), .ZN(new_n813));
  NOR3_X1   g627(.A1(new_n289), .A2(new_n290), .A3(new_n662), .ZN(new_n814));
  AND3_X1   g628(.A1(new_n813), .A2(new_n522), .A3(new_n814), .ZN(new_n815));
  AND3_X1   g629(.A1(new_n640), .A2(new_n815), .A3(new_n578), .ZN(new_n816));
  AOI21_X1  g630(.A(KEYINPUT42), .B1(new_n816), .B2(new_n802), .ZN(new_n817));
  INV_X1    g631(.A(new_n636), .ZN(new_n818));
  OAI21_X1  g632(.A(KEYINPUT107), .B1(new_n617), .B2(new_n618), .ZN(new_n819));
  OR2_X1    g633(.A1(new_n618), .A2(KEYINPUT107), .ZN(new_n820));
  NAND2_X1  g634(.A1(new_n819), .A2(new_n820), .ZN(new_n821));
  AOI21_X1  g635(.A(new_n818), .B1(new_n821), .B2(KEYINPUT108), .ZN(new_n822));
  INV_X1    g636(.A(KEYINPUT108), .ZN(new_n823));
  NAND3_X1  g637(.A1(new_n819), .A2(new_n820), .A3(new_n823), .ZN(new_n824));
  AOI21_X1  g638(.A(new_n579), .B1(new_n822), .B2(new_n824), .ZN(new_n825));
  AND3_X1   g639(.A1(new_n802), .A2(KEYINPUT42), .A3(new_n815), .ZN(new_n826));
  AOI21_X1  g640(.A(new_n817), .B1(new_n825), .B2(new_n826), .ZN(new_n827));
  XNOR2_X1  g641(.A(new_n827), .B(new_n332), .ZN(G33));
  NAND3_X1  g642(.A1(new_n725), .A2(new_n696), .A3(new_n815), .ZN(new_n829));
  XNOR2_X1  g643(.A(new_n829), .B(G134), .ZN(G36));
  NAND3_X1  g644(.A1(new_n808), .A2(KEYINPUT45), .A3(new_n811), .ZN(new_n831));
  OAI211_X1 g645(.A(new_n831), .B(G469), .C1(KEYINPUT45), .C2(new_n519), .ZN(new_n832));
  NAND2_X1  g646(.A1(new_n832), .A2(new_n512), .ZN(new_n833));
  INV_X1    g647(.A(KEYINPUT46), .ZN(new_n834));
  NAND2_X1  g648(.A1(new_n833), .A2(new_n834), .ZN(new_n835));
  NAND2_X1  g649(.A1(new_n835), .A2(new_n511), .ZN(new_n836));
  NOR2_X1   g650(.A1(new_n833), .A2(new_n834), .ZN(new_n837));
  OR2_X1    g651(.A1(new_n836), .A2(new_n837), .ZN(new_n838));
  NAND3_X1  g652(.A1(new_n838), .A2(new_n522), .A3(new_n699), .ZN(new_n839));
  INV_X1    g653(.A(new_n839), .ZN(new_n840));
  NAND2_X1  g654(.A1(new_n684), .A2(new_n718), .ZN(new_n841));
  OR2_X1    g655(.A1(new_n841), .A2(KEYINPUT43), .ZN(new_n842));
  NAND2_X1  g656(.A1(new_n841), .A2(KEYINPUT43), .ZN(new_n843));
  NAND4_X1  g657(.A1(new_n842), .A2(new_n647), .A3(new_n762), .A4(new_n843), .ZN(new_n844));
  INV_X1    g658(.A(KEYINPUT44), .ZN(new_n845));
  OR2_X1    g659(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  INV_X1    g660(.A(new_n814), .ZN(new_n847));
  AOI21_X1  g661(.A(new_n847), .B1(new_n844), .B2(new_n845), .ZN(new_n848));
  NAND3_X1  g662(.A1(new_n840), .A2(new_n846), .A3(new_n848), .ZN(new_n849));
  XNOR2_X1  g663(.A(new_n849), .B(G137), .ZN(G39));
  INV_X1    g664(.A(KEYINPUT47), .ZN(new_n851));
  NOR2_X1   g665(.A1(new_n851), .A2(KEYINPUT109), .ZN(new_n852));
  INV_X1    g666(.A(new_n852), .ZN(new_n853));
  NAND3_X1  g667(.A1(new_n838), .A2(new_n522), .A3(new_n853), .ZN(new_n854));
  OAI21_X1  g668(.A(new_n522), .B1(new_n836), .B2(new_n837), .ZN(new_n855));
  XNOR2_X1  g669(.A(KEYINPUT109), .B(KEYINPUT47), .ZN(new_n856));
  INV_X1    g670(.A(new_n856), .ZN(new_n857));
  NAND2_X1  g671(.A1(new_n855), .A2(new_n857), .ZN(new_n858));
  NOR4_X1   g672(.A1(new_n640), .A2(new_n578), .A3(new_n781), .A4(new_n847), .ZN(new_n859));
  NAND3_X1  g673(.A1(new_n854), .A2(new_n858), .A3(new_n859), .ZN(new_n860));
  XNOR2_X1  g674(.A(new_n860), .B(G140), .ZN(G42));
  NOR2_X1   g675(.A1(G952), .A2(G953), .ZN(new_n862));
  INV_X1    g676(.A(KEYINPUT52), .ZN(new_n863));
  INV_X1    g677(.A(KEYINPUT112), .ZN(new_n864));
  OAI21_X1  g678(.A(new_n522), .B1(new_n694), .B2(new_n864), .ZN(new_n865));
  AOI21_X1  g679(.A(new_n865), .B1(new_n864), .B2(new_n694), .ZN(new_n866));
  AND3_X1   g680(.A1(new_n813), .A2(new_n682), .A3(new_n866), .ZN(new_n867));
  AND3_X1   g681(.A1(new_n714), .A2(KEYINPUT102), .A3(new_n667), .ZN(new_n868));
  AOI21_X1  g682(.A(KEYINPUT102), .B1(new_n714), .B2(new_n667), .ZN(new_n869));
  OAI211_X1 g683(.A(new_n705), .B(new_n867), .C1(new_n868), .C2(new_n869), .ZN(new_n870));
  AND3_X1   g684(.A1(new_n723), .A2(new_n870), .A3(new_n697), .ZN(new_n871));
  AND3_X1   g685(.A1(new_n871), .A2(new_n806), .A3(KEYINPUT113), .ZN(new_n872));
  AOI21_X1  g686(.A(KEYINPUT113), .B1(new_n871), .B2(new_n806), .ZN(new_n873));
  OAI21_X1  g687(.A(new_n863), .B1(new_n872), .B2(new_n873), .ZN(new_n874));
  INV_X1    g688(.A(KEYINPUT113), .ZN(new_n875));
  NOR3_X1   g689(.A1(new_n785), .A2(new_n798), .A3(new_n780), .ZN(new_n876));
  AOI21_X1  g690(.A(KEYINPUT105), .B1(new_n802), .B2(new_n804), .ZN(new_n877));
  NOR2_X1   g691(.A1(new_n876), .A2(new_n877), .ZN(new_n878));
  NAND3_X1  g692(.A1(new_n723), .A2(new_n870), .A3(new_n697), .ZN(new_n879));
  OAI21_X1  g693(.A(new_n875), .B1(new_n878), .B2(new_n879), .ZN(new_n880));
  NAND3_X1  g694(.A1(new_n871), .A2(new_n806), .A3(KEYINPUT113), .ZN(new_n881));
  NAND3_X1  g695(.A1(new_n880), .A2(KEYINPUT52), .A3(new_n881), .ZN(new_n882));
  AND3_X1   g696(.A1(new_n376), .A2(new_n381), .A3(new_n439), .ZN(new_n883));
  OAI21_X1  g697(.A(new_n673), .B1(new_n883), .B2(new_n656), .ZN(new_n884));
  NAND2_X1  g698(.A1(new_n292), .A2(new_n294), .ZN(new_n885));
  NOR2_X1   g699(.A1(new_n884), .A2(new_n885), .ZN(new_n886));
  AOI22_X1  g700(.A1(new_n648), .A2(new_n886), .B1(new_n769), .B2(new_n776), .ZN(new_n887));
  NAND3_X1  g701(.A1(new_n762), .A2(new_n684), .A3(new_n685), .ZN(new_n888));
  AOI21_X1  g702(.A(new_n888), .B1(new_n619), .B2(new_n636), .ZN(new_n889));
  AOI22_X1  g703(.A1(new_n889), .A2(new_n752), .B1(new_n683), .B2(new_n686), .ZN(new_n890));
  OAI211_X1 g704(.A(new_n725), .B(new_n740), .C1(new_n658), .C2(new_n674), .ZN(new_n891));
  NAND4_X1  g705(.A1(new_n642), .A2(new_n887), .A3(new_n890), .A4(new_n891), .ZN(new_n892));
  AND4_X1   g706(.A1(new_n713), .A2(new_n672), .A3(new_n694), .A4(new_n814), .ZN(new_n893));
  NAND3_X1  g707(.A1(new_n893), .A2(new_n640), .A3(new_n690), .ZN(new_n894));
  NOR3_X1   g708(.A1(new_n682), .A2(new_n787), .A3(new_n796), .ZN(new_n895));
  NAND4_X1  g709(.A1(new_n783), .A2(new_n815), .A3(new_n895), .A4(new_n784), .ZN(new_n896));
  AND3_X1   g710(.A1(new_n829), .A2(new_n894), .A3(new_n896), .ZN(new_n897));
  INV_X1    g711(.A(new_n897), .ZN(new_n898));
  NOR3_X1   g712(.A1(new_n827), .A2(new_n892), .A3(new_n898), .ZN(new_n899));
  NAND3_X1  g713(.A1(new_n874), .A2(new_n882), .A3(new_n899), .ZN(new_n900));
  INV_X1    g714(.A(KEYINPUT53), .ZN(new_n901));
  NAND2_X1  g715(.A1(new_n900), .A2(new_n901), .ZN(new_n902));
  INV_X1    g716(.A(KEYINPUT54), .ZN(new_n903));
  NAND3_X1  g717(.A1(new_n376), .A2(new_n439), .A3(new_n381), .ZN(new_n904));
  AOI21_X1  g718(.A(new_n446), .B1(new_n657), .B2(new_n904), .ZN(new_n905));
  NOR2_X1   g719(.A1(new_n523), .A2(new_n579), .ZN(new_n906));
  INV_X1    g720(.A(new_n647), .ZN(new_n907));
  NAND4_X1  g721(.A1(new_n905), .A2(new_n906), .A3(new_n295), .A4(new_n907), .ZN(new_n908));
  AND4_X1   g722(.A1(new_n687), .A2(new_n777), .A3(new_n908), .A4(new_n763), .ZN(new_n909));
  NAND4_X1  g723(.A1(new_n909), .A2(new_n642), .A3(new_n891), .A4(new_n897), .ZN(new_n910));
  NOR3_X1   g724(.A1(new_n910), .A2(new_n901), .A3(new_n827), .ZN(new_n911));
  OAI21_X1  g725(.A(KEYINPUT52), .B1(new_n878), .B2(new_n879), .ZN(new_n912));
  NAND3_X1  g726(.A1(new_n911), .A2(new_n874), .A3(new_n912), .ZN(new_n913));
  AND3_X1   g727(.A1(new_n902), .A2(new_n903), .A3(new_n913), .ZN(new_n914));
  OAI21_X1  g728(.A(KEYINPUT111), .B1(new_n910), .B2(new_n827), .ZN(new_n915));
  NAND2_X1  g729(.A1(new_n825), .A2(new_n826), .ZN(new_n916));
  INV_X1    g730(.A(new_n817), .ZN(new_n917));
  NAND2_X1  g731(.A1(new_n916), .A2(new_n917), .ZN(new_n918));
  AND4_X1   g732(.A1(new_n642), .A2(new_n887), .A3(new_n890), .A4(new_n891), .ZN(new_n919));
  INV_X1    g733(.A(KEYINPUT111), .ZN(new_n920));
  NAND4_X1  g734(.A1(new_n918), .A2(new_n919), .A3(new_n920), .A4(new_n897), .ZN(new_n921));
  NAND4_X1  g735(.A1(new_n915), .A2(new_n921), .A3(new_n874), .A4(new_n912), .ZN(new_n922));
  NAND2_X1  g736(.A1(new_n922), .A2(new_n901), .ZN(new_n923));
  NAND3_X1  g737(.A1(new_n911), .A2(new_n874), .A3(new_n882), .ZN(new_n924));
  INV_X1    g738(.A(KEYINPUT114), .ZN(new_n925));
  NAND2_X1  g739(.A1(new_n924), .A2(new_n925), .ZN(new_n926));
  NAND4_X1  g740(.A1(new_n911), .A2(KEYINPUT114), .A3(new_n874), .A4(new_n882), .ZN(new_n927));
  NAND3_X1  g741(.A1(new_n923), .A2(new_n926), .A3(new_n927), .ZN(new_n928));
  AOI21_X1  g742(.A(new_n914), .B1(KEYINPUT54), .B2(new_n928), .ZN(new_n929));
  INV_X1    g743(.A(KEYINPUT117), .ZN(new_n930));
  NAND3_X1  g744(.A1(new_n842), .A2(new_n441), .A3(new_n843), .ZN(new_n931));
  NOR4_X1   g745(.A1(new_n931), .A2(KEYINPUT115), .A3(new_n775), .A4(new_n847), .ZN(new_n932));
  INV_X1    g746(.A(KEYINPUT115), .ZN(new_n933));
  NOR2_X1   g747(.A1(new_n931), .A2(new_n775), .ZN(new_n934));
  AOI21_X1  g748(.A(new_n933), .B1(new_n934), .B2(new_n814), .ZN(new_n935));
  NAND2_X1  g749(.A1(new_n854), .A2(new_n858), .ZN(new_n936));
  NAND2_X1  g750(.A1(new_n739), .A2(new_n737), .ZN(new_n937));
  AND2_X1   g751(.A1(new_n937), .A2(new_n511), .ZN(new_n938));
  NAND2_X1  g752(.A1(new_n938), .A2(new_n747), .ZN(new_n939));
  AOI211_X1 g753(.A(new_n932), .B(new_n935), .C1(new_n936), .C2(new_n939), .ZN(new_n940));
  AND3_X1   g754(.A1(new_n709), .A2(new_n662), .A3(new_n740), .ZN(new_n941));
  NAND2_X1  g755(.A1(new_n934), .A2(new_n941), .ZN(new_n942));
  INV_X1    g756(.A(KEYINPUT50), .ZN(new_n943));
  NAND2_X1  g757(.A1(new_n942), .A2(new_n943), .ZN(new_n944));
  NAND3_X1  g758(.A1(new_n934), .A2(KEYINPUT50), .A3(new_n941), .ZN(new_n945));
  NAND2_X1  g759(.A1(new_n944), .A2(new_n945), .ZN(new_n946));
  NAND2_X1  g760(.A1(new_n740), .A2(new_n814), .ZN(new_n947));
  NOR2_X1   g761(.A1(new_n931), .A2(new_n947), .ZN(new_n948));
  NAND3_X1  g762(.A1(new_n706), .A2(new_n578), .A3(new_n441), .ZN(new_n949));
  NOR2_X1   g763(.A1(new_n949), .A2(new_n947), .ZN(new_n950));
  NOR2_X1   g764(.A1(new_n382), .A2(new_n718), .ZN(new_n951));
  AOI22_X1  g765(.A1(new_n948), .A2(new_n895), .B1(new_n950), .B2(new_n951), .ZN(new_n952));
  NAND3_X1  g766(.A1(new_n946), .A2(KEYINPUT51), .A3(new_n952), .ZN(new_n953));
  OAI21_X1  g767(.A(new_n930), .B1(new_n940), .B2(new_n953), .ZN(new_n954));
  INV_X1    g768(.A(new_n952), .ZN(new_n955));
  AOI21_X1  g769(.A(new_n955), .B1(new_n944), .B2(new_n945), .ZN(new_n956));
  NAND2_X1  g770(.A1(new_n936), .A2(new_n939), .ZN(new_n957));
  NOR2_X1   g771(.A1(new_n935), .A2(new_n932), .ZN(new_n958));
  NAND2_X1  g772(.A1(new_n957), .A2(new_n958), .ZN(new_n959));
  NAND4_X1  g773(.A1(new_n956), .A2(new_n959), .A3(KEYINPUT117), .A4(KEYINPUT51), .ZN(new_n960));
  NAND2_X1  g774(.A1(new_n954), .A2(new_n960), .ZN(new_n961));
  INV_X1    g775(.A(KEYINPUT48), .ZN(new_n962));
  INV_X1    g776(.A(new_n825), .ZN(new_n963));
  INV_X1    g777(.A(new_n948), .ZN(new_n964));
  OAI21_X1  g778(.A(new_n962), .B1(new_n963), .B2(new_n964), .ZN(new_n965));
  NAND3_X1  g779(.A1(new_n825), .A2(new_n948), .A3(KEYINPUT48), .ZN(new_n966));
  NAND2_X1  g780(.A1(new_n950), .A2(new_n656), .ZN(new_n967));
  AOI21_X1  g781(.A(new_n440), .B1(new_n934), .B2(new_n752), .ZN(new_n968));
  NAND4_X1  g782(.A1(new_n965), .A2(new_n966), .A3(new_n967), .A4(new_n968), .ZN(new_n969));
  INV_X1    g783(.A(new_n958), .ZN(new_n970));
  XNOR2_X1  g784(.A(new_n939), .B(KEYINPUT116), .ZN(new_n971));
  AOI21_X1  g785(.A(new_n971), .B1(new_n854), .B2(new_n858), .ZN(new_n972));
  OAI21_X1  g786(.A(new_n956), .B1(new_n970), .B2(new_n972), .ZN(new_n973));
  INV_X1    g787(.A(KEYINPUT51), .ZN(new_n974));
  AOI21_X1  g788(.A(new_n969), .B1(new_n973), .B2(new_n974), .ZN(new_n975));
  AND2_X1   g789(.A1(new_n961), .A2(new_n975), .ZN(new_n976));
  AOI21_X1  g790(.A(new_n862), .B1(new_n929), .B2(new_n976), .ZN(new_n977));
  NAND3_X1  g791(.A1(new_n578), .A2(new_n187), .A3(new_n522), .ZN(new_n978));
  INV_X1    g792(.A(new_n938), .ZN(new_n979));
  AOI211_X1 g793(.A(new_n841), .B(new_n978), .C1(new_n979), .C2(KEYINPUT49), .ZN(new_n980));
  XOR2_X1   g794(.A(new_n980), .B(KEYINPUT110), .Z(new_n981));
  OAI211_X1 g795(.A(new_n706), .B(new_n709), .C1(new_n979), .C2(KEYINPUT49), .ZN(new_n982));
  NOR2_X1   g796(.A1(new_n981), .A2(new_n982), .ZN(new_n983));
  OAI21_X1  g797(.A(KEYINPUT118), .B1(new_n977), .B2(new_n983), .ZN(new_n984));
  NAND2_X1  g798(.A1(new_n928), .A2(KEYINPUT54), .ZN(new_n985));
  NAND3_X1  g799(.A1(new_n902), .A2(new_n903), .A3(new_n913), .ZN(new_n986));
  NAND3_X1  g800(.A1(new_n985), .A2(new_n976), .A3(new_n986), .ZN(new_n987));
  INV_X1    g801(.A(new_n862), .ZN(new_n988));
  NAND2_X1  g802(.A1(new_n987), .A2(new_n988), .ZN(new_n989));
  INV_X1    g803(.A(KEYINPUT118), .ZN(new_n990));
  INV_X1    g804(.A(new_n983), .ZN(new_n991));
  NAND3_X1  g805(.A1(new_n989), .A2(new_n990), .A3(new_n991), .ZN(new_n992));
  NAND2_X1  g806(.A1(new_n984), .A2(new_n992), .ZN(G75));
  OR2_X1    g807(.A1(new_n257), .A2(G952), .ZN(new_n994));
  XOR2_X1   g808(.A(new_n994), .B(KEYINPUT120), .Z(new_n995));
  AOI21_X1  g809(.A(new_n286), .B1(new_n902), .B2(new_n913), .ZN(new_n996));
  AOI21_X1  g810(.A(KEYINPUT56), .B1(new_n996), .B2(G210), .ZN(new_n997));
  NAND2_X1  g811(.A1(new_n232), .A2(new_n267), .ZN(new_n998));
  XNOR2_X1  g812(.A(new_n998), .B(new_n265), .ZN(new_n999));
  XNOR2_X1  g813(.A(new_n999), .B(KEYINPUT55), .ZN(new_n1000));
  OAI21_X1  g814(.A(new_n995), .B1(new_n997), .B2(new_n1000), .ZN(new_n1001));
  NAND2_X1  g815(.A1(new_n997), .A2(new_n1000), .ZN(new_n1002));
  INV_X1    g816(.A(KEYINPUT119), .ZN(new_n1003));
  NAND2_X1  g817(.A1(new_n1002), .A2(new_n1003), .ZN(new_n1004));
  NAND3_X1  g818(.A1(new_n997), .A2(KEYINPUT119), .A3(new_n1000), .ZN(new_n1005));
  AOI21_X1  g819(.A(new_n1001), .B1(new_n1004), .B2(new_n1005), .ZN(G51));
  INV_X1    g820(.A(new_n995), .ZN(new_n1007));
  AOI211_X1 g821(.A(new_n286), .B(new_n832), .C1(new_n902), .C2(new_n913), .ZN(new_n1008));
  INV_X1    g822(.A(new_n509), .ZN(new_n1009));
  NAND2_X1  g823(.A1(new_n902), .A2(new_n913), .ZN(new_n1010));
  NAND2_X1  g824(.A1(new_n1010), .A2(KEYINPUT54), .ZN(new_n1011));
  NAND2_X1  g825(.A1(new_n1011), .A2(new_n986), .ZN(new_n1012));
  XOR2_X1   g826(.A(new_n512), .B(KEYINPUT121), .Z(new_n1013));
  XOR2_X1   g827(.A(new_n1013), .B(KEYINPUT57), .Z(new_n1014));
  AOI21_X1  g828(.A(new_n1009), .B1(new_n1012), .B2(new_n1014), .ZN(new_n1015));
  AOI21_X1  g829(.A(new_n1008), .B1(new_n1015), .B2(KEYINPUT122), .ZN(new_n1016));
  INV_X1    g830(.A(KEYINPUT122), .ZN(new_n1017));
  INV_X1    g831(.A(new_n1014), .ZN(new_n1018));
  AOI21_X1  g832(.A(new_n1018), .B1(new_n1011), .B2(new_n986), .ZN(new_n1019));
  OAI21_X1  g833(.A(new_n1017), .B1(new_n1019), .B2(new_n1009), .ZN(new_n1020));
  AOI21_X1  g834(.A(new_n1007), .B1(new_n1016), .B2(new_n1020), .ZN(G54));
  AND3_X1   g835(.A1(new_n996), .A2(KEYINPUT58), .A3(G475), .ZN(new_n1022));
  INV_X1    g836(.A(new_n373), .ZN(new_n1023));
  OR2_X1    g837(.A1(new_n1022), .A2(new_n1023), .ZN(new_n1024));
  NAND2_X1  g838(.A1(new_n1022), .A2(new_n1023), .ZN(new_n1025));
  AOI21_X1  g839(.A(new_n1007), .B1(new_n1024), .B2(new_n1025), .ZN(G60));
  INV_X1    g840(.A(new_n1012), .ZN(new_n1027));
  AND2_X1   g841(.A1(new_n650), .A2(new_n651), .ZN(new_n1028));
  XNOR2_X1  g842(.A(new_n653), .B(KEYINPUT59), .ZN(new_n1029));
  OR2_X1    g843(.A1(new_n1028), .A2(new_n1029), .ZN(new_n1030));
  OAI21_X1  g844(.A(new_n995), .B1(new_n1027), .B2(new_n1030), .ZN(new_n1031));
  OR2_X1    g845(.A1(new_n929), .A2(new_n1029), .ZN(new_n1032));
  AOI21_X1  g846(.A(new_n1031), .B1(new_n1032), .B2(new_n1028), .ZN(G63));
  NAND2_X1  g847(.A1(G217), .A2(G902), .ZN(new_n1034));
  XOR2_X1   g848(.A(new_n1034), .B(KEYINPUT60), .Z(new_n1035));
  NAND2_X1  g849(.A1(new_n1010), .A2(new_n1035), .ZN(new_n1036));
  INV_X1    g850(.A(new_n1036), .ZN(new_n1037));
  NOR2_X1   g851(.A1(new_n679), .A2(new_n680), .ZN(new_n1038));
  AOI21_X1  g852(.A(KEYINPUT124), .B1(new_n1037), .B2(new_n1038), .ZN(new_n1039));
  NOR2_X1   g853(.A1(new_n1039), .A2(KEYINPUT61), .ZN(new_n1040));
  AOI21_X1  g854(.A(new_n1007), .B1(new_n1037), .B2(new_n1038), .ZN(new_n1041));
  XNOR2_X1  g855(.A(new_n757), .B(KEYINPUT123), .ZN(new_n1042));
  NAND2_X1  g856(.A1(new_n1036), .A2(new_n1042), .ZN(new_n1043));
  NAND2_X1  g857(.A1(new_n1041), .A2(new_n1043), .ZN(new_n1044));
  NAND2_X1  g858(.A1(new_n1040), .A2(new_n1044), .ZN(new_n1045));
  OAI211_X1 g859(.A(new_n1043), .B(new_n1041), .C1(new_n1039), .C2(KEYINPUT61), .ZN(new_n1046));
  NAND2_X1  g860(.A1(new_n1045), .A2(new_n1046), .ZN(G66));
  NAND2_X1  g861(.A1(new_n892), .A2(new_n257), .ZN(new_n1048));
  XOR2_X1   g862(.A(new_n1048), .B(KEYINPUT125), .Z(new_n1049));
  INV_X1    g863(.A(G224), .ZN(new_n1050));
  OAI21_X1  g864(.A(G953), .B1(new_n445), .B2(new_n1050), .ZN(new_n1051));
  NAND2_X1  g865(.A1(new_n1049), .A2(new_n1051), .ZN(new_n1052));
  OAI21_X1  g866(.A(new_n998), .B1(G898), .B2(new_n257), .ZN(new_n1053));
  XNOR2_X1  g867(.A(new_n1052), .B(new_n1053), .ZN(G69));
  NAND2_X1  g868(.A1(new_n602), .A2(new_n604), .ZN(new_n1055));
  XNOR2_X1  g869(.A(new_n1055), .B(new_n344), .ZN(new_n1056));
  OAI21_X1  g870(.A(new_n1056), .B1(new_n692), .B2(new_n257), .ZN(new_n1057));
  AND3_X1   g871(.A1(new_n806), .A2(new_n697), .A3(new_n723), .ZN(new_n1058));
  AND4_X1   g872(.A1(new_n829), .A2(new_n849), .A3(new_n860), .A4(new_n1058), .ZN(new_n1059));
  NAND3_X1  g873(.A1(new_n840), .A2(new_n769), .A3(new_n825), .ZN(new_n1060));
  AND3_X1   g874(.A1(new_n1059), .A2(new_n918), .A3(new_n1060), .ZN(new_n1061));
  AOI21_X1  g875(.A(new_n1057), .B1(new_n1061), .B2(new_n257), .ZN(new_n1062));
  NAND2_X1  g876(.A1(new_n716), .A2(new_n1058), .ZN(new_n1063));
  OR2_X1    g877(.A1(new_n1063), .A2(KEYINPUT62), .ZN(new_n1064));
  NAND2_X1  g878(.A1(new_n1063), .A2(KEYINPUT62), .ZN(new_n1065));
  AOI211_X1 g879(.A(new_n847), .B(new_n700), .C1(new_n657), .C2(new_n904), .ZN(new_n1066));
  OAI21_X1  g880(.A(new_n1066), .B1(new_n641), .B2(new_n637), .ZN(new_n1067));
  XNOR2_X1  g881(.A(new_n1067), .B(KEYINPUT126), .ZN(new_n1068));
  AND2_X1   g882(.A1(new_n849), .A2(new_n860), .ZN(new_n1069));
  NAND4_X1  g883(.A1(new_n1064), .A2(new_n1065), .A3(new_n1068), .A4(new_n1069), .ZN(new_n1070));
  AOI21_X1  g884(.A(new_n1056), .B1(new_n1070), .B2(new_n257), .ZN(new_n1071));
  NOR2_X1   g885(.A1(new_n1062), .A2(new_n1071), .ZN(new_n1072));
  OAI21_X1  g886(.A(G953), .B1(new_n491), .B2(new_n692), .ZN(new_n1073));
  XNOR2_X1  g887(.A(new_n1072), .B(new_n1073), .ZN(G72));
  AND2_X1   g888(.A1(new_n1061), .A2(new_n919), .ZN(new_n1075));
  NAND2_X1  g889(.A1(G472), .A2(G902), .ZN(new_n1076));
  XOR2_X1   g890(.A(new_n1076), .B(KEYINPUT63), .Z(new_n1077));
  INV_X1    g891(.A(new_n1077), .ZN(new_n1078));
  OAI21_X1  g892(.A(new_n622), .B1(new_n1075), .B2(new_n1078), .ZN(new_n1079));
  OAI21_X1  g893(.A(new_n1077), .B1(new_n1070), .B2(new_n892), .ZN(new_n1080));
  AOI21_X1  g894(.A(new_n1007), .B1(new_n1080), .B2(new_n702), .ZN(new_n1081));
  NAND2_X1  g895(.A1(new_n1079), .A2(new_n1081), .ZN(new_n1082));
  NOR3_X1   g896(.A1(new_n622), .A2(new_n702), .A3(new_n1078), .ZN(new_n1083));
  XOR2_X1   g897(.A(new_n1083), .B(KEYINPUT127), .Z(new_n1084));
  AOI21_X1  g898(.A(new_n1082), .B1(new_n928), .B2(new_n1084), .ZN(G57));
endmodule


