

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589,
         n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, n600,
         n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, n611,
         n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, n622,
         n623, n624, n625, n626, n627, n628, n629, n630, n631, n632, n633,
         n634, n635, n636, n637, n638, n639, n640, n641, n642, n643, n644,
         n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, n655,
         n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666,
         n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, n677,
         n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688,
         n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n699,
         n700, n701, n702, n703, n704, n705, n706, n707, n708, n709, n710,
         n711, n712, n713, n714, n715, n716, n717, n718, n719, n720, n721,
         n722, n723, n724, n725, n726, n727, n728, n729, n730, n731, n732,
         n733, n734, n735, n736, n737, n738, n739, n740, n741, n742, n743,
         n744, n745, n746, n747, n748, n749, n750, n751, n752, n753, n754,
         n755, n756, n757, n758, n759, n760, n761, n762, n763, n764, n765,
         n766, n767, n768, n769, n770, n771, n772, n773, n774, n775, n776,
         n777, n778, n779, n780, n781, n782, n783, n784, n785, n786, n787,
         n788, n789, n790, n791, n792, n793, n794, n795, n796, n797, n798,
         n799, n800, n801, n802, n803, n804, n805, n806, n807, n808, n809,
         n810, n811, n812, n813, n814, n815, n816, n817, n818, n819, n820,
         n821, n822, n823, n824, n825, n826, n827, n828, n829, n830, n831,
         n832, n833, n834, n835, n836, n837, n838, n839, n840, n841, n842,
         n843, n844, n845, n846, n847, n848, n849, n850, n851, n852, n853,
         n854, n855, n856, n857, n858, n859, n860, n861, n862, n863, n864,
         n865, n866, n867, n868, n869, n870, n871, n872, n873, n874, n875,
         n876, n877, n878, n879, n880, n881, n882, n883, n884, n885, n886,
         n887, n888, n889, n890, n891, n892, n893, n894, n895, n896, n897,
         n898, n899, n900, n901, n902, n903, n904, n905, n906, n907, n908,
         n909, n910, n911, n912, n913, n914, n915, n916, n917, n918, n919,
         n920, n921, n922, n923, n924, n925, n926, n927, n928, n929, n930,
         n931, n932, n933, n934, n935, n936, n937, n938, n939, n940, n941,
         n942, n943, n944, n945, n946, n947, n948, n949, n950, n951, n952,
         n953, n954, n955, n956, n957, n958, n959, n960, n961, n962, n963,
         n964, n965, n966, n967, n968, n969, n970, n971, n972, n973, n974,
         n975, n976, n977, n978, n979, n980, n981, n982, n983, n984, n985,
         n986, n987, n988, n989, n990, n991, n992, n993, n994, n995, n996,
         n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006,
         n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016,
         n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026,
         n1027, n1028, n1029, n1030, n1031, n1032;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NOR2_X2 U556 ( .A1(n790), .A2(n789), .ZN(n801) );
  OR2_X1 U557 ( .A1(n723), .A2(n722), .ZN(n721) );
  NOR2_X1 U558 ( .A1(n715), .A2(n930), .ZN(n717) );
  BUF_X1 U559 ( .A(n562), .Z(n520) );
  XNOR2_X1 U560 ( .A(KEYINPUT65), .B(n551), .ZN(n562) );
  NOR2_X1 U561 ( .A1(G1966), .A2(n797), .ZN(n769) );
  INV_X1 U562 ( .A(n936), .ZN(n777) );
  NOR2_X2 U563 ( .A1(n624), .A2(n548), .ZN(n571) );
  XNOR2_X2 U564 ( .A(n527), .B(n526), .ZN(n608) );
  XOR2_X1 U565 ( .A(KEYINPUT12), .B(n573), .Z(n521) );
  XOR2_X1 U566 ( .A(KEYINPUT14), .B(n576), .Z(n522) );
  OR2_X1 U567 ( .A1(n777), .A2(n797), .ZN(n523) );
  NAND2_X1 U568 ( .A1(n798), .A2(n797), .ZN(n524) );
  INV_X1 U569 ( .A(KEYINPUT64), .ZN(n716) );
  INV_X1 U570 ( .A(KEYINPUT29), .ZN(n738) );
  XNOR2_X1 U571 ( .A(n752), .B(KEYINPUT96), .ZN(n753) );
  XNOR2_X1 U572 ( .A(n754), .B(n753), .ZN(n755) );
  AND2_X1 U573 ( .A1(n764), .A2(n763), .ZN(n765) );
  OR2_X1 U574 ( .A1(n778), .A2(n523), .ZN(n779) );
  INV_X1 U575 ( .A(n925), .ZN(n787) );
  OR2_X1 U576 ( .A1(n788), .A2(n787), .ZN(n789) );
  INV_X1 U577 ( .A(KEYINPUT99), .ZN(n802) );
  INV_X1 U578 ( .A(KEYINPUT17), .ZN(n525) );
  XNOR2_X1 U579 ( .A(n803), .B(n802), .ZN(n804) );
  XNOR2_X1 U580 ( .A(n525), .B(KEYINPUT68), .ZN(n526) );
  NOR2_X1 U581 ( .A1(n805), .A2(n804), .ZN(n807) );
  NOR2_X1 U582 ( .A1(G651), .A2(G543), .ZN(n656) );
  AND2_X1 U583 ( .A1(n530), .A2(G2104), .ZN(n902) );
  NAND2_X1 U584 ( .A1(n580), .A2(n579), .ZN(n930) );
  NOR2_X1 U585 ( .A1(n535), .A2(n534), .ZN(G164) );
  INV_X1 U586 ( .A(G2105), .ZN(n530) );
  NAND2_X1 U587 ( .A1(n902), .A2(G102), .ZN(n529) );
  NOR2_X1 U588 ( .A1(G2104), .A2(G2105), .ZN(n527) );
  NAND2_X1 U589 ( .A1(G138), .A2(n608), .ZN(n528) );
  NAND2_X1 U590 ( .A1(n529), .A2(n528), .ZN(n535) );
  NOR2_X1 U591 ( .A1(G2104), .A2(n530), .ZN(n898) );
  NAND2_X1 U592 ( .A1(G126), .A2(n898), .ZN(n533) );
  NAND2_X1 U593 ( .A1(G2104), .A2(G2105), .ZN(n531) );
  XOR2_X1 U594 ( .A(KEYINPUT66), .B(n531), .Z(n609) );
  NAND2_X1 U595 ( .A1(G114), .A2(n609), .ZN(n532) );
  NAND2_X1 U596 ( .A1(n533), .A2(n532), .ZN(n534) );
  NAND2_X1 U597 ( .A1(n609), .A2(G113), .ZN(n536) );
  XOR2_X1 U598 ( .A(n536), .B(KEYINPUT67), .Z(n539) );
  NAND2_X1 U599 ( .A1(G101), .A2(n902), .ZN(n537) );
  XOR2_X1 U600 ( .A(KEYINPUT23), .B(n537), .Z(n538) );
  NAND2_X1 U601 ( .A1(n539), .A2(n538), .ZN(n543) );
  NAND2_X1 U602 ( .A1(n898), .A2(G125), .ZN(n541) );
  NAND2_X1 U603 ( .A1(G137), .A2(n608), .ZN(n540) );
  NAND2_X1 U604 ( .A1(n541), .A2(n540), .ZN(n542) );
  NOR2_X2 U605 ( .A1(n543), .A2(n542), .ZN(G160) );
  AND2_X1 U606 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U607 ( .A(G57), .ZN(G237) );
  XNOR2_X1 U608 ( .A(KEYINPUT71), .B(KEYINPUT1), .ZN(n545) );
  INV_X1 U609 ( .A(G651), .ZN(n548) );
  NOR2_X1 U610 ( .A1(G543), .A2(n548), .ZN(n544) );
  XNOR2_X1 U611 ( .A(n545), .B(n544), .ZN(n649) );
  NAND2_X1 U612 ( .A1(G65), .A2(n649), .ZN(n546) );
  XNOR2_X1 U613 ( .A(n546), .B(KEYINPUT72), .ZN(n556) );
  XNOR2_X1 U614 ( .A(G543), .B(KEYINPUT0), .ZN(n547) );
  XNOR2_X1 U615 ( .A(n547), .B(KEYINPUT69), .ZN(n624) );
  NAND2_X1 U616 ( .A1(G78), .A2(n571), .ZN(n550) );
  NAND2_X1 U617 ( .A1(G91), .A2(n656), .ZN(n549) );
  NAND2_X1 U618 ( .A1(n550), .A2(n549), .ZN(n554) );
  OR2_X1 U619 ( .A1(G651), .A2(n624), .ZN(n551) );
  NAND2_X1 U620 ( .A1(G53), .A2(n562), .ZN(n552) );
  XNOR2_X1 U621 ( .A(KEYINPUT73), .B(n552), .ZN(n553) );
  NOR2_X1 U622 ( .A1(n554), .A2(n553), .ZN(n555) );
  NAND2_X1 U623 ( .A1(n556), .A2(n555), .ZN(n557) );
  XNOR2_X1 U624 ( .A(KEYINPUT74), .B(n557), .ZN(G299) );
  NAND2_X1 U625 ( .A1(n656), .A2(G89), .ZN(n558) );
  XNOR2_X1 U626 ( .A(n558), .B(KEYINPUT4), .ZN(n560) );
  NAND2_X1 U627 ( .A1(G76), .A2(n571), .ZN(n559) );
  NAND2_X1 U628 ( .A1(n560), .A2(n559), .ZN(n561) );
  XNOR2_X1 U629 ( .A(n561), .B(KEYINPUT5), .ZN(n567) );
  NAND2_X1 U630 ( .A1(G63), .A2(n649), .ZN(n564) );
  NAND2_X1 U631 ( .A1(G51), .A2(n520), .ZN(n563) );
  NAND2_X1 U632 ( .A1(n564), .A2(n563), .ZN(n565) );
  XOR2_X1 U633 ( .A(KEYINPUT6), .B(n565), .Z(n566) );
  NAND2_X1 U634 ( .A1(n567), .A2(n566), .ZN(n568) );
  XNOR2_X1 U635 ( .A(n568), .B(KEYINPUT7), .ZN(G168) );
  XOR2_X1 U636 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U637 ( .A1(G7), .A2(G661), .ZN(n569) );
  XNOR2_X1 U638 ( .A(n569), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U639 ( .A(G223), .ZN(n836) );
  NAND2_X1 U640 ( .A1(n836), .A2(G567), .ZN(n570) );
  XOR2_X1 U641 ( .A(KEYINPUT11), .B(n570), .Z(G234) );
  NAND2_X1 U642 ( .A1(n571), .A2(G68), .ZN(n572) );
  XNOR2_X1 U643 ( .A(KEYINPUT75), .B(n572), .ZN(n574) );
  NAND2_X1 U644 ( .A1(n656), .A2(G81), .ZN(n573) );
  NOR2_X1 U645 ( .A1(n574), .A2(n521), .ZN(n575) );
  XNOR2_X1 U646 ( .A(n575), .B(KEYINPUT13), .ZN(n577) );
  NAND2_X1 U647 ( .A1(n649), .A2(G56), .ZN(n576) );
  NOR2_X1 U648 ( .A1(n577), .A2(n522), .ZN(n578) );
  XNOR2_X1 U649 ( .A(n578), .B(KEYINPUT76), .ZN(n580) );
  NAND2_X1 U650 ( .A1(G43), .A2(n520), .ZN(n579) );
  INV_X1 U651 ( .A(G860), .ZN(n841) );
  OR2_X1 U652 ( .A1(n930), .A2(n841), .ZN(G153) );
  NAND2_X1 U653 ( .A1(G77), .A2(n571), .ZN(n582) );
  NAND2_X1 U654 ( .A1(G90), .A2(n656), .ZN(n581) );
  NAND2_X1 U655 ( .A1(n582), .A2(n581), .ZN(n583) );
  XNOR2_X1 U656 ( .A(KEYINPUT9), .B(n583), .ZN(n587) );
  NAND2_X1 U657 ( .A1(G64), .A2(n649), .ZN(n585) );
  NAND2_X1 U658 ( .A1(G52), .A2(n520), .ZN(n584) );
  AND2_X1 U659 ( .A1(n585), .A2(n584), .ZN(n586) );
  NAND2_X1 U660 ( .A1(n587), .A2(n586), .ZN(G301) );
  NAND2_X1 U661 ( .A1(G868), .A2(G301), .ZN(n597) );
  NAND2_X1 U662 ( .A1(G92), .A2(n656), .ZN(n589) );
  NAND2_X1 U663 ( .A1(G66), .A2(n649), .ZN(n588) );
  NAND2_X1 U664 ( .A1(n589), .A2(n588), .ZN(n594) );
  NAND2_X1 U665 ( .A1(G79), .A2(n571), .ZN(n591) );
  NAND2_X1 U666 ( .A1(G54), .A2(n520), .ZN(n590) );
  NAND2_X1 U667 ( .A1(n591), .A2(n590), .ZN(n592) );
  XOR2_X1 U668 ( .A(KEYINPUT77), .B(n592), .Z(n593) );
  NOR2_X1 U669 ( .A1(n594), .A2(n593), .ZN(n595) );
  XNOR2_X1 U670 ( .A(KEYINPUT15), .B(n595), .ZN(n722) );
  INV_X1 U671 ( .A(G868), .ZN(n667) );
  NAND2_X1 U672 ( .A1(n722), .A2(n667), .ZN(n596) );
  NAND2_X1 U673 ( .A1(n597), .A2(n596), .ZN(G284) );
  NOR2_X1 U674 ( .A1(G286), .A2(n667), .ZN(n599) );
  NOR2_X1 U675 ( .A1(G299), .A2(G868), .ZN(n598) );
  NOR2_X1 U676 ( .A1(n599), .A2(n598), .ZN(G297) );
  NAND2_X1 U677 ( .A1(n841), .A2(G559), .ZN(n600) );
  INV_X1 U678 ( .A(n722), .ZN(n924) );
  NAND2_X1 U679 ( .A1(n600), .A2(n924), .ZN(n601) );
  XNOR2_X1 U680 ( .A(n601), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U681 ( .A1(G868), .A2(n930), .ZN(n604) );
  NAND2_X1 U682 ( .A1(G868), .A2(n924), .ZN(n602) );
  NOR2_X1 U683 ( .A1(G559), .A2(n602), .ZN(n603) );
  NOR2_X1 U684 ( .A1(n604), .A2(n603), .ZN(G282) );
  NAND2_X1 U685 ( .A1(G123), .A2(n898), .ZN(n605) );
  XNOR2_X1 U686 ( .A(n605), .B(KEYINPUT18), .ZN(n607) );
  NAND2_X1 U687 ( .A1(n902), .A2(G99), .ZN(n606) );
  NAND2_X1 U688 ( .A1(n607), .A2(n606), .ZN(n613) );
  NAND2_X1 U689 ( .A1(G135), .A2(n608), .ZN(n611) );
  BUF_X1 U690 ( .A(n609), .Z(n899) );
  NAND2_X1 U691 ( .A1(G111), .A2(n899), .ZN(n610) );
  NAND2_X1 U692 ( .A1(n611), .A2(n610), .ZN(n612) );
  NOR2_X1 U693 ( .A1(n613), .A2(n612), .ZN(n969) );
  XOR2_X1 U694 ( .A(n969), .B(G2096), .Z(n614) );
  NOR2_X1 U695 ( .A1(G2100), .A2(n614), .ZN(n615) );
  XOR2_X1 U696 ( .A(KEYINPUT78), .B(n615), .Z(G156) );
  NAND2_X1 U697 ( .A1(G88), .A2(n656), .ZN(n616) );
  XNOR2_X1 U698 ( .A(n616), .B(KEYINPUT86), .ZN(n623) );
  NAND2_X1 U699 ( .A1(G75), .A2(n571), .ZN(n618) );
  NAND2_X1 U700 ( .A1(G62), .A2(n649), .ZN(n617) );
  NAND2_X1 U701 ( .A1(n618), .A2(n617), .ZN(n621) );
  NAND2_X1 U702 ( .A1(G50), .A2(n520), .ZN(n619) );
  XNOR2_X1 U703 ( .A(KEYINPUT85), .B(n619), .ZN(n620) );
  NOR2_X1 U704 ( .A1(n621), .A2(n620), .ZN(n622) );
  NAND2_X1 U705 ( .A1(n623), .A2(n622), .ZN(G303) );
  INV_X1 U706 ( .A(G303), .ZN(G166) );
  NAND2_X1 U707 ( .A1(G49), .A2(n520), .ZN(n626) );
  NAND2_X1 U708 ( .A1(G87), .A2(n624), .ZN(n625) );
  NAND2_X1 U709 ( .A1(n626), .A2(n625), .ZN(n627) );
  NOR2_X1 U710 ( .A1(n649), .A2(n627), .ZN(n629) );
  NAND2_X1 U711 ( .A1(G651), .A2(G74), .ZN(n628) );
  NAND2_X1 U712 ( .A1(n629), .A2(n628), .ZN(G288) );
  NAND2_X1 U713 ( .A1(G48), .A2(n520), .ZN(n630) );
  XNOR2_X1 U714 ( .A(n630), .B(KEYINPUT84), .ZN(n638) );
  NAND2_X1 U715 ( .A1(n571), .A2(G73), .ZN(n631) );
  XNOR2_X1 U716 ( .A(n631), .B(KEYINPUT2), .ZN(n633) );
  NAND2_X1 U717 ( .A1(G61), .A2(n649), .ZN(n632) );
  NAND2_X1 U718 ( .A1(n633), .A2(n632), .ZN(n636) );
  NAND2_X1 U719 ( .A1(G86), .A2(n656), .ZN(n634) );
  XNOR2_X1 U720 ( .A(KEYINPUT83), .B(n634), .ZN(n635) );
  NOR2_X1 U721 ( .A1(n636), .A2(n635), .ZN(n637) );
  NAND2_X1 U722 ( .A1(n638), .A2(n637), .ZN(G305) );
  NAND2_X1 U723 ( .A1(G85), .A2(n656), .ZN(n640) );
  NAND2_X1 U724 ( .A1(G60), .A2(n649), .ZN(n639) );
  NAND2_X1 U725 ( .A1(n640), .A2(n639), .ZN(n643) );
  NAND2_X1 U726 ( .A1(G72), .A2(n571), .ZN(n641) );
  XOR2_X1 U727 ( .A(KEYINPUT70), .B(n641), .Z(n642) );
  NOR2_X1 U728 ( .A1(n643), .A2(n642), .ZN(n645) );
  NAND2_X1 U729 ( .A1(n520), .A2(G47), .ZN(n644) );
  NAND2_X1 U730 ( .A1(n645), .A2(n644), .ZN(G290) );
  XNOR2_X1 U731 ( .A(KEYINPUT19), .B(KEYINPUT88), .ZN(n647) );
  XNOR2_X1 U732 ( .A(G288), .B(KEYINPUT87), .ZN(n646) );
  XNOR2_X1 U733 ( .A(n647), .B(n646), .ZN(n648) );
  XNOR2_X1 U734 ( .A(n648), .B(G305), .ZN(n661) );
  NAND2_X1 U735 ( .A1(n649), .A2(G67), .ZN(n650) );
  XNOR2_X1 U736 ( .A(n650), .B(KEYINPUT80), .ZN(n652) );
  NAND2_X1 U737 ( .A1(G55), .A2(n520), .ZN(n651) );
  NAND2_X1 U738 ( .A1(n652), .A2(n651), .ZN(n653) );
  XNOR2_X1 U739 ( .A(n653), .B(KEYINPUT81), .ZN(n655) );
  NAND2_X1 U740 ( .A1(G80), .A2(n571), .ZN(n654) );
  NAND2_X1 U741 ( .A1(n655), .A2(n654), .ZN(n659) );
  NAND2_X1 U742 ( .A1(G93), .A2(n656), .ZN(n657) );
  XNOR2_X1 U743 ( .A(KEYINPUT79), .B(n657), .ZN(n658) );
  NOR2_X1 U744 ( .A1(n659), .A2(n658), .ZN(n660) );
  XOR2_X1 U745 ( .A(KEYINPUT82), .B(n660), .Z(n842) );
  XOR2_X1 U746 ( .A(n661), .B(n842), .Z(n662) );
  XNOR2_X1 U747 ( .A(G166), .B(n662), .ZN(n664) );
  XNOR2_X1 U748 ( .A(G290), .B(G299), .ZN(n663) );
  XNOR2_X1 U749 ( .A(n664), .B(n663), .ZN(n846) );
  NAND2_X1 U750 ( .A1(G559), .A2(n924), .ZN(n665) );
  XOR2_X1 U751 ( .A(n930), .B(n665), .Z(n840) );
  XOR2_X1 U752 ( .A(n846), .B(n840), .Z(n666) );
  NOR2_X1 U753 ( .A1(n667), .A2(n666), .ZN(n669) );
  NOR2_X1 U754 ( .A1(n842), .A2(G868), .ZN(n668) );
  NOR2_X1 U755 ( .A1(n669), .A2(n668), .ZN(G295) );
  NAND2_X1 U756 ( .A1(G2084), .A2(G2078), .ZN(n670) );
  XOR2_X1 U757 ( .A(KEYINPUT20), .B(n670), .Z(n671) );
  NAND2_X1 U758 ( .A1(G2090), .A2(n671), .ZN(n672) );
  XNOR2_X1 U759 ( .A(KEYINPUT21), .B(n672), .ZN(n673) );
  NAND2_X1 U760 ( .A1(n673), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U761 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  XOR2_X1 U762 ( .A(KEYINPUT89), .B(KEYINPUT22), .Z(n675) );
  NAND2_X1 U763 ( .A1(G132), .A2(G82), .ZN(n674) );
  XNOR2_X1 U764 ( .A(n675), .B(n674), .ZN(n676) );
  NOR2_X1 U765 ( .A1(n676), .A2(G218), .ZN(n677) );
  NAND2_X1 U766 ( .A1(G96), .A2(n677), .ZN(n845) );
  NAND2_X1 U767 ( .A1(n845), .A2(G2106), .ZN(n682) );
  NAND2_X1 U768 ( .A1(G120), .A2(G108), .ZN(n678) );
  NOR2_X1 U769 ( .A1(G237), .A2(n678), .ZN(n679) );
  NAND2_X1 U770 ( .A1(G69), .A2(n679), .ZN(n844) );
  NAND2_X1 U771 ( .A1(G567), .A2(n844), .ZN(n680) );
  XNOR2_X1 U772 ( .A(KEYINPUT90), .B(n680), .ZN(n681) );
  NAND2_X1 U773 ( .A1(n682), .A2(n681), .ZN(n851) );
  NAND2_X1 U774 ( .A1(G661), .A2(G483), .ZN(n683) );
  NOR2_X1 U775 ( .A1(n851), .A2(n683), .ZN(n839) );
  NAND2_X1 U776 ( .A1(n839), .A2(G36), .ZN(G176) );
  NOR2_X1 U777 ( .A1(G164), .A2(G1384), .ZN(n710) );
  NAND2_X1 U778 ( .A1(G160), .A2(G40), .ZN(n684) );
  NOR2_X1 U779 ( .A1(n710), .A2(n684), .ZN(n820) );
  NAND2_X1 U780 ( .A1(n898), .A2(G129), .ZN(n686) );
  NAND2_X1 U781 ( .A1(G141), .A2(n608), .ZN(n685) );
  NAND2_X1 U782 ( .A1(n686), .A2(n685), .ZN(n689) );
  NAND2_X1 U783 ( .A1(n902), .A2(G105), .ZN(n687) );
  XOR2_X1 U784 ( .A(KEYINPUT38), .B(n687), .Z(n688) );
  NOR2_X1 U785 ( .A1(n689), .A2(n688), .ZN(n691) );
  NAND2_X1 U786 ( .A1(G117), .A2(n899), .ZN(n690) );
  NAND2_X1 U787 ( .A1(n691), .A2(n690), .ZN(n882) );
  AND2_X1 U788 ( .A1(n882), .A2(G1996), .ZN(n972) );
  NAND2_X1 U789 ( .A1(n902), .A2(G95), .ZN(n693) );
  NAND2_X1 U790 ( .A1(G131), .A2(n608), .ZN(n692) );
  NAND2_X1 U791 ( .A1(n693), .A2(n692), .ZN(n697) );
  NAND2_X1 U792 ( .A1(G119), .A2(n898), .ZN(n695) );
  NAND2_X1 U793 ( .A1(G107), .A2(n899), .ZN(n694) );
  NAND2_X1 U794 ( .A1(n695), .A2(n694), .ZN(n696) );
  NOR2_X1 U795 ( .A1(n697), .A2(n696), .ZN(n897) );
  INV_X1 U796 ( .A(G1991), .ZN(n810) );
  NOR2_X1 U797 ( .A1(n897), .A2(n810), .ZN(n970) );
  OR2_X1 U798 ( .A1(n972), .A2(n970), .ZN(n698) );
  NAND2_X1 U799 ( .A1(n820), .A2(n698), .ZN(n809) );
  NAND2_X1 U800 ( .A1(n902), .A2(G104), .ZN(n700) );
  NAND2_X1 U801 ( .A1(G140), .A2(n608), .ZN(n699) );
  NAND2_X1 U802 ( .A1(n700), .A2(n699), .ZN(n701) );
  XNOR2_X1 U803 ( .A(KEYINPUT34), .B(n701), .ZN(n707) );
  NAND2_X1 U804 ( .A1(n898), .A2(G128), .ZN(n702) );
  XOR2_X1 U805 ( .A(KEYINPUT91), .B(n702), .Z(n704) );
  NAND2_X1 U806 ( .A1(G116), .A2(n899), .ZN(n703) );
  NAND2_X1 U807 ( .A1(n704), .A2(n703), .ZN(n705) );
  XOR2_X1 U808 ( .A(KEYINPUT35), .B(n705), .Z(n706) );
  NOR2_X1 U809 ( .A1(n707), .A2(n706), .ZN(n708) );
  XNOR2_X1 U810 ( .A(KEYINPUT36), .B(n708), .ZN(n914) );
  XNOR2_X1 U811 ( .A(G2067), .B(KEYINPUT37), .ZN(n808) );
  NOR2_X1 U812 ( .A1(n914), .A2(n808), .ZN(n991) );
  NAND2_X1 U813 ( .A1(n820), .A2(n991), .ZN(n816) );
  NAND2_X1 U814 ( .A1(n809), .A2(n816), .ZN(n709) );
  XNOR2_X1 U815 ( .A(n709), .B(KEYINPUT92), .ZN(n805) );
  AND2_X1 U816 ( .A1(G160), .A2(G40), .ZN(n711) );
  NAND2_X1 U817 ( .A1(n711), .A2(n710), .ZN(n757) );
  INV_X1 U818 ( .A(n757), .ZN(n726) );
  NAND2_X1 U819 ( .A1(n726), .A2(G1996), .ZN(n712) );
  XNOR2_X1 U820 ( .A(n712), .B(KEYINPUT26), .ZN(n714) );
  NAND2_X1 U821 ( .A1(n757), .A2(G1341), .ZN(n713) );
  NAND2_X1 U822 ( .A1(n714), .A2(n713), .ZN(n715) );
  XNOR2_X1 U823 ( .A(n717), .B(n716), .ZN(n723) );
  NOR2_X1 U824 ( .A1(n726), .A2(G1348), .ZN(n719) );
  NOR2_X1 U825 ( .A1(G2067), .A2(n757), .ZN(n718) );
  NOR2_X1 U826 ( .A1(n719), .A2(n718), .ZN(n720) );
  NAND2_X1 U827 ( .A1(n721), .A2(n720), .ZN(n725) );
  NAND2_X1 U828 ( .A1(n723), .A2(n722), .ZN(n724) );
  NAND2_X1 U829 ( .A1(n725), .A2(n724), .ZN(n732) );
  NAND2_X1 U830 ( .A1(G2072), .A2(n726), .ZN(n727) );
  XNOR2_X1 U831 ( .A(n727), .B(KEYINPUT94), .ZN(n728) );
  XNOR2_X1 U832 ( .A(KEYINPUT27), .B(n728), .ZN(n730) );
  INV_X1 U833 ( .A(G1956), .ZN(n999) );
  NOR2_X1 U834 ( .A1(n726), .A2(n999), .ZN(n729) );
  NOR2_X1 U835 ( .A1(n730), .A2(n729), .ZN(n734) );
  INV_X1 U836 ( .A(G299), .ZN(n733) );
  NAND2_X1 U837 ( .A1(n734), .A2(n733), .ZN(n731) );
  NAND2_X1 U838 ( .A1(n732), .A2(n731), .ZN(n737) );
  NOR2_X1 U839 ( .A1(n734), .A2(n733), .ZN(n735) );
  XOR2_X1 U840 ( .A(n735), .B(KEYINPUT28), .Z(n736) );
  NAND2_X1 U841 ( .A1(n737), .A2(n736), .ZN(n739) );
  XNOR2_X1 U842 ( .A(n739), .B(n738), .ZN(n744) );
  NAND2_X1 U843 ( .A1(G1961), .A2(n757), .ZN(n741) );
  XOR2_X1 U844 ( .A(KEYINPUT25), .B(G2078), .Z(n951) );
  NAND2_X1 U845 ( .A1(n726), .A2(n951), .ZN(n740) );
  NAND2_X1 U846 ( .A1(n741), .A2(n740), .ZN(n749) );
  NOR2_X1 U847 ( .A1(G301), .A2(n749), .ZN(n742) );
  XNOR2_X1 U848 ( .A(n742), .B(KEYINPUT93), .ZN(n743) );
  NAND2_X1 U849 ( .A1(n744), .A2(n743), .ZN(n756) );
  NAND2_X1 U850 ( .A1(G8), .A2(n757), .ZN(n797) );
  NOR2_X1 U851 ( .A1(G2084), .A2(n757), .ZN(n766) );
  NOR2_X1 U852 ( .A1(n769), .A2(n766), .ZN(n745) );
  XOR2_X1 U853 ( .A(KEYINPUT95), .B(n745), .Z(n746) );
  NAND2_X1 U854 ( .A1(G8), .A2(n746), .ZN(n747) );
  XNOR2_X1 U855 ( .A(KEYINPUT30), .B(n747), .ZN(n748) );
  NOR2_X1 U856 ( .A1(n748), .A2(G168), .ZN(n751) );
  AND2_X1 U857 ( .A1(G301), .A2(n749), .ZN(n750) );
  NOR2_X1 U858 ( .A1(n751), .A2(n750), .ZN(n754) );
  INV_X1 U859 ( .A(KEYINPUT31), .ZN(n752) );
  NAND2_X1 U860 ( .A1(n756), .A2(n755), .ZN(n767) );
  NAND2_X1 U861 ( .A1(n767), .A2(G286), .ZN(n764) );
  INV_X1 U862 ( .A(G8), .ZN(n762) );
  NOR2_X1 U863 ( .A1(G1971), .A2(n797), .ZN(n759) );
  NOR2_X1 U864 ( .A1(G2090), .A2(n757), .ZN(n758) );
  NOR2_X1 U865 ( .A1(n759), .A2(n758), .ZN(n760) );
  NAND2_X1 U866 ( .A1(n760), .A2(G303), .ZN(n761) );
  OR2_X1 U867 ( .A1(n762), .A2(n761), .ZN(n763) );
  XNOR2_X1 U868 ( .A(n765), .B(KEYINPUT32), .ZN(n773) );
  NAND2_X1 U869 ( .A1(G8), .A2(n766), .ZN(n771) );
  INV_X1 U870 ( .A(n767), .ZN(n768) );
  NOR2_X1 U871 ( .A1(n769), .A2(n768), .ZN(n770) );
  NAND2_X1 U872 ( .A1(n771), .A2(n770), .ZN(n772) );
  NAND2_X1 U873 ( .A1(n773), .A2(n772), .ZN(n795) );
  INV_X1 U874 ( .A(n795), .ZN(n776) );
  OR2_X1 U875 ( .A1(G303), .A2(G1971), .ZN(n775) );
  NOR2_X1 U876 ( .A1(G1976), .A2(G288), .ZN(n783) );
  INV_X1 U877 ( .A(n783), .ZN(n774) );
  NAND2_X1 U878 ( .A1(n775), .A2(n774), .ZN(n942) );
  NOR2_X1 U879 ( .A1(n776), .A2(n942), .ZN(n778) );
  NAND2_X1 U880 ( .A1(G1976), .A2(G288), .ZN(n936) );
  NOR2_X1 U881 ( .A1(KEYINPUT97), .A2(n779), .ZN(n780) );
  NOR2_X1 U882 ( .A1(KEYINPUT33), .A2(n780), .ZN(n790) );
  INV_X1 U883 ( .A(KEYINPUT97), .ZN(n782) );
  NAND2_X1 U884 ( .A1(n783), .A2(KEYINPUT33), .ZN(n781) );
  NAND2_X1 U885 ( .A1(n782), .A2(n781), .ZN(n785) );
  NAND2_X1 U886 ( .A1(n783), .A2(KEYINPUT97), .ZN(n784) );
  NAND2_X1 U887 ( .A1(n785), .A2(n784), .ZN(n786) );
  NOR2_X1 U888 ( .A1(n797), .A2(n786), .ZN(n788) );
  XOR2_X1 U889 ( .A(G1981), .B(G305), .Z(n925) );
  NOR2_X1 U890 ( .A1(G1981), .A2(G305), .ZN(n791) );
  XOR2_X1 U891 ( .A(n791), .B(KEYINPUT24), .Z(n792) );
  OR2_X1 U892 ( .A1(n797), .A2(n792), .ZN(n799) );
  NOR2_X1 U893 ( .A1(G2090), .A2(G303), .ZN(n793) );
  NAND2_X1 U894 ( .A1(G8), .A2(n793), .ZN(n794) );
  XNOR2_X1 U895 ( .A(n794), .B(KEYINPUT98), .ZN(n796) );
  NAND2_X1 U896 ( .A1(n796), .A2(n795), .ZN(n798) );
  NAND2_X1 U897 ( .A1(n799), .A2(n524), .ZN(n800) );
  NOR2_X1 U898 ( .A1(n801), .A2(n800), .ZN(n803) );
  XNOR2_X1 U899 ( .A(G1986), .B(G290), .ZN(n934) );
  NAND2_X1 U900 ( .A1(n934), .A2(n820), .ZN(n806) );
  NAND2_X1 U901 ( .A1(n807), .A2(n806), .ZN(n823) );
  NAND2_X1 U902 ( .A1(n914), .A2(n808), .ZN(n977) );
  NOR2_X1 U903 ( .A1(G1996), .A2(n882), .ZN(n980) );
  INV_X1 U904 ( .A(n809), .ZN(n813) );
  NOR2_X1 U905 ( .A1(G1986), .A2(G290), .ZN(n811) );
  AND2_X1 U906 ( .A1(n810), .A2(n897), .ZN(n971) );
  NOR2_X1 U907 ( .A1(n811), .A2(n971), .ZN(n812) );
  NOR2_X1 U908 ( .A1(n813), .A2(n812), .ZN(n814) );
  NOR2_X1 U909 ( .A1(n980), .A2(n814), .ZN(n815) );
  XNOR2_X1 U910 ( .A(n815), .B(KEYINPUT39), .ZN(n817) );
  NAND2_X1 U911 ( .A1(n817), .A2(n816), .ZN(n818) );
  NAND2_X1 U912 ( .A1(n977), .A2(n818), .ZN(n819) );
  XNOR2_X1 U913 ( .A(KEYINPUT100), .B(n819), .ZN(n821) );
  NAND2_X1 U914 ( .A1(n821), .A2(n820), .ZN(n822) );
  NAND2_X1 U915 ( .A1(n823), .A2(n822), .ZN(n824) );
  XNOR2_X1 U916 ( .A(n824), .B(KEYINPUT40), .ZN(G329) );
  INV_X1 U917 ( .A(G301), .ZN(G171) );
  XNOR2_X1 U918 ( .A(G2443), .B(G2451), .ZN(n834) );
  XOR2_X1 U919 ( .A(G2446), .B(KEYINPUT101), .Z(n826) );
  XNOR2_X1 U920 ( .A(KEYINPUT102), .B(G2438), .ZN(n825) );
  XNOR2_X1 U921 ( .A(n826), .B(n825), .ZN(n830) );
  XOR2_X1 U922 ( .A(G2435), .B(G2454), .Z(n828) );
  XNOR2_X1 U923 ( .A(G1348), .B(G1341), .ZN(n827) );
  XNOR2_X1 U924 ( .A(n828), .B(n827), .ZN(n829) );
  XOR2_X1 U925 ( .A(n830), .B(n829), .Z(n832) );
  XNOR2_X1 U926 ( .A(G2427), .B(G2430), .ZN(n831) );
  XNOR2_X1 U927 ( .A(n832), .B(n831), .ZN(n833) );
  XNOR2_X1 U928 ( .A(n834), .B(n833), .ZN(n835) );
  NAND2_X1 U929 ( .A1(n835), .A2(G14), .ZN(n917) );
  XNOR2_X1 U930 ( .A(KEYINPUT103), .B(n917), .ZN(G401) );
  NAND2_X1 U931 ( .A1(G2106), .A2(n836), .ZN(G217) );
  AND2_X1 U932 ( .A1(G15), .A2(G2), .ZN(n837) );
  NAND2_X1 U933 ( .A1(G661), .A2(n837), .ZN(G259) );
  NAND2_X1 U934 ( .A1(G3), .A2(G1), .ZN(n838) );
  NAND2_X1 U935 ( .A1(n839), .A2(n838), .ZN(G188) );
  XNOR2_X1 U936 ( .A(G108), .B(KEYINPUT115), .ZN(G238) );
  NAND2_X1 U938 ( .A1(n841), .A2(n840), .ZN(n843) );
  XNOR2_X1 U939 ( .A(n843), .B(n842), .ZN(G145) );
  INV_X1 U940 ( .A(G132), .ZN(G219) );
  INV_X1 U941 ( .A(G120), .ZN(G236) );
  INV_X1 U942 ( .A(G96), .ZN(G221) );
  INV_X1 U943 ( .A(G82), .ZN(G220) );
  NOR2_X1 U944 ( .A1(n845), .A2(n844), .ZN(G325) );
  INV_X1 U945 ( .A(G325), .ZN(G261) );
  XOR2_X1 U946 ( .A(n846), .B(G286), .Z(n848) );
  XNOR2_X1 U947 ( .A(G171), .B(n924), .ZN(n847) );
  XNOR2_X1 U948 ( .A(n848), .B(n847), .ZN(n849) );
  XNOR2_X1 U949 ( .A(n849), .B(n930), .ZN(n850) );
  NOR2_X1 U950 ( .A1(G37), .A2(n850), .ZN(G397) );
  INV_X1 U951 ( .A(n851), .ZN(G319) );
  XOR2_X1 U952 ( .A(G2096), .B(KEYINPUT104), .Z(n853) );
  XNOR2_X1 U953 ( .A(G2090), .B(KEYINPUT43), .ZN(n852) );
  XNOR2_X1 U954 ( .A(n853), .B(n852), .ZN(n854) );
  XOR2_X1 U955 ( .A(n854), .B(KEYINPUT42), .Z(n856) );
  XNOR2_X1 U956 ( .A(G2067), .B(G2072), .ZN(n855) );
  XNOR2_X1 U957 ( .A(n856), .B(n855), .ZN(n860) );
  XOR2_X1 U958 ( .A(G2678), .B(G2100), .Z(n858) );
  XNOR2_X1 U959 ( .A(G2084), .B(G2078), .ZN(n857) );
  XNOR2_X1 U960 ( .A(n858), .B(n857), .ZN(n859) );
  XNOR2_X1 U961 ( .A(n860), .B(n859), .ZN(G227) );
  XOR2_X1 U962 ( .A(KEYINPUT106), .B(G1961), .Z(n862) );
  XNOR2_X1 U963 ( .A(G1996), .B(G1991), .ZN(n861) );
  XNOR2_X1 U964 ( .A(n862), .B(n861), .ZN(n863) );
  XOR2_X1 U965 ( .A(n863), .B(KEYINPUT41), .Z(n865) );
  XNOR2_X1 U966 ( .A(G1986), .B(G1956), .ZN(n864) );
  XNOR2_X1 U967 ( .A(n865), .B(n864), .ZN(n869) );
  XOR2_X1 U968 ( .A(G1976), .B(G1981), .Z(n867) );
  XNOR2_X1 U969 ( .A(G1966), .B(G1971), .ZN(n866) );
  XNOR2_X1 U970 ( .A(n867), .B(n866), .ZN(n868) );
  XOR2_X1 U971 ( .A(n869), .B(n868), .Z(n871) );
  XNOR2_X1 U972 ( .A(G2474), .B(KEYINPUT105), .ZN(n870) );
  XNOR2_X1 U973 ( .A(n871), .B(n870), .ZN(G229) );
  NAND2_X1 U974 ( .A1(G100), .A2(n902), .ZN(n873) );
  NAND2_X1 U975 ( .A1(G112), .A2(n899), .ZN(n872) );
  NAND2_X1 U976 ( .A1(n873), .A2(n872), .ZN(n881) );
  NAND2_X1 U977 ( .A1(G136), .A2(n608), .ZN(n874) );
  XNOR2_X1 U978 ( .A(KEYINPUT108), .B(n874), .ZN(n878) );
  XOR2_X1 U979 ( .A(KEYINPUT44), .B(KEYINPUT107), .Z(n876) );
  NAND2_X1 U980 ( .A1(G124), .A2(n898), .ZN(n875) );
  XNOR2_X1 U981 ( .A(n876), .B(n875), .ZN(n877) );
  NAND2_X1 U982 ( .A1(n878), .A2(n877), .ZN(n879) );
  XOR2_X1 U983 ( .A(KEYINPUT109), .B(n879), .Z(n880) );
  NOR2_X1 U984 ( .A1(n881), .A2(n880), .ZN(G162) );
  XOR2_X1 U985 ( .A(G160), .B(n882), .Z(n891) );
  NAND2_X1 U986 ( .A1(n902), .A2(G103), .ZN(n884) );
  NAND2_X1 U987 ( .A1(G139), .A2(n608), .ZN(n883) );
  NAND2_X1 U988 ( .A1(n884), .A2(n883), .ZN(n890) );
  NAND2_X1 U989 ( .A1(G127), .A2(n898), .ZN(n886) );
  NAND2_X1 U990 ( .A1(G115), .A2(n899), .ZN(n885) );
  NAND2_X1 U991 ( .A1(n886), .A2(n885), .ZN(n887) );
  XNOR2_X1 U992 ( .A(KEYINPUT47), .B(n887), .ZN(n888) );
  XNOR2_X1 U993 ( .A(KEYINPUT111), .B(n888), .ZN(n889) );
  NOR2_X1 U994 ( .A1(n890), .A2(n889), .ZN(n984) );
  XNOR2_X1 U995 ( .A(n891), .B(n984), .ZN(n896) );
  XOR2_X1 U996 ( .A(KEYINPUT112), .B(KEYINPUT113), .Z(n893) );
  XNOR2_X1 U997 ( .A(KEYINPUT46), .B(KEYINPUT48), .ZN(n892) );
  XNOR2_X1 U998 ( .A(n893), .B(n892), .ZN(n894) );
  XOR2_X1 U999 ( .A(G164), .B(n894), .Z(n895) );
  XOR2_X1 U1000 ( .A(n896), .B(n895), .Z(n913) );
  XNOR2_X1 U1001 ( .A(n897), .B(n969), .ZN(n910) );
  NAND2_X1 U1002 ( .A1(G130), .A2(n898), .ZN(n901) );
  NAND2_X1 U1003 ( .A1(G118), .A2(n899), .ZN(n900) );
  NAND2_X1 U1004 ( .A1(n901), .A2(n900), .ZN(n908) );
  NAND2_X1 U1005 ( .A1(n902), .A2(G106), .ZN(n904) );
  NAND2_X1 U1006 ( .A1(G142), .A2(n608), .ZN(n903) );
  NAND2_X1 U1007 ( .A1(n904), .A2(n903), .ZN(n905) );
  XOR2_X1 U1008 ( .A(KEYINPUT110), .B(n905), .Z(n906) );
  XNOR2_X1 U1009 ( .A(KEYINPUT45), .B(n906), .ZN(n907) );
  NOR2_X1 U1010 ( .A1(n908), .A2(n907), .ZN(n909) );
  XNOR2_X1 U1011 ( .A(n910), .B(n909), .ZN(n911) );
  XNOR2_X1 U1012 ( .A(G162), .B(n911), .ZN(n912) );
  XNOR2_X1 U1013 ( .A(n913), .B(n912), .ZN(n915) );
  XNOR2_X1 U1014 ( .A(n915), .B(n914), .ZN(n916) );
  NOR2_X1 U1015 ( .A1(G37), .A2(n916), .ZN(G395) );
  NAND2_X1 U1016 ( .A1(G319), .A2(n917), .ZN(n918) );
  NOR2_X1 U1017 ( .A1(G397), .A2(n918), .ZN(n921) );
  NOR2_X1 U1018 ( .A1(G227), .A2(G229), .ZN(n919) );
  XOR2_X1 U1019 ( .A(KEYINPUT49), .B(n919), .Z(n920) );
  NAND2_X1 U1020 ( .A1(n921), .A2(n920), .ZN(n922) );
  NOR2_X1 U1021 ( .A1(n922), .A2(G395), .ZN(n923) );
  XNOR2_X1 U1022 ( .A(n923), .B(KEYINPUT114), .ZN(G308) );
  INV_X1 U1023 ( .A(G308), .ZN(G225) );
  INV_X1 U1024 ( .A(G69), .ZN(G235) );
  XNOR2_X1 U1025 ( .A(KEYINPUT62), .B(KEYINPUT127), .ZN(n1032) );
  XNOR2_X1 U1026 ( .A(KEYINPUT56), .B(G16), .ZN(n946) );
  XNOR2_X1 U1027 ( .A(G1348), .B(n924), .ZN(n929) );
  XNOR2_X1 U1028 ( .A(G1966), .B(G168), .ZN(n926) );
  NAND2_X1 U1029 ( .A1(n926), .A2(n925), .ZN(n927) );
  XNOR2_X1 U1030 ( .A(n927), .B(KEYINPUT57), .ZN(n928) );
  NAND2_X1 U1031 ( .A1(n929), .A2(n928), .ZN(n932) );
  XNOR2_X1 U1032 ( .A(G1341), .B(n930), .ZN(n931) );
  NOR2_X1 U1033 ( .A1(n932), .A2(n931), .ZN(n944) );
  XNOR2_X1 U1034 ( .A(G1961), .B(G301), .ZN(n933) );
  NOR2_X1 U1035 ( .A1(n934), .A2(n933), .ZN(n940) );
  NAND2_X1 U1036 ( .A1(G1971), .A2(G303), .ZN(n935) );
  NAND2_X1 U1037 ( .A1(n936), .A2(n935), .ZN(n938) );
  XNOR2_X1 U1038 ( .A(G1956), .B(G299), .ZN(n937) );
  NOR2_X1 U1039 ( .A1(n938), .A2(n937), .ZN(n939) );
  NAND2_X1 U1040 ( .A1(n940), .A2(n939), .ZN(n941) );
  NOR2_X1 U1041 ( .A1(n942), .A2(n941), .ZN(n943) );
  NAND2_X1 U1042 ( .A1(n944), .A2(n943), .ZN(n945) );
  NAND2_X1 U1043 ( .A1(n946), .A2(n945), .ZN(n947) );
  XNOR2_X1 U1044 ( .A(KEYINPUT122), .B(n947), .ZN(n1030) );
  XOR2_X1 U1045 ( .A(G2067), .B(G26), .Z(n948) );
  NAND2_X1 U1046 ( .A1(n948), .A2(G28), .ZN(n957) );
  XNOR2_X1 U1047 ( .A(G1996), .B(G32), .ZN(n950) );
  XNOR2_X1 U1048 ( .A(G33), .B(G2072), .ZN(n949) );
  NOR2_X1 U1049 ( .A1(n950), .A2(n949), .ZN(n955) );
  XNOR2_X1 U1050 ( .A(G1991), .B(G25), .ZN(n953) );
  XNOR2_X1 U1051 ( .A(G27), .B(n951), .ZN(n952) );
  NOR2_X1 U1052 ( .A1(n953), .A2(n952), .ZN(n954) );
  NAND2_X1 U1053 ( .A1(n955), .A2(n954), .ZN(n956) );
  NOR2_X1 U1054 ( .A1(n957), .A2(n956), .ZN(n958) );
  XOR2_X1 U1055 ( .A(KEYINPUT53), .B(n958), .Z(n961) );
  XOR2_X1 U1056 ( .A(G34), .B(KEYINPUT54), .Z(n959) );
  XNOR2_X1 U1057 ( .A(G2084), .B(n959), .ZN(n960) );
  NAND2_X1 U1058 ( .A1(n961), .A2(n960), .ZN(n964) );
  XNOR2_X1 U1059 ( .A(KEYINPUT120), .B(G2090), .ZN(n962) );
  XNOR2_X1 U1060 ( .A(G35), .B(n962), .ZN(n963) );
  NOR2_X1 U1061 ( .A1(n964), .A2(n963), .ZN(n965) );
  XNOR2_X1 U1062 ( .A(KEYINPUT55), .B(KEYINPUT119), .ZN(n996) );
  XOR2_X1 U1063 ( .A(n965), .B(n996), .Z(n967) );
  XNOR2_X1 U1064 ( .A(G29), .B(KEYINPUT121), .ZN(n966) );
  NAND2_X1 U1065 ( .A1(n967), .A2(n966), .ZN(n968) );
  NAND2_X1 U1066 ( .A1(G11), .A2(n968), .ZN(n1028) );
  NOR2_X1 U1067 ( .A1(n970), .A2(n969), .ZN(n974) );
  NOR2_X1 U1068 ( .A1(n972), .A2(n971), .ZN(n973) );
  NAND2_X1 U1069 ( .A1(n974), .A2(n973), .ZN(n976) );
  XOR2_X1 U1070 ( .A(G160), .B(G2084), .Z(n975) );
  NOR2_X1 U1071 ( .A1(n976), .A2(n975), .ZN(n978) );
  NAND2_X1 U1072 ( .A1(n978), .A2(n977), .ZN(n983) );
  XOR2_X1 U1073 ( .A(G2090), .B(G162), .Z(n979) );
  NOR2_X1 U1074 ( .A1(n980), .A2(n979), .ZN(n981) );
  XNOR2_X1 U1075 ( .A(n981), .B(KEYINPUT51), .ZN(n982) );
  NOR2_X1 U1076 ( .A1(n983), .A2(n982), .ZN(n993) );
  XNOR2_X1 U1077 ( .A(n984), .B(G2072), .ZN(n985) );
  XNOR2_X1 U1078 ( .A(n985), .B(KEYINPUT116), .ZN(n988) );
  XOR2_X1 U1079 ( .A(G164), .B(G2078), .Z(n986) );
  XNOR2_X1 U1080 ( .A(KEYINPUT117), .B(n986), .ZN(n987) );
  NAND2_X1 U1081 ( .A1(n988), .A2(n987), .ZN(n989) );
  XNOR2_X1 U1082 ( .A(KEYINPUT50), .B(n989), .ZN(n990) );
  NOR2_X1 U1083 ( .A1(n991), .A2(n990), .ZN(n992) );
  NAND2_X1 U1084 ( .A1(n993), .A2(n992), .ZN(n994) );
  XNOR2_X1 U1085 ( .A(KEYINPUT52), .B(n994), .ZN(n995) );
  XOR2_X1 U1086 ( .A(KEYINPUT118), .B(n995), .Z(n997) );
  NAND2_X1 U1087 ( .A1(n997), .A2(n996), .ZN(n998) );
  NAND2_X1 U1088 ( .A1(n998), .A2(G29), .ZN(n1026) );
  XNOR2_X1 U1089 ( .A(G20), .B(n999), .ZN(n1003) );
  XNOR2_X1 U1090 ( .A(G1341), .B(G19), .ZN(n1001) );
  XNOR2_X1 U1091 ( .A(G1981), .B(G6), .ZN(n1000) );
  NOR2_X1 U1092 ( .A1(n1001), .A2(n1000), .ZN(n1002) );
  NAND2_X1 U1093 ( .A1(n1003), .A2(n1002), .ZN(n1006) );
  XOR2_X1 U1094 ( .A(KEYINPUT59), .B(G1348), .Z(n1004) );
  XNOR2_X1 U1095 ( .A(G4), .B(n1004), .ZN(n1005) );
  NOR2_X1 U1096 ( .A1(n1006), .A2(n1005), .ZN(n1007) );
  XNOR2_X1 U1097 ( .A(KEYINPUT124), .B(n1007), .ZN(n1008) );
  XNOR2_X1 U1098 ( .A(n1008), .B(KEYINPUT60), .ZN(n1019) );
  XOR2_X1 U1099 ( .A(G1961), .B(KEYINPUT123), .Z(n1009) );
  XNOR2_X1 U1100 ( .A(G5), .B(n1009), .ZN(n1017) );
  XNOR2_X1 U1101 ( .A(G1986), .B(G24), .ZN(n1011) );
  XNOR2_X1 U1102 ( .A(G23), .B(G1976), .ZN(n1010) );
  NOR2_X1 U1103 ( .A1(n1011), .A2(n1010), .ZN(n1014) );
  XNOR2_X1 U1104 ( .A(G1971), .B(G22), .ZN(n1012) );
  XNOR2_X1 U1105 ( .A(n1012), .B(KEYINPUT125), .ZN(n1013) );
  NAND2_X1 U1106 ( .A1(n1014), .A2(n1013), .ZN(n1015) );
  XNOR2_X1 U1107 ( .A(KEYINPUT58), .B(n1015), .ZN(n1016) );
  NOR2_X1 U1108 ( .A1(n1017), .A2(n1016), .ZN(n1018) );
  NAND2_X1 U1109 ( .A1(n1019), .A2(n1018), .ZN(n1021) );
  XNOR2_X1 U1110 ( .A(G21), .B(G1966), .ZN(n1020) );
  NOR2_X1 U1111 ( .A1(n1021), .A2(n1020), .ZN(n1022) );
  XOR2_X1 U1112 ( .A(KEYINPUT61), .B(n1022), .Z(n1023) );
  NOR2_X1 U1113 ( .A1(G16), .A2(n1023), .ZN(n1024) );
  XOR2_X1 U1114 ( .A(KEYINPUT126), .B(n1024), .Z(n1025) );
  NAND2_X1 U1115 ( .A1(n1026), .A2(n1025), .ZN(n1027) );
  NOR2_X1 U1116 ( .A1(n1028), .A2(n1027), .ZN(n1029) );
  NAND2_X1 U1117 ( .A1(n1030), .A2(n1029), .ZN(n1031) );
  XNOR2_X1 U1118 ( .A(n1032), .B(n1031), .ZN(G311) );
  INV_X1 U1119 ( .A(G311), .ZN(G150) );
endmodule

