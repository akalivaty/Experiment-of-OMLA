//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 1 0 0 0 1 1 1 1 0 1 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 0 1 0 0 0 1 0 0 1 1 0 0 1 0 1 0 0 1 0 0 1 1 1 0 1 1 0 1 0 0 0 0 1 0 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:26:37 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n633, new_n634, new_n635, new_n636,
    new_n638, new_n639, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n681, new_n682,
    new_n683, new_n684, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n695, new_n697, new_n698, new_n699,
    new_n701, new_n702, new_n703, new_n704, new_n705, new_n706, new_n708,
    new_n709, new_n710, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n721, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n744, new_n745, new_n746, new_n747,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n884,
    new_n885, new_n886, new_n888, new_n889, new_n890, new_n891, new_n892,
    new_n893, new_n894, new_n895, new_n896, new_n897, new_n898, new_n899,
    new_n900, new_n901, new_n902, new_n903, new_n904, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n949, new_n950, new_n951, new_n952,
    new_n953, new_n954, new_n955, new_n956, new_n957, new_n958, new_n959,
    new_n960;
  XNOR2_X1  g000(.A(G113), .B(G122), .ZN(new_n187));
  XNOR2_X1  g001(.A(KEYINPUT92), .B(G104), .ZN(new_n188));
  XNOR2_X1  g002(.A(new_n187), .B(new_n188), .ZN(new_n189));
  INV_X1    g003(.A(new_n189), .ZN(new_n190));
  INV_X1    g004(.A(G237), .ZN(new_n191));
  INV_X1    g005(.A(G953), .ZN(new_n192));
  NAND3_X1  g006(.A1(new_n191), .A2(new_n192), .A3(G214), .ZN(new_n193));
  XNOR2_X1  g007(.A(new_n193), .B(G143), .ZN(new_n194));
  INV_X1    g008(.A(G131), .ZN(new_n195));
  NOR2_X1   g009(.A1(new_n194), .A2(new_n195), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n196), .A2(KEYINPUT18), .ZN(new_n197));
  INV_X1    g011(.A(KEYINPUT18), .ZN(new_n198));
  OAI21_X1  g012(.A(new_n194), .B1(new_n198), .B2(new_n195), .ZN(new_n199));
  XNOR2_X1  g013(.A(G125), .B(G140), .ZN(new_n200));
  INV_X1    g014(.A(G146), .ZN(new_n201));
  XNOR2_X1  g015(.A(new_n200), .B(new_n201), .ZN(new_n202));
  NAND3_X1  g016(.A1(new_n197), .A2(new_n199), .A3(new_n202), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n196), .A2(KEYINPUT17), .ZN(new_n204));
  XNOR2_X1  g018(.A(new_n194), .B(new_n195), .ZN(new_n205));
  OAI21_X1  g019(.A(new_n204), .B1(new_n205), .B2(KEYINPUT17), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n200), .A2(KEYINPUT16), .ZN(new_n207));
  INV_X1    g021(.A(G125), .ZN(new_n208));
  OR3_X1    g022(.A1(new_n208), .A2(KEYINPUT16), .A3(G140), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n207), .A2(new_n209), .ZN(new_n210));
  AOI21_X1  g024(.A(KEYINPUT75), .B1(new_n210), .B2(new_n201), .ZN(new_n211));
  NOR2_X1   g025(.A1(new_n210), .A2(new_n201), .ZN(new_n212));
  NOR2_X1   g026(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  NAND3_X1  g027(.A1(new_n210), .A2(KEYINPUT75), .A3(new_n201), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n213), .A2(new_n214), .ZN(new_n215));
  OAI211_X1 g029(.A(new_n190), .B(new_n203), .C1(new_n206), .C2(new_n215), .ZN(new_n216));
  INV_X1    g030(.A(KEYINPUT93), .ZN(new_n217));
  OR2_X1    g031(.A1(new_n216), .A2(new_n217), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n216), .A2(new_n217), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n218), .A2(new_n219), .ZN(new_n220));
  XNOR2_X1  g034(.A(new_n200), .B(KEYINPUT19), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n221), .A2(new_n201), .ZN(new_n222));
  OAI21_X1  g036(.A(new_n222), .B1(new_n201), .B2(new_n210), .ZN(new_n223));
  INV_X1    g037(.A(KEYINPUT91), .ZN(new_n224));
  OR2_X1    g038(.A1(new_n223), .A2(new_n224), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n223), .A2(new_n224), .ZN(new_n226));
  NAND3_X1  g040(.A1(new_n225), .A2(new_n226), .A3(new_n205), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n227), .A2(new_n203), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n228), .A2(new_n189), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n220), .A2(new_n229), .ZN(new_n230));
  INV_X1    g044(.A(KEYINPUT20), .ZN(new_n231));
  NOR2_X1   g045(.A1(G475), .A2(G902), .ZN(new_n232));
  NAND3_X1  g046(.A1(new_n230), .A2(new_n231), .A3(new_n232), .ZN(new_n233));
  AOI22_X1  g047(.A1(new_n218), .A2(new_n219), .B1(new_n189), .B2(new_n228), .ZN(new_n234));
  INV_X1    g048(.A(new_n232), .ZN(new_n235));
  OAI21_X1  g049(.A(KEYINPUT20), .B1(new_n234), .B2(new_n235), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n233), .A2(new_n236), .ZN(new_n237));
  OR2_X1    g051(.A1(new_n206), .A2(new_n215), .ZN(new_n238));
  AOI21_X1  g052(.A(new_n190), .B1(new_n238), .B2(new_n203), .ZN(new_n239));
  AOI21_X1  g053(.A(new_n239), .B1(new_n218), .B2(new_n219), .ZN(new_n240));
  OAI21_X1  g054(.A(G475), .B1(new_n240), .B2(G902), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n237), .A2(new_n241), .ZN(new_n242));
  INV_X1    g056(.A(new_n242), .ZN(new_n243));
  INV_X1    g057(.A(KEYINPUT97), .ZN(new_n244));
  NAND2_X1  g058(.A1(G234), .A2(G237), .ZN(new_n245));
  AND3_X1   g059(.A1(new_n245), .A2(G952), .A3(new_n192), .ZN(new_n246));
  NAND3_X1  g060(.A1(new_n245), .A2(G902), .A3(G953), .ZN(new_n247));
  XOR2_X1   g061(.A(new_n247), .B(KEYINPUT96), .Z(new_n248));
  XNOR2_X1  g062(.A(KEYINPUT21), .B(G898), .ZN(new_n249));
  AOI21_X1  g063(.A(new_n246), .B1(new_n248), .B2(new_n249), .ZN(new_n250));
  INV_X1    g064(.A(new_n250), .ZN(new_n251));
  INV_X1    g065(.A(G116), .ZN(new_n252));
  AND2_X1   g066(.A1(new_n252), .A2(G122), .ZN(new_n253));
  INV_X1    g067(.A(KEYINPUT14), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n253), .A2(new_n254), .ZN(new_n255));
  NOR2_X1   g069(.A1(new_n252), .A2(G122), .ZN(new_n256));
  NOR2_X1   g070(.A1(new_n256), .A2(KEYINPUT14), .ZN(new_n257));
  OAI21_X1  g071(.A(new_n255), .B1(new_n257), .B2(new_n253), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n258), .A2(G107), .ZN(new_n259));
  INV_X1    g073(.A(KEYINPUT95), .ZN(new_n260));
  XNOR2_X1  g074(.A(new_n259), .B(new_n260), .ZN(new_n261));
  NOR2_X1   g075(.A1(new_n253), .A2(new_n256), .ZN(new_n262));
  INV_X1    g076(.A(G107), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n262), .A2(new_n263), .ZN(new_n264));
  INV_X1    g078(.A(G143), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n265), .A2(G128), .ZN(new_n266));
  INV_X1    g080(.A(G128), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n267), .A2(G143), .ZN(new_n268));
  INV_X1    g082(.A(G134), .ZN(new_n269));
  NAND3_X1  g083(.A1(new_n266), .A2(new_n268), .A3(new_n269), .ZN(new_n270));
  INV_X1    g084(.A(new_n270), .ZN(new_n271));
  AOI21_X1  g085(.A(new_n269), .B1(new_n266), .B2(new_n268), .ZN(new_n272));
  OAI211_X1 g086(.A(new_n261), .B(new_n264), .C1(new_n271), .C2(new_n272), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n268), .A2(KEYINPUT13), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n274), .A2(new_n266), .ZN(new_n275));
  NAND3_X1  g089(.A1(new_n265), .A2(KEYINPUT13), .A3(G128), .ZN(new_n276));
  AOI21_X1  g090(.A(new_n269), .B1(new_n275), .B2(new_n276), .ZN(new_n277));
  INV_X1    g091(.A(KEYINPUT94), .ZN(new_n278));
  OR2_X1    g092(.A1(new_n277), .A2(new_n278), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n277), .A2(new_n278), .ZN(new_n280));
  XNOR2_X1  g094(.A(new_n262), .B(new_n263), .ZN(new_n281));
  NAND4_X1  g095(.A1(new_n279), .A2(new_n270), .A3(new_n280), .A4(new_n281), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n273), .A2(new_n282), .ZN(new_n283));
  XNOR2_X1  g097(.A(KEYINPUT9), .B(G234), .ZN(new_n284));
  INV_X1    g098(.A(G217), .ZN(new_n285));
  NOR3_X1   g099(.A1(new_n284), .A2(new_n285), .A3(G953), .ZN(new_n286));
  INV_X1    g100(.A(new_n286), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n283), .A2(new_n287), .ZN(new_n288));
  NAND3_X1  g102(.A1(new_n273), .A2(new_n282), .A3(new_n286), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n288), .A2(new_n289), .ZN(new_n290));
  INV_X1    g104(.A(G902), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n290), .A2(new_n291), .ZN(new_n292));
  INV_X1    g106(.A(G478), .ZN(new_n293));
  NOR2_X1   g107(.A1(new_n293), .A2(KEYINPUT15), .ZN(new_n294));
  AND2_X1   g108(.A1(new_n292), .A2(new_n294), .ZN(new_n295));
  NOR2_X1   g109(.A1(new_n292), .A2(new_n294), .ZN(new_n296));
  NOR2_X1   g110(.A1(new_n295), .A2(new_n296), .ZN(new_n297));
  NAND4_X1  g111(.A1(new_n243), .A2(new_n244), .A3(new_n251), .A4(new_n297), .ZN(new_n298));
  NAND3_X1  g112(.A1(new_n297), .A2(new_n237), .A3(new_n241), .ZN(new_n299));
  OAI21_X1  g113(.A(KEYINPUT97), .B1(new_n299), .B2(new_n250), .ZN(new_n300));
  NAND2_X1  g114(.A1(new_n298), .A2(new_n300), .ZN(new_n301));
  OAI21_X1  g115(.A(G221), .B1(new_n284), .B2(G902), .ZN(new_n302));
  INV_X1    g116(.A(G469), .ZN(new_n303));
  INV_X1    g117(.A(KEYINPUT67), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n201), .A2(G143), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n265), .A2(G146), .ZN(new_n306));
  AOI21_X1  g120(.A(G128), .B1(new_n305), .B2(new_n306), .ZN(new_n307));
  NAND3_X1  g121(.A1(new_n265), .A2(KEYINPUT1), .A3(G146), .ZN(new_n308));
  INV_X1    g122(.A(new_n308), .ZN(new_n309));
  OAI21_X1  g123(.A(new_n304), .B1(new_n307), .B2(new_n309), .ZN(new_n310));
  XNOR2_X1  g124(.A(G143), .B(G146), .ZN(new_n311));
  OAI211_X1 g125(.A(KEYINPUT67), .B(new_n308), .C1(new_n311), .C2(G128), .ZN(new_n312));
  INV_X1    g126(.A(KEYINPUT1), .ZN(new_n313));
  NAND3_X1  g127(.A1(new_n311), .A2(new_n313), .A3(G128), .ZN(new_n314));
  NAND3_X1  g128(.A1(new_n310), .A2(new_n312), .A3(new_n314), .ZN(new_n315));
  AND2_X1   g129(.A1(KEYINPUT79), .A2(G104), .ZN(new_n316));
  NOR2_X1   g130(.A1(KEYINPUT79), .A2(G104), .ZN(new_n317));
  OAI21_X1  g131(.A(new_n263), .B1(new_n316), .B2(new_n317), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n318), .A2(KEYINPUT3), .ZN(new_n319));
  INV_X1    g133(.A(KEYINPUT3), .ZN(new_n320));
  NAND3_X1  g134(.A1(new_n320), .A2(new_n263), .A3(G104), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n321), .A2(KEYINPUT80), .ZN(new_n322));
  INV_X1    g136(.A(KEYINPUT80), .ZN(new_n323));
  NAND4_X1  g137(.A1(new_n323), .A2(new_n320), .A3(new_n263), .A4(G104), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n322), .A2(new_n324), .ZN(new_n325));
  INV_X1    g139(.A(G101), .ZN(new_n326));
  NOR2_X1   g140(.A1(new_n316), .A2(new_n317), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n327), .A2(G107), .ZN(new_n328));
  NAND4_X1  g142(.A1(new_n319), .A2(new_n325), .A3(new_n326), .A4(new_n328), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n329), .A2(KEYINPUT81), .ZN(new_n330));
  AOI22_X1  g144(.A1(new_n322), .A2(new_n324), .B1(new_n327), .B2(G107), .ZN(new_n331));
  INV_X1    g145(.A(KEYINPUT81), .ZN(new_n332));
  NAND4_X1  g146(.A1(new_n331), .A2(new_n332), .A3(new_n326), .A4(new_n319), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n330), .A2(new_n333), .ZN(new_n334));
  OR2_X1    g148(.A1(new_n263), .A2(G104), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n318), .A2(new_n335), .ZN(new_n336));
  INV_X1    g150(.A(new_n336), .ZN(new_n337));
  OAI21_X1  g151(.A(KEYINPUT82), .B1(new_n337), .B2(new_n326), .ZN(new_n338));
  INV_X1    g152(.A(KEYINPUT82), .ZN(new_n339));
  NAND3_X1  g153(.A1(new_n336), .A2(new_n339), .A3(G101), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n338), .A2(new_n340), .ZN(new_n341));
  AND3_X1   g155(.A1(new_n334), .A2(KEYINPUT83), .A3(new_n341), .ZN(new_n342));
  AOI21_X1  g156(.A(KEYINPUT83), .B1(new_n334), .B2(new_n341), .ZN(new_n343));
  OAI211_X1 g157(.A(KEYINPUT10), .B(new_n315), .C1(new_n342), .C2(new_n343), .ZN(new_n344));
  NAND2_X1  g158(.A1(KEYINPUT65), .A2(G131), .ZN(new_n345));
  INV_X1    g159(.A(new_n345), .ZN(new_n346));
  INV_X1    g160(.A(KEYINPUT11), .ZN(new_n347));
  OAI211_X1 g161(.A(KEYINPUT64), .B(new_n347), .C1(new_n269), .C2(G137), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n269), .A2(G137), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n348), .A2(new_n349), .ZN(new_n350));
  INV_X1    g164(.A(G137), .ZN(new_n351));
  NAND2_X1  g165(.A1(new_n351), .A2(G134), .ZN(new_n352));
  AOI21_X1  g166(.A(new_n347), .B1(new_n352), .B2(KEYINPUT64), .ZN(new_n353));
  OAI21_X1  g167(.A(new_n346), .B1(new_n350), .B2(new_n353), .ZN(new_n354));
  OAI21_X1  g168(.A(KEYINPUT64), .B1(new_n269), .B2(G137), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n355), .A2(KEYINPUT11), .ZN(new_n356));
  NAND4_X1  g170(.A1(new_n356), .A2(new_n348), .A3(new_n349), .A4(new_n345), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n354), .A2(new_n357), .ZN(new_n358));
  INV_X1    g172(.A(new_n358), .ZN(new_n359));
  NOR2_X1   g173(.A1(new_n307), .A2(new_n309), .ZN(new_n360));
  NAND2_X1  g174(.A1(new_n360), .A2(new_n314), .ZN(new_n361));
  NAND3_X1  g175(.A1(new_n334), .A2(new_n341), .A3(new_n361), .ZN(new_n362));
  INV_X1    g176(.A(KEYINPUT10), .ZN(new_n363));
  AOI21_X1  g177(.A(new_n326), .B1(new_n331), .B2(new_n319), .ZN(new_n364));
  INV_X1    g178(.A(KEYINPUT4), .ZN(new_n365));
  NOR2_X1   g179(.A1(new_n364), .A2(new_n365), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n334), .A2(new_n366), .ZN(new_n367));
  INV_X1    g181(.A(KEYINPUT0), .ZN(new_n368));
  OAI21_X1  g182(.A(new_n311), .B1(new_n368), .B2(new_n267), .ZN(new_n369));
  XOR2_X1   g183(.A(KEYINPUT0), .B(G128), .Z(new_n370));
  OAI21_X1  g184(.A(new_n369), .B1(new_n311), .B2(new_n370), .ZN(new_n371));
  INV_X1    g185(.A(new_n371), .ZN(new_n372));
  AOI21_X1  g186(.A(new_n372), .B1(new_n364), .B2(new_n365), .ZN(new_n373));
  AOI22_X1  g187(.A1(new_n362), .A2(new_n363), .B1(new_n367), .B2(new_n373), .ZN(new_n374));
  NAND3_X1  g188(.A1(new_n344), .A2(new_n359), .A3(new_n374), .ZN(new_n375));
  XNOR2_X1  g189(.A(G110), .B(G140), .ZN(new_n376));
  INV_X1    g190(.A(G227), .ZN(new_n377));
  NOR2_X1   g191(.A1(new_n377), .A2(G953), .ZN(new_n378));
  XOR2_X1   g192(.A(new_n376), .B(new_n378), .Z(new_n379));
  AND2_X1   g193(.A1(new_n375), .A2(new_n379), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n344), .A2(new_n374), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n381), .A2(new_n358), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n380), .A2(new_n382), .ZN(new_n383));
  INV_X1    g197(.A(new_n375), .ZN(new_n384));
  INV_X1    g198(.A(KEYINPUT12), .ZN(new_n385));
  INV_X1    g199(.A(new_n362), .ZN(new_n386));
  NOR2_X1   g200(.A1(new_n342), .A2(new_n343), .ZN(new_n387));
  AND3_X1   g201(.A1(new_n310), .A2(new_n312), .A3(new_n314), .ZN(new_n388));
  AOI21_X1  g202(.A(new_n386), .B1(new_n387), .B2(new_n388), .ZN(new_n389));
  OAI21_X1  g203(.A(new_n385), .B1(new_n389), .B2(new_n359), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n334), .A2(new_n341), .ZN(new_n391));
  INV_X1    g205(.A(KEYINPUT83), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n391), .A2(new_n392), .ZN(new_n393));
  NAND3_X1  g207(.A1(new_n334), .A2(KEYINPUT83), .A3(new_n341), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n393), .A2(new_n394), .ZN(new_n395));
  OAI21_X1  g209(.A(new_n362), .B1(new_n395), .B2(new_n315), .ZN(new_n396));
  NAND3_X1  g210(.A1(new_n396), .A2(KEYINPUT12), .A3(new_n358), .ZN(new_n397));
  AOI21_X1  g211(.A(new_n384), .B1(new_n390), .B2(new_n397), .ZN(new_n398));
  OAI21_X1  g212(.A(new_n383), .B1(new_n398), .B2(new_n379), .ZN(new_n399));
  AOI21_X1  g213(.A(new_n303), .B1(new_n399), .B2(new_n291), .ZN(new_n400));
  XNOR2_X1  g214(.A(KEYINPUT84), .B(G469), .ZN(new_n401));
  INV_X1    g215(.A(new_n401), .ZN(new_n402));
  INV_X1    g216(.A(new_n397), .ZN(new_n403));
  AOI21_X1  g217(.A(KEYINPUT12), .B1(new_n396), .B2(new_n358), .ZN(new_n404));
  OAI21_X1  g218(.A(new_n380), .B1(new_n403), .B2(new_n404), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n382), .A2(new_n375), .ZN(new_n406));
  INV_X1    g220(.A(new_n379), .ZN(new_n407));
  NAND2_X1  g221(.A1(new_n406), .A2(new_n407), .ZN(new_n408));
  AOI211_X1 g222(.A(G902), .B(new_n402), .C1(new_n405), .C2(new_n408), .ZN(new_n409));
  OAI21_X1  g223(.A(new_n302), .B1(new_n400), .B2(new_n409), .ZN(new_n410));
  INV_X1    g224(.A(new_n410), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n301), .A2(new_n411), .ZN(new_n412));
  INV_X1    g226(.A(new_n412), .ZN(new_n413));
  INV_X1    g227(.A(KEYINPUT78), .ZN(new_n414));
  NAND2_X1  g228(.A1(new_n267), .A2(G119), .ZN(new_n415));
  INV_X1    g229(.A(G119), .ZN(new_n416));
  NAND2_X1  g230(.A1(new_n416), .A2(G128), .ZN(new_n417));
  NAND2_X1  g231(.A1(new_n415), .A2(new_n417), .ZN(new_n418));
  XNOR2_X1  g232(.A(KEYINPUT24), .B(G110), .ZN(new_n419));
  NOR2_X1   g233(.A1(new_n418), .A2(new_n419), .ZN(new_n420));
  OR2_X1    g234(.A1(new_n420), .A2(KEYINPUT74), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n420), .A2(KEYINPUT74), .ZN(new_n422));
  INV_X1    g236(.A(KEYINPUT23), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n415), .A2(new_n423), .ZN(new_n424));
  NAND3_X1  g238(.A1(new_n267), .A2(KEYINPUT23), .A3(G119), .ZN(new_n425));
  NAND3_X1  g239(.A1(new_n424), .A2(new_n425), .A3(new_n417), .ZN(new_n426));
  AOI22_X1  g240(.A1(new_n421), .A2(new_n422), .B1(G110), .B2(new_n426), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n215), .A2(new_n427), .ZN(new_n428));
  AOI21_X1  g242(.A(new_n212), .B1(new_n201), .B2(new_n200), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n418), .A2(new_n419), .ZN(new_n430));
  OAI21_X1  g244(.A(new_n430), .B1(new_n426), .B2(G110), .ZN(new_n431));
  OR2_X1    g245(.A1(new_n431), .A2(KEYINPUT76), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n431), .A2(KEYINPUT76), .ZN(new_n433));
  NAND3_X1  g247(.A1(new_n429), .A2(new_n432), .A3(new_n433), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n428), .A2(new_n434), .ZN(new_n435));
  XNOR2_X1  g249(.A(KEYINPUT22), .B(G137), .ZN(new_n436));
  AND3_X1   g250(.A1(new_n192), .A2(G221), .A3(G234), .ZN(new_n437));
  XOR2_X1   g251(.A(new_n436), .B(new_n437), .Z(new_n438));
  NOR2_X1   g252(.A1(new_n435), .A2(new_n438), .ZN(new_n439));
  INV_X1    g253(.A(new_n438), .ZN(new_n440));
  AOI21_X1  g254(.A(new_n440), .B1(new_n428), .B2(new_n434), .ZN(new_n441));
  OAI21_X1  g255(.A(new_n291), .B1(new_n439), .B2(new_n441), .ZN(new_n442));
  OAI21_X1  g256(.A(new_n442), .B1(KEYINPUT77), .B2(KEYINPUT25), .ZN(new_n443));
  NOR2_X1   g257(.A1(KEYINPUT77), .A2(KEYINPUT25), .ZN(new_n444));
  OAI211_X1 g258(.A(new_n291), .B(new_n444), .C1(new_n439), .C2(new_n441), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n443), .A2(new_n445), .ZN(new_n446));
  NAND2_X1  g260(.A1(KEYINPUT77), .A2(KEYINPUT25), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n446), .A2(new_n447), .ZN(new_n448));
  AOI21_X1  g262(.A(new_n285), .B1(G234), .B2(new_n291), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n448), .A2(new_n449), .ZN(new_n450));
  OR2_X1    g264(.A1(new_n439), .A2(new_n441), .ZN(new_n451));
  NOR2_X1   g265(.A1(new_n449), .A2(G902), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n451), .A2(new_n452), .ZN(new_n453));
  AOI21_X1  g267(.A(new_n414), .B1(new_n450), .B2(new_n453), .ZN(new_n454));
  AOI22_X1  g268(.A1(new_n443), .A2(new_n445), .B1(KEYINPUT77), .B2(KEYINPUT25), .ZN(new_n455));
  INV_X1    g269(.A(new_n449), .ZN(new_n456));
  OAI211_X1 g270(.A(new_n414), .B(new_n453), .C1(new_n455), .C2(new_n456), .ZN(new_n457));
  INV_X1    g271(.A(new_n457), .ZN(new_n458));
  OR2_X1    g272(.A1(new_n454), .A2(new_n458), .ZN(new_n459));
  INV_X1    g273(.A(KEYINPUT29), .ZN(new_n460));
  XNOR2_X1  g274(.A(KEYINPUT26), .B(G101), .ZN(new_n461));
  NAND3_X1  g275(.A1(new_n191), .A2(new_n192), .A3(G210), .ZN(new_n462));
  XNOR2_X1  g276(.A(new_n461), .B(new_n462), .ZN(new_n463));
  XNOR2_X1  g277(.A(KEYINPUT70), .B(KEYINPUT27), .ZN(new_n464));
  XNOR2_X1  g278(.A(new_n463), .B(new_n464), .ZN(new_n465));
  INV_X1    g279(.A(new_n465), .ZN(new_n466));
  XNOR2_X1  g280(.A(G116), .B(G119), .ZN(new_n467));
  NOR2_X1   g281(.A1(new_n467), .A2(KEYINPUT69), .ZN(new_n468));
  XOR2_X1   g282(.A(KEYINPUT2), .B(G113), .Z(new_n469));
  XNOR2_X1  g283(.A(new_n468), .B(new_n469), .ZN(new_n470));
  INV_X1    g284(.A(KEYINPUT66), .ZN(new_n471));
  AOI21_X1  g285(.A(new_n471), .B1(new_n269), .B2(G137), .ZN(new_n472));
  INV_X1    g286(.A(new_n352), .ZN(new_n473));
  NOR2_X1   g287(.A1(new_n472), .A2(new_n473), .ZN(new_n474));
  NOR2_X1   g288(.A1(new_n352), .A2(new_n471), .ZN(new_n475));
  OAI21_X1  g289(.A(G131), .B1(new_n474), .B2(new_n475), .ZN(new_n476));
  NAND4_X1  g290(.A1(new_n356), .A2(new_n195), .A3(new_n348), .A4(new_n349), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  OAI21_X1  g292(.A(KEYINPUT68), .B1(new_n388), .B2(new_n478), .ZN(new_n479));
  INV_X1    g293(.A(KEYINPUT30), .ZN(new_n480));
  NAND2_X1  g294(.A1(new_n358), .A2(new_n371), .ZN(new_n481));
  INV_X1    g295(.A(KEYINPUT68), .ZN(new_n482));
  NAND4_X1  g296(.A1(new_n315), .A2(new_n482), .A3(new_n476), .A4(new_n477), .ZN(new_n483));
  NAND4_X1  g297(.A1(new_n479), .A2(new_n480), .A3(new_n481), .A4(new_n483), .ZN(new_n484));
  OAI21_X1  g298(.A(new_n481), .B1(new_n388), .B2(new_n478), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n485), .A2(KEYINPUT30), .ZN(new_n486));
  AOI21_X1  g300(.A(new_n470), .B1(new_n484), .B2(new_n486), .ZN(new_n487));
  OAI211_X1 g301(.A(new_n481), .B(new_n470), .C1(new_n388), .C2(new_n478), .ZN(new_n488));
  INV_X1    g302(.A(new_n488), .ZN(new_n489));
  OAI21_X1  g303(.A(new_n466), .B1(new_n487), .B2(new_n489), .ZN(new_n490));
  NOR2_X1   g304(.A1(new_n489), .A2(KEYINPUT28), .ZN(new_n491));
  INV_X1    g305(.A(new_n491), .ZN(new_n492));
  INV_X1    g306(.A(new_n470), .ZN(new_n493));
  NAND3_X1  g307(.A1(new_n479), .A2(new_n481), .A3(new_n483), .ZN(new_n494));
  AOI21_X1  g308(.A(new_n489), .B1(new_n493), .B2(new_n494), .ZN(new_n495));
  INV_X1    g309(.A(KEYINPUT28), .ZN(new_n496));
  OAI21_X1  g310(.A(new_n492), .B1(new_n495), .B2(new_n496), .ZN(new_n497));
  OAI211_X1 g311(.A(new_n460), .B(new_n490), .C1(new_n497), .C2(new_n466), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n485), .A2(new_n493), .ZN(new_n499));
  NAND2_X1  g313(.A1(new_n499), .A2(new_n488), .ZN(new_n500));
  AOI21_X1  g314(.A(new_n491), .B1(new_n500), .B2(KEYINPUT28), .ZN(new_n501));
  NOR2_X1   g315(.A1(new_n466), .A2(new_n460), .ZN(new_n502));
  AOI21_X1  g316(.A(G902), .B1(new_n501), .B2(new_n502), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n498), .A2(new_n503), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n504), .A2(G472), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n494), .A2(new_n493), .ZN(new_n506));
  AOI21_X1  g320(.A(new_n496), .B1(new_n506), .B2(new_n488), .ZN(new_n507));
  OAI21_X1  g321(.A(new_n466), .B1(new_n507), .B2(new_n491), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n488), .A2(new_n465), .ZN(new_n509));
  NAND2_X1  g323(.A1(new_n509), .A2(KEYINPUT71), .ZN(new_n510));
  INV_X1    g324(.A(KEYINPUT71), .ZN(new_n511));
  NAND3_X1  g325(.A1(new_n488), .A2(new_n511), .A3(new_n465), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n510), .A2(new_n512), .ZN(new_n513));
  OAI21_X1  g327(.A(KEYINPUT31), .B1(new_n513), .B2(new_n487), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n484), .A2(new_n486), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n515), .A2(new_n493), .ZN(new_n516));
  INV_X1    g330(.A(KEYINPUT31), .ZN(new_n517));
  NAND4_X1  g331(.A1(new_n516), .A2(new_n517), .A3(new_n510), .A4(new_n512), .ZN(new_n518));
  NAND3_X1  g332(.A1(new_n508), .A2(new_n514), .A3(new_n518), .ZN(new_n519));
  INV_X1    g333(.A(KEYINPUT32), .ZN(new_n520));
  NOR2_X1   g334(.A1(G472), .A2(G902), .ZN(new_n521));
  XNOR2_X1  g335(.A(new_n521), .B(KEYINPUT72), .ZN(new_n522));
  AND3_X1   g336(.A1(new_n519), .A2(new_n520), .A3(new_n522), .ZN(new_n523));
  AOI21_X1  g337(.A(new_n520), .B1(new_n519), .B2(new_n522), .ZN(new_n524));
  OAI21_X1  g338(.A(new_n505), .B1(new_n523), .B2(new_n524), .ZN(new_n525));
  INV_X1    g339(.A(KEYINPUT73), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  OAI211_X1 g341(.A(new_n505), .B(KEYINPUT73), .C1(new_n523), .C2(new_n524), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  NOR2_X1   g343(.A1(new_n459), .A2(new_n529), .ZN(new_n530));
  INV_X1    g344(.A(G113), .ZN(new_n531));
  XNOR2_X1  g345(.A(KEYINPUT85), .B(KEYINPUT5), .ZN(new_n532));
  NOR2_X1   g346(.A1(new_n252), .A2(G119), .ZN(new_n533));
  AOI21_X1  g347(.A(new_n531), .B1(new_n532), .B2(new_n533), .ZN(new_n534));
  INV_X1    g348(.A(new_n467), .ZN(new_n535));
  OAI21_X1  g349(.A(new_n534), .B1(new_n535), .B2(new_n532), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n469), .A2(new_n467), .ZN(new_n537));
  NAND2_X1  g351(.A1(new_n536), .A2(new_n537), .ZN(new_n538));
  AOI21_X1  g352(.A(new_n538), .B1(new_n393), .B2(new_n394), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n364), .A2(new_n365), .ZN(new_n540));
  NAND3_X1  g354(.A1(new_n367), .A2(new_n493), .A3(new_n540), .ZN(new_n541));
  INV_X1    g355(.A(new_n541), .ZN(new_n542));
  OAI21_X1  g356(.A(KEYINPUT86), .B1(new_n539), .B2(new_n542), .ZN(new_n543));
  INV_X1    g357(.A(KEYINPUT6), .ZN(new_n544));
  INV_X1    g358(.A(new_n538), .ZN(new_n545));
  OAI21_X1  g359(.A(new_n545), .B1(new_n342), .B2(new_n343), .ZN(new_n546));
  INV_X1    g360(.A(KEYINPUT86), .ZN(new_n547));
  NAND3_X1  g361(.A1(new_n546), .A2(new_n547), .A3(new_n541), .ZN(new_n548));
  XNOR2_X1  g362(.A(G110), .B(G122), .ZN(new_n549));
  XOR2_X1   g363(.A(new_n549), .B(KEYINPUT87), .Z(new_n550));
  NAND4_X1  g364(.A1(new_n543), .A2(new_n544), .A3(new_n548), .A4(new_n550), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n551), .A2(KEYINPUT88), .ZN(new_n552));
  INV_X1    g366(.A(new_n550), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n546), .A2(new_n541), .ZN(new_n554));
  AOI21_X1  g368(.A(new_n553), .B1(new_n554), .B2(KEYINPUT86), .ZN(new_n555));
  INV_X1    g369(.A(KEYINPUT88), .ZN(new_n556));
  NAND4_X1  g370(.A1(new_n555), .A2(new_n556), .A3(new_n544), .A4(new_n548), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n552), .A2(new_n557), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n555), .A2(new_n548), .ZN(new_n559));
  NAND3_X1  g373(.A1(new_n546), .A2(new_n541), .A3(new_n549), .ZN(new_n560));
  AND2_X1   g374(.A1(new_n560), .A2(KEYINPUT6), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n559), .A2(new_n561), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n372), .A2(G125), .ZN(new_n563));
  OR2_X1    g377(.A1(new_n563), .A2(KEYINPUT89), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n388), .A2(new_n208), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n563), .A2(KEYINPUT89), .ZN(new_n566));
  AND3_X1   g380(.A1(new_n564), .A2(new_n565), .A3(new_n566), .ZN(new_n567));
  INV_X1    g381(.A(G224), .ZN(new_n568));
  NOR2_X1   g382(.A1(new_n568), .A2(G953), .ZN(new_n569));
  XOR2_X1   g383(.A(new_n567), .B(new_n569), .Z(new_n570));
  NAND3_X1  g384(.A1(new_n558), .A2(new_n562), .A3(new_n570), .ZN(new_n571));
  INV_X1    g385(.A(KEYINPUT7), .ZN(new_n572));
  NOR2_X1   g386(.A1(new_n569), .A2(new_n572), .ZN(new_n573));
  AOI21_X1  g387(.A(new_n573), .B1(new_n565), .B2(new_n563), .ZN(new_n574));
  AOI21_X1  g388(.A(new_n574), .B1(new_n567), .B2(new_n573), .ZN(new_n575));
  AND2_X1   g389(.A1(new_n560), .A2(new_n575), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n391), .A2(new_n538), .ZN(new_n577));
  INV_X1    g391(.A(KEYINPUT5), .ZN(new_n578));
  OAI21_X1  g392(.A(new_n534), .B1(new_n578), .B2(new_n535), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n579), .A2(new_n537), .ZN(new_n580));
  OAI21_X1  g394(.A(new_n577), .B1(new_n387), .B2(new_n580), .ZN(new_n581));
  NOR2_X1   g395(.A1(new_n549), .A2(KEYINPUT8), .ZN(new_n582));
  AND2_X1   g396(.A1(new_n549), .A2(KEYINPUT8), .ZN(new_n583));
  OAI21_X1  g397(.A(new_n581), .B1(new_n582), .B2(new_n583), .ZN(new_n584));
  AOI21_X1  g398(.A(G902), .B1(new_n576), .B2(new_n584), .ZN(new_n585));
  OAI21_X1  g399(.A(G210), .B1(G237), .B2(G902), .ZN(new_n586));
  INV_X1    g400(.A(new_n586), .ZN(new_n587));
  NAND2_X1  g401(.A1(new_n587), .A2(KEYINPUT90), .ZN(new_n588));
  AND3_X1   g402(.A1(new_n571), .A2(new_n585), .A3(new_n588), .ZN(new_n589));
  AOI21_X1  g403(.A(new_n588), .B1(new_n571), .B2(new_n585), .ZN(new_n590));
  NOR2_X1   g404(.A1(new_n589), .A2(new_n590), .ZN(new_n591));
  OAI21_X1  g405(.A(G214), .B1(G237), .B2(G902), .ZN(new_n592));
  INV_X1    g406(.A(new_n592), .ZN(new_n593));
  NOR2_X1   g407(.A1(new_n591), .A2(new_n593), .ZN(new_n594));
  NAND3_X1  g408(.A1(new_n413), .A2(new_n530), .A3(new_n594), .ZN(new_n595));
  XNOR2_X1  g409(.A(new_n595), .B(G101), .ZN(G3));
  INV_X1    g410(.A(new_n585), .ZN(new_n597));
  AOI22_X1  g411(.A1(new_n552), .A2(new_n557), .B1(new_n559), .B2(new_n561), .ZN(new_n598));
  AOI211_X1 g412(.A(new_n587), .B(new_n597), .C1(new_n598), .C2(new_n570), .ZN(new_n599));
  AOI21_X1  g413(.A(new_n586), .B1(new_n571), .B2(new_n585), .ZN(new_n600));
  OAI21_X1  g414(.A(new_n592), .B1(new_n599), .B2(new_n600), .ZN(new_n601));
  INV_X1    g415(.A(KEYINPUT98), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n601), .A2(new_n602), .ZN(new_n603));
  OAI211_X1 g417(.A(KEYINPUT98), .B(new_n592), .C1(new_n599), .C2(new_n600), .ZN(new_n604));
  AND2_X1   g418(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  NAND2_X1  g419(.A1(new_n292), .A2(new_n293), .ZN(new_n606));
  NOR2_X1   g420(.A1(new_n290), .A2(KEYINPUT33), .ZN(new_n607));
  INV_X1    g421(.A(KEYINPUT99), .ZN(new_n608));
  AOI21_X1  g422(.A(new_n608), .B1(new_n273), .B2(new_n282), .ZN(new_n609));
  NAND2_X1  g423(.A1(new_n609), .A2(new_n287), .ZN(new_n610));
  INV_X1    g424(.A(KEYINPUT100), .ZN(new_n611));
  NAND2_X1  g425(.A1(new_n289), .A2(new_n611), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n286), .A2(KEYINPUT100), .ZN(new_n613));
  OAI211_X1 g427(.A(new_n610), .B(new_n612), .C1(new_n609), .C2(new_n613), .ZN(new_n614));
  AOI21_X1  g428(.A(new_n607), .B1(new_n614), .B2(KEYINPUT33), .ZN(new_n615));
  NOR2_X1   g429(.A1(new_n293), .A2(G902), .ZN(new_n616));
  INV_X1    g430(.A(new_n616), .ZN(new_n617));
  OAI21_X1  g431(.A(new_n606), .B1(new_n615), .B2(new_n617), .ZN(new_n618));
  INV_X1    g432(.A(new_n618), .ZN(new_n619));
  NOR2_X1   g433(.A1(new_n243), .A2(new_n619), .ZN(new_n620));
  NAND3_X1  g434(.A1(new_n605), .A2(new_n251), .A3(new_n620), .ZN(new_n621));
  NAND2_X1  g435(.A1(new_n519), .A2(new_n522), .ZN(new_n622));
  INV_X1    g436(.A(new_n622), .ZN(new_n623));
  INV_X1    g437(.A(G472), .ZN(new_n624));
  AOI21_X1  g438(.A(new_n624), .B1(new_n519), .B2(new_n291), .ZN(new_n625));
  NOR2_X1   g439(.A1(new_n623), .A2(new_n625), .ZN(new_n626));
  INV_X1    g440(.A(new_n626), .ZN(new_n627));
  NOR3_X1   g441(.A1(new_n459), .A2(new_n410), .A3(new_n627), .ZN(new_n628));
  INV_X1    g442(.A(new_n628), .ZN(new_n629));
  NOR2_X1   g443(.A1(new_n621), .A2(new_n629), .ZN(new_n630));
  XNOR2_X1  g444(.A(KEYINPUT34), .B(G104), .ZN(new_n631));
  XNOR2_X1  g445(.A(new_n630), .B(new_n631), .ZN(G6));
  INV_X1    g446(.A(new_n297), .ZN(new_n633));
  NAND4_X1  g447(.A1(new_n605), .A2(new_n251), .A3(new_n243), .A4(new_n633), .ZN(new_n634));
  NOR2_X1   g448(.A1(new_n634), .A2(new_n629), .ZN(new_n635));
  XNOR2_X1  g449(.A(KEYINPUT35), .B(G107), .ZN(new_n636));
  XNOR2_X1  g450(.A(new_n635), .B(new_n636), .ZN(G9));
  INV_X1    g451(.A(KEYINPUT102), .ZN(new_n638));
  AOI21_X1  g452(.A(KEYINPUT101), .B1(new_n428), .B2(new_n434), .ZN(new_n639));
  INV_X1    g453(.A(new_n639), .ZN(new_n640));
  NAND3_X1  g454(.A1(new_n428), .A2(KEYINPUT101), .A3(new_n434), .ZN(new_n641));
  OAI211_X1 g455(.A(new_n640), .B(new_n641), .C1(KEYINPUT36), .C2(new_n440), .ZN(new_n642));
  NOR2_X1   g456(.A1(new_n440), .A2(KEYINPUT36), .ZN(new_n643));
  INV_X1    g457(.A(new_n641), .ZN(new_n644));
  OAI21_X1  g458(.A(new_n643), .B1(new_n644), .B2(new_n639), .ZN(new_n645));
  NAND2_X1  g459(.A1(new_n642), .A2(new_n645), .ZN(new_n646));
  INV_X1    g460(.A(new_n646), .ZN(new_n647));
  INV_X1    g461(.A(new_n452), .ZN(new_n648));
  OAI21_X1  g462(.A(new_n638), .B1(new_n647), .B2(new_n648), .ZN(new_n649));
  NAND3_X1  g463(.A1(new_n646), .A2(KEYINPUT102), .A3(new_n452), .ZN(new_n650));
  NAND2_X1  g464(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  NAND2_X1  g465(.A1(new_n651), .A2(new_n450), .ZN(new_n652));
  NAND4_X1  g466(.A1(new_n413), .A2(new_n594), .A3(new_n626), .A4(new_n652), .ZN(new_n653));
  XOR2_X1   g467(.A(KEYINPUT37), .B(G110), .Z(new_n654));
  XNOR2_X1  g468(.A(new_n653), .B(new_n654), .ZN(G12));
  NAND3_X1  g469(.A1(new_n527), .A2(new_n528), .A3(new_n652), .ZN(new_n656));
  NOR2_X1   g470(.A1(new_n656), .A2(new_n410), .ZN(new_n657));
  NAND2_X1  g471(.A1(new_n243), .A2(new_n633), .ZN(new_n658));
  INV_X1    g472(.A(G900), .ZN(new_n659));
  AOI21_X1  g473(.A(new_n246), .B1(new_n248), .B2(new_n659), .ZN(new_n660));
  NOR2_X1   g474(.A1(new_n658), .A2(new_n660), .ZN(new_n661));
  NAND4_X1  g475(.A1(new_n603), .A2(new_n657), .A3(new_n604), .A4(new_n661), .ZN(new_n662));
  XNOR2_X1  g476(.A(new_n662), .B(G128), .ZN(G30));
  NOR2_X1   g477(.A1(new_n513), .A2(new_n487), .ZN(new_n664));
  AOI21_X1  g478(.A(new_n664), .B1(new_n466), .B2(new_n500), .ZN(new_n665));
  OAI21_X1  g479(.A(G472), .B1(new_n665), .B2(G902), .ZN(new_n666));
  OAI21_X1  g480(.A(new_n666), .B1(new_n523), .B2(new_n524), .ZN(new_n667));
  INV_X1    g481(.A(new_n667), .ZN(new_n668));
  NOR2_X1   g482(.A1(new_n243), .A2(new_n297), .ZN(new_n669));
  AOI22_X1  g483(.A1(new_n649), .A2(new_n650), .B1(new_n448), .B2(new_n449), .ZN(new_n670));
  NAND3_X1  g484(.A1(new_n669), .A2(new_n592), .A3(new_n670), .ZN(new_n671));
  XOR2_X1   g485(.A(new_n660), .B(KEYINPUT39), .Z(new_n672));
  NAND2_X1  g486(.A1(new_n411), .A2(new_n672), .ZN(new_n673));
  AOI211_X1 g487(.A(new_n668), .B(new_n671), .C1(new_n673), .C2(KEYINPUT40), .ZN(new_n674));
  OAI21_X1  g488(.A(new_n674), .B1(KEYINPUT40), .B2(new_n673), .ZN(new_n675));
  XOR2_X1   g489(.A(KEYINPUT103), .B(KEYINPUT38), .Z(new_n676));
  XOR2_X1   g490(.A(new_n591), .B(new_n676), .Z(new_n677));
  NOR2_X1   g491(.A1(new_n675), .A2(new_n677), .ZN(new_n678));
  XNOR2_X1  g492(.A(new_n678), .B(KEYINPUT104), .ZN(new_n679));
  XNOR2_X1  g493(.A(new_n679), .B(G143), .ZN(G45));
  INV_X1    g494(.A(new_n660), .ZN(new_n681));
  NAND3_X1  g495(.A1(new_n242), .A2(new_n618), .A3(new_n681), .ZN(new_n682));
  NOR3_X1   g496(.A1(new_n656), .A2(new_n410), .A3(new_n682), .ZN(new_n683));
  NAND3_X1  g497(.A1(new_n683), .A2(new_n603), .A3(new_n604), .ZN(new_n684));
  XNOR2_X1  g498(.A(new_n684), .B(G146), .ZN(G48));
  AOI21_X1  g499(.A(G902), .B1(new_n405), .B2(new_n408), .ZN(new_n686));
  NOR2_X1   g500(.A1(new_n686), .A2(new_n303), .ZN(new_n687));
  NOR2_X1   g501(.A1(new_n687), .A2(new_n409), .ZN(new_n688));
  NAND2_X1  g502(.A1(new_n688), .A2(new_n302), .ZN(new_n689));
  INV_X1    g503(.A(new_n689), .ZN(new_n690));
  NAND2_X1  g504(.A1(new_n530), .A2(new_n690), .ZN(new_n691));
  NOR2_X1   g505(.A1(new_n621), .A2(new_n691), .ZN(new_n692));
  XOR2_X1   g506(.A(KEYINPUT41), .B(G113), .Z(new_n693));
  XNOR2_X1  g507(.A(new_n692), .B(new_n693), .ZN(G15));
  OR2_X1    g508(.A1(new_n634), .A2(new_n691), .ZN(new_n695));
  XNOR2_X1  g509(.A(new_n695), .B(G116), .ZN(G18));
  AOI21_X1  g510(.A(new_n656), .B1(new_n298), .B2(new_n300), .ZN(new_n697));
  NAND3_X1  g511(.A1(new_n605), .A2(new_n690), .A3(new_n697), .ZN(new_n698));
  XNOR2_X1  g512(.A(new_n698), .B(KEYINPUT105), .ZN(new_n699));
  XNOR2_X1  g513(.A(new_n699), .B(G119), .ZN(G21));
  AND2_X1   g514(.A1(new_n450), .A2(new_n453), .ZN(new_n701));
  OAI211_X1 g515(.A(new_n518), .B(new_n514), .C1(new_n465), .C2(new_n501), .ZN(new_n702));
  AOI21_X1  g516(.A(new_n625), .B1(new_n522), .B2(new_n702), .ZN(new_n703));
  NAND2_X1  g517(.A1(new_n701), .A2(new_n703), .ZN(new_n704));
  NOR3_X1   g518(.A1(new_n689), .A2(new_n704), .A3(new_n250), .ZN(new_n705));
  NAND3_X1  g519(.A1(new_n605), .A2(new_n669), .A3(new_n705), .ZN(new_n706));
  XNOR2_X1  g520(.A(new_n706), .B(G122), .ZN(G24));
  INV_X1    g521(.A(new_n682), .ZN(new_n708));
  AND3_X1   g522(.A1(new_n708), .A2(new_n652), .A3(new_n703), .ZN(new_n709));
  NAND4_X1  g523(.A1(new_n603), .A2(new_n690), .A3(new_n709), .A4(new_n604), .ZN(new_n710));
  XNOR2_X1  g524(.A(new_n710), .B(G125), .ZN(G27));
  NOR3_X1   g525(.A1(new_n589), .A2(new_n590), .A3(new_n593), .ZN(new_n712));
  NAND2_X1  g526(.A1(new_n712), .A2(new_n411), .ZN(new_n713));
  AND2_X1   g527(.A1(new_n701), .A2(new_n525), .ZN(new_n714));
  NAND2_X1  g528(.A1(new_n714), .A2(new_n708), .ZN(new_n715));
  OAI21_X1  g529(.A(KEYINPUT42), .B1(new_n713), .B2(new_n715), .ZN(new_n716));
  NOR2_X1   g530(.A1(new_n682), .A2(KEYINPUT42), .ZN(new_n717));
  NAND4_X1  g531(.A1(new_n530), .A2(new_n712), .A3(new_n411), .A4(new_n717), .ZN(new_n718));
  AND2_X1   g532(.A1(new_n716), .A2(new_n718), .ZN(new_n719));
  XNOR2_X1  g533(.A(new_n719), .B(G131), .ZN(G33));
  NAND4_X1  g534(.A1(new_n530), .A2(new_n712), .A3(new_n411), .A4(new_n661), .ZN(new_n721));
  XNOR2_X1  g535(.A(new_n721), .B(G134), .ZN(G36));
  NOR2_X1   g536(.A1(new_n619), .A2(new_n242), .ZN(new_n723));
  XNOR2_X1  g537(.A(new_n723), .B(KEYINPUT43), .ZN(new_n724));
  INV_X1    g538(.A(KEYINPUT106), .ZN(new_n725));
  XNOR2_X1  g539(.A(new_n724), .B(new_n725), .ZN(new_n726));
  NAND3_X1  g540(.A1(new_n726), .A2(new_n627), .A3(new_n652), .ZN(new_n727));
  INV_X1    g541(.A(KEYINPUT44), .ZN(new_n728));
  NOR2_X1   g542(.A1(new_n727), .A2(new_n728), .ZN(new_n729));
  XNOR2_X1  g543(.A(new_n729), .B(KEYINPUT107), .ZN(new_n730));
  XNOR2_X1  g544(.A(new_n712), .B(KEYINPUT108), .ZN(new_n731));
  NAND2_X1  g545(.A1(new_n727), .A2(new_n728), .ZN(new_n732));
  NAND3_X1  g546(.A1(new_n730), .A2(new_n731), .A3(new_n732), .ZN(new_n733));
  INV_X1    g547(.A(new_n302), .ZN(new_n734));
  XNOR2_X1  g548(.A(new_n399), .B(KEYINPUT45), .ZN(new_n735));
  OAI21_X1  g549(.A(G469), .B1(new_n735), .B2(G902), .ZN(new_n736));
  OR2_X1    g550(.A1(new_n736), .A2(KEYINPUT46), .ZN(new_n737));
  AOI21_X1  g551(.A(new_n409), .B1(new_n736), .B2(KEYINPUT46), .ZN(new_n738));
  AOI21_X1  g552(.A(new_n734), .B1(new_n737), .B2(new_n738), .ZN(new_n739));
  AND2_X1   g553(.A1(new_n739), .A2(new_n672), .ZN(new_n740));
  INV_X1    g554(.A(new_n740), .ZN(new_n741));
  OR2_X1    g555(.A1(new_n733), .A2(new_n741), .ZN(new_n742));
  XNOR2_X1  g556(.A(new_n742), .B(G137), .ZN(G39));
  XNOR2_X1  g557(.A(new_n739), .B(KEYINPUT47), .ZN(new_n744));
  INV_X1    g558(.A(new_n459), .ZN(new_n745));
  NOR2_X1   g559(.A1(new_n745), .A2(new_n682), .ZN(new_n746));
  NAND4_X1  g560(.A1(new_n744), .A2(new_n529), .A3(new_n712), .A4(new_n746), .ZN(new_n747));
  XNOR2_X1  g561(.A(new_n747), .B(G140), .ZN(G42));
  OAI21_X1  g562(.A(new_n658), .B1(new_n243), .B2(new_n619), .ZN(new_n749));
  NAND4_X1  g563(.A1(new_n628), .A2(new_n594), .A3(new_n251), .A4(new_n749), .ZN(new_n750));
  NAND4_X1  g564(.A1(new_n706), .A2(new_n595), .A3(new_n653), .A4(new_n750), .ZN(new_n751));
  NOR2_X1   g565(.A1(new_n751), .A2(new_n692), .ZN(new_n752));
  NAND3_X1  g566(.A1(new_n709), .A2(new_n411), .A3(new_n712), .ZN(new_n753));
  NAND4_X1  g567(.A1(new_n716), .A2(new_n718), .A3(new_n721), .A4(new_n753), .ZN(new_n754));
  NOR2_X1   g568(.A1(new_n299), .A2(new_n660), .ZN(new_n755));
  NAND3_X1  g569(.A1(new_n712), .A2(KEYINPUT110), .A3(new_n755), .ZN(new_n756));
  NAND2_X1  g570(.A1(new_n756), .A2(new_n657), .ZN(new_n757));
  AOI21_X1  g571(.A(KEYINPUT110), .B1(new_n712), .B2(new_n755), .ZN(new_n758));
  NOR2_X1   g572(.A1(new_n757), .A2(new_n758), .ZN(new_n759));
  NOR2_X1   g573(.A1(new_n754), .A2(new_n759), .ZN(new_n760));
  NAND4_X1  g574(.A1(new_n752), .A2(new_n699), .A3(new_n760), .A4(new_n695), .ZN(new_n761));
  NAND3_X1  g575(.A1(new_n670), .A2(new_n681), .A3(new_n667), .ZN(new_n762));
  NOR2_X1   g576(.A1(new_n410), .A2(new_n762), .ZN(new_n763));
  NAND4_X1  g577(.A1(new_n603), .A2(new_n604), .A3(new_n669), .A4(new_n763), .ZN(new_n764));
  NAND4_X1  g578(.A1(new_n662), .A2(new_n710), .A3(new_n764), .A4(new_n684), .ZN(new_n765));
  INV_X1    g579(.A(KEYINPUT52), .ZN(new_n766));
  NAND2_X1  g580(.A1(new_n765), .A2(new_n766), .ZN(new_n767));
  INV_X1    g581(.A(KEYINPUT111), .ZN(new_n768));
  NAND2_X1  g582(.A1(new_n767), .A2(new_n768), .ZN(new_n769));
  AND3_X1   g583(.A1(new_n662), .A2(new_n710), .A3(new_n684), .ZN(new_n770));
  NAND3_X1  g584(.A1(new_n770), .A2(KEYINPUT52), .A3(new_n764), .ZN(new_n771));
  NAND3_X1  g585(.A1(new_n765), .A2(KEYINPUT111), .A3(new_n766), .ZN(new_n772));
  NAND3_X1  g586(.A1(new_n769), .A2(new_n771), .A3(new_n772), .ZN(new_n773));
  NAND2_X1  g587(.A1(new_n773), .A2(KEYINPUT112), .ZN(new_n774));
  INV_X1    g588(.A(KEYINPUT112), .ZN(new_n775));
  NAND4_X1  g589(.A1(new_n769), .A2(new_n771), .A3(new_n775), .A4(new_n772), .ZN(new_n776));
  AOI21_X1  g590(.A(new_n761), .B1(new_n774), .B2(new_n776), .ZN(new_n777));
  INV_X1    g591(.A(KEYINPUT53), .ZN(new_n778));
  NAND2_X1  g592(.A1(new_n777), .A2(new_n778), .ZN(new_n779));
  INV_X1    g593(.A(new_n761), .ZN(new_n780));
  NAND2_X1  g594(.A1(new_n771), .A2(new_n767), .ZN(new_n781));
  NAND2_X1  g595(.A1(new_n780), .A2(new_n781), .ZN(new_n782));
  NAND2_X1  g596(.A1(new_n782), .A2(KEYINPUT53), .ZN(new_n783));
  AND3_X1   g597(.A1(new_n779), .A2(KEYINPUT54), .A3(new_n783), .ZN(new_n784));
  AOI21_X1  g598(.A(KEYINPUT53), .B1(new_n780), .B2(new_n781), .ZN(new_n785));
  NOR2_X1   g599(.A1(new_n765), .A2(new_n766), .ZN(new_n786));
  AOI21_X1  g600(.A(new_n786), .B1(new_n768), .B2(new_n767), .ZN(new_n787));
  AOI21_X1  g601(.A(new_n775), .B1(new_n787), .B2(new_n772), .ZN(new_n788));
  INV_X1    g602(.A(new_n776), .ZN(new_n789));
  OAI211_X1 g603(.A(KEYINPUT53), .B(new_n780), .C1(new_n788), .C2(new_n789), .ZN(new_n790));
  NAND2_X1  g604(.A1(new_n790), .A2(KEYINPUT113), .ZN(new_n791));
  INV_X1    g605(.A(KEYINPUT113), .ZN(new_n792));
  NAND3_X1  g606(.A1(new_n777), .A2(new_n792), .A3(KEYINPUT53), .ZN(new_n793));
  AOI211_X1 g607(.A(KEYINPUT54), .B(new_n785), .C1(new_n791), .C2(new_n793), .ZN(new_n794));
  INV_X1    g608(.A(KEYINPUT114), .ZN(new_n795));
  AOI21_X1  g609(.A(new_n784), .B1(new_n794), .B2(new_n795), .ZN(new_n796));
  INV_X1    g610(.A(KEYINPUT54), .ZN(new_n797));
  INV_X1    g611(.A(new_n785), .ZN(new_n798));
  NOR2_X1   g612(.A1(new_n790), .A2(KEYINPUT113), .ZN(new_n799));
  AOI21_X1  g613(.A(new_n792), .B1(new_n777), .B2(KEYINPUT53), .ZN(new_n800));
  OAI211_X1 g614(.A(new_n797), .B(new_n798), .C1(new_n799), .C2(new_n800), .ZN(new_n801));
  NAND2_X1  g615(.A1(new_n801), .A2(KEYINPUT114), .ZN(new_n802));
  NAND3_X1  g616(.A1(new_n745), .A2(new_n246), .A3(new_n668), .ZN(new_n803));
  NAND2_X1  g617(.A1(new_n690), .A2(new_n712), .ZN(new_n804));
  NOR2_X1   g618(.A1(new_n803), .A2(new_n804), .ZN(new_n805));
  XNOR2_X1  g619(.A(new_n805), .B(KEYINPUT116), .ZN(new_n806));
  NAND2_X1  g620(.A1(new_n806), .A2(new_n620), .ZN(new_n807));
  NAND2_X1  g621(.A1(new_n724), .A2(new_n246), .ZN(new_n808));
  NOR2_X1   g622(.A1(new_n808), .A2(new_n704), .ZN(new_n809));
  NAND3_X1  g623(.A1(new_n809), .A2(new_n605), .A3(new_n690), .ZN(new_n810));
  NAND4_X1  g624(.A1(new_n807), .A2(G952), .A3(new_n192), .A4(new_n810), .ZN(new_n811));
  NOR2_X1   g625(.A1(new_n808), .A2(new_n804), .ZN(new_n812));
  NAND2_X1  g626(.A1(new_n812), .A2(new_n714), .ZN(new_n813));
  NOR2_X1   g627(.A1(new_n813), .A2(KEYINPUT48), .ZN(new_n814));
  XNOR2_X1  g628(.A(new_n814), .B(KEYINPUT117), .ZN(new_n815));
  NAND2_X1  g629(.A1(new_n813), .A2(KEYINPUT48), .ZN(new_n816));
  XNOR2_X1  g630(.A(new_n816), .B(KEYINPUT118), .ZN(new_n817));
  AOI21_X1  g631(.A(new_n811), .B1(new_n815), .B2(new_n817), .ZN(new_n818));
  XOR2_X1   g632(.A(new_n818), .B(KEYINPUT119), .Z(new_n819));
  NAND4_X1  g633(.A1(new_n809), .A2(new_n593), .A3(new_n677), .A4(new_n690), .ZN(new_n820));
  XOR2_X1   g634(.A(new_n820), .B(KEYINPUT50), .Z(new_n821));
  NAND3_X1  g635(.A1(new_n806), .A2(new_n243), .A3(new_n619), .ZN(new_n822));
  NAND3_X1  g636(.A1(new_n812), .A2(new_n652), .A3(new_n703), .ZN(new_n823));
  NAND3_X1  g637(.A1(new_n821), .A2(new_n822), .A3(new_n823), .ZN(new_n824));
  NAND2_X1  g638(.A1(new_n809), .A2(new_n731), .ZN(new_n825));
  INV_X1    g639(.A(new_n744), .ZN(new_n826));
  NAND2_X1  g640(.A1(new_n688), .A2(new_n734), .ZN(new_n827));
  AOI21_X1  g641(.A(new_n825), .B1(new_n826), .B2(new_n827), .ZN(new_n828));
  INV_X1    g642(.A(KEYINPUT51), .ZN(new_n829));
  NOR3_X1   g643(.A1(new_n824), .A2(new_n828), .A3(new_n829), .ZN(new_n830));
  XNOR2_X1  g644(.A(new_n827), .B(KEYINPUT115), .ZN(new_n831));
  AOI21_X1  g645(.A(new_n825), .B1(new_n826), .B2(new_n831), .ZN(new_n832));
  OR2_X1    g646(.A1(new_n824), .A2(new_n832), .ZN(new_n833));
  AOI21_X1  g647(.A(new_n830), .B1(new_n829), .B2(new_n833), .ZN(new_n834));
  NAND4_X1  g648(.A1(new_n796), .A2(new_n802), .A3(new_n819), .A4(new_n834), .ZN(new_n835));
  OAI21_X1  g649(.A(new_n835), .B1(G952), .B2(G953), .ZN(new_n836));
  NAND4_X1  g650(.A1(new_n723), .A2(new_n701), .A3(new_n592), .A4(new_n302), .ZN(new_n837));
  XOR2_X1   g651(.A(new_n837), .B(KEYINPUT109), .Z(new_n838));
  NOR2_X1   g652(.A1(new_n838), .A2(new_n667), .ZN(new_n839));
  OR3_X1    g653(.A1(new_n687), .A2(new_n409), .A3(KEYINPUT49), .ZN(new_n840));
  OAI21_X1  g654(.A(KEYINPUT49), .B1(new_n687), .B2(new_n409), .ZN(new_n841));
  NAND4_X1  g655(.A1(new_n839), .A2(new_n677), .A3(new_n840), .A4(new_n841), .ZN(new_n842));
  NAND2_X1  g656(.A1(new_n836), .A2(new_n842), .ZN(G75));
  INV_X1    g657(.A(KEYINPUT120), .ZN(new_n844));
  NAND2_X1  g658(.A1(new_n791), .A2(new_n793), .ZN(new_n845));
  AOI21_X1  g659(.A(new_n291), .B1(new_n845), .B2(new_n798), .ZN(new_n846));
  AOI21_X1  g660(.A(new_n844), .B1(new_n846), .B2(G210), .ZN(new_n847));
  AOI21_X1  g661(.A(new_n785), .B1(new_n791), .B2(new_n793), .ZN(new_n848));
  INV_X1    g662(.A(G210), .ZN(new_n849));
  NOR4_X1   g663(.A1(new_n848), .A2(KEYINPUT120), .A3(new_n849), .A4(new_n291), .ZN(new_n850));
  OR2_X1    g664(.A1(new_n598), .A2(new_n570), .ZN(new_n851));
  AND2_X1   g665(.A1(new_n851), .A2(new_n571), .ZN(new_n852));
  XOR2_X1   g666(.A(new_n852), .B(KEYINPUT55), .Z(new_n853));
  INV_X1    g667(.A(new_n853), .ZN(new_n854));
  INV_X1    g668(.A(KEYINPUT56), .ZN(new_n855));
  NAND2_X1  g669(.A1(new_n854), .A2(new_n855), .ZN(new_n856));
  NOR3_X1   g670(.A1(new_n847), .A2(new_n850), .A3(new_n856), .ZN(new_n857));
  NOR2_X1   g671(.A1(new_n192), .A2(G952), .ZN(new_n858));
  XNOR2_X1  g672(.A(new_n858), .B(KEYINPUT121), .ZN(new_n859));
  AOI21_X1  g673(.A(KEYINPUT56), .B1(new_n846), .B2(G210), .ZN(new_n860));
  OAI21_X1  g674(.A(new_n859), .B1(new_n860), .B2(new_n854), .ZN(new_n861));
  OAI21_X1  g675(.A(KEYINPUT122), .B1(new_n857), .B2(new_n861), .ZN(new_n862));
  INV_X1    g676(.A(new_n859), .ZN(new_n863));
  OAI21_X1  g677(.A(new_n798), .B1(new_n799), .B2(new_n800), .ZN(new_n864));
  NAND3_X1  g678(.A1(new_n864), .A2(G210), .A3(G902), .ZN(new_n865));
  NAND2_X1  g679(.A1(new_n865), .A2(new_n855), .ZN(new_n866));
  AOI21_X1  g680(.A(new_n863), .B1(new_n866), .B2(new_n853), .ZN(new_n867));
  NAND2_X1  g681(.A1(new_n865), .A2(KEYINPUT120), .ZN(new_n868));
  NAND3_X1  g682(.A1(new_n846), .A2(new_n844), .A3(G210), .ZN(new_n869));
  NAND4_X1  g683(.A1(new_n868), .A2(new_n869), .A3(new_n855), .A4(new_n854), .ZN(new_n870));
  INV_X1    g684(.A(KEYINPUT122), .ZN(new_n871));
  NAND3_X1  g685(.A1(new_n867), .A2(new_n870), .A3(new_n871), .ZN(new_n872));
  NAND2_X1  g686(.A1(new_n862), .A2(new_n872), .ZN(G51));
  NAND2_X1  g687(.A1(new_n864), .A2(KEYINPUT54), .ZN(new_n874));
  NAND2_X1  g688(.A1(new_n874), .A2(new_n801), .ZN(new_n875));
  INV_X1    g689(.A(new_n875), .ZN(new_n876));
  NAND2_X1  g690(.A1(G469), .A2(G902), .ZN(new_n877));
  XNOR2_X1  g691(.A(new_n877), .B(KEYINPUT57), .ZN(new_n878));
  INV_X1    g692(.A(new_n408), .ZN(new_n879));
  INV_X1    g693(.A(new_n405), .ZN(new_n880));
  OAI22_X1  g694(.A1(new_n876), .A2(new_n878), .B1(new_n879), .B2(new_n880), .ZN(new_n881));
  NAND3_X1  g695(.A1(new_n846), .A2(G469), .A3(new_n735), .ZN(new_n882));
  AOI21_X1  g696(.A(new_n858), .B1(new_n881), .B2(new_n882), .ZN(G54));
  INV_X1    g697(.A(new_n858), .ZN(new_n884));
  AND3_X1   g698(.A1(new_n846), .A2(KEYINPUT58), .A3(G475), .ZN(new_n885));
  OAI21_X1  g699(.A(new_n884), .B1(new_n885), .B2(new_n230), .ZN(new_n886));
  AOI21_X1  g700(.A(new_n886), .B1(new_n230), .B2(new_n885), .ZN(G60));
  INV_X1    g701(.A(KEYINPUT123), .ZN(new_n888));
  INV_X1    g702(.A(new_n615), .ZN(new_n889));
  NAND3_X1  g703(.A1(new_n848), .A2(new_n795), .A3(new_n797), .ZN(new_n890));
  INV_X1    g704(.A(new_n784), .ZN(new_n891));
  NAND3_X1  g705(.A1(new_n802), .A2(new_n890), .A3(new_n891), .ZN(new_n892));
  NAND2_X1  g706(.A1(G478), .A2(G902), .ZN(new_n893));
  XOR2_X1   g707(.A(new_n893), .B(KEYINPUT59), .Z(new_n894));
  INV_X1    g708(.A(new_n894), .ZN(new_n895));
  AOI21_X1  g709(.A(new_n889), .B1(new_n892), .B2(new_n895), .ZN(new_n896));
  NOR2_X1   g710(.A1(new_n615), .A2(new_n894), .ZN(new_n897));
  NOR2_X1   g711(.A1(new_n848), .A2(new_n797), .ZN(new_n898));
  OAI21_X1  g712(.A(new_n897), .B1(new_n898), .B2(new_n794), .ZN(new_n899));
  NAND2_X1  g713(.A1(new_n899), .A2(new_n859), .ZN(new_n900));
  OAI21_X1  g714(.A(new_n888), .B1(new_n896), .B2(new_n900), .ZN(new_n901));
  AOI21_X1  g715(.A(new_n863), .B1(new_n875), .B2(new_n897), .ZN(new_n902));
  AOI21_X1  g716(.A(new_n894), .B1(new_n796), .B2(new_n802), .ZN(new_n903));
  OAI211_X1 g717(.A(KEYINPUT123), .B(new_n902), .C1(new_n903), .C2(new_n889), .ZN(new_n904));
  NAND2_X1  g718(.A1(new_n901), .A2(new_n904), .ZN(G63));
  INV_X1    g719(.A(new_n451), .ZN(new_n906));
  NAND2_X1  g720(.A1(G217), .A2(G902), .ZN(new_n907));
  OR2_X1    g721(.A1(new_n907), .A2(KEYINPUT60), .ZN(new_n908));
  NAND2_X1  g722(.A1(new_n907), .A2(KEYINPUT60), .ZN(new_n909));
  NAND2_X1  g723(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  OAI21_X1  g724(.A(new_n906), .B1(new_n848), .B2(new_n910), .ZN(new_n911));
  NAND3_X1  g725(.A1(new_n864), .A2(new_n909), .A3(new_n908), .ZN(new_n912));
  OAI211_X1 g726(.A(new_n859), .B(new_n911), .C1(new_n912), .C2(new_n647), .ZN(new_n913));
  XNOR2_X1  g727(.A(KEYINPUT124), .B(KEYINPUT61), .ZN(new_n914));
  NAND2_X1  g728(.A1(new_n913), .A2(new_n914), .ZN(new_n915));
  INV_X1    g729(.A(KEYINPUT125), .ZN(new_n916));
  NAND2_X1  g730(.A1(new_n915), .A2(new_n916), .ZN(new_n917));
  NAND3_X1  g731(.A1(new_n913), .A2(KEYINPUT125), .A3(new_n914), .ZN(new_n918));
  INV_X1    g732(.A(KEYINPUT61), .ZN(new_n919));
  OR2_X1    g733(.A1(new_n913), .A2(new_n919), .ZN(new_n920));
  NAND3_X1  g734(.A1(new_n917), .A2(new_n918), .A3(new_n920), .ZN(G66));
  OAI21_X1  g735(.A(G953), .B1(new_n249), .B2(new_n568), .ZN(new_n922));
  XNOR2_X1  g736(.A(new_n922), .B(KEYINPUT126), .ZN(new_n923));
  NAND2_X1  g737(.A1(new_n752), .A2(new_n695), .ZN(new_n924));
  INV_X1    g738(.A(new_n699), .ZN(new_n925));
  NOR2_X1   g739(.A1(new_n924), .A2(new_n925), .ZN(new_n926));
  OAI21_X1  g740(.A(new_n923), .B1(new_n926), .B2(G953), .ZN(new_n927));
  INV_X1    g741(.A(G898), .ZN(new_n928));
  AOI21_X1  g742(.A(new_n598), .B1(new_n928), .B2(G953), .ZN(new_n929));
  XOR2_X1   g743(.A(new_n927), .B(new_n929), .Z(G69));
  AND2_X1   g744(.A1(new_n411), .A2(new_n672), .ZN(new_n931));
  NAND4_X1  g745(.A1(new_n931), .A2(new_n530), .A3(new_n712), .A4(new_n749), .ZN(new_n932));
  NAND3_X1  g746(.A1(new_n742), .A2(new_n747), .A3(new_n932), .ZN(new_n933));
  NAND2_X1  g747(.A1(new_n679), .A2(new_n770), .ZN(new_n934));
  XNOR2_X1  g748(.A(new_n934), .B(KEYINPUT62), .ZN(new_n935));
  NOR2_X1   g749(.A1(new_n933), .A2(new_n935), .ZN(new_n936));
  NAND2_X1  g750(.A1(new_n936), .A2(new_n192), .ZN(new_n937));
  NAND3_X1  g751(.A1(G227), .A2(G900), .A3(G953), .ZN(new_n938));
  XNOR2_X1  g752(.A(new_n515), .B(new_n221), .ZN(new_n939));
  INV_X1    g753(.A(new_n939), .ZN(new_n940));
  NAND3_X1  g754(.A1(new_n937), .A2(new_n938), .A3(new_n940), .ZN(new_n941));
  NAND4_X1  g755(.A1(new_n740), .A2(new_n605), .A3(new_n669), .A4(new_n714), .ZN(new_n942));
  AND3_X1   g756(.A1(new_n747), .A2(new_n770), .A3(new_n942), .ZN(new_n943));
  NAND4_X1  g757(.A1(new_n742), .A2(new_n719), .A3(new_n721), .A4(new_n943), .ZN(new_n944));
  NAND2_X1  g758(.A1(new_n944), .A2(new_n192), .ZN(new_n945));
  NAND3_X1  g759(.A1(new_n377), .A2(G900), .A3(G953), .ZN(new_n946));
  NAND3_X1  g760(.A1(new_n945), .A2(new_n939), .A3(new_n946), .ZN(new_n947));
  NAND2_X1  g761(.A1(new_n941), .A2(new_n947), .ZN(G72));
  NAND2_X1  g762(.A1(G472), .A2(G902), .ZN(new_n949));
  XOR2_X1   g763(.A(new_n949), .B(KEYINPUT63), .Z(new_n950));
  INV_X1    g764(.A(new_n926), .ZN(new_n951));
  OAI21_X1  g765(.A(new_n950), .B1(new_n944), .B2(new_n951), .ZN(new_n952));
  NAND4_X1  g766(.A1(new_n952), .A2(new_n466), .A3(new_n488), .A4(new_n516), .ZN(new_n953));
  INV_X1    g767(.A(new_n950), .ZN(new_n954));
  AOI21_X1  g768(.A(new_n954), .B1(new_n936), .B2(new_n926), .ZN(new_n955));
  OAI21_X1  g769(.A(new_n465), .B1(new_n487), .B2(new_n489), .ZN(new_n956));
  OAI211_X1 g770(.A(new_n953), .B(new_n884), .C1(new_n955), .C2(new_n956), .ZN(new_n957));
  AND2_X1   g771(.A1(new_n779), .A2(new_n783), .ZN(new_n958));
  INV_X1    g772(.A(new_n664), .ZN(new_n959));
  AOI21_X1  g773(.A(new_n954), .B1(new_n959), .B2(new_n490), .ZN(new_n960));
  AOI21_X1  g774(.A(new_n957), .B1(new_n958), .B2(new_n960), .ZN(G57));
endmodule


