//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 1 1 0 1 1 0 1 0 0 1 1 0 1 0 0 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 1 1 1 1 1 1 1 1 0 1 1 0 1 0 1 0 0 1 0 0 1 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:28:48 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n446, new_n448, new_n452, new_n453, new_n454, new_n455,
    new_n456, new_n459, new_n460, new_n461, new_n462, new_n463, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n531, new_n532,
    new_n533, new_n534, new_n535, new_n536, new_n537, new_n538, new_n539,
    new_n540, new_n541, new_n542, new_n545, new_n546, new_n547, new_n548,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n560, new_n561, new_n562, new_n564, new_n565, new_n566, new_n567,
    new_n568, new_n569, new_n570, new_n571, new_n572, new_n573, new_n574,
    new_n575, new_n576, new_n577, new_n578, new_n579, new_n580, new_n581,
    new_n584, new_n585, new_n586, new_n588, new_n589, new_n590, new_n591,
    new_n592, new_n593, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n615, new_n618,
    new_n619, new_n621, new_n622, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n832, new_n833, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1195, new_n1196,
    new_n1198, new_n1199;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  XOR2_X1   g006(.A(KEYINPUT64), .B(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(new_n436));
  XNOR2_X1  g011(.A(new_n436), .B(KEYINPUT65), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  INV_X1    g015(.A(G57), .ZN(G237));
  XOR2_X1   g016(.A(KEYINPUT66), .B(G108), .Z(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  NAND2_X1  g020(.A1(G94), .A2(G452), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT67), .Z(G173));
  NAND2_X1  g022(.A1(G7), .A2(G661), .ZN(new_n448));
  XOR2_X1   g023(.A(new_n448), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g024(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g025(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  OR4_X1    g026(.A1(G218), .A2(G220), .A3(G221), .A4(G219), .ZN(new_n452));
  XOR2_X1   g027(.A(new_n452), .B(KEYINPUT2), .Z(new_n453));
  NOR4_X1   g028(.A1(G238), .A2(G237), .A3(G235), .A4(G236), .ZN(new_n454));
  XOR2_X1   g029(.A(new_n454), .B(KEYINPUT68), .Z(new_n455));
  NAND2_X1  g030(.A1(new_n453), .A2(new_n455), .ZN(new_n456));
  INV_X1    g031(.A(new_n456), .ZN(G325));
  XNOR2_X1  g032(.A(new_n456), .B(KEYINPUT69), .ZN(G261));
  INV_X1    g033(.A(new_n453), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n459), .A2(G2106), .ZN(new_n460));
  INV_X1    g035(.A(G567), .ZN(new_n461));
  OR2_X1    g036(.A1(new_n455), .A2(new_n461), .ZN(new_n462));
  NAND2_X1  g037(.A1(new_n460), .A2(new_n462), .ZN(new_n463));
  INV_X1    g038(.A(new_n463), .ZN(G319));
  INV_X1    g039(.A(G2105), .ZN(new_n465));
  NAND3_X1  g040(.A1(new_n465), .A2(G101), .A3(G2104), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n466), .A2(KEYINPUT70), .ZN(new_n467));
  INV_X1    g042(.A(KEYINPUT70), .ZN(new_n468));
  NAND4_X1  g043(.A1(new_n468), .A2(new_n465), .A3(G101), .A4(G2104), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n467), .A2(new_n469), .ZN(new_n470));
  AND2_X1   g045(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n471));
  NOR2_X1   g046(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n472));
  OAI211_X1 g047(.A(G137), .B(new_n465), .C1(new_n471), .C2(new_n472), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n470), .A2(new_n473), .ZN(new_n474));
  OAI21_X1  g049(.A(G125), .B1(new_n471), .B2(new_n472), .ZN(new_n475));
  NAND2_X1  g050(.A1(G113), .A2(G2104), .ZN(new_n476));
  AOI21_X1  g051(.A(new_n465), .B1(new_n475), .B2(new_n476), .ZN(new_n477));
  NOR2_X1   g052(.A1(new_n474), .A2(new_n477), .ZN(G160));
  INV_X1    g053(.A(KEYINPUT3), .ZN(new_n479));
  INV_X1    g054(.A(G2104), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n479), .A2(new_n480), .ZN(new_n481));
  NAND2_X1  g056(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n482));
  AOI21_X1  g057(.A(G2105), .B1(new_n481), .B2(new_n482), .ZN(new_n483));
  NAND2_X1  g058(.A1(new_n483), .A2(G136), .ZN(new_n484));
  NOR2_X1   g059(.A1(new_n465), .A2(G112), .ZN(new_n485));
  OAI21_X1  g060(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n486));
  OAI21_X1  g061(.A(new_n484), .B1(new_n485), .B2(new_n486), .ZN(new_n487));
  NAND2_X1  g062(.A1(new_n481), .A2(new_n482), .ZN(new_n488));
  INV_X1    g063(.A(KEYINPUT71), .ZN(new_n489));
  NAND3_X1  g064(.A1(new_n488), .A2(new_n489), .A3(G2105), .ZN(new_n490));
  INV_X1    g065(.A(new_n490), .ZN(new_n491));
  AOI21_X1  g066(.A(new_n489), .B1(new_n488), .B2(G2105), .ZN(new_n492));
  NOR2_X1   g067(.A1(new_n491), .A2(new_n492), .ZN(new_n493));
  INV_X1    g068(.A(new_n493), .ZN(new_n494));
  AOI21_X1  g069(.A(new_n487), .B1(new_n494), .B2(G124), .ZN(G162));
  OAI211_X1 g070(.A(G138), .B(new_n465), .C1(new_n471), .C2(new_n472), .ZN(new_n496));
  INV_X1    g071(.A(KEYINPUT4), .ZN(new_n497));
  NOR2_X1   g072(.A1(new_n497), .A2(KEYINPUT73), .ZN(new_n498));
  INV_X1    g073(.A(new_n498), .ZN(new_n499));
  NAND2_X1  g074(.A1(new_n496), .A2(new_n499), .ZN(new_n500));
  INV_X1    g075(.A(KEYINPUT73), .ZN(new_n501));
  NAND4_X1  g076(.A1(new_n501), .A2(new_n465), .A3(KEYINPUT4), .A4(G138), .ZN(new_n502));
  NAND2_X1  g077(.A1(G126), .A2(G2105), .ZN(new_n503));
  NAND2_X1  g078(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  NAND2_X1  g079(.A1(new_n504), .A2(new_n488), .ZN(new_n505));
  OR2_X1    g080(.A1(G102), .A2(G2105), .ZN(new_n506));
  OAI21_X1  g081(.A(G2105), .B1(KEYINPUT72), .B2(G114), .ZN(new_n507));
  AND2_X1   g082(.A1(KEYINPUT72), .A2(G114), .ZN(new_n508));
  OAI211_X1 g083(.A(G2104), .B(new_n506), .C1(new_n507), .C2(new_n508), .ZN(new_n509));
  NAND3_X1  g084(.A1(new_n500), .A2(new_n505), .A3(new_n509), .ZN(new_n510));
  INV_X1    g085(.A(new_n510), .ZN(G164));
  INV_X1    g086(.A(KEYINPUT5), .ZN(new_n512));
  INV_X1    g087(.A(G543), .ZN(new_n513));
  OAI21_X1  g088(.A(new_n512), .B1(new_n513), .B2(KEYINPUT74), .ZN(new_n514));
  INV_X1    g089(.A(KEYINPUT74), .ZN(new_n515));
  NAND3_X1  g090(.A1(new_n515), .A2(KEYINPUT5), .A3(G543), .ZN(new_n516));
  NAND2_X1  g091(.A1(new_n514), .A2(new_n516), .ZN(new_n517));
  AOI22_X1  g092(.A1(new_n517), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n518));
  INV_X1    g093(.A(G651), .ZN(new_n519));
  NOR2_X1   g094(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  INV_X1    g095(.A(KEYINPUT6), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n521), .A2(new_n519), .ZN(new_n522));
  NAND2_X1  g097(.A1(KEYINPUT6), .A2(G651), .ZN(new_n523));
  AOI21_X1  g098(.A(new_n513), .B1(new_n522), .B2(new_n523), .ZN(new_n524));
  NAND2_X1  g099(.A1(new_n524), .A2(G50), .ZN(new_n525));
  NAND2_X1  g100(.A1(new_n522), .A2(new_n523), .ZN(new_n526));
  NAND2_X1  g101(.A1(new_n517), .A2(new_n526), .ZN(new_n527));
  INV_X1    g102(.A(G88), .ZN(new_n528));
  OAI21_X1  g103(.A(new_n525), .B1(new_n527), .B2(new_n528), .ZN(new_n529));
  NOR2_X1   g104(.A1(new_n520), .A2(new_n529), .ZN(G166));
  NAND3_X1  g105(.A1(new_n517), .A2(G63), .A3(G651), .ZN(new_n531));
  INV_X1    g106(.A(new_n524), .ZN(new_n532));
  INV_X1    g107(.A(G51), .ZN(new_n533));
  OAI21_X1  g108(.A(new_n531), .B1(new_n532), .B2(new_n533), .ZN(new_n534));
  NAND2_X1  g109(.A1(new_n534), .A2(KEYINPUT75), .ZN(new_n535));
  INV_X1    g110(.A(KEYINPUT75), .ZN(new_n536));
  OAI211_X1 g111(.A(new_n531), .B(new_n536), .C1(new_n533), .C2(new_n532), .ZN(new_n537));
  AOI22_X1  g112(.A1(new_n514), .A2(new_n516), .B1(new_n522), .B2(new_n523), .ZN(new_n538));
  NAND3_X1  g113(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n539));
  NAND2_X1  g114(.A1(new_n539), .A2(KEYINPUT7), .ZN(new_n540));
  OR2_X1    g115(.A1(new_n539), .A2(KEYINPUT7), .ZN(new_n541));
  AOI22_X1  g116(.A1(new_n538), .A2(G89), .B1(new_n540), .B2(new_n541), .ZN(new_n542));
  NAND3_X1  g117(.A1(new_n535), .A2(new_n537), .A3(new_n542), .ZN(G286));
  INV_X1    g118(.A(G286), .ZN(G168));
  AOI22_X1  g119(.A1(new_n538), .A2(G90), .B1(new_n524), .B2(G52), .ZN(new_n545));
  XNOR2_X1  g120(.A(new_n545), .B(KEYINPUT76), .ZN(new_n546));
  AOI22_X1  g121(.A1(new_n517), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n547));
  OR2_X1    g122(.A1(new_n547), .A2(new_n519), .ZN(new_n548));
  NAND2_X1  g123(.A1(new_n546), .A2(new_n548), .ZN(G301));
  INV_X1    g124(.A(G301), .ZN(G171));
  AOI22_X1  g125(.A1(new_n517), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n551));
  NOR2_X1   g126(.A1(new_n551), .A2(new_n519), .ZN(new_n552));
  NAND2_X1  g127(.A1(new_n524), .A2(G43), .ZN(new_n553));
  XNOR2_X1  g128(.A(KEYINPUT77), .B(G81), .ZN(new_n554));
  OAI21_X1  g129(.A(new_n553), .B1(new_n527), .B2(new_n554), .ZN(new_n555));
  NOR2_X1   g130(.A1(new_n552), .A2(new_n555), .ZN(new_n556));
  NAND2_X1  g131(.A1(new_n556), .A2(G860), .ZN(new_n557));
  XNOR2_X1  g132(.A(new_n557), .B(KEYINPUT78), .ZN(G153));
  NAND4_X1  g133(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g134(.A1(G1), .A2(G3), .ZN(new_n560));
  XNOR2_X1  g135(.A(new_n560), .B(KEYINPUT8), .ZN(new_n561));
  NAND4_X1  g136(.A1(G319), .A2(G483), .A3(G661), .A4(new_n561), .ZN(new_n562));
  XOR2_X1   g137(.A(new_n562), .B(KEYINPUT79), .Z(G188));
  INV_X1    g138(.A(KEYINPUT81), .ZN(new_n564));
  INV_X1    g139(.A(G91), .ZN(new_n565));
  OAI21_X1  g140(.A(new_n564), .B1(new_n527), .B2(new_n565), .ZN(new_n566));
  NAND3_X1  g141(.A1(new_n538), .A2(KEYINPUT81), .A3(G91), .ZN(new_n567));
  NAND2_X1  g142(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  INV_X1    g143(.A(new_n568), .ZN(new_n569));
  NAND3_X1  g144(.A1(new_n526), .A2(G53), .A3(G543), .ZN(new_n570));
  XOR2_X1   g145(.A(KEYINPUT80), .B(KEYINPUT9), .Z(new_n571));
  NAND2_X1  g146(.A1(new_n570), .A2(new_n571), .ZN(new_n572));
  INV_X1    g147(.A(KEYINPUT9), .ZN(new_n573));
  OAI211_X1 g148(.A(new_n524), .B(G53), .C1(KEYINPUT80), .C2(new_n573), .ZN(new_n574));
  NAND2_X1  g149(.A1(new_n572), .A2(new_n574), .ZN(new_n575));
  INV_X1    g150(.A(G65), .ZN(new_n576));
  AOI21_X1  g151(.A(new_n576), .B1(new_n514), .B2(new_n516), .ZN(new_n577));
  AND2_X1   g152(.A1(G78), .A2(G543), .ZN(new_n578));
  OAI21_X1  g153(.A(G651), .B1(new_n577), .B2(new_n578), .ZN(new_n579));
  NAND2_X1  g154(.A1(new_n575), .A2(new_n579), .ZN(new_n580));
  NOR2_X1   g155(.A1(new_n569), .A2(new_n580), .ZN(new_n581));
  INV_X1    g156(.A(new_n581), .ZN(G299));
  INV_X1    g157(.A(G166), .ZN(G303));
  OAI21_X1  g158(.A(G651), .B1(new_n517), .B2(G74), .ZN(new_n584));
  NAND3_X1  g159(.A1(new_n517), .A2(G87), .A3(new_n526), .ZN(new_n585));
  NAND2_X1  g160(.A1(new_n524), .A2(G49), .ZN(new_n586));
  NAND3_X1  g161(.A1(new_n584), .A2(new_n585), .A3(new_n586), .ZN(G288));
  AOI22_X1  g162(.A1(new_n538), .A2(G86), .B1(new_n524), .B2(G48), .ZN(new_n588));
  INV_X1    g163(.A(G61), .ZN(new_n589));
  AOI21_X1  g164(.A(new_n589), .B1(new_n514), .B2(new_n516), .ZN(new_n590));
  NAND2_X1  g165(.A1(G73), .A2(G543), .ZN(new_n591));
  INV_X1    g166(.A(new_n591), .ZN(new_n592));
  OAI21_X1  g167(.A(G651), .B1(new_n590), .B2(new_n592), .ZN(new_n593));
  NAND2_X1  g168(.A1(new_n588), .A2(new_n593), .ZN(G305));
  NAND2_X1  g169(.A1(new_n517), .A2(G60), .ZN(new_n595));
  INV_X1    g170(.A(G72), .ZN(new_n596));
  OAI21_X1  g171(.A(new_n595), .B1(new_n596), .B2(new_n513), .ZN(new_n597));
  INV_X1    g172(.A(KEYINPUT82), .ZN(new_n598));
  AOI21_X1  g173(.A(new_n519), .B1(new_n597), .B2(new_n598), .ZN(new_n599));
  OAI21_X1  g174(.A(new_n599), .B1(new_n598), .B2(new_n597), .ZN(new_n600));
  AOI22_X1  g175(.A1(new_n538), .A2(G85), .B1(new_n524), .B2(G47), .ZN(new_n601));
  NAND2_X1  g176(.A1(new_n600), .A2(new_n601), .ZN(G290));
  AOI22_X1  g177(.A1(new_n517), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n603));
  AOI21_X1  g178(.A(new_n519), .B1(new_n603), .B2(KEYINPUT83), .ZN(new_n604));
  OAI21_X1  g179(.A(new_n604), .B1(KEYINPUT83), .B2(new_n603), .ZN(new_n605));
  NAND2_X1  g180(.A1(new_n524), .A2(G54), .ZN(new_n606));
  NAND2_X1  g181(.A1(new_n538), .A2(G92), .ZN(new_n607));
  INV_X1    g182(.A(KEYINPUT10), .ZN(new_n608));
  XNOR2_X1  g183(.A(new_n607), .B(new_n608), .ZN(new_n609));
  NAND3_X1  g184(.A1(new_n605), .A2(new_n606), .A3(new_n609), .ZN(new_n610));
  INV_X1    g185(.A(G868), .ZN(new_n611));
  NAND2_X1  g186(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  OAI21_X1  g187(.A(new_n612), .B1(G171), .B2(new_n611), .ZN(G284));
  OAI21_X1  g188(.A(new_n612), .B1(G171), .B2(new_n611), .ZN(G321));
  NAND2_X1  g189(.A1(G286), .A2(G868), .ZN(new_n615));
  OAI21_X1  g190(.A(new_n615), .B1(new_n581), .B2(G868), .ZN(G280));
  XOR2_X1   g191(.A(G280), .B(KEYINPUT84), .Z(G297));
  INV_X1    g192(.A(new_n610), .ZN(new_n618));
  INV_X1    g193(.A(G559), .ZN(new_n619));
  OAI21_X1  g194(.A(new_n618), .B1(new_n619), .B2(G860), .ZN(G148));
  OAI21_X1  g195(.A(new_n611), .B1(new_n552), .B2(new_n555), .ZN(new_n621));
  NOR2_X1   g196(.A1(new_n610), .A2(G559), .ZN(new_n622));
  OAI21_X1  g197(.A(new_n621), .B1(new_n622), .B2(new_n611), .ZN(G323));
  XNOR2_X1  g198(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NOR2_X1   g199(.A1(new_n480), .A2(G2105), .ZN(new_n625));
  NAND2_X1  g200(.A1(new_n488), .A2(new_n625), .ZN(new_n626));
  XNOR2_X1  g201(.A(new_n626), .B(KEYINPUT12), .ZN(new_n627));
  XNOR2_X1  g202(.A(new_n627), .B(KEYINPUT13), .ZN(new_n628));
  INV_X1    g203(.A(new_n628), .ZN(new_n629));
  OR2_X1    g204(.A1(new_n629), .A2(G2100), .ZN(new_n630));
  OAI21_X1  g205(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n631));
  INV_X1    g206(.A(G111), .ZN(new_n632));
  AOI21_X1  g207(.A(new_n631), .B1(new_n632), .B2(G2105), .ZN(new_n633));
  AOI21_X1  g208(.A(new_n633), .B1(G135), .B2(new_n483), .ZN(new_n634));
  INV_X1    g209(.A(new_n634), .ZN(new_n635));
  AOI21_X1  g210(.A(new_n635), .B1(new_n494), .B2(G123), .ZN(new_n636));
  INV_X1    g211(.A(new_n636), .ZN(new_n637));
  OR2_X1    g212(.A1(new_n637), .A2(G2096), .ZN(new_n638));
  NAND2_X1  g213(.A1(new_n629), .A2(G2100), .ZN(new_n639));
  NAND2_X1  g214(.A1(new_n637), .A2(G2096), .ZN(new_n640));
  NAND4_X1  g215(.A1(new_n630), .A2(new_n638), .A3(new_n639), .A4(new_n640), .ZN(G156));
  XNOR2_X1  g216(.A(G2427), .B(G2438), .ZN(new_n642));
  XNOR2_X1  g217(.A(new_n642), .B(G2430), .ZN(new_n643));
  XNOR2_X1  g218(.A(KEYINPUT15), .B(G2435), .ZN(new_n644));
  OR2_X1    g219(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  NAND2_X1  g220(.A1(new_n643), .A2(new_n644), .ZN(new_n646));
  NAND3_X1  g221(.A1(new_n645), .A2(KEYINPUT14), .A3(new_n646), .ZN(new_n647));
  XOR2_X1   g222(.A(G1341), .B(G1348), .Z(new_n648));
  XNOR2_X1  g223(.A(KEYINPUT85), .B(KEYINPUT16), .ZN(new_n649));
  XNOR2_X1  g224(.A(new_n648), .B(new_n649), .ZN(new_n650));
  XNOR2_X1  g225(.A(new_n647), .B(new_n650), .ZN(new_n651));
  XOR2_X1   g226(.A(G2451), .B(G2454), .Z(new_n652));
  XNOR2_X1  g227(.A(G2443), .B(G2446), .ZN(new_n653));
  XNOR2_X1  g228(.A(new_n652), .B(new_n653), .ZN(new_n654));
  OR2_X1    g229(.A1(new_n651), .A2(new_n654), .ZN(new_n655));
  NAND2_X1  g230(.A1(new_n651), .A2(new_n654), .ZN(new_n656));
  NAND3_X1  g231(.A1(new_n655), .A2(G14), .A3(new_n656), .ZN(new_n657));
  XOR2_X1   g232(.A(new_n657), .B(KEYINPUT86), .Z(G401));
  XOR2_X1   g233(.A(G2084), .B(G2090), .Z(new_n659));
  INV_X1    g234(.A(new_n659), .ZN(new_n660));
  XNOR2_X1  g235(.A(G2067), .B(G2678), .ZN(new_n661));
  XNOR2_X1  g236(.A(G2072), .B(G2078), .ZN(new_n662));
  OAI21_X1  g237(.A(new_n660), .B1(new_n661), .B2(new_n662), .ZN(new_n663));
  XOR2_X1   g238(.A(new_n662), .B(KEYINPUT17), .Z(new_n664));
  INV_X1    g239(.A(new_n664), .ZN(new_n665));
  AOI21_X1  g240(.A(new_n663), .B1(new_n665), .B2(new_n661), .ZN(new_n666));
  XNOR2_X1  g241(.A(new_n666), .B(KEYINPUT87), .ZN(new_n667));
  NAND3_X1  g242(.A1(new_n659), .A2(new_n661), .A3(new_n662), .ZN(new_n668));
  XOR2_X1   g243(.A(new_n668), .B(KEYINPUT18), .Z(new_n669));
  OR2_X1    g244(.A1(new_n660), .A2(new_n661), .ZN(new_n670));
  OAI211_X1 g245(.A(new_n667), .B(new_n669), .C1(new_n665), .C2(new_n670), .ZN(new_n671));
  XOR2_X1   g246(.A(G2096), .B(G2100), .Z(new_n672));
  XNOR2_X1  g247(.A(new_n671), .B(new_n672), .ZN(G227));
  XNOR2_X1  g248(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n674));
  XNOR2_X1  g249(.A(new_n674), .B(KEYINPUT91), .ZN(new_n675));
  INV_X1    g250(.A(new_n675), .ZN(new_n676));
  XNOR2_X1  g251(.A(G1961), .B(G1966), .ZN(new_n677));
  XNOR2_X1  g252(.A(new_n677), .B(KEYINPUT88), .ZN(new_n678));
  XNOR2_X1  g253(.A(G1971), .B(G1976), .ZN(new_n679));
  XNOR2_X1  g254(.A(new_n679), .B(KEYINPUT19), .ZN(new_n680));
  XOR2_X1   g255(.A(G1956), .B(G2474), .Z(new_n681));
  NAND3_X1  g256(.A1(new_n678), .A2(new_n680), .A3(new_n681), .ZN(new_n682));
  OAI21_X1  g257(.A(new_n682), .B1(new_n678), .B2(new_n681), .ZN(new_n683));
  INV_X1    g258(.A(KEYINPUT90), .ZN(new_n684));
  NAND2_X1  g259(.A1(new_n680), .A2(new_n684), .ZN(new_n685));
  XOR2_X1   g260(.A(new_n683), .B(new_n685), .Z(new_n686));
  NAND2_X1  g261(.A1(new_n678), .A2(new_n681), .ZN(new_n687));
  NOR2_X1   g262(.A1(new_n687), .A2(new_n680), .ZN(new_n688));
  XNOR2_X1  g263(.A(KEYINPUT89), .B(KEYINPUT20), .ZN(new_n689));
  XNOR2_X1  g264(.A(new_n688), .B(new_n689), .ZN(new_n690));
  NAND2_X1  g265(.A1(new_n686), .A2(new_n690), .ZN(new_n691));
  INV_X1    g266(.A(G1981), .ZN(new_n692));
  XNOR2_X1  g267(.A(new_n691), .B(new_n692), .ZN(new_n693));
  OR2_X1    g268(.A1(new_n693), .A2(G1986), .ZN(new_n694));
  NAND2_X1  g269(.A1(new_n693), .A2(G1986), .ZN(new_n695));
  AOI21_X1  g270(.A(new_n676), .B1(new_n694), .B2(new_n695), .ZN(new_n696));
  INV_X1    g271(.A(new_n696), .ZN(new_n697));
  XNOR2_X1  g272(.A(G1991), .B(G1996), .ZN(new_n698));
  NAND3_X1  g273(.A1(new_n694), .A2(new_n676), .A3(new_n695), .ZN(new_n699));
  NAND3_X1  g274(.A1(new_n697), .A2(new_n698), .A3(new_n699), .ZN(new_n700));
  INV_X1    g275(.A(new_n698), .ZN(new_n701));
  AND3_X1   g276(.A1(new_n694), .A2(new_n676), .A3(new_n695), .ZN(new_n702));
  OAI21_X1  g277(.A(new_n701), .B1(new_n702), .B2(new_n696), .ZN(new_n703));
  NAND2_X1  g278(.A1(new_n700), .A2(new_n703), .ZN(G229));
  NAND2_X1  g279(.A1(G171), .A2(G16), .ZN(new_n705));
  OAI21_X1  g280(.A(new_n705), .B1(G5), .B2(G16), .ZN(new_n706));
  INV_X1    g281(.A(G1961), .ZN(new_n707));
  OR2_X1    g282(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  NAND2_X1  g283(.A1(new_n706), .A2(new_n707), .ZN(new_n709));
  XNOR2_X1  g284(.A(KEYINPUT27), .B(G1996), .ZN(new_n710));
  XNOR2_X1  g285(.A(KEYINPUT97), .B(KEYINPUT26), .ZN(new_n711));
  NAND3_X1  g286(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n712));
  XNOR2_X1  g287(.A(new_n711), .B(new_n712), .ZN(new_n713));
  AOI21_X1  g288(.A(new_n713), .B1(G105), .B2(new_n625), .ZN(new_n714));
  INV_X1    g289(.A(G141), .ZN(new_n715));
  INV_X1    g290(.A(new_n483), .ZN(new_n716));
  OAI21_X1  g291(.A(new_n714), .B1(new_n715), .B2(new_n716), .ZN(new_n717));
  AND2_X1   g292(.A1(new_n494), .A2(G129), .ZN(new_n718));
  OAI21_X1  g293(.A(G29), .B1(new_n717), .B2(new_n718), .ZN(new_n719));
  INV_X1    g294(.A(KEYINPUT98), .ZN(new_n720));
  INV_X1    g295(.A(G29), .ZN(new_n721));
  NAND2_X1  g296(.A1(new_n721), .A2(G32), .ZN(new_n722));
  AND3_X1   g297(.A1(new_n719), .A2(new_n720), .A3(new_n722), .ZN(new_n723));
  AOI21_X1  g298(.A(new_n720), .B1(new_n719), .B2(new_n722), .ZN(new_n724));
  OAI21_X1  g299(.A(new_n710), .B1(new_n723), .B2(new_n724), .ZN(new_n725));
  AND3_X1   g300(.A1(new_n708), .A2(new_n709), .A3(new_n725), .ZN(new_n726));
  INV_X1    g301(.A(G16), .ZN(new_n727));
  NAND2_X1  g302(.A1(new_n727), .A2(G21), .ZN(new_n728));
  OAI21_X1  g303(.A(new_n728), .B1(G168), .B2(new_n727), .ZN(new_n729));
  NOR2_X1   g304(.A1(new_n729), .A2(G1966), .ZN(new_n730));
  NAND2_X1  g305(.A1(new_n729), .A2(G1966), .ZN(new_n731));
  NAND2_X1  g306(.A1(new_n721), .A2(G27), .ZN(new_n732));
  OAI21_X1  g307(.A(new_n732), .B1(G164), .B2(new_n721), .ZN(new_n733));
  XOR2_X1   g308(.A(new_n733), .B(KEYINPUT99), .Z(new_n734));
  OAI21_X1  g309(.A(new_n731), .B1(new_n734), .B2(G2078), .ZN(new_n735));
  AOI211_X1 g310(.A(new_n730), .B(new_n735), .C1(G2078), .C2(new_n734), .ZN(new_n736));
  NOR3_X1   g311(.A1(new_n723), .A2(new_n724), .A3(new_n710), .ZN(new_n737));
  XNOR2_X1  g312(.A(KEYINPUT30), .B(G28), .ZN(new_n738));
  OR2_X1    g313(.A1(KEYINPUT31), .A2(G11), .ZN(new_n739));
  NAND2_X1  g314(.A1(KEYINPUT31), .A2(G11), .ZN(new_n740));
  AOI22_X1  g315(.A1(new_n738), .A2(new_n721), .B1(new_n739), .B2(new_n740), .ZN(new_n741));
  NAND2_X1  g316(.A1(new_n721), .A2(G33), .ZN(new_n742));
  NAND3_X1  g317(.A1(new_n465), .A2(G103), .A3(G2104), .ZN(new_n743));
  XNOR2_X1  g318(.A(new_n743), .B(KEYINPUT25), .ZN(new_n744));
  NAND2_X1  g319(.A1(new_n488), .A2(G127), .ZN(new_n745));
  NAND2_X1  g320(.A1(G115), .A2(G2104), .ZN(new_n746));
  AOI21_X1  g321(.A(new_n465), .B1(new_n745), .B2(new_n746), .ZN(new_n747));
  AOI211_X1 g322(.A(new_n744), .B(new_n747), .C1(G139), .C2(new_n483), .ZN(new_n748));
  OAI21_X1  g323(.A(new_n742), .B1(new_n748), .B2(new_n721), .ZN(new_n749));
  OAI221_X1 g324(.A(new_n741), .B1(new_n637), .B2(new_n721), .C1(new_n749), .C2(G2072), .ZN(new_n750));
  NAND2_X1  g325(.A1(G160), .A2(G29), .ZN(new_n751));
  INV_X1    g326(.A(G34), .ZN(new_n752));
  AOI21_X1  g327(.A(G29), .B1(new_n752), .B2(KEYINPUT24), .ZN(new_n753));
  OAI21_X1  g328(.A(new_n753), .B1(KEYINPUT24), .B2(new_n752), .ZN(new_n754));
  AOI21_X1  g329(.A(G2084), .B1(new_n751), .B2(new_n754), .ZN(new_n755));
  AOI21_X1  g330(.A(new_n755), .B1(new_n749), .B2(G2072), .ZN(new_n756));
  NAND3_X1  g331(.A1(new_n751), .A2(G2084), .A3(new_n754), .ZN(new_n757));
  NAND2_X1  g332(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  NOR3_X1   g333(.A1(new_n737), .A2(new_n750), .A3(new_n758), .ZN(new_n759));
  NAND3_X1  g334(.A1(new_n726), .A2(new_n736), .A3(new_n759), .ZN(new_n760));
  AND2_X1   g335(.A1(new_n760), .A2(KEYINPUT100), .ZN(new_n761));
  NOR2_X1   g336(.A1(new_n760), .A2(KEYINPUT100), .ZN(new_n762));
  NAND2_X1  g337(.A1(new_n721), .A2(G35), .ZN(new_n763));
  OAI21_X1  g338(.A(new_n763), .B1(G162), .B2(new_n721), .ZN(new_n764));
  XNOR2_X1  g339(.A(new_n764), .B(KEYINPUT29), .ZN(new_n765));
  NOR2_X1   g340(.A1(new_n765), .A2(G2090), .ZN(new_n766));
  XNOR2_X1  g341(.A(new_n766), .B(KEYINPUT101), .ZN(new_n767));
  NAND2_X1  g342(.A1(new_n727), .A2(G19), .ZN(new_n768));
  OAI21_X1  g343(.A(new_n768), .B1(new_n556), .B2(new_n727), .ZN(new_n769));
  XNOR2_X1  g344(.A(new_n769), .B(G1341), .ZN(new_n770));
  NAND2_X1  g345(.A1(new_n721), .A2(G26), .ZN(new_n771));
  XNOR2_X1  g346(.A(new_n771), .B(KEYINPUT28), .ZN(new_n772));
  NAND2_X1  g347(.A1(new_n483), .A2(G140), .ZN(new_n773));
  NOR2_X1   g348(.A1(new_n465), .A2(G116), .ZN(new_n774));
  OAI21_X1  g349(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n775));
  OAI21_X1  g350(.A(new_n773), .B1(new_n774), .B2(new_n775), .ZN(new_n776));
  AOI21_X1  g351(.A(new_n776), .B1(new_n494), .B2(G128), .ZN(new_n777));
  OAI21_X1  g352(.A(new_n772), .B1(new_n777), .B2(new_n721), .ZN(new_n778));
  XNOR2_X1  g353(.A(new_n778), .B(G2067), .ZN(new_n779));
  AOI211_X1 g354(.A(new_n770), .B(new_n779), .C1(G2090), .C2(new_n765), .ZN(new_n780));
  NAND2_X1  g355(.A1(new_n618), .A2(G16), .ZN(new_n781));
  OAI21_X1  g356(.A(new_n781), .B1(G4), .B2(G16), .ZN(new_n782));
  INV_X1    g357(.A(G1348), .ZN(new_n783));
  OR2_X1    g358(.A1(new_n782), .A2(new_n783), .ZN(new_n784));
  NAND2_X1  g359(.A1(new_n727), .A2(G20), .ZN(new_n785));
  XNOR2_X1  g360(.A(new_n785), .B(KEYINPUT102), .ZN(new_n786));
  XNOR2_X1  g361(.A(new_n786), .B(KEYINPUT23), .ZN(new_n787));
  OAI21_X1  g362(.A(new_n787), .B1(new_n581), .B2(new_n727), .ZN(new_n788));
  XNOR2_X1  g363(.A(new_n788), .B(G1956), .ZN(new_n789));
  AOI21_X1  g364(.A(new_n789), .B1(new_n782), .B2(new_n783), .ZN(new_n790));
  NAND4_X1  g365(.A1(new_n767), .A2(new_n780), .A3(new_n784), .A4(new_n790), .ZN(new_n791));
  NOR3_X1   g366(.A1(new_n761), .A2(new_n762), .A3(new_n791), .ZN(new_n792));
  NAND2_X1  g367(.A1(new_n727), .A2(G23), .ZN(new_n793));
  INV_X1    g368(.A(G288), .ZN(new_n794));
  OAI21_X1  g369(.A(new_n793), .B1(new_n794), .B2(new_n727), .ZN(new_n795));
  XNOR2_X1  g370(.A(new_n795), .B(KEYINPUT33), .ZN(new_n796));
  XNOR2_X1  g371(.A(new_n796), .B(G1976), .ZN(new_n797));
  MUX2_X1   g372(.A(G6), .B(G305), .S(G16), .Z(new_n798));
  XOR2_X1   g373(.A(KEYINPUT32), .B(G1981), .Z(new_n799));
  XNOR2_X1  g374(.A(new_n799), .B(KEYINPUT93), .ZN(new_n800));
  XNOR2_X1  g375(.A(new_n798), .B(new_n800), .ZN(new_n801));
  NAND2_X1  g376(.A1(new_n727), .A2(G22), .ZN(new_n802));
  XNOR2_X1  g377(.A(new_n802), .B(KEYINPUT94), .ZN(new_n803));
  OAI21_X1  g378(.A(new_n803), .B1(G166), .B2(new_n727), .ZN(new_n804));
  XNOR2_X1  g379(.A(new_n804), .B(KEYINPUT95), .ZN(new_n805));
  AOI21_X1  g380(.A(new_n801), .B1(new_n805), .B2(G1971), .ZN(new_n806));
  OR2_X1    g381(.A1(new_n805), .A2(G1971), .ZN(new_n807));
  NAND3_X1  g382(.A1(new_n797), .A2(new_n806), .A3(new_n807), .ZN(new_n808));
  OR2_X1    g383(.A1(new_n808), .A2(KEYINPUT34), .ZN(new_n809));
  NAND2_X1  g384(.A1(new_n808), .A2(KEYINPUT34), .ZN(new_n810));
  NAND2_X1  g385(.A1(new_n721), .A2(G25), .ZN(new_n811));
  OR2_X1    g386(.A1(G95), .A2(G2105), .ZN(new_n812));
  OAI211_X1 g387(.A(new_n812), .B(G2104), .C1(G107), .C2(new_n465), .ZN(new_n813));
  XNOR2_X1  g388(.A(new_n813), .B(KEYINPUT92), .ZN(new_n814));
  INV_X1    g389(.A(G131), .ZN(new_n815));
  OAI21_X1  g390(.A(new_n814), .B1(new_n815), .B2(new_n716), .ZN(new_n816));
  AOI21_X1  g391(.A(new_n816), .B1(G119), .B2(new_n494), .ZN(new_n817));
  OAI21_X1  g392(.A(new_n811), .B1(new_n817), .B2(new_n721), .ZN(new_n818));
  XOR2_X1   g393(.A(KEYINPUT35), .B(G1991), .Z(new_n819));
  INV_X1    g394(.A(new_n819), .ZN(new_n820));
  XNOR2_X1  g395(.A(new_n818), .B(new_n820), .ZN(new_n821));
  AND2_X1   g396(.A1(new_n727), .A2(G24), .ZN(new_n822));
  AOI21_X1  g397(.A(new_n822), .B1(G290), .B2(G16), .ZN(new_n823));
  INV_X1    g398(.A(new_n823), .ZN(new_n824));
  AND2_X1   g399(.A1(new_n824), .A2(G1986), .ZN(new_n825));
  NOR2_X1   g400(.A1(new_n824), .A2(G1986), .ZN(new_n826));
  NOR3_X1   g401(.A1(new_n821), .A2(new_n825), .A3(new_n826), .ZN(new_n827));
  NAND3_X1  g402(.A1(new_n809), .A2(new_n810), .A3(new_n827), .ZN(new_n828));
  AND2_X1   g403(.A1(KEYINPUT96), .A2(KEYINPUT36), .ZN(new_n829));
  XNOR2_X1  g404(.A(new_n828), .B(new_n829), .ZN(new_n830));
  AND2_X1   g405(.A1(new_n792), .A2(new_n830), .ZN(G311));
  AND3_X1   g406(.A1(new_n792), .A2(new_n830), .A3(KEYINPUT103), .ZN(new_n832));
  AOI21_X1  g407(.A(KEYINPUT103), .B1(new_n792), .B2(new_n830), .ZN(new_n833));
  NOR2_X1   g408(.A1(new_n832), .A2(new_n833), .ZN(G150));
  AOI22_X1  g409(.A1(new_n517), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n835));
  NOR2_X1   g410(.A1(new_n835), .A2(new_n519), .ZN(new_n836));
  NAND2_X1  g411(.A1(new_n524), .A2(G55), .ZN(new_n837));
  INV_X1    g412(.A(G93), .ZN(new_n838));
  OAI21_X1  g413(.A(new_n837), .B1(new_n527), .B2(new_n838), .ZN(new_n839));
  OR2_X1    g414(.A1(new_n836), .A2(new_n839), .ZN(new_n840));
  INV_X1    g415(.A(KEYINPUT104), .ZN(new_n841));
  AOI21_X1  g416(.A(new_n556), .B1(new_n840), .B2(new_n841), .ZN(new_n842));
  NOR2_X1   g417(.A1(new_n836), .A2(new_n839), .ZN(new_n843));
  NAND2_X1  g418(.A1(new_n843), .A2(KEYINPUT104), .ZN(new_n844));
  NAND2_X1  g419(.A1(new_n842), .A2(new_n844), .ZN(new_n845));
  NAND3_X1  g420(.A1(new_n556), .A2(new_n843), .A3(KEYINPUT104), .ZN(new_n846));
  AND2_X1   g421(.A1(new_n845), .A2(new_n846), .ZN(new_n847));
  XNOR2_X1  g422(.A(new_n847), .B(KEYINPUT38), .ZN(new_n848));
  NOR2_X1   g423(.A1(new_n610), .A2(new_n619), .ZN(new_n849));
  XNOR2_X1  g424(.A(new_n848), .B(new_n849), .ZN(new_n850));
  INV_X1    g425(.A(KEYINPUT39), .ZN(new_n851));
  AOI21_X1  g426(.A(G860), .B1(new_n850), .B2(new_n851), .ZN(new_n852));
  OAI21_X1  g427(.A(new_n852), .B1(new_n851), .B2(new_n850), .ZN(new_n853));
  NAND2_X1  g428(.A1(new_n840), .A2(G860), .ZN(new_n854));
  XOR2_X1   g429(.A(KEYINPUT105), .B(KEYINPUT37), .Z(new_n855));
  XNOR2_X1  g430(.A(new_n854), .B(new_n855), .ZN(new_n856));
  NAND2_X1  g431(.A1(new_n853), .A2(new_n856), .ZN(G145));
  XOR2_X1   g432(.A(G162), .B(new_n636), .Z(new_n858));
  XNOR2_X1  g433(.A(new_n858), .B(G160), .ZN(new_n859));
  INV_X1    g434(.A(new_n859), .ZN(new_n860));
  NOR2_X1   g435(.A1(new_n717), .A2(new_n718), .ZN(new_n861));
  XNOR2_X1  g436(.A(new_n861), .B(new_n748), .ZN(new_n862));
  XOR2_X1   g437(.A(new_n817), .B(new_n627), .Z(new_n863));
  XNOR2_X1  g438(.A(new_n862), .B(new_n863), .ZN(new_n864));
  XNOR2_X1  g439(.A(new_n777), .B(G164), .ZN(new_n865));
  NAND2_X1  g440(.A1(new_n483), .A2(G142), .ZN(new_n866));
  NOR2_X1   g441(.A1(new_n465), .A2(G118), .ZN(new_n867));
  OAI21_X1  g442(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n868));
  OAI21_X1  g443(.A(new_n866), .B1(new_n867), .B2(new_n868), .ZN(new_n869));
  AOI21_X1  g444(.A(new_n869), .B1(new_n494), .B2(G130), .ZN(new_n870));
  XNOR2_X1  g445(.A(new_n865), .B(new_n870), .ZN(new_n871));
  NAND2_X1  g446(.A1(new_n864), .A2(new_n871), .ZN(new_n872));
  INV_X1    g447(.A(new_n872), .ZN(new_n873));
  NOR2_X1   g448(.A1(new_n864), .A2(new_n871), .ZN(new_n874));
  OAI21_X1  g449(.A(new_n860), .B1(new_n873), .B2(new_n874), .ZN(new_n875));
  INV_X1    g450(.A(new_n874), .ZN(new_n876));
  NAND3_X1  g451(.A1(new_n876), .A2(new_n859), .A3(new_n872), .ZN(new_n877));
  INV_X1    g452(.A(G37), .ZN(new_n878));
  NAND3_X1  g453(.A1(new_n875), .A2(new_n877), .A3(new_n878), .ZN(new_n879));
  XNOR2_X1  g454(.A(new_n879), .B(KEYINPUT40), .ZN(G395));
  XNOR2_X1  g455(.A(new_n847), .B(new_n622), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n618), .A2(G299), .ZN(new_n882));
  NAND2_X1  g457(.A1(new_n610), .A2(new_n581), .ZN(new_n883));
  NAND3_X1  g458(.A1(new_n882), .A2(KEYINPUT106), .A3(new_n883), .ZN(new_n884));
  OR3_X1    g459(.A1(new_n610), .A2(new_n581), .A3(KEYINPUT106), .ZN(new_n885));
  NAND2_X1  g460(.A1(new_n884), .A2(new_n885), .ZN(new_n886));
  INV_X1    g461(.A(new_n886), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n881), .A2(new_n887), .ZN(new_n888));
  OR3_X1    g463(.A1(new_n618), .A2(G299), .A3(KEYINPUT107), .ZN(new_n889));
  NAND3_X1  g464(.A1(new_n882), .A2(KEYINPUT107), .A3(new_n883), .ZN(new_n890));
  INV_X1    g465(.A(KEYINPUT41), .ZN(new_n891));
  NAND3_X1  g466(.A1(new_n889), .A2(new_n890), .A3(new_n891), .ZN(new_n892));
  INV_X1    g467(.A(new_n892), .ZN(new_n893));
  AOI21_X1  g468(.A(new_n891), .B1(new_n884), .B2(new_n885), .ZN(new_n894));
  NOR2_X1   g469(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  OAI21_X1  g470(.A(new_n888), .B1(new_n895), .B2(new_n881), .ZN(new_n896));
  OR2_X1    g471(.A1(new_n896), .A2(KEYINPUT42), .ZN(new_n897));
  XOR2_X1   g472(.A(G166), .B(G305), .Z(new_n898));
  NAND2_X1  g473(.A1(G290), .A2(G288), .ZN(new_n899));
  NAND3_X1  g474(.A1(new_n600), .A2(new_n794), .A3(new_n601), .ZN(new_n900));
  NAND2_X1  g475(.A1(new_n899), .A2(new_n900), .ZN(new_n901));
  INV_X1    g476(.A(KEYINPUT108), .ZN(new_n902));
  AOI21_X1  g477(.A(new_n898), .B1(new_n901), .B2(new_n902), .ZN(new_n903));
  NAND3_X1  g478(.A1(new_n899), .A2(KEYINPUT108), .A3(new_n900), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n903), .A2(new_n904), .ZN(new_n905));
  NAND4_X1  g480(.A1(new_n898), .A2(new_n899), .A3(KEYINPUT108), .A4(new_n900), .ZN(new_n906));
  NAND2_X1  g481(.A1(new_n905), .A2(new_n906), .ZN(new_n907));
  INV_X1    g482(.A(new_n907), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n896), .A2(KEYINPUT42), .ZN(new_n909));
  AND3_X1   g484(.A1(new_n897), .A2(new_n908), .A3(new_n909), .ZN(new_n910));
  AOI21_X1  g485(.A(new_n908), .B1(new_n897), .B2(new_n909), .ZN(new_n911));
  OAI21_X1  g486(.A(G868), .B1(new_n910), .B2(new_n911), .ZN(new_n912));
  OAI21_X1  g487(.A(new_n912), .B1(G868), .B2(new_n843), .ZN(G295));
  OAI21_X1  g488(.A(new_n912), .B1(G868), .B2(new_n843), .ZN(G331));
  NAND2_X1  g489(.A1(G301), .A2(G286), .ZN(new_n915));
  NAND2_X1  g490(.A1(G171), .A2(G168), .ZN(new_n916));
  NAND3_X1  g491(.A1(new_n847), .A2(new_n915), .A3(new_n916), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n916), .A2(new_n915), .ZN(new_n918));
  NAND2_X1  g493(.A1(new_n845), .A2(new_n846), .ZN(new_n919));
  NAND2_X1  g494(.A1(new_n918), .A2(new_n919), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n917), .A2(new_n920), .ZN(new_n921));
  OAI21_X1  g496(.A(new_n921), .B1(new_n893), .B2(new_n894), .ZN(new_n922));
  OAI211_X1 g497(.A(new_n908), .B(new_n922), .C1(new_n886), .C2(new_n921), .ZN(new_n923));
  NAND2_X1  g498(.A1(new_n886), .A2(KEYINPUT41), .ZN(new_n924));
  AOI22_X1  g499(.A1(new_n924), .A2(new_n892), .B1(new_n917), .B2(new_n920), .ZN(new_n925));
  NOR2_X1   g500(.A1(new_n921), .A2(new_n886), .ZN(new_n926));
  OAI21_X1  g501(.A(new_n907), .B1(new_n925), .B2(new_n926), .ZN(new_n927));
  NAND3_X1  g502(.A1(new_n923), .A2(new_n927), .A3(new_n878), .ZN(new_n928));
  INV_X1    g503(.A(KEYINPUT43), .ZN(new_n929));
  AND2_X1   g504(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  AOI21_X1  g505(.A(new_n891), .B1(new_n917), .B2(new_n920), .ZN(new_n931));
  NAND3_X1  g506(.A1(new_n931), .A2(new_n889), .A3(new_n890), .ZN(new_n932));
  OAI211_X1 g507(.A(new_n932), .B(new_n907), .C1(new_n887), .C2(new_n931), .ZN(new_n933));
  AND4_X1   g508(.A1(KEYINPUT43), .A2(new_n933), .A3(new_n923), .A4(new_n878), .ZN(new_n934));
  OAI21_X1  g509(.A(KEYINPUT44), .B1(new_n930), .B2(new_n934), .ZN(new_n935));
  AOI21_X1  g510(.A(KEYINPUT109), .B1(new_n928), .B2(KEYINPUT43), .ZN(new_n936));
  NAND2_X1  g511(.A1(new_n928), .A2(KEYINPUT43), .ZN(new_n937));
  NAND4_X1  g512(.A1(new_n933), .A2(new_n923), .A3(new_n929), .A4(new_n878), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n937), .A2(new_n938), .ZN(new_n939));
  AOI21_X1  g514(.A(new_n936), .B1(new_n939), .B2(KEYINPUT109), .ZN(new_n940));
  OAI21_X1  g515(.A(new_n935), .B1(new_n940), .B2(KEYINPUT44), .ZN(G397));
  INV_X1    g516(.A(KEYINPUT72), .ZN(new_n942));
  INV_X1    g517(.A(G114), .ZN(new_n943));
  NAND2_X1  g518(.A1(new_n942), .A2(new_n943), .ZN(new_n944));
  NAND2_X1  g519(.A1(KEYINPUT72), .A2(G114), .ZN(new_n945));
  NAND3_X1  g520(.A1(new_n944), .A2(G2105), .A3(new_n945), .ZN(new_n946));
  OAI21_X1  g521(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n947));
  INV_X1    g522(.A(new_n947), .ZN(new_n948));
  AOI22_X1  g523(.A1(new_n504), .A2(new_n488), .B1(new_n946), .B2(new_n948), .ZN(new_n949));
  AOI21_X1  g524(.A(G1384), .B1(new_n949), .B2(new_n500), .ZN(new_n950));
  INV_X1    g525(.A(G125), .ZN(new_n951));
  AOI21_X1  g526(.A(new_n951), .B1(new_n481), .B2(new_n482), .ZN(new_n952));
  INV_X1    g527(.A(new_n476), .ZN(new_n953));
  OAI21_X1  g528(.A(G2105), .B1(new_n952), .B2(new_n953), .ZN(new_n954));
  NAND4_X1  g529(.A1(new_n954), .A2(G40), .A3(new_n473), .A4(new_n470), .ZN(new_n955));
  XNOR2_X1  g530(.A(KEYINPUT110), .B(KEYINPUT45), .ZN(new_n956));
  NOR3_X1   g531(.A1(new_n950), .A2(new_n955), .A3(new_n956), .ZN(new_n957));
  XNOR2_X1  g532(.A(new_n817), .B(new_n820), .ZN(new_n958));
  XNOR2_X1  g533(.A(new_n958), .B(KEYINPUT111), .ZN(new_n959));
  XNOR2_X1  g534(.A(new_n777), .B(G2067), .ZN(new_n960));
  XNOR2_X1  g535(.A(new_n861), .B(G1996), .ZN(new_n961));
  NAND3_X1  g536(.A1(new_n959), .A2(new_n960), .A3(new_n961), .ZN(new_n962));
  XNOR2_X1  g537(.A(G290), .B(G1986), .ZN(new_n963));
  OAI21_X1  g538(.A(new_n957), .B1(new_n962), .B2(new_n963), .ZN(new_n964));
  XOR2_X1   g539(.A(KEYINPUT114), .B(G8), .Z(new_n965));
  INV_X1    g540(.A(new_n965), .ZN(new_n966));
  INV_X1    g541(.A(G40), .ZN(new_n967));
  NOR3_X1   g542(.A1(new_n474), .A2(new_n477), .A3(new_n967), .ZN(new_n968));
  INV_X1    g543(.A(KEYINPUT50), .ZN(new_n969));
  OAI21_X1  g544(.A(new_n968), .B1(new_n950), .B2(new_n969), .ZN(new_n970));
  AOI211_X1 g545(.A(KEYINPUT50), .B(G1384), .C1(new_n949), .C2(new_n500), .ZN(new_n971));
  NOR3_X1   g546(.A1(new_n970), .A2(G2090), .A3(new_n971), .ZN(new_n972));
  XOR2_X1   g547(.A(KEYINPUT112), .B(G1971), .Z(new_n973));
  INV_X1    g548(.A(new_n973), .ZN(new_n974));
  INV_X1    g549(.A(G1384), .ZN(new_n975));
  INV_X1    g550(.A(new_n503), .ZN(new_n976));
  INV_X1    g551(.A(G138), .ZN(new_n977));
  NOR2_X1   g552(.A1(new_n977), .A2(G2105), .ZN(new_n978));
  AOI21_X1  g553(.A(new_n976), .B1(new_n498), .B2(new_n978), .ZN(new_n979));
  NOR2_X1   g554(.A1(new_n471), .A2(new_n472), .ZN(new_n980));
  OAI21_X1  g555(.A(new_n509), .B1(new_n979), .B2(new_n980), .ZN(new_n981));
  AOI21_X1  g556(.A(new_n498), .B1(new_n483), .B2(G138), .ZN(new_n982));
  OAI21_X1  g557(.A(new_n975), .B1(new_n981), .B2(new_n982), .ZN(new_n983));
  INV_X1    g558(.A(new_n956), .ZN(new_n984));
  AOI21_X1  g559(.A(new_n955), .B1(new_n983), .B2(new_n984), .ZN(new_n985));
  OAI211_X1 g560(.A(KEYINPUT45), .B(new_n975), .C1(new_n981), .C2(new_n982), .ZN(new_n986));
  AOI21_X1  g561(.A(new_n974), .B1(new_n985), .B2(new_n986), .ZN(new_n987));
  OAI21_X1  g562(.A(new_n966), .B1(new_n972), .B2(new_n987), .ZN(new_n988));
  OAI21_X1  g563(.A(G8), .B1(new_n520), .B2(new_n529), .ZN(new_n989));
  XNOR2_X1  g564(.A(KEYINPUT113), .B(KEYINPUT55), .ZN(new_n990));
  XNOR2_X1  g565(.A(new_n989), .B(new_n990), .ZN(new_n991));
  INV_X1    g566(.A(new_n991), .ZN(new_n992));
  NAND2_X1  g567(.A1(new_n988), .A2(new_n992), .ZN(new_n993));
  OAI211_X1 g568(.A(new_n986), .B(new_n968), .C1(new_n950), .C2(new_n956), .ZN(new_n994));
  NAND2_X1  g569(.A1(new_n994), .A2(new_n973), .ZN(new_n995));
  AOI21_X1  g570(.A(new_n955), .B1(new_n983), .B2(KEYINPUT50), .ZN(new_n996));
  NAND2_X1  g571(.A1(new_n950), .A2(new_n969), .ZN(new_n997));
  NAND2_X1  g572(.A1(new_n996), .A2(new_n997), .ZN(new_n998));
  OAI21_X1  g573(.A(new_n995), .B1(G2090), .B2(new_n998), .ZN(new_n999));
  NAND3_X1  g574(.A1(new_n999), .A2(G8), .A3(new_n991), .ZN(new_n1000));
  NAND4_X1  g575(.A1(G160), .A2(G40), .A3(new_n975), .A4(new_n510), .ZN(new_n1001));
  NAND4_X1  g576(.A1(new_n584), .A2(new_n585), .A3(G1976), .A4(new_n586), .ZN(new_n1002));
  INV_X1    g577(.A(KEYINPUT115), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n1002), .A2(new_n1003), .ZN(new_n1004));
  AOI22_X1  g579(.A1(new_n538), .A2(G87), .B1(new_n524), .B2(G49), .ZN(new_n1005));
  NAND4_X1  g580(.A1(new_n1005), .A2(KEYINPUT115), .A3(G1976), .A4(new_n584), .ZN(new_n1006));
  NAND4_X1  g581(.A1(new_n1001), .A2(new_n966), .A3(new_n1004), .A4(new_n1006), .ZN(new_n1007));
  NAND2_X1  g582(.A1(new_n1007), .A2(KEYINPUT52), .ZN(new_n1008));
  INV_X1    g583(.A(KEYINPUT49), .ZN(new_n1009));
  AND3_X1   g584(.A1(new_n588), .A2(new_n692), .A3(new_n593), .ZN(new_n1010));
  AOI21_X1  g585(.A(new_n692), .B1(new_n588), .B2(new_n593), .ZN(new_n1011));
  OAI21_X1  g586(.A(new_n1009), .B1(new_n1010), .B2(new_n1011), .ZN(new_n1012));
  AOI21_X1  g587(.A(new_n965), .B1(new_n968), .B2(new_n950), .ZN(new_n1013));
  NAND2_X1  g588(.A1(new_n517), .A2(G61), .ZN(new_n1014));
  AOI21_X1  g589(.A(new_n519), .B1(new_n1014), .B2(new_n591), .ZN(new_n1015));
  NAND3_X1  g590(.A1(new_n517), .A2(G86), .A3(new_n526), .ZN(new_n1016));
  NAND2_X1  g591(.A1(new_n524), .A2(G48), .ZN(new_n1017));
  NAND2_X1  g592(.A1(new_n1016), .A2(new_n1017), .ZN(new_n1018));
  OAI21_X1  g593(.A(G1981), .B1(new_n1015), .B2(new_n1018), .ZN(new_n1019));
  NAND3_X1  g594(.A1(new_n588), .A2(new_n692), .A3(new_n593), .ZN(new_n1020));
  NAND3_X1  g595(.A1(new_n1019), .A2(KEYINPUT49), .A3(new_n1020), .ZN(new_n1021));
  NAND3_X1  g596(.A1(new_n1012), .A2(new_n1013), .A3(new_n1021), .ZN(new_n1022));
  INV_X1    g597(.A(G1976), .ZN(new_n1023));
  AOI21_X1  g598(.A(KEYINPUT52), .B1(G288), .B2(new_n1023), .ZN(new_n1024));
  NAND4_X1  g599(.A1(new_n1013), .A2(new_n1004), .A3(new_n1006), .A4(new_n1024), .ZN(new_n1025));
  AND3_X1   g600(.A1(new_n1008), .A2(new_n1022), .A3(new_n1025), .ZN(new_n1026));
  INV_X1    g601(.A(G1966), .ZN(new_n1027));
  NAND3_X1  g602(.A1(new_n510), .A2(new_n975), .A3(new_n956), .ZN(new_n1028));
  NAND2_X1  g603(.A1(new_n1028), .A2(new_n968), .ZN(new_n1029));
  AOI21_X1  g604(.A(KEYINPUT45), .B1(new_n510), .B2(new_n975), .ZN(new_n1030));
  OAI21_X1  g605(.A(new_n1027), .B1(new_n1029), .B2(new_n1030), .ZN(new_n1031));
  INV_X1    g606(.A(G2084), .ZN(new_n1032));
  NAND3_X1  g607(.A1(new_n996), .A2(new_n1032), .A3(new_n997), .ZN(new_n1033));
  AOI211_X1 g608(.A(G286), .B(new_n965), .C1(new_n1031), .C2(new_n1033), .ZN(new_n1034));
  NAND4_X1  g609(.A1(new_n993), .A2(new_n1000), .A3(new_n1026), .A4(new_n1034), .ZN(new_n1035));
  INV_X1    g610(.A(KEYINPUT63), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n1035), .A2(new_n1036), .ZN(new_n1037));
  INV_X1    g612(.A(KEYINPUT117), .ZN(new_n1038));
  NAND2_X1  g613(.A1(new_n1037), .A2(new_n1038), .ZN(new_n1039));
  NAND3_X1  g614(.A1(new_n1035), .A2(KEYINPUT117), .A3(new_n1036), .ZN(new_n1040));
  NAND3_X1  g615(.A1(new_n1008), .A2(new_n1022), .A3(new_n1025), .ZN(new_n1041));
  XNOR2_X1  g616(.A(new_n1041), .B(KEYINPUT116), .ZN(new_n1042));
  AND3_X1   g617(.A1(new_n999), .A2(G8), .A3(new_n991), .ZN(new_n1043));
  NOR2_X1   g618(.A1(new_n1043), .A2(new_n1036), .ZN(new_n1044));
  NAND2_X1  g619(.A1(new_n999), .A2(G8), .ZN(new_n1045));
  NAND2_X1  g620(.A1(new_n1045), .A2(new_n992), .ZN(new_n1046));
  NAND4_X1  g621(.A1(new_n1042), .A2(new_n1044), .A3(new_n1034), .A4(new_n1046), .ZN(new_n1047));
  NAND3_X1  g622(.A1(new_n1039), .A2(new_n1040), .A3(new_n1047), .ZN(new_n1048));
  NAND3_X1  g623(.A1(new_n1022), .A2(new_n1023), .A3(new_n794), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n1049), .A2(new_n1020), .ZN(new_n1050));
  AOI22_X1  g625(.A1(new_n1042), .A2(new_n1043), .B1(new_n1013), .B2(new_n1050), .ZN(new_n1051));
  NAND2_X1  g626(.A1(new_n1048), .A2(new_n1051), .ZN(new_n1052));
  NAND2_X1  g627(.A1(new_n1031), .A2(new_n1033), .ZN(new_n1053));
  NAND3_X1  g628(.A1(new_n1053), .A2(KEYINPUT122), .A3(new_n966), .ZN(new_n1054));
  NAND2_X1  g629(.A1(G286), .A2(new_n966), .ZN(new_n1055));
  INV_X1    g630(.A(KEYINPUT51), .ZN(new_n1056));
  NAND2_X1  g631(.A1(new_n1055), .A2(new_n1056), .ZN(new_n1057));
  INV_X1    g632(.A(new_n1057), .ZN(new_n1058));
  NAND2_X1  g633(.A1(new_n1054), .A2(new_n1058), .ZN(new_n1059));
  AOI21_X1  g634(.A(new_n965), .B1(new_n1031), .B2(new_n1033), .ZN(new_n1060));
  NOR2_X1   g635(.A1(new_n1060), .A2(KEYINPUT122), .ZN(new_n1061));
  OAI21_X1  g636(.A(KEYINPUT123), .B1(new_n1059), .B2(new_n1061), .ZN(new_n1062));
  NAND2_X1  g637(.A1(new_n1053), .A2(new_n966), .ZN(new_n1063));
  INV_X1    g638(.A(KEYINPUT122), .ZN(new_n1064));
  NAND2_X1  g639(.A1(new_n1063), .A2(new_n1064), .ZN(new_n1065));
  AOI21_X1  g640(.A(new_n1057), .B1(new_n1060), .B2(KEYINPUT122), .ZN(new_n1066));
  INV_X1    g641(.A(KEYINPUT123), .ZN(new_n1067));
  NAND3_X1  g642(.A1(new_n1065), .A2(new_n1066), .A3(new_n1067), .ZN(new_n1068));
  NAND2_X1  g643(.A1(new_n1053), .A2(G8), .ZN(new_n1069));
  AOI21_X1  g644(.A(new_n1056), .B1(new_n1069), .B2(new_n1055), .ZN(new_n1070));
  INV_X1    g645(.A(new_n1070), .ZN(new_n1071));
  NAND3_X1  g646(.A1(new_n1062), .A2(new_n1068), .A3(new_n1071), .ZN(new_n1072));
  INV_X1    g647(.A(new_n1055), .ZN(new_n1073));
  NAND2_X1  g648(.A1(new_n1053), .A2(new_n1073), .ZN(new_n1074));
  NAND2_X1  g649(.A1(new_n1072), .A2(new_n1074), .ZN(new_n1075));
  OAI21_X1  g650(.A(new_n707), .B1(new_n970), .B2(new_n971), .ZN(new_n1076));
  INV_X1    g651(.A(KEYINPUT124), .ZN(new_n1077));
  NAND2_X1  g652(.A1(new_n1076), .A2(new_n1077), .ZN(new_n1078));
  NAND3_X1  g653(.A1(new_n998), .A2(KEYINPUT124), .A3(new_n707), .ZN(new_n1079));
  NAND2_X1  g654(.A1(new_n1078), .A2(new_n1079), .ZN(new_n1080));
  INV_X1    g655(.A(KEYINPUT53), .ZN(new_n1081));
  OAI21_X1  g656(.A(new_n1081), .B1(new_n994), .B2(G2078), .ZN(new_n1082));
  INV_X1    g657(.A(G2078), .ZN(new_n1083));
  NAND4_X1  g658(.A1(new_n985), .A2(KEYINPUT53), .A3(new_n1083), .A4(new_n986), .ZN(new_n1084));
  AND2_X1   g659(.A1(new_n1082), .A2(new_n1084), .ZN(new_n1085));
  NAND2_X1  g660(.A1(new_n1080), .A2(new_n1085), .ZN(new_n1086));
  NAND2_X1  g661(.A1(new_n1086), .A2(G171), .ZN(new_n1087));
  INV_X1    g662(.A(new_n1030), .ZN(new_n1088));
  NOR2_X1   g663(.A1(new_n1081), .A2(G2078), .ZN(new_n1089));
  NAND4_X1  g664(.A1(new_n1088), .A2(new_n968), .A3(new_n1028), .A4(new_n1089), .ZN(new_n1090));
  NAND4_X1  g665(.A1(new_n1082), .A2(G301), .A3(new_n1090), .A4(new_n1076), .ZN(new_n1091));
  AND2_X1   g666(.A1(new_n1091), .A2(KEYINPUT54), .ZN(new_n1092));
  NAND2_X1  g667(.A1(new_n1087), .A2(new_n1092), .ZN(new_n1093));
  AND3_X1   g668(.A1(new_n993), .A2(new_n1000), .A3(new_n1026), .ZN(new_n1094));
  NAND3_X1  g669(.A1(new_n1080), .A2(new_n1085), .A3(G301), .ZN(new_n1095));
  INV_X1    g670(.A(KEYINPUT125), .ZN(new_n1096));
  NAND3_X1  g671(.A1(new_n1082), .A2(new_n1090), .A3(new_n1076), .ZN(new_n1097));
  AOI21_X1  g672(.A(new_n1096), .B1(new_n1097), .B2(G171), .ZN(new_n1098));
  AND2_X1   g673(.A1(new_n1095), .A2(new_n1098), .ZN(new_n1099));
  NAND4_X1  g674(.A1(new_n1080), .A2(new_n1085), .A3(new_n1096), .A4(G301), .ZN(new_n1100));
  INV_X1    g675(.A(KEYINPUT54), .ZN(new_n1101));
  NAND2_X1  g676(.A1(new_n1100), .A2(new_n1101), .ZN(new_n1102));
  OAI211_X1 g677(.A(new_n1093), .B(new_n1094), .C1(new_n1099), .C2(new_n1102), .ZN(new_n1103));
  AOI21_X1  g678(.A(G1348), .B1(new_n996), .B2(new_n997), .ZN(new_n1104));
  NOR2_X1   g679(.A1(new_n1001), .A2(G2067), .ZN(new_n1105));
  NOR2_X1   g680(.A1(new_n1104), .A2(new_n1105), .ZN(new_n1106));
  NAND2_X1  g681(.A1(new_n1106), .A2(KEYINPUT60), .ZN(new_n1107));
  INV_X1    g682(.A(KEYINPUT60), .ZN(new_n1108));
  OAI21_X1  g683(.A(new_n1108), .B1(new_n1104), .B2(new_n1105), .ZN(new_n1109));
  NAND3_X1  g684(.A1(new_n1107), .A2(new_n1109), .A3(new_n618), .ZN(new_n1110));
  OR2_X1    g685(.A1(new_n577), .A2(new_n578), .ZN(new_n1111));
  AOI22_X1  g686(.A1(new_n1111), .A2(G651), .B1(new_n572), .B2(new_n574), .ZN(new_n1112));
  INV_X1    g687(.A(KEYINPUT118), .ZN(new_n1113));
  AOI21_X1  g688(.A(new_n1113), .B1(new_n572), .B2(new_n574), .ZN(new_n1114));
  OAI211_X1 g689(.A(new_n1112), .B(new_n568), .C1(KEYINPUT57), .C2(new_n1114), .ZN(new_n1115));
  AOI21_X1  g690(.A(KEYINPUT57), .B1(new_n575), .B2(KEYINPUT118), .ZN(new_n1116));
  OAI21_X1  g691(.A(new_n1116), .B1(new_n569), .B2(new_n580), .ZN(new_n1117));
  XNOR2_X1  g692(.A(KEYINPUT56), .B(G2072), .ZN(new_n1118));
  XNOR2_X1  g693(.A(new_n1118), .B(KEYINPUT119), .ZN(new_n1119));
  INV_X1    g694(.A(new_n1119), .ZN(new_n1120));
  NOR2_X1   g695(.A1(new_n994), .A2(new_n1120), .ZN(new_n1121));
  AOI21_X1  g696(.A(G1956), .B1(new_n996), .B2(new_n997), .ZN(new_n1122));
  OAI211_X1 g697(.A(new_n1115), .B(new_n1117), .C1(new_n1121), .C2(new_n1122), .ZN(new_n1123));
  INV_X1    g698(.A(G1956), .ZN(new_n1124));
  NAND2_X1  g699(.A1(new_n998), .A2(new_n1124), .ZN(new_n1125));
  NAND2_X1  g700(.A1(new_n1117), .A2(new_n1115), .ZN(new_n1126));
  NAND3_X1  g701(.A1(new_n985), .A2(new_n986), .A3(new_n1119), .ZN(new_n1127));
  NAND3_X1  g702(.A1(new_n1125), .A2(new_n1126), .A3(new_n1127), .ZN(new_n1128));
  NAND3_X1  g703(.A1(new_n1123), .A2(new_n1128), .A3(KEYINPUT61), .ZN(new_n1129));
  NAND2_X1  g704(.A1(new_n1110), .A2(new_n1129), .ZN(new_n1130));
  NOR2_X1   g705(.A1(new_n983), .A2(new_n955), .ZN(new_n1131));
  XNOR2_X1  g706(.A(KEYINPUT58), .B(G1341), .ZN(new_n1132));
  OAI22_X1  g707(.A1(new_n994), .A2(G1996), .B1(new_n1131), .B2(new_n1132), .ZN(new_n1133));
  NAND2_X1  g708(.A1(new_n1133), .A2(new_n556), .ZN(new_n1134));
  INV_X1    g709(.A(KEYINPUT59), .ZN(new_n1135));
  NAND2_X1  g710(.A1(new_n1134), .A2(new_n1135), .ZN(new_n1136));
  NAND3_X1  g711(.A1(new_n1133), .A2(KEYINPUT59), .A3(new_n556), .ZN(new_n1137));
  OAI211_X1 g712(.A(new_n1136), .B(new_n1137), .C1(new_n1107), .C2(new_n618), .ZN(new_n1138));
  NOR2_X1   g713(.A1(new_n1130), .A2(new_n1138), .ZN(new_n1139));
  INV_X1    g714(.A(KEYINPUT120), .ZN(new_n1140));
  NAND2_X1  g715(.A1(new_n1128), .A2(new_n1140), .ZN(new_n1141));
  AOI21_X1  g716(.A(new_n1126), .B1(new_n1125), .B2(new_n1127), .ZN(new_n1142));
  NOR2_X1   g717(.A1(new_n1141), .A2(new_n1142), .ZN(new_n1143));
  INV_X1    g718(.A(KEYINPUT61), .ZN(new_n1144));
  OAI21_X1  g719(.A(new_n1144), .B1(new_n1123), .B2(new_n1140), .ZN(new_n1145));
  OAI21_X1  g720(.A(KEYINPUT121), .B1(new_n1143), .B2(new_n1145), .ZN(new_n1146));
  AOI21_X1  g721(.A(KEYINPUT61), .B1(new_n1142), .B2(KEYINPUT120), .ZN(new_n1147));
  INV_X1    g722(.A(KEYINPUT121), .ZN(new_n1148));
  OAI211_X1 g723(.A(new_n1147), .B(new_n1148), .C1(new_n1142), .C2(new_n1141), .ZN(new_n1149));
  NAND3_X1  g724(.A1(new_n1139), .A2(new_n1146), .A3(new_n1149), .ZN(new_n1150));
  NOR2_X1   g725(.A1(new_n1106), .A2(new_n610), .ZN(new_n1151));
  AOI21_X1  g726(.A(new_n1142), .B1(new_n1151), .B2(new_n1128), .ZN(new_n1152));
  AOI21_X1  g727(.A(new_n1103), .B1(new_n1150), .B2(new_n1152), .ZN(new_n1153));
  AOI21_X1  g728(.A(new_n1052), .B1(new_n1075), .B2(new_n1153), .ZN(new_n1154));
  INV_X1    g729(.A(KEYINPUT62), .ZN(new_n1155));
  NAND3_X1  g730(.A1(new_n1072), .A2(new_n1155), .A3(new_n1074), .ZN(new_n1156));
  AND3_X1   g731(.A1(new_n1094), .A2(G171), .A3(new_n1097), .ZN(new_n1157));
  NAND2_X1  g732(.A1(new_n1156), .A2(new_n1157), .ZN(new_n1158));
  INV_X1    g733(.A(KEYINPUT126), .ZN(new_n1159));
  INV_X1    g734(.A(new_n1074), .ZN(new_n1160));
  NAND2_X1  g735(.A1(new_n1065), .A2(new_n1066), .ZN(new_n1161));
  AOI21_X1  g736(.A(new_n1070), .B1(new_n1161), .B2(KEYINPUT123), .ZN(new_n1162));
  AOI21_X1  g737(.A(new_n1160), .B1(new_n1162), .B2(new_n1068), .ZN(new_n1163));
  OAI21_X1  g738(.A(new_n1159), .B1(new_n1163), .B2(new_n1155), .ZN(new_n1164));
  NAND3_X1  g739(.A1(new_n1075), .A2(KEYINPUT126), .A3(KEYINPUT62), .ZN(new_n1165));
  AOI21_X1  g740(.A(new_n1158), .B1(new_n1164), .B2(new_n1165), .ZN(new_n1166));
  INV_X1    g741(.A(KEYINPUT127), .ZN(new_n1167));
  OAI21_X1  g742(.A(new_n1154), .B1(new_n1166), .B2(new_n1167), .ZN(new_n1168));
  AND2_X1   g743(.A1(new_n1156), .A2(new_n1157), .ZN(new_n1169));
  AOI21_X1  g744(.A(KEYINPUT126), .B1(new_n1075), .B2(KEYINPUT62), .ZN(new_n1170));
  AOI211_X1 g745(.A(new_n1159), .B(new_n1155), .C1(new_n1072), .C2(new_n1074), .ZN(new_n1171));
  OAI211_X1 g746(.A(new_n1169), .B(new_n1167), .C1(new_n1170), .C2(new_n1171), .ZN(new_n1172));
  INV_X1    g747(.A(new_n1172), .ZN(new_n1173));
  OAI21_X1  g748(.A(new_n964), .B1(new_n1168), .B2(new_n1173), .ZN(new_n1174));
  NAND2_X1  g749(.A1(new_n960), .A2(new_n861), .ZN(new_n1175));
  INV_X1    g750(.A(G1996), .ZN(new_n1176));
  NAND2_X1  g751(.A1(new_n957), .A2(new_n1176), .ZN(new_n1177));
  NAND2_X1  g752(.A1(new_n1177), .A2(KEYINPUT46), .ZN(new_n1178));
  OR2_X1    g753(.A1(new_n1177), .A2(KEYINPUT46), .ZN(new_n1179));
  AOI22_X1  g754(.A1(new_n1175), .A2(new_n957), .B1(new_n1178), .B2(new_n1179), .ZN(new_n1180));
  XNOR2_X1  g755(.A(new_n1180), .B(KEYINPUT47), .ZN(new_n1181));
  INV_X1    g756(.A(G2067), .ZN(new_n1182));
  NAND2_X1  g757(.A1(new_n777), .A2(new_n1182), .ZN(new_n1183));
  NAND2_X1  g758(.A1(new_n961), .A2(new_n960), .ZN(new_n1184));
  NAND2_X1  g759(.A1(new_n817), .A2(new_n819), .ZN(new_n1185));
  OAI21_X1  g760(.A(new_n1183), .B1(new_n1184), .B2(new_n1185), .ZN(new_n1186));
  AND2_X1   g761(.A1(new_n1186), .A2(new_n957), .ZN(new_n1187));
  NAND2_X1  g762(.A1(new_n962), .A2(new_n957), .ZN(new_n1188));
  NOR2_X1   g763(.A1(G290), .A2(G1986), .ZN(new_n1189));
  NAND2_X1  g764(.A1(new_n1189), .A2(new_n957), .ZN(new_n1190));
  XNOR2_X1  g765(.A(new_n1190), .B(KEYINPUT48), .ZN(new_n1191));
  AOI211_X1 g766(.A(new_n1181), .B(new_n1187), .C1(new_n1188), .C2(new_n1191), .ZN(new_n1192));
  NAND2_X1  g767(.A1(new_n1174), .A2(new_n1192), .ZN(G329));
  assign    G231 = 1'b0;
  NOR3_X1   g768(.A1(G401), .A2(new_n463), .A3(G227), .ZN(new_n1195));
  NAND4_X1  g769(.A1(new_n700), .A2(new_n703), .A3(new_n879), .A4(new_n1195), .ZN(new_n1196));
  NOR2_X1   g770(.A1(new_n940), .A2(new_n1196), .ZN(G308));
  AND4_X1   g771(.A1(new_n700), .A2(new_n703), .A3(new_n879), .A4(new_n1195), .ZN(new_n1198));
  AND2_X1   g772(.A1(new_n939), .A2(KEYINPUT109), .ZN(new_n1199));
  OAI21_X1  g773(.A(new_n1198), .B1(new_n1199), .B2(new_n936), .ZN(G225));
endmodule


