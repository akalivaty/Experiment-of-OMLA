//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 1 1 1 1 0 0 0 0 0 0 1 0 1 1 1 1 1 1 1 1 1 1 1 0 0 1 1 0 0 0 1 1 0 1 0 1 1 0 0 0 0 1 0 1 0 1 0 0 1 1 1 0 1 0 1 0 1 1 0 0 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:41:59 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n245, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1246, new_n1247,
    new_n1248, new_n1249, new_n1251, new_n1252, new_n1253, new_n1254,
    new_n1256, new_n1257, new_n1258, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1321, new_n1322, new_n1323,
    new_n1324, new_n1325, new_n1326, new_n1327, new_n1328, new_n1329;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0005(.A1(G1), .A2(G20), .ZN(new_n206));
  XOR2_X1   g0006(.A(new_n206), .B(KEYINPUT64), .Z(new_n207));
  NOR2_X1   g0007(.A1(new_n207), .A2(G13), .ZN(new_n208));
  OAI211_X1 g0008(.A(new_n208), .B(G250), .C1(G257), .C2(G264), .ZN(new_n209));
  INV_X1    g0009(.A(KEYINPUT0), .ZN(new_n210));
  NAND2_X1  g0010(.A1(G1), .A2(G13), .ZN(new_n211));
  INV_X1    g0011(.A(G20), .ZN(new_n212));
  NOR2_X1   g0012(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  INV_X1    g0013(.A(new_n201), .ZN(new_n214));
  NAND2_X1  g0014(.A1(new_n214), .A2(G50), .ZN(new_n215));
  INV_X1    g0015(.A(new_n215), .ZN(new_n216));
  AOI22_X1  g0016(.A1(new_n209), .A2(new_n210), .B1(new_n213), .B2(new_n216), .ZN(new_n217));
  OAI21_X1  g0017(.A(new_n217), .B1(new_n210), .B2(new_n209), .ZN(new_n218));
  AOI22_X1  g0018(.A1(G50), .A2(G226), .B1(G77), .B2(G244), .ZN(new_n219));
  AOI22_X1  g0019(.A1(G68), .A2(G238), .B1(G116), .B2(G270), .ZN(new_n220));
  NAND2_X1  g0020(.A1(new_n219), .A2(new_n220), .ZN(new_n221));
  NAND2_X1  g0021(.A1(new_n221), .A2(KEYINPUT65), .ZN(new_n222));
  AOI22_X1  g0022(.A1(G87), .A2(G250), .B1(G107), .B2(G264), .ZN(new_n223));
  AOI22_X1  g0023(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n224));
  NAND3_X1  g0024(.A1(new_n222), .A2(new_n223), .A3(new_n224), .ZN(new_n225));
  NOR2_X1   g0025(.A1(new_n221), .A2(KEYINPUT65), .ZN(new_n226));
  OAI21_X1  g0026(.A(new_n207), .B1(new_n225), .B2(new_n226), .ZN(new_n227));
  AND2_X1   g0027(.A1(new_n227), .A2(KEYINPUT1), .ZN(new_n228));
  NOR2_X1   g0028(.A1(new_n227), .A2(KEYINPUT1), .ZN(new_n229));
  NOR3_X1   g0029(.A1(new_n218), .A2(new_n228), .A3(new_n229), .ZN(G361));
  XNOR2_X1  g0030(.A(G238), .B(G244), .ZN(new_n231));
  XNOR2_X1  g0031(.A(new_n231), .B(KEYINPUT2), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n232), .B(G226), .ZN(new_n233));
  INV_X1    g0033(.A(G232), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n233), .B(new_n234), .ZN(new_n235));
  XOR2_X1   g0035(.A(G250), .B(G257), .Z(new_n236));
  XNOR2_X1  g0036(.A(G264), .B(G270), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XOR2_X1   g0038(.A(new_n235), .B(new_n238), .Z(G358));
  XOR2_X1   g0039(.A(G68), .B(G77), .Z(new_n240));
  XNOR2_X1  g0040(.A(G50), .B(G58), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XOR2_X1   g0042(.A(G87), .B(G97), .Z(new_n243));
  XNOR2_X1  g0043(.A(G107), .B(G116), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n242), .B(new_n245), .ZN(G351));
  OR2_X1    g0046(.A1(KEYINPUT3), .A2(G33), .ZN(new_n247));
  NAND2_X1  g0047(.A1(KEYINPUT3), .A2(G33), .ZN(new_n248));
  NAND2_X1  g0048(.A1(new_n247), .A2(new_n248), .ZN(new_n249));
  INV_X1    g0049(.A(G1698), .ZN(new_n250));
  NAND3_X1  g0050(.A1(new_n249), .A2(G222), .A3(new_n250), .ZN(new_n251));
  INV_X1    g0051(.A(G77), .ZN(new_n252));
  NAND2_X1  g0052(.A1(new_n249), .A2(G1698), .ZN(new_n253));
  INV_X1    g0053(.A(G223), .ZN(new_n254));
  OAI221_X1 g0054(.A(new_n251), .B1(new_n252), .B2(new_n249), .C1(new_n253), .C2(new_n254), .ZN(new_n255));
  AOI21_X1  g0055(.A(new_n211), .B1(G33), .B2(G41), .ZN(new_n256));
  NAND2_X1  g0056(.A1(new_n255), .A2(new_n256), .ZN(new_n257));
  NOR2_X1   g0057(.A1(G41), .A2(G45), .ZN(new_n258));
  INV_X1    g0058(.A(G274), .ZN(new_n259));
  NOR3_X1   g0059(.A1(new_n258), .A2(G1), .A3(new_n259), .ZN(new_n260));
  OAI21_X1  g0060(.A(KEYINPUT66), .B1(new_n258), .B2(G1), .ZN(new_n261));
  INV_X1    g0061(.A(KEYINPUT66), .ZN(new_n262));
  INV_X1    g0062(.A(G1), .ZN(new_n263));
  OAI211_X1 g0063(.A(new_n262), .B(new_n263), .C1(G41), .C2(G45), .ZN(new_n264));
  AOI21_X1  g0064(.A(new_n256), .B1(new_n261), .B2(new_n264), .ZN(new_n265));
  AOI21_X1  g0065(.A(new_n260), .B1(new_n265), .B2(G226), .ZN(new_n266));
  NAND2_X1  g0066(.A1(new_n257), .A2(new_n266), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n267), .A2(G169), .ZN(new_n268));
  INV_X1    g0068(.A(G179), .ZN(new_n269));
  OAI21_X1  g0069(.A(new_n268), .B1(new_n269), .B2(new_n267), .ZN(new_n270));
  NAND3_X1  g0070(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n271), .A2(new_n211), .ZN(new_n272));
  INV_X1    g0072(.A(new_n272), .ZN(new_n273));
  XNOR2_X1  g0073(.A(KEYINPUT8), .B(G58), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n212), .A2(G33), .ZN(new_n275));
  OR2_X1    g0075(.A1(new_n274), .A2(new_n275), .ZN(new_n276));
  NOR2_X1   g0076(.A1(G20), .A2(G33), .ZN(new_n277));
  AOI22_X1  g0077(.A1(new_n203), .A2(G20), .B1(G150), .B2(new_n277), .ZN(new_n278));
  AOI21_X1  g0078(.A(new_n273), .B1(new_n276), .B2(new_n278), .ZN(new_n279));
  OR2_X1    g0079(.A1(new_n279), .A2(KEYINPUT67), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n279), .A2(KEYINPUT67), .ZN(new_n281));
  NAND3_X1  g0081(.A1(new_n263), .A2(G13), .A3(G20), .ZN(new_n282));
  INV_X1    g0082(.A(new_n282), .ZN(new_n283));
  NOR2_X1   g0083(.A1(new_n283), .A2(new_n272), .ZN(new_n284));
  AOI21_X1  g0084(.A(new_n202), .B1(new_n263), .B2(G20), .ZN(new_n285));
  AOI22_X1  g0085(.A1(new_n284), .A2(new_n285), .B1(new_n202), .B2(new_n283), .ZN(new_n286));
  NAND3_X1  g0086(.A1(new_n280), .A2(new_n281), .A3(new_n286), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n270), .A2(new_n287), .ZN(new_n288));
  NAND2_X1  g0088(.A1(G20), .A2(G77), .ZN(new_n289));
  INV_X1    g0089(.A(new_n277), .ZN(new_n290));
  XNOR2_X1  g0090(.A(KEYINPUT15), .B(G87), .ZN(new_n291));
  OAI221_X1 g0091(.A(new_n289), .B1(new_n274), .B2(new_n290), .C1(new_n275), .C2(new_n291), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n292), .A2(new_n272), .ZN(new_n293));
  INV_X1    g0093(.A(G13), .ZN(new_n294));
  NOR2_X1   g0094(.A1(new_n294), .A2(G1), .ZN(new_n295));
  INV_X1    g0095(.A(KEYINPUT68), .ZN(new_n296));
  NAND3_X1  g0096(.A1(new_n295), .A2(new_n296), .A3(G20), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n282), .A2(KEYINPUT68), .ZN(new_n298));
  AOI21_X1  g0098(.A(new_n272), .B1(new_n297), .B2(new_n298), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n263), .A2(G20), .ZN(new_n300));
  NAND3_X1  g0100(.A1(new_n299), .A2(G77), .A3(new_n300), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n297), .A2(new_n298), .ZN(new_n302));
  INV_X1    g0102(.A(new_n302), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n303), .A2(new_n252), .ZN(new_n304));
  NAND3_X1  g0104(.A1(new_n293), .A2(new_n301), .A3(new_n304), .ZN(new_n305));
  NAND3_X1  g0105(.A1(new_n249), .A2(G232), .A3(new_n250), .ZN(new_n306));
  AND2_X1   g0106(.A1(KEYINPUT3), .A2(G33), .ZN(new_n307));
  NOR2_X1   g0107(.A1(KEYINPUT3), .A2(G33), .ZN(new_n308));
  NOR2_X1   g0108(.A1(new_n307), .A2(new_n308), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n309), .A2(G107), .ZN(new_n310));
  INV_X1    g0110(.A(G238), .ZN(new_n311));
  OAI211_X1 g0111(.A(new_n306), .B(new_n310), .C1(new_n253), .C2(new_n311), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n312), .A2(new_n256), .ZN(new_n313));
  AOI21_X1  g0113(.A(new_n260), .B1(new_n265), .B2(G244), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n313), .A2(new_n314), .ZN(new_n315));
  INV_X1    g0115(.A(new_n315), .ZN(new_n316));
  INV_X1    g0116(.A(G190), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n316), .A2(new_n317), .ZN(new_n318));
  INV_X1    g0118(.A(G200), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n315), .A2(new_n319), .ZN(new_n320));
  AOI21_X1  g0120(.A(new_n305), .B1(new_n318), .B2(new_n320), .ZN(new_n321));
  INV_X1    g0121(.A(new_n305), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n316), .A2(G179), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n315), .A2(G169), .ZN(new_n324));
  AOI21_X1  g0124(.A(new_n322), .B1(new_n323), .B2(new_n324), .ZN(new_n325));
  NOR2_X1   g0125(.A1(new_n321), .A2(new_n325), .ZN(new_n326));
  INV_X1    g0126(.A(KEYINPUT9), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n287), .A2(new_n327), .ZN(new_n328));
  NAND4_X1  g0128(.A1(new_n280), .A2(KEYINPUT9), .A3(new_n281), .A4(new_n286), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n267), .A2(G200), .ZN(new_n330));
  NAND3_X1  g0130(.A1(new_n257), .A2(G190), .A3(new_n266), .ZN(new_n331));
  NAND4_X1  g0131(.A1(new_n328), .A2(new_n329), .A3(new_n330), .A4(new_n331), .ZN(new_n332));
  AND2_X1   g0132(.A1(new_n332), .A2(KEYINPUT10), .ZN(new_n333));
  NOR2_X1   g0133(.A1(new_n332), .A2(KEYINPUT10), .ZN(new_n334));
  OAI211_X1 g0134(.A(new_n288), .B(new_n326), .C1(new_n333), .C2(new_n334), .ZN(new_n335));
  INV_X1    g0135(.A(new_n284), .ZN(new_n336));
  INV_X1    g0136(.A(new_n274), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n337), .A2(new_n300), .ZN(new_n338));
  OAI22_X1  g0138(.A1(new_n336), .A2(new_n338), .B1(new_n282), .B2(new_n337), .ZN(new_n339));
  INV_X1    g0139(.A(G58), .ZN(new_n340));
  INV_X1    g0140(.A(G68), .ZN(new_n341));
  NOR2_X1   g0141(.A1(new_n340), .A2(new_n341), .ZN(new_n342));
  OAI21_X1  g0142(.A(G20), .B1(new_n342), .B2(new_n201), .ZN(new_n343));
  NAND2_X1  g0143(.A1(new_n277), .A2(G159), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n343), .A2(new_n344), .ZN(new_n345));
  NOR3_X1   g0145(.A1(new_n307), .A2(new_n308), .A3(G20), .ZN(new_n346));
  OAI21_X1  g0146(.A(KEYINPUT72), .B1(new_n346), .B2(KEYINPUT7), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n346), .A2(KEYINPUT7), .ZN(new_n348));
  NAND3_X1  g0148(.A1(new_n247), .A2(new_n212), .A3(new_n248), .ZN(new_n349));
  INV_X1    g0149(.A(KEYINPUT72), .ZN(new_n350));
  INV_X1    g0150(.A(KEYINPUT7), .ZN(new_n351));
  NAND3_X1  g0151(.A1(new_n349), .A2(new_n350), .A3(new_n351), .ZN(new_n352));
  NAND3_X1  g0152(.A1(new_n347), .A2(new_n348), .A3(new_n352), .ZN(new_n353));
  AOI21_X1  g0153(.A(new_n345), .B1(new_n353), .B2(G68), .ZN(new_n354));
  AOI21_X1  g0154(.A(new_n273), .B1(new_n354), .B2(KEYINPUT16), .ZN(new_n355));
  INV_X1    g0155(.A(KEYINPUT16), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n349), .A2(new_n351), .ZN(new_n357));
  AOI21_X1  g0157(.A(new_n341), .B1(new_n348), .B2(new_n357), .ZN(new_n358));
  OAI21_X1  g0158(.A(new_n356), .B1(new_n358), .B2(new_n345), .ZN(new_n359));
  AOI21_X1  g0159(.A(new_n339), .B1(new_n355), .B2(new_n359), .ZN(new_n360));
  INV_X1    g0160(.A(G169), .ZN(new_n361));
  INV_X1    g0161(.A(new_n211), .ZN(new_n362));
  NAND2_X1  g0162(.A1(G33), .A2(G41), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n362), .A2(new_n363), .ZN(new_n364));
  INV_X1    g0164(.A(G33), .ZN(new_n365));
  INV_X1    g0165(.A(G87), .ZN(new_n366));
  NOR2_X1   g0166(.A1(new_n365), .A2(new_n366), .ZN(new_n367));
  NOR2_X1   g0167(.A1(new_n309), .A2(new_n250), .ZN(new_n368));
  AOI21_X1  g0168(.A(new_n367), .B1(new_n368), .B2(G226), .ZN(new_n369));
  NAND3_X1  g0169(.A1(new_n249), .A2(G223), .A3(new_n250), .ZN(new_n370));
  AOI21_X1  g0170(.A(new_n364), .B1(new_n369), .B2(new_n370), .ZN(new_n371));
  AOI21_X1  g0171(.A(new_n260), .B1(new_n265), .B2(G232), .ZN(new_n372));
  INV_X1    g0172(.A(new_n372), .ZN(new_n373));
  OAI21_X1  g0173(.A(new_n361), .B1(new_n371), .B2(new_n373), .ZN(new_n374));
  INV_X1    g0174(.A(G226), .ZN(new_n375));
  OAI22_X1  g0175(.A1(new_n253), .A2(new_n375), .B1(new_n365), .B2(new_n366), .ZN(new_n376));
  INV_X1    g0176(.A(new_n370), .ZN(new_n377));
  OAI21_X1  g0177(.A(new_n256), .B1(new_n376), .B2(new_n377), .ZN(new_n378));
  NAND3_X1  g0178(.A1(new_n378), .A2(new_n269), .A3(new_n372), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n374), .A2(new_n379), .ZN(new_n380));
  OAI21_X1  g0180(.A(KEYINPUT18), .B1(new_n360), .B2(new_n380), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n353), .A2(G68), .ZN(new_n382));
  INV_X1    g0182(.A(new_n345), .ZN(new_n383));
  NAND3_X1  g0183(.A1(new_n382), .A2(KEYINPUT16), .A3(new_n383), .ZN(new_n384));
  NAND3_X1  g0184(.A1(new_n384), .A2(new_n272), .A3(new_n359), .ZN(new_n385));
  OAI21_X1  g0185(.A(new_n319), .B1(new_n371), .B2(new_n373), .ZN(new_n386));
  NAND3_X1  g0186(.A1(new_n378), .A2(new_n317), .A3(new_n372), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n386), .A2(new_n387), .ZN(new_n388));
  INV_X1    g0188(.A(new_n339), .ZN(new_n389));
  NAND3_X1  g0189(.A1(new_n385), .A2(new_n388), .A3(new_n389), .ZN(new_n390));
  INV_X1    g0190(.A(KEYINPUT17), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n390), .A2(new_n391), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n385), .A2(new_n389), .ZN(new_n393));
  INV_X1    g0193(.A(new_n380), .ZN(new_n394));
  INV_X1    g0194(.A(KEYINPUT18), .ZN(new_n395));
  NAND3_X1  g0195(.A1(new_n393), .A2(new_n394), .A3(new_n395), .ZN(new_n396));
  NAND3_X1  g0196(.A1(new_n360), .A2(KEYINPUT17), .A3(new_n388), .ZN(new_n397));
  NAND4_X1  g0197(.A1(new_n381), .A2(new_n392), .A3(new_n396), .A4(new_n397), .ZN(new_n398));
  NOR2_X1   g0198(.A1(new_n335), .A2(new_n398), .ZN(new_n399));
  OAI21_X1  g0199(.A(KEYINPUT12), .B1(new_n302), .B2(G68), .ZN(new_n400));
  AND2_X1   g0200(.A1(new_n400), .A2(KEYINPUT71), .ZN(new_n401));
  NOR2_X1   g0201(.A1(new_n400), .A2(KEYINPUT71), .ZN(new_n402));
  NOR3_X1   g0202(.A1(new_n282), .A2(KEYINPUT12), .A3(G68), .ZN(new_n403));
  NOR3_X1   g0203(.A1(new_n401), .A2(new_n402), .A3(new_n403), .ZN(new_n404));
  OAI22_X1  g0204(.A1(new_n290), .A2(new_n202), .B1(new_n212), .B2(G68), .ZN(new_n405));
  NOR2_X1   g0205(.A1(new_n275), .A2(new_n252), .ZN(new_n406));
  OAI21_X1  g0206(.A(new_n272), .B1(new_n405), .B2(new_n406), .ZN(new_n407));
  XNOR2_X1  g0207(.A(new_n407), .B(KEYINPUT11), .ZN(new_n408));
  NAND3_X1  g0208(.A1(new_n299), .A2(G68), .A3(new_n300), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n408), .A2(new_n409), .ZN(new_n410));
  NOR2_X1   g0210(.A1(new_n404), .A2(new_n410), .ZN(new_n411));
  INV_X1    g0211(.A(new_n411), .ZN(new_n412));
  INV_X1    g0212(.A(KEYINPUT69), .ZN(new_n413));
  AOI221_X4 g0213(.A(new_n413), .B1(new_n362), .B2(new_n363), .C1(new_n261), .C2(new_n264), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n261), .A2(new_n264), .ZN(new_n415));
  AOI21_X1  g0215(.A(KEYINPUT69), .B1(new_n415), .B2(new_n364), .ZN(new_n416));
  OAI21_X1  g0216(.A(G238), .B1(new_n414), .B2(new_n416), .ZN(new_n417));
  INV_X1    g0217(.A(new_n260), .ZN(new_n418));
  NAND3_X1  g0218(.A1(new_n417), .A2(KEYINPUT70), .A3(new_n418), .ZN(new_n419));
  AOI22_X1  g0219(.A1(new_n368), .A2(G232), .B1(G33), .B2(G97), .ZN(new_n420));
  NAND3_X1  g0220(.A1(new_n249), .A2(G226), .A3(new_n250), .ZN(new_n421));
  AOI21_X1  g0221(.A(new_n364), .B1(new_n420), .B2(new_n421), .ZN(new_n422));
  INV_X1    g0222(.A(new_n422), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n419), .A2(new_n423), .ZN(new_n424));
  AOI21_X1  g0224(.A(KEYINPUT70), .B1(new_n417), .B2(new_n418), .ZN(new_n425));
  OAI21_X1  g0225(.A(KEYINPUT13), .B1(new_n424), .B2(new_n425), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n417), .A2(new_n418), .ZN(new_n427));
  INV_X1    g0227(.A(KEYINPUT70), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n427), .A2(new_n428), .ZN(new_n429));
  INV_X1    g0229(.A(KEYINPUT13), .ZN(new_n430));
  NAND4_X1  g0230(.A1(new_n429), .A2(new_n430), .A3(new_n419), .A4(new_n423), .ZN(new_n431));
  NAND3_X1  g0231(.A1(new_n426), .A2(G179), .A3(new_n431), .ZN(new_n432));
  AOI21_X1  g0232(.A(new_n361), .B1(new_n426), .B2(new_n431), .ZN(new_n433));
  INV_X1    g0233(.A(KEYINPUT14), .ZN(new_n434));
  OAI21_X1  g0234(.A(new_n432), .B1(new_n433), .B2(new_n434), .ZN(new_n435));
  AOI211_X1 g0235(.A(KEYINPUT14), .B(new_n361), .C1(new_n426), .C2(new_n431), .ZN(new_n436));
  OAI21_X1  g0236(.A(new_n412), .B1(new_n435), .B2(new_n436), .ZN(new_n437));
  NAND3_X1  g0237(.A1(new_n426), .A2(new_n317), .A3(new_n431), .ZN(new_n438));
  INV_X1    g0238(.A(new_n438), .ZN(new_n439));
  AOI21_X1  g0239(.A(G200), .B1(new_n426), .B2(new_n431), .ZN(new_n440));
  OAI21_X1  g0240(.A(new_n411), .B1(new_n439), .B2(new_n440), .ZN(new_n441));
  NAND3_X1  g0241(.A1(new_n399), .A2(new_n437), .A3(new_n441), .ZN(new_n442));
  INV_X1    g0242(.A(new_n442), .ZN(new_n443));
  INV_X1    g0243(.A(G45), .ZN(new_n444));
  OAI21_X1  g0244(.A(G250), .B1(new_n444), .B2(G1), .ZN(new_n445));
  NOR2_X1   g0245(.A1(new_n444), .A2(G1), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n446), .A2(G274), .ZN(new_n447));
  AOI21_X1  g0247(.A(new_n256), .B1(new_n445), .B2(new_n447), .ZN(new_n448));
  OAI211_X1 g0248(.A(G244), .B(G1698), .C1(new_n307), .C2(new_n308), .ZN(new_n449));
  OAI211_X1 g0249(.A(G238), .B(new_n250), .C1(new_n307), .C2(new_n308), .ZN(new_n450));
  NAND2_X1  g0250(.A1(G33), .A2(G116), .ZN(new_n451));
  NAND3_X1  g0251(.A1(new_n449), .A2(new_n450), .A3(new_n451), .ZN(new_n452));
  AOI21_X1  g0252(.A(new_n448), .B1(new_n452), .B2(new_n256), .ZN(new_n453));
  OAI21_X1  g0253(.A(KEYINPUT78), .B1(new_n453), .B2(G169), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n453), .A2(new_n269), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n454), .A2(new_n455), .ZN(new_n456));
  INV_X1    g0256(.A(KEYINPUT79), .ZN(new_n457));
  NAND3_X1  g0257(.A1(new_n453), .A2(KEYINPUT78), .A3(new_n269), .ZN(new_n458));
  AND3_X1   g0258(.A1(new_n456), .A2(new_n457), .A3(new_n458), .ZN(new_n459));
  AOI21_X1  g0259(.A(new_n457), .B1(new_n456), .B2(new_n458), .ZN(new_n460));
  NOR2_X1   g0260(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  NAND3_X1  g0261(.A1(KEYINPUT19), .A2(G33), .A3(G97), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n462), .A2(new_n212), .ZN(new_n463));
  NOR2_X1   g0263(.A1(G87), .A2(G97), .ZN(new_n464));
  INV_X1    g0264(.A(G107), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  NAND3_X1  g0266(.A1(new_n212), .A2(G33), .A3(G97), .ZN(new_n467));
  INV_X1    g0267(.A(KEYINPUT19), .ZN(new_n468));
  AOI22_X1  g0268(.A1(new_n463), .A2(new_n466), .B1(new_n467), .B2(new_n468), .ZN(new_n469));
  NAND3_X1  g0269(.A1(new_n249), .A2(new_n212), .A3(G68), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n469), .A2(new_n470), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n471), .A2(new_n272), .ZN(new_n472));
  NAND2_X1  g0272(.A1(new_n303), .A2(new_n291), .ZN(new_n473));
  NAND3_X1  g0273(.A1(new_n472), .A2(KEYINPUT80), .A3(new_n473), .ZN(new_n474));
  INV_X1    g0274(.A(KEYINPUT80), .ZN(new_n475));
  AOI21_X1  g0275(.A(new_n273), .B1(new_n469), .B2(new_n470), .ZN(new_n476));
  INV_X1    g0276(.A(new_n291), .ZN(new_n477));
  NOR2_X1   g0277(.A1(new_n302), .A2(new_n477), .ZN(new_n478));
  OAI21_X1  g0278(.A(new_n475), .B1(new_n476), .B2(new_n478), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n474), .A2(new_n479), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n263), .A2(G33), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n284), .A2(new_n481), .ZN(new_n482));
  INV_X1    g0282(.A(new_n482), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n483), .A2(new_n477), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n480), .A2(new_n484), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n485), .A2(KEYINPUT81), .ZN(new_n486));
  INV_X1    g0286(.A(KEYINPUT81), .ZN(new_n487));
  NAND3_X1  g0287(.A1(new_n480), .A2(new_n487), .A3(new_n484), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n486), .A2(new_n488), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n483), .A2(G87), .ZN(new_n490));
  OAI211_X1 g0290(.A(new_n480), .B(new_n490), .C1(new_n319), .C2(new_n453), .ZN(new_n491));
  INV_X1    g0291(.A(new_n491), .ZN(new_n492));
  AND2_X1   g0292(.A1(new_n453), .A2(G190), .ZN(new_n493));
  XOR2_X1   g0293(.A(new_n493), .B(KEYINPUT82), .Z(new_n494));
  AOI22_X1  g0294(.A1(new_n461), .A2(new_n489), .B1(new_n492), .B2(new_n494), .ZN(new_n495));
  NOR2_X1   g0295(.A1(new_n482), .A2(new_n465), .ZN(new_n496));
  NAND3_X1  g0296(.A1(new_n295), .A2(G20), .A3(new_n465), .ZN(new_n497));
  XNOR2_X1  g0297(.A(new_n497), .B(KEYINPUT25), .ZN(new_n498));
  NOR2_X1   g0298(.A1(new_n496), .A2(new_n498), .ZN(new_n499));
  INV_X1    g0299(.A(new_n499), .ZN(new_n500));
  OAI211_X1 g0300(.A(new_n212), .B(G87), .C1(new_n307), .C2(new_n308), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n501), .A2(KEYINPUT83), .ZN(new_n502));
  INV_X1    g0302(.A(KEYINPUT83), .ZN(new_n503));
  NAND4_X1  g0303(.A1(new_n249), .A2(new_n503), .A3(new_n212), .A4(G87), .ZN(new_n504));
  NAND3_X1  g0304(.A1(new_n502), .A2(new_n504), .A3(KEYINPUT22), .ZN(new_n505));
  INV_X1    g0305(.A(KEYINPUT22), .ZN(new_n506));
  NAND3_X1  g0306(.A1(new_n501), .A2(KEYINPUT83), .A3(new_n506), .ZN(new_n507));
  INV_X1    g0307(.A(KEYINPUT23), .ZN(new_n508));
  AOI21_X1  g0308(.A(new_n508), .B1(G20), .B2(new_n465), .ZN(new_n509));
  NOR3_X1   g0309(.A1(new_n212), .A2(KEYINPUT23), .A3(G107), .ZN(new_n510));
  NOR2_X1   g0310(.A1(new_n451), .A2(G20), .ZN(new_n511));
  NOR3_X1   g0311(.A1(new_n509), .A2(new_n510), .A3(new_n511), .ZN(new_n512));
  NAND4_X1  g0312(.A1(new_n505), .A2(KEYINPUT24), .A3(new_n507), .A4(new_n512), .ZN(new_n513));
  AND2_X1   g0313(.A1(new_n513), .A2(new_n272), .ZN(new_n514));
  NAND3_X1  g0314(.A1(new_n505), .A2(new_n507), .A3(new_n512), .ZN(new_n515));
  INV_X1    g0315(.A(KEYINPUT24), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  AOI21_X1  g0317(.A(new_n500), .B1(new_n514), .B2(new_n517), .ZN(new_n518));
  OAI211_X1 g0318(.A(G250), .B(new_n250), .C1(new_n307), .C2(new_n308), .ZN(new_n519));
  OAI211_X1 g0319(.A(G257), .B(G1698), .C1(new_n307), .C2(new_n308), .ZN(new_n520));
  INV_X1    g0320(.A(G294), .ZN(new_n521));
  OAI211_X1 g0321(.A(new_n519), .B(new_n520), .C1(new_n365), .C2(new_n521), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n522), .A2(new_n256), .ZN(new_n523));
  INV_X1    g0323(.A(KEYINPUT5), .ZN(new_n524));
  INV_X1    g0324(.A(KEYINPUT76), .ZN(new_n525));
  OAI21_X1  g0325(.A(new_n524), .B1(new_n525), .B2(G41), .ZN(new_n526));
  INV_X1    g0326(.A(G41), .ZN(new_n527));
  NAND3_X1  g0327(.A1(new_n527), .A2(KEYINPUT76), .A3(KEYINPUT5), .ZN(new_n528));
  NAND3_X1  g0328(.A1(new_n526), .A2(new_n446), .A3(new_n528), .ZN(new_n529));
  NAND3_X1  g0329(.A1(new_n529), .A2(new_n364), .A3(G264), .ZN(new_n530));
  INV_X1    g0330(.A(KEYINPUT84), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n530), .A2(new_n531), .ZN(new_n532));
  NAND4_X1  g0332(.A1(new_n529), .A2(new_n364), .A3(KEYINPUT84), .A4(G264), .ZN(new_n533));
  NAND4_X1  g0333(.A1(new_n526), .A2(new_n528), .A3(new_n446), .A4(G274), .ZN(new_n534));
  NAND4_X1  g0334(.A1(new_n523), .A2(new_n532), .A3(new_n533), .A4(new_n534), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n535), .A2(new_n319), .ZN(new_n536));
  OAI21_X1  g0336(.A(new_n536), .B1(G190), .B2(new_n535), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n518), .A2(new_n537), .ZN(new_n538));
  NAND3_X1  g0338(.A1(new_n517), .A2(new_n272), .A3(new_n513), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n539), .A2(new_n499), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n535), .A2(G169), .ZN(new_n541));
  AOI22_X1  g0341(.A1(new_n522), .A2(new_n256), .B1(new_n530), .B2(new_n531), .ZN(new_n542));
  NAND4_X1  g0342(.A1(new_n542), .A2(G179), .A3(new_n533), .A4(new_n534), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n541), .A2(new_n543), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n540), .A2(new_n544), .ZN(new_n545));
  AND2_X1   g0345(.A1(new_n538), .A2(new_n545), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n365), .A2(G97), .ZN(new_n547));
  NAND2_X1  g0347(.A1(G33), .A2(G283), .ZN(new_n548));
  AOI21_X1  g0348(.A(G20), .B1(new_n547), .B2(new_n548), .ZN(new_n549));
  INV_X1    g0349(.A(G116), .ZN(new_n550));
  NOR2_X1   g0350(.A1(new_n212), .A2(new_n550), .ZN(new_n551));
  OAI21_X1  g0351(.A(new_n272), .B1(new_n549), .B2(new_n551), .ZN(new_n552));
  INV_X1    g0352(.A(KEYINPUT20), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n552), .A2(new_n553), .ZN(new_n554));
  OAI211_X1 g0354(.A(KEYINPUT20), .B(new_n272), .C1(new_n549), .C2(new_n551), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n303), .A2(new_n550), .ZN(new_n557));
  NAND4_X1  g0357(.A1(new_n302), .A2(G116), .A3(new_n273), .A4(new_n481), .ZN(new_n558));
  NAND3_X1  g0358(.A1(new_n556), .A2(new_n557), .A3(new_n558), .ZN(new_n559));
  INV_X1    g0359(.A(new_n559), .ZN(new_n560));
  NAND3_X1  g0360(.A1(new_n529), .A2(new_n364), .A3(G270), .ZN(new_n561));
  AND2_X1   g0361(.A1(new_n561), .A2(new_n534), .ZN(new_n562));
  OAI211_X1 g0362(.A(G264), .B(G1698), .C1(new_n307), .C2(new_n308), .ZN(new_n563));
  OAI211_X1 g0363(.A(G257), .B(new_n250), .C1(new_n307), .C2(new_n308), .ZN(new_n564));
  INV_X1    g0364(.A(G303), .ZN(new_n565));
  OAI211_X1 g0365(.A(new_n563), .B(new_n564), .C1(new_n565), .C2(new_n249), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n566), .A2(new_n256), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n562), .A2(new_n567), .ZN(new_n568));
  NAND3_X1  g0368(.A1(new_n568), .A2(KEYINPUT21), .A3(G169), .ZN(new_n569));
  NAND3_X1  g0369(.A1(new_n562), .A2(new_n567), .A3(G179), .ZN(new_n570));
  AOI21_X1  g0370(.A(new_n560), .B1(new_n569), .B2(new_n570), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n568), .A2(new_n319), .ZN(new_n572));
  NAND3_X1  g0372(.A1(new_n562), .A2(new_n567), .A3(new_n317), .ZN(new_n573));
  AOI21_X1  g0373(.A(new_n559), .B1(new_n572), .B2(new_n573), .ZN(new_n574));
  AOI21_X1  g0374(.A(new_n361), .B1(new_n562), .B2(new_n567), .ZN(new_n575));
  AOI21_X1  g0375(.A(KEYINPUT21), .B1(new_n559), .B2(new_n575), .ZN(new_n576));
  NOR3_X1   g0376(.A1(new_n571), .A2(new_n574), .A3(new_n576), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n348), .A2(new_n357), .ZN(new_n578));
  AOI22_X1  g0378(.A1(new_n578), .A2(G107), .B1(G77), .B2(new_n277), .ZN(new_n579));
  XNOR2_X1  g0379(.A(KEYINPUT73), .B(G107), .ZN(new_n580));
  INV_X1    g0380(.A(new_n580), .ZN(new_n581));
  INV_X1    g0381(.A(G97), .ZN(new_n582));
  NAND3_X1  g0382(.A1(new_n582), .A2(new_n465), .A3(KEYINPUT6), .ZN(new_n583));
  OR2_X1    g0383(.A1(new_n582), .A2(KEYINPUT6), .ZN(new_n584));
  NAND3_X1  g0384(.A1(new_n581), .A2(new_n583), .A3(new_n584), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n584), .A2(new_n583), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n586), .A2(new_n580), .ZN(new_n587));
  NAND3_X1  g0387(.A1(new_n585), .A2(new_n587), .A3(G20), .ZN(new_n588));
  AOI21_X1  g0388(.A(new_n273), .B1(new_n579), .B2(new_n588), .ZN(new_n589));
  NOR2_X1   g0389(.A1(new_n282), .A2(G97), .ZN(new_n590));
  AOI21_X1  g0390(.A(new_n590), .B1(new_n483), .B2(G97), .ZN(new_n591));
  INV_X1    g0391(.A(new_n591), .ZN(new_n592));
  OAI21_X1  g0392(.A(KEYINPUT77), .B1(new_n589), .B2(new_n592), .ZN(new_n593));
  OAI211_X1 g0393(.A(G244), .B(new_n250), .C1(new_n307), .C2(new_n308), .ZN(new_n594));
  INV_X1    g0394(.A(KEYINPUT74), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n594), .A2(new_n595), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n596), .A2(KEYINPUT4), .ZN(new_n597));
  INV_X1    g0397(.A(KEYINPUT4), .ZN(new_n598));
  NAND3_X1  g0398(.A1(new_n594), .A2(new_n595), .A3(new_n598), .ZN(new_n599));
  AND2_X1   g0399(.A1(new_n597), .A2(new_n599), .ZN(new_n600));
  OAI211_X1 g0400(.A(G250), .B(G1698), .C1(new_n307), .C2(new_n308), .ZN(new_n601));
  INV_X1    g0401(.A(KEYINPUT75), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n601), .A2(new_n602), .ZN(new_n603));
  NAND4_X1  g0403(.A1(new_n249), .A2(KEYINPUT75), .A3(G250), .A4(G1698), .ZN(new_n604));
  AOI22_X1  g0404(.A1(new_n603), .A2(new_n604), .B1(G33), .B2(G283), .ZN(new_n605));
  AOI21_X1  g0405(.A(new_n364), .B1(new_n600), .B2(new_n605), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n529), .A2(new_n364), .ZN(new_n607));
  INV_X1    g0407(.A(G257), .ZN(new_n608));
  OAI21_X1  g0408(.A(new_n534), .B1(new_n607), .B2(new_n608), .ZN(new_n609));
  OAI21_X1  g0409(.A(new_n361), .B1(new_n606), .B2(new_n609), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n578), .A2(G107), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n277), .A2(G77), .ZN(new_n612));
  NAND3_X1  g0412(.A1(new_n611), .A2(new_n588), .A3(new_n612), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n613), .A2(new_n272), .ZN(new_n614));
  INV_X1    g0414(.A(KEYINPUT77), .ZN(new_n615));
  NAND3_X1  g0415(.A1(new_n614), .A2(new_n615), .A3(new_n591), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n603), .A2(new_n604), .ZN(new_n617));
  NAND4_X1  g0417(.A1(new_n617), .A2(new_n597), .A3(new_n548), .A4(new_n599), .ZN(new_n618));
  AOI21_X1  g0418(.A(new_n609), .B1(new_n618), .B2(new_n256), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n619), .A2(new_n269), .ZN(new_n620));
  NAND4_X1  g0420(.A1(new_n593), .A2(new_n610), .A3(new_n616), .A4(new_n620), .ZN(new_n621));
  NOR2_X1   g0421(.A1(new_n589), .A2(new_n592), .ZN(new_n622));
  NOR2_X1   g0422(.A1(new_n619), .A2(G200), .ZN(new_n623));
  AOI211_X1 g0423(.A(G190), .B(new_n609), .C1(new_n618), .C2(new_n256), .ZN(new_n624));
  OAI21_X1  g0424(.A(new_n622), .B1(new_n623), .B2(new_n624), .ZN(new_n625));
  AND3_X1   g0425(.A1(new_n577), .A2(new_n621), .A3(new_n625), .ZN(new_n626));
  AND4_X1   g0426(.A1(new_n443), .A2(new_n495), .A3(new_n546), .A4(new_n626), .ZN(G372));
  AND2_X1   g0427(.A1(new_n381), .A2(new_n396), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n415), .A2(new_n364), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n629), .A2(new_n413), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n265), .A2(KEYINPUT69), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n630), .A2(new_n631), .ZN(new_n632));
  AOI21_X1  g0432(.A(new_n260), .B1(new_n632), .B2(G238), .ZN(new_n633));
  AOI21_X1  g0433(.A(new_n422), .B1(new_n633), .B2(KEYINPUT70), .ZN(new_n634));
  AOI21_X1  g0434(.A(new_n430), .B1(new_n634), .B2(new_n429), .ZN(new_n635));
  NOR3_X1   g0435(.A1(new_n424), .A2(KEYINPUT13), .A3(new_n425), .ZN(new_n636));
  OAI21_X1  g0436(.A(G169), .B1(new_n635), .B2(new_n636), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n637), .A2(KEYINPUT14), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n433), .A2(new_n434), .ZN(new_n639));
  NAND3_X1  g0439(.A1(new_n638), .A2(new_n639), .A3(new_n432), .ZN(new_n640));
  AOI21_X1  g0440(.A(new_n325), .B1(new_n640), .B2(new_n412), .ZN(new_n641));
  NAND3_X1  g0441(.A1(new_n441), .A2(new_n392), .A3(new_n397), .ZN(new_n642));
  OAI21_X1  g0442(.A(new_n628), .B1(new_n641), .B2(new_n642), .ZN(new_n643));
  NOR2_X1   g0443(.A1(new_n333), .A2(new_n334), .ZN(new_n644));
  INV_X1    g0444(.A(new_n644), .ZN(new_n645));
  AOI22_X1  g0445(.A1(new_n643), .A2(new_n645), .B1(new_n287), .B2(new_n270), .ZN(new_n646));
  INV_X1    g0446(.A(KEYINPUT26), .ZN(new_n647));
  INV_X1    g0447(.A(new_n621), .ZN(new_n648));
  AOI21_X1  g0448(.A(new_n647), .B1(new_n495), .B2(new_n648), .ZN(new_n649));
  NOR2_X1   g0449(.A1(new_n453), .A2(G169), .ZN(new_n650));
  AOI21_X1  g0450(.A(new_n650), .B1(new_n269), .B2(new_n453), .ZN(new_n651));
  AND3_X1   g0451(.A1(new_n480), .A2(new_n487), .A3(new_n484), .ZN(new_n652));
  AOI21_X1  g0452(.A(new_n487), .B1(new_n480), .B2(new_n484), .ZN(new_n653));
  OAI21_X1  g0453(.A(new_n651), .B1(new_n652), .B2(new_n653), .ZN(new_n654));
  NOR2_X1   g0454(.A1(new_n491), .A2(new_n493), .ZN(new_n655));
  INV_X1    g0455(.A(new_n655), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n614), .A2(new_n591), .ZN(new_n657));
  AND3_X1   g0457(.A1(new_n610), .A2(new_n657), .A3(new_n620), .ZN(new_n658));
  NAND4_X1  g0458(.A1(new_n656), .A2(new_n654), .A3(new_n658), .A4(new_n647), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n569), .A2(new_n570), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n660), .A2(new_n559), .ZN(new_n661));
  INV_X1    g0461(.A(new_n576), .ZN(new_n662));
  AND2_X1   g0462(.A1(new_n541), .A2(new_n543), .ZN(new_n663));
  OAI211_X1 g0463(.A(new_n661), .B(new_n662), .C1(new_n518), .C2(new_n663), .ZN(new_n664));
  NAND4_X1  g0464(.A1(new_n664), .A2(new_n538), .A3(new_n625), .A4(new_n621), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n656), .A2(new_n654), .ZN(new_n666));
  OAI211_X1 g0466(.A(new_n654), .B(new_n659), .C1(new_n665), .C2(new_n666), .ZN(new_n667));
  OAI21_X1  g0467(.A(new_n443), .B1(new_n649), .B2(new_n667), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n646), .A2(new_n668), .ZN(new_n669));
  XNOR2_X1  g0469(.A(new_n669), .B(KEYINPUT85), .ZN(G369));
  NAND2_X1  g0470(.A1(new_n661), .A2(new_n662), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n295), .A2(new_n212), .ZN(new_n672));
  OR2_X1    g0472(.A1(new_n672), .A2(KEYINPUT27), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n672), .A2(KEYINPUT27), .ZN(new_n674));
  NAND3_X1  g0474(.A1(new_n673), .A2(G213), .A3(new_n674), .ZN(new_n675));
  INV_X1    g0475(.A(G343), .ZN(new_n676));
  NOR2_X1   g0476(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  INV_X1    g0477(.A(new_n677), .ZN(new_n678));
  NOR2_X1   g0478(.A1(new_n560), .A2(new_n678), .ZN(new_n679));
  MUX2_X1   g0479(.A(new_n577), .B(new_n671), .S(new_n679), .Z(new_n680));
  INV_X1    g0480(.A(new_n545), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n681), .A2(new_n677), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n540), .A2(new_n677), .ZN(new_n683));
  NAND3_X1  g0483(.A1(new_n545), .A2(new_n538), .A3(new_n683), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n682), .A2(new_n684), .ZN(new_n685));
  NAND3_X1  g0485(.A1(new_n680), .A2(new_n685), .A3(G330), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n681), .A2(new_n678), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n671), .A2(new_n678), .ZN(new_n688));
  OAI21_X1  g0488(.A(new_n687), .B1(new_n684), .B2(new_n688), .ZN(new_n689));
  INV_X1    g0489(.A(new_n689), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n686), .A2(new_n690), .ZN(G399));
  INV_X1    g0491(.A(new_n208), .ZN(new_n692));
  NOR2_X1   g0492(.A1(new_n692), .A2(G41), .ZN(new_n693));
  INV_X1    g0493(.A(new_n693), .ZN(new_n694));
  OAI21_X1  g0494(.A(KEYINPUT86), .B1(new_n694), .B2(new_n215), .ZN(new_n695));
  NAND3_X1  g0495(.A1(new_n464), .A2(new_n465), .A3(new_n550), .ZN(new_n696));
  NOR3_X1   g0496(.A1(new_n693), .A2(new_n263), .A3(new_n696), .ZN(new_n697));
  MUX2_X1   g0497(.A(new_n695), .B(KEYINPUT86), .S(new_n697), .Z(new_n698));
  XNOR2_X1  g0498(.A(new_n698), .B(KEYINPUT28), .ZN(new_n699));
  INV_X1    g0499(.A(G330), .ZN(new_n700));
  NOR2_X1   g0500(.A1(new_n453), .A2(G179), .ZN(new_n701));
  NAND3_X1  g0501(.A1(new_n701), .A2(new_n535), .A3(new_n568), .ZN(new_n702));
  NOR2_X1   g0502(.A1(new_n702), .A2(new_n619), .ZN(new_n703));
  NAND3_X1  g0503(.A1(new_n542), .A2(new_n453), .A3(new_n533), .ZN(new_n704));
  NOR2_X1   g0504(.A1(new_n704), .A2(new_n570), .ZN(new_n705));
  NAND2_X1  g0505(.A1(new_n705), .A2(new_n619), .ZN(new_n706));
  INV_X1    g0506(.A(KEYINPUT87), .ZN(new_n707));
  OR2_X1    g0507(.A1(new_n707), .A2(KEYINPUT30), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n706), .A2(new_n708), .ZN(new_n709));
  NOR2_X1   g0509(.A1(new_n707), .A2(KEYINPUT30), .ZN(new_n710));
  NAND3_X1  g0510(.A1(new_n705), .A2(new_n619), .A3(new_n710), .ZN(new_n711));
  AOI21_X1  g0511(.A(new_n703), .B1(new_n709), .B2(new_n711), .ZN(new_n712));
  INV_X1    g0512(.A(KEYINPUT31), .ZN(new_n713));
  NOR3_X1   g0513(.A1(new_n712), .A2(new_n713), .A3(new_n678), .ZN(new_n714));
  AND3_X1   g0514(.A1(new_n705), .A2(new_n619), .A3(new_n710), .ZN(new_n715));
  AOI21_X1  g0515(.A(new_n710), .B1(new_n705), .B2(new_n619), .ZN(new_n716));
  OAI22_X1  g0516(.A1(new_n715), .A2(new_n716), .B1(new_n619), .B2(new_n702), .ZN(new_n717));
  AOI21_X1  g0517(.A(KEYINPUT31), .B1(new_n717), .B2(new_n677), .ZN(new_n718));
  NOR2_X1   g0518(.A1(new_n714), .A2(new_n718), .ZN(new_n719));
  NAND4_X1  g0519(.A1(new_n626), .A2(new_n495), .A3(new_n546), .A4(new_n678), .ZN(new_n720));
  AOI21_X1  g0520(.A(new_n700), .B1(new_n719), .B2(new_n720), .ZN(new_n721));
  INV_X1    g0521(.A(KEYINPUT88), .ZN(new_n722));
  OAI21_X1  g0522(.A(new_n722), .B1(new_n665), .B2(new_n666), .ZN(new_n723));
  AND3_X1   g0523(.A1(new_n621), .A2(new_n538), .A3(new_n625), .ZN(new_n724));
  AOI21_X1  g0524(.A(new_n655), .B1(new_n489), .B2(new_n651), .ZN(new_n725));
  NAND4_X1  g0525(.A1(new_n724), .A2(new_n725), .A3(KEYINPUT88), .A4(new_n664), .ZN(new_n726));
  INV_X1    g0526(.A(new_n654), .ZN(new_n727));
  NAND3_X1  g0527(.A1(new_n656), .A2(new_n654), .A3(new_n658), .ZN(new_n728));
  AOI21_X1  g0528(.A(new_n727), .B1(new_n728), .B2(KEYINPUT26), .ZN(new_n729));
  NAND3_X1  g0529(.A1(new_n495), .A2(new_n647), .A3(new_n648), .ZN(new_n730));
  NAND4_X1  g0530(.A1(new_n723), .A2(new_n726), .A3(new_n729), .A4(new_n730), .ZN(new_n731));
  NAND3_X1  g0531(.A1(new_n731), .A2(KEYINPUT29), .A3(new_n678), .ZN(new_n732));
  OAI21_X1  g0532(.A(new_n678), .B1(new_n667), .B2(new_n649), .ZN(new_n733));
  INV_X1    g0533(.A(KEYINPUT29), .ZN(new_n734));
  NAND2_X1  g0534(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  AOI21_X1  g0535(.A(new_n721), .B1(new_n732), .B2(new_n735), .ZN(new_n736));
  OAI21_X1  g0536(.A(new_n699), .B1(new_n736), .B2(G1), .ZN(G364));
  NOR2_X1   g0537(.A1(new_n294), .A2(G20), .ZN(new_n738));
  NAND2_X1  g0538(.A1(new_n738), .A2(G45), .ZN(new_n739));
  NOR2_X1   g0539(.A1(new_n739), .A2(KEYINPUT89), .ZN(new_n740));
  NOR2_X1   g0540(.A1(new_n740), .A2(new_n263), .ZN(new_n741));
  NAND2_X1  g0541(.A1(new_n739), .A2(KEYINPUT89), .ZN(new_n742));
  NAND2_X1  g0542(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  NOR2_X1   g0543(.A1(new_n693), .A2(new_n743), .ZN(new_n744));
  NOR2_X1   g0544(.A1(G13), .A2(G33), .ZN(new_n745));
  INV_X1    g0545(.A(new_n745), .ZN(new_n746));
  NOR2_X1   g0546(.A1(new_n746), .A2(G20), .ZN(new_n747));
  AOI21_X1  g0547(.A(new_n211), .B1(G20), .B2(new_n361), .ZN(new_n748));
  NOR2_X1   g0548(.A1(new_n747), .A2(new_n748), .ZN(new_n749));
  INV_X1    g0549(.A(new_n749), .ZN(new_n750));
  NAND3_X1  g0550(.A1(new_n208), .A2(G355), .A3(new_n249), .ZN(new_n751));
  OAI21_X1  g0551(.A(new_n751), .B1(G116), .B2(new_n208), .ZN(new_n752));
  NOR2_X1   g0552(.A1(new_n692), .A2(new_n249), .ZN(new_n753));
  NAND2_X1  g0553(.A1(new_n242), .A2(G45), .ZN(new_n754));
  OAI21_X1  g0554(.A(new_n754), .B1(G45), .B2(new_n216), .ZN(new_n755));
  AOI21_X1  g0555(.A(new_n752), .B1(new_n753), .B2(new_n755), .ZN(new_n756));
  NOR2_X1   g0556(.A1(new_n212), .A2(G190), .ZN(new_n757));
  XNOR2_X1  g0557(.A(new_n757), .B(KEYINPUT90), .ZN(new_n758));
  NOR3_X1   g0558(.A1(new_n758), .A2(G179), .A3(G200), .ZN(new_n759));
  XOR2_X1   g0559(.A(KEYINPUT91), .B(G159), .Z(new_n760));
  INV_X1    g0560(.A(new_n760), .ZN(new_n761));
  NAND2_X1  g0561(.A1(new_n759), .A2(new_n761), .ZN(new_n762));
  XNOR2_X1  g0562(.A(new_n762), .B(KEYINPUT32), .ZN(new_n763));
  NOR2_X1   g0563(.A1(G179), .A2(G200), .ZN(new_n764));
  AOI21_X1  g0564(.A(new_n212), .B1(new_n764), .B2(G190), .ZN(new_n765));
  NOR2_X1   g0565(.A1(new_n765), .A2(new_n582), .ZN(new_n766));
  NOR2_X1   g0566(.A1(new_n212), .A2(new_n317), .ZN(new_n767));
  NOR2_X1   g0567(.A1(new_n269), .A2(new_n319), .ZN(new_n768));
  NAND2_X1  g0568(.A1(new_n767), .A2(new_n768), .ZN(new_n769));
  NOR2_X1   g0569(.A1(new_n269), .A2(G200), .ZN(new_n770));
  NAND2_X1  g0570(.A1(new_n767), .A2(new_n770), .ZN(new_n771));
  OAI22_X1  g0571(.A1(new_n769), .A2(new_n202), .B1(new_n771), .B2(new_n340), .ZN(new_n772));
  NAND2_X1  g0572(.A1(new_n768), .A2(new_n757), .ZN(new_n773));
  NAND2_X1  g0573(.A1(new_n757), .A2(new_n770), .ZN(new_n774));
  OAI22_X1  g0574(.A1(new_n773), .A2(new_n341), .B1(new_n774), .B2(new_n252), .ZN(new_n775));
  NOR4_X1   g0575(.A1(new_n763), .A2(new_n766), .A3(new_n772), .A4(new_n775), .ZN(new_n776));
  NOR3_X1   g0576(.A1(new_n758), .A2(G179), .A3(new_n319), .ZN(new_n777));
  NAND2_X1  g0577(.A1(new_n777), .A2(G107), .ZN(new_n778));
  NAND3_X1  g0578(.A1(new_n767), .A2(new_n269), .A3(G200), .ZN(new_n779));
  OR2_X1    g0579(.A1(new_n779), .A2(KEYINPUT92), .ZN(new_n780));
  NAND2_X1  g0580(.A1(new_n779), .A2(KEYINPUT92), .ZN(new_n781));
  NAND2_X1  g0581(.A1(new_n780), .A2(new_n781), .ZN(new_n782));
  OAI211_X1 g0582(.A(new_n778), .B(new_n249), .C1(new_n366), .C2(new_n782), .ZN(new_n783));
  XNOR2_X1  g0583(.A(new_n783), .B(KEYINPUT93), .ZN(new_n784));
  INV_X1    g0584(.A(new_n777), .ZN(new_n785));
  INV_X1    g0585(.A(G283), .ZN(new_n786));
  NOR2_X1   g0586(.A1(new_n785), .A2(new_n786), .ZN(new_n787));
  INV_X1    g0587(.A(G311), .ZN(new_n788));
  OAI221_X1 g0588(.A(new_n309), .B1(new_n788), .B2(new_n774), .C1(new_n782), .C2(new_n565), .ZN(new_n789));
  AOI211_X1 g0589(.A(new_n787), .B(new_n789), .C1(G329), .C2(new_n759), .ZN(new_n790));
  XOR2_X1   g0590(.A(KEYINPUT33), .B(G317), .Z(new_n791));
  INV_X1    g0591(.A(G322), .ZN(new_n792));
  OAI22_X1  g0592(.A1(new_n791), .A2(new_n773), .B1(new_n771), .B2(new_n792), .ZN(new_n793));
  XNOR2_X1  g0593(.A(new_n793), .B(KEYINPUT95), .ZN(new_n794));
  INV_X1    g0594(.A(G326), .ZN(new_n795));
  OAI22_X1  g0595(.A1(new_n769), .A2(new_n795), .B1(new_n765), .B2(new_n521), .ZN(new_n796));
  INV_X1    g0596(.A(KEYINPUT94), .ZN(new_n797));
  OR2_X1    g0597(.A1(new_n796), .A2(new_n797), .ZN(new_n798));
  NAND2_X1  g0598(.A1(new_n796), .A2(new_n797), .ZN(new_n799));
  NAND3_X1  g0599(.A1(new_n794), .A2(new_n798), .A3(new_n799), .ZN(new_n800));
  INV_X1    g0600(.A(new_n800), .ZN(new_n801));
  AOI22_X1  g0601(.A1(new_n776), .A2(new_n784), .B1(new_n790), .B2(new_n801), .ZN(new_n802));
  INV_X1    g0602(.A(new_n748), .ZN(new_n803));
  OAI221_X1 g0603(.A(new_n744), .B1(new_n750), .B2(new_n756), .C1(new_n802), .C2(new_n803), .ZN(new_n804));
  INV_X1    g0604(.A(new_n747), .ZN(new_n805));
  NOR2_X1   g0605(.A1(new_n680), .A2(new_n805), .ZN(new_n806));
  NOR2_X1   g0606(.A1(new_n804), .A2(new_n806), .ZN(new_n807));
  XOR2_X1   g0607(.A(new_n807), .B(KEYINPUT96), .Z(new_n808));
  NOR2_X1   g0608(.A1(new_n680), .A2(G330), .ZN(new_n809));
  NAND2_X1  g0609(.A1(new_n680), .A2(G330), .ZN(new_n810));
  INV_X1    g0610(.A(new_n744), .ZN(new_n811));
  NAND2_X1  g0611(.A1(new_n810), .A2(new_n811), .ZN(new_n812));
  OAI21_X1  g0612(.A(new_n808), .B1(new_n809), .B2(new_n812), .ZN(G396));
  OAI21_X1  g0613(.A(new_n324), .B1(new_n269), .B2(new_n315), .ZN(new_n814));
  NAND2_X1  g0614(.A1(new_n814), .A2(new_n305), .ZN(new_n815));
  NOR2_X1   g0615(.A1(new_n322), .A2(new_n678), .ZN(new_n816));
  OAI21_X1  g0616(.A(new_n815), .B1(new_n321), .B2(new_n816), .ZN(new_n817));
  INV_X1    g0617(.A(KEYINPUT99), .ZN(new_n818));
  NAND2_X1  g0618(.A1(new_n325), .A2(new_n678), .ZN(new_n819));
  AND3_X1   g0619(.A1(new_n817), .A2(new_n818), .A3(new_n819), .ZN(new_n820));
  AOI21_X1  g0620(.A(new_n818), .B1(new_n817), .B2(new_n819), .ZN(new_n821));
  OR2_X1    g0621(.A1(new_n820), .A2(new_n821), .ZN(new_n822));
  NAND2_X1  g0622(.A1(new_n733), .A2(new_n822), .ZN(new_n823));
  NOR2_X1   g0623(.A1(new_n820), .A2(new_n821), .ZN(new_n824));
  OAI211_X1 g0624(.A(new_n824), .B(new_n678), .C1(new_n667), .C2(new_n649), .ZN(new_n825));
  NAND2_X1  g0625(.A1(new_n823), .A2(new_n825), .ZN(new_n826));
  INV_X1    g0626(.A(new_n721), .ZN(new_n827));
  OAI21_X1  g0627(.A(new_n811), .B1(new_n826), .B2(new_n827), .ZN(new_n828));
  INV_X1    g0628(.A(new_n828), .ZN(new_n829));
  NAND2_X1  g0629(.A1(new_n826), .A2(new_n827), .ZN(new_n830));
  NAND2_X1  g0630(.A1(new_n822), .A2(new_n745), .ZN(new_n831));
  NOR2_X1   g0631(.A1(new_n748), .A2(new_n745), .ZN(new_n832));
  INV_X1    g0632(.A(new_n832), .ZN(new_n833));
  OAI21_X1  g0633(.A(new_n744), .B1(G77), .B2(new_n833), .ZN(new_n834));
  AOI22_X1  g0634(.A1(G87), .A2(new_n777), .B1(new_n759), .B2(G311), .ZN(new_n835));
  OAI22_X1  g0635(.A1(new_n773), .A2(new_n786), .B1(new_n774), .B2(new_n550), .ZN(new_n836));
  INV_X1    g0636(.A(new_n771), .ZN(new_n837));
  AOI21_X1  g0637(.A(new_n836), .B1(G294), .B2(new_n837), .ZN(new_n838));
  INV_X1    g0638(.A(new_n782), .ZN(new_n839));
  NAND2_X1  g0639(.A1(new_n839), .A2(G107), .ZN(new_n840));
  INV_X1    g0640(.A(new_n769), .ZN(new_n841));
  AOI211_X1 g0641(.A(new_n249), .B(new_n766), .C1(G303), .C2(new_n841), .ZN(new_n842));
  NAND4_X1  g0642(.A1(new_n835), .A2(new_n838), .A3(new_n840), .A4(new_n842), .ZN(new_n843));
  AOI21_X1  g0643(.A(new_n309), .B1(new_n759), .B2(G132), .ZN(new_n844));
  XOR2_X1   g0644(.A(new_n844), .B(KEYINPUT98), .Z(new_n845));
  INV_X1    g0645(.A(new_n773), .ZN(new_n846));
  AOI22_X1  g0646(.A1(G143), .A2(new_n837), .B1(new_n846), .B2(G150), .ZN(new_n847));
  INV_X1    g0647(.A(G137), .ZN(new_n848));
  OAI221_X1 g0648(.A(new_n847), .B1(new_n848), .B2(new_n769), .C1(new_n774), .C2(new_n760), .ZN(new_n849));
  INV_X1    g0649(.A(KEYINPUT34), .ZN(new_n850));
  INV_X1    g0650(.A(new_n765), .ZN(new_n851));
  AOI22_X1  g0651(.A1(new_n849), .A2(new_n850), .B1(G58), .B2(new_n851), .ZN(new_n852));
  OAI211_X1 g0652(.A(new_n845), .B(new_n852), .C1(new_n850), .C2(new_n849), .ZN(new_n853));
  NAND2_X1  g0653(.A1(new_n777), .A2(G68), .ZN(new_n854));
  OAI21_X1  g0654(.A(new_n854), .B1(new_n202), .B2(new_n782), .ZN(new_n855));
  XNOR2_X1  g0655(.A(new_n855), .B(KEYINPUT97), .ZN(new_n856));
  OAI21_X1  g0656(.A(new_n843), .B1(new_n853), .B2(new_n856), .ZN(new_n857));
  AOI21_X1  g0657(.A(new_n834), .B1(new_n857), .B2(new_n748), .ZN(new_n858));
  AOI22_X1  g0658(.A1(new_n829), .A2(new_n830), .B1(new_n831), .B2(new_n858), .ZN(new_n859));
  INV_X1    g0659(.A(new_n859), .ZN(G384));
  NOR2_X1   g0660(.A1(new_n738), .A2(new_n263), .ZN(new_n861));
  NAND3_X1  g0661(.A1(new_n443), .A2(new_n732), .A3(new_n735), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n646), .A2(new_n862), .ZN(new_n863));
  XOR2_X1   g0663(.A(new_n863), .B(KEYINPUT102), .Z(new_n864));
  OAI21_X1  g0664(.A(new_n355), .B1(KEYINPUT16), .B2(new_n354), .ZN(new_n865));
  AOI21_X1  g0665(.A(new_n675), .B1(new_n865), .B2(new_n389), .ZN(new_n866));
  NAND2_X1  g0666(.A1(new_n398), .A2(new_n866), .ZN(new_n867));
  AOI22_X1  g0667(.A1(new_n865), .A2(new_n389), .B1(new_n380), .B2(new_n675), .ZN(new_n868));
  INV_X1    g0668(.A(new_n390), .ZN(new_n869));
  OAI21_X1  g0669(.A(KEYINPUT37), .B1(new_n868), .B2(new_n869), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n393), .A2(new_n394), .ZN(new_n871));
  INV_X1    g0671(.A(new_n675), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n393), .A2(new_n872), .ZN(new_n873));
  INV_X1    g0673(.A(KEYINPUT37), .ZN(new_n874));
  NAND4_X1  g0674(.A1(new_n871), .A2(new_n873), .A3(new_n874), .A4(new_n390), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n870), .A2(new_n875), .ZN(new_n876));
  NAND3_X1  g0676(.A1(new_n867), .A2(new_n876), .A3(KEYINPUT38), .ZN(new_n877));
  INV_X1    g0677(.A(new_n877), .ZN(new_n878));
  AOI21_X1  g0678(.A(KEYINPUT38), .B1(new_n867), .B2(new_n876), .ZN(new_n879));
  OAI21_X1  g0679(.A(KEYINPUT39), .B1(new_n878), .B2(new_n879), .ZN(new_n880));
  OAI21_X1  g0680(.A(new_n390), .B1(new_n360), .B2(new_n380), .ZN(new_n881));
  NOR2_X1   g0681(.A1(new_n360), .A2(new_n675), .ZN(new_n882));
  OAI21_X1  g0682(.A(KEYINPUT37), .B1(new_n881), .B2(new_n882), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n883), .A2(new_n875), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n398), .A2(new_n882), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n884), .A2(new_n885), .ZN(new_n886));
  INV_X1    g0686(.A(KEYINPUT38), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n886), .A2(new_n887), .ZN(new_n888));
  INV_X1    g0688(.A(KEYINPUT39), .ZN(new_n889));
  NAND3_X1  g0689(.A1(new_n888), .A2(new_n889), .A3(new_n877), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n880), .A2(new_n890), .ZN(new_n891));
  NAND3_X1  g0691(.A1(new_n640), .A2(new_n412), .A3(new_n678), .ZN(new_n892));
  INV_X1    g0692(.A(new_n892), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n891), .A2(new_n893), .ZN(new_n894));
  OAI21_X1  g0694(.A(new_n894), .B1(new_n628), .B2(new_n872), .ZN(new_n895));
  INV_X1    g0695(.A(new_n440), .ZN(new_n896));
  AOI21_X1  g0696(.A(new_n412), .B1(new_n896), .B2(new_n438), .ZN(new_n897));
  OAI211_X1 g0697(.A(new_n412), .B(new_n677), .C1(new_n640), .C2(new_n897), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n412), .A2(new_n677), .ZN(new_n899));
  NAND3_X1  g0699(.A1(new_n437), .A2(new_n441), .A3(new_n899), .ZN(new_n900));
  AOI22_X1  g0700(.A1(new_n825), .A2(new_n819), .B1(new_n898), .B2(new_n900), .ZN(new_n901));
  XNOR2_X1  g0701(.A(new_n901), .B(KEYINPUT101), .ZN(new_n902));
  INV_X1    g0702(.A(new_n879), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n903), .A2(new_n877), .ZN(new_n904));
  AOI21_X1  g0704(.A(new_n895), .B1(new_n902), .B2(new_n904), .ZN(new_n905));
  XNOR2_X1  g0705(.A(new_n864), .B(new_n905), .ZN(new_n906));
  AOI21_X1  g0706(.A(new_n822), .B1(new_n898), .B2(new_n900), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n719), .A2(new_n720), .ZN(new_n908));
  NAND3_X1  g0708(.A1(new_n907), .A2(new_n908), .A3(new_n904), .ZN(new_n909));
  INV_X1    g0709(.A(KEYINPUT40), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n909), .A2(new_n910), .ZN(new_n911));
  AOI221_X4 g0711(.A(new_n822), .B1(new_n720), .B2(new_n719), .C1(new_n898), .C2(new_n900), .ZN(new_n912));
  AOI21_X1  g0712(.A(new_n910), .B1(new_n888), .B2(new_n877), .ZN(new_n913));
  AOI21_X1  g0713(.A(KEYINPUT103), .B1(new_n912), .B2(new_n913), .ZN(new_n914));
  AND4_X1   g0714(.A1(KEYINPUT103), .A2(new_n913), .A3(new_n907), .A4(new_n908), .ZN(new_n915));
  OAI211_X1 g0715(.A(G330), .B(new_n911), .C1(new_n914), .C2(new_n915), .ZN(new_n916));
  OAI21_X1  g0716(.A(new_n916), .B1(new_n442), .B2(new_n827), .ZN(new_n917));
  INV_X1    g0717(.A(KEYINPUT103), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n898), .A2(new_n900), .ZN(new_n919));
  NAND3_X1  g0719(.A1(new_n919), .A2(new_n908), .A3(new_n824), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n888), .A2(new_n877), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n921), .A2(KEYINPUT40), .ZN(new_n922));
  OAI21_X1  g0722(.A(new_n918), .B1(new_n920), .B2(new_n922), .ZN(new_n923));
  NAND4_X1  g0723(.A1(new_n913), .A2(new_n907), .A3(KEYINPUT103), .A4(new_n908), .ZN(new_n924));
  AOI22_X1  g0724(.A1(new_n923), .A2(new_n924), .B1(new_n910), .B2(new_n909), .ZN(new_n925));
  NAND3_X1  g0725(.A1(new_n925), .A2(new_n443), .A3(new_n908), .ZN(new_n926));
  NAND2_X1  g0726(.A1(new_n917), .A2(new_n926), .ZN(new_n927));
  AOI21_X1  g0727(.A(new_n861), .B1(new_n906), .B2(new_n927), .ZN(new_n928));
  OAI21_X1  g0728(.A(new_n928), .B1(new_n906), .B2(new_n927), .ZN(new_n929));
  NOR3_X1   g0729(.A1(new_n215), .A2(new_n252), .A3(new_n342), .ZN(new_n930));
  NOR2_X1   g0730(.A1(new_n341), .A2(G50), .ZN(new_n931));
  XOR2_X1   g0731(.A(new_n931), .B(KEYINPUT100), .Z(new_n932));
  OAI211_X1 g0732(.A(G1), .B(new_n294), .C1(new_n930), .C2(new_n932), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n585), .A2(new_n587), .ZN(new_n934));
  INV_X1    g0734(.A(KEYINPUT35), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n934), .A2(new_n935), .ZN(new_n936));
  NAND3_X1  g0736(.A1(new_n585), .A2(new_n587), .A3(KEYINPUT35), .ZN(new_n937));
  NAND4_X1  g0737(.A1(new_n936), .A2(G116), .A3(new_n213), .A4(new_n937), .ZN(new_n938));
  XNOR2_X1  g0738(.A(new_n938), .B(KEYINPUT36), .ZN(new_n939));
  NAND3_X1  g0739(.A1(new_n929), .A2(new_n933), .A3(new_n939), .ZN(G367));
  INV_X1    g0740(.A(new_n686), .ZN(new_n941));
  NAND2_X1  g0741(.A1(new_n658), .A2(new_n677), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n621), .A2(new_n625), .ZN(new_n943));
  NOR2_X1   g0743(.A1(new_n622), .A2(new_n678), .ZN(new_n944));
  OAI21_X1  g0744(.A(new_n942), .B1(new_n943), .B2(new_n944), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n941), .A2(new_n945), .ZN(new_n946));
  XNOR2_X1  g0746(.A(new_n946), .B(KEYINPUT105), .ZN(new_n947));
  AOI21_X1  g0747(.A(new_n678), .B1(new_n480), .B2(new_n490), .ZN(new_n948));
  NOR2_X1   g0748(.A1(new_n666), .A2(new_n948), .ZN(new_n949));
  NAND2_X1  g0749(.A1(new_n727), .A2(new_n948), .ZN(new_n950));
  AOI21_X1  g0750(.A(new_n949), .B1(KEYINPUT104), .B2(new_n950), .ZN(new_n951));
  OAI21_X1  g0751(.A(new_n951), .B1(KEYINPUT104), .B2(new_n950), .ZN(new_n952));
  NOR2_X1   g0752(.A1(new_n952), .A2(KEYINPUT43), .ZN(new_n953));
  XNOR2_X1  g0753(.A(new_n947), .B(new_n953), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n952), .A2(KEYINPUT43), .ZN(new_n955));
  AOI21_X1  g0755(.A(new_n648), .B1(new_n945), .B2(new_n681), .ZN(new_n956));
  NOR3_X1   g0756(.A1(new_n684), .A2(new_n943), .A3(new_n688), .ZN(new_n957));
  INV_X1    g0757(.A(KEYINPUT42), .ZN(new_n958));
  OAI22_X1  g0758(.A1(new_n956), .A2(new_n677), .B1(new_n957), .B2(new_n958), .ZN(new_n959));
  INV_X1    g0759(.A(new_n957), .ZN(new_n960));
  NOR2_X1   g0760(.A1(new_n960), .A2(KEYINPUT42), .ZN(new_n961));
  OAI21_X1  g0761(.A(new_n955), .B1(new_n959), .B2(new_n961), .ZN(new_n962));
  XNOR2_X1  g0762(.A(new_n954), .B(new_n962), .ZN(new_n963));
  NOR2_X1   g0763(.A1(new_n684), .A2(new_n688), .ZN(new_n964));
  INV_X1    g0764(.A(new_n685), .ZN(new_n965));
  NAND2_X1  g0765(.A1(new_n810), .A2(new_n965), .ZN(new_n966));
  NAND2_X1  g0766(.A1(new_n966), .A2(new_n686), .ZN(new_n967));
  AOI21_X1  g0767(.A(new_n964), .B1(new_n967), .B2(new_n688), .ZN(new_n968));
  AND3_X1   g0768(.A1(new_n736), .A2(KEYINPUT106), .A3(new_n968), .ZN(new_n969));
  AOI21_X1  g0769(.A(KEYINPUT106), .B1(new_n736), .B2(new_n968), .ZN(new_n970));
  OAI21_X1  g0770(.A(KEYINPUT107), .B1(new_n969), .B2(new_n970), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n732), .A2(new_n735), .ZN(new_n972));
  NAND3_X1  g0772(.A1(new_n972), .A2(new_n968), .A3(new_n827), .ZN(new_n973));
  INV_X1    g0773(.A(KEYINPUT106), .ZN(new_n974));
  NAND2_X1  g0774(.A1(new_n973), .A2(new_n974), .ZN(new_n975));
  INV_X1    g0775(.A(KEYINPUT107), .ZN(new_n976));
  NAND3_X1  g0776(.A1(new_n736), .A2(KEYINPUT106), .A3(new_n968), .ZN(new_n977));
  NAND3_X1  g0777(.A1(new_n975), .A2(new_n976), .A3(new_n977), .ZN(new_n978));
  INV_X1    g0778(.A(new_n945), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n979), .A2(new_n689), .ZN(new_n980));
  NAND2_X1  g0780(.A1(new_n980), .A2(KEYINPUT44), .ZN(new_n981));
  INV_X1    g0781(.A(KEYINPUT44), .ZN(new_n982));
  NAND3_X1  g0782(.A1(new_n979), .A2(new_n982), .A3(new_n689), .ZN(new_n983));
  AND2_X1   g0783(.A1(new_n981), .A2(new_n983), .ZN(new_n984));
  INV_X1    g0784(.A(KEYINPUT45), .ZN(new_n985));
  OAI21_X1  g0785(.A(new_n985), .B1(new_n979), .B2(new_n689), .ZN(new_n986));
  NAND3_X1  g0786(.A1(new_n690), .A2(KEYINPUT45), .A3(new_n945), .ZN(new_n987));
  NAND2_X1  g0787(.A1(new_n986), .A2(new_n987), .ZN(new_n988));
  NAND4_X1  g0788(.A1(new_n984), .A2(KEYINPUT108), .A3(new_n686), .A4(new_n988), .ZN(new_n989));
  NAND4_X1  g0789(.A1(new_n988), .A2(new_n981), .A3(new_n686), .A4(new_n983), .ZN(new_n990));
  INV_X1    g0790(.A(KEYINPUT108), .ZN(new_n991));
  NAND2_X1  g0791(.A1(new_n990), .A2(new_n991), .ZN(new_n992));
  NAND2_X1  g0792(.A1(new_n989), .A2(new_n992), .ZN(new_n993));
  NAND2_X1  g0793(.A1(new_n984), .A2(new_n988), .ZN(new_n994));
  NAND2_X1  g0794(.A1(new_n994), .A2(new_n941), .ZN(new_n995));
  AND2_X1   g0795(.A1(new_n993), .A2(new_n995), .ZN(new_n996));
  NAND3_X1  g0796(.A1(new_n971), .A2(new_n978), .A3(new_n996), .ZN(new_n997));
  NAND2_X1  g0797(.A1(new_n997), .A2(new_n736), .ZN(new_n998));
  XOR2_X1   g0798(.A(new_n693), .B(KEYINPUT41), .Z(new_n999));
  INV_X1    g0799(.A(new_n999), .ZN(new_n1000));
  NAND3_X1  g0800(.A1(new_n998), .A2(KEYINPUT109), .A3(new_n1000), .ZN(new_n1001));
  INV_X1    g0801(.A(new_n743), .ZN(new_n1002));
  NAND2_X1  g0802(.A1(new_n1001), .A2(new_n1002), .ZN(new_n1003));
  AOI21_X1  g0803(.A(new_n999), .B1(new_n997), .B2(new_n736), .ZN(new_n1004));
  NOR2_X1   g0804(.A1(new_n1004), .A2(KEYINPUT109), .ZN(new_n1005));
  OAI21_X1  g0805(.A(new_n963), .B1(new_n1003), .B2(new_n1005), .ZN(new_n1006));
  OR2_X1    g0806(.A1(new_n952), .A2(new_n805), .ZN(new_n1007));
  INV_X1    g0807(.A(new_n753), .ZN(new_n1008));
  NOR2_X1   g0808(.A1(new_n1008), .A2(new_n238), .ZN(new_n1009));
  OAI21_X1  g0809(.A(new_n749), .B1(new_n208), .B2(new_n291), .ZN(new_n1010));
  OAI21_X1  g0810(.A(new_n744), .B1(new_n1009), .B2(new_n1010), .ZN(new_n1011));
  AOI22_X1  g0811(.A1(new_n839), .A2(G58), .B1(new_n759), .B2(G137), .ZN(new_n1012));
  OAI21_X1  g0812(.A(new_n1012), .B1(new_n252), .B2(new_n785), .ZN(new_n1013));
  OAI22_X1  g0813(.A1(new_n760), .A2(new_n773), .B1(new_n774), .B2(new_n202), .ZN(new_n1014));
  XNOR2_X1  g0814(.A(new_n1014), .B(KEYINPUT111), .ZN(new_n1015));
  NOR2_X1   g0815(.A1(new_n765), .A2(new_n341), .ZN(new_n1016));
  AOI21_X1  g0816(.A(new_n309), .B1(new_n841), .B2(G143), .ZN(new_n1017));
  INV_X1    g0817(.A(G150), .ZN(new_n1018));
  OAI21_X1  g0818(.A(new_n1017), .B1(new_n1018), .B2(new_n771), .ZN(new_n1019));
  NOR4_X1   g0819(.A1(new_n1013), .A2(new_n1015), .A3(new_n1016), .A4(new_n1019), .ZN(new_n1020));
  NAND2_X1  g0820(.A1(new_n839), .A2(G116), .ZN(new_n1021));
  INV_X1    g0821(.A(KEYINPUT46), .ZN(new_n1022));
  OAI22_X1  g0822(.A1(new_n1021), .A2(new_n1022), .B1(new_n521), .B2(new_n773), .ZN(new_n1023));
  AOI21_X1  g0823(.A(new_n1023), .B1(new_n1022), .B2(new_n1021), .ZN(new_n1024));
  XOR2_X1   g0824(.A(new_n1024), .B(KEYINPUT110), .Z(new_n1025));
  INV_X1    g0825(.A(new_n774), .ZN(new_n1026));
  AOI21_X1  g0826(.A(new_n249), .B1(new_n1026), .B2(G283), .ZN(new_n1027));
  OAI221_X1 g0827(.A(new_n1027), .B1(new_n565), .B2(new_n771), .C1(new_n788), .C2(new_n769), .ZN(new_n1028));
  NAND2_X1  g0828(.A1(new_n777), .A2(G97), .ZN(new_n1029));
  INV_X1    g0829(.A(new_n759), .ZN(new_n1030));
  INV_X1    g0830(.A(G317), .ZN(new_n1031));
  OAI21_X1  g0831(.A(new_n1029), .B1(new_n1030), .B2(new_n1031), .ZN(new_n1032));
  AOI211_X1 g0832(.A(new_n1028), .B(new_n1032), .C1(G107), .C2(new_n851), .ZN(new_n1033));
  AOI21_X1  g0833(.A(new_n1020), .B1(new_n1025), .B2(new_n1033), .ZN(new_n1034));
  OR2_X1    g0834(.A1(new_n1034), .A2(KEYINPUT47), .ZN(new_n1035));
  AOI21_X1  g0835(.A(new_n803), .B1(new_n1034), .B2(KEYINPUT47), .ZN(new_n1036));
  AOI21_X1  g0836(.A(new_n1011), .B1(new_n1035), .B2(new_n1036), .ZN(new_n1037));
  NAND2_X1  g0837(.A1(new_n1007), .A2(new_n1037), .ZN(new_n1038));
  NAND2_X1  g0838(.A1(new_n1006), .A2(new_n1038), .ZN(G387));
  NAND2_X1  g0839(.A1(new_n975), .A2(new_n977), .ZN(new_n1040));
  OAI211_X1 g0840(.A(new_n1040), .B(new_n693), .C1(new_n736), .C2(new_n968), .ZN(new_n1041));
  OAI21_X1  g0841(.A(new_n309), .B1(new_n785), .B2(new_n550), .ZN(new_n1042));
  OAI22_X1  g0842(.A1(new_n782), .A2(new_n521), .B1(new_n786), .B2(new_n765), .ZN(new_n1043));
  NOR2_X1   g0843(.A1(new_n774), .A2(new_n565), .ZN(new_n1044));
  OAI22_X1  g0844(.A1(new_n788), .A2(new_n773), .B1(new_n771), .B2(new_n1031), .ZN(new_n1045));
  AOI211_X1 g0845(.A(new_n1044), .B(new_n1045), .C1(G322), .C2(new_n841), .ZN(new_n1046));
  AOI21_X1  g0846(.A(new_n1043), .B1(new_n1046), .B2(KEYINPUT48), .ZN(new_n1047));
  XOR2_X1   g0847(.A(new_n1047), .B(KEYINPUT112), .Z(new_n1048));
  OAI21_X1  g0848(.A(new_n1048), .B1(KEYINPUT48), .B2(new_n1046), .ZN(new_n1049));
  XOR2_X1   g0849(.A(new_n1049), .B(KEYINPUT49), .Z(new_n1050));
  AOI211_X1 g0850(.A(new_n1042), .B(new_n1050), .C1(G326), .C2(new_n759), .ZN(new_n1051));
  NAND2_X1  g0851(.A1(new_n839), .A2(G77), .ZN(new_n1052));
  OAI211_X1 g0852(.A(new_n1052), .B(new_n1029), .C1(new_n1018), .C2(new_n1030), .ZN(new_n1053));
  AOI22_X1  g0853(.A1(new_n841), .A2(G159), .B1(new_n846), .B2(new_n337), .ZN(new_n1054));
  OAI21_X1  g0854(.A(new_n1054), .B1(new_n341), .B2(new_n774), .ZN(new_n1055));
  NOR2_X1   g0855(.A1(new_n765), .A2(new_n291), .ZN(new_n1056));
  OAI21_X1  g0856(.A(new_n249), .B1(new_n771), .B2(new_n202), .ZN(new_n1057));
  NOR4_X1   g0857(.A1(new_n1053), .A2(new_n1055), .A3(new_n1056), .A4(new_n1057), .ZN(new_n1058));
  OAI21_X1  g0858(.A(new_n748), .B1(new_n1051), .B2(new_n1058), .ZN(new_n1059));
  NAND3_X1  g0859(.A1(new_n235), .A2(G45), .A3(new_n309), .ZN(new_n1060));
  NAND3_X1  g0860(.A1(new_n337), .A2(KEYINPUT50), .A3(new_n202), .ZN(new_n1061));
  INV_X1    g0861(.A(KEYINPUT50), .ZN(new_n1062));
  OAI21_X1  g0862(.A(new_n1062), .B1(new_n274), .B2(G50), .ZN(new_n1063));
  NAND2_X1  g0863(.A1(new_n1061), .A2(new_n1063), .ZN(new_n1064));
  AOI21_X1  g0864(.A(G45), .B1(G68), .B2(G77), .ZN(new_n1065));
  AOI21_X1  g0865(.A(new_n249), .B1(new_n1064), .B2(new_n1065), .ZN(new_n1066));
  OAI21_X1  g0866(.A(new_n1060), .B1(new_n696), .B2(new_n1066), .ZN(new_n1067));
  NAND2_X1  g0867(.A1(new_n1067), .A2(new_n208), .ZN(new_n1068));
  AOI21_X1  g0868(.A(new_n750), .B1(new_n692), .B2(G107), .ZN(new_n1069));
  AOI21_X1  g0869(.A(new_n811), .B1(new_n1068), .B2(new_n1069), .ZN(new_n1070));
  OAI211_X1 g0870(.A(new_n1059), .B(new_n1070), .C1(new_n685), .C2(new_n805), .ZN(new_n1071));
  NAND2_X1  g0871(.A1(new_n968), .A2(new_n743), .ZN(new_n1072));
  NAND3_X1  g0872(.A1(new_n1041), .A2(new_n1071), .A3(new_n1072), .ZN(G393));
  NOR2_X1   g0873(.A1(new_n1008), .A2(new_n245), .ZN(new_n1074));
  OAI21_X1  g0874(.A(new_n749), .B1(new_n208), .B2(new_n582), .ZN(new_n1075));
  OAI21_X1  g0875(.A(new_n744), .B1(new_n1074), .B2(new_n1075), .ZN(new_n1076));
  AOI22_X1  g0876(.A1(new_n839), .A2(G68), .B1(new_n759), .B2(G143), .ZN(new_n1077));
  AOI21_X1  g0877(.A(new_n309), .B1(new_n851), .B2(G77), .ZN(new_n1078));
  OAI211_X1 g0878(.A(new_n1077), .B(new_n1078), .C1(new_n366), .C2(new_n785), .ZN(new_n1079));
  OAI22_X1  g0879(.A1(new_n773), .A2(new_n202), .B1(new_n774), .B2(new_n274), .ZN(new_n1080));
  XOR2_X1   g0880(.A(new_n1080), .B(KEYINPUT114), .Z(new_n1081));
  INV_X1    g0881(.A(G159), .ZN(new_n1082));
  OAI22_X1  g0882(.A1(new_n769), .A2(new_n1018), .B1(new_n771), .B2(new_n1082), .ZN(new_n1083));
  XNOR2_X1  g0883(.A(new_n1083), .B(KEYINPUT51), .ZN(new_n1084));
  NAND2_X1  g0884(.A1(new_n1081), .A2(new_n1084), .ZN(new_n1085));
  NAND2_X1  g0885(.A1(new_n759), .A2(G322), .ZN(new_n1086));
  OAI22_X1  g0886(.A1(new_n769), .A2(new_n1031), .B1(new_n771), .B2(new_n788), .ZN(new_n1087));
  INV_X1    g0887(.A(KEYINPUT52), .ZN(new_n1088));
  OAI221_X1 g0888(.A(new_n1086), .B1(new_n1087), .B2(new_n1088), .C1(new_n786), .C2(new_n782), .ZN(new_n1089));
  NAND2_X1  g0889(.A1(new_n851), .A2(G116), .ZN(new_n1090));
  OAI21_X1  g0890(.A(new_n309), .B1(new_n773), .B2(new_n565), .ZN(new_n1091));
  AOI21_X1  g0891(.A(new_n1091), .B1(G294), .B2(new_n1026), .ZN(new_n1092));
  NAND2_X1  g0892(.A1(new_n1087), .A2(new_n1088), .ZN(new_n1093));
  NAND4_X1  g0893(.A1(new_n778), .A2(new_n1090), .A3(new_n1092), .A4(new_n1093), .ZN(new_n1094));
  OAI22_X1  g0894(.A1(new_n1079), .A2(new_n1085), .B1(new_n1089), .B2(new_n1094), .ZN(new_n1095));
  AOI21_X1  g0895(.A(new_n1076), .B1(new_n1095), .B2(new_n748), .ZN(new_n1096));
  OAI21_X1  g0896(.A(new_n1096), .B1(new_n945), .B2(new_n805), .ZN(new_n1097));
  XOR2_X1   g0897(.A(new_n995), .B(KEYINPUT113), .Z(new_n1098));
  NAND2_X1  g0898(.A1(new_n1098), .A2(new_n993), .ZN(new_n1099));
  OAI21_X1  g0899(.A(new_n1097), .B1(new_n1099), .B2(new_n1002), .ZN(new_n1100));
  AOI21_X1  g0900(.A(new_n694), .B1(new_n1099), .B2(new_n1040), .ZN(new_n1101));
  AOI21_X1  g0901(.A(new_n1100), .B1(new_n997), .B2(new_n1101), .ZN(new_n1102));
  INV_X1    g0902(.A(new_n1102), .ZN(G390));
  NAND2_X1  g0903(.A1(new_n825), .A2(new_n819), .ZN(new_n1104));
  AOI21_X1  g0904(.A(new_n893), .B1(new_n1104), .B2(new_n919), .ZN(new_n1105));
  NOR2_X1   g0905(.A1(new_n1105), .A2(new_n891), .ZN(new_n1106));
  NAND2_X1  g0906(.A1(new_n921), .A2(new_n892), .ZN(new_n1107));
  NAND3_X1  g0907(.A1(new_n731), .A2(new_n678), .A3(new_n824), .ZN(new_n1108));
  NAND2_X1  g0908(.A1(new_n1108), .A2(new_n819), .ZN(new_n1109));
  AOI21_X1  g0909(.A(new_n1107), .B1(new_n1109), .B2(new_n919), .ZN(new_n1110));
  OAI211_X1 g0910(.A(new_n721), .B(new_n907), .C1(new_n1106), .C2(new_n1110), .ZN(new_n1111));
  INV_X1    g0911(.A(new_n1107), .ZN(new_n1112));
  INV_X1    g0912(.A(new_n1109), .ZN(new_n1113));
  INV_X1    g0913(.A(new_n919), .ZN(new_n1114));
  OAI21_X1  g0914(.A(new_n1112), .B1(new_n1113), .B2(new_n1114), .ZN(new_n1115));
  OAI211_X1 g0915(.A(new_n880), .B(new_n890), .C1(new_n901), .C2(new_n893), .ZN(new_n1116));
  AND3_X1   g0916(.A1(new_n437), .A2(new_n441), .A3(new_n899), .ZN(new_n1117));
  AOI21_X1  g0917(.A(new_n899), .B1(new_n437), .B2(new_n441), .ZN(new_n1118));
  OAI211_X1 g0918(.A(new_n721), .B(new_n824), .C1(new_n1117), .C2(new_n1118), .ZN(new_n1119));
  INV_X1    g0919(.A(KEYINPUT115), .ZN(new_n1120));
  NAND2_X1  g0920(.A1(new_n1119), .A2(new_n1120), .ZN(new_n1121));
  NAND3_X1  g0921(.A1(new_n907), .A2(KEYINPUT115), .A3(new_n721), .ZN(new_n1122));
  NAND4_X1  g0922(.A1(new_n1115), .A2(new_n1116), .A3(new_n1121), .A4(new_n1122), .ZN(new_n1123));
  AND2_X1   g0923(.A1(new_n1111), .A2(new_n1123), .ZN(new_n1124));
  NAND2_X1  g0924(.A1(new_n1124), .A2(new_n743), .ZN(new_n1125));
  AOI21_X1  g0925(.A(new_n811), .B1(new_n274), .B2(new_n832), .ZN(new_n1126));
  INV_X1    g0926(.A(G125), .ZN(new_n1127));
  OAI22_X1  g0927(.A1(new_n202), .A2(new_n785), .B1(new_n1030), .B2(new_n1127), .ZN(new_n1128));
  NAND2_X1  g0928(.A1(new_n837), .A2(G132), .ZN(new_n1129));
  XNOR2_X1  g0929(.A(KEYINPUT54), .B(G143), .ZN(new_n1130));
  OAI221_X1 g0930(.A(new_n1129), .B1(new_n774), .B2(new_n1130), .C1(new_n848), .C2(new_n773), .ZN(new_n1131));
  INV_X1    g0931(.A(G128), .ZN(new_n1132));
  OAI221_X1 g0932(.A(new_n249), .B1(new_n765), .B2(new_n1082), .C1(new_n769), .C2(new_n1132), .ZN(new_n1133));
  NOR3_X1   g0933(.A1(new_n1128), .A2(new_n1131), .A3(new_n1133), .ZN(new_n1134));
  NOR2_X1   g0934(.A1(new_n782), .A2(new_n1018), .ZN(new_n1135));
  XNOR2_X1  g0935(.A(new_n1135), .B(KEYINPUT53), .ZN(new_n1136));
  OAI22_X1  g0936(.A1(new_n769), .A2(new_n786), .B1(new_n774), .B2(new_n582), .ZN(new_n1137));
  AOI21_X1  g0937(.A(new_n1137), .B1(G107), .B2(new_n846), .ZN(new_n1138));
  XNOR2_X1  g0938(.A(new_n1138), .B(KEYINPUT118), .ZN(new_n1139));
  OAI221_X1 g0939(.A(new_n309), .B1(new_n765), .B2(new_n252), .C1(new_n550), .C2(new_n771), .ZN(new_n1140));
  AOI21_X1  g0940(.A(new_n1140), .B1(new_n839), .B2(G87), .ZN(new_n1141));
  NAND2_X1  g0941(.A1(new_n759), .A2(G294), .ZN(new_n1142));
  AND3_X1   g0942(.A1(new_n1141), .A2(new_n854), .A3(new_n1142), .ZN(new_n1143));
  AOI22_X1  g0943(.A1(new_n1134), .A2(new_n1136), .B1(new_n1139), .B2(new_n1143), .ZN(new_n1144));
  OAI221_X1 g0944(.A(new_n1126), .B1(new_n803), .B2(new_n1144), .C1(new_n891), .C2(new_n746), .ZN(new_n1145));
  NAND2_X1  g0945(.A1(new_n1125), .A2(new_n1145), .ZN(new_n1146));
  INV_X1    g0946(.A(KEYINPUT116), .ZN(new_n1147));
  OAI21_X1  g0947(.A(new_n1147), .B1(new_n827), .B2(new_n442), .ZN(new_n1148));
  NAND3_X1  g0948(.A1(new_n443), .A2(KEYINPUT116), .A3(new_n721), .ZN(new_n1149));
  NAND4_X1  g0949(.A1(new_n646), .A2(new_n862), .A3(new_n1148), .A4(new_n1149), .ZN(new_n1150));
  NAND3_X1  g0950(.A1(new_n908), .A2(G330), .A3(new_n824), .ZN(new_n1151));
  NAND3_X1  g0951(.A1(new_n1151), .A2(new_n900), .A3(new_n898), .ZN(new_n1152));
  NAND4_X1  g0952(.A1(new_n1121), .A2(new_n1113), .A3(new_n1122), .A4(new_n1152), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n1152), .A2(new_n1119), .ZN(new_n1154));
  NAND2_X1  g0954(.A1(new_n1154), .A2(new_n1104), .ZN(new_n1155));
  AOI21_X1  g0955(.A(new_n1150), .B1(new_n1153), .B2(new_n1155), .ZN(new_n1156));
  NAND3_X1  g0956(.A1(new_n1156), .A2(new_n1111), .A3(new_n1123), .ZN(new_n1157));
  AND2_X1   g0957(.A1(new_n1157), .A2(new_n693), .ZN(new_n1158));
  OR2_X1    g0958(.A1(new_n1158), .A2(KEYINPUT117), .ZN(new_n1159));
  NOR2_X1   g0959(.A1(new_n1124), .A2(new_n1156), .ZN(new_n1160));
  AOI21_X1  g0960(.A(new_n1160), .B1(new_n1158), .B2(KEYINPUT117), .ZN(new_n1161));
  AOI21_X1  g0961(.A(new_n1146), .B1(new_n1159), .B2(new_n1161), .ZN(new_n1162));
  INV_X1    g0962(.A(new_n1162), .ZN(G378));
  XOR2_X1   g0963(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1164));
  NAND3_X1  g0964(.A1(new_n645), .A2(new_n288), .A3(new_n1164), .ZN(new_n1165));
  INV_X1    g0965(.A(new_n1165), .ZN(new_n1166));
  NAND2_X1  g0966(.A1(new_n287), .A2(new_n872), .ZN(new_n1167));
  XOR2_X1   g0967(.A(new_n1167), .B(KEYINPUT121), .Z(new_n1168));
  INV_X1    g0968(.A(new_n1168), .ZN(new_n1169));
  AOI21_X1  g0969(.A(new_n1164), .B1(new_n645), .B2(new_n288), .ZN(new_n1170));
  OR3_X1    g0970(.A1(new_n1166), .A2(new_n1169), .A3(new_n1170), .ZN(new_n1171));
  OAI21_X1  g0971(.A(new_n1169), .B1(new_n1166), .B2(new_n1170), .ZN(new_n1172));
  NAND2_X1  g0972(.A1(new_n1171), .A2(new_n1172), .ZN(new_n1173));
  INV_X1    g0973(.A(new_n1173), .ZN(new_n1174));
  NAND2_X1  g0974(.A1(new_n916), .A2(new_n1174), .ZN(new_n1175));
  NAND3_X1  g0975(.A1(new_n925), .A2(G330), .A3(new_n1173), .ZN(new_n1176));
  AND3_X1   g0976(.A1(new_n1175), .A2(new_n905), .A3(new_n1176), .ZN(new_n1177));
  AOI21_X1  g0977(.A(new_n905), .B1(new_n1175), .B2(new_n1176), .ZN(new_n1178));
  OAI21_X1  g0978(.A(KEYINPUT122), .B1(new_n1177), .B2(new_n1178), .ZN(new_n1179));
  INV_X1    g0979(.A(new_n1150), .ZN(new_n1180));
  NAND2_X1  g0980(.A1(new_n1157), .A2(new_n1180), .ZN(new_n1181));
  INV_X1    g0981(.A(new_n905), .ZN(new_n1182));
  NOR2_X1   g0982(.A1(new_n916), .A2(new_n1174), .ZN(new_n1183));
  AOI21_X1  g0983(.A(new_n1173), .B1(new_n925), .B2(G330), .ZN(new_n1184));
  OAI21_X1  g0984(.A(new_n1182), .B1(new_n1183), .B2(new_n1184), .ZN(new_n1185));
  INV_X1    g0985(.A(KEYINPUT122), .ZN(new_n1186));
  NAND3_X1  g0986(.A1(new_n1175), .A2(new_n1176), .A3(new_n905), .ZN(new_n1187));
  NAND3_X1  g0987(.A1(new_n1185), .A2(new_n1186), .A3(new_n1187), .ZN(new_n1188));
  NAND3_X1  g0988(.A1(new_n1179), .A2(new_n1181), .A3(new_n1188), .ZN(new_n1189));
  INV_X1    g0989(.A(KEYINPUT57), .ZN(new_n1190));
  NAND2_X1  g0990(.A1(new_n1189), .A2(new_n1190), .ZN(new_n1191));
  AOI21_X1  g0991(.A(new_n1190), .B1(new_n1157), .B2(new_n1180), .ZN(new_n1192));
  NAND3_X1  g0992(.A1(new_n1192), .A2(new_n1185), .A3(new_n1187), .ZN(new_n1193));
  NAND2_X1  g0993(.A1(new_n1193), .A2(new_n693), .ZN(new_n1194));
  INV_X1    g0994(.A(new_n1194), .ZN(new_n1195));
  NAND2_X1  g0995(.A1(new_n1191), .A2(new_n1195), .ZN(new_n1196));
  NAND3_X1  g0996(.A1(new_n1179), .A2(new_n743), .A3(new_n1188), .ZN(new_n1197));
  NOR2_X1   g0997(.A1(new_n1174), .A2(new_n746), .ZN(new_n1198));
  NAND2_X1  g0998(.A1(new_n777), .A2(G58), .ZN(new_n1199));
  XOR2_X1   g0999(.A(new_n1199), .B(KEYINPUT119), .Z(new_n1200));
  NOR2_X1   g1000(.A1(new_n249), .A2(G41), .ZN(new_n1201));
  OAI221_X1 g1001(.A(new_n1201), .B1(new_n582), .B2(new_n773), .C1(new_n550), .C2(new_n769), .ZN(new_n1202));
  OAI22_X1  g1002(.A1(new_n771), .A2(new_n465), .B1(new_n774), .B2(new_n291), .ZN(new_n1203));
  NOR3_X1   g1003(.A1(new_n1202), .A2(new_n1016), .A3(new_n1203), .ZN(new_n1204));
  NAND2_X1  g1004(.A1(new_n759), .A2(G283), .ZN(new_n1205));
  NAND4_X1  g1005(.A1(new_n1200), .A2(new_n1052), .A3(new_n1204), .A4(new_n1205), .ZN(new_n1206));
  XOR2_X1   g1006(.A(new_n1206), .B(KEYINPUT120), .Z(new_n1207));
  NAND2_X1  g1007(.A1(new_n1207), .A2(KEYINPUT58), .ZN(new_n1208));
  AOI211_X1 g1008(.A(G50), .B(new_n1201), .C1(new_n365), .C2(new_n527), .ZN(new_n1209));
  OAI211_X1 g1009(.A(new_n365), .B(new_n527), .C1(new_n785), .C2(new_n760), .ZN(new_n1210));
  INV_X1    g1010(.A(G132), .ZN(new_n1211));
  OAI22_X1  g1011(.A1(new_n773), .A2(new_n1211), .B1(new_n774), .B2(new_n848), .ZN(new_n1212));
  OAI22_X1  g1012(.A1(new_n769), .A2(new_n1127), .B1(new_n771), .B2(new_n1132), .ZN(new_n1213));
  AOI211_X1 g1013(.A(new_n1212), .B(new_n1213), .C1(G150), .C2(new_n851), .ZN(new_n1214));
  OAI21_X1  g1014(.A(new_n1214), .B1(new_n782), .B2(new_n1130), .ZN(new_n1215));
  AND2_X1   g1015(.A1(new_n1215), .A2(KEYINPUT59), .ZN(new_n1216));
  AOI211_X1 g1016(.A(new_n1210), .B(new_n1216), .C1(G124), .C2(new_n759), .ZN(new_n1217));
  OR2_X1    g1017(.A1(new_n1215), .A2(KEYINPUT59), .ZN(new_n1218));
  AOI21_X1  g1018(.A(new_n1209), .B1(new_n1217), .B2(new_n1218), .ZN(new_n1219));
  NAND2_X1  g1019(.A1(new_n1208), .A2(new_n1219), .ZN(new_n1220));
  NOR2_X1   g1020(.A1(new_n1207), .A2(KEYINPUT58), .ZN(new_n1221));
  OAI21_X1  g1021(.A(new_n748), .B1(new_n1220), .B2(new_n1221), .ZN(new_n1222));
  OAI211_X1 g1022(.A(new_n1222), .B(new_n744), .C1(G50), .C2(new_n833), .ZN(new_n1223));
  NOR2_X1   g1023(.A1(new_n1198), .A2(new_n1223), .ZN(new_n1224));
  INV_X1    g1024(.A(new_n1224), .ZN(new_n1225));
  NAND2_X1  g1025(.A1(new_n1197), .A2(new_n1225), .ZN(new_n1226));
  INV_X1    g1026(.A(new_n1226), .ZN(new_n1227));
  NAND2_X1  g1027(.A1(new_n1196), .A2(new_n1227), .ZN(G375));
  NAND2_X1  g1028(.A1(new_n1153), .A2(new_n1155), .ZN(new_n1229));
  NAND2_X1  g1029(.A1(new_n1229), .A2(new_n1180), .ZN(new_n1230));
  NAND3_X1  g1030(.A1(new_n1153), .A2(new_n1150), .A3(new_n1155), .ZN(new_n1231));
  NAND3_X1  g1031(.A1(new_n1230), .A2(new_n1000), .A3(new_n1231), .ZN(new_n1232));
  NAND2_X1  g1032(.A1(new_n1114), .A2(new_n745), .ZN(new_n1233));
  OAI21_X1  g1033(.A(new_n744), .B1(G68), .B2(new_n833), .ZN(new_n1234));
  AOI22_X1  g1034(.A1(G77), .A2(new_n777), .B1(new_n759), .B2(G303), .ZN(new_n1235));
  OAI22_X1  g1035(.A1(new_n773), .A2(new_n550), .B1(new_n774), .B2(new_n465), .ZN(new_n1236));
  AOI21_X1  g1036(.A(new_n1236), .B1(G283), .B2(new_n837), .ZN(new_n1237));
  NAND2_X1  g1037(.A1(new_n839), .A2(G97), .ZN(new_n1238));
  AOI211_X1 g1038(.A(new_n249), .B(new_n1056), .C1(G294), .C2(new_n841), .ZN(new_n1239));
  NAND4_X1  g1039(.A1(new_n1235), .A2(new_n1237), .A3(new_n1238), .A4(new_n1239), .ZN(new_n1240));
  INV_X1    g1040(.A(new_n1200), .ZN(new_n1241));
  OAI22_X1  g1041(.A1(new_n769), .A2(new_n1211), .B1(new_n773), .B2(new_n1130), .ZN(new_n1242));
  OAI221_X1 g1042(.A(new_n249), .B1(new_n765), .B2(new_n202), .C1(new_n848), .C2(new_n771), .ZN(new_n1243));
  AOI211_X1 g1043(.A(new_n1242), .B(new_n1243), .C1(G150), .C2(new_n1026), .ZN(new_n1244));
  OAI221_X1 g1044(.A(new_n1244), .B1(new_n1132), .B2(new_n1030), .C1(new_n1082), .C2(new_n782), .ZN(new_n1245));
  OAI21_X1  g1045(.A(new_n1240), .B1(new_n1241), .B2(new_n1245), .ZN(new_n1246));
  AOI21_X1  g1046(.A(new_n1234), .B1(new_n1246), .B2(new_n748), .ZN(new_n1247));
  AOI22_X1  g1047(.A1(new_n1229), .A2(new_n743), .B1(new_n1233), .B2(new_n1247), .ZN(new_n1248));
  NAND2_X1  g1048(.A1(new_n1232), .A2(new_n1248), .ZN(new_n1249));
  XNOR2_X1  g1049(.A(new_n1249), .B(KEYINPUT123), .ZN(G381));
  NOR2_X1   g1050(.A1(G375), .A2(G378), .ZN(new_n1251));
  NAND3_X1  g1051(.A1(new_n1006), .A2(new_n1038), .A3(new_n1102), .ZN(new_n1252));
  OR2_X1    g1052(.A1(G393), .A2(G396), .ZN(new_n1253));
  NOR4_X1   g1053(.A1(new_n1252), .A2(G381), .A3(G384), .A4(new_n1253), .ZN(new_n1254));
  NAND2_X1  g1054(.A1(new_n1251), .A2(new_n1254), .ZN(G407));
  NAND2_X1  g1055(.A1(new_n676), .A2(G213), .ZN(new_n1256));
  INV_X1    g1056(.A(new_n1256), .ZN(new_n1257));
  NAND2_X1  g1057(.A1(new_n1251), .A2(new_n1257), .ZN(new_n1258));
  NAND3_X1  g1058(.A1(G407), .A2(new_n1258), .A3(G213), .ZN(G409));
  INV_X1    g1059(.A(new_n963), .ZN(new_n1260));
  AOI21_X1  g1060(.A(new_n743), .B1(new_n1004), .B2(KEYINPUT109), .ZN(new_n1261));
  INV_X1    g1061(.A(KEYINPUT109), .ZN(new_n1262));
  INV_X1    g1062(.A(new_n736), .ZN(new_n1263));
  NAND2_X1  g1063(.A1(new_n993), .A2(new_n995), .ZN(new_n1264));
  AOI21_X1  g1064(.A(new_n1264), .B1(new_n1040), .B2(KEYINPUT107), .ZN(new_n1265));
  AOI21_X1  g1065(.A(new_n1263), .B1(new_n1265), .B2(new_n978), .ZN(new_n1266));
  OAI21_X1  g1066(.A(new_n1262), .B1(new_n1266), .B2(new_n999), .ZN(new_n1267));
  AOI21_X1  g1067(.A(new_n1260), .B1(new_n1261), .B2(new_n1267), .ZN(new_n1268));
  INV_X1    g1068(.A(new_n1038), .ZN(new_n1269));
  OAI21_X1  g1069(.A(G390), .B1(new_n1268), .B2(new_n1269), .ZN(new_n1270));
  XNOR2_X1  g1070(.A(G393), .B(G396), .ZN(new_n1271));
  AND3_X1   g1071(.A1(new_n1252), .A2(new_n1270), .A3(new_n1271), .ZN(new_n1272));
  AOI21_X1  g1072(.A(new_n1271), .B1(new_n1252), .B2(new_n1270), .ZN(new_n1273));
  NOR2_X1   g1073(.A1(new_n1272), .A2(new_n1273), .ZN(new_n1274));
  INV_X1    g1074(.A(new_n1274), .ZN(new_n1275));
  INV_X1    g1075(.A(KEYINPUT60), .ZN(new_n1276));
  NAND2_X1  g1076(.A1(new_n1231), .A2(new_n1276), .ZN(new_n1277));
  NAND3_X1  g1077(.A1(new_n1277), .A2(KEYINPUT124), .A3(new_n1230), .ZN(new_n1278));
  NAND4_X1  g1078(.A1(new_n1153), .A2(new_n1150), .A3(new_n1155), .A4(KEYINPUT60), .ZN(new_n1279));
  AND2_X1   g1079(.A1(new_n1279), .A2(new_n693), .ZN(new_n1280));
  NAND2_X1  g1080(.A1(new_n1278), .A2(new_n1280), .ZN(new_n1281));
  AOI21_X1  g1081(.A(KEYINPUT124), .B1(new_n1277), .B2(new_n1230), .ZN(new_n1282));
  OAI21_X1  g1082(.A(new_n1248), .B1(new_n1281), .B2(new_n1282), .ZN(new_n1283));
  NAND2_X1  g1083(.A1(new_n1283), .A2(new_n859), .ZN(new_n1284));
  OAI211_X1 g1084(.A(G384), .B(new_n1248), .C1(new_n1281), .C2(new_n1282), .ZN(new_n1285));
  AND2_X1   g1085(.A1(new_n1284), .A2(new_n1285), .ZN(new_n1286));
  AOI21_X1  g1086(.A(new_n1194), .B1(new_n1189), .B2(new_n1190), .ZN(new_n1287));
  NOR3_X1   g1087(.A1(new_n1287), .A2(new_n1226), .A3(new_n1162), .ZN(new_n1288));
  NAND4_X1  g1088(.A1(new_n1179), .A2(new_n1188), .A3(new_n1000), .A4(new_n1181), .ZN(new_n1289));
  NOR2_X1   g1089(.A1(new_n1177), .A2(new_n1178), .ZN(new_n1290));
  AOI21_X1  g1090(.A(new_n1224), .B1(new_n1290), .B2(new_n743), .ZN(new_n1291));
  NAND2_X1  g1091(.A1(new_n1289), .A2(new_n1291), .ZN(new_n1292));
  AND2_X1   g1092(.A1(new_n1292), .A2(new_n1162), .ZN(new_n1293));
  OAI211_X1 g1093(.A(new_n1256), .B(new_n1286), .C1(new_n1288), .C2(new_n1293), .ZN(new_n1294));
  NAND2_X1  g1094(.A1(new_n1294), .A2(KEYINPUT125), .ZN(new_n1295));
  NAND3_X1  g1095(.A1(new_n1196), .A2(new_n1227), .A3(G378), .ZN(new_n1296));
  NAND2_X1  g1096(.A1(new_n1292), .A2(new_n1162), .ZN(new_n1297));
  NAND2_X1  g1097(.A1(new_n1296), .A2(new_n1297), .ZN(new_n1298));
  INV_X1    g1098(.A(KEYINPUT125), .ZN(new_n1299));
  NAND4_X1  g1099(.A1(new_n1298), .A2(new_n1299), .A3(new_n1256), .A4(new_n1286), .ZN(new_n1300));
  AOI21_X1  g1100(.A(KEYINPUT62), .B1(new_n1295), .B2(new_n1300), .ZN(new_n1301));
  NAND2_X1  g1101(.A1(new_n1294), .A2(KEYINPUT62), .ZN(new_n1302));
  OAI21_X1  g1102(.A(new_n1256), .B1(new_n1288), .B2(new_n1293), .ZN(new_n1303));
  AOI21_X1  g1103(.A(KEYINPUT126), .B1(new_n1284), .B2(new_n1285), .ZN(new_n1304));
  NAND3_X1  g1104(.A1(new_n1284), .A2(KEYINPUT126), .A3(new_n1285), .ZN(new_n1305));
  NAND2_X1  g1105(.A1(new_n1257), .A2(G2897), .ZN(new_n1306));
  INV_X1    g1106(.A(new_n1306), .ZN(new_n1307));
  AOI21_X1  g1107(.A(new_n1304), .B1(new_n1305), .B2(new_n1307), .ZN(new_n1308));
  AOI211_X1 g1108(.A(KEYINPUT126), .B(new_n1306), .C1(new_n1284), .C2(new_n1285), .ZN(new_n1309));
  NOR2_X1   g1109(.A1(new_n1308), .A2(new_n1309), .ZN(new_n1310));
  NAND2_X1  g1110(.A1(new_n1303), .A2(new_n1310), .ZN(new_n1311));
  INV_X1    g1111(.A(KEYINPUT61), .ZN(new_n1312));
  NAND3_X1  g1112(.A1(new_n1302), .A2(new_n1311), .A3(new_n1312), .ZN(new_n1313));
  OAI21_X1  g1113(.A(new_n1275), .B1(new_n1301), .B2(new_n1313), .ZN(new_n1314));
  INV_X1    g1114(.A(KEYINPUT63), .ZN(new_n1315));
  NAND3_X1  g1115(.A1(new_n1295), .A2(new_n1300), .A3(new_n1315), .ZN(new_n1316));
  OR2_X1    g1116(.A1(new_n1294), .A2(new_n1315), .ZN(new_n1317));
  AOI21_X1  g1117(.A(KEYINPUT61), .B1(new_n1303), .B2(new_n1310), .ZN(new_n1318));
  NAND4_X1  g1118(.A1(new_n1316), .A2(new_n1317), .A3(new_n1318), .A4(new_n1274), .ZN(new_n1319));
  NAND2_X1  g1119(.A1(new_n1314), .A2(new_n1319), .ZN(G405));
  OAI21_X1  g1120(.A(new_n1162), .B1(new_n1287), .B2(new_n1226), .ZN(new_n1321));
  INV_X1    g1121(.A(KEYINPUT127), .ZN(new_n1322));
  NAND2_X1  g1122(.A1(new_n1286), .A2(new_n1322), .ZN(new_n1323));
  NAND3_X1  g1123(.A1(new_n1296), .A2(new_n1321), .A3(new_n1323), .ZN(new_n1324));
  OR2_X1    g1124(.A1(new_n1274), .A2(new_n1324), .ZN(new_n1325));
  NOR2_X1   g1125(.A1(new_n1286), .A2(new_n1322), .ZN(new_n1326));
  NAND2_X1  g1126(.A1(new_n1274), .A2(new_n1324), .ZN(new_n1327));
  AND3_X1   g1127(.A1(new_n1325), .A2(new_n1326), .A3(new_n1327), .ZN(new_n1328));
  AOI21_X1  g1128(.A(new_n1326), .B1(new_n1325), .B2(new_n1327), .ZN(new_n1329));
  NOR2_X1   g1129(.A1(new_n1328), .A2(new_n1329), .ZN(G402));
endmodule


