

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n513, n514, n515, n516,
         n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527,
         n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538,
         n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549,
         n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560,
         n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571,
         n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582,
         n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593,
         n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604,
         n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615,
         n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626,
         n627, n628, n629, n630, n631, n632, n633, n634, n635, n636, n637,
         n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, n648,
         n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659,
         n660, n661, n662, n663, n664, n665, n666, n667, n668, n669, n670,
         n671, n672, n673, n674, n675, n676, n677, n678, n679, n680, n681,
         n682, n683, n684, n685, n686, n687, n688, n689, n690, n691, n692,
         n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, n703,
         n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, n714,
         n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, n725,
         n726, n727, n728, n729, n730, n731, n732, n733, n734, n735, n736,
         n737, n738, n739, n740, n741, n742, n743, n744, n745, n746, n747,
         n748, n749, n750, n751, n752, n753, n754, n755, n756, n757, n758,
         n759, n760, n761, n762, n763, n764, n765, n766, n767, n768, n769,
         n770, n771, n772, n773, n774, n775, n776, n777, n778, n779, n780,
         n781, n782, n783, n784, n785, n786, n787, n788, n789, n790, n791,
         n792, n793, n794, n795, n796, n797, n798, n799, n800, n801, n802,
         n803, n804, n805, n806, n807, n808, n809, n810, n811, n812, n813,
         n814, n815, n816, n817, n818, n819, n820, n821, n822, n823, n824,
         n825, n826, n827, n828, n829, n830, n831, n832, n833, n834, n835,
         n836, n837, n838, n839, n840, n841, n842, n843, n844, n845, n846,
         n847, n848, n849, n850, n851, n852, n853, n854, n855, n856, n857,
         n858, n859, n860, n861, n862, n863, n864, n865, n866, n867, n868,
         n869, n870, n871, n872, n873, n874, n875, n876, n877, n878, n879,
         n880, n881, n882, n883, n884, n885, n886, n887, n888, n889, n890,
         n891, n892, n893, n894, n895, n896, n897, n898, n899, n900, n901,
         n902, n903, n904, n905, n906, n907, n908, n909, n910, n911, n912,
         n913, n914, n915, n916, n917, n918, n919, n920, n921, n922, n923,
         n924, n925, n926, n927, n928, n929, n930, n931, n932, n933, n934,
         n935, n936, n937, n938, n939, n940, n941, n942, n943, n944, n945,
         n946, n947, n948, n949, n950, n951, n952, n953, n954, n955, n956,
         n957, n958, n959, n960, n961, n962, n963, n964, n965, n966, n967,
         n968, n969, n970, n971, n972, n973, n974, n975, n976, n977, n978,
         n979, n980, n981, n982, n983, n984, n985, n986, n987, n988, n989,
         n990, n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000,
         n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010,
         n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020,
         n1021, n1022;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NOR2_X1 U548 ( .A1(G651), .A2(n610), .ZN(n636) );
  NOR2_X2 U549 ( .A1(n666), .A2(G1384), .ZN(n667) );
  BUF_X1 U550 ( .A(n592), .Z(n593) );
  XNOR2_X1 U551 ( .A(n530), .B(KEYINPUT66), .ZN(n592) );
  NOR2_X1 U552 ( .A1(G651), .A2(G543), .ZN(n630) );
  NOR2_X2 U553 ( .A1(G2104), .A2(G2105), .ZN(n536) );
  NAND2_X1 U554 ( .A1(n761), .A2(n760), .ZN(n763) );
  NOR2_X1 U555 ( .A1(n570), .A2(n569), .ZN(n571) );
  XNOR2_X1 U556 ( .A(KEYINPUT67), .B(KEYINPUT23), .ZN(n531) );
  XOR2_X1 U557 ( .A(KEYINPUT14), .B(n559), .Z(n513) );
  NOR2_X1 U558 ( .A1(n752), .A2(n755), .ZN(n514) );
  INV_X1 U559 ( .A(KEYINPUT86), .ZN(n674) );
  INV_X1 U560 ( .A(KEYINPUT30), .ZN(n706) );
  XNOR2_X1 U561 ( .A(n706), .B(KEYINPUT87), .ZN(n707) );
  XNOR2_X1 U562 ( .A(n708), .B(n707), .ZN(n709) );
  INV_X1 U563 ( .A(KEYINPUT29), .ZN(n697) );
  XNOR2_X1 U564 ( .A(n698), .B(n697), .ZN(n703) );
  INV_X1 U565 ( .A(KEYINPUT92), .ZN(n739) );
  AND2_X1 U566 ( .A1(G2104), .A2(n535), .ZN(n530) );
  INV_X1 U567 ( .A(KEYINPUT93), .ZN(n762) );
  XOR2_X1 U568 ( .A(KEYINPUT0), .B(G543), .Z(n610) );
  XNOR2_X1 U569 ( .A(n523), .B(n522), .ZN(n631) );
  XNOR2_X1 U570 ( .A(n532), .B(n531), .ZN(n533) );
  NAND2_X1 U571 ( .A1(G89), .A2(n630), .ZN(n515) );
  XOR2_X1 U572 ( .A(KEYINPUT75), .B(n515), .Z(n516) );
  XNOR2_X1 U573 ( .A(n516), .B(KEYINPUT4), .ZN(n519) );
  INV_X1 U574 ( .A(G651), .ZN(n521) );
  OR2_X1 U575 ( .A1(n521), .A2(n610), .ZN(n517) );
  XOR2_X2 U576 ( .A(KEYINPUT68), .B(n517), .Z(n629) );
  NAND2_X1 U577 ( .A1(G76), .A2(n629), .ZN(n518) );
  NAND2_X1 U578 ( .A1(n519), .A2(n518), .ZN(n520) );
  XNOR2_X1 U579 ( .A(n520), .B(KEYINPUT5), .ZN(n528) );
  NOR2_X1 U580 ( .A1(G543), .A2(n521), .ZN(n523) );
  XNOR2_X1 U581 ( .A(KEYINPUT69), .B(KEYINPUT1), .ZN(n522) );
  NAND2_X1 U582 ( .A1(G63), .A2(n631), .ZN(n525) );
  NAND2_X1 U583 ( .A1(G51), .A2(n636), .ZN(n524) );
  NAND2_X1 U584 ( .A1(n525), .A2(n524), .ZN(n526) );
  XOR2_X1 U585 ( .A(KEYINPUT6), .B(n526), .Z(n527) );
  NAND2_X1 U586 ( .A1(n528), .A2(n527), .ZN(n529) );
  XNOR2_X1 U587 ( .A(n529), .B(KEYINPUT7), .ZN(G168) );
  XOR2_X1 U588 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  INV_X1 U589 ( .A(G2105), .ZN(n535) );
  AND2_X1 U590 ( .A1(G2105), .A2(G2104), .ZN(n867) );
  NAND2_X1 U591 ( .A1(G113), .A2(n867), .ZN(n534) );
  NAND2_X1 U592 ( .A1(n592), .A2(G101), .ZN(n532) );
  AND2_X1 U593 ( .A1(n534), .A2(n533), .ZN(n664) );
  NOR2_X2 U594 ( .A1(G2104), .A2(n535), .ZN(n869) );
  NAND2_X1 U595 ( .A1(G125), .A2(n869), .ZN(n538) );
  XOR2_X2 U596 ( .A(KEYINPUT17), .B(n536), .Z(n864) );
  NAND2_X1 U597 ( .A1(G137), .A2(n864), .ZN(n537) );
  AND2_X1 U598 ( .A1(n538), .A2(n537), .ZN(n663) );
  AND2_X1 U599 ( .A1(n664), .A2(n663), .ZN(G160) );
  AND2_X1 U600 ( .A1(G452), .A2(G94), .ZN(G173) );
  NAND2_X1 U601 ( .A1(G138), .A2(n864), .ZN(n540) );
  NAND2_X1 U602 ( .A1(G102), .A2(n592), .ZN(n539) );
  NAND2_X1 U603 ( .A1(n540), .A2(n539), .ZN(n544) );
  NAND2_X1 U604 ( .A1(G114), .A2(n867), .ZN(n542) );
  NAND2_X1 U605 ( .A1(G126), .A2(n869), .ZN(n541) );
  NAND2_X1 U606 ( .A1(n542), .A2(n541), .ZN(n543) );
  NOR2_X1 U607 ( .A1(n544), .A2(n543), .ZN(n666) );
  BUF_X1 U608 ( .A(n666), .Z(G164) );
  INV_X1 U609 ( .A(G57), .ZN(G237) );
  INV_X1 U610 ( .A(G132), .ZN(G219) );
  NAND2_X1 U611 ( .A1(G64), .A2(n631), .ZN(n546) );
  NAND2_X1 U612 ( .A1(G52), .A2(n636), .ZN(n545) );
  NAND2_X1 U613 ( .A1(n546), .A2(n545), .ZN(n552) );
  NAND2_X1 U614 ( .A1(G90), .A2(n630), .ZN(n548) );
  NAND2_X1 U615 ( .A1(G77), .A2(n629), .ZN(n547) );
  NAND2_X1 U616 ( .A1(n548), .A2(n547), .ZN(n549) );
  XOR2_X1 U617 ( .A(KEYINPUT70), .B(n549), .Z(n550) );
  XNOR2_X1 U618 ( .A(KEYINPUT9), .B(n550), .ZN(n551) );
  NOR2_X1 U619 ( .A1(n552), .A2(n551), .ZN(G171) );
  INV_X1 U620 ( .A(G171), .ZN(G301) );
  NAND2_X1 U621 ( .A1(G7), .A2(G661), .ZN(n553) );
  XOR2_X1 U622 ( .A(n553), .B(KEYINPUT10), .Z(n913) );
  NAND2_X1 U623 ( .A1(n913), .A2(G567), .ZN(n554) );
  XOR2_X1 U624 ( .A(KEYINPUT11), .B(n554), .Z(G234) );
  NAND2_X1 U625 ( .A1(n630), .A2(G81), .ZN(n555) );
  XNOR2_X1 U626 ( .A(n555), .B(KEYINPUT12), .ZN(n557) );
  NAND2_X1 U627 ( .A1(G68), .A2(n629), .ZN(n556) );
  NAND2_X1 U628 ( .A1(n557), .A2(n556), .ZN(n558) );
  XNOR2_X1 U629 ( .A(KEYINPUT13), .B(n558), .ZN(n563) );
  NAND2_X1 U630 ( .A1(G56), .A2(n631), .ZN(n559) );
  NAND2_X1 U631 ( .A1(G43), .A2(n636), .ZN(n560) );
  XNOR2_X1 U632 ( .A(KEYINPUT73), .B(n560), .ZN(n561) );
  NOR2_X1 U633 ( .A1(n513), .A2(n561), .ZN(n562) );
  NAND2_X1 U634 ( .A1(n563), .A2(n562), .ZN(n939) );
  INV_X1 U635 ( .A(G860), .ZN(n601) );
  OR2_X1 U636 ( .A1(n939), .A2(n601), .ZN(G153) );
  NAND2_X1 U637 ( .A1(G868), .A2(G301), .ZN(n573) );
  NAND2_X1 U638 ( .A1(G92), .A2(n630), .ZN(n565) );
  NAND2_X1 U639 ( .A1(G66), .A2(n631), .ZN(n564) );
  NAND2_X1 U640 ( .A1(n565), .A2(n564), .ZN(n570) );
  NAND2_X1 U641 ( .A1(n636), .A2(G54), .ZN(n567) );
  NAND2_X1 U642 ( .A1(G79), .A2(n629), .ZN(n566) );
  NAND2_X1 U643 ( .A1(n567), .A2(n566), .ZN(n568) );
  XNOR2_X1 U644 ( .A(KEYINPUT74), .B(n568), .ZN(n569) );
  XOR2_X2 U645 ( .A(n571), .B(KEYINPUT15), .Z(n942) );
  OR2_X1 U646 ( .A1(n942), .A2(G868), .ZN(n572) );
  NAND2_X1 U647 ( .A1(n573), .A2(n572), .ZN(G284) );
  NAND2_X1 U648 ( .A1(G65), .A2(n631), .ZN(n575) );
  NAND2_X1 U649 ( .A1(G53), .A2(n636), .ZN(n574) );
  NAND2_X1 U650 ( .A1(n575), .A2(n574), .ZN(n576) );
  XNOR2_X1 U651 ( .A(KEYINPUT71), .B(n576), .ZN(n580) );
  NAND2_X1 U652 ( .A1(n629), .A2(G78), .ZN(n578) );
  NAND2_X1 U653 ( .A1(G91), .A2(n630), .ZN(n577) );
  AND2_X1 U654 ( .A1(n578), .A2(n577), .ZN(n579) );
  NAND2_X1 U655 ( .A1(n580), .A2(n579), .ZN(G299) );
  XOR2_X1 U656 ( .A(KEYINPUT76), .B(G868), .Z(n581) );
  NOR2_X1 U657 ( .A1(G286), .A2(n581), .ZN(n583) );
  NOR2_X1 U658 ( .A1(G868), .A2(G299), .ZN(n582) );
  NOR2_X1 U659 ( .A1(n583), .A2(n582), .ZN(G297) );
  NAND2_X1 U660 ( .A1(n601), .A2(G559), .ZN(n584) );
  NAND2_X1 U661 ( .A1(n584), .A2(n942), .ZN(n585) );
  XNOR2_X1 U662 ( .A(n585), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U663 ( .A1(G868), .A2(n939), .ZN(n588) );
  NAND2_X1 U664 ( .A1(n942), .A2(G868), .ZN(n586) );
  NOR2_X1 U665 ( .A1(G559), .A2(n586), .ZN(n587) );
  NOR2_X1 U666 ( .A1(n588), .A2(n587), .ZN(G282) );
  NAND2_X1 U667 ( .A1(G123), .A2(n869), .ZN(n589) );
  XNOR2_X1 U668 ( .A(n589), .B(KEYINPUT18), .ZN(n591) );
  NAND2_X1 U669 ( .A1(n867), .A2(G111), .ZN(n590) );
  NAND2_X1 U670 ( .A1(n591), .A2(n590), .ZN(n597) );
  NAND2_X1 U671 ( .A1(G135), .A2(n864), .ZN(n595) );
  NAND2_X1 U672 ( .A1(G99), .A2(n593), .ZN(n594) );
  NAND2_X1 U673 ( .A1(n595), .A2(n594), .ZN(n596) );
  NOR2_X1 U674 ( .A1(n597), .A2(n596), .ZN(n927) );
  XOR2_X1 U675 ( .A(n927), .B(G2096), .Z(n598) );
  NOR2_X1 U676 ( .A1(G2100), .A2(n598), .ZN(n599) );
  XNOR2_X1 U677 ( .A(KEYINPUT77), .B(n599), .ZN(G156) );
  NAND2_X1 U678 ( .A1(G559), .A2(n942), .ZN(n600) );
  XOR2_X1 U679 ( .A(n939), .B(n600), .Z(n645) );
  NAND2_X1 U680 ( .A1(n601), .A2(n645), .ZN(n608) );
  NAND2_X1 U681 ( .A1(G67), .A2(n631), .ZN(n603) );
  NAND2_X1 U682 ( .A1(G55), .A2(n636), .ZN(n602) );
  NAND2_X1 U683 ( .A1(n603), .A2(n602), .ZN(n607) );
  NAND2_X1 U684 ( .A1(G93), .A2(n630), .ZN(n605) );
  NAND2_X1 U685 ( .A1(G80), .A2(n629), .ZN(n604) );
  NAND2_X1 U686 ( .A1(n605), .A2(n604), .ZN(n606) );
  NOR2_X1 U687 ( .A1(n607), .A2(n606), .ZN(n647) );
  XOR2_X1 U688 ( .A(n608), .B(n647), .Z(G145) );
  NAND2_X1 U689 ( .A1(G49), .A2(n636), .ZN(n609) );
  XNOR2_X1 U690 ( .A(n609), .B(KEYINPUT78), .ZN(n615) );
  NAND2_X1 U691 ( .A1(G87), .A2(n610), .ZN(n612) );
  NAND2_X1 U692 ( .A1(G74), .A2(G651), .ZN(n611) );
  NAND2_X1 U693 ( .A1(n612), .A2(n611), .ZN(n613) );
  NOR2_X1 U694 ( .A1(n631), .A2(n613), .ZN(n614) );
  NAND2_X1 U695 ( .A1(n615), .A2(n614), .ZN(G288) );
  NAND2_X1 U696 ( .A1(G88), .A2(n630), .ZN(n617) );
  NAND2_X1 U697 ( .A1(G75), .A2(n629), .ZN(n616) );
  NAND2_X1 U698 ( .A1(n617), .A2(n616), .ZN(n621) );
  NAND2_X1 U699 ( .A1(G62), .A2(n631), .ZN(n619) );
  NAND2_X1 U700 ( .A1(G50), .A2(n636), .ZN(n618) );
  NAND2_X1 U701 ( .A1(n619), .A2(n618), .ZN(n620) );
  NOR2_X1 U702 ( .A1(n621), .A2(n620), .ZN(G166) );
  INV_X1 U703 ( .A(G166), .ZN(G303) );
  NAND2_X1 U704 ( .A1(G86), .A2(n630), .ZN(n623) );
  NAND2_X1 U705 ( .A1(G61), .A2(n631), .ZN(n622) );
  NAND2_X1 U706 ( .A1(n623), .A2(n622), .ZN(n626) );
  NAND2_X1 U707 ( .A1(n629), .A2(G73), .ZN(n624) );
  XOR2_X1 U708 ( .A(KEYINPUT2), .B(n624), .Z(n625) );
  NOR2_X1 U709 ( .A1(n626), .A2(n625), .ZN(n628) );
  NAND2_X1 U710 ( .A1(n636), .A2(G48), .ZN(n627) );
  NAND2_X1 U711 ( .A1(n628), .A2(n627), .ZN(G305) );
  AND2_X1 U712 ( .A1(G72), .A2(n629), .ZN(n635) );
  NAND2_X1 U713 ( .A1(G85), .A2(n630), .ZN(n633) );
  NAND2_X1 U714 ( .A1(G60), .A2(n631), .ZN(n632) );
  NAND2_X1 U715 ( .A1(n633), .A2(n632), .ZN(n634) );
  NOR2_X1 U716 ( .A1(n635), .A2(n634), .ZN(n638) );
  NAND2_X1 U717 ( .A1(n636), .A2(G47), .ZN(n637) );
  NAND2_X1 U718 ( .A1(n638), .A2(n637), .ZN(G290) );
  XNOR2_X1 U719 ( .A(KEYINPUT19), .B(G288), .ZN(n643) );
  XNOR2_X1 U720 ( .A(n647), .B(G305), .ZN(n639) );
  INV_X1 U721 ( .A(G299), .ZN(n948) );
  XOR2_X1 U722 ( .A(n639), .B(n948), .Z(n640) );
  XOR2_X1 U723 ( .A(G303), .B(n640), .Z(n641) );
  XNOR2_X1 U724 ( .A(n641), .B(G290), .ZN(n642) );
  XNOR2_X1 U725 ( .A(n643), .B(n642), .ZN(n881) );
  XOR2_X1 U726 ( .A(n881), .B(KEYINPUT79), .Z(n644) );
  XNOR2_X1 U727 ( .A(n645), .B(n644), .ZN(n646) );
  NAND2_X1 U728 ( .A1(n646), .A2(G868), .ZN(n649) );
  OR2_X1 U729 ( .A1(G868), .A2(n647), .ZN(n648) );
  NAND2_X1 U730 ( .A1(n649), .A2(n648), .ZN(G295) );
  NAND2_X1 U731 ( .A1(G2078), .A2(G2084), .ZN(n650) );
  XOR2_X1 U732 ( .A(KEYINPUT20), .B(n650), .Z(n651) );
  NAND2_X1 U733 ( .A1(G2090), .A2(n651), .ZN(n653) );
  XNOR2_X1 U734 ( .A(KEYINPUT21), .B(KEYINPUT80), .ZN(n652) );
  XNOR2_X1 U735 ( .A(n653), .B(n652), .ZN(n654) );
  NAND2_X1 U736 ( .A1(G2072), .A2(n654), .ZN(G158) );
  XNOR2_X1 U737 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  XOR2_X1 U738 ( .A(KEYINPUT72), .B(G82), .Z(G220) );
  NOR2_X1 U739 ( .A1(G220), .A2(G219), .ZN(n655) );
  XOR2_X1 U740 ( .A(KEYINPUT22), .B(n655), .Z(n656) );
  NOR2_X1 U741 ( .A1(G218), .A2(n656), .ZN(n657) );
  NAND2_X1 U742 ( .A1(G96), .A2(n657), .ZN(n820) );
  NAND2_X1 U743 ( .A1(n820), .A2(G2106), .ZN(n661) );
  NAND2_X1 U744 ( .A1(G69), .A2(G120), .ZN(n658) );
  NOR2_X1 U745 ( .A1(G237), .A2(n658), .ZN(n659) );
  NAND2_X1 U746 ( .A1(G108), .A2(n659), .ZN(n821) );
  NAND2_X1 U747 ( .A1(n821), .A2(G567), .ZN(n660) );
  NAND2_X1 U748 ( .A1(n661), .A2(n660), .ZN(n835) );
  NAND2_X1 U749 ( .A1(G661), .A2(G483), .ZN(n662) );
  NOR2_X1 U750 ( .A1(n835), .A2(n662), .ZN(n819) );
  NAND2_X1 U751 ( .A1(n819), .A2(G36), .ZN(G176) );
  INV_X1 U752 ( .A(n942), .ZN(n682) );
  AND2_X1 U753 ( .A1(G40), .A2(n663), .ZN(n665) );
  NAND2_X1 U754 ( .A1(n665), .A2(n664), .ZN(n794) );
  XOR2_X1 U755 ( .A(n667), .B(KEYINPUT64), .Z(n795) );
  NOR2_X1 U756 ( .A1(n794), .A2(n795), .ZN(n683) );
  AND2_X1 U757 ( .A1(n683), .A2(G1996), .ZN(n668) );
  XNOR2_X1 U758 ( .A(n668), .B(KEYINPUT26), .ZN(n672) );
  INV_X1 U759 ( .A(n683), .ZN(n676) );
  NAND2_X1 U760 ( .A1(n676), .A2(G1341), .ZN(n670) );
  INV_X1 U761 ( .A(n939), .ZN(n669) );
  NAND2_X1 U762 ( .A1(n670), .A2(n669), .ZN(n671) );
  NOR2_X1 U763 ( .A1(n672), .A2(n671), .ZN(n673) );
  XNOR2_X1 U764 ( .A(KEYINPUT65), .B(n673), .ZN(n681) );
  NOR2_X1 U765 ( .A1(n682), .A2(n681), .ZN(n675) );
  XNOR2_X1 U766 ( .A(n675), .B(n674), .ZN(n680) );
  BUF_X1 U767 ( .A(n683), .Z(n699) );
  NOR2_X1 U768 ( .A1(n699), .A2(G1348), .ZN(n678) );
  NOR2_X1 U769 ( .A1(G2067), .A2(n676), .ZN(n677) );
  NOR2_X1 U770 ( .A1(n678), .A2(n677), .ZN(n679) );
  NAND2_X1 U771 ( .A1(n680), .A2(n679), .ZN(n690) );
  NAND2_X1 U772 ( .A1(n682), .A2(n681), .ZN(n688) );
  NAND2_X1 U773 ( .A1(n683), .A2(G2072), .ZN(n684) );
  XNOR2_X1 U774 ( .A(n684), .B(KEYINPUT27), .ZN(n686) );
  INV_X1 U775 ( .A(G1956), .ZN(n949) );
  NOR2_X1 U776 ( .A1(n949), .A2(n699), .ZN(n685) );
  NOR2_X1 U777 ( .A1(n686), .A2(n685), .ZN(n692) );
  NOR2_X1 U778 ( .A1(n948), .A2(n692), .ZN(n687) );
  XOR2_X1 U779 ( .A(n687), .B(KEYINPUT28), .Z(n691) );
  AND2_X1 U780 ( .A1(n688), .A2(n691), .ZN(n689) );
  NAND2_X1 U781 ( .A1(n690), .A2(n689), .ZN(n696) );
  INV_X1 U782 ( .A(n691), .ZN(n694) );
  NAND2_X1 U783 ( .A1(n948), .A2(n692), .ZN(n693) );
  OR2_X1 U784 ( .A1(n694), .A2(n693), .ZN(n695) );
  NAND2_X1 U785 ( .A1(n696), .A2(n695), .ZN(n698) );
  XOR2_X1 U786 ( .A(G2078), .B(KEYINPUT25), .Z(n998) );
  NOR2_X1 U787 ( .A1(n998), .A2(n676), .ZN(n701) );
  NOR2_X1 U788 ( .A1(n699), .A2(G1961), .ZN(n700) );
  NOR2_X1 U789 ( .A1(n701), .A2(n700), .ZN(n710) );
  NOR2_X1 U790 ( .A1(G301), .A2(n710), .ZN(n702) );
  NOR2_X1 U791 ( .A1(n703), .A2(n702), .ZN(n715) );
  NAND2_X1 U792 ( .A1(G8), .A2(n676), .ZN(n755) );
  NOR2_X1 U793 ( .A1(G1966), .A2(n755), .ZN(n730) );
  NOR2_X1 U794 ( .A1(G2084), .A2(n676), .ZN(n728) );
  INV_X1 U795 ( .A(n728), .ZN(n704) );
  NAND2_X1 U796 ( .A1(G8), .A2(n704), .ZN(n705) );
  OR2_X1 U797 ( .A1(n730), .A2(n705), .ZN(n708) );
  NOR2_X1 U798 ( .A1(G168), .A2(n709), .ZN(n712) );
  AND2_X1 U799 ( .A1(G301), .A2(n710), .ZN(n711) );
  NOR2_X1 U800 ( .A1(n712), .A2(n711), .ZN(n713) );
  XNOR2_X1 U801 ( .A(n713), .B(KEYINPUT31), .ZN(n714) );
  NOR2_X1 U802 ( .A1(n715), .A2(n714), .ZN(n716) );
  XNOR2_X1 U803 ( .A(n716), .B(KEYINPUT88), .ZN(n729) );
  INV_X1 U804 ( .A(G286), .ZN(n717) );
  OR2_X1 U805 ( .A1(n729), .A2(n717), .ZN(n725) );
  NOR2_X1 U806 ( .A1(n676), .A2(G2090), .ZN(n718) );
  XOR2_X1 U807 ( .A(KEYINPUT90), .B(n718), .Z(n719) );
  NAND2_X1 U808 ( .A1(G303), .A2(n719), .ZN(n722) );
  NOR2_X1 U809 ( .A1(G1971), .A2(n755), .ZN(n720) );
  XOR2_X1 U810 ( .A(KEYINPUT89), .B(n720), .Z(n721) );
  NOR2_X1 U811 ( .A1(n722), .A2(n721), .ZN(n723) );
  XNOR2_X1 U812 ( .A(n723), .B(KEYINPUT91), .ZN(n724) );
  NAND2_X1 U813 ( .A1(n725), .A2(n724), .ZN(n726) );
  NAND2_X1 U814 ( .A1(n726), .A2(G8), .ZN(n727) );
  XNOR2_X1 U815 ( .A(n727), .B(KEYINPUT32), .ZN(n745) );
  NAND2_X1 U816 ( .A1(G8), .A2(n728), .ZN(n732) );
  NOR2_X1 U817 ( .A1(n730), .A2(n729), .ZN(n731) );
  NAND2_X1 U818 ( .A1(n732), .A2(n731), .ZN(n746) );
  AND2_X1 U819 ( .A1(n746), .A2(n755), .ZN(n733) );
  NAND2_X1 U820 ( .A1(n745), .A2(n733), .ZN(n738) );
  INV_X1 U821 ( .A(n755), .ZN(n736) );
  NOR2_X1 U822 ( .A1(G2090), .A2(G303), .ZN(n734) );
  NAND2_X1 U823 ( .A1(G8), .A2(n734), .ZN(n735) );
  OR2_X1 U824 ( .A1(n736), .A2(n735), .ZN(n737) );
  NAND2_X1 U825 ( .A1(n738), .A2(n737), .ZN(n740) );
  XNOR2_X1 U826 ( .A(n740), .B(n739), .ZN(n744) );
  NOR2_X1 U827 ( .A1(G1981), .A2(G305), .ZN(n741) );
  XOR2_X1 U828 ( .A(n741), .B(KEYINPUT24), .Z(n742) );
  OR2_X1 U829 ( .A1(n755), .A2(n742), .ZN(n743) );
  AND2_X1 U830 ( .A1(n744), .A2(n743), .ZN(n761) );
  NAND2_X1 U831 ( .A1(n746), .A2(n745), .ZN(n751) );
  NOR2_X1 U832 ( .A1(G1971), .A2(G303), .ZN(n747) );
  NOR2_X1 U833 ( .A1(G1976), .A2(G288), .ZN(n953) );
  NOR2_X1 U834 ( .A1(n747), .A2(n953), .ZN(n749) );
  INV_X1 U835 ( .A(KEYINPUT33), .ZN(n748) );
  AND2_X1 U836 ( .A1(n749), .A2(n748), .ZN(n750) );
  NAND2_X1 U837 ( .A1(n751), .A2(n750), .ZN(n754) );
  NAND2_X1 U838 ( .A1(G1976), .A2(G288), .ZN(n950) );
  INV_X1 U839 ( .A(n950), .ZN(n752) );
  OR2_X1 U840 ( .A1(KEYINPUT33), .A2(n514), .ZN(n753) );
  NAND2_X1 U841 ( .A1(n754), .A2(n753), .ZN(n758) );
  NAND2_X1 U842 ( .A1(n953), .A2(KEYINPUT33), .ZN(n756) );
  NOR2_X1 U843 ( .A1(n756), .A2(n755), .ZN(n757) );
  NOR2_X1 U844 ( .A1(n758), .A2(n757), .ZN(n759) );
  XOR2_X1 U845 ( .A(G1981), .B(G305), .Z(n956) );
  NAND2_X1 U846 ( .A1(n759), .A2(n956), .ZN(n760) );
  XNOR2_X1 U847 ( .A(n763), .B(n762), .ZN(n799) );
  NAND2_X1 U848 ( .A1(G140), .A2(n864), .ZN(n765) );
  NAND2_X1 U849 ( .A1(G104), .A2(n593), .ZN(n764) );
  NAND2_X1 U850 ( .A1(n765), .A2(n764), .ZN(n766) );
  XNOR2_X1 U851 ( .A(KEYINPUT34), .B(n766), .ZN(n771) );
  NAND2_X1 U852 ( .A1(G116), .A2(n867), .ZN(n768) );
  NAND2_X1 U853 ( .A1(G128), .A2(n869), .ZN(n767) );
  NAND2_X1 U854 ( .A1(n768), .A2(n767), .ZN(n769) );
  XOR2_X1 U855 ( .A(n769), .B(KEYINPUT35), .Z(n770) );
  NOR2_X1 U856 ( .A1(n771), .A2(n770), .ZN(n772) );
  XOR2_X1 U857 ( .A(KEYINPUT36), .B(n772), .Z(n773) );
  XOR2_X1 U858 ( .A(KEYINPUT82), .B(n773), .Z(n877) );
  XNOR2_X1 U859 ( .A(G2067), .B(KEYINPUT37), .ZN(n774) );
  XOR2_X1 U860 ( .A(n774), .B(KEYINPUT81), .Z(n800) );
  OR2_X1 U861 ( .A1(n877), .A2(n800), .ZN(n775) );
  XOR2_X1 U862 ( .A(n775), .B(KEYINPUT83), .Z(n809) );
  INV_X1 U863 ( .A(n809), .ZN(n793) );
  NAND2_X1 U864 ( .A1(G107), .A2(n867), .ZN(n777) );
  NAND2_X1 U865 ( .A1(G119), .A2(n869), .ZN(n776) );
  NAND2_X1 U866 ( .A1(n777), .A2(n776), .ZN(n781) );
  NAND2_X1 U867 ( .A1(G131), .A2(n864), .ZN(n779) );
  NAND2_X1 U868 ( .A1(G95), .A2(n593), .ZN(n778) );
  NAND2_X1 U869 ( .A1(n779), .A2(n778), .ZN(n780) );
  NOR2_X1 U870 ( .A1(n781), .A2(n780), .ZN(n782) );
  XOR2_X1 U871 ( .A(KEYINPUT84), .B(n782), .Z(n855) );
  NAND2_X1 U872 ( .A1(n855), .A2(G1991), .ZN(n792) );
  NAND2_X1 U873 ( .A1(G117), .A2(n867), .ZN(n784) );
  NAND2_X1 U874 ( .A1(G129), .A2(n869), .ZN(n783) );
  NAND2_X1 U875 ( .A1(n784), .A2(n783), .ZN(n787) );
  NAND2_X1 U876 ( .A1(G105), .A2(n593), .ZN(n785) );
  XOR2_X1 U877 ( .A(KEYINPUT38), .B(n785), .Z(n786) );
  NOR2_X1 U878 ( .A1(n787), .A2(n786), .ZN(n788) );
  XOR2_X1 U879 ( .A(KEYINPUT85), .B(n788), .Z(n790) );
  NAND2_X1 U880 ( .A1(n864), .A2(G141), .ZN(n789) );
  NAND2_X1 U881 ( .A1(n790), .A2(n789), .ZN(n854) );
  NAND2_X1 U882 ( .A1(G1996), .A2(n854), .ZN(n791) );
  NAND2_X1 U883 ( .A1(n792), .A2(n791), .ZN(n804) );
  NOR2_X1 U884 ( .A1(n793), .A2(n804), .ZN(n923) );
  XOR2_X1 U885 ( .A(G1986), .B(G290), .Z(n955) );
  NAND2_X1 U886 ( .A1(n923), .A2(n955), .ZN(n797) );
  INV_X1 U887 ( .A(n795), .ZN(n796) );
  NOR2_X1 U888 ( .A1(n794), .A2(n796), .ZN(n812) );
  NAND2_X1 U889 ( .A1(n797), .A2(n812), .ZN(n798) );
  NAND2_X1 U890 ( .A1(n799), .A2(n798), .ZN(n815) );
  NAND2_X1 U891 ( .A1(n877), .A2(n800), .ZN(n928) );
  NOR2_X1 U892 ( .A1(G1996), .A2(n854), .ZN(n920) );
  NOR2_X1 U893 ( .A1(n855), .A2(G1991), .ZN(n930) );
  NOR2_X1 U894 ( .A1(G1986), .A2(G290), .ZN(n801) );
  NOR2_X1 U895 ( .A1(n930), .A2(n801), .ZN(n802) );
  XNOR2_X1 U896 ( .A(n802), .B(KEYINPUT94), .ZN(n803) );
  NOR2_X1 U897 ( .A1(n804), .A2(n803), .ZN(n805) );
  XOR2_X1 U898 ( .A(KEYINPUT95), .B(n805), .Z(n806) );
  NOR2_X1 U899 ( .A1(n920), .A2(n806), .ZN(n807) );
  XNOR2_X1 U900 ( .A(KEYINPUT39), .B(n807), .ZN(n808) );
  XNOR2_X1 U901 ( .A(n808), .B(KEYINPUT96), .ZN(n810) );
  NAND2_X1 U902 ( .A1(n810), .A2(n809), .ZN(n811) );
  NAND2_X1 U903 ( .A1(n928), .A2(n811), .ZN(n813) );
  NAND2_X1 U904 ( .A1(n813), .A2(n812), .ZN(n814) );
  NAND2_X1 U905 ( .A1(n815), .A2(n814), .ZN(n816) );
  XNOR2_X1 U906 ( .A(n816), .B(KEYINPUT40), .ZN(G329) );
  NAND2_X1 U907 ( .A1(G2106), .A2(n913), .ZN(G217) );
  AND2_X1 U908 ( .A1(G15), .A2(G2), .ZN(n817) );
  NAND2_X1 U909 ( .A1(G661), .A2(n817), .ZN(G259) );
  NAND2_X1 U910 ( .A1(G3), .A2(G1), .ZN(n818) );
  NAND2_X1 U911 ( .A1(n819), .A2(n818), .ZN(G188) );
  INV_X1 U913 ( .A(G120), .ZN(G236) );
  INV_X1 U914 ( .A(G96), .ZN(G221) );
  INV_X1 U915 ( .A(G69), .ZN(G235) );
  NOR2_X1 U916 ( .A1(n821), .A2(n820), .ZN(G325) );
  INV_X1 U917 ( .A(G325), .ZN(G261) );
  XOR2_X1 U918 ( .A(G2443), .B(G2451), .Z(n823) );
  XNOR2_X1 U919 ( .A(G2454), .B(G2427), .ZN(n822) );
  XNOR2_X1 U920 ( .A(n823), .B(n822), .ZN(n824) );
  XOR2_X1 U921 ( .A(n824), .B(G2430), .Z(n826) );
  XNOR2_X1 U922 ( .A(G1348), .B(G1341), .ZN(n825) );
  XNOR2_X1 U923 ( .A(n826), .B(n825), .ZN(n830) );
  XOR2_X1 U924 ( .A(KEYINPUT98), .B(G2435), .Z(n828) );
  XNOR2_X1 U925 ( .A(KEYINPUT99), .B(G2438), .ZN(n827) );
  XNOR2_X1 U926 ( .A(n828), .B(n827), .ZN(n829) );
  XOR2_X1 U927 ( .A(n830), .B(n829), .Z(n832) );
  XNOR2_X1 U928 ( .A(G2446), .B(KEYINPUT97), .ZN(n831) );
  XNOR2_X1 U929 ( .A(n832), .B(n831), .ZN(n833) );
  NAND2_X1 U930 ( .A1(G14), .A2(n833), .ZN(n834) );
  XNOR2_X1 U931 ( .A(n834), .B(KEYINPUT100), .ZN(n908) );
  XNOR2_X1 U932 ( .A(n908), .B(KEYINPUT101), .ZN(G401) );
  INV_X1 U933 ( .A(n835), .ZN(G319) );
  XOR2_X1 U934 ( .A(KEYINPUT44), .B(KEYINPUT104), .Z(n837) );
  NAND2_X1 U935 ( .A1(G124), .A2(n869), .ZN(n836) );
  XNOR2_X1 U936 ( .A(n837), .B(n836), .ZN(n844) );
  NAND2_X1 U937 ( .A1(G112), .A2(n867), .ZN(n839) );
  NAND2_X1 U938 ( .A1(G100), .A2(n593), .ZN(n838) );
  NAND2_X1 U939 ( .A1(n839), .A2(n838), .ZN(n840) );
  XNOR2_X1 U940 ( .A(n840), .B(KEYINPUT105), .ZN(n842) );
  NAND2_X1 U941 ( .A1(G136), .A2(n864), .ZN(n841) );
  NAND2_X1 U942 ( .A1(n842), .A2(n841), .ZN(n843) );
  NOR2_X1 U943 ( .A1(n844), .A2(n843), .ZN(G162) );
  NAND2_X1 U944 ( .A1(G118), .A2(n867), .ZN(n846) );
  NAND2_X1 U945 ( .A1(G130), .A2(n869), .ZN(n845) );
  NAND2_X1 U946 ( .A1(n846), .A2(n845), .ZN(n851) );
  NAND2_X1 U947 ( .A1(G142), .A2(n864), .ZN(n848) );
  NAND2_X1 U948 ( .A1(G106), .A2(n593), .ZN(n847) );
  NAND2_X1 U949 ( .A1(n848), .A2(n847), .ZN(n849) );
  XOR2_X1 U950 ( .A(KEYINPUT45), .B(n849), .Z(n850) );
  NOR2_X1 U951 ( .A1(n851), .A2(n850), .ZN(n852) );
  XOR2_X1 U952 ( .A(G162), .B(n852), .Z(n853) );
  XNOR2_X1 U953 ( .A(n854), .B(n853), .ZN(n858) );
  XNOR2_X1 U954 ( .A(n855), .B(G160), .ZN(n856) );
  XNOR2_X1 U955 ( .A(n856), .B(n927), .ZN(n857) );
  XOR2_X1 U956 ( .A(n858), .B(n857), .Z(n863) );
  XOR2_X1 U957 ( .A(KEYINPUT109), .B(KEYINPUT48), .Z(n860) );
  XNOR2_X1 U958 ( .A(KEYINPUT110), .B(KEYINPUT46), .ZN(n859) );
  XNOR2_X1 U959 ( .A(n860), .B(n859), .ZN(n861) );
  XNOR2_X1 U960 ( .A(G164), .B(n861), .ZN(n862) );
  XNOR2_X1 U961 ( .A(n863), .B(n862), .ZN(n879) );
  NAND2_X1 U962 ( .A1(G139), .A2(n864), .ZN(n866) );
  NAND2_X1 U963 ( .A1(G103), .A2(n593), .ZN(n865) );
  NAND2_X1 U964 ( .A1(n866), .A2(n865), .ZN(n875) );
  NAND2_X1 U965 ( .A1(n867), .A2(G115), .ZN(n868) );
  XNOR2_X1 U966 ( .A(n868), .B(KEYINPUT106), .ZN(n871) );
  NAND2_X1 U967 ( .A1(G127), .A2(n869), .ZN(n870) );
  NAND2_X1 U968 ( .A1(n871), .A2(n870), .ZN(n872) );
  XNOR2_X1 U969 ( .A(KEYINPUT47), .B(n872), .ZN(n873) );
  XNOR2_X1 U970 ( .A(KEYINPUT107), .B(n873), .ZN(n874) );
  NOR2_X1 U971 ( .A1(n875), .A2(n874), .ZN(n876) );
  XOR2_X1 U972 ( .A(KEYINPUT108), .B(n876), .Z(n914) );
  XOR2_X1 U973 ( .A(n914), .B(n877), .Z(n878) );
  XNOR2_X1 U974 ( .A(n879), .B(n878), .ZN(n880) );
  NOR2_X1 U975 ( .A1(G37), .A2(n880), .ZN(G395) );
  XNOR2_X1 U976 ( .A(G286), .B(n881), .ZN(n884) );
  XOR2_X1 U977 ( .A(KEYINPUT111), .B(G171), .Z(n882) );
  XNOR2_X1 U978 ( .A(n882), .B(n939), .ZN(n883) );
  XNOR2_X1 U979 ( .A(n884), .B(n883), .ZN(n885) );
  XNOR2_X1 U980 ( .A(n885), .B(n942), .ZN(n886) );
  NOR2_X1 U981 ( .A1(G37), .A2(n886), .ZN(G397) );
  XOR2_X1 U982 ( .A(G2096), .B(KEYINPUT102), .Z(n888) );
  XNOR2_X1 U983 ( .A(G2072), .B(KEYINPUT43), .ZN(n887) );
  XNOR2_X1 U984 ( .A(n888), .B(n887), .ZN(n889) );
  XOR2_X1 U985 ( .A(n889), .B(KEYINPUT42), .Z(n891) );
  XNOR2_X1 U986 ( .A(G2067), .B(G2090), .ZN(n890) );
  XNOR2_X1 U987 ( .A(n891), .B(n890), .ZN(n895) );
  XOR2_X1 U988 ( .A(G2678), .B(G2100), .Z(n893) );
  XNOR2_X1 U989 ( .A(G2078), .B(G2084), .ZN(n892) );
  XNOR2_X1 U990 ( .A(n893), .B(n892), .ZN(n894) );
  XNOR2_X1 U991 ( .A(n895), .B(n894), .ZN(G227) );
  XOR2_X1 U992 ( .A(G1966), .B(G1971), .Z(n897) );
  XNOR2_X1 U993 ( .A(G1986), .B(G1976), .ZN(n896) );
  XNOR2_X1 U994 ( .A(n897), .B(n896), .ZN(n901) );
  XNOR2_X1 U995 ( .A(n949), .B(G1981), .ZN(n899) );
  XNOR2_X1 U996 ( .A(G1996), .B(G1991), .ZN(n898) );
  XNOR2_X1 U997 ( .A(n899), .B(n898), .ZN(n900) );
  XOR2_X1 U998 ( .A(n901), .B(n900), .Z(n903) );
  XNOR2_X1 U999 ( .A(KEYINPUT103), .B(G2474), .ZN(n902) );
  XNOR2_X1 U1000 ( .A(n903), .B(n902), .ZN(n905) );
  XOR2_X1 U1001 ( .A(G1961), .B(KEYINPUT41), .Z(n904) );
  XNOR2_X1 U1002 ( .A(n905), .B(n904), .ZN(G229) );
  NOR2_X1 U1003 ( .A1(G395), .A2(G397), .ZN(n906) );
  XNOR2_X1 U1004 ( .A(n906), .B(KEYINPUT112), .ZN(n907) );
  NAND2_X1 U1005 ( .A1(n908), .A2(n907), .ZN(n911) );
  NOR2_X1 U1006 ( .A1(G227), .A2(G229), .ZN(n909) );
  XNOR2_X1 U1007 ( .A(KEYINPUT49), .B(n909), .ZN(n910) );
  NOR2_X1 U1008 ( .A1(n911), .A2(n910), .ZN(n912) );
  NAND2_X1 U1009 ( .A1(G319), .A2(n912), .ZN(G225) );
  INV_X1 U1010 ( .A(G225), .ZN(G308) );
  INV_X1 U1011 ( .A(G108), .ZN(G238) );
  INV_X1 U1012 ( .A(n913), .ZN(G223) );
  INV_X1 U1013 ( .A(KEYINPUT55), .ZN(n1016) );
  XNOR2_X1 U1014 ( .A(G164), .B(G2078), .ZN(n917) );
  XNOR2_X1 U1015 ( .A(G2072), .B(n914), .ZN(n915) );
  XNOR2_X1 U1016 ( .A(n915), .B(KEYINPUT113), .ZN(n916) );
  NAND2_X1 U1017 ( .A1(n917), .A2(n916), .ZN(n918) );
  XNOR2_X1 U1018 ( .A(n918), .B(KEYINPUT50), .ZN(n925) );
  XOR2_X1 U1019 ( .A(G2090), .B(G162), .Z(n919) );
  NOR2_X1 U1020 ( .A1(n920), .A2(n919), .ZN(n921) );
  XOR2_X1 U1021 ( .A(KEYINPUT51), .B(n921), .Z(n922) );
  NAND2_X1 U1022 ( .A1(n923), .A2(n922), .ZN(n924) );
  NOR2_X1 U1023 ( .A1(n925), .A2(n924), .ZN(n933) );
  XOR2_X1 U1024 ( .A(G2084), .B(G160), .Z(n926) );
  NOR2_X1 U1025 ( .A1(n927), .A2(n926), .ZN(n929) );
  NAND2_X1 U1026 ( .A1(n929), .A2(n928), .ZN(n931) );
  NOR2_X1 U1027 ( .A1(n931), .A2(n930), .ZN(n932) );
  NAND2_X1 U1028 ( .A1(n933), .A2(n932), .ZN(n934) );
  XNOR2_X1 U1029 ( .A(KEYINPUT114), .B(n934), .ZN(n935) );
  XOR2_X1 U1030 ( .A(KEYINPUT52), .B(n935), .Z(n936) );
  NAND2_X1 U1031 ( .A1(n1016), .A2(n936), .ZN(n937) );
  NAND2_X1 U1032 ( .A1(n937), .A2(G29), .ZN(n994) );
  XNOR2_X1 U1033 ( .A(KEYINPUT56), .B(G16), .ZN(n965) );
  XOR2_X1 U1034 ( .A(G303), .B(G1971), .Z(n938) );
  XNOR2_X1 U1035 ( .A(n938), .B(KEYINPUT122), .ZN(n941) );
  XOR2_X1 U1036 ( .A(G1341), .B(n939), .Z(n940) );
  NAND2_X1 U1037 ( .A1(n941), .A2(n940), .ZN(n947) );
  XNOR2_X1 U1038 ( .A(G1348), .B(n942), .ZN(n944) );
  XOR2_X1 U1039 ( .A(G301), .B(G1961), .Z(n943) );
  NAND2_X1 U1040 ( .A1(n944), .A2(n943), .ZN(n945) );
  XOR2_X1 U1041 ( .A(KEYINPUT121), .B(n945), .Z(n946) );
  NOR2_X1 U1042 ( .A1(n947), .A2(n946), .ZN(n963) );
  XOR2_X1 U1043 ( .A(n949), .B(n948), .Z(n951) );
  NAND2_X1 U1044 ( .A1(n951), .A2(n950), .ZN(n952) );
  NOR2_X1 U1045 ( .A1(n953), .A2(n952), .ZN(n954) );
  NAND2_X1 U1046 ( .A1(n955), .A2(n954), .ZN(n961) );
  XNOR2_X1 U1047 ( .A(G1966), .B(G168), .ZN(n957) );
  NAND2_X1 U1048 ( .A1(n957), .A2(n956), .ZN(n958) );
  XNOR2_X1 U1049 ( .A(n958), .B(KEYINPUT120), .ZN(n959) );
  XOR2_X1 U1050 ( .A(KEYINPUT57), .B(n959), .Z(n960) );
  NOR2_X1 U1051 ( .A1(n961), .A2(n960), .ZN(n962) );
  NAND2_X1 U1052 ( .A1(n963), .A2(n962), .ZN(n964) );
  NAND2_X1 U1053 ( .A1(n965), .A2(n964), .ZN(n966) );
  XNOR2_X1 U1054 ( .A(n966), .B(KEYINPUT123), .ZN(n992) );
  XOR2_X1 U1055 ( .A(G1341), .B(G19), .Z(n968) );
  XOR2_X1 U1056 ( .A(G1956), .B(G20), .Z(n967) );
  NAND2_X1 U1057 ( .A1(n968), .A2(n967), .ZN(n970) );
  XNOR2_X1 U1058 ( .A(G6), .B(G1981), .ZN(n969) );
  NOR2_X1 U1059 ( .A1(n970), .A2(n969), .ZN(n971) );
  XOR2_X1 U1060 ( .A(KEYINPUT124), .B(n971), .Z(n975) );
  XNOR2_X1 U1061 ( .A(KEYINPUT59), .B(KEYINPUT125), .ZN(n972) );
  XNOR2_X1 U1062 ( .A(n972), .B(G4), .ZN(n973) );
  XNOR2_X1 U1063 ( .A(G1348), .B(n973), .ZN(n974) );
  NOR2_X1 U1064 ( .A1(n975), .A2(n974), .ZN(n976) );
  XOR2_X1 U1065 ( .A(KEYINPUT60), .B(n976), .Z(n978) );
  XNOR2_X1 U1066 ( .A(G1966), .B(G21), .ZN(n977) );
  NOR2_X1 U1067 ( .A1(n978), .A2(n977), .ZN(n979) );
  XNOR2_X1 U1068 ( .A(KEYINPUT126), .B(n979), .ZN(n988) );
  XNOR2_X1 U1069 ( .A(G1961), .B(G5), .ZN(n986) );
  XNOR2_X1 U1070 ( .A(G1976), .B(G23), .ZN(n981) );
  XNOR2_X1 U1071 ( .A(G1971), .B(G22), .ZN(n980) );
  NOR2_X1 U1072 ( .A1(n981), .A2(n980), .ZN(n983) );
  XOR2_X1 U1073 ( .A(G1986), .B(G24), .Z(n982) );
  NAND2_X1 U1074 ( .A1(n983), .A2(n982), .ZN(n984) );
  XNOR2_X1 U1075 ( .A(KEYINPUT58), .B(n984), .ZN(n985) );
  NOR2_X1 U1076 ( .A1(n986), .A2(n985), .ZN(n987) );
  NAND2_X1 U1077 ( .A1(n988), .A2(n987), .ZN(n989) );
  XNOR2_X1 U1078 ( .A(KEYINPUT61), .B(n989), .ZN(n990) );
  NOR2_X1 U1079 ( .A1(n990), .A2(G16), .ZN(n991) );
  NOR2_X1 U1080 ( .A1(n992), .A2(n991), .ZN(n993) );
  NAND2_X1 U1081 ( .A1(n994), .A2(n993), .ZN(n1021) );
  XNOR2_X1 U1082 ( .A(KEYINPUT119), .B(G29), .ZN(n1018) );
  XOR2_X1 U1083 ( .A(KEYINPUT118), .B(G34), .Z(n996) );
  XNOR2_X1 U1084 ( .A(G2084), .B(KEYINPUT54), .ZN(n995) );
  XNOR2_X1 U1085 ( .A(n996), .B(n995), .ZN(n1014) );
  XNOR2_X1 U1086 ( .A(G2090), .B(G35), .ZN(n1012) );
  XNOR2_X1 U1087 ( .A(KEYINPUT117), .B(G1996), .ZN(n997) );
  XNOR2_X1 U1088 ( .A(n997), .B(G32), .ZN(n1006) );
  XNOR2_X1 U1089 ( .A(G1991), .B(G25), .ZN(n1000) );
  XNOR2_X1 U1090 ( .A(G27), .B(n998), .ZN(n999) );
  NOR2_X1 U1091 ( .A1(n1000), .A2(n999), .ZN(n1001) );
  NAND2_X1 U1092 ( .A1(G28), .A2(n1001), .ZN(n1004) );
  XNOR2_X1 U1093 ( .A(KEYINPUT116), .B(G2072), .ZN(n1002) );
  XNOR2_X1 U1094 ( .A(G33), .B(n1002), .ZN(n1003) );
  NOR2_X1 U1095 ( .A1(n1004), .A2(n1003), .ZN(n1005) );
  NAND2_X1 U1096 ( .A1(n1006), .A2(n1005), .ZN(n1009) );
  XOR2_X1 U1097 ( .A(KEYINPUT115), .B(G2067), .Z(n1007) );
  XNOR2_X1 U1098 ( .A(G26), .B(n1007), .ZN(n1008) );
  NOR2_X1 U1099 ( .A1(n1009), .A2(n1008), .ZN(n1010) );
  XNOR2_X1 U1100 ( .A(KEYINPUT53), .B(n1010), .ZN(n1011) );
  NOR2_X1 U1101 ( .A1(n1012), .A2(n1011), .ZN(n1013) );
  NAND2_X1 U1102 ( .A1(n1014), .A2(n1013), .ZN(n1015) );
  XNOR2_X1 U1103 ( .A(n1016), .B(n1015), .ZN(n1017) );
  NAND2_X1 U1104 ( .A1(n1018), .A2(n1017), .ZN(n1019) );
  NAND2_X1 U1105 ( .A1(n1019), .A2(G11), .ZN(n1020) );
  NOR2_X1 U1106 ( .A1(n1021), .A2(n1020), .ZN(n1022) );
  XOR2_X1 U1107 ( .A(n1022), .B(KEYINPUT62), .Z(G150) );
  INV_X1 U1108 ( .A(G150), .ZN(G311) );
endmodule

