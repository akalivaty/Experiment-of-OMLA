//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 0 0 1 0 0 0 1 1 1 0 0 1 0 1 0 1 1 1 1 0 1 0 0 0 1 1 0 0 0 1 0 0 1 1 0 1 0 0 0 0 0 0 1 1 1 1 1 0 1 1 0 1 1 1 1 0 1 1 0 0 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:31:34 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n454, new_n455,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n492, new_n493, new_n494, new_n495, new_n496,
    new_n497, new_n498, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n508, new_n509, new_n510, new_n511,
    new_n512, new_n513, new_n514, new_n515, new_n516, new_n518, new_n519,
    new_n520, new_n521, new_n522, new_n523, new_n524, new_n525, new_n526,
    new_n527, new_n528, new_n529, new_n530, new_n531, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n543, new_n545, new_n546, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n563, new_n564, new_n565, new_n567, new_n569,
    new_n570, new_n571, new_n573, new_n574, new_n575, new_n576, new_n577,
    new_n578, new_n579, new_n580, new_n581, new_n582, new_n583, new_n584,
    new_n585, new_n586, new_n587, new_n588, new_n589, new_n590, new_n592,
    new_n593, new_n594, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n611, new_n612, new_n613, new_n614, new_n617, new_n618,
    new_n620, new_n621, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n851, new_n852, new_n853, new_n854, new_n855, new_n856,
    new_n857, new_n858, new_n859, new_n860, new_n861, new_n862, new_n863,
    new_n865, new_n866, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n942, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1196,
    new_n1197, new_n1198, new_n1199, new_n1200, new_n1201, new_n1202,
    new_n1203, new_n1204, new_n1205, new_n1206, new_n1207, new_n1208,
    new_n1209, new_n1210, new_n1211, new_n1212;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  XOR2_X1   g002(.A(KEYINPUT64), .B(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  XOR2_X1   g005(.A(KEYINPUT65), .B(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  XOR2_X1   g018(.A(KEYINPUT66), .B(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n450));
  XNOR2_X1  g025(.A(new_n450), .B(KEYINPUT68), .ZN(new_n451));
  XNOR2_X1  g026(.A(KEYINPUT67), .B(KEYINPUT2), .ZN(new_n452));
  XNOR2_X1  g027(.A(new_n451), .B(new_n452), .ZN(new_n453));
  NAND4_X1  g028(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n454));
  OR2_X1    g029(.A1(new_n453), .A2(new_n454), .ZN(new_n455));
  XOR2_X1   g030(.A(new_n455), .B(KEYINPUT69), .Z(G261));
  INV_X1    g031(.A(G261), .ZN(G325));
  AOI22_X1  g032(.A1(new_n453), .A2(G2106), .B1(G567), .B2(new_n454), .ZN(G319));
  INV_X1    g033(.A(G2105), .ZN(new_n459));
  NAND3_X1  g034(.A1(new_n459), .A2(G101), .A3(G2104), .ZN(new_n460));
  OR2_X1    g035(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n461));
  NAND2_X1  g036(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n462));
  AOI21_X1  g037(.A(G2105), .B1(new_n461), .B2(new_n462), .ZN(new_n463));
  INV_X1    g038(.A(new_n463), .ZN(new_n464));
  INV_X1    g039(.A(G137), .ZN(new_n465));
  OAI21_X1  g040(.A(new_n460), .B1(new_n464), .B2(new_n465), .ZN(new_n466));
  XNOR2_X1  g041(.A(KEYINPUT3), .B(G2104), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n467), .A2(G125), .ZN(new_n468));
  NAND2_X1  g043(.A1(G113), .A2(G2104), .ZN(new_n469));
  AOI21_X1  g044(.A(new_n459), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  NOR2_X1   g045(.A1(new_n466), .A2(new_n470), .ZN(G160));
  OAI21_X1  g046(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n472));
  INV_X1    g047(.A(G112), .ZN(new_n473));
  AOI21_X1  g048(.A(new_n472), .B1(new_n473), .B2(G2105), .ZN(new_n474));
  AOI21_X1  g049(.A(new_n459), .B1(new_n461), .B2(new_n462), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n475), .A2(G124), .ZN(new_n476));
  XNOR2_X1  g051(.A(new_n476), .B(KEYINPUT70), .ZN(new_n477));
  AOI211_X1 g052(.A(new_n474), .B(new_n477), .C1(G136), .C2(new_n463), .ZN(G162));
  OR2_X1    g053(.A1(new_n459), .A2(G114), .ZN(new_n479));
  OAI21_X1  g054(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n480));
  INV_X1    g055(.A(new_n480), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n479), .A2(new_n481), .ZN(new_n482));
  AND2_X1   g057(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n483));
  NOR2_X1   g058(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n484));
  OAI211_X1 g059(.A(G126), .B(G2105), .C1(new_n483), .C2(new_n484), .ZN(new_n485));
  NAND2_X1  g060(.A1(new_n482), .A2(new_n485), .ZN(new_n486));
  OAI211_X1 g061(.A(G138), .B(new_n459), .C1(new_n483), .C2(new_n484), .ZN(new_n487));
  NAND2_X1  g062(.A1(new_n487), .A2(KEYINPUT4), .ZN(new_n488));
  INV_X1    g063(.A(KEYINPUT4), .ZN(new_n489));
  NAND4_X1  g064(.A1(new_n467), .A2(new_n489), .A3(G138), .A4(new_n459), .ZN(new_n490));
  AOI21_X1  g065(.A(new_n486), .B1(new_n488), .B2(new_n490), .ZN(G164));
  INV_X1    g066(.A(KEYINPUT71), .ZN(new_n492));
  INV_X1    g067(.A(KEYINPUT6), .ZN(new_n493));
  OAI21_X1  g068(.A(new_n492), .B1(new_n493), .B2(G651), .ZN(new_n494));
  INV_X1    g069(.A(G651), .ZN(new_n495));
  NAND3_X1  g070(.A1(new_n495), .A2(KEYINPUT71), .A3(KEYINPUT6), .ZN(new_n496));
  NAND2_X1  g071(.A1(new_n494), .A2(new_n496), .ZN(new_n497));
  OR2_X1    g072(.A1(KEYINPUT5), .A2(G543), .ZN(new_n498));
  NAND2_X1  g073(.A1(KEYINPUT5), .A2(G543), .ZN(new_n499));
  NAND2_X1  g074(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  NAND2_X1  g075(.A1(new_n493), .A2(G651), .ZN(new_n501));
  NAND4_X1  g076(.A1(new_n497), .A2(G88), .A3(new_n500), .A4(new_n501), .ZN(new_n502));
  AOI22_X1  g077(.A1(new_n500), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n503));
  OAI21_X1  g078(.A(new_n502), .B1(new_n503), .B2(new_n495), .ZN(new_n504));
  NAND3_X1  g079(.A1(new_n497), .A2(G543), .A3(new_n501), .ZN(new_n505));
  INV_X1    g080(.A(new_n505), .ZN(new_n506));
  AOI21_X1  g081(.A(new_n504), .B1(G50), .B2(new_n506), .ZN(G166));
  NAND4_X1  g082(.A1(new_n497), .A2(G89), .A3(new_n500), .A4(new_n501), .ZN(new_n508));
  NAND4_X1  g083(.A1(new_n497), .A2(G51), .A3(G543), .A4(new_n501), .ZN(new_n509));
  AND2_X1   g084(.A1(G63), .A2(G651), .ZN(new_n510));
  NAND3_X1  g085(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n511));
  NAND2_X1  g086(.A1(new_n511), .A2(KEYINPUT7), .ZN(new_n512));
  INV_X1    g087(.A(KEYINPUT7), .ZN(new_n513));
  NAND4_X1  g088(.A1(new_n513), .A2(G76), .A3(G543), .A4(G651), .ZN(new_n514));
  AOI22_X1  g089(.A1(new_n500), .A2(new_n510), .B1(new_n512), .B2(new_n514), .ZN(new_n515));
  NAND3_X1  g090(.A1(new_n508), .A2(new_n509), .A3(new_n515), .ZN(new_n516));
  INV_X1    g091(.A(new_n516), .ZN(G168));
  NAND4_X1  g092(.A1(new_n497), .A2(G52), .A3(G543), .A4(new_n501), .ZN(new_n518));
  NAND4_X1  g093(.A1(new_n497), .A2(G90), .A3(new_n500), .A4(new_n501), .ZN(new_n519));
  AND2_X1   g094(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  INV_X1    g095(.A(KEYINPUT72), .ZN(new_n521));
  INV_X1    g096(.A(G64), .ZN(new_n522));
  AOI21_X1  g097(.A(new_n522), .B1(new_n498), .B2(new_n499), .ZN(new_n523));
  NAND2_X1  g098(.A1(G77), .A2(G543), .ZN(new_n524));
  INV_X1    g099(.A(new_n524), .ZN(new_n525));
  OAI21_X1  g100(.A(new_n521), .B1(new_n523), .B2(new_n525), .ZN(new_n526));
  AND2_X1   g101(.A1(KEYINPUT5), .A2(G543), .ZN(new_n527));
  NOR2_X1   g102(.A1(KEYINPUT5), .A2(G543), .ZN(new_n528));
  NOR2_X1   g103(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  OAI211_X1 g104(.A(KEYINPUT72), .B(new_n524), .C1(new_n529), .C2(new_n522), .ZN(new_n530));
  NAND3_X1  g105(.A1(new_n526), .A2(G651), .A3(new_n530), .ZN(new_n531));
  AND2_X1   g106(.A1(new_n520), .A2(new_n531), .ZN(G171));
  INV_X1    g107(.A(G56), .ZN(new_n533));
  AOI21_X1  g108(.A(new_n533), .B1(new_n498), .B2(new_n499), .ZN(new_n534));
  AND2_X1   g109(.A1(G68), .A2(G543), .ZN(new_n535));
  OAI21_X1  g110(.A(G651), .B1(new_n534), .B2(new_n535), .ZN(new_n536));
  NAND4_X1  g111(.A1(new_n497), .A2(G81), .A3(new_n500), .A4(new_n501), .ZN(new_n537));
  INV_X1    g112(.A(G43), .ZN(new_n538));
  OAI211_X1 g113(.A(new_n536), .B(new_n537), .C1(new_n538), .C2(new_n505), .ZN(new_n539));
  INV_X1    g114(.A(new_n539), .ZN(new_n540));
  NAND2_X1  g115(.A1(new_n540), .A2(G860), .ZN(new_n541));
  XNOR2_X1  g116(.A(new_n541), .B(KEYINPUT73), .ZN(G153));
  NAND4_X1  g117(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(new_n543));
  XNOR2_X1  g118(.A(new_n543), .B(KEYINPUT74), .ZN(G176));
  NAND2_X1  g119(.A1(G1), .A2(G3), .ZN(new_n545));
  XNOR2_X1  g120(.A(new_n545), .B(KEYINPUT8), .ZN(new_n546));
  NAND4_X1  g121(.A1(G319), .A2(G483), .A3(G661), .A4(new_n546), .ZN(G188));
  NAND4_X1  g122(.A1(new_n497), .A2(G53), .A3(G543), .A4(new_n501), .ZN(new_n548));
  INV_X1    g123(.A(KEYINPUT9), .ZN(new_n549));
  NOR2_X1   g124(.A1(new_n549), .A2(KEYINPUT75), .ZN(new_n550));
  XNOR2_X1  g125(.A(new_n548), .B(new_n550), .ZN(new_n551));
  XNOR2_X1  g126(.A(KEYINPUT77), .B(G65), .ZN(new_n552));
  NAND2_X1  g127(.A1(new_n500), .A2(new_n552), .ZN(new_n553));
  NAND2_X1  g128(.A1(G78), .A2(G543), .ZN(new_n554));
  INV_X1    g129(.A(KEYINPUT76), .ZN(new_n555));
  XNOR2_X1  g130(.A(new_n554), .B(new_n555), .ZN(new_n556));
  AOI21_X1  g131(.A(new_n495), .B1(new_n553), .B2(new_n556), .ZN(new_n557));
  NAND3_X1  g132(.A1(new_n497), .A2(new_n501), .A3(new_n500), .ZN(new_n558));
  INV_X1    g133(.A(new_n558), .ZN(new_n559));
  AOI21_X1  g134(.A(new_n557), .B1(G91), .B2(new_n559), .ZN(new_n560));
  NAND2_X1  g135(.A1(new_n551), .A2(new_n560), .ZN(G299));
  NAND2_X1  g136(.A1(new_n520), .A2(new_n531), .ZN(G301));
  OR2_X1    g137(.A1(new_n516), .A2(KEYINPUT78), .ZN(new_n563));
  NAND2_X1  g138(.A1(new_n516), .A2(KEYINPUT78), .ZN(new_n564));
  NAND2_X1  g139(.A1(new_n563), .A2(new_n564), .ZN(new_n565));
  INV_X1    g140(.A(new_n565), .ZN(G286));
  INV_X1    g141(.A(G50), .ZN(new_n567));
  OAI221_X1 g142(.A(new_n502), .B1(new_n505), .B2(new_n567), .C1(new_n495), .C2(new_n503), .ZN(G303));
  NAND4_X1  g143(.A1(new_n497), .A2(G49), .A3(G543), .A4(new_n501), .ZN(new_n569));
  OAI21_X1  g144(.A(G651), .B1(new_n500), .B2(G74), .ZN(new_n570));
  INV_X1    g145(.A(G87), .ZN(new_n571));
  OAI211_X1 g146(.A(new_n569), .B(new_n570), .C1(new_n558), .C2(new_n571), .ZN(G288));
  INV_X1    g147(.A(KEYINPUT79), .ZN(new_n573));
  OAI21_X1  g148(.A(G61), .B1(new_n527), .B2(new_n528), .ZN(new_n574));
  NAND2_X1  g149(.A1(G73), .A2(G543), .ZN(new_n575));
  NAND2_X1  g150(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  AOI21_X1  g151(.A(new_n573), .B1(new_n576), .B2(G651), .ZN(new_n577));
  AOI211_X1 g152(.A(KEYINPUT79), .B(new_n495), .C1(new_n574), .C2(new_n575), .ZN(new_n578));
  NOR2_X1   g153(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  NAND4_X1  g154(.A1(new_n497), .A2(G48), .A3(G543), .A4(new_n501), .ZN(new_n580));
  NAND4_X1  g155(.A1(new_n497), .A2(G86), .A3(new_n500), .A4(new_n501), .ZN(new_n581));
  NAND2_X1  g156(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  NOR3_X1   g157(.A1(new_n579), .A2(KEYINPUT80), .A3(new_n582), .ZN(new_n583));
  INV_X1    g158(.A(KEYINPUT80), .ZN(new_n584));
  AOI22_X1  g159(.A1(new_n500), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n585));
  OAI21_X1  g160(.A(KEYINPUT79), .B1(new_n585), .B2(new_n495), .ZN(new_n586));
  NAND3_X1  g161(.A1(new_n576), .A2(new_n573), .A3(G651), .ZN(new_n587));
  NAND2_X1  g162(.A1(new_n586), .A2(new_n587), .ZN(new_n588));
  INV_X1    g163(.A(new_n582), .ZN(new_n589));
  AOI21_X1  g164(.A(new_n584), .B1(new_n588), .B2(new_n589), .ZN(new_n590));
  NOR2_X1   g165(.A1(new_n583), .A2(new_n590), .ZN(G305));
  NAND4_X1  g166(.A1(new_n497), .A2(G47), .A3(G543), .A4(new_n501), .ZN(new_n592));
  INV_X1    g167(.A(G85), .ZN(new_n593));
  AOI22_X1  g168(.A1(new_n500), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n594));
  OAI221_X1 g169(.A(new_n592), .B1(new_n558), .B2(new_n593), .C1(new_n495), .C2(new_n594), .ZN(G290));
  NAND2_X1  g170(.A1(G171), .A2(G868), .ZN(new_n596));
  NAND4_X1  g171(.A1(new_n497), .A2(G92), .A3(new_n500), .A4(new_n501), .ZN(new_n597));
  INV_X1    g172(.A(KEYINPUT10), .ZN(new_n598));
  XNOR2_X1  g173(.A(new_n597), .B(new_n598), .ZN(new_n599));
  NAND2_X1  g174(.A1(G79), .A2(G543), .ZN(new_n600));
  INV_X1    g175(.A(G66), .ZN(new_n601));
  OAI21_X1  g176(.A(new_n600), .B1(new_n529), .B2(new_n601), .ZN(new_n602));
  AOI22_X1  g177(.A1(new_n506), .A2(G54), .B1(new_n602), .B2(G651), .ZN(new_n603));
  NAND2_X1  g178(.A1(new_n599), .A2(new_n603), .ZN(new_n604));
  OR2_X1    g179(.A1(new_n604), .A2(KEYINPUT81), .ZN(new_n605));
  NAND2_X1  g180(.A1(new_n604), .A2(KEYINPUT81), .ZN(new_n606));
  NAND2_X1  g181(.A1(new_n605), .A2(new_n606), .ZN(new_n607));
  OAI21_X1  g182(.A(new_n596), .B1(new_n607), .B2(G868), .ZN(new_n608));
  XOR2_X1   g183(.A(new_n608), .B(KEYINPUT82), .Z(G284));
  XOR2_X1   g184(.A(new_n608), .B(KEYINPUT83), .Z(G321));
  INV_X1    g185(.A(G299), .ZN(new_n611));
  OAI21_X1  g186(.A(KEYINPUT84), .B1(new_n611), .B2(G868), .ZN(new_n612));
  INV_X1    g187(.A(G868), .ZN(new_n613));
  NOR2_X1   g188(.A1(new_n565), .A2(new_n613), .ZN(new_n614));
  MUX2_X1   g189(.A(new_n612), .B(KEYINPUT84), .S(new_n614), .Z(G297));
  MUX2_X1   g190(.A(new_n612), .B(KEYINPUT84), .S(new_n614), .Z(G280));
  INV_X1    g191(.A(new_n607), .ZN(new_n617));
  INV_X1    g192(.A(G559), .ZN(new_n618));
  OAI21_X1  g193(.A(new_n617), .B1(new_n618), .B2(G860), .ZN(G148));
  NAND2_X1  g194(.A1(new_n539), .A2(new_n613), .ZN(new_n620));
  NOR2_X1   g195(.A1(new_n607), .A2(G559), .ZN(new_n621));
  OAI21_X1  g196(.A(new_n620), .B1(new_n621), .B2(new_n613), .ZN(G323));
  XNOR2_X1  g197(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g198(.A1(new_n463), .A2(G135), .ZN(new_n624));
  NOR2_X1   g199(.A1(new_n459), .A2(G111), .ZN(new_n625));
  OAI21_X1  g200(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n626));
  AND3_X1   g201(.A1(new_n475), .A2(KEYINPUT85), .A3(G123), .ZN(new_n627));
  AOI21_X1  g202(.A(KEYINPUT85), .B1(new_n475), .B2(G123), .ZN(new_n628));
  OAI221_X1 g203(.A(new_n624), .B1(new_n625), .B2(new_n626), .C1(new_n627), .C2(new_n628), .ZN(new_n629));
  OR2_X1    g204(.A1(new_n629), .A2(G2096), .ZN(new_n630));
  NAND3_X1  g205(.A1(new_n459), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n631));
  XNOR2_X1  g206(.A(new_n631), .B(KEYINPUT12), .ZN(new_n632));
  XNOR2_X1  g207(.A(new_n632), .B(KEYINPUT13), .ZN(new_n633));
  INV_X1    g208(.A(G2100), .ZN(new_n634));
  NAND2_X1  g209(.A1(new_n633), .A2(new_n634), .ZN(new_n635));
  OR2_X1    g210(.A1(new_n633), .A2(new_n634), .ZN(new_n636));
  NAND2_X1  g211(.A1(new_n629), .A2(G2096), .ZN(new_n637));
  NAND4_X1  g212(.A1(new_n630), .A2(new_n635), .A3(new_n636), .A4(new_n637), .ZN(G156));
  INV_X1    g213(.A(G14), .ZN(new_n639));
  XNOR2_X1  g214(.A(G2427), .B(G2438), .ZN(new_n640));
  XNOR2_X1  g215(.A(new_n640), .B(G2430), .ZN(new_n641));
  XNOR2_X1  g216(.A(KEYINPUT15), .B(G2435), .ZN(new_n642));
  OR2_X1    g217(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  NAND2_X1  g218(.A1(new_n641), .A2(new_n642), .ZN(new_n644));
  NAND3_X1  g219(.A1(new_n643), .A2(KEYINPUT14), .A3(new_n644), .ZN(new_n645));
  XNOR2_X1  g220(.A(G2451), .B(G2454), .ZN(new_n646));
  XNOR2_X1  g221(.A(new_n646), .B(KEYINPUT16), .ZN(new_n647));
  XNOR2_X1  g222(.A(new_n645), .B(new_n647), .ZN(new_n648));
  XNOR2_X1  g223(.A(G2443), .B(G2446), .ZN(new_n649));
  XNOR2_X1  g224(.A(new_n648), .B(new_n649), .ZN(new_n650));
  XNOR2_X1  g225(.A(G1341), .B(G1348), .ZN(new_n651));
  XOR2_X1   g226(.A(new_n651), .B(KEYINPUT86), .Z(new_n652));
  INV_X1    g227(.A(new_n652), .ZN(new_n653));
  AOI21_X1  g228(.A(new_n639), .B1(new_n650), .B2(new_n653), .ZN(new_n654));
  INV_X1    g229(.A(new_n650), .ZN(new_n655));
  AOI21_X1  g230(.A(KEYINPUT87), .B1(new_n655), .B2(new_n652), .ZN(new_n656));
  INV_X1    g231(.A(KEYINPUT87), .ZN(new_n657));
  NOR3_X1   g232(.A1(new_n650), .A2(new_n657), .A3(new_n653), .ZN(new_n658));
  OAI21_X1  g233(.A(new_n654), .B1(new_n656), .B2(new_n658), .ZN(new_n659));
  INV_X1    g234(.A(new_n659), .ZN(G401));
  XNOR2_X1  g235(.A(G2067), .B(G2678), .ZN(new_n661));
  XOR2_X1   g236(.A(new_n661), .B(KEYINPUT89), .Z(new_n662));
  XNOR2_X1  g237(.A(G2084), .B(G2090), .ZN(new_n663));
  INV_X1    g238(.A(new_n663), .ZN(new_n664));
  OAI21_X1  g239(.A(KEYINPUT17), .B1(new_n662), .B2(new_n664), .ZN(new_n665));
  XOR2_X1   g240(.A(G2072), .B(G2078), .Z(new_n666));
  AOI22_X1  g241(.A1(new_n665), .A2(new_n666), .B1(new_n664), .B2(new_n662), .ZN(new_n667));
  OAI21_X1  g242(.A(new_n667), .B1(new_n666), .B2(new_n665), .ZN(new_n668));
  INV_X1    g243(.A(new_n666), .ZN(new_n669));
  NAND3_X1  g244(.A1(new_n669), .A2(new_n664), .A3(new_n661), .ZN(new_n670));
  XNOR2_X1  g245(.A(KEYINPUT88), .B(KEYINPUT18), .ZN(new_n671));
  XNOR2_X1  g246(.A(new_n670), .B(new_n671), .ZN(new_n672));
  NAND2_X1  g247(.A1(new_n668), .A2(new_n672), .ZN(new_n673));
  XNOR2_X1  g248(.A(new_n673), .B(new_n634), .ZN(new_n674));
  XNOR2_X1  g249(.A(KEYINPUT90), .B(G2096), .ZN(new_n675));
  NAND2_X1  g250(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  XNOR2_X1  g251(.A(new_n673), .B(G2100), .ZN(new_n677));
  INV_X1    g252(.A(new_n675), .ZN(new_n678));
  NAND2_X1  g253(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  NAND2_X1  g254(.A1(new_n676), .A2(new_n679), .ZN(G227));
  XNOR2_X1  g255(.A(G1981), .B(G1986), .ZN(new_n681));
  INV_X1    g256(.A(new_n681), .ZN(new_n682));
  XNOR2_X1  g257(.A(G1971), .B(G1976), .ZN(new_n683));
  INV_X1    g258(.A(KEYINPUT19), .ZN(new_n684));
  XNOR2_X1  g259(.A(new_n683), .B(new_n684), .ZN(new_n685));
  XOR2_X1   g260(.A(G1956), .B(G2474), .Z(new_n686));
  XOR2_X1   g261(.A(G1961), .B(G1966), .Z(new_n687));
  AND2_X1   g262(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  NAND2_X1  g263(.A1(new_n685), .A2(new_n688), .ZN(new_n689));
  XNOR2_X1  g264(.A(new_n689), .B(KEYINPUT20), .ZN(new_n690));
  NOR2_X1   g265(.A1(new_n686), .A2(new_n687), .ZN(new_n691));
  NOR3_X1   g266(.A1(new_n685), .A2(new_n688), .A3(new_n691), .ZN(new_n692));
  AOI21_X1  g267(.A(new_n692), .B1(new_n685), .B2(new_n691), .ZN(new_n693));
  AND2_X1   g268(.A1(new_n690), .A2(new_n693), .ZN(new_n694));
  XNOR2_X1  g269(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n695));
  INV_X1    g270(.A(new_n695), .ZN(new_n696));
  XNOR2_X1  g271(.A(new_n694), .B(new_n696), .ZN(new_n697));
  XOR2_X1   g272(.A(G1991), .B(G1996), .Z(new_n698));
  INV_X1    g273(.A(new_n698), .ZN(new_n699));
  NOR2_X1   g274(.A1(new_n697), .A2(new_n699), .ZN(new_n700));
  XNOR2_X1  g275(.A(new_n694), .B(new_n695), .ZN(new_n701));
  NOR2_X1   g276(.A1(new_n701), .A2(new_n698), .ZN(new_n702));
  OAI21_X1  g277(.A(new_n682), .B1(new_n700), .B2(new_n702), .ZN(new_n703));
  NAND2_X1  g278(.A1(new_n701), .A2(new_n698), .ZN(new_n704));
  NAND2_X1  g279(.A1(new_n697), .A2(new_n699), .ZN(new_n705));
  NAND3_X1  g280(.A1(new_n704), .A2(new_n705), .A3(new_n681), .ZN(new_n706));
  NAND2_X1  g281(.A1(new_n703), .A2(new_n706), .ZN(new_n707));
  INV_X1    g282(.A(new_n707), .ZN(G229));
  NAND2_X1  g283(.A1(new_n540), .A2(G16), .ZN(new_n709));
  OAI21_X1  g284(.A(new_n709), .B1(G16), .B2(G19), .ZN(new_n710));
  INV_X1    g285(.A(G1341), .ZN(new_n711));
  OR2_X1    g286(.A1(new_n710), .A2(new_n711), .ZN(new_n712));
  INV_X1    g287(.A(G1966), .ZN(new_n713));
  NAND2_X1  g288(.A1(new_n516), .A2(G16), .ZN(new_n714));
  INV_X1    g289(.A(G16), .ZN(new_n715));
  NAND2_X1  g290(.A1(new_n715), .A2(G21), .ZN(new_n716));
  AND2_X1   g291(.A1(new_n714), .A2(new_n716), .ZN(new_n717));
  OAI21_X1  g292(.A(new_n712), .B1(new_n713), .B2(new_n717), .ZN(new_n718));
  AOI21_X1  g293(.A(new_n718), .B1(new_n711), .B2(new_n710), .ZN(new_n719));
  NAND2_X1  g294(.A1(new_n717), .A2(new_n713), .ZN(new_n720));
  INV_X1    g295(.A(G29), .ZN(new_n721));
  NAND2_X1  g296(.A1(new_n721), .A2(G26), .ZN(new_n722));
  XOR2_X1   g297(.A(new_n722), .B(KEYINPUT28), .Z(new_n723));
  NAND2_X1  g298(.A1(new_n475), .A2(G128), .ZN(new_n724));
  INV_X1    g299(.A(G140), .ZN(new_n725));
  OAI21_X1  g300(.A(new_n724), .B1(new_n725), .B2(new_n464), .ZN(new_n726));
  NOR2_X1   g301(.A1(G104), .A2(G2105), .ZN(new_n727));
  XNOR2_X1  g302(.A(new_n727), .B(KEYINPUT92), .ZN(new_n728));
  INV_X1    g303(.A(G2104), .ZN(new_n729));
  INV_X1    g304(.A(G116), .ZN(new_n730));
  AOI21_X1  g305(.A(new_n729), .B1(new_n730), .B2(G2105), .ZN(new_n731));
  NAND2_X1  g306(.A1(new_n728), .A2(new_n731), .ZN(new_n732));
  INV_X1    g307(.A(KEYINPUT93), .ZN(new_n733));
  NAND2_X1  g308(.A1(new_n732), .A2(new_n733), .ZN(new_n734));
  NAND3_X1  g309(.A1(new_n728), .A2(KEYINPUT93), .A3(new_n731), .ZN(new_n735));
  AOI21_X1  g310(.A(new_n726), .B1(new_n734), .B2(new_n735), .ZN(new_n736));
  INV_X1    g311(.A(new_n736), .ZN(new_n737));
  AOI21_X1  g312(.A(new_n723), .B1(new_n737), .B2(G29), .ZN(new_n738));
  XNOR2_X1  g313(.A(new_n738), .B(G2067), .ZN(new_n739));
  NAND2_X1  g314(.A1(new_n715), .A2(G5), .ZN(new_n740));
  OAI21_X1  g315(.A(new_n740), .B1(G171), .B2(new_n715), .ZN(new_n741));
  INV_X1    g316(.A(G1961), .ZN(new_n742));
  XNOR2_X1  g317(.A(new_n741), .B(new_n742), .ZN(new_n743));
  AND4_X1   g318(.A1(new_n719), .A2(new_n720), .A3(new_n739), .A4(new_n743), .ZN(new_n744));
  NAND2_X1  g319(.A1(new_n715), .A2(G4), .ZN(new_n745));
  OAI21_X1  g320(.A(new_n745), .B1(new_n617), .B2(new_n715), .ZN(new_n746));
  INV_X1    g321(.A(G1348), .ZN(new_n747));
  XNOR2_X1  g322(.A(new_n746), .B(new_n747), .ZN(new_n748));
  NAND2_X1  g323(.A1(G162), .A2(G29), .ZN(new_n749));
  OR2_X1    g324(.A1(G29), .A2(G35), .ZN(new_n750));
  XNOR2_X1  g325(.A(KEYINPUT99), .B(KEYINPUT29), .ZN(new_n751));
  AND3_X1   g326(.A1(new_n749), .A2(new_n750), .A3(new_n751), .ZN(new_n752));
  AOI21_X1  g327(.A(new_n751), .B1(new_n749), .B2(new_n750), .ZN(new_n753));
  NOR3_X1   g328(.A1(new_n752), .A2(new_n753), .A3(G2090), .ZN(new_n754));
  INV_X1    g329(.A(G34), .ZN(new_n755));
  AND2_X1   g330(.A1(new_n755), .A2(KEYINPUT24), .ZN(new_n756));
  NOR2_X1   g331(.A1(new_n755), .A2(KEYINPUT24), .ZN(new_n757));
  OAI21_X1  g332(.A(new_n721), .B1(new_n756), .B2(new_n757), .ZN(new_n758));
  OAI21_X1  g333(.A(new_n758), .B1(G160), .B2(new_n721), .ZN(new_n759));
  XNOR2_X1  g334(.A(new_n759), .B(G2084), .ZN(new_n760));
  NOR2_X1   g335(.A1(G27), .A2(G29), .ZN(new_n761));
  AOI21_X1  g336(.A(new_n761), .B1(G164), .B2(G29), .ZN(new_n762));
  XNOR2_X1  g337(.A(new_n762), .B(G2078), .ZN(new_n763));
  NOR2_X1   g338(.A1(new_n629), .A2(new_n721), .ZN(new_n764));
  INV_X1    g339(.A(KEYINPUT31), .ZN(new_n765));
  OR2_X1    g340(.A1(new_n765), .A2(G11), .ZN(new_n766));
  NAND2_X1  g341(.A1(new_n765), .A2(G11), .ZN(new_n767));
  INV_X1    g342(.A(KEYINPUT30), .ZN(new_n768));
  AND2_X1   g343(.A1(new_n768), .A2(G28), .ZN(new_n769));
  OAI21_X1  g344(.A(new_n721), .B1(new_n768), .B2(G28), .ZN(new_n770));
  OAI211_X1 g345(.A(new_n766), .B(new_n767), .C1(new_n769), .C2(new_n770), .ZN(new_n771));
  OR4_X1    g346(.A1(new_n760), .A2(new_n763), .A3(new_n764), .A4(new_n771), .ZN(new_n772));
  NAND2_X1  g347(.A1(new_n721), .A2(G32), .ZN(new_n773));
  NAND3_X1  g348(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n774));
  XOR2_X1   g349(.A(new_n774), .B(KEYINPUT26), .Z(new_n775));
  NAND2_X1  g350(.A1(new_n463), .A2(G141), .ZN(new_n776));
  NAND2_X1  g351(.A1(new_n475), .A2(G129), .ZN(new_n777));
  NAND3_X1  g352(.A1(new_n459), .A2(G105), .A3(G2104), .ZN(new_n778));
  NAND4_X1  g353(.A1(new_n775), .A2(new_n776), .A3(new_n777), .A4(new_n778), .ZN(new_n779));
  INV_X1    g354(.A(new_n779), .ZN(new_n780));
  OAI21_X1  g355(.A(new_n773), .B1(new_n780), .B2(new_n721), .ZN(new_n781));
  XNOR2_X1  g356(.A(new_n781), .B(KEYINPUT27), .ZN(new_n782));
  INV_X1    g357(.A(G1996), .ZN(new_n783));
  XNOR2_X1  g358(.A(new_n782), .B(new_n783), .ZN(new_n784));
  NOR3_X1   g359(.A1(new_n754), .A2(new_n772), .A3(new_n784), .ZN(new_n785));
  NAND3_X1  g360(.A1(new_n744), .A2(new_n748), .A3(new_n785), .ZN(new_n786));
  INV_X1    g361(.A(new_n786), .ZN(new_n787));
  OAI21_X1  g362(.A(G2090), .B1(new_n752), .B2(new_n753), .ZN(new_n788));
  XNOR2_X1  g363(.A(KEYINPUT100), .B(KEYINPUT23), .ZN(new_n789));
  NAND2_X1  g364(.A1(new_n715), .A2(G20), .ZN(new_n790));
  XNOR2_X1  g365(.A(new_n789), .B(new_n790), .ZN(new_n791));
  AOI21_X1  g366(.A(new_n791), .B1(G299), .B2(G16), .ZN(new_n792));
  XNOR2_X1  g367(.A(new_n792), .B(G1956), .ZN(new_n793));
  NAND2_X1  g368(.A1(new_n788), .A2(new_n793), .ZN(new_n794));
  OR2_X1    g369(.A1(new_n794), .A2(KEYINPUT101), .ZN(new_n795));
  NOR2_X1   g370(.A1(G29), .A2(G33), .ZN(new_n796));
  XOR2_X1   g371(.A(new_n796), .B(KEYINPUT94), .Z(new_n797));
  NAND2_X1  g372(.A1(new_n467), .A2(G127), .ZN(new_n798));
  NAND2_X1  g373(.A1(G115), .A2(G2104), .ZN(new_n799));
  AOI21_X1  g374(.A(new_n459), .B1(new_n798), .B2(new_n799), .ZN(new_n800));
  INV_X1    g375(.A(new_n800), .ZN(new_n801));
  INV_X1    g376(.A(KEYINPUT95), .ZN(new_n802));
  INV_X1    g377(.A(KEYINPUT25), .ZN(new_n803));
  NAND2_X1  g378(.A1(G103), .A2(G2104), .ZN(new_n804));
  OAI21_X1  g379(.A(new_n803), .B1(new_n804), .B2(G2105), .ZN(new_n805));
  NAND4_X1  g380(.A1(new_n459), .A2(KEYINPUT25), .A3(G103), .A4(G2104), .ZN(new_n806));
  AOI22_X1  g381(.A1(new_n463), .A2(G139), .B1(new_n805), .B2(new_n806), .ZN(new_n807));
  NAND3_X1  g382(.A1(new_n801), .A2(new_n802), .A3(new_n807), .ZN(new_n808));
  INV_X1    g383(.A(new_n807), .ZN(new_n809));
  OAI21_X1  g384(.A(KEYINPUT95), .B1(new_n809), .B2(new_n800), .ZN(new_n810));
  AND3_X1   g385(.A1(new_n808), .A2(new_n810), .A3(KEYINPUT96), .ZN(new_n811));
  AOI21_X1  g386(.A(KEYINPUT96), .B1(new_n808), .B2(new_n810), .ZN(new_n812));
  NOR2_X1   g387(.A1(new_n811), .A2(new_n812), .ZN(new_n813));
  AOI21_X1  g388(.A(new_n797), .B1(new_n813), .B2(G29), .ZN(new_n814));
  NAND2_X1  g389(.A1(new_n814), .A2(G2072), .ZN(new_n815));
  XNOR2_X1  g390(.A(new_n815), .B(KEYINPUT98), .ZN(new_n816));
  AND2_X1   g391(.A1(new_n795), .A2(new_n816), .ZN(new_n817));
  INV_X1    g392(.A(KEYINPUT102), .ZN(new_n818));
  NAND2_X1  g393(.A1(new_n794), .A2(KEYINPUT101), .ZN(new_n819));
  NOR2_X1   g394(.A1(new_n814), .A2(G2072), .ZN(new_n820));
  XNOR2_X1  g395(.A(new_n820), .B(KEYINPUT97), .ZN(new_n821));
  AND2_X1   g396(.A1(new_n819), .A2(new_n821), .ZN(new_n822));
  NAND4_X1  g397(.A1(new_n787), .A2(new_n817), .A3(new_n818), .A4(new_n822), .ZN(new_n823));
  NAND4_X1  g398(.A1(new_n795), .A2(new_n816), .A3(new_n819), .A4(new_n821), .ZN(new_n824));
  OAI21_X1  g399(.A(KEYINPUT102), .B1(new_n824), .B2(new_n786), .ZN(new_n825));
  NAND2_X1  g400(.A1(G305), .A2(G16), .ZN(new_n826));
  XNOR2_X1  g401(.A(KEYINPUT32), .B(G1981), .ZN(new_n827));
  INV_X1    g402(.A(new_n827), .ZN(new_n828));
  NAND2_X1  g403(.A1(new_n715), .A2(G6), .ZN(new_n829));
  NAND3_X1  g404(.A1(new_n826), .A2(new_n828), .A3(new_n829), .ZN(new_n830));
  NAND2_X1  g405(.A1(new_n715), .A2(G22), .ZN(new_n831));
  OAI21_X1  g406(.A(new_n831), .B1(G166), .B2(new_n715), .ZN(new_n832));
  INV_X1    g407(.A(G1971), .ZN(new_n833));
  XNOR2_X1  g408(.A(new_n832), .B(new_n833), .ZN(new_n834));
  MUX2_X1   g409(.A(G23), .B(G288), .S(G16), .Z(new_n835));
  XNOR2_X1  g410(.A(KEYINPUT33), .B(G1976), .ZN(new_n836));
  XNOR2_X1  g411(.A(new_n835), .B(new_n836), .ZN(new_n837));
  NAND3_X1  g412(.A1(new_n830), .A2(new_n834), .A3(new_n837), .ZN(new_n838));
  AOI21_X1  g413(.A(new_n828), .B1(new_n826), .B2(new_n829), .ZN(new_n839));
  NOR2_X1   g414(.A1(new_n838), .A2(new_n839), .ZN(new_n840));
  INV_X1    g415(.A(KEYINPUT34), .ZN(new_n841));
  NAND2_X1  g416(.A1(new_n840), .A2(new_n841), .ZN(new_n842));
  NAND2_X1  g417(.A1(new_n463), .A2(G131), .ZN(new_n843));
  NAND2_X1  g418(.A1(new_n475), .A2(G119), .ZN(new_n844));
  NOR2_X1   g419(.A1(new_n459), .A2(G107), .ZN(new_n845));
  OAI21_X1  g420(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n846));
  OAI211_X1 g421(.A(new_n843), .B(new_n844), .C1(new_n845), .C2(new_n846), .ZN(new_n847));
  MUX2_X1   g422(.A(G25), .B(new_n847), .S(G29), .Z(new_n848));
  XOR2_X1   g423(.A(KEYINPUT35), .B(G1991), .Z(new_n849));
  XNOR2_X1  g424(.A(new_n848), .B(new_n849), .ZN(new_n850));
  INV_X1    g425(.A(G1986), .ZN(new_n851));
  AND2_X1   g426(.A1(new_n715), .A2(G24), .ZN(new_n852));
  AOI21_X1  g427(.A(new_n852), .B1(G290), .B2(G16), .ZN(new_n853));
  OAI21_X1  g428(.A(new_n850), .B1(new_n851), .B2(new_n853), .ZN(new_n854));
  AOI21_X1  g429(.A(new_n854), .B1(new_n851), .B2(new_n853), .ZN(new_n855));
  NAND2_X1  g430(.A1(new_n842), .A2(new_n855), .ZN(new_n856));
  INV_X1    g431(.A(KEYINPUT91), .ZN(new_n857));
  NOR2_X1   g432(.A1(new_n857), .A2(KEYINPUT36), .ZN(new_n858));
  NOR2_X1   g433(.A1(new_n840), .A2(new_n841), .ZN(new_n859));
  OR3_X1    g434(.A1(new_n856), .A2(new_n858), .A3(new_n859), .ZN(new_n860));
  OAI21_X1  g435(.A(new_n858), .B1(new_n856), .B2(new_n859), .ZN(new_n861));
  NAND2_X1  g436(.A1(new_n860), .A2(new_n861), .ZN(new_n862));
  NAND2_X1  g437(.A1(new_n857), .A2(KEYINPUT36), .ZN(new_n863));
  AOI22_X1  g438(.A1(new_n823), .A2(new_n825), .B1(new_n862), .B2(new_n863), .ZN(G311));
  NAND2_X1  g439(.A1(new_n823), .A2(new_n825), .ZN(new_n865));
  NAND2_X1  g440(.A1(new_n862), .A2(new_n863), .ZN(new_n866));
  NAND2_X1  g441(.A1(new_n865), .A2(new_n866), .ZN(G150));
  INV_X1    g442(.A(G860), .ZN(new_n868));
  INV_X1    g443(.A(KEYINPUT39), .ZN(new_n869));
  NOR2_X1   g444(.A1(new_n607), .A2(new_n618), .ZN(new_n870));
  XNOR2_X1  g445(.A(new_n870), .B(KEYINPUT38), .ZN(new_n871));
  INV_X1    g446(.A(G67), .ZN(new_n872));
  AOI21_X1  g447(.A(new_n872), .B1(new_n498), .B2(new_n499), .ZN(new_n873));
  AND2_X1   g448(.A1(G80), .A2(G543), .ZN(new_n874));
  OAI21_X1  g449(.A(G651), .B1(new_n873), .B2(new_n874), .ZN(new_n875));
  NAND4_X1  g450(.A1(new_n497), .A2(G55), .A3(G543), .A4(new_n501), .ZN(new_n876));
  INV_X1    g451(.A(G93), .ZN(new_n877));
  OAI211_X1 g452(.A(new_n875), .B(new_n876), .C1(new_n877), .C2(new_n558), .ZN(new_n878));
  AND2_X1   g453(.A1(new_n539), .A2(new_n878), .ZN(new_n879));
  NOR2_X1   g454(.A1(new_n539), .A2(new_n878), .ZN(new_n880));
  NOR2_X1   g455(.A1(new_n879), .A2(new_n880), .ZN(new_n881));
  XNOR2_X1  g456(.A(new_n871), .B(new_n881), .ZN(new_n882));
  AND3_X1   g457(.A1(new_n882), .A2(KEYINPUT103), .A3(new_n869), .ZN(new_n883));
  AOI21_X1  g458(.A(KEYINPUT103), .B1(new_n882), .B2(new_n869), .ZN(new_n884));
  OAI221_X1 g459(.A(new_n868), .B1(new_n869), .B2(new_n882), .C1(new_n883), .C2(new_n884), .ZN(new_n885));
  NAND2_X1  g460(.A1(new_n878), .A2(G860), .ZN(new_n886));
  XOR2_X1   g461(.A(new_n886), .B(KEYINPUT37), .Z(new_n887));
  NAND2_X1  g462(.A1(new_n885), .A2(new_n887), .ZN(G145));
  NAND2_X1  g463(.A1(new_n475), .A2(G130), .ZN(new_n889));
  NOR2_X1   g464(.A1(new_n459), .A2(G118), .ZN(new_n890));
  OAI21_X1  g465(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n891));
  OAI21_X1  g466(.A(new_n889), .B1(new_n890), .B2(new_n891), .ZN(new_n892));
  AOI21_X1  g467(.A(new_n892), .B1(G142), .B2(new_n463), .ZN(new_n893));
  XNOR2_X1  g468(.A(new_n893), .B(new_n632), .ZN(new_n894));
  XNOR2_X1  g469(.A(new_n894), .B(new_n847), .ZN(new_n895));
  NAND2_X1  g470(.A1(new_n808), .A2(new_n810), .ZN(new_n896));
  NAND2_X1  g471(.A1(new_n488), .A2(new_n490), .ZN(new_n897));
  INV_X1    g472(.A(KEYINPUT104), .ZN(new_n898));
  AOI22_X1  g473(.A1(new_n475), .A2(G126), .B1(new_n479), .B2(new_n481), .ZN(new_n899));
  AND3_X1   g474(.A1(new_n897), .A2(new_n898), .A3(new_n899), .ZN(new_n900));
  AOI21_X1  g475(.A(new_n898), .B1(new_n897), .B2(new_n899), .ZN(new_n901));
  OAI21_X1  g476(.A(new_n780), .B1(new_n900), .B2(new_n901), .ZN(new_n902));
  AOI21_X1  g477(.A(new_n489), .B1(new_n463), .B2(G138), .ZN(new_n903));
  NOR2_X1   g478(.A1(new_n487), .A2(KEYINPUT4), .ZN(new_n904));
  OAI21_X1  g479(.A(new_n899), .B1(new_n903), .B2(new_n904), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n905), .A2(KEYINPUT104), .ZN(new_n906));
  NAND3_X1  g481(.A1(new_n897), .A2(new_n898), .A3(new_n899), .ZN(new_n907));
  NAND3_X1  g482(.A1(new_n906), .A2(new_n779), .A3(new_n907), .ZN(new_n908));
  AND3_X1   g483(.A1(new_n902), .A2(new_n908), .A3(new_n736), .ZN(new_n909));
  AOI21_X1  g484(.A(new_n736), .B1(new_n902), .B2(new_n908), .ZN(new_n910));
  OAI21_X1  g485(.A(new_n896), .B1(new_n909), .B2(new_n910), .ZN(new_n911));
  NOR3_X1   g486(.A1(new_n900), .A2(new_n780), .A3(new_n901), .ZN(new_n912));
  AOI21_X1  g487(.A(new_n779), .B1(new_n906), .B2(new_n907), .ZN(new_n913));
  OAI21_X1  g488(.A(new_n737), .B1(new_n912), .B2(new_n913), .ZN(new_n914));
  NAND3_X1  g489(.A1(new_n902), .A2(new_n908), .A3(new_n736), .ZN(new_n915));
  NAND3_X1  g490(.A1(new_n914), .A2(new_n813), .A3(new_n915), .ZN(new_n916));
  NAND3_X1  g491(.A1(new_n895), .A2(new_n911), .A3(new_n916), .ZN(new_n917));
  XNOR2_X1  g492(.A(new_n629), .B(G160), .ZN(new_n918));
  XNOR2_X1  g493(.A(new_n918), .B(G162), .ZN(new_n919));
  INV_X1    g494(.A(new_n919), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n917), .A2(new_n920), .ZN(new_n921));
  INV_X1    g496(.A(new_n921), .ZN(new_n922));
  NAND2_X1  g497(.A1(new_n911), .A2(new_n916), .ZN(new_n923));
  NAND2_X1  g498(.A1(new_n923), .A2(KEYINPUT105), .ZN(new_n924));
  INV_X1    g499(.A(KEYINPUT105), .ZN(new_n925));
  NAND3_X1  g500(.A1(new_n911), .A2(new_n916), .A3(new_n925), .ZN(new_n926));
  INV_X1    g501(.A(new_n895), .ZN(new_n927));
  AND4_X1   g502(.A1(KEYINPUT106), .A2(new_n924), .A3(new_n926), .A4(new_n927), .ZN(new_n928));
  AOI21_X1  g503(.A(new_n895), .B1(new_n923), .B2(KEYINPUT105), .ZN(new_n929));
  AOI21_X1  g504(.A(KEYINPUT106), .B1(new_n929), .B2(new_n926), .ZN(new_n930));
  OAI21_X1  g505(.A(new_n922), .B1(new_n928), .B2(new_n930), .ZN(new_n931));
  INV_X1    g506(.A(KEYINPUT107), .ZN(new_n932));
  NAND2_X1  g507(.A1(new_n931), .A2(new_n932), .ZN(new_n933));
  OAI211_X1 g508(.A(new_n922), .B(KEYINPUT107), .C1(new_n928), .C2(new_n930), .ZN(new_n934));
  NAND2_X1  g509(.A1(new_n933), .A2(new_n934), .ZN(new_n935));
  NAND2_X1  g510(.A1(new_n927), .A2(new_n923), .ZN(new_n936));
  NAND2_X1  g511(.A1(new_n936), .A2(new_n917), .ZN(new_n937));
  AOI21_X1  g512(.A(G37), .B1(new_n937), .B2(new_n919), .ZN(new_n938));
  AOI21_X1  g513(.A(KEYINPUT40), .B1(new_n935), .B2(new_n938), .ZN(new_n939));
  INV_X1    g514(.A(KEYINPUT40), .ZN(new_n940));
  INV_X1    g515(.A(new_n938), .ZN(new_n941));
  AOI211_X1 g516(.A(new_n940), .B(new_n941), .C1(new_n933), .C2(new_n934), .ZN(new_n942));
  NOR2_X1   g517(.A1(new_n939), .A2(new_n942), .ZN(G395));
  NAND2_X1  g518(.A1(new_n878), .A2(new_n613), .ZN(new_n944));
  XNOR2_X1  g519(.A(new_n621), .B(new_n881), .ZN(new_n945));
  NAND2_X1  g520(.A1(G299), .A2(new_n604), .ZN(new_n946));
  NAND4_X1  g521(.A1(new_n551), .A2(new_n599), .A3(new_n560), .A4(new_n603), .ZN(new_n947));
  NAND2_X1  g522(.A1(new_n946), .A2(new_n947), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n945), .A2(new_n948), .ZN(new_n949));
  AND3_X1   g524(.A1(new_n946), .A2(KEYINPUT41), .A3(new_n947), .ZN(new_n950));
  AOI21_X1  g525(.A(KEYINPUT41), .B1(new_n946), .B2(new_n947), .ZN(new_n951));
  NOR2_X1   g526(.A1(new_n950), .A2(new_n951), .ZN(new_n952));
  OAI21_X1  g527(.A(new_n949), .B1(new_n945), .B2(new_n952), .ZN(new_n953));
  OAI21_X1  g528(.A(G166), .B1(new_n583), .B2(new_n590), .ZN(new_n954));
  OAI21_X1  g529(.A(KEYINPUT80), .B1(new_n579), .B2(new_n582), .ZN(new_n955));
  NAND3_X1  g530(.A1(new_n588), .A2(new_n584), .A3(new_n589), .ZN(new_n956));
  NAND3_X1  g531(.A1(new_n955), .A2(new_n956), .A3(G303), .ZN(new_n957));
  NAND2_X1  g532(.A1(new_n954), .A2(new_n957), .ZN(new_n958));
  OR2_X1    g533(.A1(G290), .A2(G288), .ZN(new_n959));
  NAND2_X1  g534(.A1(G290), .A2(G288), .ZN(new_n960));
  NAND3_X1  g535(.A1(new_n959), .A2(KEYINPUT108), .A3(new_n960), .ZN(new_n961));
  INV_X1    g536(.A(new_n961), .ZN(new_n962));
  NAND2_X1  g537(.A1(new_n958), .A2(new_n962), .ZN(new_n963));
  INV_X1    g538(.A(KEYINPUT108), .ZN(new_n964));
  INV_X1    g539(.A(new_n960), .ZN(new_n965));
  NOR2_X1   g540(.A1(G290), .A2(G288), .ZN(new_n966));
  OAI21_X1  g541(.A(new_n964), .B1(new_n965), .B2(new_n966), .ZN(new_n967));
  NAND4_X1  g542(.A1(new_n967), .A2(new_n961), .A3(new_n954), .A4(new_n957), .ZN(new_n968));
  AND2_X1   g543(.A1(new_n963), .A2(new_n968), .ZN(new_n969));
  XOR2_X1   g544(.A(new_n969), .B(KEYINPUT42), .Z(new_n970));
  XNOR2_X1  g545(.A(new_n953), .B(new_n970), .ZN(new_n971));
  OAI21_X1  g546(.A(new_n944), .B1(new_n971), .B2(new_n613), .ZN(G295));
  OAI21_X1  g547(.A(new_n944), .B1(new_n971), .B2(new_n613), .ZN(G331));
  INV_X1    g548(.A(KEYINPUT44), .ZN(new_n974));
  INV_X1    g549(.A(new_n969), .ZN(new_n975));
  INV_X1    g550(.A(KEYINPUT109), .ZN(new_n976));
  OAI21_X1  g551(.A(new_n976), .B1(G171), .B2(new_n516), .ZN(new_n977));
  NAND3_X1  g552(.A1(G301), .A2(KEYINPUT109), .A3(G168), .ZN(new_n978));
  AND2_X1   g553(.A1(new_n977), .A2(new_n978), .ZN(new_n979));
  OAI21_X1  g554(.A(KEYINPUT110), .B1(new_n879), .B2(new_n880), .ZN(new_n980));
  INV_X1    g555(.A(new_n880), .ZN(new_n981));
  INV_X1    g556(.A(KEYINPUT110), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n539), .A2(new_n878), .ZN(new_n983));
  NAND3_X1  g558(.A1(new_n981), .A2(new_n982), .A3(new_n983), .ZN(new_n984));
  NAND3_X1  g559(.A1(G171), .A2(new_n563), .A3(new_n564), .ZN(new_n985));
  NAND4_X1  g560(.A1(new_n979), .A2(new_n980), .A3(new_n984), .A4(new_n985), .ZN(new_n986));
  NAND2_X1  g561(.A1(new_n984), .A2(new_n980), .ZN(new_n987));
  NAND3_X1  g562(.A1(new_n977), .A2(new_n985), .A3(new_n978), .ZN(new_n988));
  NAND2_X1  g563(.A1(new_n987), .A2(new_n988), .ZN(new_n989));
  AND3_X1   g564(.A1(new_n986), .A2(new_n952), .A3(new_n989), .ZN(new_n990));
  AOI21_X1  g565(.A(new_n948), .B1(new_n986), .B2(new_n989), .ZN(new_n991));
  OAI21_X1  g566(.A(new_n975), .B1(new_n990), .B2(new_n991), .ZN(new_n992));
  INV_X1    g567(.A(KEYINPUT43), .ZN(new_n993));
  INV_X1    g568(.A(G37), .ZN(new_n994));
  INV_X1    g569(.A(new_n948), .ZN(new_n995));
  AND2_X1   g570(.A1(new_n987), .A2(new_n988), .ZN(new_n996));
  NOR2_X1   g571(.A1(new_n987), .A2(new_n988), .ZN(new_n997));
  OAI21_X1  g572(.A(new_n995), .B1(new_n996), .B2(new_n997), .ZN(new_n998));
  NAND3_X1  g573(.A1(new_n986), .A2(new_n952), .A3(new_n989), .ZN(new_n999));
  NAND3_X1  g574(.A1(new_n998), .A2(new_n999), .A3(new_n969), .ZN(new_n1000));
  NAND4_X1  g575(.A1(new_n992), .A2(new_n993), .A3(new_n994), .A4(new_n1000), .ZN(new_n1001));
  INV_X1    g576(.A(KEYINPUT112), .ZN(new_n1002));
  XNOR2_X1  g577(.A(new_n1001), .B(new_n1002), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n1000), .A2(new_n994), .ZN(new_n1004));
  AOI21_X1  g579(.A(new_n969), .B1(new_n998), .B2(new_n999), .ZN(new_n1005));
  OAI21_X1  g580(.A(KEYINPUT43), .B1(new_n1004), .B2(new_n1005), .ZN(new_n1006));
  INV_X1    g581(.A(KEYINPUT111), .ZN(new_n1007));
  NAND2_X1  g582(.A1(new_n1006), .A2(new_n1007), .ZN(new_n1008));
  OAI211_X1 g583(.A(KEYINPUT111), .B(KEYINPUT43), .C1(new_n1004), .C2(new_n1005), .ZN(new_n1009));
  NAND2_X1  g584(.A1(new_n1008), .A2(new_n1009), .ZN(new_n1010));
  OAI21_X1  g585(.A(new_n974), .B1(new_n1003), .B2(new_n1010), .ZN(new_n1011));
  NAND3_X1  g586(.A1(new_n1006), .A2(KEYINPUT44), .A3(new_n1001), .ZN(new_n1012));
  NAND2_X1  g587(.A1(new_n1011), .A2(new_n1012), .ZN(G397));
  INV_X1    g588(.A(G1384), .ZN(new_n1014));
  NAND3_X1  g589(.A1(new_n906), .A2(new_n1014), .A3(new_n907), .ZN(new_n1015));
  INV_X1    g590(.A(KEYINPUT45), .ZN(new_n1016));
  NAND2_X1  g591(.A1(new_n1015), .A2(new_n1016), .ZN(new_n1017));
  INV_X1    g592(.A(G40), .ZN(new_n1018));
  NOR3_X1   g593(.A1(new_n466), .A2(new_n470), .A3(new_n1018), .ZN(new_n1019));
  INV_X1    g594(.A(new_n1019), .ZN(new_n1020));
  NOR2_X1   g595(.A1(new_n1017), .A2(new_n1020), .ZN(new_n1021));
  XNOR2_X1  g596(.A(new_n736), .B(G2067), .ZN(new_n1022));
  XNOR2_X1  g597(.A(new_n779), .B(new_n783), .ZN(new_n1023));
  AND2_X1   g598(.A1(new_n1022), .A2(new_n1023), .ZN(new_n1024));
  XNOR2_X1  g599(.A(new_n847), .B(new_n849), .ZN(new_n1025));
  NAND2_X1  g600(.A1(new_n1024), .A2(new_n1025), .ZN(new_n1026));
  XNOR2_X1  g601(.A(G290), .B(G1986), .ZN(new_n1027));
  OAI21_X1  g602(.A(new_n1021), .B1(new_n1026), .B2(new_n1027), .ZN(new_n1028));
  NAND4_X1  g603(.A1(new_n906), .A2(KEYINPUT45), .A3(new_n1014), .A4(new_n907), .ZN(new_n1029));
  NAND2_X1  g604(.A1(new_n905), .A2(new_n1014), .ZN(new_n1030));
  INV_X1    g605(.A(KEYINPUT113), .ZN(new_n1031));
  NAND3_X1  g606(.A1(new_n1030), .A2(new_n1031), .A3(new_n1016), .ZN(new_n1032));
  AOI21_X1  g607(.A(G1384), .B1(new_n897), .B2(new_n899), .ZN(new_n1033));
  OAI21_X1  g608(.A(KEYINPUT113), .B1(new_n1033), .B2(KEYINPUT45), .ZN(new_n1034));
  NAND4_X1  g609(.A1(new_n1029), .A2(new_n1032), .A3(new_n1019), .A4(new_n1034), .ZN(new_n1035));
  XOR2_X1   g610(.A(KEYINPUT56), .B(G2072), .Z(new_n1036));
  INV_X1    g611(.A(KEYINPUT50), .ZN(new_n1037));
  NAND2_X1  g612(.A1(new_n1033), .A2(new_n1037), .ZN(new_n1038));
  OAI21_X1  g613(.A(KEYINPUT50), .B1(G164), .B2(G1384), .ZN(new_n1039));
  NAND3_X1  g614(.A1(new_n1038), .A2(new_n1039), .A3(new_n1019), .ZN(new_n1040));
  INV_X1    g615(.A(new_n1040), .ZN(new_n1041));
  XNOR2_X1  g616(.A(KEYINPUT118), .B(G1956), .ZN(new_n1042));
  OAI22_X1  g617(.A1(new_n1035), .A2(new_n1036), .B1(new_n1041), .B2(new_n1042), .ZN(new_n1043));
  INV_X1    g618(.A(KEYINPUT119), .ZN(new_n1044));
  AOI21_X1  g619(.A(KEYINPUT57), .B1(new_n551), .B2(new_n1044), .ZN(new_n1045));
  XNOR2_X1  g620(.A(new_n611), .B(new_n1045), .ZN(new_n1046));
  OR2_X1    g621(.A1(new_n1043), .A2(new_n1046), .ZN(new_n1047));
  INV_X1    g622(.A(KEYINPUT120), .ZN(new_n1048));
  NAND2_X1  g623(.A1(new_n1040), .A2(new_n1048), .ZN(new_n1049));
  NAND4_X1  g624(.A1(new_n1038), .A2(new_n1039), .A3(KEYINPUT120), .A4(new_n1019), .ZN(new_n1050));
  NAND3_X1  g625(.A1(new_n1049), .A2(new_n747), .A3(new_n1050), .ZN(new_n1051));
  INV_X1    g626(.A(G2067), .ZN(new_n1052));
  NAND3_X1  g627(.A1(new_n1019), .A2(new_n1052), .A3(new_n1033), .ZN(new_n1053));
  AOI21_X1  g628(.A(new_n604), .B1(new_n1051), .B2(new_n1053), .ZN(new_n1054));
  NAND2_X1  g629(.A1(new_n1047), .A2(new_n1054), .ZN(new_n1055));
  NAND2_X1  g630(.A1(new_n1043), .A2(new_n1046), .ZN(new_n1056));
  NAND2_X1  g631(.A1(new_n1055), .A2(new_n1056), .ZN(new_n1057));
  XNOR2_X1  g632(.A(KEYINPUT122), .B(KEYINPUT59), .ZN(new_n1058));
  NOR2_X1   g633(.A1(new_n1020), .A2(G1996), .ZN(new_n1059));
  NAND4_X1  g634(.A1(new_n1059), .A2(new_n1029), .A3(new_n1034), .A4(new_n1032), .ZN(new_n1060));
  XOR2_X1   g635(.A(KEYINPUT58), .B(G1341), .Z(new_n1061));
  OAI21_X1  g636(.A(new_n1061), .B1(new_n1020), .B2(new_n1030), .ZN(new_n1062));
  AND3_X1   g637(.A1(new_n1060), .A2(KEYINPUT121), .A3(new_n1062), .ZN(new_n1063));
  AOI21_X1  g638(.A(KEYINPUT121), .B1(new_n1060), .B2(new_n1062), .ZN(new_n1064));
  OAI211_X1 g639(.A(new_n540), .B(new_n1058), .C1(new_n1063), .C2(new_n1064), .ZN(new_n1065));
  OAI21_X1  g640(.A(new_n540), .B1(new_n1063), .B2(new_n1064), .ZN(new_n1066));
  INV_X1    g641(.A(new_n1058), .ZN(new_n1067));
  NAND2_X1  g642(.A1(new_n1066), .A2(new_n1067), .ZN(new_n1068));
  NAND3_X1  g643(.A1(new_n1047), .A2(new_n1056), .A3(KEYINPUT61), .ZN(new_n1069));
  AND3_X1   g644(.A1(new_n1051), .A2(new_n604), .A3(new_n1053), .ZN(new_n1070));
  OAI21_X1  g645(.A(KEYINPUT60), .B1(new_n1070), .B2(new_n1054), .ZN(new_n1071));
  AND4_X1   g646(.A1(new_n1065), .A2(new_n1068), .A3(new_n1069), .A4(new_n1071), .ZN(new_n1072));
  AOI21_X1  g647(.A(KEYINPUT61), .B1(new_n1047), .B2(new_n1056), .ZN(new_n1073));
  NAND2_X1  g648(.A1(new_n1051), .A2(new_n1053), .ZN(new_n1074));
  NOR3_X1   g649(.A1(new_n1074), .A2(KEYINPUT60), .A3(new_n604), .ZN(new_n1075));
  NOR2_X1   g650(.A1(new_n1073), .A2(new_n1075), .ZN(new_n1076));
  AOI21_X1  g651(.A(new_n1057), .B1(new_n1072), .B2(new_n1076), .ZN(new_n1077));
  INV_X1    g652(.A(G2084), .ZN(new_n1078));
  NAND2_X1  g653(.A1(new_n1033), .A2(KEYINPUT45), .ZN(new_n1079));
  OAI21_X1  g654(.A(new_n1016), .B1(G164), .B2(G1384), .ZN(new_n1080));
  NAND3_X1  g655(.A1(new_n1079), .A2(new_n1080), .A3(new_n1019), .ZN(new_n1081));
  AOI22_X1  g656(.A1(new_n1041), .A2(new_n1078), .B1(new_n1081), .B2(new_n713), .ZN(new_n1082));
  INV_X1    g657(.A(G8), .ZN(new_n1083));
  NOR2_X1   g658(.A1(G168), .A2(new_n1083), .ZN(new_n1084));
  INV_X1    g659(.A(new_n1084), .ZN(new_n1085));
  OAI21_X1  g660(.A(KEYINPUT123), .B1(new_n1082), .B2(new_n1085), .ZN(new_n1086));
  NAND2_X1  g661(.A1(new_n1081), .A2(new_n713), .ZN(new_n1087));
  OAI21_X1  g662(.A(new_n1087), .B1(G2084), .B2(new_n1040), .ZN(new_n1088));
  INV_X1    g663(.A(KEYINPUT123), .ZN(new_n1089));
  NAND3_X1  g664(.A1(new_n1088), .A2(new_n1089), .A3(new_n1084), .ZN(new_n1090));
  AOI21_X1  g665(.A(new_n1083), .B1(new_n1082), .B2(G168), .ZN(new_n1091));
  INV_X1    g666(.A(KEYINPUT51), .ZN(new_n1092));
  AOI22_X1  g667(.A1(new_n1086), .A2(new_n1090), .B1(new_n1091), .B2(new_n1092), .ZN(new_n1093));
  OAI211_X1 g668(.A(KEYINPUT51), .B(new_n1085), .C1(new_n1082), .C2(new_n1083), .ZN(new_n1094));
  INV_X1    g669(.A(KEYINPUT53), .ZN(new_n1095));
  OAI21_X1  g670(.A(new_n1095), .B1(new_n1035), .B2(G2078), .ZN(new_n1096));
  NAND3_X1  g671(.A1(new_n1049), .A2(new_n742), .A3(new_n1050), .ZN(new_n1097));
  NOR2_X1   g672(.A1(new_n1095), .A2(G2078), .ZN(new_n1098));
  NAND4_X1  g673(.A1(new_n1079), .A2(new_n1080), .A3(new_n1019), .A4(new_n1098), .ZN(new_n1099));
  NAND3_X1  g674(.A1(new_n1096), .A2(new_n1097), .A3(new_n1099), .ZN(new_n1100));
  OR2_X1    g675(.A1(new_n1100), .A2(G171), .ZN(new_n1101));
  INV_X1    g676(.A(KEYINPUT54), .ZN(new_n1102));
  NAND4_X1  g677(.A1(new_n1017), .A2(new_n1019), .A3(new_n1029), .A4(new_n1098), .ZN(new_n1103));
  NAND3_X1  g678(.A1(new_n1096), .A2(new_n1097), .A3(new_n1103), .ZN(new_n1104));
  AOI21_X1  g679(.A(new_n1102), .B1(new_n1104), .B2(G171), .ZN(new_n1105));
  AOI22_X1  g680(.A1(new_n1093), .A2(new_n1094), .B1(new_n1101), .B2(new_n1105), .ZN(new_n1106));
  INV_X1    g681(.A(KEYINPUT52), .ZN(new_n1107));
  AOI21_X1  g682(.A(new_n1083), .B1(new_n1019), .B2(new_n1033), .ZN(new_n1108));
  INV_X1    g683(.A(G1976), .ZN(new_n1109));
  OR2_X1    g684(.A1(G288), .A2(new_n1109), .ZN(new_n1110));
  AOI21_X1  g685(.A(new_n1107), .B1(new_n1108), .B2(new_n1110), .ZN(new_n1111));
  AND2_X1   g686(.A1(new_n1108), .A2(new_n1110), .ZN(new_n1112));
  AOI21_X1  g687(.A(KEYINPUT52), .B1(G288), .B2(new_n1109), .ZN(new_n1113));
  AOI21_X1  g688(.A(new_n1111), .B1(new_n1112), .B2(new_n1113), .ZN(new_n1114));
  OAI21_X1  g689(.A(G1981), .B1(new_n579), .B2(new_n582), .ZN(new_n1115));
  XOR2_X1   g690(.A(KEYINPUT115), .B(G1981), .Z(new_n1116));
  NAND3_X1  g691(.A1(new_n588), .A2(new_n589), .A3(new_n1116), .ZN(new_n1117));
  NAND3_X1  g692(.A1(new_n1115), .A2(new_n1117), .A3(KEYINPUT49), .ZN(new_n1118));
  AOI21_X1  g693(.A(KEYINPUT49), .B1(new_n1115), .B2(new_n1117), .ZN(new_n1119));
  INV_X1    g694(.A(KEYINPUT116), .ZN(new_n1120));
  OAI211_X1 g695(.A(new_n1108), .B(new_n1118), .C1(new_n1119), .C2(new_n1120), .ZN(new_n1121));
  AND2_X1   g696(.A1(new_n1119), .A2(new_n1120), .ZN(new_n1122));
  OAI21_X1  g697(.A(new_n1114), .B1(new_n1121), .B2(new_n1122), .ZN(new_n1123));
  NAND2_X1  g698(.A1(new_n1123), .A2(KEYINPUT117), .ZN(new_n1124));
  NAND3_X1  g699(.A1(G303), .A2(KEYINPUT55), .A3(G8), .ZN(new_n1125));
  INV_X1    g700(.A(KEYINPUT114), .ZN(new_n1126));
  OR2_X1    g701(.A1(new_n1125), .A2(new_n1126), .ZN(new_n1127));
  NAND2_X1  g702(.A1(new_n1125), .A2(new_n1126), .ZN(new_n1128));
  INV_X1    g703(.A(KEYINPUT55), .ZN(new_n1129));
  OAI21_X1  g704(.A(new_n1129), .B1(G166), .B2(new_n1083), .ZN(new_n1130));
  NAND3_X1  g705(.A1(new_n1127), .A2(new_n1128), .A3(new_n1130), .ZN(new_n1131));
  AND2_X1   g706(.A1(new_n1035), .A2(new_n833), .ZN(new_n1132));
  NOR2_X1   g707(.A1(new_n1040), .A2(G2090), .ZN(new_n1133));
  OAI211_X1 g708(.A(G8), .B(new_n1131), .C1(new_n1132), .C2(new_n1133), .ZN(new_n1134));
  AND3_X1   g709(.A1(new_n1127), .A2(new_n1128), .A3(new_n1130), .ZN(new_n1135));
  INV_X1    g710(.A(G2090), .ZN(new_n1136));
  AOI22_X1  g711(.A1(new_n1035), .A2(new_n833), .B1(new_n1041), .B2(new_n1136), .ZN(new_n1137));
  OAI21_X1  g712(.A(new_n1135), .B1(new_n1137), .B2(new_n1083), .ZN(new_n1138));
  INV_X1    g713(.A(KEYINPUT117), .ZN(new_n1139));
  OAI211_X1 g714(.A(new_n1114), .B(new_n1139), .C1(new_n1121), .C2(new_n1122), .ZN(new_n1140));
  NAND4_X1  g715(.A1(new_n1124), .A2(new_n1134), .A3(new_n1138), .A4(new_n1140), .ZN(new_n1141));
  INV_X1    g716(.A(KEYINPUT124), .ZN(new_n1142));
  NAND2_X1  g717(.A1(new_n1141), .A2(new_n1142), .ZN(new_n1143));
  AND2_X1   g718(.A1(new_n1134), .A2(new_n1138), .ZN(new_n1144));
  NAND4_X1  g719(.A1(new_n1144), .A2(KEYINPUT124), .A3(new_n1124), .A4(new_n1140), .ZN(new_n1145));
  NAND2_X1  g720(.A1(new_n1100), .A2(G171), .ZN(new_n1146));
  OAI21_X1  g721(.A(new_n1146), .B1(G171), .B2(new_n1104), .ZN(new_n1147));
  NAND2_X1  g722(.A1(new_n1147), .A2(new_n1102), .ZN(new_n1148));
  NAND4_X1  g723(.A1(new_n1106), .A2(new_n1143), .A3(new_n1145), .A4(new_n1148), .ZN(new_n1149));
  NOR2_X1   g724(.A1(new_n1077), .A2(new_n1149), .ZN(new_n1150));
  NAND2_X1  g725(.A1(new_n1086), .A2(new_n1090), .ZN(new_n1151));
  OAI211_X1 g726(.A(new_n1092), .B(G8), .C1(new_n1088), .C2(new_n516), .ZN(new_n1152));
  NAND3_X1  g727(.A1(new_n1151), .A2(new_n1094), .A3(new_n1152), .ZN(new_n1153));
  AOI21_X1  g728(.A(new_n1146), .B1(new_n1153), .B2(KEYINPUT62), .ZN(new_n1154));
  INV_X1    g729(.A(KEYINPUT62), .ZN(new_n1155));
  NAND3_X1  g730(.A1(new_n1093), .A2(new_n1155), .A3(new_n1094), .ZN(new_n1156));
  NAND4_X1  g731(.A1(new_n1154), .A2(new_n1143), .A3(new_n1145), .A4(new_n1156), .ZN(new_n1157));
  INV_X1    g732(.A(KEYINPUT63), .ZN(new_n1158));
  NAND3_X1  g733(.A1(new_n1088), .A2(G8), .A3(new_n565), .ZN(new_n1159));
  OAI21_X1  g734(.A(new_n1158), .B1(new_n1141), .B2(new_n1159), .ZN(new_n1160));
  NOR3_X1   g735(.A1(new_n1123), .A2(new_n1159), .A3(new_n1158), .ZN(new_n1161));
  NAND2_X1  g736(.A1(new_n1144), .A2(new_n1161), .ZN(new_n1162));
  NAND2_X1  g737(.A1(new_n1160), .A2(new_n1162), .ZN(new_n1163));
  NOR2_X1   g738(.A1(new_n1134), .A2(new_n1123), .ZN(new_n1164));
  NOR2_X1   g739(.A1(new_n1121), .A2(new_n1122), .ZN(new_n1165));
  OR2_X1    g740(.A1(G288), .A2(G1976), .ZN(new_n1166));
  OAI21_X1  g741(.A(new_n1117), .B1(new_n1165), .B2(new_n1166), .ZN(new_n1167));
  AOI21_X1  g742(.A(new_n1164), .B1(new_n1108), .B2(new_n1167), .ZN(new_n1168));
  NAND3_X1  g743(.A1(new_n1157), .A2(new_n1163), .A3(new_n1168), .ZN(new_n1169));
  OAI21_X1  g744(.A(new_n1028), .B1(new_n1150), .B2(new_n1169), .ZN(new_n1170));
  AOI21_X1  g745(.A(new_n779), .B1(KEYINPUT46), .B2(new_n783), .ZN(new_n1171));
  AND2_X1   g746(.A1(new_n1022), .A2(new_n1171), .ZN(new_n1172));
  INV_X1    g747(.A(new_n1021), .ZN(new_n1173));
  NOR2_X1   g748(.A1(new_n1172), .A2(new_n1173), .ZN(new_n1174));
  AOI21_X1  g749(.A(KEYINPUT46), .B1(new_n1021), .B2(new_n783), .ZN(new_n1175));
  INV_X1    g750(.A(new_n1175), .ZN(new_n1176));
  AOI21_X1  g751(.A(new_n1174), .B1(KEYINPUT125), .B2(new_n1176), .ZN(new_n1177));
  OAI21_X1  g752(.A(new_n1177), .B1(KEYINPUT125), .B2(new_n1176), .ZN(new_n1178));
  INV_X1    g753(.A(KEYINPUT47), .ZN(new_n1179));
  OR2_X1    g754(.A1(new_n1178), .A2(new_n1179), .ZN(new_n1180));
  INV_X1    g755(.A(new_n849), .ZN(new_n1181));
  NOR2_X1   g756(.A1(new_n847), .A2(new_n1181), .ZN(new_n1182));
  NAND2_X1  g757(.A1(new_n1024), .A2(new_n1182), .ZN(new_n1183));
  NAND2_X1  g758(.A1(new_n736), .A2(new_n1052), .ZN(new_n1184));
  AOI21_X1  g759(.A(new_n1173), .B1(new_n1183), .B2(new_n1184), .ZN(new_n1185));
  OR3_X1    g760(.A1(new_n1173), .A2(G1986), .A3(G290), .ZN(new_n1186));
  INV_X1    g761(.A(new_n1186), .ZN(new_n1187));
  XOR2_X1   g762(.A(KEYINPUT126), .B(KEYINPUT48), .Z(new_n1188));
  OR2_X1    g763(.A1(new_n1187), .A2(new_n1188), .ZN(new_n1189));
  AOI22_X1  g764(.A1(new_n1187), .A2(new_n1188), .B1(new_n1021), .B2(new_n1026), .ZN(new_n1190));
  AOI21_X1  g765(.A(new_n1185), .B1(new_n1189), .B2(new_n1190), .ZN(new_n1191));
  NAND2_X1  g766(.A1(new_n1178), .A2(new_n1179), .ZN(new_n1192));
  AND3_X1   g767(.A1(new_n1180), .A2(new_n1191), .A3(new_n1192), .ZN(new_n1193));
  NAND2_X1  g768(.A1(new_n1170), .A2(new_n1193), .ZN(G329));
  assign    G231 = 1'b0;
  AND2_X1   g769(.A1(new_n1001), .A2(KEYINPUT112), .ZN(new_n1196));
  NOR2_X1   g770(.A1(new_n1001), .A2(KEYINPUT112), .ZN(new_n1197));
  OAI211_X1 g771(.A(new_n1009), .B(new_n1008), .C1(new_n1196), .C2(new_n1197), .ZN(new_n1198));
  NAND3_X1  g772(.A1(new_n924), .A2(new_n926), .A3(new_n927), .ZN(new_n1199));
  INV_X1    g773(.A(KEYINPUT106), .ZN(new_n1200));
  NAND2_X1  g774(.A1(new_n1199), .A2(new_n1200), .ZN(new_n1201));
  NAND3_X1  g775(.A1(new_n929), .A2(KEYINPUT106), .A3(new_n926), .ZN(new_n1202));
  NAND2_X1  g776(.A1(new_n1201), .A2(new_n1202), .ZN(new_n1203));
  AOI21_X1  g777(.A(KEYINPUT107), .B1(new_n1203), .B2(new_n922), .ZN(new_n1204));
  INV_X1    g778(.A(new_n934), .ZN(new_n1205));
  OAI21_X1  g779(.A(new_n938), .B1(new_n1204), .B2(new_n1205), .ZN(new_n1206));
  AND3_X1   g780(.A1(new_n676), .A2(new_n679), .A3(G319), .ZN(new_n1207));
  NAND3_X1  g781(.A1(new_n659), .A2(new_n707), .A3(new_n1207), .ZN(new_n1208));
  INV_X1    g782(.A(KEYINPUT127), .ZN(new_n1209));
  NAND2_X1  g783(.A1(new_n1208), .A2(new_n1209), .ZN(new_n1210));
  NAND4_X1  g784(.A1(new_n659), .A2(new_n707), .A3(new_n1207), .A4(KEYINPUT127), .ZN(new_n1211));
  NAND2_X1  g785(.A1(new_n1210), .A2(new_n1211), .ZN(new_n1212));
  AND3_X1   g786(.A1(new_n1198), .A2(new_n1206), .A3(new_n1212), .ZN(G308));
  NAND3_X1  g787(.A1(new_n1198), .A2(new_n1206), .A3(new_n1212), .ZN(G225));
endmodule


