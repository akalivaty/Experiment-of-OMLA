//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 1 1 1 1 0 0 1 1 1 0 0 0 0 1 0 0 0 1 0 1 0 0 0 1 1 1 1 1 1 0 1 1 0 0 0 1 1 1 1 0 0 0 1 1 1 1 1 0 1 1 0 1 1 0 0 1 0 1 1 0 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:37:11 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n202, new_n203, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1247,
    new_n1248, new_n1249, new_n1250, new_n1251, new_n1252, new_n1253,
    new_n1254, new_n1255, new_n1256, new_n1257, new_n1258, new_n1259,
    new_n1260, new_n1261, new_n1262, new_n1263, new_n1264, new_n1265,
    new_n1266, new_n1267, new_n1268, new_n1269, new_n1270, new_n1271,
    new_n1272, new_n1274, new_n1275, new_n1276, new_n1277, new_n1279,
    new_n1280, new_n1281, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1346,
    new_n1347, new_n1348, new_n1349, new_n1350, new_n1351, new_n1352,
    new_n1353, new_n1354, new_n1355, new_n1356, new_n1357, new_n1358,
    new_n1359, new_n1361, new_n1362, new_n1363, new_n1364, new_n1365;
  NOR4_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .A4(G77), .ZN(G353));
  NOR2_X1   g0001(.A1(G97), .A2(G107), .ZN(new_n202));
  INV_X1    g0002(.A(new_n202), .ZN(new_n203));
  NAND2_X1  g0003(.A1(new_n203), .A2(G87), .ZN(G355));
  INV_X1    g0004(.A(G1), .ZN(new_n205));
  INV_X1    g0005(.A(G20), .ZN(new_n206));
  NOR2_X1   g0006(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  INV_X1    g0007(.A(new_n207), .ZN(new_n208));
  NOR2_X1   g0008(.A1(new_n208), .A2(G13), .ZN(new_n209));
  INV_X1    g0009(.A(new_n209), .ZN(new_n210));
  OAI21_X1  g0010(.A(G250), .B1(G257), .B2(G264), .ZN(new_n211));
  NOR2_X1   g0011(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  XNOR2_X1  g0012(.A(KEYINPUT64), .B(KEYINPUT0), .ZN(new_n213));
  NAND2_X1  g0013(.A1(G1), .A2(G13), .ZN(new_n214));
  NOR2_X1   g0014(.A1(new_n214), .A2(new_n206), .ZN(new_n215));
  OAI21_X1  g0015(.A(G50), .B1(G58), .B2(G68), .ZN(new_n216));
  INV_X1    g0016(.A(new_n216), .ZN(new_n217));
  AOI22_X1  g0017(.A1(new_n212), .A2(new_n213), .B1(new_n215), .B2(new_n217), .ZN(new_n218));
  OAI21_X1  g0018(.A(new_n218), .B1(new_n212), .B2(new_n213), .ZN(new_n219));
  AOI22_X1  g0019(.A1(G87), .A2(G250), .B1(G116), .B2(G270), .ZN(new_n220));
  INV_X1    g0020(.A(G58), .ZN(new_n221));
  INV_X1    g0021(.A(G232), .ZN(new_n222));
  INV_X1    g0022(.A(G97), .ZN(new_n223));
  INV_X1    g0023(.A(G257), .ZN(new_n224));
  OAI221_X1 g0024(.A(new_n220), .B1(new_n221), .B2(new_n222), .C1(new_n223), .C2(new_n224), .ZN(new_n225));
  AOI22_X1  g0025(.A1(G50), .A2(G226), .B1(G68), .B2(G238), .ZN(new_n226));
  AOI22_X1  g0026(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n227));
  NAND2_X1  g0027(.A1(new_n226), .A2(new_n227), .ZN(new_n228));
  OAI21_X1  g0028(.A(new_n208), .B1(new_n225), .B2(new_n228), .ZN(new_n229));
  XNOR2_X1  g0029(.A(new_n229), .B(KEYINPUT1), .ZN(new_n230));
  NOR2_X1   g0030(.A1(new_n219), .A2(new_n230), .ZN(G361));
  XOR2_X1   g0031(.A(G250), .B(G257), .Z(new_n232));
  XNOR2_X1  g0032(.A(G264), .B(G270), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n232), .B(new_n233), .ZN(new_n234));
  XNOR2_X1  g0034(.A(KEYINPUT65), .B(KEYINPUT66), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XNOR2_X1  g0036(.A(G238), .B(G244), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n237), .B(new_n222), .ZN(new_n238));
  XOR2_X1   g0038(.A(KEYINPUT2), .B(G226), .Z(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XOR2_X1   g0040(.A(new_n236), .B(new_n240), .Z(G358));
  XOR2_X1   g0041(.A(G68), .B(G77), .Z(new_n242));
  XOR2_X1   g0042(.A(G50), .B(G58), .Z(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XOR2_X1   g0044(.A(G87), .B(G97), .Z(new_n245));
  XNOR2_X1  g0045(.A(G107), .B(G116), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n245), .B(new_n246), .ZN(new_n247));
  XOR2_X1   g0047(.A(new_n244), .B(new_n247), .Z(G351));
  XNOR2_X1  g0048(.A(KEYINPUT3), .B(G33), .ZN(new_n249));
  INV_X1    g0049(.A(G1698), .ZN(new_n250));
  NAND3_X1  g0050(.A1(new_n249), .A2(G222), .A3(new_n250), .ZN(new_n251));
  NAND3_X1  g0051(.A1(new_n249), .A2(G223), .A3(G1698), .ZN(new_n252));
  INV_X1    g0052(.A(G77), .ZN(new_n253));
  OAI211_X1 g0053(.A(new_n251), .B(new_n252), .C1(new_n253), .C2(new_n249), .ZN(new_n254));
  NAND2_X1  g0054(.A1(G33), .A2(G41), .ZN(new_n255));
  NAND3_X1  g0055(.A1(new_n255), .A2(G1), .A3(G13), .ZN(new_n256));
  INV_X1    g0056(.A(new_n256), .ZN(new_n257));
  NAND2_X1  g0057(.A1(new_n254), .A2(new_n257), .ZN(new_n258));
  INV_X1    g0058(.A(G41), .ZN(new_n259));
  INV_X1    g0059(.A(G45), .ZN(new_n260));
  AOI21_X1  g0060(.A(G1), .B1(new_n259), .B2(new_n260), .ZN(new_n261));
  NAND3_X1  g0061(.A1(new_n261), .A2(new_n256), .A3(G274), .ZN(new_n262));
  INV_X1    g0062(.A(new_n262), .ZN(new_n263));
  NOR2_X1   g0063(.A1(new_n257), .A2(new_n261), .ZN(new_n264));
  AOI21_X1  g0064(.A(new_n263), .B1(G226), .B2(new_n264), .ZN(new_n265));
  AND2_X1   g0065(.A1(new_n258), .A2(new_n265), .ZN(new_n266));
  INV_X1    g0066(.A(G200), .ZN(new_n267));
  NOR2_X1   g0067(.A1(new_n266), .A2(new_n267), .ZN(new_n268));
  NAND3_X1  g0068(.A1(new_n205), .A2(G13), .A3(G20), .ZN(new_n269));
  INV_X1    g0069(.A(new_n269), .ZN(new_n270));
  NAND3_X1  g0070(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n271), .A2(new_n214), .ZN(new_n272));
  NOR2_X1   g0072(.A1(new_n270), .A2(new_n272), .ZN(new_n273));
  INV_X1    g0073(.A(G50), .ZN(new_n274));
  AOI21_X1  g0074(.A(new_n274), .B1(new_n205), .B2(G20), .ZN(new_n275));
  AOI22_X1  g0075(.A1(new_n273), .A2(new_n275), .B1(new_n274), .B2(new_n270), .ZN(new_n276));
  XNOR2_X1  g0076(.A(KEYINPUT8), .B(G58), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n206), .A2(G33), .ZN(new_n278));
  INV_X1    g0078(.A(G150), .ZN(new_n279));
  NOR2_X1   g0079(.A1(G20), .A2(G33), .ZN(new_n280));
  INV_X1    g0080(.A(new_n280), .ZN(new_n281));
  OAI22_X1  g0081(.A1(new_n277), .A2(new_n278), .B1(new_n279), .B2(new_n281), .ZN(new_n282));
  NOR2_X1   g0082(.A1(G50), .A2(G58), .ZN(new_n283));
  INV_X1    g0083(.A(G68), .ZN(new_n284));
  AOI21_X1  g0084(.A(new_n206), .B1(new_n283), .B2(new_n284), .ZN(new_n285));
  NOR2_X1   g0085(.A1(new_n282), .A2(new_n285), .ZN(new_n286));
  AND2_X1   g0086(.A1(new_n271), .A2(new_n214), .ZN(new_n287));
  OAI21_X1  g0087(.A(new_n276), .B1(new_n286), .B2(new_n287), .ZN(new_n288));
  INV_X1    g0088(.A(KEYINPUT9), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n288), .A2(new_n289), .ZN(new_n290));
  NAND3_X1  g0090(.A1(new_n258), .A2(G190), .A3(new_n265), .ZN(new_n291));
  OAI211_X1 g0091(.A(KEYINPUT9), .B(new_n276), .C1(new_n286), .C2(new_n287), .ZN(new_n292));
  NAND3_X1  g0092(.A1(new_n290), .A2(new_n291), .A3(new_n292), .ZN(new_n293));
  OR3_X1    g0093(.A1(new_n268), .A2(new_n293), .A3(KEYINPUT10), .ZN(new_n294));
  OAI21_X1  g0094(.A(KEYINPUT10), .B1(new_n268), .B2(new_n293), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n294), .A2(new_n295), .ZN(new_n296));
  AOI21_X1  g0096(.A(new_n263), .B1(G244), .B2(new_n264), .ZN(new_n297));
  AND2_X1   g0097(.A1(KEYINPUT3), .A2(G33), .ZN(new_n298));
  NOR2_X1   g0098(.A1(KEYINPUT3), .A2(G33), .ZN(new_n299));
  OAI211_X1 g0099(.A(G238), .B(G1698), .C1(new_n298), .C2(new_n299), .ZN(new_n300));
  OR2_X1    g0100(.A1(KEYINPUT3), .A2(G33), .ZN(new_n301));
  NAND2_X1  g0101(.A1(KEYINPUT3), .A2(G33), .ZN(new_n302));
  NAND3_X1  g0102(.A1(new_n301), .A2(G107), .A3(new_n302), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n300), .A2(new_n303), .ZN(new_n304));
  OAI211_X1 g0104(.A(G232), .B(new_n250), .C1(new_n298), .C2(new_n299), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n305), .A2(KEYINPUT67), .ZN(new_n306));
  INV_X1    g0106(.A(KEYINPUT67), .ZN(new_n307));
  NAND4_X1  g0107(.A1(new_n249), .A2(new_n307), .A3(G232), .A4(new_n250), .ZN(new_n308));
  AOI21_X1  g0108(.A(new_n304), .B1(new_n306), .B2(new_n308), .ZN(new_n309));
  OAI21_X1  g0109(.A(new_n257), .B1(new_n309), .B2(KEYINPUT68), .ZN(new_n310));
  INV_X1    g0110(.A(KEYINPUT68), .ZN(new_n311));
  AOI211_X1 g0111(.A(new_n311), .B(new_n304), .C1(new_n306), .C2(new_n308), .ZN(new_n312));
  OAI21_X1  g0112(.A(new_n297), .B1(new_n310), .B2(new_n312), .ZN(new_n313));
  AND2_X1   g0113(.A1(new_n313), .A2(G200), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n205), .A2(G20), .ZN(new_n315));
  NAND3_X1  g0115(.A1(new_n273), .A2(G77), .A3(new_n315), .ZN(new_n316));
  OAI21_X1  g0116(.A(new_n316), .B1(G77), .B2(new_n269), .ZN(new_n317));
  NAND2_X1  g0117(.A1(G20), .A2(G77), .ZN(new_n318));
  XOR2_X1   g0118(.A(KEYINPUT15), .B(G87), .Z(new_n319));
  INV_X1    g0119(.A(new_n319), .ZN(new_n320));
  OAI221_X1 g0120(.A(new_n318), .B1(new_n277), .B2(new_n281), .C1(new_n278), .C2(new_n320), .ZN(new_n321));
  AOI21_X1  g0121(.A(new_n317), .B1(new_n321), .B2(new_n272), .ZN(new_n322));
  INV_X1    g0122(.A(G190), .ZN(new_n323));
  OAI21_X1  g0123(.A(new_n322), .B1(new_n313), .B2(new_n323), .ZN(new_n324));
  OR2_X1    g0124(.A1(new_n314), .A2(new_n324), .ZN(new_n325));
  INV_X1    g0125(.A(G179), .ZN(new_n326));
  AND2_X1   g0126(.A1(new_n266), .A2(new_n326), .ZN(new_n327));
  OAI21_X1  g0127(.A(new_n288), .B1(new_n266), .B2(G169), .ZN(new_n328));
  OR2_X1    g0128(.A1(new_n327), .A2(new_n328), .ZN(new_n329));
  AND3_X1   g0129(.A1(new_n296), .A2(new_n325), .A3(new_n329), .ZN(new_n330));
  OR2_X1    g0130(.A1(new_n313), .A2(G179), .ZN(new_n331));
  INV_X1    g0131(.A(G169), .ZN(new_n332));
  AOI21_X1  g0132(.A(new_n322), .B1(new_n313), .B2(new_n332), .ZN(new_n333));
  INV_X1    g0133(.A(KEYINPUT69), .ZN(new_n334));
  OAI21_X1  g0134(.A(new_n331), .B1(new_n333), .B2(new_n334), .ZN(new_n335));
  AND2_X1   g0135(.A1(new_n333), .A2(new_n334), .ZN(new_n336));
  NOR2_X1   g0136(.A1(new_n335), .A2(new_n336), .ZN(new_n337));
  INV_X1    g0137(.A(new_n337), .ZN(new_n338));
  INV_X1    g0138(.A(G226), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n339), .A2(new_n250), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n222), .A2(G1698), .ZN(new_n341));
  OAI211_X1 g0141(.A(new_n340), .B(new_n341), .C1(new_n298), .C2(new_n299), .ZN(new_n342));
  NAND2_X1  g0142(.A1(G33), .A2(G97), .ZN(new_n343));
  NAND2_X1  g0143(.A1(new_n342), .A2(new_n343), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n344), .A2(new_n257), .ZN(new_n345));
  OAI21_X1  g0145(.A(new_n205), .B1(G41), .B2(G45), .ZN(new_n346));
  NAND3_X1  g0146(.A1(new_n256), .A2(G238), .A3(new_n346), .ZN(new_n347));
  AND2_X1   g0147(.A1(new_n262), .A2(new_n347), .ZN(new_n348));
  XNOR2_X1  g0148(.A(KEYINPUT70), .B(KEYINPUT13), .ZN(new_n349));
  NAND3_X1  g0149(.A1(new_n345), .A2(new_n348), .A3(new_n349), .ZN(new_n350));
  INV_X1    g0150(.A(new_n349), .ZN(new_n351));
  AOI21_X1  g0151(.A(new_n256), .B1(new_n342), .B2(new_n343), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n262), .A2(new_n347), .ZN(new_n353));
  OAI21_X1  g0153(.A(new_n351), .B1(new_n352), .B2(new_n353), .ZN(new_n354));
  AOI21_X1  g0154(.A(new_n267), .B1(new_n350), .B2(new_n354), .ZN(new_n355));
  OAI22_X1  g0155(.A1(new_n281), .A2(new_n274), .B1(new_n206), .B2(G68), .ZN(new_n356));
  NOR2_X1   g0156(.A1(new_n278), .A2(new_n253), .ZN(new_n357));
  OAI21_X1  g0157(.A(new_n272), .B1(new_n356), .B2(new_n357), .ZN(new_n358));
  XNOR2_X1  g0158(.A(new_n358), .B(KEYINPUT11), .ZN(new_n359));
  NOR2_X1   g0159(.A1(new_n269), .A2(G68), .ZN(new_n360));
  XNOR2_X1  g0160(.A(KEYINPUT71), .B(KEYINPUT12), .ZN(new_n361));
  NOR2_X1   g0161(.A1(new_n360), .A2(new_n361), .ZN(new_n362));
  INV_X1    g0162(.A(KEYINPUT12), .ZN(new_n363));
  AOI22_X1  g0163(.A1(new_n362), .A2(KEYINPUT72), .B1(new_n363), .B2(new_n360), .ZN(new_n364));
  OAI21_X1  g0164(.A(new_n364), .B1(KEYINPUT72), .B2(new_n362), .ZN(new_n365));
  NAND3_X1  g0165(.A1(new_n273), .A2(G68), .A3(new_n315), .ZN(new_n366));
  NAND3_X1  g0166(.A1(new_n359), .A2(new_n365), .A3(new_n366), .ZN(new_n367));
  OAI21_X1  g0167(.A(KEYINPUT13), .B1(new_n352), .B2(new_n353), .ZN(new_n368));
  AND2_X1   g0168(.A1(new_n350), .A2(new_n368), .ZN(new_n369));
  AOI211_X1 g0169(.A(new_n355), .B(new_n367), .C1(G190), .C2(new_n369), .ZN(new_n370));
  INV_X1    g0170(.A(KEYINPUT14), .ZN(new_n371));
  AOI21_X1  g0171(.A(new_n349), .B1(new_n345), .B2(new_n348), .ZN(new_n372));
  NOR3_X1   g0172(.A1(new_n352), .A2(new_n353), .A3(new_n351), .ZN(new_n373));
  OAI211_X1 g0173(.A(new_n371), .B(G169), .C1(new_n372), .C2(new_n373), .ZN(new_n374));
  NAND3_X1  g0174(.A1(new_n350), .A2(G179), .A3(new_n368), .ZN(new_n375));
  AND2_X1   g0175(.A1(new_n374), .A2(new_n375), .ZN(new_n376));
  INV_X1    g0176(.A(KEYINPUT73), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n350), .A2(new_n354), .ZN(new_n378));
  AOI21_X1  g0178(.A(new_n371), .B1(new_n378), .B2(G169), .ZN(new_n379));
  INV_X1    g0179(.A(new_n379), .ZN(new_n380));
  NAND3_X1  g0180(.A1(new_n376), .A2(new_n377), .A3(new_n380), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n374), .A2(new_n375), .ZN(new_n382));
  OAI21_X1  g0182(.A(KEYINPUT73), .B1(new_n382), .B2(new_n379), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n381), .A2(new_n383), .ZN(new_n384));
  XNOR2_X1  g0184(.A(new_n367), .B(KEYINPUT74), .ZN(new_n385));
  AOI21_X1  g0185(.A(new_n370), .B1(new_n384), .B2(new_n385), .ZN(new_n386));
  AOI21_X1  g0186(.A(new_n277), .B1(new_n205), .B2(G20), .ZN(new_n387));
  AOI22_X1  g0187(.A1(new_n387), .A2(new_n273), .B1(new_n277), .B2(new_n270), .ZN(new_n388));
  INV_X1    g0188(.A(new_n388), .ZN(new_n389));
  NOR2_X1   g0189(.A1(new_n298), .A2(new_n299), .ZN(new_n390));
  AOI21_X1  g0190(.A(KEYINPUT7), .B1(new_n390), .B2(new_n206), .ZN(new_n391));
  INV_X1    g0191(.A(KEYINPUT7), .ZN(new_n392));
  NOR4_X1   g0192(.A1(new_n298), .A2(new_n299), .A3(new_n392), .A4(G20), .ZN(new_n393));
  OAI21_X1  g0193(.A(G68), .B1(new_n391), .B2(new_n393), .ZN(new_n394));
  NOR2_X1   g0194(.A1(new_n221), .A2(new_n284), .ZN(new_n395));
  NOR2_X1   g0195(.A1(G58), .A2(G68), .ZN(new_n396));
  OAI21_X1  g0196(.A(G20), .B1(new_n395), .B2(new_n396), .ZN(new_n397));
  NAND2_X1  g0197(.A1(new_n280), .A2(G159), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n397), .A2(new_n398), .ZN(new_n399));
  INV_X1    g0199(.A(new_n399), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n394), .A2(new_n400), .ZN(new_n401));
  INV_X1    g0201(.A(KEYINPUT16), .ZN(new_n402));
  AOI21_X1  g0202(.A(new_n287), .B1(new_n401), .B2(new_n402), .ZN(new_n403));
  NAND3_X1  g0203(.A1(new_n394), .A2(KEYINPUT16), .A3(new_n400), .ZN(new_n404));
  AOI21_X1  g0204(.A(new_n389), .B1(new_n403), .B2(new_n404), .ZN(new_n405));
  OR2_X1    g0205(.A1(G223), .A2(G1698), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n339), .A2(G1698), .ZN(new_n407));
  OAI211_X1 g0207(.A(new_n406), .B(new_n407), .C1(new_n298), .C2(new_n299), .ZN(new_n408));
  NAND2_X1  g0208(.A1(G33), .A2(G87), .ZN(new_n409));
  AOI21_X1  g0209(.A(new_n256), .B1(new_n408), .B2(new_n409), .ZN(new_n410));
  INV_X1    g0210(.A(new_n410), .ZN(new_n411));
  NAND3_X1  g0211(.A1(new_n256), .A2(G232), .A3(new_n346), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n262), .A2(new_n412), .ZN(new_n413));
  INV_X1    g0213(.A(new_n413), .ZN(new_n414));
  NAND3_X1  g0214(.A1(new_n411), .A2(new_n414), .A3(new_n326), .ZN(new_n415));
  OAI21_X1  g0215(.A(new_n332), .B1(new_n410), .B2(new_n413), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n415), .A2(new_n416), .ZN(new_n417));
  OAI21_X1  g0217(.A(KEYINPUT18), .B1(new_n405), .B2(new_n417), .ZN(new_n418));
  NAND3_X1  g0218(.A1(new_n301), .A2(new_n206), .A3(new_n302), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n419), .A2(new_n392), .ZN(new_n420));
  NAND4_X1  g0220(.A1(new_n301), .A2(KEYINPUT7), .A3(new_n206), .A4(new_n302), .ZN(new_n421));
  AOI21_X1  g0221(.A(new_n284), .B1(new_n420), .B2(new_n421), .ZN(new_n422));
  OAI21_X1  g0222(.A(new_n402), .B1(new_n422), .B2(new_n399), .ZN(new_n423));
  NAND3_X1  g0223(.A1(new_n423), .A2(new_n404), .A3(new_n272), .ZN(new_n424));
  AOI21_X1  g0224(.A(new_n417), .B1(new_n424), .B2(new_n388), .ZN(new_n425));
  INV_X1    g0225(.A(KEYINPUT18), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n425), .A2(new_n426), .ZN(new_n427));
  NAND3_X1  g0227(.A1(new_n411), .A2(new_n414), .A3(new_n323), .ZN(new_n428));
  OAI21_X1  g0228(.A(new_n267), .B1(new_n410), .B2(new_n413), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n428), .A2(new_n429), .ZN(new_n430));
  NAND3_X1  g0230(.A1(new_n424), .A2(new_n430), .A3(new_n388), .ZN(new_n431));
  INV_X1    g0231(.A(KEYINPUT17), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n431), .A2(new_n432), .ZN(new_n433));
  NAND4_X1  g0233(.A1(new_n424), .A2(new_n430), .A3(KEYINPUT17), .A4(new_n388), .ZN(new_n434));
  NAND4_X1  g0234(.A1(new_n418), .A2(new_n427), .A3(new_n433), .A4(new_n434), .ZN(new_n435));
  INV_X1    g0235(.A(new_n435), .ZN(new_n436));
  NAND4_X1  g0236(.A1(new_n330), .A2(new_n338), .A3(new_n386), .A4(new_n436), .ZN(new_n437));
  NAND2_X1  g0237(.A1(new_n437), .A2(KEYINPUT75), .ZN(new_n438));
  AND4_X1   g0238(.A1(new_n436), .A2(new_n325), .A3(new_n296), .A4(new_n329), .ZN(new_n439));
  INV_X1    g0239(.A(KEYINPUT75), .ZN(new_n440));
  NAND4_X1  g0240(.A1(new_n439), .A2(new_n440), .A3(new_n338), .A4(new_n386), .ZN(new_n441));
  NAND2_X1  g0241(.A1(new_n438), .A2(new_n441), .ZN(new_n442));
  INV_X1    g0242(.A(new_n442), .ZN(new_n443));
  OAI211_X1 g0243(.A(G244), .B(G1698), .C1(new_n298), .C2(new_n299), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n444), .A2(KEYINPUT80), .ZN(new_n445));
  INV_X1    g0245(.A(KEYINPUT80), .ZN(new_n446));
  NAND4_X1  g0246(.A1(new_n249), .A2(new_n446), .A3(G244), .A4(G1698), .ZN(new_n447));
  NAND2_X1  g0247(.A1(G33), .A2(G116), .ZN(new_n448));
  NAND3_X1  g0248(.A1(new_n249), .A2(G238), .A3(new_n250), .ZN(new_n449));
  NAND4_X1  g0249(.A1(new_n445), .A2(new_n447), .A3(new_n448), .A4(new_n449), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n450), .A2(new_n257), .ZN(new_n451));
  NOR2_X1   g0251(.A1(new_n260), .A2(G1), .ZN(new_n452));
  INV_X1    g0252(.A(G274), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n452), .A2(new_n453), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n205), .A2(G45), .ZN(new_n455));
  INV_X1    g0255(.A(G250), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n455), .A2(new_n456), .ZN(new_n457));
  NAND3_X1  g0257(.A1(new_n454), .A2(new_n256), .A3(new_n457), .ZN(new_n458));
  NAND3_X1  g0258(.A1(new_n451), .A2(G190), .A3(new_n458), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n459), .A2(KEYINPUT83), .ZN(new_n460));
  INV_X1    g0260(.A(new_n458), .ZN(new_n461));
  AOI21_X1  g0261(.A(new_n461), .B1(new_n450), .B2(new_n257), .ZN(new_n462));
  INV_X1    g0262(.A(KEYINPUT83), .ZN(new_n463));
  NAND3_X1  g0263(.A1(new_n462), .A2(new_n463), .A3(G190), .ZN(new_n464));
  NAND2_X1  g0264(.A1(new_n460), .A2(new_n464), .ZN(new_n465));
  NOR2_X1   g0265(.A1(new_n319), .A2(new_n269), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n205), .A2(G33), .ZN(new_n467));
  NAND4_X1  g0267(.A1(new_n269), .A2(new_n467), .A3(new_n214), .A4(new_n271), .ZN(new_n468));
  INV_X1    g0268(.A(G87), .ZN(new_n469));
  NOR2_X1   g0269(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  INV_X1    g0270(.A(KEYINPUT19), .ZN(new_n471));
  OAI21_X1  g0271(.A(new_n206), .B1(new_n343), .B2(new_n471), .ZN(new_n472));
  OAI21_X1  g0272(.A(new_n472), .B1(G87), .B2(new_n203), .ZN(new_n473));
  OAI21_X1  g0273(.A(new_n471), .B1(new_n278), .B2(new_n223), .ZN(new_n474));
  OAI211_X1 g0274(.A(new_n206), .B(G68), .C1(new_n298), .C2(new_n299), .ZN(new_n475));
  NAND3_X1  g0275(.A1(new_n473), .A2(new_n474), .A3(new_n475), .ZN(new_n476));
  AOI211_X1 g0276(.A(new_n466), .B(new_n470), .C1(new_n476), .C2(new_n272), .ZN(new_n477));
  OAI21_X1  g0277(.A(new_n477), .B1(new_n462), .B2(new_n267), .ZN(new_n478));
  INV_X1    g0278(.A(KEYINPUT82), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n478), .A2(new_n479), .ZN(new_n480));
  OAI211_X1 g0280(.A(new_n477), .B(KEYINPUT82), .C1(new_n462), .C2(new_n267), .ZN(new_n481));
  NAND3_X1  g0281(.A1(new_n465), .A2(new_n480), .A3(new_n481), .ZN(new_n482));
  NOR2_X1   g0282(.A1(new_n462), .A2(new_n332), .ZN(new_n483));
  AOI211_X1 g0283(.A(new_n326), .B(new_n461), .C1(new_n450), .C2(new_n257), .ZN(new_n484));
  OAI21_X1  g0284(.A(KEYINPUT81), .B1(new_n483), .B2(new_n484), .ZN(new_n485));
  NAND3_X1  g0285(.A1(new_n451), .A2(G179), .A3(new_n458), .ZN(new_n486));
  INV_X1    g0286(.A(KEYINPUT81), .ZN(new_n487));
  OAI211_X1 g0287(.A(new_n486), .B(new_n487), .C1(new_n332), .C2(new_n462), .ZN(new_n488));
  AOI21_X1  g0288(.A(new_n466), .B1(new_n476), .B2(new_n272), .ZN(new_n489));
  OAI21_X1  g0289(.A(new_n489), .B1(new_n320), .B2(new_n468), .ZN(new_n490));
  NAND3_X1  g0290(.A1(new_n485), .A2(new_n488), .A3(new_n490), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n482), .A2(new_n491), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n270), .A2(new_n223), .ZN(new_n493));
  OAI21_X1  g0293(.A(new_n493), .B1(new_n468), .B2(new_n223), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n280), .A2(G77), .ZN(new_n495));
  INV_X1    g0295(.A(G107), .ZN(new_n496));
  AND3_X1   g0296(.A1(new_n496), .A2(KEYINPUT6), .A3(G97), .ZN(new_n497));
  XNOR2_X1  g0297(.A(G97), .B(G107), .ZN(new_n498));
  INV_X1    g0298(.A(KEYINPUT6), .ZN(new_n499));
  AOI21_X1  g0299(.A(new_n497), .B1(new_n498), .B2(new_n499), .ZN(new_n500));
  OAI21_X1  g0300(.A(new_n495), .B1(new_n500), .B2(new_n206), .ZN(new_n501));
  AOI21_X1  g0301(.A(new_n496), .B1(new_n420), .B2(new_n421), .ZN(new_n502));
  OAI21_X1  g0302(.A(new_n272), .B1(new_n501), .B2(new_n502), .ZN(new_n503));
  INV_X1    g0303(.A(KEYINPUT76), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  OAI21_X1  g0305(.A(G107), .B1(new_n391), .B2(new_n393), .ZN(new_n506));
  AND2_X1   g0306(.A1(G97), .A2(G107), .ZN(new_n507));
  OAI21_X1  g0307(.A(new_n499), .B1(new_n507), .B2(new_n202), .ZN(new_n508));
  NAND3_X1  g0308(.A1(new_n496), .A2(KEYINPUT6), .A3(G97), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  AOI22_X1  g0310(.A1(new_n510), .A2(G20), .B1(G77), .B2(new_n280), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n506), .A2(new_n511), .ZN(new_n512));
  NAND3_X1  g0312(.A1(new_n512), .A2(KEYINPUT76), .A3(new_n272), .ZN(new_n513));
  AOI21_X1  g0313(.A(new_n494), .B1(new_n505), .B2(new_n513), .ZN(new_n514));
  INV_X1    g0314(.A(KEYINPUT5), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n515), .A2(G41), .ZN(new_n516));
  NAND4_X1  g0316(.A1(new_n256), .A2(G274), .A3(new_n452), .A4(new_n516), .ZN(new_n517));
  INV_X1    g0317(.A(KEYINPUT78), .ZN(new_n518));
  OAI21_X1  g0318(.A(new_n518), .B1(new_n515), .B2(G41), .ZN(new_n519));
  NAND3_X1  g0319(.A1(new_n259), .A2(KEYINPUT78), .A3(KEYINPUT5), .ZN(new_n520));
  AND2_X1   g0320(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  OAI21_X1  g0321(.A(KEYINPUT79), .B1(new_n517), .B2(new_n521), .ZN(new_n522));
  INV_X1    g0322(.A(new_n214), .ZN(new_n523));
  AOI21_X1  g0323(.A(new_n453), .B1(new_n523), .B2(new_n255), .ZN(new_n524));
  OAI211_X1 g0324(.A(new_n205), .B(G45), .C1(new_n259), .C2(KEYINPUT5), .ZN(new_n525));
  INV_X1    g0325(.A(new_n525), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n519), .A2(new_n520), .ZN(new_n527));
  INV_X1    g0327(.A(KEYINPUT79), .ZN(new_n528));
  NAND4_X1  g0328(.A1(new_n524), .A2(new_n526), .A3(new_n527), .A4(new_n528), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n259), .A2(KEYINPUT5), .ZN(new_n530));
  NAND3_X1  g0330(.A1(new_n452), .A2(new_n530), .A3(new_n516), .ZN(new_n531));
  AND2_X1   g0331(.A1(new_n531), .A2(new_n256), .ZN(new_n532));
  AOI22_X1  g0332(.A1(new_n522), .A2(new_n529), .B1(new_n532), .B2(G257), .ZN(new_n533));
  OAI21_X1  g0333(.A(G244), .B1(new_n298), .B2(new_n299), .ZN(new_n534));
  INV_X1    g0334(.A(KEYINPUT4), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n534), .A2(new_n535), .ZN(new_n536));
  NOR2_X1   g0336(.A1(new_n535), .A2(G1698), .ZN(new_n537));
  NAND3_X1  g0337(.A1(new_n249), .A2(G244), .A3(new_n537), .ZN(new_n538));
  NAND2_X1  g0338(.A1(G33), .A2(G283), .ZN(new_n539));
  NAND3_X1  g0339(.A1(new_n536), .A2(new_n538), .A3(new_n539), .ZN(new_n540));
  OAI21_X1  g0340(.A(G250), .B1(new_n298), .B2(new_n299), .ZN(new_n541));
  AOI21_X1  g0341(.A(new_n250), .B1(new_n541), .B2(KEYINPUT4), .ZN(new_n542));
  OAI21_X1  g0342(.A(new_n257), .B1(new_n540), .B2(new_n542), .ZN(new_n543));
  AND2_X1   g0343(.A1(new_n533), .A2(new_n543), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n544), .A2(G190), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n522), .A2(new_n529), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n532), .A2(G257), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n546), .A2(new_n547), .ZN(new_n548));
  INV_X1    g0348(.A(KEYINPUT77), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n543), .A2(new_n549), .ZN(new_n550));
  OAI211_X1 g0350(.A(KEYINPUT77), .B(new_n257), .C1(new_n540), .C2(new_n542), .ZN(new_n551));
  AOI21_X1  g0351(.A(new_n548), .B1(new_n550), .B2(new_n551), .ZN(new_n552));
  OAI211_X1 g0352(.A(new_n514), .B(new_n545), .C1(new_n267), .C2(new_n552), .ZN(new_n553));
  INV_X1    g0353(.A(new_n494), .ZN(new_n554));
  AOI21_X1  g0354(.A(KEYINPUT76), .B1(new_n512), .B2(new_n272), .ZN(new_n555));
  AOI211_X1 g0355(.A(new_n504), .B(new_n287), .C1(new_n506), .C2(new_n511), .ZN(new_n556));
  OAI21_X1  g0356(.A(new_n554), .B1(new_n555), .B2(new_n556), .ZN(new_n557));
  INV_X1    g0357(.A(new_n551), .ZN(new_n558));
  AOI21_X1  g0358(.A(new_n456), .B1(new_n301), .B2(new_n302), .ZN(new_n559));
  OAI21_X1  g0359(.A(G1698), .B1(new_n559), .B2(new_n535), .ZN(new_n560));
  AOI22_X1  g0360(.A1(new_n534), .A2(new_n535), .B1(G33), .B2(G283), .ZN(new_n561));
  NAND3_X1  g0361(.A1(new_n560), .A2(new_n561), .A3(new_n538), .ZN(new_n562));
  AOI21_X1  g0362(.A(KEYINPUT77), .B1(new_n562), .B2(new_n257), .ZN(new_n563));
  OAI211_X1 g0363(.A(new_n326), .B(new_n533), .C1(new_n558), .C2(new_n563), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n533), .A2(new_n543), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n565), .A2(new_n332), .ZN(new_n566));
  NAND3_X1  g0366(.A1(new_n557), .A2(new_n564), .A3(new_n566), .ZN(new_n567));
  INV_X1    g0367(.A(G13), .ZN(new_n568));
  NOR2_X1   g0368(.A1(new_n568), .A2(G1), .ZN(new_n569));
  INV_X1    g0369(.A(KEYINPUT25), .ZN(new_n570));
  NAND4_X1  g0370(.A1(new_n569), .A2(new_n570), .A3(G20), .A4(new_n496), .ZN(new_n571));
  OAI21_X1  g0371(.A(KEYINPUT25), .B1(new_n269), .B2(G107), .ZN(new_n572));
  OAI211_X1 g0372(.A(new_n571), .B(new_n572), .C1(new_n468), .C2(new_n496), .ZN(new_n573));
  INV_X1    g0373(.A(KEYINPUT86), .ZN(new_n574));
  XNOR2_X1  g0374(.A(new_n573), .B(new_n574), .ZN(new_n575));
  OAI21_X1  g0375(.A(KEYINPUT23), .B1(new_n206), .B2(G107), .ZN(new_n576));
  INV_X1    g0376(.A(KEYINPUT23), .ZN(new_n577));
  NAND3_X1  g0377(.A1(new_n577), .A2(new_n496), .A3(G20), .ZN(new_n578));
  NAND3_X1  g0378(.A1(new_n206), .A2(G33), .A3(G116), .ZN(new_n579));
  NAND3_X1  g0379(.A1(new_n576), .A2(new_n578), .A3(new_n579), .ZN(new_n580));
  INV_X1    g0380(.A(KEYINPUT85), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  NAND4_X1  g0382(.A1(new_n576), .A2(new_n578), .A3(new_n579), .A4(KEYINPUT85), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  OAI211_X1 g0384(.A(new_n206), .B(G87), .C1(new_n298), .C2(new_n299), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n585), .A2(KEYINPUT22), .ZN(new_n586));
  INV_X1    g0386(.A(KEYINPUT22), .ZN(new_n587));
  NAND4_X1  g0387(.A1(new_n249), .A2(new_n587), .A3(new_n206), .A4(G87), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n586), .A2(new_n588), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n584), .A2(new_n589), .ZN(new_n590));
  INV_X1    g0390(.A(KEYINPUT24), .ZN(new_n591));
  AOI21_X1  g0391(.A(new_n287), .B1(new_n590), .B2(new_n591), .ZN(new_n592));
  AOI22_X1  g0392(.A1(new_n582), .A2(new_n583), .B1(new_n586), .B2(new_n588), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n593), .A2(KEYINPUT24), .ZN(new_n594));
  AOI21_X1  g0394(.A(new_n575), .B1(new_n592), .B2(new_n594), .ZN(new_n595));
  NOR2_X1   g0395(.A1(new_n515), .A2(G41), .ZN(new_n596));
  OAI211_X1 g0396(.A(G264), .B(new_n256), .C1(new_n525), .C2(new_n596), .ZN(new_n597));
  INV_X1    g0397(.A(KEYINPUT87), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n597), .A2(new_n598), .ZN(new_n599));
  NAND4_X1  g0399(.A1(new_n531), .A2(KEYINPUT87), .A3(G264), .A4(new_n256), .ZN(new_n600));
  OAI211_X1 g0400(.A(G257), .B(G1698), .C1(new_n298), .C2(new_n299), .ZN(new_n601));
  OAI211_X1 g0401(.A(G250), .B(new_n250), .C1(new_n298), .C2(new_n299), .ZN(new_n602));
  INV_X1    g0402(.A(G33), .ZN(new_n603));
  INV_X1    g0403(.A(G294), .ZN(new_n604));
  OAI211_X1 g0404(.A(new_n601), .B(new_n602), .C1(new_n603), .C2(new_n604), .ZN(new_n605));
  AOI22_X1  g0405(.A1(new_n599), .A2(new_n600), .B1(new_n605), .B2(new_n257), .ZN(new_n606));
  NAND3_X1  g0406(.A1(new_n606), .A2(G190), .A3(new_n546), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n605), .A2(new_n257), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n599), .A2(new_n600), .ZN(new_n609));
  NAND3_X1  g0409(.A1(new_n546), .A2(new_n608), .A3(new_n609), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n610), .A2(G200), .ZN(new_n611));
  NAND3_X1  g0411(.A1(new_n595), .A2(new_n607), .A3(new_n611), .ZN(new_n612));
  NAND3_X1  g0412(.A1(new_n553), .A2(new_n567), .A3(new_n612), .ZN(new_n613));
  AOI22_X1  g0413(.A1(new_n522), .A2(new_n529), .B1(new_n532), .B2(G270), .ZN(new_n614));
  OAI211_X1 g0414(.A(G264), .B(G1698), .C1(new_n298), .C2(new_n299), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n615), .A2(KEYINPUT84), .ZN(new_n616));
  INV_X1    g0416(.A(KEYINPUT84), .ZN(new_n617));
  NAND4_X1  g0417(.A1(new_n249), .A2(new_n617), .A3(G264), .A4(G1698), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n390), .A2(G303), .ZN(new_n619));
  NAND3_X1  g0419(.A1(new_n249), .A2(G257), .A3(new_n250), .ZN(new_n620));
  NAND4_X1  g0420(.A1(new_n616), .A2(new_n618), .A3(new_n619), .A4(new_n620), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n621), .A2(new_n257), .ZN(new_n622));
  AND3_X1   g0422(.A1(new_n614), .A2(G190), .A3(new_n622), .ZN(new_n623));
  AOI21_X1  g0423(.A(new_n267), .B1(new_n614), .B2(new_n622), .ZN(new_n624));
  OAI211_X1 g0424(.A(new_n539), .B(new_n206), .C1(G33), .C2(new_n223), .ZN(new_n625));
  INV_X1    g0425(.A(G116), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n626), .A2(G20), .ZN(new_n627));
  NAND3_X1  g0427(.A1(new_n625), .A2(new_n272), .A3(new_n627), .ZN(new_n628));
  INV_X1    g0428(.A(KEYINPUT20), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  NAND4_X1  g0430(.A1(new_n625), .A2(KEYINPUT20), .A3(new_n272), .A4(new_n627), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n630), .A2(new_n631), .ZN(new_n632));
  MUX2_X1   g0432(.A(new_n269), .B(new_n468), .S(G116), .Z(new_n633));
  NAND2_X1  g0433(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  OR3_X1    g0434(.A1(new_n623), .A2(new_n624), .A3(new_n634), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n614), .A2(new_n622), .ZN(new_n636));
  AOI21_X1  g0436(.A(new_n332), .B1(new_n632), .B2(new_n633), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n638), .A2(KEYINPUT21), .ZN(new_n639));
  INV_X1    g0439(.A(KEYINPUT21), .ZN(new_n640));
  NAND3_X1  g0440(.A1(new_n636), .A2(new_n640), .A3(new_n637), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n639), .A2(new_n641), .ZN(new_n642));
  AND2_X1   g0442(.A1(new_n614), .A2(new_n622), .ZN(new_n643));
  NAND3_X1  g0443(.A1(new_n643), .A2(G179), .A3(new_n634), .ZN(new_n644));
  XNOR2_X1  g0444(.A(new_n573), .B(KEYINPUT86), .ZN(new_n645));
  OAI21_X1  g0445(.A(new_n272), .B1(new_n593), .B2(KEYINPUT24), .ZN(new_n646));
  NOR2_X1   g0446(.A1(new_n590), .A2(new_n591), .ZN(new_n647));
  OAI21_X1  g0447(.A(new_n645), .B1(new_n646), .B2(new_n647), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n610), .A2(new_n332), .ZN(new_n649));
  NAND3_X1  g0449(.A1(new_n606), .A2(new_n326), .A3(new_n546), .ZN(new_n650));
  NAND3_X1  g0450(.A1(new_n648), .A2(new_n649), .A3(new_n650), .ZN(new_n651));
  NAND4_X1  g0451(.A1(new_n635), .A2(new_n642), .A3(new_n644), .A4(new_n651), .ZN(new_n652));
  NOR4_X1   g0452(.A1(new_n443), .A2(new_n492), .A3(new_n613), .A4(new_n652), .ZN(G372));
  INV_X1    g0453(.A(new_n329), .ZN(new_n654));
  AOI211_X1 g0454(.A(KEYINPUT18), .B(new_n417), .C1(new_n424), .C2(new_n388), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n424), .A2(new_n388), .ZN(new_n656));
  INV_X1    g0456(.A(new_n417), .ZN(new_n657));
  AOI21_X1  g0457(.A(new_n426), .B1(new_n656), .B2(new_n657), .ZN(new_n658));
  NOR2_X1   g0458(.A1(new_n655), .A2(new_n658), .ZN(new_n659));
  AOI21_X1  g0459(.A(new_n377), .B1(new_n376), .B2(new_n380), .ZN(new_n660));
  NOR3_X1   g0460(.A1(new_n382), .A2(KEYINPUT73), .A3(new_n379), .ZN(new_n661));
  OAI21_X1  g0461(.A(new_n385), .B1(new_n660), .B2(new_n661), .ZN(new_n662));
  INV_X1    g0462(.A(new_n662), .ZN(new_n663));
  INV_X1    g0463(.A(new_n370), .ZN(new_n664));
  AOI21_X1  g0464(.A(new_n663), .B1(new_n337), .B2(new_n664), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n433), .A2(new_n434), .ZN(new_n666));
  OAI21_X1  g0466(.A(new_n659), .B1(new_n665), .B2(new_n666), .ZN(new_n667));
  AOI21_X1  g0467(.A(new_n654), .B1(new_n667), .B2(new_n296), .ZN(new_n668));
  AND3_X1   g0468(.A1(new_n553), .A2(new_n567), .A3(new_n612), .ZN(new_n669));
  NAND3_X1  g0469(.A1(new_n642), .A2(new_n644), .A3(new_n651), .ZN(new_n670));
  INV_X1    g0470(.A(KEYINPUT88), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n478), .A2(new_n671), .ZN(new_n672));
  OAI211_X1 g0472(.A(new_n477), .B(KEYINPUT88), .C1(new_n462), .C2(new_n267), .ZN(new_n673));
  NAND3_X1  g0473(.A1(new_n465), .A2(new_n672), .A3(new_n673), .ZN(new_n674));
  OAI21_X1  g0474(.A(new_n490), .B1(new_n483), .B2(new_n484), .ZN(new_n675));
  AND2_X1   g0475(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  NAND3_X1  g0476(.A1(new_n669), .A2(new_n670), .A3(new_n676), .ZN(new_n677));
  AND3_X1   g0477(.A1(new_n557), .A2(new_n564), .A3(new_n566), .ZN(new_n678));
  AOI21_X1  g0478(.A(KEYINPUT26), .B1(new_n676), .B2(new_n678), .ZN(new_n679));
  NAND3_X1  g0479(.A1(new_n678), .A2(new_n482), .A3(new_n491), .ZN(new_n680));
  XOR2_X1   g0480(.A(KEYINPUT89), .B(KEYINPUT26), .Z(new_n681));
  NOR2_X1   g0481(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  OAI211_X1 g0482(.A(new_n677), .B(new_n675), .C1(new_n679), .C2(new_n682), .ZN(new_n683));
  INV_X1    g0483(.A(new_n683), .ZN(new_n684));
  OAI21_X1  g0484(.A(new_n668), .B1(new_n443), .B2(new_n684), .ZN(G369));
  NOR3_X1   g0485(.A1(new_n623), .A2(new_n624), .A3(new_n634), .ZN(new_n686));
  AND3_X1   g0486(.A1(new_n636), .A2(new_n640), .A3(new_n637), .ZN(new_n687));
  AOI21_X1  g0487(.A(new_n640), .B1(new_n636), .B2(new_n637), .ZN(new_n688));
  OAI21_X1  g0488(.A(new_n644), .B1(new_n687), .B2(new_n688), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n569), .A2(new_n206), .ZN(new_n690));
  OR2_X1    g0490(.A1(new_n690), .A2(KEYINPUT27), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n690), .A2(KEYINPUT27), .ZN(new_n692));
  NAND3_X1  g0492(.A1(new_n691), .A2(G213), .A3(new_n692), .ZN(new_n693));
  INV_X1    g0493(.A(new_n693), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n694), .A2(G343), .ZN(new_n695));
  INV_X1    g0495(.A(new_n695), .ZN(new_n696));
  NAND3_X1  g0496(.A1(new_n689), .A2(new_n634), .A3(new_n696), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n696), .A2(new_n634), .ZN(new_n698));
  NAND3_X1  g0498(.A1(new_n642), .A2(new_n644), .A3(new_n698), .ZN(new_n699));
  AOI21_X1  g0499(.A(new_n686), .B1(new_n697), .B2(new_n699), .ZN(new_n700));
  NAND2_X1  g0500(.A1(new_n700), .A2(G330), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n649), .A2(new_n650), .ZN(new_n702));
  NOR3_X1   g0502(.A1(new_n702), .A2(new_n595), .A3(new_n696), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n648), .A2(new_n696), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n612), .A2(new_n704), .ZN(new_n705));
  AOI21_X1  g0505(.A(new_n703), .B1(new_n705), .B2(new_n651), .ZN(new_n706));
  INV_X1    g0506(.A(new_n706), .ZN(new_n707));
  NOR2_X1   g0507(.A1(new_n701), .A2(new_n707), .ZN(new_n708));
  INV_X1    g0508(.A(new_n708), .ZN(new_n709));
  NAND2_X1  g0509(.A1(new_n689), .A2(new_n695), .ZN(new_n710));
  INV_X1    g0510(.A(KEYINPUT90), .ZN(new_n711));
  NAND2_X1  g0511(.A1(new_n710), .A2(new_n711), .ZN(new_n712));
  NAND3_X1  g0512(.A1(new_n689), .A2(KEYINPUT90), .A3(new_n695), .ZN(new_n713));
  NAND2_X1  g0513(.A1(new_n712), .A2(new_n713), .ZN(new_n714));
  AOI21_X1  g0514(.A(new_n703), .B1(new_n714), .B2(new_n706), .ZN(new_n715));
  NAND2_X1  g0515(.A1(new_n709), .A2(new_n715), .ZN(G399));
  NOR2_X1   g0516(.A1(new_n210), .A2(G41), .ZN(new_n717));
  INV_X1    g0517(.A(new_n717), .ZN(new_n718));
  NOR3_X1   g0518(.A1(new_n203), .A2(G87), .A3(G116), .ZN(new_n719));
  NAND3_X1  g0519(.A1(new_n718), .A2(G1), .A3(new_n719), .ZN(new_n720));
  OAI21_X1  g0520(.A(new_n720), .B1(new_n216), .B2(new_n718), .ZN(new_n721));
  XNOR2_X1  g0521(.A(new_n721), .B(KEYINPUT28), .ZN(new_n722));
  NAND4_X1  g0522(.A1(new_n484), .A2(new_n606), .A3(new_n622), .A4(new_n614), .ZN(new_n723));
  AND3_X1   g0523(.A1(new_n533), .A2(KEYINPUT30), .A3(new_n543), .ZN(new_n724));
  INV_X1    g0524(.A(new_n724), .ZN(new_n725));
  NAND2_X1  g0525(.A1(new_n451), .A2(new_n458), .ZN(new_n726));
  NAND4_X1  g0526(.A1(new_n636), .A2(new_n726), .A3(new_n326), .A4(new_n610), .ZN(new_n727));
  OAI22_X1  g0527(.A1(new_n723), .A2(new_n725), .B1(new_n727), .B2(new_n552), .ZN(new_n728));
  XNOR2_X1  g0528(.A(KEYINPUT91), .B(KEYINPUT30), .ZN(new_n729));
  NAND3_X1  g0529(.A1(new_n614), .A2(new_n606), .A3(new_n622), .ZN(new_n730));
  NOR2_X1   g0530(.A1(new_n730), .A2(new_n486), .ZN(new_n731));
  AOI21_X1  g0531(.A(new_n729), .B1(new_n731), .B2(new_n544), .ZN(new_n732));
  OAI211_X1 g0532(.A(KEYINPUT31), .B(new_n696), .C1(new_n728), .C2(new_n732), .ZN(new_n733));
  INV_X1    g0533(.A(new_n733), .ZN(new_n734));
  OAI21_X1  g0534(.A(new_n533), .B1(new_n558), .B2(new_n563), .ZN(new_n735));
  AOI21_X1  g0535(.A(G179), .B1(new_n606), .B2(new_n546), .ZN(new_n736));
  AOI21_X1  g0536(.A(new_n462), .B1(new_n622), .B2(new_n614), .ZN(new_n737));
  NAND3_X1  g0537(.A1(new_n735), .A2(new_n736), .A3(new_n737), .ZN(new_n738));
  NAND4_X1  g0538(.A1(new_n724), .A2(new_n643), .A3(new_n484), .A4(new_n606), .ZN(new_n739));
  NOR3_X1   g0539(.A1(new_n730), .A2(new_n486), .A3(new_n565), .ZN(new_n740));
  OAI211_X1 g0540(.A(new_n738), .B(new_n739), .C1(new_n740), .C2(new_n729), .ZN(new_n741));
  AOI21_X1  g0541(.A(KEYINPUT31), .B1(new_n741), .B2(new_n696), .ZN(new_n742));
  OAI21_X1  g0542(.A(KEYINPUT92), .B1(new_n734), .B2(new_n742), .ZN(new_n743));
  OAI21_X1  g0543(.A(new_n696), .B1(new_n728), .B2(new_n732), .ZN(new_n744));
  INV_X1    g0544(.A(KEYINPUT31), .ZN(new_n745));
  NAND2_X1  g0545(.A1(new_n744), .A2(new_n745), .ZN(new_n746));
  INV_X1    g0546(.A(KEYINPUT92), .ZN(new_n747));
  NAND3_X1  g0547(.A1(new_n746), .A2(new_n747), .A3(new_n733), .ZN(new_n748));
  NOR2_X1   g0548(.A1(new_n702), .A2(new_n595), .ZN(new_n749));
  NOR3_X1   g0549(.A1(new_n689), .A2(new_n749), .A3(new_n686), .ZN(new_n750));
  AND2_X1   g0550(.A1(new_n482), .A2(new_n491), .ZN(new_n751));
  NAND4_X1  g0551(.A1(new_n669), .A2(new_n750), .A3(new_n751), .A4(new_n695), .ZN(new_n752));
  NAND3_X1  g0552(.A1(new_n743), .A2(new_n748), .A3(new_n752), .ZN(new_n753));
  NAND2_X1  g0553(.A1(new_n753), .A2(G330), .ZN(new_n754));
  INV_X1    g0554(.A(new_n754), .ZN(new_n755));
  INV_X1    g0555(.A(KEYINPUT29), .ZN(new_n756));
  AND3_X1   g0556(.A1(new_n683), .A2(new_n756), .A3(new_n695), .ZN(new_n757));
  AND3_X1   g0557(.A1(new_n678), .A2(new_n482), .A3(new_n491), .ZN(new_n758));
  INV_X1    g0558(.A(new_n681), .ZN(new_n759));
  INV_X1    g0559(.A(KEYINPUT26), .ZN(new_n760));
  NAND3_X1  g0560(.A1(new_n678), .A2(new_n675), .A3(new_n674), .ZN(new_n761));
  OAI22_X1  g0561(.A1(new_n758), .A2(new_n759), .B1(new_n760), .B2(new_n761), .ZN(new_n762));
  NAND3_X1  g0562(.A1(new_n762), .A2(new_n675), .A3(new_n677), .ZN(new_n763));
  AOI21_X1  g0563(.A(new_n756), .B1(new_n763), .B2(new_n695), .ZN(new_n764));
  NOR3_X1   g0564(.A1(new_n755), .A2(new_n757), .A3(new_n764), .ZN(new_n765));
  OAI21_X1  g0565(.A(new_n722), .B1(new_n765), .B2(G1), .ZN(G364));
  INV_X1    g0566(.A(new_n701), .ZN(new_n767));
  NOR2_X1   g0567(.A1(new_n568), .A2(G20), .ZN(new_n768));
  AOI21_X1  g0568(.A(new_n205), .B1(new_n768), .B2(G45), .ZN(new_n769));
  INV_X1    g0569(.A(new_n769), .ZN(new_n770));
  NOR2_X1   g0570(.A1(new_n717), .A2(new_n770), .ZN(new_n771));
  NOR2_X1   g0571(.A1(new_n767), .A2(new_n771), .ZN(new_n772));
  NOR2_X1   g0572(.A1(new_n700), .A2(G330), .ZN(new_n773));
  INV_X1    g0573(.A(new_n773), .ZN(new_n774));
  NOR2_X1   g0574(.A1(G13), .A2(G33), .ZN(new_n775));
  INV_X1    g0575(.A(new_n775), .ZN(new_n776));
  NOR2_X1   g0576(.A1(new_n776), .A2(G20), .ZN(new_n777));
  INV_X1    g0577(.A(new_n777), .ZN(new_n778));
  OR2_X1    g0578(.A1(new_n700), .A2(new_n778), .ZN(new_n779));
  NOR2_X1   g0579(.A1(new_n210), .A2(new_n390), .ZN(new_n780));
  NAND2_X1  g0580(.A1(new_n780), .A2(G355), .ZN(new_n781));
  OAI21_X1  g0581(.A(new_n781), .B1(G116), .B2(new_n209), .ZN(new_n782));
  NOR2_X1   g0582(.A1(new_n210), .A2(new_n249), .ZN(new_n783));
  INV_X1    g0583(.A(new_n783), .ZN(new_n784));
  AOI21_X1  g0584(.A(new_n784), .B1(new_n260), .B2(new_n217), .ZN(new_n785));
  NAND2_X1  g0585(.A1(new_n244), .A2(G45), .ZN(new_n786));
  AOI21_X1  g0586(.A(new_n782), .B1(new_n785), .B2(new_n786), .ZN(new_n787));
  AOI21_X1  g0587(.A(new_n214), .B1(G20), .B2(new_n332), .ZN(new_n788));
  NOR2_X1   g0588(.A1(new_n777), .A2(new_n788), .ZN(new_n789));
  INV_X1    g0589(.A(new_n789), .ZN(new_n790));
  OAI21_X1  g0590(.A(new_n771), .B1(new_n787), .B2(new_n790), .ZN(new_n791));
  NOR2_X1   g0591(.A1(new_n206), .A2(G190), .ZN(new_n792));
  NOR2_X1   g0592(.A1(new_n267), .A2(G179), .ZN(new_n793));
  NAND2_X1  g0593(.A1(new_n792), .A2(new_n793), .ZN(new_n794));
  INV_X1    g0594(.A(G283), .ZN(new_n795));
  OAI21_X1  g0595(.A(new_n390), .B1(new_n794), .B2(new_n795), .ZN(new_n796));
  NOR2_X1   g0596(.A1(new_n206), .A2(new_n326), .ZN(new_n797));
  NAND2_X1  g0597(.A1(new_n797), .A2(G190), .ZN(new_n798));
  NOR2_X1   g0598(.A1(new_n798), .A2(G200), .ZN(new_n799));
  AOI21_X1  g0599(.A(new_n796), .B1(G322), .B2(new_n799), .ZN(new_n800));
  NAND3_X1  g0600(.A1(new_n797), .A2(new_n323), .A3(new_n267), .ZN(new_n801));
  INV_X1    g0601(.A(new_n801), .ZN(new_n802));
  NAND3_X1  g0602(.A1(new_n793), .A2(G20), .A3(G190), .ZN(new_n803));
  INV_X1    g0603(.A(new_n803), .ZN(new_n804));
  AOI22_X1  g0604(.A1(G311), .A2(new_n802), .B1(new_n804), .B2(G303), .ZN(new_n805));
  NOR2_X1   g0605(.A1(new_n798), .A2(new_n267), .ZN(new_n806));
  NOR2_X1   g0606(.A1(G179), .A2(G200), .ZN(new_n807));
  AOI21_X1  g0607(.A(new_n206), .B1(new_n807), .B2(G190), .ZN(new_n808));
  INV_X1    g0608(.A(new_n808), .ZN(new_n809));
  AOI22_X1  g0609(.A1(new_n806), .A2(G326), .B1(G294), .B2(new_n809), .ZN(new_n810));
  NAND3_X1  g0610(.A1(new_n792), .A2(G179), .A3(G200), .ZN(new_n811));
  INV_X1    g0611(.A(new_n811), .ZN(new_n812));
  XNOR2_X1  g0612(.A(KEYINPUT33), .B(G317), .ZN(new_n813));
  NAND2_X1  g0613(.A1(new_n792), .A2(new_n807), .ZN(new_n814));
  INV_X1    g0614(.A(new_n814), .ZN(new_n815));
  AOI22_X1  g0615(.A1(new_n812), .A2(new_n813), .B1(new_n815), .B2(G329), .ZN(new_n816));
  NAND4_X1  g0616(.A1(new_n800), .A2(new_n805), .A3(new_n810), .A4(new_n816), .ZN(new_n817));
  OAI221_X1 g0617(.A(new_n249), .B1(new_n794), .B2(new_n496), .C1(new_n469), .C2(new_n803), .ZN(new_n818));
  XNOR2_X1  g0618(.A(new_n818), .B(KEYINPUT93), .ZN(new_n819));
  AOI22_X1  g0619(.A1(G50), .A2(new_n806), .B1(new_n799), .B2(G58), .ZN(new_n820));
  INV_X1    g0620(.A(G159), .ZN(new_n821));
  OAI21_X1  g0621(.A(KEYINPUT32), .B1(new_n814), .B2(new_n821), .ZN(new_n822));
  AOI22_X1  g0622(.A1(G77), .A2(new_n802), .B1(new_n812), .B2(G68), .ZN(new_n823));
  NOR3_X1   g0623(.A1(new_n814), .A2(KEYINPUT32), .A3(new_n821), .ZN(new_n824));
  NOR2_X1   g0624(.A1(new_n808), .A2(new_n223), .ZN(new_n825));
  NOR2_X1   g0625(.A1(new_n824), .A2(new_n825), .ZN(new_n826));
  NAND4_X1  g0626(.A1(new_n820), .A2(new_n822), .A3(new_n823), .A4(new_n826), .ZN(new_n827));
  OAI21_X1  g0627(.A(new_n817), .B1(new_n819), .B2(new_n827), .ZN(new_n828));
  AOI21_X1  g0628(.A(new_n791), .B1(new_n828), .B2(new_n788), .ZN(new_n829));
  AOI22_X1  g0629(.A1(new_n772), .A2(new_n774), .B1(new_n779), .B2(new_n829), .ZN(new_n830));
  INV_X1    g0630(.A(new_n830), .ZN(G396));
  OR2_X1    g0631(.A1(new_n322), .A2(new_n695), .ZN(new_n832));
  OAI21_X1  g0632(.A(new_n832), .B1(new_n314), .B2(new_n324), .ZN(new_n833));
  OAI21_X1  g0633(.A(new_n833), .B1(new_n335), .B2(new_n336), .ZN(new_n834));
  AND2_X1   g0634(.A1(new_n313), .A2(new_n332), .ZN(new_n835));
  OAI21_X1  g0635(.A(KEYINPUT69), .B1(new_n835), .B2(new_n322), .ZN(new_n836));
  NAND2_X1  g0636(.A1(new_n333), .A2(new_n334), .ZN(new_n837));
  NAND4_X1  g0637(.A1(new_n836), .A2(new_n837), .A3(new_n331), .A4(new_n832), .ZN(new_n838));
  AND2_X1   g0638(.A1(new_n834), .A2(new_n838), .ZN(new_n839));
  AOI21_X1  g0639(.A(new_n839), .B1(new_n683), .B2(new_n695), .ZN(new_n840));
  AND3_X1   g0640(.A1(new_n834), .A2(new_n838), .A3(new_n695), .ZN(new_n841));
  AOI21_X1  g0641(.A(new_n840), .B1(new_n683), .B2(new_n841), .ZN(new_n842));
  AND2_X1   g0642(.A1(new_n842), .A2(new_n755), .ZN(new_n843));
  NOR2_X1   g0643(.A1(new_n842), .A2(new_n755), .ZN(new_n844));
  AOI211_X1 g0644(.A(new_n771), .B(new_n843), .C1(new_n844), .C2(KEYINPUT97), .ZN(new_n845));
  OAI21_X1  g0645(.A(new_n845), .B1(KEYINPUT97), .B2(new_n844), .ZN(new_n846));
  INV_X1    g0646(.A(new_n771), .ZN(new_n847));
  NOR2_X1   g0647(.A1(new_n788), .A2(new_n775), .ZN(new_n848));
  XOR2_X1   g0648(.A(new_n848), .B(KEYINPUT94), .Z(new_n849));
  INV_X1    g0649(.A(new_n849), .ZN(new_n850));
  AOI21_X1  g0650(.A(new_n847), .B1(new_n850), .B2(new_n253), .ZN(new_n851));
  INV_X1    g0651(.A(new_n794), .ZN(new_n852));
  AOI22_X1  g0652(.A1(new_n852), .A2(G87), .B1(new_n815), .B2(G311), .ZN(new_n853));
  OAI221_X1 g0653(.A(new_n853), .B1(new_n496), .B2(new_n803), .C1(new_n626), .C2(new_n801), .ZN(new_n854));
  INV_X1    g0654(.A(new_n799), .ZN(new_n855));
  INV_X1    g0655(.A(new_n806), .ZN(new_n856));
  INV_X1    g0656(.A(G303), .ZN(new_n857));
  OAI22_X1  g0657(.A1(new_n855), .A2(new_n604), .B1(new_n856), .B2(new_n857), .ZN(new_n858));
  OAI21_X1  g0658(.A(new_n390), .B1(new_n811), .B2(new_n795), .ZN(new_n859));
  NOR4_X1   g0659(.A1(new_n854), .A2(new_n825), .A3(new_n858), .A4(new_n859), .ZN(new_n860));
  XOR2_X1   g0660(.A(new_n860), .B(KEYINPUT95), .Z(new_n861));
  AOI22_X1  g0661(.A1(G159), .A2(new_n802), .B1(new_n812), .B2(G150), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n799), .A2(G143), .ZN(new_n863));
  INV_X1    g0663(.A(G137), .ZN(new_n864));
  OAI211_X1 g0664(.A(new_n862), .B(new_n863), .C1(new_n864), .C2(new_n856), .ZN(new_n865));
  XOR2_X1   g0665(.A(new_n865), .B(KEYINPUT34), .Z(new_n866));
  OR2_X1    g0666(.A1(new_n866), .A2(KEYINPUT96), .ZN(new_n867));
  AOI22_X1  g0667(.A1(new_n804), .A2(G50), .B1(new_n852), .B2(G68), .ZN(new_n868));
  AOI21_X1  g0668(.A(new_n390), .B1(new_n815), .B2(G132), .ZN(new_n869));
  OAI211_X1 g0669(.A(new_n868), .B(new_n869), .C1(new_n221), .C2(new_n808), .ZN(new_n870));
  AOI21_X1  g0670(.A(new_n870), .B1(new_n866), .B2(KEYINPUT96), .ZN(new_n871));
  AOI21_X1  g0671(.A(new_n861), .B1(new_n867), .B2(new_n871), .ZN(new_n872));
  INV_X1    g0672(.A(new_n788), .ZN(new_n873));
  OAI221_X1 g0673(.A(new_n851), .B1(new_n872), .B2(new_n873), .C1(new_n839), .C2(new_n776), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n846), .A2(new_n874), .ZN(G384));
  OR2_X1    g0675(.A1(new_n510), .A2(KEYINPUT35), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n510), .A2(KEYINPUT35), .ZN(new_n877));
  NAND4_X1  g0677(.A1(new_n876), .A2(new_n877), .A3(G116), .A4(new_n215), .ZN(new_n878));
  XOR2_X1   g0678(.A(new_n878), .B(KEYINPUT36), .Z(new_n879));
  OAI211_X1 g0679(.A(new_n217), .B(G77), .C1(new_n221), .C2(new_n284), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n274), .A2(G68), .ZN(new_n881));
  AOI211_X1 g0681(.A(new_n205), .B(G13), .C1(new_n880), .C2(new_n881), .ZN(new_n882));
  NOR2_X1   g0682(.A1(new_n879), .A2(new_n882), .ZN(new_n883));
  INV_X1    g0683(.A(KEYINPUT98), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n656), .A2(new_n657), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n656), .A2(new_n694), .ZN(new_n886));
  NAND3_X1  g0686(.A1(new_n885), .A2(new_n886), .A3(new_n431), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n887), .A2(KEYINPUT37), .ZN(new_n888));
  INV_X1    g0688(.A(KEYINPUT37), .ZN(new_n889));
  NAND4_X1  g0689(.A1(new_n885), .A2(new_n886), .A3(new_n889), .A4(new_n431), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n888), .A2(new_n890), .ZN(new_n891));
  INV_X1    g0691(.A(new_n886), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n435), .A2(new_n892), .ZN(new_n893));
  AND3_X1   g0693(.A1(new_n891), .A2(new_n893), .A3(KEYINPUT38), .ZN(new_n894));
  AOI21_X1  g0694(.A(KEYINPUT38), .B1(new_n891), .B2(new_n893), .ZN(new_n895));
  OAI21_X1  g0695(.A(new_n884), .B1(new_n894), .B2(new_n895), .ZN(new_n896));
  INV_X1    g0696(.A(KEYINPUT38), .ZN(new_n897));
  AND3_X1   g0697(.A1(new_n424), .A2(new_n388), .A3(new_n430), .ZN(new_n898));
  NOR2_X1   g0698(.A1(new_n898), .A2(new_n425), .ZN(new_n899));
  AOI21_X1  g0699(.A(new_n889), .B1(new_n899), .B2(new_n886), .ZN(new_n900));
  AND4_X1   g0700(.A1(new_n889), .A2(new_n885), .A3(new_n886), .A4(new_n431), .ZN(new_n901));
  NOR2_X1   g0701(.A1(new_n900), .A2(new_n901), .ZN(new_n902));
  INV_X1    g0702(.A(new_n666), .ZN(new_n903));
  AOI21_X1  g0703(.A(new_n886), .B1(new_n903), .B2(new_n659), .ZN(new_n904));
  OAI21_X1  g0704(.A(new_n897), .B1(new_n902), .B2(new_n904), .ZN(new_n905));
  NAND3_X1  g0705(.A1(new_n891), .A2(new_n893), .A3(KEYINPUT38), .ZN(new_n906));
  NAND3_X1  g0706(.A1(new_n905), .A2(KEYINPUT98), .A3(new_n906), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n896), .A2(new_n907), .ZN(new_n908));
  NAND3_X1  g0708(.A1(new_n752), .A2(new_n746), .A3(new_n733), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n385), .A2(new_n696), .ZN(new_n910));
  NAND3_X1  g0710(.A1(new_n662), .A2(new_n664), .A3(new_n910), .ZN(new_n911));
  OAI211_X1 g0711(.A(new_n385), .B(new_n696), .C1(new_n384), .C2(new_n370), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n911), .A2(new_n912), .ZN(new_n913));
  AND3_X1   g0713(.A1(new_n909), .A2(new_n839), .A3(new_n913), .ZN(new_n914));
  AOI21_X1  g0714(.A(KEYINPUT40), .B1(new_n908), .B2(new_n914), .ZN(new_n915));
  INV_X1    g0715(.A(new_n915), .ZN(new_n916));
  INV_X1    g0716(.A(KEYINPUT40), .ZN(new_n917));
  AOI21_X1  g0717(.A(new_n917), .B1(new_n905), .B2(new_n906), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n914), .A2(new_n918), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n916), .A2(new_n919), .ZN(new_n920));
  INV_X1    g0720(.A(new_n909), .ZN(new_n921));
  NOR3_X1   g0721(.A1(new_n920), .A2(new_n443), .A3(new_n921), .ZN(new_n922));
  INV_X1    g0722(.A(G330), .ZN(new_n923));
  AOI22_X1  g0723(.A1(new_n916), .A2(new_n919), .B1(new_n442), .B2(new_n909), .ZN(new_n924));
  NOR3_X1   g0724(.A1(new_n922), .A2(new_n923), .A3(new_n924), .ZN(new_n925));
  AND3_X1   g0725(.A1(new_n905), .A2(KEYINPUT39), .A3(new_n906), .ZN(new_n926));
  AOI21_X1  g0726(.A(KEYINPUT39), .B1(new_n905), .B2(new_n906), .ZN(new_n927));
  OR2_X1    g0727(.A1(new_n926), .A2(new_n927), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n663), .A2(new_n695), .ZN(new_n929));
  INV_X1    g0729(.A(KEYINPUT99), .ZN(new_n930));
  XNOR2_X1  g0730(.A(new_n929), .B(new_n930), .ZN(new_n931));
  OAI22_X1  g0731(.A1(new_n928), .A2(new_n931), .B1(new_n659), .B2(new_n694), .ZN(new_n932));
  INV_X1    g0732(.A(new_n913), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n677), .A2(new_n675), .ZN(new_n934));
  AOI22_X1  g0734(.A1(new_n758), .A2(new_n759), .B1(new_n761), .B2(new_n760), .ZN(new_n935));
  OAI21_X1  g0735(.A(new_n841), .B1(new_n934), .B2(new_n935), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n337), .A2(new_n695), .ZN(new_n937));
  AOI21_X1  g0737(.A(new_n933), .B1(new_n936), .B2(new_n937), .ZN(new_n938));
  AND2_X1   g0738(.A1(new_n938), .A2(new_n908), .ZN(new_n939));
  NOR2_X1   g0739(.A1(new_n932), .A2(new_n939), .ZN(new_n940));
  OAI21_X1  g0740(.A(new_n442), .B1(new_n757), .B2(new_n764), .ZN(new_n941));
  NAND2_X1  g0741(.A1(new_n941), .A2(new_n668), .ZN(new_n942));
  XNOR2_X1  g0742(.A(new_n940), .B(new_n942), .ZN(new_n943));
  OAI22_X1  g0743(.A1(new_n925), .A2(new_n943), .B1(new_n205), .B2(new_n768), .ZN(new_n944));
  AND2_X1   g0744(.A1(new_n925), .A2(new_n943), .ZN(new_n945));
  OAI21_X1  g0745(.A(new_n883), .B1(new_n944), .B2(new_n945), .ZN(G367));
  OAI211_X1 g0746(.A(new_n553), .B(new_n567), .C1(new_n514), .C2(new_n695), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n678), .A2(new_n696), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n947), .A2(new_n948), .ZN(new_n949));
  INV_X1    g0749(.A(new_n949), .ZN(new_n950));
  AND3_X1   g0750(.A1(new_n689), .A2(KEYINPUT90), .A3(new_n695), .ZN(new_n951));
  AOI21_X1  g0751(.A(KEYINPUT90), .B1(new_n689), .B2(new_n695), .ZN(new_n952));
  OAI21_X1  g0752(.A(new_n706), .B1(new_n951), .B2(new_n952), .ZN(new_n953));
  NOR2_X1   g0753(.A1(new_n950), .A2(new_n953), .ZN(new_n954));
  XNOR2_X1  g0754(.A(new_n954), .B(KEYINPUT42), .ZN(new_n955));
  OR2_X1    g0755(.A1(new_n695), .A2(new_n477), .ZN(new_n956));
  NAND2_X1  g0756(.A1(new_n676), .A2(new_n956), .ZN(new_n957));
  OR2_X1    g0757(.A1(new_n675), .A2(new_n956), .ZN(new_n958));
  OR2_X1    g0758(.A1(new_n958), .A2(KEYINPUT100), .ZN(new_n959));
  NAND2_X1  g0759(.A1(new_n958), .A2(KEYINPUT100), .ZN(new_n960));
  NAND3_X1  g0760(.A1(new_n957), .A2(new_n959), .A3(new_n960), .ZN(new_n961));
  AND2_X1   g0761(.A1(new_n961), .A2(KEYINPUT101), .ZN(new_n962));
  NOR2_X1   g0762(.A1(new_n961), .A2(KEYINPUT101), .ZN(new_n963));
  NOR3_X1   g0763(.A1(new_n962), .A2(new_n963), .A3(KEYINPUT43), .ZN(new_n964));
  OAI21_X1  g0764(.A(new_n567), .B1(new_n947), .B2(new_n651), .ZN(new_n965));
  NAND2_X1  g0765(.A1(new_n965), .A2(new_n695), .ZN(new_n966));
  NAND3_X1  g0766(.A1(new_n955), .A2(new_n964), .A3(new_n966), .ZN(new_n967));
  XNOR2_X1  g0767(.A(new_n967), .B(KEYINPUT102), .ZN(new_n968));
  NOR2_X1   g0768(.A1(new_n709), .A2(new_n950), .ZN(new_n969));
  AOI21_X1  g0769(.A(new_n964), .B1(KEYINPUT43), .B2(new_n961), .ZN(new_n970));
  NAND2_X1  g0770(.A1(new_n955), .A2(new_n966), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n970), .A2(new_n971), .ZN(new_n972));
  NAND3_X1  g0772(.A1(new_n968), .A2(new_n969), .A3(new_n972), .ZN(new_n973));
  INV_X1    g0773(.A(new_n973), .ZN(new_n974));
  AOI21_X1  g0774(.A(new_n969), .B1(new_n968), .B2(new_n972), .ZN(new_n975));
  NOR2_X1   g0775(.A1(new_n974), .A2(new_n975), .ZN(new_n976));
  XOR2_X1   g0776(.A(new_n717), .B(KEYINPUT41), .Z(new_n977));
  NOR2_X1   g0777(.A1(new_n757), .A2(new_n764), .ZN(new_n978));
  NAND3_X1  g0778(.A1(new_n707), .A2(new_n712), .A3(new_n713), .ZN(new_n979));
  AND3_X1   g0779(.A1(new_n767), .A2(new_n953), .A3(new_n979), .ZN(new_n980));
  AOI21_X1  g0780(.A(new_n767), .B1(new_n953), .B2(new_n979), .ZN(new_n981));
  NOR2_X1   g0781(.A1(new_n980), .A2(new_n981), .ZN(new_n982));
  AND3_X1   g0782(.A1(new_n978), .A2(new_n754), .A3(new_n982), .ZN(new_n983));
  INV_X1    g0783(.A(KEYINPUT45), .ZN(new_n984));
  INV_X1    g0784(.A(new_n703), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n953), .A2(new_n985), .ZN(new_n986));
  OAI21_X1  g0786(.A(new_n984), .B1(new_n986), .B2(new_n950), .ZN(new_n987));
  NAND3_X1  g0787(.A1(new_n715), .A2(KEYINPUT45), .A3(new_n949), .ZN(new_n988));
  NAND2_X1  g0788(.A1(new_n987), .A2(new_n988), .ZN(new_n989));
  XOR2_X1   g0789(.A(KEYINPUT103), .B(KEYINPUT44), .Z(new_n990));
  NAND3_X1  g0790(.A1(new_n986), .A2(new_n950), .A3(new_n990), .ZN(new_n991));
  INV_X1    g0791(.A(new_n990), .ZN(new_n992));
  OAI21_X1  g0792(.A(new_n992), .B1(new_n715), .B2(new_n949), .ZN(new_n993));
  NAND4_X1  g0793(.A1(new_n989), .A2(KEYINPUT104), .A3(new_n991), .A4(new_n993), .ZN(new_n994));
  INV_X1    g0794(.A(KEYINPUT105), .ZN(new_n995));
  AOI21_X1  g0795(.A(new_n709), .B1(new_n994), .B2(new_n995), .ZN(new_n996));
  AOI21_X1  g0796(.A(KEYINPUT45), .B1(new_n715), .B2(new_n949), .ZN(new_n997));
  AND4_X1   g0797(.A1(KEYINPUT45), .A2(new_n953), .A3(new_n985), .A4(new_n949), .ZN(new_n998));
  OAI211_X1 g0798(.A(new_n991), .B(new_n993), .C1(new_n997), .C2(new_n998), .ZN(new_n999));
  OAI21_X1  g0799(.A(KEYINPUT104), .B1(new_n708), .B2(KEYINPUT105), .ZN(new_n1000));
  NAND2_X1  g0800(.A1(new_n999), .A2(new_n1000), .ZN(new_n1001));
  INV_X1    g0801(.A(new_n1001), .ZN(new_n1002));
  OAI21_X1  g0802(.A(new_n983), .B1(new_n996), .B2(new_n1002), .ZN(new_n1003));
  AOI21_X1  g0803(.A(new_n977), .B1(new_n1003), .B2(new_n765), .ZN(new_n1004));
  INV_X1    g0804(.A(KEYINPUT106), .ZN(new_n1005));
  OAI21_X1  g0805(.A(new_n769), .B1(new_n1004), .B2(new_n1005), .ZN(new_n1006));
  AOI211_X1 g0806(.A(KEYINPUT106), .B(new_n977), .C1(new_n1003), .C2(new_n765), .ZN(new_n1007));
  OAI21_X1  g0807(.A(new_n976), .B1(new_n1006), .B2(new_n1007), .ZN(new_n1008));
  NOR2_X1   g0808(.A1(new_n808), .A2(new_n284), .ZN(new_n1009));
  AOI211_X1 g0809(.A(new_n390), .B(new_n1009), .C1(G50), .C2(new_n802), .ZN(new_n1010));
  AOI22_X1  g0810(.A1(new_n804), .A2(G58), .B1(new_n852), .B2(G77), .ZN(new_n1011));
  AOI22_X1  g0811(.A1(new_n812), .A2(G159), .B1(new_n815), .B2(G137), .ZN(new_n1012));
  AOI22_X1  g0812(.A1(G143), .A2(new_n806), .B1(new_n799), .B2(G150), .ZN(new_n1013));
  NAND4_X1  g0813(.A1(new_n1010), .A2(new_n1011), .A3(new_n1012), .A4(new_n1013), .ZN(new_n1014));
  INV_X1    g0814(.A(G311), .ZN(new_n1015));
  OAI221_X1 g0815(.A(new_n390), .B1(new_n604), .B2(new_n811), .C1(new_n856), .C2(new_n1015), .ZN(new_n1016));
  NOR2_X1   g0816(.A1(new_n794), .A2(new_n223), .ZN(new_n1017));
  INV_X1    g0817(.A(G317), .ZN(new_n1018));
  OAI22_X1  g0818(.A1(new_n801), .A2(new_n795), .B1(new_n814), .B2(new_n1018), .ZN(new_n1019));
  NOR3_X1   g0819(.A1(new_n1016), .A2(new_n1017), .A3(new_n1019), .ZN(new_n1020));
  NAND3_X1  g0820(.A1(new_n804), .A2(KEYINPUT46), .A3(G116), .ZN(new_n1021));
  AOI22_X1  g0821(.A1(new_n799), .A2(G303), .B1(G107), .B2(new_n809), .ZN(new_n1022));
  NAND3_X1  g0822(.A1(new_n1020), .A2(new_n1021), .A3(new_n1022), .ZN(new_n1023));
  AOI21_X1  g0823(.A(KEYINPUT46), .B1(new_n804), .B2(G116), .ZN(new_n1024));
  XOR2_X1   g0824(.A(new_n1024), .B(KEYINPUT107), .Z(new_n1025));
  OAI21_X1  g0825(.A(new_n1014), .B1(new_n1023), .B2(new_n1025), .ZN(new_n1026));
  XNOR2_X1  g0826(.A(new_n1026), .B(KEYINPUT47), .ZN(new_n1027));
  NAND2_X1  g0827(.A1(new_n1027), .A2(new_n788), .ZN(new_n1028));
  NAND2_X1  g0828(.A1(new_n236), .A2(new_n783), .ZN(new_n1029));
  AOI21_X1  g0829(.A(new_n790), .B1(new_n210), .B2(new_n319), .ZN(new_n1030));
  AOI21_X1  g0830(.A(new_n847), .B1(new_n1029), .B2(new_n1030), .ZN(new_n1031));
  OAI211_X1 g0831(.A(new_n1028), .B(new_n1031), .C1(new_n961), .C2(new_n778), .ZN(new_n1032));
  NAND2_X1  g0832(.A1(new_n1008), .A2(new_n1032), .ZN(G387));
  INV_X1    g0833(.A(new_n765), .ZN(new_n1034));
  INV_X1    g0834(.A(new_n982), .ZN(new_n1035));
  NAND2_X1  g0835(.A1(new_n1034), .A2(new_n1035), .ZN(new_n1036));
  NAND2_X1  g0836(.A1(new_n765), .A2(new_n982), .ZN(new_n1037));
  XNOR2_X1  g0837(.A(new_n717), .B(KEYINPUT108), .ZN(new_n1038));
  NAND3_X1  g0838(.A1(new_n1036), .A2(new_n1037), .A3(new_n1038), .ZN(new_n1039));
  AOI211_X1 g0839(.A(new_n390), .B(new_n1017), .C1(G50), .C2(new_n799), .ZN(new_n1040));
  INV_X1    g0840(.A(new_n277), .ZN(new_n1041));
  AOI22_X1  g0841(.A1(new_n812), .A2(new_n1041), .B1(new_n815), .B2(G150), .ZN(new_n1042));
  AOI22_X1  g0842(.A1(G68), .A2(new_n802), .B1(new_n804), .B2(G77), .ZN(new_n1043));
  AOI22_X1  g0843(.A1(new_n806), .A2(G159), .B1(new_n319), .B2(new_n809), .ZN(new_n1044));
  NAND4_X1  g0844(.A1(new_n1040), .A2(new_n1042), .A3(new_n1043), .A4(new_n1044), .ZN(new_n1045));
  AOI21_X1  g0845(.A(new_n249), .B1(new_n815), .B2(G326), .ZN(new_n1046));
  OAI22_X1  g0846(.A1(new_n803), .A2(new_n604), .B1(new_n808), .B2(new_n795), .ZN(new_n1047));
  AOI22_X1  g0847(.A1(G303), .A2(new_n802), .B1(new_n812), .B2(G311), .ZN(new_n1048));
  INV_X1    g0848(.A(G322), .ZN(new_n1049));
  OAI221_X1 g0849(.A(new_n1048), .B1(new_n1018), .B2(new_n855), .C1(new_n1049), .C2(new_n856), .ZN(new_n1050));
  INV_X1    g0850(.A(KEYINPUT48), .ZN(new_n1051));
  AOI21_X1  g0851(.A(new_n1047), .B1(new_n1050), .B2(new_n1051), .ZN(new_n1052));
  OAI21_X1  g0852(.A(new_n1052), .B1(new_n1051), .B2(new_n1050), .ZN(new_n1053));
  INV_X1    g0853(.A(KEYINPUT49), .ZN(new_n1054));
  OAI221_X1 g0854(.A(new_n1046), .B1(new_n626), .B2(new_n794), .C1(new_n1053), .C2(new_n1054), .ZN(new_n1055));
  AND2_X1   g0855(.A1(new_n1053), .A2(new_n1054), .ZN(new_n1056));
  OAI21_X1  g0856(.A(new_n1045), .B1(new_n1055), .B2(new_n1056), .ZN(new_n1057));
  NAND2_X1  g0857(.A1(new_n1057), .A2(new_n788), .ZN(new_n1058));
  INV_X1    g0858(.A(new_n719), .ZN(new_n1059));
  AOI22_X1  g0859(.A1(new_n780), .A2(new_n1059), .B1(new_n496), .B2(new_n210), .ZN(new_n1060));
  NOR2_X1   g0860(.A1(new_n240), .A2(new_n260), .ZN(new_n1061));
  NAND2_X1  g0861(.A1(new_n1041), .A2(new_n274), .ZN(new_n1062));
  XNOR2_X1  g0862(.A(new_n1062), .B(KEYINPUT50), .ZN(new_n1063));
  OAI211_X1 g0863(.A(new_n719), .B(new_n260), .C1(new_n284), .C2(new_n253), .ZN(new_n1064));
  OAI21_X1  g0864(.A(new_n783), .B1(new_n1063), .B2(new_n1064), .ZN(new_n1065));
  OAI21_X1  g0865(.A(new_n1060), .B1(new_n1061), .B2(new_n1065), .ZN(new_n1066));
  AOI21_X1  g0866(.A(new_n847), .B1(new_n1066), .B2(new_n789), .ZN(new_n1067));
  OAI211_X1 g0867(.A(new_n1058), .B(new_n1067), .C1(new_n706), .C2(new_n778), .ZN(new_n1068));
  OAI211_X1 g0868(.A(new_n1039), .B(new_n1068), .C1(new_n769), .C2(new_n1035), .ZN(G393));
  INV_X1    g0869(.A(new_n999), .ZN(new_n1070));
  NAND3_X1  g0870(.A1(new_n1070), .A2(KEYINPUT109), .A3(new_n708), .ZN(new_n1071));
  NAND2_X1  g0871(.A1(new_n708), .A2(KEYINPUT109), .ZN(new_n1072));
  OR2_X1    g0872(.A1(new_n708), .A2(KEYINPUT109), .ZN(new_n1073));
  NAND3_X1  g0873(.A1(new_n999), .A2(new_n1072), .A3(new_n1073), .ZN(new_n1074));
  NAND2_X1  g0874(.A1(new_n1071), .A2(new_n1074), .ZN(new_n1075));
  OAI211_X1 g0875(.A(new_n1003), .B(new_n1038), .C1(new_n983), .C2(new_n1075), .ZN(new_n1076));
  NAND2_X1  g0876(.A1(new_n1075), .A2(new_n770), .ZN(new_n1077));
  OAI221_X1 g0877(.A(new_n789), .B1(new_n223), .B2(new_n209), .C1(new_n784), .C2(new_n247), .ZN(new_n1078));
  NAND2_X1  g0878(.A1(new_n1078), .A2(new_n771), .ZN(new_n1079));
  AOI22_X1  g0879(.A1(G311), .A2(new_n799), .B1(new_n806), .B2(G317), .ZN(new_n1080));
  XNOR2_X1  g0880(.A(new_n1080), .B(KEYINPUT52), .ZN(new_n1081));
  OAI22_X1  g0881(.A1(new_n811), .A2(new_n857), .B1(new_n808), .B2(new_n626), .ZN(new_n1082));
  NOR2_X1   g0882(.A1(new_n1082), .A2(KEYINPUT110), .ZN(new_n1083));
  OAI22_X1  g0883(.A1(new_n801), .A2(new_n604), .B1(new_n814), .B2(new_n1049), .ZN(new_n1084));
  AOI21_X1  g0884(.A(new_n1084), .B1(G283), .B2(new_n804), .ZN(new_n1085));
  NAND2_X1  g0885(.A1(new_n1082), .A2(KEYINPUT110), .ZN(new_n1086));
  AOI21_X1  g0886(.A(new_n249), .B1(new_n852), .B2(G107), .ZN(new_n1087));
  NAND3_X1  g0887(.A1(new_n1085), .A2(new_n1086), .A3(new_n1087), .ZN(new_n1088));
  NOR3_X1   g0888(.A1(new_n1081), .A2(new_n1083), .A3(new_n1088), .ZN(new_n1089));
  OR2_X1    g0889(.A1(new_n1089), .A2(KEYINPUT111), .ZN(new_n1090));
  NAND2_X1  g0890(.A1(new_n1089), .A2(KEYINPUT111), .ZN(new_n1091));
  AOI22_X1  g0891(.A1(G150), .A2(new_n806), .B1(new_n799), .B2(G159), .ZN(new_n1092));
  XOR2_X1   g0892(.A(new_n1092), .B(KEYINPUT51), .Z(new_n1093));
  AOI22_X1  g0893(.A1(G50), .A2(new_n812), .B1(new_n804), .B2(G68), .ZN(new_n1094));
  AOI22_X1  g0894(.A1(new_n802), .A2(new_n1041), .B1(new_n815), .B2(G143), .ZN(new_n1095));
  NOR2_X1   g0895(.A1(new_n808), .A2(new_n253), .ZN(new_n1096));
  AOI211_X1 g0896(.A(new_n390), .B(new_n1096), .C1(G87), .C2(new_n852), .ZN(new_n1097));
  NAND4_X1  g0897(.A1(new_n1093), .A2(new_n1094), .A3(new_n1095), .A4(new_n1097), .ZN(new_n1098));
  NAND3_X1  g0898(.A1(new_n1090), .A2(new_n1091), .A3(new_n1098), .ZN(new_n1099));
  AOI21_X1  g0899(.A(new_n1079), .B1(new_n1099), .B2(new_n788), .ZN(new_n1100));
  OAI21_X1  g0900(.A(new_n1100), .B1(new_n949), .B2(new_n778), .ZN(new_n1101));
  NAND3_X1  g0901(.A1(new_n1076), .A2(new_n1077), .A3(new_n1101), .ZN(G390));
  XNOR2_X1  g0902(.A(new_n929), .B(KEYINPUT99), .ZN(new_n1103));
  NAND2_X1  g0903(.A1(new_n936), .A2(new_n937), .ZN(new_n1104));
  AOI21_X1  g0904(.A(new_n1103), .B1(new_n1104), .B2(new_n913), .ZN(new_n1105));
  NOR2_X1   g0905(.A1(new_n926), .A2(new_n927), .ZN(new_n1106));
  INV_X1    g0906(.A(new_n761), .ZN(new_n1107));
  AOI22_X1  g0907(.A1(new_n1107), .A2(KEYINPUT26), .B1(new_n680), .B2(new_n681), .ZN(new_n1108));
  OAI211_X1 g0908(.A(new_n695), .B(new_n839), .C1(new_n934), .C2(new_n1108), .ZN(new_n1109));
  AOI21_X1  g0909(.A(new_n933), .B1(new_n1109), .B2(new_n937), .ZN(new_n1110));
  NAND2_X1  g0910(.A1(new_n905), .A2(new_n906), .ZN(new_n1111));
  NAND2_X1  g0911(.A1(new_n931), .A2(new_n1111), .ZN(new_n1112));
  OAI22_X1  g0912(.A1(new_n1105), .A2(new_n1106), .B1(new_n1110), .B2(new_n1112), .ZN(new_n1113));
  NAND4_X1  g0913(.A1(new_n753), .A2(G330), .A3(new_n839), .A4(new_n913), .ZN(new_n1114));
  INV_X1    g0914(.A(KEYINPUT112), .ZN(new_n1115));
  XNOR2_X1  g0915(.A(new_n1114), .B(new_n1115), .ZN(new_n1116));
  OAI21_X1  g0916(.A(KEYINPUT113), .B1(new_n1113), .B2(new_n1116), .ZN(new_n1117));
  XNOR2_X1  g0917(.A(new_n1114), .B(KEYINPUT112), .ZN(new_n1118));
  OR2_X1    g0918(.A1(new_n1110), .A2(new_n1112), .ZN(new_n1119));
  OAI21_X1  g0919(.A(new_n928), .B1(new_n938), .B2(new_n1103), .ZN(new_n1120));
  INV_X1    g0920(.A(KEYINPUT113), .ZN(new_n1121));
  NAND4_X1  g0921(.A1(new_n1118), .A2(new_n1119), .A3(new_n1120), .A4(new_n1121), .ZN(new_n1122));
  NAND2_X1  g0922(.A1(new_n834), .A2(new_n838), .ZN(new_n1123));
  NOR2_X1   g0923(.A1(new_n734), .A2(new_n742), .ZN(new_n1124));
  AOI21_X1  g0924(.A(new_n1123), .B1(new_n1124), .B2(new_n752), .ZN(new_n1125));
  NAND3_X1  g0925(.A1(new_n1125), .A2(G330), .A3(new_n913), .ZN(new_n1126));
  INV_X1    g0926(.A(new_n1126), .ZN(new_n1127));
  NAND2_X1  g0927(.A1(new_n1113), .A2(new_n1127), .ZN(new_n1128));
  NAND4_X1  g0928(.A1(new_n1117), .A2(new_n1122), .A3(new_n770), .A4(new_n1128), .ZN(new_n1129));
  AOI21_X1  g0929(.A(new_n847), .B1(new_n850), .B2(new_n277), .ZN(new_n1130));
  NOR2_X1   g0930(.A1(new_n856), .A2(new_n795), .ZN(new_n1131));
  AOI211_X1 g0931(.A(new_n1096), .B(new_n1131), .C1(G116), .C2(new_n799), .ZN(new_n1132));
  OAI22_X1  g0932(.A1(new_n801), .A2(new_n223), .B1(new_n811), .B2(new_n496), .ZN(new_n1133));
  OR2_X1    g0933(.A1(new_n1133), .A2(KEYINPUT114), .ZN(new_n1134));
  NAND2_X1  g0934(.A1(new_n1133), .A2(KEYINPUT114), .ZN(new_n1135));
  OAI22_X1  g0935(.A1(new_n794), .A2(new_n284), .B1(new_n814), .B2(new_n604), .ZN(new_n1136));
  AOI211_X1 g0936(.A(new_n249), .B(new_n1136), .C1(G87), .C2(new_n804), .ZN(new_n1137));
  NAND4_X1  g0937(.A1(new_n1132), .A2(new_n1134), .A3(new_n1135), .A4(new_n1137), .ZN(new_n1138));
  NOR2_X1   g0938(.A1(new_n803), .A2(new_n279), .ZN(new_n1139));
  XNOR2_X1  g0939(.A(new_n1139), .B(KEYINPUT53), .ZN(new_n1140));
  OAI21_X1  g0940(.A(new_n249), .B1(new_n794), .B2(new_n274), .ZN(new_n1141));
  AOI21_X1  g0941(.A(new_n1141), .B1(G128), .B2(new_n806), .ZN(new_n1142));
  AOI22_X1  g0942(.A1(new_n799), .A2(G132), .B1(G159), .B2(new_n809), .ZN(new_n1143));
  INV_X1    g0943(.A(G125), .ZN(new_n1144));
  OAI22_X1  g0944(.A1(new_n811), .A2(new_n864), .B1(new_n814), .B2(new_n1144), .ZN(new_n1145));
  XNOR2_X1  g0945(.A(KEYINPUT54), .B(G143), .ZN(new_n1146));
  INV_X1    g0946(.A(new_n1146), .ZN(new_n1147));
  AOI21_X1  g0947(.A(new_n1145), .B1(new_n802), .B2(new_n1147), .ZN(new_n1148));
  NAND4_X1  g0948(.A1(new_n1140), .A2(new_n1142), .A3(new_n1143), .A4(new_n1148), .ZN(new_n1149));
  AND2_X1   g0949(.A1(new_n1138), .A2(new_n1149), .ZN(new_n1150));
  OAI221_X1 g0950(.A(new_n1130), .B1(new_n873), .B2(new_n1150), .C1(new_n1106), .C2(new_n776), .ZN(new_n1151));
  NAND2_X1  g0951(.A1(new_n1129), .A2(new_n1151), .ZN(new_n1152));
  NOR2_X1   g0952(.A1(new_n921), .A2(new_n923), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n442), .A2(new_n1153), .ZN(new_n1154));
  NAND3_X1  g0954(.A1(new_n941), .A2(new_n668), .A3(new_n1154), .ZN(new_n1155));
  NAND2_X1  g0955(.A1(new_n1109), .A2(new_n937), .ZN(new_n1156));
  AOI21_X1  g0956(.A(new_n913), .B1(new_n1125), .B2(G330), .ZN(new_n1157));
  NOR2_X1   g0957(.A1(new_n1156), .A2(new_n1157), .ZN(new_n1158));
  AND2_X1   g0958(.A1(new_n1114), .A2(KEYINPUT112), .ZN(new_n1159));
  NOR2_X1   g0959(.A1(new_n1114), .A2(KEYINPUT112), .ZN(new_n1160));
  OAI21_X1  g0960(.A(new_n1158), .B1(new_n1159), .B2(new_n1160), .ZN(new_n1161));
  NAND3_X1  g0961(.A1(new_n753), .A2(G330), .A3(new_n839), .ZN(new_n1162));
  AND2_X1   g0962(.A1(new_n1162), .A2(new_n933), .ZN(new_n1163));
  OAI21_X1  g0963(.A(new_n1104), .B1(new_n1163), .B2(new_n1127), .ZN(new_n1164));
  AOI21_X1  g0964(.A(new_n1155), .B1(new_n1161), .B2(new_n1164), .ZN(new_n1165));
  NAND4_X1  g0965(.A1(new_n1165), .A2(new_n1117), .A3(new_n1122), .A4(new_n1128), .ZN(new_n1166));
  AND2_X1   g0966(.A1(new_n1166), .A2(new_n1038), .ZN(new_n1167));
  NAND3_X1  g0967(.A1(new_n1117), .A2(new_n1122), .A3(new_n1128), .ZN(new_n1168));
  INV_X1    g0968(.A(new_n1165), .ZN(new_n1169));
  NAND2_X1  g0969(.A1(new_n1168), .A2(new_n1169), .ZN(new_n1170));
  AOI21_X1  g0970(.A(new_n1152), .B1(new_n1167), .B2(new_n1170), .ZN(new_n1171));
  INV_X1    g0971(.A(new_n1171), .ZN(G378));
  INV_X1    g0972(.A(new_n1038), .ZN(new_n1173));
  INV_X1    g0973(.A(KEYINPUT120), .ZN(new_n1174));
  NOR4_X1   g0974(.A1(new_n613), .A2(new_n652), .A3(new_n492), .A4(new_n696), .ZN(new_n1175));
  NAND2_X1  g0975(.A1(new_n746), .A2(new_n733), .ZN(new_n1176));
  OAI211_X1 g0976(.A(new_n913), .B(new_n839), .C1(new_n1175), .C2(new_n1176), .ZN(new_n1177));
  OAI21_X1  g0977(.A(KEYINPUT40), .B1(new_n894), .B2(new_n895), .ZN(new_n1178));
  OAI21_X1  g0978(.A(G330), .B1(new_n1177), .B2(new_n1178), .ZN(new_n1179));
  OAI21_X1  g0979(.A(new_n1174), .B1(new_n915), .B2(new_n1179), .ZN(new_n1180));
  AOI21_X1  g0980(.A(new_n923), .B1(new_n914), .B2(new_n918), .ZN(new_n1181));
  AOI21_X1  g0981(.A(new_n1177), .B1(new_n896), .B2(new_n907), .ZN(new_n1182));
  OAI211_X1 g0982(.A(new_n1181), .B(KEYINPUT120), .C1(KEYINPUT40), .C2(new_n1182), .ZN(new_n1183));
  NAND2_X1  g0983(.A1(new_n296), .A2(new_n329), .ZN(new_n1184));
  AND2_X1   g0984(.A1(new_n288), .A2(new_n694), .ZN(new_n1185));
  AND2_X1   g0985(.A1(new_n1184), .A2(new_n1185), .ZN(new_n1186));
  NOR2_X1   g0986(.A1(new_n1184), .A2(new_n1185), .ZN(new_n1187));
  XNOR2_X1  g0987(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1188));
  INV_X1    g0988(.A(new_n1188), .ZN(new_n1189));
  OR3_X1    g0989(.A1(new_n1186), .A2(new_n1187), .A3(new_n1189), .ZN(new_n1190));
  OAI21_X1  g0990(.A(new_n1189), .B1(new_n1186), .B2(new_n1187), .ZN(new_n1191));
  NAND2_X1  g0991(.A1(new_n1190), .A2(new_n1191), .ZN(new_n1192));
  INV_X1    g0992(.A(new_n1192), .ZN(new_n1193));
  NAND3_X1  g0993(.A1(new_n1180), .A2(new_n1183), .A3(new_n1193), .ZN(new_n1194));
  OAI211_X1 g0994(.A(new_n1174), .B(new_n1192), .C1(new_n915), .C2(new_n1179), .ZN(new_n1195));
  AND3_X1   g0995(.A1(new_n1194), .A2(new_n940), .A3(new_n1195), .ZN(new_n1196));
  AOI21_X1  g0996(.A(new_n940), .B1(new_n1194), .B2(new_n1195), .ZN(new_n1197));
  NOR2_X1   g0997(.A1(new_n1196), .A2(new_n1197), .ZN(new_n1198));
  INV_X1    g0998(.A(new_n1155), .ZN(new_n1199));
  NAND2_X1  g0999(.A1(new_n1166), .A2(new_n1199), .ZN(new_n1200));
  NAND2_X1  g1000(.A1(new_n1198), .A2(new_n1200), .ZN(new_n1201));
  INV_X1    g1001(.A(KEYINPUT57), .ZN(new_n1202));
  AOI21_X1  g1002(.A(new_n1173), .B1(new_n1201), .B2(new_n1202), .ZN(new_n1203));
  AND2_X1   g1003(.A1(new_n1166), .A2(new_n1199), .ZN(new_n1204));
  NAND2_X1  g1004(.A1(new_n1194), .A2(new_n1195), .ZN(new_n1205));
  INV_X1    g1005(.A(new_n940), .ZN(new_n1206));
  NAND2_X1  g1006(.A1(new_n1205), .A2(new_n1206), .ZN(new_n1207));
  NAND3_X1  g1007(.A1(new_n1194), .A2(new_n940), .A3(new_n1195), .ZN(new_n1208));
  NAND3_X1  g1008(.A1(new_n1207), .A2(KEYINPUT57), .A3(new_n1208), .ZN(new_n1209));
  NOR3_X1   g1009(.A1(new_n1204), .A2(new_n1209), .A3(KEYINPUT121), .ZN(new_n1210));
  INV_X1    g1010(.A(KEYINPUT121), .ZN(new_n1211));
  NOR3_X1   g1011(.A1(new_n1196), .A2(new_n1197), .A3(new_n1202), .ZN(new_n1212));
  AOI21_X1  g1012(.A(new_n1211), .B1(new_n1212), .B2(new_n1200), .ZN(new_n1213));
  OAI21_X1  g1013(.A(new_n1203), .B1(new_n1210), .B2(new_n1213), .ZN(new_n1214));
  NOR3_X1   g1014(.A1(new_n1196), .A2(new_n1197), .A3(new_n769), .ZN(new_n1215));
  AOI21_X1  g1015(.A(new_n847), .B1(new_n274), .B2(new_n848), .ZN(new_n1216));
  XNOR2_X1  g1016(.A(new_n1216), .B(KEYINPUT118), .ZN(new_n1217));
  AOI22_X1  g1017(.A1(new_n806), .A2(G125), .B1(G150), .B2(new_n809), .ZN(new_n1218));
  XOR2_X1   g1018(.A(new_n1218), .B(KEYINPUT116), .Z(new_n1219));
  AOI22_X1  g1019(.A1(G137), .A2(new_n802), .B1(new_n812), .B2(G132), .ZN(new_n1220));
  OAI21_X1  g1020(.A(new_n1220), .B1(new_n803), .B2(new_n1146), .ZN(new_n1221));
  AOI21_X1  g1021(.A(new_n1221), .B1(G128), .B2(new_n799), .ZN(new_n1222));
  NAND2_X1  g1022(.A1(new_n1219), .A2(new_n1222), .ZN(new_n1223));
  OR2_X1    g1023(.A1(new_n1223), .A2(KEYINPUT59), .ZN(new_n1224));
  NAND2_X1  g1024(.A1(new_n1223), .A2(KEYINPUT59), .ZN(new_n1225));
  NOR2_X1   g1025(.A1(new_n794), .A2(new_n821), .ZN(new_n1226));
  NAND2_X1  g1026(.A1(new_n603), .A2(new_n259), .ZN(new_n1227));
  XNOR2_X1  g1027(.A(new_n1227), .B(KEYINPUT115), .ZN(new_n1228));
  XNOR2_X1  g1028(.A(KEYINPUT117), .B(G124), .ZN(new_n1229));
  AOI211_X1 g1029(.A(new_n1226), .B(new_n1228), .C1(new_n815), .C2(new_n1229), .ZN(new_n1230));
  NAND3_X1  g1030(.A1(new_n1224), .A2(new_n1225), .A3(new_n1230), .ZN(new_n1231));
  NOR2_X1   g1031(.A1(new_n249), .A2(G41), .ZN(new_n1232));
  INV_X1    g1032(.A(new_n1232), .ZN(new_n1233));
  AOI211_X1 g1033(.A(new_n1009), .B(new_n1233), .C1(G77), .C2(new_n804), .ZN(new_n1234));
  OAI221_X1 g1034(.A(new_n1234), .B1(new_n496), .B2(new_n855), .C1(new_n626), .C2(new_n856), .ZN(new_n1235));
  OAI22_X1  g1035(.A1(new_n811), .A2(new_n223), .B1(new_n814), .B2(new_n795), .ZN(new_n1236));
  OAI22_X1  g1036(.A1(new_n320), .A2(new_n801), .B1(new_n221), .B2(new_n794), .ZN(new_n1237));
  NOR3_X1   g1037(.A1(new_n1235), .A2(new_n1236), .A3(new_n1237), .ZN(new_n1238));
  OR2_X1    g1038(.A1(new_n1238), .A2(KEYINPUT58), .ZN(new_n1239));
  NAND2_X1  g1039(.A1(new_n1238), .A2(KEYINPUT58), .ZN(new_n1240));
  NAND3_X1  g1040(.A1(new_n1233), .A2(new_n274), .A3(new_n1228), .ZN(new_n1241));
  AND4_X1   g1041(.A1(new_n1231), .A2(new_n1239), .A3(new_n1240), .A4(new_n1241), .ZN(new_n1242));
  OAI221_X1 g1042(.A(new_n1217), .B1(new_n873), .B2(new_n1242), .C1(new_n1192), .C2(new_n776), .ZN(new_n1243));
  XNOR2_X1  g1043(.A(new_n1243), .B(KEYINPUT119), .ZN(new_n1244));
  NOR2_X1   g1044(.A1(new_n1215), .A2(new_n1244), .ZN(new_n1245));
  NAND2_X1  g1045(.A1(new_n1214), .A2(new_n1245), .ZN(G375));
  NAND2_X1  g1046(.A1(new_n1161), .A2(new_n1164), .ZN(new_n1247));
  NAND2_X1  g1047(.A1(new_n1247), .A2(new_n770), .ZN(new_n1248));
  AOI21_X1  g1048(.A(new_n847), .B1(new_n850), .B2(new_n284), .ZN(new_n1249));
  OAI22_X1  g1049(.A1(new_n801), .A2(new_n496), .B1(new_n811), .B2(new_n626), .ZN(new_n1250));
  XNOR2_X1  g1050(.A(new_n1250), .B(KEYINPUT123), .ZN(new_n1251));
  AOI22_X1  g1051(.A1(new_n804), .A2(G97), .B1(new_n815), .B2(G303), .ZN(new_n1252));
  OAI211_X1 g1052(.A(new_n1252), .B(new_n390), .C1(new_n253), .C2(new_n794), .ZN(new_n1253));
  AOI22_X1  g1053(.A1(new_n799), .A2(G283), .B1(new_n319), .B2(new_n809), .ZN(new_n1254));
  OAI21_X1  g1054(.A(new_n1254), .B1(new_n604), .B2(new_n856), .ZN(new_n1255));
  NOR3_X1   g1055(.A1(new_n1251), .A2(new_n1253), .A3(new_n1255), .ZN(new_n1256));
  OR2_X1    g1056(.A1(new_n1256), .A2(KEYINPUT124), .ZN(new_n1257));
  NAND2_X1  g1057(.A1(new_n1256), .A2(KEYINPUT124), .ZN(new_n1258));
  OAI21_X1  g1058(.A(new_n249), .B1(new_n794), .B2(new_n221), .ZN(new_n1259));
  AOI21_X1  g1059(.A(new_n1259), .B1(G137), .B2(new_n799), .ZN(new_n1260));
  AOI22_X1  g1060(.A1(G150), .A2(new_n802), .B1(new_n812), .B2(new_n1147), .ZN(new_n1261));
  AOI22_X1  g1061(.A1(new_n806), .A2(G132), .B1(G50), .B2(new_n809), .ZN(new_n1262));
  AOI22_X1  g1062(.A1(new_n804), .A2(G159), .B1(new_n815), .B2(G128), .ZN(new_n1263));
  NAND4_X1  g1063(.A1(new_n1260), .A2(new_n1261), .A3(new_n1262), .A4(new_n1263), .ZN(new_n1264));
  AND3_X1   g1064(.A1(new_n1257), .A2(new_n1258), .A3(new_n1264), .ZN(new_n1265));
  OAI221_X1 g1065(.A(new_n1249), .B1(new_n873), .B2(new_n1265), .C1(new_n913), .C2(new_n776), .ZN(new_n1266));
  NAND2_X1  g1066(.A1(new_n1248), .A2(new_n1266), .ZN(new_n1267));
  INV_X1    g1067(.A(new_n1267), .ZN(new_n1268));
  NAND3_X1  g1068(.A1(new_n1161), .A2(new_n1155), .A3(new_n1164), .ZN(new_n1269));
  XOR2_X1   g1069(.A(new_n977), .B(KEYINPUT122), .Z(new_n1270));
  INV_X1    g1070(.A(new_n1270), .ZN(new_n1271));
  NAND3_X1  g1071(.A1(new_n1169), .A2(new_n1269), .A3(new_n1271), .ZN(new_n1272));
  NAND2_X1  g1072(.A1(new_n1268), .A2(new_n1272), .ZN(G381));
  INV_X1    g1073(.A(G375), .ZN(new_n1274));
  INV_X1    g1074(.A(G390), .ZN(new_n1275));
  AND3_X1   g1075(.A1(new_n1008), .A2(new_n1032), .A3(new_n1275), .ZN(new_n1276));
  NOR4_X1   g1076(.A1(G384), .A2(G381), .A3(G396), .A4(G393), .ZN(new_n1277));
  NAND4_X1  g1077(.A1(new_n1274), .A2(new_n1171), .A3(new_n1276), .A4(new_n1277), .ZN(G407));
  INV_X1    g1078(.A(G213), .ZN(new_n1279));
  NOR2_X1   g1079(.A1(new_n1279), .A2(G343), .ZN(new_n1280));
  NAND3_X1  g1080(.A1(new_n1274), .A2(new_n1171), .A3(new_n1280), .ZN(new_n1281));
  NAND3_X1  g1081(.A1(G407), .A2(new_n1281), .A3(G213), .ZN(G409));
  INV_X1    g1082(.A(KEYINPUT61), .ZN(new_n1283));
  NAND3_X1  g1083(.A1(new_n1214), .A2(G378), .A3(new_n1245), .ZN(new_n1284));
  NAND3_X1  g1084(.A1(new_n1198), .A2(new_n1200), .A3(new_n1271), .ZN(new_n1285));
  AND2_X1   g1085(.A1(new_n1285), .A2(new_n1243), .ZN(new_n1286));
  NAND2_X1  g1086(.A1(new_n1198), .A2(KEYINPUT125), .ZN(new_n1287));
  INV_X1    g1087(.A(KEYINPUT125), .ZN(new_n1288));
  OAI21_X1  g1088(.A(new_n1288), .B1(new_n1196), .B2(new_n1197), .ZN(new_n1289));
  NAND3_X1  g1089(.A1(new_n1287), .A2(new_n770), .A3(new_n1289), .ZN(new_n1290));
  NAND2_X1  g1090(.A1(new_n1286), .A2(new_n1290), .ZN(new_n1291));
  NAND2_X1  g1091(.A1(new_n1291), .A2(new_n1171), .ZN(new_n1292));
  AOI21_X1  g1092(.A(new_n1280), .B1(new_n1284), .B2(new_n1292), .ZN(new_n1293));
  NAND2_X1  g1093(.A1(new_n1280), .A2(G2897), .ZN(new_n1294));
  INV_X1    g1094(.A(G384), .ZN(new_n1295));
  OR2_X1    g1095(.A1(new_n1269), .A2(KEYINPUT60), .ZN(new_n1296));
  NAND2_X1  g1096(.A1(new_n1269), .A2(KEYINPUT60), .ZN(new_n1297));
  AOI211_X1 g1097(.A(new_n1173), .B(new_n1165), .C1(new_n1296), .C2(new_n1297), .ZN(new_n1298));
  OAI21_X1  g1098(.A(new_n1295), .B1(new_n1298), .B2(new_n1267), .ZN(new_n1299));
  NAND2_X1  g1099(.A1(new_n1296), .A2(new_n1297), .ZN(new_n1300));
  NAND3_X1  g1100(.A1(new_n1300), .A2(new_n1038), .A3(new_n1169), .ZN(new_n1301));
  NAND3_X1  g1101(.A1(new_n1301), .A2(G384), .A3(new_n1268), .ZN(new_n1302));
  AOI21_X1  g1102(.A(new_n1294), .B1(new_n1299), .B2(new_n1302), .ZN(new_n1303));
  INV_X1    g1103(.A(new_n1303), .ZN(new_n1304));
  NAND3_X1  g1104(.A1(new_n1299), .A2(new_n1302), .A3(new_n1294), .ZN(new_n1305));
  NAND2_X1  g1105(.A1(new_n1304), .A2(new_n1305), .ZN(new_n1306));
  OAI21_X1  g1106(.A(new_n1283), .B1(new_n1293), .B2(new_n1306), .ZN(new_n1307));
  XNOR2_X1  g1107(.A(G393), .B(new_n830), .ZN(new_n1308));
  INV_X1    g1108(.A(new_n1308), .ZN(new_n1309));
  AOI21_X1  g1109(.A(new_n1275), .B1(new_n1008), .B2(new_n1032), .ZN(new_n1310));
  NOR3_X1   g1110(.A1(new_n1276), .A2(new_n1310), .A3(KEYINPUT127), .ZN(new_n1311));
  INV_X1    g1111(.A(KEYINPUT127), .ZN(new_n1312));
  INV_X1    g1112(.A(new_n975), .ZN(new_n1313));
  NAND2_X1  g1113(.A1(new_n1313), .A2(new_n973), .ZN(new_n1314));
  INV_X1    g1114(.A(new_n977), .ZN(new_n1315));
  INV_X1    g1115(.A(KEYINPUT104), .ZN(new_n1316));
  OAI21_X1  g1116(.A(new_n995), .B1(new_n999), .B2(new_n1316), .ZN(new_n1317));
  NAND2_X1  g1117(.A1(new_n1317), .A2(new_n708), .ZN(new_n1318));
  AOI21_X1  g1118(.A(new_n1037), .B1(new_n1318), .B2(new_n1001), .ZN(new_n1319));
  OAI21_X1  g1119(.A(new_n1315), .B1(new_n1319), .B2(new_n1034), .ZN(new_n1320));
  AOI21_X1  g1120(.A(new_n770), .B1(new_n1320), .B2(KEYINPUT106), .ZN(new_n1321));
  INV_X1    g1121(.A(new_n1007), .ZN(new_n1322));
  AOI21_X1  g1122(.A(new_n1314), .B1(new_n1321), .B2(new_n1322), .ZN(new_n1323));
  INV_X1    g1123(.A(new_n1032), .ZN(new_n1324));
  OAI21_X1  g1124(.A(G390), .B1(new_n1323), .B2(new_n1324), .ZN(new_n1325));
  NAND3_X1  g1125(.A1(new_n1008), .A2(new_n1032), .A3(new_n1275), .ZN(new_n1326));
  AOI21_X1  g1126(.A(new_n1312), .B1(new_n1325), .B2(new_n1326), .ZN(new_n1327));
  OAI21_X1  g1127(.A(new_n1309), .B1(new_n1311), .B2(new_n1327), .ZN(new_n1328));
  OAI21_X1  g1128(.A(KEYINPUT127), .B1(new_n1276), .B2(new_n1310), .ZN(new_n1329));
  NAND3_X1  g1129(.A1(new_n1325), .A2(new_n1312), .A3(new_n1326), .ZN(new_n1330));
  NAND3_X1  g1130(.A1(new_n1329), .A2(new_n1330), .A3(new_n1308), .ZN(new_n1331));
  NAND2_X1  g1131(.A1(new_n1328), .A2(new_n1331), .ZN(new_n1332));
  NOR2_X1   g1132(.A1(new_n1307), .A2(new_n1332), .ZN(new_n1333));
  NAND2_X1  g1133(.A1(new_n1299), .A2(new_n1302), .ZN(new_n1334));
  AOI211_X1 g1134(.A(new_n1280), .B(new_n1334), .C1(new_n1284), .C2(new_n1292), .ZN(new_n1335));
  NAND2_X1  g1135(.A1(new_n1335), .A2(KEYINPUT63), .ZN(new_n1336));
  INV_X1    g1136(.A(KEYINPUT126), .ZN(new_n1337));
  OAI21_X1  g1137(.A(new_n1337), .B1(new_n1335), .B2(KEYINPUT63), .ZN(new_n1338));
  INV_X1    g1138(.A(new_n1280), .ZN(new_n1339));
  INV_X1    g1139(.A(new_n1334), .ZN(new_n1340));
  INV_X1    g1140(.A(new_n1245), .ZN(new_n1341));
  OAI21_X1  g1141(.A(KEYINPUT121), .B1(new_n1204), .B2(new_n1209), .ZN(new_n1342));
  NAND3_X1  g1142(.A1(new_n1212), .A2(new_n1211), .A3(new_n1200), .ZN(new_n1343));
  NAND2_X1  g1143(.A1(new_n1342), .A2(new_n1343), .ZN(new_n1344));
  AOI211_X1 g1144(.A(new_n1171), .B(new_n1341), .C1(new_n1344), .C2(new_n1203), .ZN(new_n1345));
  AOI21_X1  g1145(.A(G378), .B1(new_n1286), .B2(new_n1290), .ZN(new_n1346));
  OAI211_X1 g1146(.A(new_n1339), .B(new_n1340), .C1(new_n1345), .C2(new_n1346), .ZN(new_n1347));
  INV_X1    g1147(.A(KEYINPUT63), .ZN(new_n1348));
  NAND3_X1  g1148(.A1(new_n1347), .A2(KEYINPUT126), .A3(new_n1348), .ZN(new_n1349));
  NAND4_X1  g1149(.A1(new_n1333), .A2(new_n1336), .A3(new_n1338), .A4(new_n1349), .ZN(new_n1350));
  OAI21_X1  g1150(.A(new_n1339), .B1(new_n1345), .B2(new_n1346), .ZN(new_n1351));
  INV_X1    g1151(.A(new_n1305), .ZN(new_n1352));
  NOR2_X1   g1152(.A1(new_n1352), .A2(new_n1303), .ZN(new_n1353));
  AOI21_X1  g1153(.A(KEYINPUT61), .B1(new_n1351), .B2(new_n1353), .ZN(new_n1354));
  INV_X1    g1154(.A(KEYINPUT62), .ZN(new_n1355));
  NAND3_X1  g1155(.A1(new_n1293), .A2(new_n1355), .A3(new_n1340), .ZN(new_n1356));
  NAND2_X1  g1156(.A1(new_n1347), .A2(KEYINPUT62), .ZN(new_n1357));
  NAND3_X1  g1157(.A1(new_n1354), .A2(new_n1356), .A3(new_n1357), .ZN(new_n1358));
  NAND2_X1  g1158(.A1(new_n1358), .A2(new_n1332), .ZN(new_n1359));
  NAND2_X1  g1159(.A1(new_n1350), .A2(new_n1359), .ZN(G405));
  NAND2_X1  g1160(.A1(G375), .A2(new_n1171), .ZN(new_n1361));
  NAND2_X1  g1161(.A1(new_n1361), .A2(new_n1284), .ZN(new_n1362));
  NAND2_X1  g1162(.A1(new_n1362), .A2(new_n1340), .ZN(new_n1363));
  NAND3_X1  g1163(.A1(new_n1361), .A2(new_n1284), .A3(new_n1334), .ZN(new_n1364));
  NAND2_X1  g1164(.A1(new_n1363), .A2(new_n1364), .ZN(new_n1365));
  XNOR2_X1  g1165(.A(new_n1365), .B(new_n1332), .ZN(G402));
endmodule


