//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 1 1 1 1 1 0 1 1 0 1 1 0 0 0 1 1 1 1 1 0 1 1 0 1 1 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 0 0 0 0 1 1 1 0 1 1 0 1 0 1 0 1 1 1 1 0 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:34:59 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n236, new_n237,
    new_n238, new_n240, new_n241, new_n242, new_n243, new_n244, new_n245,
    new_n246, new_n247, new_n248, new_n250, new_n251, new_n252, new_n253,
    new_n254, new_n255, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n692, new_n693, new_n694, new_n695, new_n696,
    new_n697, new_n698, new_n699, new_n700, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n772, new_n773, new_n774, new_n775,
    new_n776, new_n777, new_n778, new_n779, new_n780, new_n781, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1087,
    new_n1088, new_n1089, new_n1090, new_n1091, new_n1092, new_n1093,
    new_n1094, new_n1095, new_n1096, new_n1097, new_n1098, new_n1099,
    new_n1100, new_n1101, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1108, new_n1109, new_n1110, new_n1111, new_n1112,
    new_n1113, new_n1114, new_n1115, new_n1116, new_n1117, new_n1118,
    new_n1119, new_n1120, new_n1121, new_n1122, new_n1123, new_n1124,
    new_n1125, new_n1126, new_n1127, new_n1128, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1186, new_n1187, new_n1188, new_n1189, new_n1190, new_n1191,
    new_n1192, new_n1193, new_n1194, new_n1195, new_n1196, new_n1197,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1251, new_n1252,
    new_n1253, new_n1254, new_n1255, new_n1256, new_n1257, new_n1258,
    new_n1260, new_n1261, new_n1262, new_n1263, new_n1264, new_n1265,
    new_n1266, new_n1267, new_n1268, new_n1269, new_n1270, new_n1271,
    new_n1272, new_n1273, new_n1274, new_n1275, new_n1276, new_n1277,
    new_n1278, new_n1279, new_n1280, new_n1281, new_n1282, new_n1283,
    new_n1284, new_n1285, new_n1286, new_n1287, new_n1289, new_n1290,
    new_n1291, new_n1292, new_n1293, new_n1294, new_n1295, new_n1296,
    new_n1297, new_n1298, new_n1300, new_n1301, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1346,
    new_n1347, new_n1348, new_n1349, new_n1350, new_n1351, new_n1352,
    new_n1353, new_n1354, new_n1355, new_n1356, new_n1357, new_n1358,
    new_n1359, new_n1361, new_n1362, new_n1363, new_n1364, new_n1365,
    new_n1366, new_n1367;
  XNOR2_X1  g0000(.A(KEYINPUT64), .B(G50), .ZN(new_n201));
  NOR2_X1   g0001(.A1(G58), .A2(G68), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0005(.A(G1), .ZN(new_n206));
  INV_X1    g0006(.A(G20), .ZN(new_n207));
  NOR2_X1   g0007(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  NAND2_X1  g0008(.A1(G116), .A2(G270), .ZN(new_n209));
  INV_X1    g0009(.A(G107), .ZN(new_n210));
  INV_X1    g0010(.A(G264), .ZN(new_n211));
  OAI21_X1  g0011(.A(new_n209), .B1(new_n210), .B2(new_n211), .ZN(new_n212));
  AOI22_X1  g0012(.A1(G50), .A2(G226), .B1(G77), .B2(G244), .ZN(new_n213));
  INV_X1    g0013(.A(G87), .ZN(new_n214));
  INV_X1    g0014(.A(G250), .ZN(new_n215));
  INV_X1    g0015(.A(G97), .ZN(new_n216));
  INV_X1    g0016(.A(G257), .ZN(new_n217));
  OAI221_X1 g0017(.A(new_n213), .B1(new_n214), .B2(new_n215), .C1(new_n216), .C2(new_n217), .ZN(new_n218));
  AOI211_X1 g0018(.A(new_n212), .B(new_n218), .C1(G58), .C2(G232), .ZN(new_n219));
  XNOR2_X1  g0019(.A(KEYINPUT66), .B(G68), .ZN(new_n220));
  NAND2_X1  g0020(.A1(new_n220), .A2(G238), .ZN(new_n221));
  AOI21_X1  g0021(.A(new_n208), .B1(new_n219), .B2(new_n221), .ZN(new_n222));
  INV_X1    g0022(.A(KEYINPUT1), .ZN(new_n223));
  NAND2_X1  g0023(.A1(new_n222), .A2(new_n223), .ZN(new_n224));
  XOR2_X1   g0024(.A(new_n224), .B(KEYINPUT67), .Z(new_n225));
  INV_X1    g0025(.A(G13), .ZN(new_n226));
  NAND2_X1  g0026(.A1(new_n208), .A2(new_n226), .ZN(new_n227));
  INV_X1    g0027(.A(new_n227), .ZN(new_n228));
  OAI211_X1 g0028(.A(new_n228), .B(G250), .C1(G257), .C2(G264), .ZN(new_n229));
  XNOR2_X1  g0029(.A(new_n229), .B(KEYINPUT0), .ZN(new_n230));
  NAND2_X1  g0030(.A1(G1), .A2(G13), .ZN(new_n231));
  INV_X1    g0031(.A(new_n231), .ZN(new_n232));
  NAND2_X1  g0032(.A1(new_n232), .A2(G20), .ZN(new_n233));
  INV_X1    g0033(.A(G50), .ZN(new_n234));
  INV_X1    g0034(.A(new_n202), .ZN(new_n235));
  AOI21_X1  g0035(.A(new_n234), .B1(new_n235), .B2(KEYINPUT65), .ZN(new_n236));
  OAI21_X1  g0036(.A(new_n236), .B1(KEYINPUT65), .B2(new_n235), .ZN(new_n237));
  OAI221_X1 g0037(.A(new_n230), .B1(new_n233), .B2(new_n237), .C1(new_n222), .C2(new_n223), .ZN(new_n238));
  NOR2_X1   g0038(.A1(new_n225), .A2(new_n238), .ZN(G361));
  XOR2_X1   g0039(.A(G238), .B(G244), .Z(new_n240));
  XNOR2_X1  g0040(.A(KEYINPUT68), .B(KEYINPUT2), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XNOR2_X1  g0042(.A(G226), .B(G232), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XNOR2_X1  g0044(.A(G250), .B(G257), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n245), .B(KEYINPUT69), .ZN(new_n246));
  XOR2_X1   g0046(.A(G264), .B(G270), .Z(new_n247));
  XNOR2_X1  g0047(.A(new_n246), .B(new_n247), .ZN(new_n248));
  XOR2_X1   g0048(.A(new_n244), .B(new_n248), .Z(G358));
  XOR2_X1   g0049(.A(G87), .B(G97), .Z(new_n250));
  XNOR2_X1  g0050(.A(G107), .B(G116), .ZN(new_n251));
  XNOR2_X1  g0051(.A(new_n250), .B(new_n251), .ZN(new_n252));
  XOR2_X1   g0052(.A(G68), .B(G77), .Z(new_n253));
  XNOR2_X1  g0053(.A(G50), .B(G58), .ZN(new_n254));
  XNOR2_X1  g0054(.A(new_n253), .B(new_n254), .ZN(new_n255));
  XNOR2_X1  g0055(.A(new_n252), .B(new_n255), .ZN(G351));
  NAND2_X1  g0056(.A1(G33), .A2(G41), .ZN(new_n257));
  NAND2_X1  g0057(.A1(new_n232), .A2(new_n257), .ZN(new_n258));
  INV_X1    g0058(.A(G77), .ZN(new_n259));
  INV_X1    g0059(.A(G33), .ZN(new_n260));
  NAND2_X1  g0060(.A1(new_n260), .A2(KEYINPUT3), .ZN(new_n261));
  INV_X1    g0061(.A(KEYINPUT3), .ZN(new_n262));
  NAND2_X1  g0062(.A1(new_n262), .A2(G33), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n261), .A2(new_n263), .ZN(new_n264));
  AOI21_X1  g0064(.A(new_n258), .B1(new_n259), .B2(new_n264), .ZN(new_n265));
  MUX2_X1   g0065(.A(G222), .B(G223), .S(G1698), .Z(new_n266));
  OAI21_X1  g0066(.A(new_n265), .B1(new_n264), .B2(new_n266), .ZN(new_n267));
  INV_X1    g0067(.A(KEYINPUT70), .ZN(new_n268));
  NAND2_X1  g0068(.A1(new_n257), .A2(new_n268), .ZN(new_n269));
  NAND3_X1  g0069(.A1(KEYINPUT70), .A2(G33), .A3(G41), .ZN(new_n270));
  NAND3_X1  g0070(.A1(new_n269), .A2(new_n232), .A3(new_n270), .ZN(new_n271));
  INV_X1    g0071(.A(G41), .ZN(new_n272));
  INV_X1    g0072(.A(G45), .ZN(new_n273));
  AOI21_X1  g0073(.A(G1), .B1(new_n272), .B2(new_n273), .ZN(new_n274));
  NAND3_X1  g0074(.A1(new_n271), .A2(G274), .A3(new_n274), .ZN(new_n275));
  INV_X1    g0075(.A(new_n274), .ZN(new_n276));
  NAND3_X1  g0076(.A1(new_n271), .A2(new_n276), .A3(G226), .ZN(new_n277));
  NAND3_X1  g0077(.A1(new_n267), .A2(new_n275), .A3(new_n277), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n278), .A2(G200), .ZN(new_n279));
  INV_X1    g0079(.A(G190), .ZN(new_n280));
  OAI21_X1  g0080(.A(new_n279), .B1(new_n280), .B2(new_n278), .ZN(new_n281));
  NAND3_X1  g0081(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n282), .A2(new_n231), .ZN(new_n283));
  INV_X1    g0083(.A(new_n283), .ZN(new_n284));
  INV_X1    g0084(.A(KEYINPUT8), .ZN(new_n285));
  NAND2_X1  g0085(.A1(new_n285), .A2(G58), .ZN(new_n286));
  XNOR2_X1  g0086(.A(new_n286), .B(KEYINPUT72), .ZN(new_n287));
  NOR2_X1   g0087(.A1(new_n285), .A2(G58), .ZN(new_n288));
  INV_X1    g0088(.A(new_n288), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n289), .A2(KEYINPUT71), .ZN(new_n290));
  OR3_X1    g0090(.A1(new_n285), .A2(KEYINPUT71), .A3(G58), .ZN(new_n291));
  NAND3_X1  g0091(.A1(new_n287), .A2(new_n290), .A3(new_n291), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n207), .A2(G33), .ZN(new_n293));
  INV_X1    g0093(.A(new_n293), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n292), .A2(new_n294), .ZN(new_n295));
  NOR2_X1   g0095(.A1(G20), .A2(G33), .ZN(new_n296));
  AOI22_X1  g0096(.A1(new_n203), .A2(G20), .B1(G150), .B2(new_n296), .ZN(new_n297));
  AOI21_X1  g0097(.A(new_n284), .B1(new_n295), .B2(new_n297), .ZN(new_n298));
  NAND3_X1  g0098(.A1(new_n206), .A2(G13), .A3(G20), .ZN(new_n299));
  INV_X1    g0099(.A(new_n299), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n300), .A2(new_n234), .ZN(new_n301));
  AOI21_X1  g0101(.A(new_n283), .B1(new_n206), .B2(G20), .ZN(new_n302));
  INV_X1    g0102(.A(new_n302), .ZN(new_n303));
  OAI21_X1  g0103(.A(new_n301), .B1(new_n303), .B2(new_n234), .ZN(new_n304));
  OR2_X1    g0104(.A1(new_n298), .A2(new_n304), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n305), .A2(KEYINPUT9), .ZN(new_n306));
  OR3_X1    g0106(.A1(new_n298), .A2(KEYINPUT9), .A3(new_n304), .ZN(new_n307));
  AOI21_X1  g0107(.A(new_n281), .B1(new_n306), .B2(new_n307), .ZN(new_n308));
  NOR2_X1   g0108(.A1(new_n281), .A2(KEYINPUT75), .ZN(new_n309));
  NOR2_X1   g0109(.A1(new_n309), .A2(KEYINPUT10), .ZN(new_n310));
  XNOR2_X1  g0110(.A(new_n308), .B(new_n310), .ZN(new_n311));
  NAND3_X1  g0111(.A1(new_n271), .A2(new_n276), .A3(G244), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n312), .A2(new_n275), .ZN(new_n313));
  INV_X1    g0113(.A(new_n258), .ZN(new_n314));
  XNOR2_X1  g0114(.A(KEYINPUT3), .B(G33), .ZN(new_n315));
  NAND3_X1  g0115(.A1(new_n315), .A2(G238), .A3(G1698), .ZN(new_n316));
  INV_X1    g0116(.A(G1698), .ZN(new_n317));
  NAND3_X1  g0117(.A1(new_n315), .A2(G232), .A3(new_n317), .ZN(new_n318));
  OAI211_X1 g0118(.A(new_n316), .B(new_n318), .C1(new_n210), .C2(new_n315), .ZN(new_n319));
  AOI21_X1  g0119(.A(new_n313), .B1(new_n314), .B2(new_n319), .ZN(new_n320));
  NOR2_X1   g0120(.A1(new_n320), .A2(G169), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n302), .A2(G77), .ZN(new_n322));
  OAI21_X1  g0122(.A(new_n322), .B1(G77), .B2(new_n299), .ZN(new_n323));
  XOR2_X1   g0123(.A(KEYINPUT15), .B(G87), .Z(new_n324));
  NAND2_X1  g0124(.A1(new_n324), .A2(new_n294), .ZN(new_n325));
  AND2_X1   g0125(.A1(new_n289), .A2(new_n286), .ZN(new_n326));
  INV_X1    g0126(.A(new_n296), .ZN(new_n327));
  OAI221_X1 g0127(.A(new_n325), .B1(new_n207), .B2(new_n259), .C1(new_n326), .C2(new_n327), .ZN(new_n328));
  AOI21_X1  g0128(.A(new_n323), .B1(new_n283), .B2(new_n328), .ZN(new_n329));
  OR3_X1    g0129(.A1(new_n321), .A2(new_n329), .A3(KEYINPUT73), .ZN(new_n330));
  INV_X1    g0130(.A(G179), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n320), .A2(new_n331), .ZN(new_n332));
  OAI21_X1  g0132(.A(KEYINPUT73), .B1(new_n321), .B2(new_n329), .ZN(new_n333));
  NAND3_X1  g0133(.A1(new_n330), .A2(new_n332), .A3(new_n333), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n320), .A2(G190), .ZN(new_n335));
  INV_X1    g0135(.A(G200), .ZN(new_n336));
  OAI211_X1 g0136(.A(new_n335), .B(new_n329), .C1(new_n336), .C2(new_n320), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n334), .A2(new_n337), .ZN(new_n338));
  INV_X1    g0138(.A(KEYINPUT74), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n338), .A2(new_n339), .ZN(new_n340));
  OR2_X1    g0140(.A1(new_n278), .A2(G179), .ZN(new_n341));
  INV_X1    g0141(.A(G169), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n278), .A2(new_n342), .ZN(new_n343));
  NAND3_X1  g0143(.A1(new_n305), .A2(new_n341), .A3(new_n343), .ZN(new_n344));
  NAND3_X1  g0144(.A1(new_n311), .A2(new_n340), .A3(new_n344), .ZN(new_n345));
  NOR2_X1   g0145(.A1(new_n292), .A2(new_n300), .ZN(new_n346));
  AOI21_X1  g0146(.A(new_n346), .B1(new_n292), .B2(new_n303), .ZN(new_n347));
  AND3_X1   g0147(.A1(new_n262), .A2(KEYINPUT79), .A3(G33), .ZN(new_n348));
  AOI21_X1  g0148(.A(KEYINPUT79), .B1(new_n262), .B2(G33), .ZN(new_n349));
  OAI21_X1  g0149(.A(new_n261), .B1(new_n348), .B2(new_n349), .ZN(new_n350));
  INV_X1    g0150(.A(KEYINPUT7), .ZN(new_n351));
  NAND3_X1  g0151(.A1(new_n350), .A2(new_n351), .A3(new_n207), .ZN(new_n352));
  NOR2_X1   g0152(.A1(new_n262), .A2(G33), .ZN(new_n353));
  INV_X1    g0153(.A(KEYINPUT79), .ZN(new_n354));
  OAI21_X1  g0154(.A(new_n354), .B1(new_n260), .B2(KEYINPUT3), .ZN(new_n355));
  NAND3_X1  g0155(.A1(new_n262), .A2(KEYINPUT79), .A3(G33), .ZN(new_n356));
  AOI21_X1  g0156(.A(new_n353), .B1(new_n355), .B2(new_n356), .ZN(new_n357));
  OAI21_X1  g0157(.A(KEYINPUT7), .B1(new_n357), .B2(G20), .ZN(new_n358));
  NAND3_X1  g0158(.A1(new_n352), .A2(new_n358), .A3(G68), .ZN(new_n359));
  INV_X1    g0159(.A(KEYINPUT80), .ZN(new_n360));
  INV_X1    g0160(.A(G159), .ZN(new_n361));
  NOR2_X1   g0161(.A1(new_n327), .A2(new_n361), .ZN(new_n362));
  INV_X1    g0162(.A(new_n362), .ZN(new_n363));
  AOI21_X1  g0163(.A(new_n202), .B1(new_n220), .B2(G58), .ZN(new_n364));
  OAI211_X1 g0164(.A(new_n360), .B(new_n363), .C1(new_n364), .C2(new_n207), .ZN(new_n365));
  AND2_X1   g0165(.A1(KEYINPUT66), .A2(G68), .ZN(new_n366));
  NOR2_X1   g0166(.A1(KEYINPUT66), .A2(G68), .ZN(new_n367));
  OAI21_X1  g0167(.A(G58), .B1(new_n366), .B2(new_n367), .ZN(new_n368));
  AOI21_X1  g0168(.A(new_n207), .B1(new_n368), .B2(new_n235), .ZN(new_n369));
  OAI21_X1  g0169(.A(KEYINPUT80), .B1(new_n369), .B2(new_n362), .ZN(new_n370));
  NAND4_X1  g0170(.A1(new_n359), .A2(KEYINPUT16), .A3(new_n365), .A4(new_n370), .ZN(new_n371));
  AND2_X1   g0171(.A1(new_n371), .A2(new_n283), .ZN(new_n372));
  INV_X1    g0172(.A(KEYINPUT16), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n370), .A2(new_n365), .ZN(new_n374));
  INV_X1    g0174(.A(KEYINPUT81), .ZN(new_n375));
  OAI21_X1  g0175(.A(new_n375), .B1(new_n262), .B2(G33), .ZN(new_n376));
  NAND3_X1  g0176(.A1(new_n260), .A2(KEYINPUT81), .A3(KEYINPUT3), .ZN(new_n377));
  NAND3_X1  g0177(.A1(new_n376), .A2(new_n263), .A3(new_n377), .ZN(new_n378));
  AOI21_X1  g0178(.A(new_n351), .B1(new_n378), .B2(new_n207), .ZN(new_n379));
  NOR2_X1   g0179(.A1(new_n366), .A2(new_n367), .ZN(new_n380));
  NOR3_X1   g0180(.A1(new_n315), .A2(KEYINPUT7), .A3(G20), .ZN(new_n381));
  NOR3_X1   g0181(.A1(new_n379), .A2(new_n380), .A3(new_n381), .ZN(new_n382));
  OAI21_X1  g0182(.A(new_n373), .B1(new_n374), .B2(new_n382), .ZN(new_n383));
  AOI21_X1  g0183(.A(new_n347), .B1(new_n372), .B2(new_n383), .ZN(new_n384));
  NAND3_X1  g0184(.A1(new_n271), .A2(new_n276), .A3(G232), .ZN(new_n385));
  NAND2_X1  g0185(.A1(new_n275), .A2(new_n385), .ZN(new_n386));
  NOR2_X1   g0186(.A1(G223), .A2(G1698), .ZN(new_n387));
  INV_X1    g0187(.A(G226), .ZN(new_n388));
  AOI21_X1  g0188(.A(new_n387), .B1(new_n388), .B2(G1698), .ZN(new_n389));
  AOI22_X1  g0189(.A1(new_n357), .A2(new_n389), .B1(G33), .B2(G87), .ZN(new_n390));
  AOI21_X1  g0190(.A(new_n258), .B1(new_n390), .B2(KEYINPUT82), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n357), .A2(new_n389), .ZN(new_n392));
  NAND2_X1  g0192(.A1(G33), .A2(G87), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n392), .A2(new_n393), .ZN(new_n394));
  INV_X1    g0194(.A(KEYINPUT82), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n394), .A2(new_n395), .ZN(new_n396));
  AOI21_X1  g0196(.A(new_n386), .B1(new_n391), .B2(new_n396), .ZN(new_n397));
  NOR2_X1   g0197(.A1(new_n397), .A2(new_n342), .ZN(new_n398));
  AOI211_X1 g0198(.A(new_n331), .B(new_n386), .C1(new_n391), .C2(new_n396), .ZN(new_n399));
  NOR2_X1   g0199(.A1(new_n398), .A2(new_n399), .ZN(new_n400));
  OAI21_X1  g0200(.A(KEYINPUT18), .B1(new_n384), .B2(new_n400), .ZN(new_n401));
  NAND3_X1  g0201(.A1(new_n383), .A2(new_n283), .A3(new_n371), .ZN(new_n402));
  INV_X1    g0202(.A(new_n347), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n402), .A2(new_n403), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n397), .A2(G179), .ZN(new_n405));
  OAI21_X1  g0205(.A(new_n405), .B1(new_n342), .B2(new_n397), .ZN(new_n406));
  INV_X1    g0206(.A(KEYINPUT18), .ZN(new_n407));
  NAND3_X1  g0207(.A1(new_n404), .A2(new_n406), .A3(new_n407), .ZN(new_n408));
  INV_X1    g0208(.A(new_n386), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n388), .A2(G1698), .ZN(new_n410));
  OAI21_X1  g0210(.A(new_n410), .B1(G223), .B2(G1698), .ZN(new_n411));
  OAI211_X1 g0211(.A(KEYINPUT82), .B(new_n393), .C1(new_n350), .C2(new_n411), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n412), .A2(new_n314), .ZN(new_n413));
  AOI21_X1  g0213(.A(KEYINPUT82), .B1(new_n392), .B2(new_n393), .ZN(new_n414));
  OAI211_X1 g0214(.A(new_n280), .B(new_n409), .C1(new_n413), .C2(new_n414), .ZN(new_n415));
  OAI21_X1  g0215(.A(new_n415), .B1(new_n397), .B2(G200), .ZN(new_n416));
  NAND3_X1  g0216(.A1(new_n402), .A2(new_n416), .A3(new_n403), .ZN(new_n417));
  INV_X1    g0217(.A(KEYINPUT17), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n417), .A2(new_n418), .ZN(new_n419));
  NAND4_X1  g0219(.A1(new_n402), .A2(new_n416), .A3(KEYINPUT17), .A4(new_n403), .ZN(new_n420));
  NAND4_X1  g0220(.A1(new_n401), .A2(new_n408), .A3(new_n419), .A4(new_n420), .ZN(new_n421));
  INV_X1    g0221(.A(KEYINPUT12), .ZN(new_n422));
  AOI21_X1  g0222(.A(new_n422), .B1(new_n380), .B2(new_n300), .ZN(new_n423));
  XNOR2_X1  g0223(.A(new_n423), .B(KEYINPUT77), .ZN(new_n424));
  INV_X1    g0224(.A(G68), .ZN(new_n425));
  NAND3_X1  g0225(.A1(new_n300), .A2(new_n422), .A3(new_n425), .ZN(new_n426));
  AOI22_X1  g0226(.A1(new_n424), .A2(new_n426), .B1(G68), .B2(new_n302), .ZN(new_n427));
  NOR2_X1   g0227(.A1(new_n220), .A2(new_n207), .ZN(new_n428));
  OAI22_X1  g0228(.A1(new_n327), .A2(new_n234), .B1(new_n293), .B2(new_n259), .ZN(new_n429));
  OAI21_X1  g0229(.A(new_n283), .B1(new_n428), .B2(new_n429), .ZN(new_n430));
  XNOR2_X1  g0230(.A(new_n430), .B(KEYINPUT11), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n427), .A2(new_n431), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n432), .A2(KEYINPUT78), .ZN(new_n433));
  AND2_X1   g0233(.A1(new_n427), .A2(new_n431), .ZN(new_n434));
  INV_X1    g0234(.A(KEYINPUT78), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n434), .A2(new_n435), .ZN(new_n436));
  NAND4_X1  g0236(.A1(new_n261), .A2(new_n263), .A3(G232), .A4(G1698), .ZN(new_n437));
  NAND2_X1  g0237(.A1(new_n437), .A2(KEYINPUT76), .ZN(new_n438));
  INV_X1    g0238(.A(KEYINPUT76), .ZN(new_n439));
  NAND4_X1  g0239(.A1(new_n315), .A2(new_n439), .A3(G232), .A4(G1698), .ZN(new_n440));
  NAND2_X1  g0240(.A1(new_n438), .A2(new_n440), .ZN(new_n441));
  NAND4_X1  g0241(.A1(new_n261), .A2(new_n263), .A3(G226), .A4(new_n317), .ZN(new_n442));
  NAND2_X1  g0242(.A1(G33), .A2(G97), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  INV_X1    g0244(.A(new_n444), .ZN(new_n445));
  AOI21_X1  g0245(.A(new_n258), .B1(new_n441), .B2(new_n445), .ZN(new_n446));
  NAND3_X1  g0246(.A1(new_n271), .A2(new_n276), .A3(G238), .ZN(new_n447));
  NAND2_X1  g0247(.A1(new_n275), .A2(new_n447), .ZN(new_n448));
  OAI21_X1  g0248(.A(KEYINPUT13), .B1(new_n446), .B2(new_n448), .ZN(new_n449));
  INV_X1    g0249(.A(new_n448), .ZN(new_n450));
  INV_X1    g0250(.A(KEYINPUT13), .ZN(new_n451));
  AOI21_X1  g0251(.A(new_n444), .B1(new_n440), .B2(new_n438), .ZN(new_n452));
  OAI211_X1 g0252(.A(new_n450), .B(new_n451), .C1(new_n452), .C2(new_n258), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n449), .A2(new_n453), .ZN(new_n454));
  INV_X1    g0254(.A(KEYINPUT14), .ZN(new_n455));
  NAND3_X1  g0255(.A1(new_n454), .A2(new_n455), .A3(G169), .ZN(new_n456));
  NAND3_X1  g0256(.A1(new_n449), .A2(new_n453), .A3(G179), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n456), .A2(new_n457), .ZN(new_n458));
  AOI21_X1  g0258(.A(new_n455), .B1(new_n454), .B2(G169), .ZN(new_n459));
  OAI211_X1 g0259(.A(new_n433), .B(new_n436), .C1(new_n458), .C2(new_n459), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n454), .A2(G200), .ZN(new_n461));
  NAND3_X1  g0261(.A1(new_n449), .A2(new_n453), .A3(G190), .ZN(new_n462));
  NAND3_X1  g0262(.A1(new_n461), .A2(new_n434), .A3(new_n462), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n460), .A2(new_n463), .ZN(new_n464));
  NOR2_X1   g0264(.A1(new_n338), .A2(new_n339), .ZN(new_n465));
  NOR4_X1   g0265(.A1(new_n345), .A2(new_n421), .A3(new_n464), .A4(new_n465), .ZN(new_n466));
  NOR2_X1   g0266(.A1(new_n299), .A2(G116), .ZN(new_n467));
  OAI21_X1  g0267(.A(new_n299), .B1(G1), .B2(new_n260), .ZN(new_n468));
  NOR2_X1   g0268(.A1(new_n468), .A2(new_n283), .ZN(new_n469));
  AOI21_X1  g0269(.A(new_n467), .B1(new_n469), .B2(G116), .ZN(new_n470));
  NAND2_X1  g0270(.A1(G33), .A2(G283), .ZN(new_n471));
  OAI211_X1 g0271(.A(new_n471), .B(new_n207), .C1(G33), .C2(new_n216), .ZN(new_n472));
  INV_X1    g0272(.A(G116), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n473), .A2(G20), .ZN(new_n474));
  NAND3_X1  g0274(.A1(new_n472), .A2(new_n283), .A3(new_n474), .ZN(new_n475));
  INV_X1    g0275(.A(KEYINPUT20), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n475), .A2(new_n476), .ZN(new_n477));
  NAND4_X1  g0277(.A1(new_n472), .A2(KEYINPUT20), .A3(new_n283), .A4(new_n474), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  AOI21_X1  g0279(.A(new_n342), .B1(new_n470), .B2(new_n479), .ZN(new_n480));
  NOR2_X1   g0280(.A1(new_n217), .A2(G1698), .ZN(new_n481));
  OAI211_X1 g0281(.A(new_n261), .B(new_n481), .C1(new_n348), .C2(new_n349), .ZN(new_n482));
  INV_X1    g0282(.A(KEYINPUT88), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n482), .A2(new_n483), .ZN(new_n484));
  NAND3_X1  g0284(.A1(new_n357), .A2(KEYINPUT88), .A3(new_n481), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n484), .A2(new_n485), .ZN(new_n486));
  NOR2_X1   g0286(.A1(new_n211), .A2(new_n317), .ZN(new_n487));
  OAI211_X1 g0287(.A(new_n261), .B(new_n487), .C1(new_n348), .C2(new_n349), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n264), .A2(G303), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  INV_X1    g0290(.A(new_n490), .ZN(new_n491));
  AOI21_X1  g0291(.A(new_n258), .B1(new_n486), .B2(new_n491), .ZN(new_n492));
  INV_X1    g0292(.A(KEYINPUT5), .ZN(new_n493));
  OAI21_X1  g0293(.A(KEYINPUT84), .B1(new_n493), .B2(G41), .ZN(new_n494));
  INV_X1    g0294(.A(KEYINPUT84), .ZN(new_n495));
  NAND3_X1  g0295(.A1(new_n495), .A2(new_n272), .A3(KEYINPUT5), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n494), .A2(new_n496), .ZN(new_n497));
  NOR2_X1   g0297(.A1(new_n272), .A2(KEYINPUT5), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n206), .A2(G45), .ZN(new_n499));
  NOR2_X1   g0299(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  NAND4_X1  g0300(.A1(new_n271), .A2(new_n497), .A3(new_n500), .A4(G274), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n493), .A2(G41), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n272), .A2(KEYINPUT5), .ZN(new_n503));
  NAND4_X1  g0303(.A1(new_n502), .A2(new_n503), .A3(new_n206), .A4(G45), .ZN(new_n504));
  NAND3_X1  g0304(.A1(new_n504), .A2(new_n271), .A3(G270), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n501), .A2(new_n505), .ZN(new_n506));
  OAI211_X1 g0306(.A(new_n480), .B(KEYINPUT21), .C1(new_n492), .C2(new_n506), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n507), .A2(KEYINPUT89), .ZN(new_n508));
  INV_X1    g0308(.A(new_n506), .ZN(new_n509));
  AOI21_X1  g0309(.A(new_n490), .B1(new_n484), .B2(new_n485), .ZN(new_n510));
  OAI21_X1  g0310(.A(new_n509), .B1(new_n510), .B2(new_n258), .ZN(new_n511));
  INV_X1    g0311(.A(KEYINPUT89), .ZN(new_n512));
  NAND4_X1  g0312(.A1(new_n511), .A2(new_n512), .A3(KEYINPUT21), .A4(new_n480), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n508), .A2(new_n513), .ZN(new_n514));
  AOI21_X1  g0314(.A(KEYINPUT21), .B1(new_n511), .B2(new_n480), .ZN(new_n515));
  OAI211_X1 g0315(.A(G179), .B(new_n509), .C1(new_n510), .C2(new_n258), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n470), .A2(new_n479), .ZN(new_n517));
  INV_X1    g0317(.A(new_n517), .ZN(new_n518));
  NOR2_X1   g0318(.A1(new_n516), .A2(new_n518), .ZN(new_n519));
  NOR2_X1   g0319(.A1(new_n515), .A2(new_n519), .ZN(new_n520));
  AOI21_X1  g0320(.A(new_n517), .B1(new_n511), .B2(G200), .ZN(new_n521));
  OAI21_X1  g0321(.A(new_n521), .B1(new_n280), .B2(new_n511), .ZN(new_n522));
  AND3_X1   g0322(.A1(new_n514), .A2(new_n520), .A3(new_n522), .ZN(new_n523));
  NAND3_X1  g0323(.A1(new_n504), .A2(new_n271), .A3(G264), .ZN(new_n524));
  NOR2_X1   g0324(.A1(G250), .A2(G1698), .ZN(new_n525));
  AOI21_X1  g0325(.A(new_n525), .B1(new_n217), .B2(G1698), .ZN(new_n526));
  AOI22_X1  g0326(.A1(new_n357), .A2(new_n526), .B1(G33), .B2(G294), .ZN(new_n527));
  OAI211_X1 g0327(.A(new_n501), .B(new_n524), .C1(new_n527), .C2(new_n258), .ZN(new_n528));
  NOR2_X1   g0328(.A1(new_n528), .A2(G179), .ZN(new_n529));
  AOI21_X1  g0329(.A(new_n529), .B1(new_n342), .B2(new_n528), .ZN(new_n530));
  NAND3_X1  g0330(.A1(new_n357), .A2(new_n207), .A3(G87), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n531), .A2(KEYINPUT22), .ZN(new_n532));
  NAND4_X1  g0332(.A1(new_n261), .A2(new_n263), .A3(new_n207), .A4(G87), .ZN(new_n533));
  XNOR2_X1  g0333(.A(KEYINPUT90), .B(KEYINPUT22), .ZN(new_n534));
  NOR2_X1   g0334(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  INV_X1    g0335(.A(new_n535), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n532), .A2(new_n536), .ZN(new_n537));
  INV_X1    g0337(.A(KEYINPUT24), .ZN(new_n538));
  AOI21_X1  g0338(.A(KEYINPUT23), .B1(new_n210), .B2(G20), .ZN(new_n539));
  INV_X1    g0339(.A(new_n539), .ZN(new_n540));
  NAND3_X1  g0340(.A1(new_n210), .A2(KEYINPUT23), .A3(G20), .ZN(new_n541));
  NOR2_X1   g0341(.A1(new_n260), .A2(new_n473), .ZN(new_n542));
  AOI22_X1  g0342(.A1(new_n540), .A2(new_n541), .B1(new_n542), .B2(new_n207), .ZN(new_n543));
  NAND3_X1  g0343(.A1(new_n537), .A2(new_n538), .A3(new_n543), .ZN(new_n544));
  AOI21_X1  g0344(.A(new_n535), .B1(new_n531), .B2(KEYINPUT22), .ZN(new_n545));
  INV_X1    g0345(.A(new_n543), .ZN(new_n546));
  OAI21_X1  g0346(.A(KEYINPUT24), .B1(new_n545), .B2(new_n546), .ZN(new_n547));
  AOI21_X1  g0347(.A(new_n284), .B1(new_n544), .B2(new_n547), .ZN(new_n548));
  AOI21_X1  g0348(.A(KEYINPUT25), .B1(new_n300), .B2(new_n210), .ZN(new_n549));
  INV_X1    g0349(.A(new_n549), .ZN(new_n550));
  NAND3_X1  g0350(.A1(new_n300), .A2(KEYINPUT25), .A3(new_n210), .ZN(new_n551));
  AOI22_X1  g0351(.A1(new_n550), .A2(new_n551), .B1(new_n469), .B2(G107), .ZN(new_n552));
  INV_X1    g0352(.A(new_n552), .ZN(new_n553));
  OAI21_X1  g0353(.A(new_n530), .B1(new_n548), .B2(new_n553), .ZN(new_n554));
  AOI21_X1  g0354(.A(new_n538), .B1(new_n537), .B2(new_n543), .ZN(new_n555));
  NOR3_X1   g0355(.A1(new_n545), .A2(KEYINPUT24), .A3(new_n546), .ZN(new_n556));
  OAI21_X1  g0356(.A(new_n283), .B1(new_n555), .B2(new_n556), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n528), .A2(new_n336), .ZN(new_n558));
  OAI21_X1  g0358(.A(new_n558), .B1(G190), .B2(new_n528), .ZN(new_n559));
  NAND3_X1  g0359(.A1(new_n557), .A2(new_n552), .A3(new_n559), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n554), .A2(new_n560), .ZN(new_n561));
  INV_X1    g0361(.A(G244), .ZN(new_n562));
  NOR2_X1   g0362(.A1(new_n562), .A2(G1698), .ZN(new_n563));
  AOI21_X1  g0363(.A(KEYINPUT4), .B1(new_n357), .B2(new_n563), .ZN(new_n564));
  NAND4_X1  g0364(.A1(new_n261), .A2(new_n263), .A3(G250), .A4(G1698), .ZN(new_n565));
  AND2_X1   g0365(.A1(KEYINPUT4), .A2(G244), .ZN(new_n566));
  NAND4_X1  g0366(.A1(new_n261), .A2(new_n263), .A3(new_n566), .A4(new_n317), .ZN(new_n567));
  NAND3_X1  g0367(.A1(new_n565), .A2(new_n567), .A3(new_n471), .ZN(new_n568));
  OAI21_X1  g0368(.A(new_n314), .B1(new_n564), .B2(new_n568), .ZN(new_n569));
  NAND3_X1  g0369(.A1(new_n504), .A2(new_n271), .A3(G257), .ZN(new_n570));
  AND2_X1   g0370(.A1(new_n501), .A2(new_n570), .ZN(new_n571));
  NAND3_X1  g0371(.A1(new_n569), .A2(new_n571), .A3(new_n280), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n501), .A2(new_n570), .ZN(new_n573));
  AND3_X1   g0373(.A1(new_n565), .A2(new_n567), .A3(new_n471), .ZN(new_n574));
  OAI211_X1 g0374(.A(new_n261), .B(new_n563), .C1(new_n348), .C2(new_n349), .ZN(new_n575));
  INV_X1    g0375(.A(KEYINPUT4), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n575), .A2(new_n576), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n574), .A2(new_n577), .ZN(new_n578));
  AOI21_X1  g0378(.A(new_n573), .B1(new_n578), .B2(new_n314), .ZN(new_n579));
  OAI21_X1  g0379(.A(new_n572), .B1(new_n579), .B2(G200), .ZN(new_n580));
  NOR2_X1   g0380(.A1(new_n299), .A2(G97), .ZN(new_n581));
  AOI21_X1  g0381(.A(new_n581), .B1(new_n469), .B2(G97), .ZN(new_n582));
  INV_X1    g0382(.A(KEYINPUT83), .ZN(new_n583));
  NAND3_X1  g0383(.A1(new_n264), .A2(new_n351), .A3(new_n207), .ZN(new_n584));
  AOI21_X1  g0384(.A(KEYINPUT81), .B1(new_n260), .B2(KEYINPUT3), .ZN(new_n585));
  NOR2_X1   g0385(.A1(new_n260), .A2(KEYINPUT3), .ZN(new_n586));
  NOR2_X1   g0386(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  AOI21_X1  g0387(.A(G20), .B1(new_n587), .B2(new_n377), .ZN(new_n588));
  OAI211_X1 g0388(.A(G107), .B(new_n584), .C1(new_n588), .C2(new_n351), .ZN(new_n589));
  XNOR2_X1  g0389(.A(G97), .B(G107), .ZN(new_n590));
  INV_X1    g0390(.A(KEYINPUT6), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  NOR3_X1   g0392(.A1(new_n591), .A2(new_n216), .A3(G107), .ZN(new_n593));
  INV_X1    g0393(.A(new_n593), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n592), .A2(new_n594), .ZN(new_n595));
  AOI22_X1  g0395(.A1(new_n595), .A2(G20), .B1(G77), .B2(new_n296), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n589), .A2(new_n596), .ZN(new_n597));
  AOI21_X1  g0397(.A(new_n583), .B1(new_n597), .B2(new_n283), .ZN(new_n598));
  AOI211_X1 g0398(.A(KEYINPUT83), .B(new_n284), .C1(new_n589), .C2(new_n596), .ZN(new_n599));
  OAI211_X1 g0399(.A(new_n580), .B(new_n582), .C1(new_n598), .C2(new_n599), .ZN(new_n600));
  INV_X1    g0400(.A(new_n582), .ZN(new_n601));
  NOR3_X1   g0401(.A1(new_n379), .A2(new_n210), .A3(new_n381), .ZN(new_n602));
  AOI21_X1  g0402(.A(new_n593), .B1(new_n591), .B2(new_n590), .ZN(new_n603));
  OAI22_X1  g0403(.A1(new_n603), .A2(new_n207), .B1(new_n259), .B2(new_n327), .ZN(new_n604));
  NOR2_X1   g0404(.A1(new_n602), .A2(new_n604), .ZN(new_n605));
  OAI21_X1  g0405(.A(KEYINPUT83), .B1(new_n605), .B2(new_n284), .ZN(new_n606));
  NAND3_X1  g0406(.A1(new_n597), .A2(new_n583), .A3(new_n283), .ZN(new_n607));
  AOI21_X1  g0407(.A(new_n601), .B1(new_n606), .B2(new_n607), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n579), .A2(new_n331), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n569), .A2(new_n571), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n610), .A2(new_n342), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n609), .A2(new_n611), .ZN(new_n612));
  OAI21_X1  g0412(.A(new_n600), .B1(new_n608), .B2(new_n612), .ZN(new_n613));
  NOR2_X1   g0413(.A1(new_n324), .A2(new_n299), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n355), .A2(new_n356), .ZN(new_n615));
  NAND4_X1  g0415(.A1(new_n615), .A2(new_n207), .A3(G68), .A4(new_n261), .ZN(new_n616));
  INV_X1    g0416(.A(KEYINPUT19), .ZN(new_n617));
  OAI21_X1  g0417(.A(new_n617), .B1(new_n293), .B2(new_n216), .ZN(new_n618));
  NAND3_X1  g0418(.A1(KEYINPUT19), .A2(G33), .A3(G97), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n619), .A2(new_n207), .ZN(new_n620));
  INV_X1    g0420(.A(KEYINPUT86), .ZN(new_n621));
  NAND3_X1  g0421(.A1(new_n214), .A2(new_n216), .A3(new_n210), .ZN(new_n622));
  AND3_X1   g0422(.A1(new_n620), .A2(new_n621), .A3(new_n622), .ZN(new_n623));
  AOI21_X1  g0423(.A(new_n621), .B1(new_n620), .B2(new_n622), .ZN(new_n624));
  OAI211_X1 g0424(.A(new_n616), .B(new_n618), .C1(new_n623), .C2(new_n624), .ZN(new_n625));
  INV_X1    g0425(.A(KEYINPUT87), .ZN(new_n626));
  AOI21_X1  g0426(.A(new_n284), .B1(new_n625), .B2(new_n626), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n620), .A2(new_n622), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n628), .A2(KEYINPUT86), .ZN(new_n629));
  NAND3_X1  g0429(.A1(new_n620), .A2(new_n621), .A3(new_n622), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  NAND4_X1  g0431(.A1(new_n631), .A2(KEYINPUT87), .A3(new_n616), .A4(new_n618), .ZN(new_n632));
  AOI21_X1  g0432(.A(new_n614), .B1(new_n627), .B2(new_n632), .ZN(new_n633));
  INV_X1    g0433(.A(new_n469), .ZN(new_n634));
  NOR2_X1   g0434(.A1(new_n634), .A2(new_n214), .ZN(new_n635));
  INV_X1    g0435(.A(new_n635), .ZN(new_n636));
  NOR2_X1   g0436(.A1(G238), .A2(G1698), .ZN(new_n637));
  AOI21_X1  g0437(.A(new_n637), .B1(new_n562), .B2(G1698), .ZN(new_n638));
  AOI21_X1  g0438(.A(new_n542), .B1(new_n357), .B2(new_n638), .ZN(new_n639));
  INV_X1    g0439(.A(KEYINPUT85), .ZN(new_n640));
  AOI21_X1  g0440(.A(new_n258), .B1(new_n639), .B2(new_n640), .ZN(new_n641));
  INV_X1    g0441(.A(new_n542), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n562), .A2(G1698), .ZN(new_n643));
  OAI21_X1  g0443(.A(new_n643), .B1(G238), .B2(G1698), .ZN(new_n644));
  OAI21_X1  g0444(.A(new_n642), .B1(new_n350), .B2(new_n644), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n645), .A2(KEYINPUT85), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n641), .A2(new_n646), .ZN(new_n647));
  OR2_X1    g0447(.A1(new_n499), .A2(G274), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n499), .A2(new_n215), .ZN(new_n649));
  NAND3_X1  g0449(.A1(new_n648), .A2(new_n271), .A3(new_n649), .ZN(new_n650));
  AOI21_X1  g0450(.A(G200), .B1(new_n647), .B2(new_n650), .ZN(new_n651));
  INV_X1    g0451(.A(new_n650), .ZN(new_n652));
  AOI211_X1 g0452(.A(G190), .B(new_n652), .C1(new_n641), .C2(new_n646), .ZN(new_n653));
  OAI211_X1 g0453(.A(new_n633), .B(new_n636), .C1(new_n651), .C2(new_n653), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n616), .A2(new_n618), .ZN(new_n655));
  NOR2_X1   g0455(.A1(new_n623), .A2(new_n624), .ZN(new_n656));
  OAI21_X1  g0456(.A(new_n626), .B1(new_n655), .B2(new_n656), .ZN(new_n657));
  NAND3_X1  g0457(.A1(new_n657), .A2(new_n283), .A3(new_n632), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n469), .A2(new_n324), .ZN(new_n659));
  INV_X1    g0459(.A(new_n614), .ZN(new_n660));
  NAND3_X1  g0460(.A1(new_n658), .A2(new_n659), .A3(new_n660), .ZN(new_n661));
  AOI21_X1  g0461(.A(new_n652), .B1(new_n641), .B2(new_n646), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n662), .A2(new_n331), .ZN(new_n663));
  OAI211_X1 g0463(.A(new_n640), .B(new_n642), .C1(new_n350), .C2(new_n644), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n664), .A2(new_n314), .ZN(new_n665));
  NOR2_X1   g0465(.A1(new_n639), .A2(new_n640), .ZN(new_n666));
  OAI21_X1  g0466(.A(new_n650), .B1(new_n665), .B2(new_n666), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n667), .A2(new_n342), .ZN(new_n668));
  NAND3_X1  g0468(.A1(new_n661), .A2(new_n663), .A3(new_n668), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n654), .A2(new_n669), .ZN(new_n670));
  NOR3_X1   g0470(.A1(new_n561), .A2(new_n613), .A3(new_n670), .ZN(new_n671));
  AND3_X1   g0471(.A1(new_n466), .A2(new_n523), .A3(new_n671), .ZN(G372));
  INV_X1    g0472(.A(new_n344), .ZN(new_n673));
  AND3_X1   g0473(.A1(new_n404), .A2(new_n407), .A3(new_n406), .ZN(new_n674));
  AOI21_X1  g0474(.A(new_n407), .B1(new_n404), .B2(new_n406), .ZN(new_n675));
  NOR2_X1   g0475(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  NAND4_X1  g0476(.A1(new_n463), .A2(new_n330), .A3(new_n332), .A4(new_n333), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n460), .A2(new_n677), .ZN(new_n678));
  INV_X1    g0478(.A(KEYINPUT91), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  AND2_X1   g0480(.A1(new_n419), .A2(new_n420), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  NOR2_X1   g0482(.A1(new_n678), .A2(new_n679), .ZN(new_n683));
  OAI21_X1  g0483(.A(new_n676), .B1(new_n682), .B2(new_n683), .ZN(new_n684));
  AOI21_X1  g0484(.A(new_n673), .B1(new_n684), .B2(new_n311), .ZN(new_n685));
  INV_X1    g0485(.A(new_n669), .ZN(new_n686));
  INV_X1    g0486(.A(KEYINPUT26), .ZN(new_n687));
  OAI21_X1  g0487(.A(new_n582), .B1(new_n598), .B2(new_n599), .ZN(new_n688));
  INV_X1    g0488(.A(new_n612), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  OAI21_X1  g0490(.A(new_n687), .B1(new_n670), .B2(new_n690), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n606), .A2(new_n607), .ZN(new_n692));
  AOI21_X1  g0492(.A(new_n612), .B1(new_n692), .B2(new_n582), .ZN(new_n693));
  NAND4_X1  g0493(.A1(new_n693), .A2(KEYINPUT26), .A3(new_n669), .A4(new_n654), .ZN(new_n694));
  AOI21_X1  g0494(.A(new_n686), .B1(new_n691), .B2(new_n694), .ZN(new_n695));
  NOR2_X1   g0495(.A1(new_n613), .A2(new_n670), .ZN(new_n696));
  NAND3_X1  g0496(.A1(new_n514), .A2(new_n520), .A3(new_n554), .ZN(new_n697));
  NAND3_X1  g0497(.A1(new_n696), .A2(new_n560), .A3(new_n697), .ZN(new_n698));
  NAND2_X1  g0498(.A1(new_n695), .A2(new_n698), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n466), .A2(new_n699), .ZN(new_n700));
  NAND2_X1  g0500(.A1(new_n685), .A2(new_n700), .ZN(G369));
  NAND3_X1  g0501(.A1(new_n206), .A2(new_n207), .A3(G13), .ZN(new_n702));
  OR2_X1    g0502(.A1(new_n702), .A2(KEYINPUT27), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n702), .A2(KEYINPUT27), .ZN(new_n704));
  NAND3_X1  g0504(.A1(new_n703), .A2(G213), .A3(new_n704), .ZN(new_n705));
  INV_X1    g0505(.A(G343), .ZN(new_n706));
  NOR2_X1   g0506(.A1(new_n705), .A2(new_n706), .ZN(new_n707));
  INV_X1    g0507(.A(new_n707), .ZN(new_n708));
  NOR2_X1   g0508(.A1(new_n518), .A2(new_n708), .ZN(new_n709));
  INV_X1    g0509(.A(new_n709), .ZN(new_n710));
  NAND2_X1  g0510(.A1(new_n523), .A2(new_n710), .ZN(new_n711));
  AND2_X1   g0511(.A1(new_n514), .A2(new_n520), .ZN(new_n712));
  OAI21_X1  g0512(.A(new_n711), .B1(new_n712), .B2(new_n710), .ZN(new_n713));
  XNOR2_X1  g0513(.A(KEYINPUT92), .B(G330), .ZN(new_n714));
  AND2_X1   g0514(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  AOI21_X1  g0515(.A(new_n708), .B1(new_n557), .B2(new_n552), .ZN(new_n716));
  OAI22_X1  g0516(.A1(new_n561), .A2(new_n716), .B1(new_n554), .B2(new_n708), .ZN(new_n717));
  NAND2_X1  g0517(.A1(new_n715), .A2(new_n717), .ZN(new_n718));
  NOR2_X1   g0518(.A1(new_n712), .A2(new_n707), .ZN(new_n719));
  INV_X1    g0519(.A(new_n561), .ZN(new_n720));
  INV_X1    g0520(.A(new_n554), .ZN(new_n721));
  AOI22_X1  g0521(.A1(new_n719), .A2(new_n720), .B1(new_n721), .B2(new_n708), .ZN(new_n722));
  NAND2_X1  g0522(.A1(new_n718), .A2(new_n722), .ZN(G399));
  NOR2_X1   g0523(.A1(new_n227), .A2(G41), .ZN(new_n724));
  INV_X1    g0524(.A(new_n724), .ZN(new_n725));
  NOR2_X1   g0525(.A1(new_n622), .A2(G116), .ZN(new_n726));
  NAND3_X1  g0526(.A1(new_n725), .A2(G1), .A3(new_n726), .ZN(new_n727));
  OAI21_X1  g0527(.A(new_n727), .B1(new_n237), .B2(new_n725), .ZN(new_n728));
  XNOR2_X1  g0528(.A(new_n728), .B(KEYINPUT28), .ZN(new_n729));
  AOI21_X1  g0529(.A(new_n707), .B1(new_n695), .B2(new_n698), .ZN(new_n730));
  INV_X1    g0530(.A(new_n730), .ZN(new_n731));
  NOR2_X1   g0531(.A1(new_n731), .A2(KEYINPUT29), .ZN(new_n732));
  INV_X1    g0532(.A(KEYINPUT29), .ZN(new_n733));
  INV_X1    g0533(.A(KEYINPUT96), .ZN(new_n734));
  NOR2_X1   g0534(.A1(new_n662), .A2(G169), .ZN(new_n735));
  AOI211_X1 g0535(.A(G179), .B(new_n652), .C1(new_n641), .C2(new_n646), .ZN(new_n736));
  NOR2_X1   g0536(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  AOI211_X1 g0537(.A(new_n614), .B(new_n635), .C1(new_n627), .C2(new_n632), .ZN(new_n738));
  OAI211_X1 g0538(.A(new_n280), .B(new_n650), .C1(new_n665), .C2(new_n666), .ZN(new_n739));
  OAI21_X1  g0539(.A(new_n739), .B1(new_n662), .B2(G200), .ZN(new_n740));
  AOI22_X1  g0540(.A1(new_n737), .A2(new_n661), .B1(new_n738), .B2(new_n740), .ZN(new_n741));
  NAND4_X1  g0541(.A1(new_n741), .A2(new_n560), .A3(new_n690), .A4(new_n600), .ZN(new_n742));
  AND3_X1   g0542(.A1(new_n514), .A2(new_n520), .A3(new_n554), .ZN(new_n743));
  OAI21_X1  g0543(.A(new_n734), .B1(new_n742), .B2(new_n743), .ZN(new_n744));
  NAND4_X1  g0544(.A1(new_n696), .A2(KEYINPUT96), .A3(new_n560), .A4(new_n697), .ZN(new_n745));
  NAND3_X1  g0545(.A1(new_n744), .A2(new_n745), .A3(new_n695), .ZN(new_n746));
  AOI21_X1  g0546(.A(new_n733), .B1(new_n746), .B2(new_n708), .ZN(new_n747));
  NOR2_X1   g0547(.A1(new_n732), .A2(new_n747), .ZN(new_n748));
  INV_X1    g0548(.A(KEYINPUT31), .ZN(new_n749));
  NOR2_X1   g0549(.A1(new_n516), .A2(new_n610), .ZN(new_n750));
  INV_X1    g0550(.A(KEYINPUT93), .ZN(new_n751));
  NAND2_X1  g0551(.A1(new_n357), .A2(new_n526), .ZN(new_n752));
  INV_X1    g0552(.A(G294), .ZN(new_n753));
  OAI21_X1  g0553(.A(new_n752), .B1(new_n260), .B2(new_n753), .ZN(new_n754));
  NAND2_X1  g0554(.A1(new_n754), .A2(new_n314), .ZN(new_n755));
  NAND4_X1  g0555(.A1(new_n662), .A2(new_n751), .A3(new_n524), .A4(new_n755), .ZN(new_n756));
  NAND2_X1  g0556(.A1(new_n755), .A2(new_n524), .ZN(new_n757));
  OAI21_X1  g0557(.A(KEYINPUT93), .B1(new_n667), .B2(new_n757), .ZN(new_n758));
  NAND3_X1  g0558(.A1(new_n750), .A2(new_n756), .A3(new_n758), .ZN(new_n759));
  INV_X1    g0559(.A(KEYINPUT94), .ZN(new_n760));
  INV_X1    g0560(.A(KEYINPUT30), .ZN(new_n761));
  AND3_X1   g0561(.A1(new_n759), .A2(new_n760), .A3(new_n761), .ZN(new_n762));
  AOI21_X1  g0562(.A(new_n760), .B1(new_n759), .B2(new_n761), .ZN(new_n763));
  NAND4_X1  g0563(.A1(new_n750), .A2(new_n758), .A3(new_n756), .A4(KEYINPUT30), .ZN(new_n764));
  AND2_X1   g0564(.A1(new_n528), .A2(new_n331), .ZN(new_n765));
  NAND4_X1  g0565(.A1(new_n765), .A2(new_n511), .A3(new_n610), .A4(new_n667), .ZN(new_n766));
  NAND2_X1  g0566(.A1(new_n764), .A2(new_n766), .ZN(new_n767));
  NOR3_X1   g0567(.A1(new_n762), .A2(new_n763), .A3(new_n767), .ZN(new_n768));
  OAI21_X1  g0568(.A(new_n749), .B1(new_n768), .B2(new_n708), .ZN(new_n769));
  NAND4_X1  g0569(.A1(new_n696), .A2(new_n523), .A3(new_n720), .A4(new_n708), .ZN(new_n770));
  NAND2_X1  g0570(.A1(new_n770), .A2(KEYINPUT95), .ZN(new_n771));
  INV_X1    g0571(.A(new_n767), .ZN(new_n772));
  NAND2_X1  g0572(.A1(new_n759), .A2(new_n761), .ZN(new_n773));
  NAND2_X1  g0573(.A1(new_n772), .A2(new_n773), .ZN(new_n774));
  NAND3_X1  g0574(.A1(new_n774), .A2(KEYINPUT31), .A3(new_n707), .ZN(new_n775));
  INV_X1    g0575(.A(KEYINPUT95), .ZN(new_n776));
  NAND4_X1  g0576(.A1(new_n671), .A2(new_n776), .A3(new_n523), .A4(new_n708), .ZN(new_n777));
  NAND4_X1  g0577(.A1(new_n769), .A2(new_n771), .A3(new_n775), .A4(new_n777), .ZN(new_n778));
  NAND2_X1  g0578(.A1(new_n778), .A2(new_n714), .ZN(new_n779));
  NAND2_X1  g0579(.A1(new_n748), .A2(new_n779), .ZN(new_n780));
  INV_X1    g0580(.A(new_n780), .ZN(new_n781));
  OAI21_X1  g0581(.A(new_n729), .B1(new_n781), .B2(G1), .ZN(G364));
  NOR2_X1   g0582(.A1(new_n226), .A2(G20), .ZN(new_n783));
  AOI21_X1  g0583(.A(new_n206), .B1(new_n783), .B2(G45), .ZN(new_n784));
  INV_X1    g0584(.A(new_n784), .ZN(new_n785));
  NOR2_X1   g0585(.A1(new_n724), .A2(new_n785), .ZN(new_n786));
  NOR2_X1   g0586(.A1(new_n715), .A2(new_n786), .ZN(new_n787));
  OAI21_X1  g0587(.A(new_n787), .B1(new_n714), .B2(new_n713), .ZN(new_n788));
  INV_X1    g0588(.A(new_n786), .ZN(new_n789));
  OAI21_X1  g0589(.A(G20), .B1(KEYINPUT98), .B2(G169), .ZN(new_n790));
  INV_X1    g0590(.A(new_n790), .ZN(new_n791));
  NAND2_X1  g0591(.A1(KEYINPUT98), .A2(G169), .ZN(new_n792));
  AOI21_X1  g0592(.A(new_n231), .B1(new_n791), .B2(new_n792), .ZN(new_n793));
  INV_X1    g0593(.A(new_n793), .ZN(new_n794));
  NOR3_X1   g0594(.A1(new_n207), .A2(new_n331), .A3(KEYINPUT99), .ZN(new_n795));
  INV_X1    g0595(.A(KEYINPUT99), .ZN(new_n796));
  AOI21_X1  g0596(.A(new_n796), .B1(G20), .B2(G179), .ZN(new_n797));
  NOR2_X1   g0597(.A1(new_n795), .A2(new_n797), .ZN(new_n798));
  NOR2_X1   g0598(.A1(new_n280), .A2(new_n336), .ZN(new_n799));
  INV_X1    g0599(.A(new_n799), .ZN(new_n800));
  NOR2_X1   g0600(.A1(new_n798), .A2(new_n800), .ZN(new_n801));
  NOR2_X1   g0601(.A1(new_n280), .A2(G200), .ZN(new_n802));
  NAND2_X1  g0602(.A1(new_n802), .A2(new_n331), .ZN(new_n803));
  NAND2_X1  g0603(.A1(new_n803), .A2(G20), .ZN(new_n804));
  AOI22_X1  g0604(.A1(new_n801), .A2(G326), .B1(G294), .B2(new_n804), .ZN(new_n805));
  INV_X1    g0605(.A(G311), .ZN(new_n806));
  INV_X1    g0606(.A(new_n798), .ZN(new_n807));
  NOR2_X1   g0607(.A1(G190), .A2(G200), .ZN(new_n808));
  NAND2_X1  g0608(.A1(new_n807), .A2(new_n808), .ZN(new_n809));
  OAI21_X1  g0609(.A(new_n805), .B1(new_n806), .B2(new_n809), .ZN(new_n810));
  XOR2_X1   g0610(.A(new_n810), .B(KEYINPUT101), .Z(new_n811));
  INV_X1    g0611(.A(G283), .ZN(new_n812));
  NOR2_X1   g0612(.A1(new_n207), .A2(G179), .ZN(new_n813));
  NOR2_X1   g0613(.A1(new_n336), .A2(G190), .ZN(new_n814));
  NAND2_X1  g0614(.A1(new_n813), .A2(new_n814), .ZN(new_n815));
  INV_X1    g0615(.A(new_n813), .ZN(new_n816));
  NOR2_X1   g0616(.A1(new_n800), .A2(new_n816), .ZN(new_n817));
  INV_X1    g0617(.A(new_n817), .ZN(new_n818));
  INV_X1    g0618(.A(G303), .ZN(new_n819));
  OAI221_X1 g0619(.A(new_n264), .B1(new_n812), .B2(new_n815), .C1(new_n818), .C2(new_n819), .ZN(new_n820));
  NAND2_X1  g0620(.A1(new_n807), .A2(new_n802), .ZN(new_n821));
  INV_X1    g0621(.A(new_n821), .ZN(new_n822));
  AOI21_X1  g0622(.A(new_n820), .B1(G322), .B2(new_n822), .ZN(new_n823));
  AND2_X1   g0623(.A1(new_n813), .A2(new_n808), .ZN(new_n824));
  OR2_X1    g0624(.A1(new_n824), .A2(KEYINPUT100), .ZN(new_n825));
  NAND2_X1  g0625(.A1(new_n824), .A2(KEYINPUT100), .ZN(new_n826));
  NAND2_X1  g0626(.A1(new_n825), .A2(new_n826), .ZN(new_n827));
  INV_X1    g0627(.A(new_n827), .ZN(new_n828));
  NAND2_X1  g0628(.A1(new_n807), .A2(new_n814), .ZN(new_n829));
  INV_X1    g0629(.A(new_n829), .ZN(new_n830));
  XNOR2_X1  g0630(.A(KEYINPUT33), .B(G317), .ZN(new_n831));
  AOI22_X1  g0631(.A1(new_n828), .A2(G329), .B1(new_n830), .B2(new_n831), .ZN(new_n832));
  NAND3_X1  g0632(.A1(new_n811), .A2(new_n823), .A3(new_n832), .ZN(new_n833));
  OAI22_X1  g0633(.A1(new_n425), .A2(new_n829), .B1(new_n809), .B2(new_n259), .ZN(new_n834));
  INV_X1    g0634(.A(new_n801), .ZN(new_n835));
  INV_X1    g0635(.A(G58), .ZN(new_n836));
  OAI22_X1  g0636(.A1(new_n835), .A2(new_n234), .B1(new_n821), .B2(new_n836), .ZN(new_n837));
  NOR2_X1   g0637(.A1(new_n834), .A2(new_n837), .ZN(new_n838));
  OR3_X1    g0638(.A1(new_n827), .A2(KEYINPUT32), .A3(new_n361), .ZN(new_n839));
  OAI21_X1  g0639(.A(KEYINPUT32), .B1(new_n827), .B2(new_n361), .ZN(new_n840));
  NOR2_X1   g0640(.A1(new_n818), .A2(new_n214), .ZN(new_n841));
  INV_X1    g0641(.A(new_n804), .ZN(new_n842));
  NOR2_X1   g0642(.A1(new_n842), .A2(new_n216), .ZN(new_n843));
  OAI21_X1  g0643(.A(new_n315), .B1(new_n815), .B2(new_n210), .ZN(new_n844));
  NOR3_X1   g0644(.A1(new_n841), .A2(new_n843), .A3(new_n844), .ZN(new_n845));
  NAND4_X1  g0645(.A1(new_n838), .A2(new_n839), .A3(new_n840), .A4(new_n845), .ZN(new_n846));
  AOI21_X1  g0646(.A(new_n794), .B1(new_n833), .B2(new_n846), .ZN(new_n847));
  NOR2_X1   g0647(.A1(G13), .A2(G33), .ZN(new_n848));
  INV_X1    g0648(.A(new_n848), .ZN(new_n849));
  NOR2_X1   g0649(.A1(new_n849), .A2(G20), .ZN(new_n850));
  NOR2_X1   g0650(.A1(new_n793), .A2(new_n850), .ZN(new_n851));
  NAND3_X1  g0651(.A1(new_n228), .A2(G355), .A3(new_n315), .ZN(new_n852));
  NOR2_X1   g0652(.A1(new_n357), .A2(new_n227), .ZN(new_n853));
  OAI21_X1  g0653(.A(new_n853), .B1(new_n237), .B2(G45), .ZN(new_n854));
  INV_X1    g0654(.A(KEYINPUT97), .ZN(new_n855));
  OAI22_X1  g0655(.A1(new_n854), .A2(new_n855), .B1(new_n255), .B2(new_n273), .ZN(new_n856));
  AND2_X1   g0656(.A1(new_n854), .A2(new_n855), .ZN(new_n857));
  OAI221_X1 g0657(.A(new_n852), .B1(G116), .B2(new_n228), .C1(new_n856), .C2(new_n857), .ZN(new_n858));
  AOI211_X1 g0658(.A(new_n789), .B(new_n847), .C1(new_n851), .C2(new_n858), .ZN(new_n859));
  INV_X1    g0659(.A(new_n850), .ZN(new_n860));
  OAI21_X1  g0660(.A(new_n859), .B1(new_n713), .B2(new_n860), .ZN(new_n861));
  AND2_X1   g0661(.A1(new_n788), .A2(new_n861), .ZN(new_n862));
  INV_X1    g0662(.A(new_n862), .ZN(G396));
  OR2_X1    g0663(.A1(new_n329), .A2(new_n708), .ZN(new_n864));
  NAND3_X1  g0664(.A1(new_n334), .A2(new_n337), .A3(new_n864), .ZN(new_n865));
  NAND2_X1  g0665(.A1(new_n865), .A2(KEYINPUT103), .ZN(new_n866));
  OR2_X1    g0666(.A1(new_n334), .A2(new_n864), .ZN(new_n867));
  INV_X1    g0667(.A(KEYINPUT103), .ZN(new_n868));
  NAND4_X1  g0668(.A1(new_n334), .A2(new_n868), .A3(new_n337), .A4(new_n864), .ZN(new_n869));
  NAND3_X1  g0669(.A1(new_n866), .A2(new_n867), .A3(new_n869), .ZN(new_n870));
  XNOR2_X1  g0670(.A(new_n730), .B(new_n870), .ZN(new_n871));
  AOI21_X1  g0671(.A(new_n786), .B1(new_n871), .B2(new_n779), .ZN(new_n872));
  OAI21_X1  g0672(.A(new_n872), .B1(new_n779), .B2(new_n871), .ZN(new_n873));
  NOR2_X1   g0673(.A1(new_n793), .A2(new_n848), .ZN(new_n874));
  AOI21_X1  g0674(.A(new_n789), .B1(new_n874), .B2(new_n259), .ZN(new_n875));
  INV_X1    g0675(.A(new_n809), .ZN(new_n876));
  AOI22_X1  g0676(.A1(new_n876), .A2(G116), .B1(new_n801), .B2(G303), .ZN(new_n877));
  OAI21_X1  g0677(.A(new_n877), .B1(new_n806), .B2(new_n827), .ZN(new_n878));
  INV_X1    g0678(.A(new_n815), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n879), .A2(G87), .ZN(new_n880));
  OAI211_X1 g0680(.A(new_n264), .B(new_n880), .C1(new_n818), .C2(new_n210), .ZN(new_n881));
  OAI22_X1  g0681(.A1(new_n812), .A2(new_n829), .B1(new_n821), .B2(new_n753), .ZN(new_n882));
  NOR4_X1   g0682(.A1(new_n878), .A2(new_n843), .A3(new_n881), .A4(new_n882), .ZN(new_n883));
  XNOR2_X1  g0683(.A(new_n883), .B(KEYINPUT102), .ZN(new_n884));
  AOI22_X1  g0684(.A1(new_n830), .A2(G150), .B1(new_n801), .B2(G137), .ZN(new_n885));
  INV_X1    g0685(.A(G143), .ZN(new_n886));
  OAI221_X1 g0686(.A(new_n885), .B1(new_n886), .B2(new_n821), .C1(new_n361), .C2(new_n809), .ZN(new_n887));
  INV_X1    g0687(.A(KEYINPUT34), .ZN(new_n888));
  OR2_X1    g0688(.A1(new_n887), .A2(new_n888), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n887), .A2(new_n888), .ZN(new_n890));
  AOI22_X1  g0690(.A1(new_n817), .A2(G50), .B1(new_n879), .B2(G68), .ZN(new_n891));
  OAI211_X1 g0691(.A(new_n891), .B(new_n357), .C1(new_n836), .C2(new_n842), .ZN(new_n892));
  AOI21_X1  g0692(.A(new_n892), .B1(G132), .B2(new_n828), .ZN(new_n893));
  AND2_X1   g0693(.A1(new_n890), .A2(new_n893), .ZN(new_n894));
  AOI21_X1  g0694(.A(new_n884), .B1(new_n889), .B2(new_n894), .ZN(new_n895));
  OAI221_X1 g0695(.A(new_n875), .B1(new_n870), .B2(new_n849), .C1(new_n895), .C2(new_n794), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n873), .A2(new_n896), .ZN(G384));
  AOI211_X1 g0697(.A(new_n473), .B(new_n233), .C1(new_n595), .C2(KEYINPUT35), .ZN(new_n898));
  OAI21_X1  g0698(.A(new_n898), .B1(KEYINPUT35), .B2(new_n595), .ZN(new_n899));
  XNOR2_X1  g0699(.A(new_n899), .B(KEYINPUT36), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n368), .A2(G77), .ZN(new_n901));
  INV_X1    g0701(.A(new_n201), .ZN(new_n902));
  OAI22_X1  g0702(.A1(new_n237), .A2(new_n901), .B1(new_n425), .B2(new_n902), .ZN(new_n903));
  NAND3_X1  g0703(.A1(new_n903), .A2(G1), .A3(new_n226), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n900), .A2(new_n904), .ZN(new_n905));
  XOR2_X1   g0705(.A(new_n905), .B(KEYINPUT104), .Z(new_n906));
  NAND3_X1  g0706(.A1(new_n359), .A2(new_n365), .A3(new_n370), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n907), .A2(new_n373), .ZN(new_n908));
  AOI21_X1  g0708(.A(new_n347), .B1(new_n372), .B2(new_n908), .ZN(new_n909));
  OAI21_X1  g0709(.A(new_n417), .B1(new_n909), .B2(new_n705), .ZN(new_n910));
  NOR2_X1   g0710(.A1(new_n909), .A2(new_n400), .ZN(new_n911));
  OAI21_X1  g0711(.A(KEYINPUT37), .B1(new_n910), .B2(new_n911), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n404), .A2(new_n406), .ZN(new_n913));
  INV_X1    g0713(.A(new_n705), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n404), .A2(new_n914), .ZN(new_n915));
  INV_X1    g0715(.A(KEYINPUT37), .ZN(new_n916));
  NAND4_X1  g0716(.A1(new_n913), .A2(new_n915), .A3(new_n916), .A4(new_n417), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n912), .A2(new_n917), .ZN(new_n918));
  NOR2_X1   g0718(.A1(new_n909), .A2(new_n705), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n421), .A2(new_n919), .ZN(new_n920));
  NAND3_X1  g0720(.A1(new_n918), .A2(new_n920), .A3(KEYINPUT38), .ZN(new_n921));
  INV_X1    g0721(.A(KEYINPUT39), .ZN(new_n922));
  OAI21_X1  g0722(.A(new_n417), .B1(new_n384), .B2(new_n400), .ZN(new_n923));
  NOR2_X1   g0723(.A1(new_n384), .A2(new_n705), .ZN(new_n924));
  OAI21_X1  g0724(.A(KEYINPUT37), .B1(new_n923), .B2(new_n924), .ZN(new_n925));
  AOI22_X1  g0725(.A1(new_n917), .A2(new_n925), .B1(new_n421), .B2(new_n924), .ZN(new_n926));
  OAI211_X1 g0726(.A(new_n921), .B(new_n922), .C1(KEYINPUT38), .C2(new_n926), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n927), .A2(KEYINPUT106), .ZN(new_n928));
  AND3_X1   g0728(.A1(new_n918), .A2(new_n920), .A3(KEYINPUT38), .ZN(new_n929));
  AOI21_X1  g0729(.A(KEYINPUT38), .B1(new_n918), .B2(new_n920), .ZN(new_n930));
  OAI21_X1  g0730(.A(KEYINPUT39), .B1(new_n929), .B2(new_n930), .ZN(new_n931));
  INV_X1    g0731(.A(KEYINPUT38), .ZN(new_n932));
  AND2_X1   g0732(.A1(new_n925), .A2(new_n917), .ZN(new_n933));
  AOI21_X1  g0733(.A(new_n915), .B1(new_n676), .B2(new_n681), .ZN(new_n934));
  OAI21_X1  g0734(.A(new_n932), .B1(new_n933), .B2(new_n934), .ZN(new_n935));
  INV_X1    g0735(.A(KEYINPUT106), .ZN(new_n936));
  NAND4_X1  g0736(.A1(new_n935), .A2(new_n936), .A3(new_n922), .A4(new_n921), .ZN(new_n937));
  NAND3_X1  g0737(.A1(new_n928), .A2(new_n931), .A3(new_n937), .ZN(new_n938));
  INV_X1    g0738(.A(new_n460), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n939), .A2(new_n708), .ZN(new_n940));
  INV_X1    g0740(.A(new_n940), .ZN(new_n941));
  NAND2_X1  g0741(.A1(new_n938), .A2(new_n941), .ZN(new_n942));
  INV_X1    g0742(.A(KEYINPUT107), .ZN(new_n943));
  NOR2_X1   g0743(.A1(new_n676), .A2(new_n914), .ZN(new_n944));
  NOR2_X1   g0744(.A1(new_n334), .A2(new_n707), .ZN(new_n945));
  AOI21_X1  g0745(.A(new_n945), .B1(new_n730), .B2(new_n870), .ZN(new_n946));
  NAND3_X1  g0746(.A1(new_n436), .A2(new_n433), .A3(new_n707), .ZN(new_n947));
  NAND3_X1  g0747(.A1(new_n460), .A2(new_n463), .A3(new_n947), .ZN(new_n948));
  INV_X1    g0748(.A(KEYINPUT105), .ZN(new_n949));
  NAND2_X1  g0749(.A1(new_n454), .A2(G169), .ZN(new_n950));
  NAND2_X1  g0750(.A1(new_n950), .A2(KEYINPUT14), .ZN(new_n951));
  NAND4_X1  g0751(.A1(new_n463), .A2(new_n951), .A3(new_n457), .A4(new_n456), .ZN(new_n952));
  AND3_X1   g0752(.A1(new_n436), .A2(new_n433), .A3(new_n707), .ZN(new_n953));
  AOI21_X1  g0753(.A(new_n949), .B1(new_n952), .B2(new_n953), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n948), .A2(new_n954), .ZN(new_n955));
  NAND3_X1  g0755(.A1(new_n952), .A2(new_n953), .A3(new_n949), .ZN(new_n956));
  NAND2_X1  g0756(.A1(new_n955), .A2(new_n956), .ZN(new_n957));
  NOR2_X1   g0757(.A1(new_n946), .A2(new_n957), .ZN(new_n958));
  NOR2_X1   g0758(.A1(new_n929), .A2(new_n930), .ZN(new_n959));
  INV_X1    g0759(.A(new_n959), .ZN(new_n960));
  AOI21_X1  g0760(.A(new_n944), .B1(new_n958), .B2(new_n960), .ZN(new_n961));
  AND3_X1   g0761(.A1(new_n942), .A2(new_n943), .A3(new_n961), .ZN(new_n962));
  AOI21_X1  g0762(.A(new_n943), .B1(new_n942), .B2(new_n961), .ZN(new_n963));
  NOR2_X1   g0763(.A1(new_n962), .A2(new_n963), .ZN(new_n964));
  OAI21_X1  g0764(.A(new_n466), .B1(new_n732), .B2(new_n747), .ZN(new_n965));
  NAND2_X1  g0765(.A1(new_n965), .A2(new_n685), .ZN(new_n966));
  XNOR2_X1  g0766(.A(new_n964), .B(new_n966), .ZN(new_n967));
  INV_X1    g0767(.A(new_n870), .ZN(new_n968));
  NOR2_X1   g0768(.A1(new_n957), .A2(new_n968), .ZN(new_n969));
  NAND2_X1  g0769(.A1(new_n773), .A2(KEYINPUT94), .ZN(new_n970));
  NAND3_X1  g0770(.A1(new_n759), .A2(new_n760), .A3(new_n761), .ZN(new_n971));
  NAND3_X1  g0771(.A1(new_n970), .A2(new_n772), .A3(new_n971), .ZN(new_n972));
  NAND3_X1  g0772(.A1(new_n972), .A2(KEYINPUT31), .A3(new_n707), .ZN(new_n973));
  NAND4_X1  g0773(.A1(new_n769), .A2(new_n771), .A3(new_n777), .A4(new_n973), .ZN(new_n974));
  AND2_X1   g0774(.A1(new_n969), .A2(new_n974), .ZN(new_n975));
  OAI21_X1  g0775(.A(new_n921), .B1(new_n926), .B2(KEYINPUT38), .ZN(new_n976));
  NAND3_X1  g0776(.A1(new_n975), .A2(KEYINPUT40), .A3(new_n976), .ZN(new_n977));
  INV_X1    g0777(.A(KEYINPUT40), .ZN(new_n978));
  NAND2_X1  g0778(.A1(new_n969), .A2(new_n974), .ZN(new_n979));
  OAI21_X1  g0779(.A(new_n978), .B1(new_n979), .B2(new_n959), .ZN(new_n980));
  NAND2_X1  g0780(.A1(new_n977), .A2(new_n980), .ZN(new_n981));
  NAND2_X1  g0781(.A1(new_n466), .A2(new_n974), .ZN(new_n982));
  OR2_X1    g0782(.A1(new_n981), .A2(new_n982), .ZN(new_n983));
  NAND2_X1  g0783(.A1(new_n981), .A2(new_n982), .ZN(new_n984));
  NAND3_X1  g0784(.A1(new_n983), .A2(new_n714), .A3(new_n984), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n967), .A2(new_n985), .ZN(new_n986));
  OAI21_X1  g0786(.A(new_n986), .B1(new_n206), .B2(new_n783), .ZN(new_n987));
  NOR2_X1   g0787(.A1(new_n967), .A2(new_n985), .ZN(new_n988));
  OAI21_X1  g0788(.A(new_n906), .B1(new_n987), .B2(new_n988), .ZN(G367));
  NAND2_X1  g0789(.A1(new_n719), .A2(new_n720), .ZN(new_n990));
  OAI211_X1 g0790(.A(new_n690), .B(new_n600), .C1(new_n608), .C2(new_n708), .ZN(new_n991));
  NAND2_X1  g0791(.A1(new_n693), .A2(new_n707), .ZN(new_n992));
  NAND2_X1  g0792(.A1(new_n991), .A2(new_n992), .ZN(new_n993));
  INV_X1    g0793(.A(new_n993), .ZN(new_n994));
  NOR2_X1   g0794(.A1(new_n990), .A2(new_n994), .ZN(new_n995));
  XNOR2_X1  g0795(.A(new_n995), .B(KEYINPUT42), .ZN(new_n996));
  OAI21_X1  g0796(.A(new_n690), .B1(new_n991), .B2(new_n554), .ZN(new_n997));
  NAND2_X1  g0797(.A1(new_n997), .A2(new_n708), .ZN(new_n998));
  NAND2_X1  g0798(.A1(new_n996), .A2(new_n998), .ZN(new_n999));
  OAI21_X1  g0799(.A(new_n741), .B1(new_n738), .B2(new_n708), .ZN(new_n1000));
  OR3_X1    g0800(.A1(new_n669), .A2(new_n738), .A3(new_n708), .ZN(new_n1001));
  NAND2_X1  g0801(.A1(new_n1000), .A2(new_n1001), .ZN(new_n1002));
  NOR3_X1   g0802(.A1(new_n999), .A2(KEYINPUT43), .A3(new_n1002), .ZN(new_n1003));
  XNOR2_X1  g0803(.A(new_n1003), .B(KEYINPUT108), .ZN(new_n1004));
  XOR2_X1   g0804(.A(new_n1002), .B(KEYINPUT43), .Z(new_n1005));
  NAND2_X1  g0805(.A1(new_n999), .A2(new_n1005), .ZN(new_n1006));
  NAND2_X1  g0806(.A1(new_n1004), .A2(new_n1006), .ZN(new_n1007));
  OAI21_X1  g0807(.A(new_n1007), .B1(new_n718), .B2(new_n994), .ZN(new_n1008));
  INV_X1    g0808(.A(new_n718), .ZN(new_n1009));
  NAND4_X1  g0809(.A1(new_n1004), .A2(new_n1009), .A3(new_n993), .A4(new_n1006), .ZN(new_n1010));
  NAND2_X1  g0810(.A1(new_n1008), .A2(new_n1010), .ZN(new_n1011));
  XOR2_X1   g0811(.A(new_n724), .B(KEYINPUT41), .Z(new_n1012));
  INV_X1    g0812(.A(new_n1012), .ZN(new_n1013));
  OAI21_X1  g0813(.A(new_n990), .B1(new_n717), .B2(new_n719), .ZN(new_n1014));
  XOR2_X1   g0814(.A(new_n715), .B(new_n1014), .Z(new_n1015));
  NOR2_X1   g0815(.A1(new_n780), .A2(new_n1015), .ZN(new_n1016));
  INV_X1    g0816(.A(new_n1016), .ZN(new_n1017));
  NOR2_X1   g0817(.A1(new_n722), .A2(new_n993), .ZN(new_n1018));
  XOR2_X1   g0818(.A(new_n1018), .B(KEYINPUT109), .Z(new_n1019));
  INV_X1    g0819(.A(KEYINPUT44), .ZN(new_n1020));
  OR2_X1    g0820(.A1(new_n1019), .A2(new_n1020), .ZN(new_n1021));
  NAND2_X1  g0821(.A1(new_n1019), .A2(new_n1020), .ZN(new_n1022));
  NAND2_X1  g0822(.A1(new_n722), .A2(new_n993), .ZN(new_n1023));
  XNOR2_X1  g0823(.A(new_n1023), .B(KEYINPUT45), .ZN(new_n1024));
  INV_X1    g0824(.A(KEYINPUT110), .ZN(new_n1025));
  AOI21_X1  g0825(.A(new_n1024), .B1(new_n1025), .B2(new_n1009), .ZN(new_n1026));
  NAND3_X1  g0826(.A1(new_n1021), .A2(new_n1022), .A3(new_n1026), .ZN(new_n1027));
  NOR2_X1   g0827(.A1(new_n1009), .A2(new_n1025), .ZN(new_n1028));
  OR2_X1    g0828(.A1(new_n1027), .A2(new_n1028), .ZN(new_n1029));
  NAND2_X1  g0829(.A1(new_n1027), .A2(new_n1028), .ZN(new_n1030));
  AOI21_X1  g0830(.A(new_n1017), .B1(new_n1029), .B2(new_n1030), .ZN(new_n1031));
  OAI21_X1  g0831(.A(new_n1013), .B1(new_n1031), .B2(new_n780), .ZN(new_n1032));
  AOI21_X1  g0832(.A(new_n1011), .B1(new_n1032), .B2(new_n784), .ZN(new_n1033));
  INV_X1    g0833(.A(new_n1033), .ZN(new_n1034));
  INV_X1    g0834(.A(new_n324), .ZN(new_n1035));
  INV_X1    g0835(.A(new_n853), .ZN(new_n1036));
  OAI221_X1 g0836(.A(new_n851), .B1(new_n228), .B2(new_n1035), .C1(new_n248), .C2(new_n1036), .ZN(new_n1037));
  INV_X1    g0837(.A(KEYINPUT111), .ZN(new_n1038));
  AOI21_X1  g0838(.A(new_n789), .B1(new_n1037), .B2(new_n1038), .ZN(new_n1039));
  OAI21_X1  g0839(.A(new_n1039), .B1(new_n1038), .B2(new_n1037), .ZN(new_n1040));
  AOI22_X1  g0840(.A1(new_n828), .A2(G137), .B1(new_n801), .B2(G143), .ZN(new_n1041));
  OAI21_X1  g0841(.A(new_n1041), .B1(new_n201), .B2(new_n809), .ZN(new_n1042));
  AOI21_X1  g0842(.A(new_n264), .B1(new_n879), .B2(G77), .ZN(new_n1043));
  OAI221_X1 g0843(.A(new_n1043), .B1(new_n842), .B2(new_n425), .C1(new_n836), .C2(new_n818), .ZN(new_n1044));
  INV_X1    g0844(.A(G150), .ZN(new_n1045));
  OAI22_X1  g0845(.A1(new_n1045), .A2(new_n821), .B1(new_n829), .B2(new_n361), .ZN(new_n1046));
  NOR3_X1   g0846(.A1(new_n1042), .A2(new_n1044), .A3(new_n1046), .ZN(new_n1047));
  INV_X1    g0847(.A(G317), .ZN(new_n1048));
  OAI22_X1  g0848(.A1(new_n827), .A2(new_n1048), .B1(new_n829), .B2(new_n753), .ZN(new_n1049));
  INV_X1    g0849(.A(KEYINPUT46), .ZN(new_n1050));
  OAI21_X1  g0850(.A(new_n1050), .B1(new_n818), .B2(new_n473), .ZN(new_n1051));
  NAND3_X1  g0851(.A1(new_n817), .A2(KEYINPUT46), .A3(G116), .ZN(new_n1052));
  OAI211_X1 g0852(.A(new_n1051), .B(new_n1052), .C1(new_n210), .C2(new_n842), .ZN(new_n1053));
  NAND2_X1  g0853(.A1(new_n879), .A2(G97), .ZN(new_n1054));
  OAI211_X1 g0854(.A(new_n350), .B(new_n1054), .C1(new_n835), .C2(new_n806), .ZN(new_n1055));
  OAI22_X1  g0855(.A1(new_n812), .A2(new_n809), .B1(new_n821), .B2(new_n819), .ZN(new_n1056));
  NOR4_X1   g0856(.A1(new_n1049), .A2(new_n1053), .A3(new_n1055), .A4(new_n1056), .ZN(new_n1057));
  NOR2_X1   g0857(.A1(new_n1047), .A2(new_n1057), .ZN(new_n1058));
  XOR2_X1   g0858(.A(new_n1058), .B(KEYINPUT47), .Z(new_n1059));
  AOI21_X1  g0859(.A(new_n1040), .B1(new_n1059), .B2(new_n793), .ZN(new_n1060));
  NAND3_X1  g0860(.A1(new_n1000), .A2(new_n1001), .A3(new_n850), .ZN(new_n1061));
  NAND2_X1  g0861(.A1(new_n1060), .A2(new_n1061), .ZN(new_n1062));
  NAND2_X1  g0862(.A1(new_n1034), .A2(new_n1062), .ZN(G387));
  INV_X1    g0863(.A(new_n1015), .ZN(new_n1064));
  OR2_X1    g0864(.A1(new_n717), .A2(new_n860), .ZN(new_n1065));
  INV_X1    g0865(.A(new_n726), .ZN(new_n1066));
  NAND3_X1  g0866(.A1(new_n1066), .A2(new_n228), .A3(new_n315), .ZN(new_n1067));
  OAI21_X1  g0867(.A(new_n1067), .B1(G107), .B2(new_n228), .ZN(new_n1068));
  NOR2_X1   g0868(.A1(new_n326), .A2(G50), .ZN(new_n1069));
  XNOR2_X1  g0869(.A(KEYINPUT112), .B(KEYINPUT50), .ZN(new_n1070));
  XNOR2_X1  g0870(.A(new_n1069), .B(new_n1070), .ZN(new_n1071));
  AOI211_X1 g0871(.A(G45), .B(new_n1066), .C1(G68), .C2(G77), .ZN(new_n1072));
  AOI21_X1  g0872(.A(new_n1036), .B1(new_n1071), .B2(new_n1072), .ZN(new_n1073));
  NAND2_X1  g0873(.A1(new_n244), .A2(G45), .ZN(new_n1074));
  AOI21_X1  g0874(.A(new_n1068), .B1(new_n1073), .B2(new_n1074), .ZN(new_n1075));
  INV_X1    g0875(.A(new_n851), .ZN(new_n1076));
  OAI21_X1  g0876(.A(new_n786), .B1(new_n1075), .B2(new_n1076), .ZN(new_n1077));
  OAI22_X1  g0877(.A1(new_n835), .A2(new_n361), .B1(new_n821), .B2(new_n234), .ZN(new_n1078));
  AOI21_X1  g0878(.A(new_n1078), .B1(G68), .B2(new_n876), .ZN(new_n1079));
  NAND2_X1  g0879(.A1(new_n817), .A2(G77), .ZN(new_n1080));
  NAND2_X1  g0880(.A1(new_n804), .A2(new_n324), .ZN(new_n1081));
  AND4_X1   g0881(.A1(new_n357), .A2(new_n1080), .A3(new_n1054), .A4(new_n1081), .ZN(new_n1082));
  AOI22_X1  g0882(.A1(new_n828), .A2(G150), .B1(new_n830), .B2(new_n292), .ZN(new_n1083));
  NAND3_X1  g0883(.A1(new_n1079), .A2(new_n1082), .A3(new_n1083), .ZN(new_n1084));
  OAI22_X1  g0884(.A1(new_n818), .A2(new_n753), .B1(new_n842), .B2(new_n812), .ZN(new_n1085));
  AOI22_X1  g0885(.A1(new_n830), .A2(G311), .B1(new_n801), .B2(G322), .ZN(new_n1086));
  OAI221_X1 g0886(.A(new_n1086), .B1(new_n819), .B2(new_n809), .C1(new_n1048), .C2(new_n821), .ZN(new_n1087));
  INV_X1    g0887(.A(KEYINPUT48), .ZN(new_n1088));
  AOI21_X1  g0888(.A(new_n1085), .B1(new_n1087), .B2(new_n1088), .ZN(new_n1089));
  OAI21_X1  g0889(.A(new_n1089), .B1(new_n1088), .B2(new_n1087), .ZN(new_n1090));
  INV_X1    g0890(.A(KEYINPUT49), .ZN(new_n1091));
  AND2_X1   g0891(.A1(new_n1090), .A2(new_n1091), .ZN(new_n1092));
  OAI21_X1  g0892(.A(new_n350), .B1(new_n473), .B2(new_n815), .ZN(new_n1093));
  AOI21_X1  g0893(.A(new_n1093), .B1(new_n828), .B2(G326), .ZN(new_n1094));
  OAI21_X1  g0894(.A(new_n1094), .B1(new_n1090), .B2(new_n1091), .ZN(new_n1095));
  OAI21_X1  g0895(.A(new_n1084), .B1(new_n1092), .B2(new_n1095), .ZN(new_n1096));
  AOI21_X1  g0896(.A(new_n1077), .B1(new_n1096), .B2(new_n793), .ZN(new_n1097));
  AOI22_X1  g0897(.A1(new_n1064), .A2(new_n785), .B1(new_n1065), .B2(new_n1097), .ZN(new_n1098));
  NAND3_X1  g0898(.A1(new_n1017), .A2(KEYINPUT113), .A3(new_n724), .ZN(new_n1099));
  OAI21_X1  g0899(.A(new_n1099), .B1(new_n781), .B2(new_n1064), .ZN(new_n1100));
  AOI21_X1  g0900(.A(KEYINPUT113), .B1(new_n1017), .B2(new_n724), .ZN(new_n1101));
  OAI21_X1  g0901(.A(new_n1098), .B1(new_n1100), .B2(new_n1101), .ZN(G393));
  NAND2_X1  g0902(.A1(new_n1029), .A2(new_n1030), .ZN(new_n1103));
  NAND2_X1  g0903(.A1(new_n1103), .A2(new_n1016), .ZN(new_n1104));
  NAND3_X1  g0904(.A1(new_n1029), .A2(new_n1017), .A3(new_n1030), .ZN(new_n1105));
  NAND3_X1  g0905(.A1(new_n1104), .A2(new_n724), .A3(new_n1105), .ZN(new_n1106));
  NAND2_X1  g0906(.A1(new_n994), .A2(new_n850), .ZN(new_n1107));
  AOI22_X1  g0907(.A1(new_n822), .A2(G159), .B1(new_n801), .B2(G150), .ZN(new_n1108));
  XNOR2_X1  g0908(.A(new_n1108), .B(KEYINPUT51), .ZN(new_n1109));
  NAND2_X1  g0909(.A1(new_n817), .A2(new_n220), .ZN(new_n1110));
  NAND2_X1  g0910(.A1(new_n804), .A2(G77), .ZN(new_n1111));
  NAND4_X1  g0911(.A1(new_n1110), .A2(new_n1111), .A3(new_n880), .A4(new_n357), .ZN(new_n1112));
  NOR2_X1   g0912(.A1(new_n827), .A2(new_n886), .ZN(new_n1113));
  OAI22_X1  g0913(.A1(new_n201), .A2(new_n829), .B1(new_n809), .B2(new_n326), .ZN(new_n1114));
  OR4_X1    g0914(.A1(new_n1109), .A2(new_n1112), .A3(new_n1113), .A4(new_n1114), .ZN(new_n1115));
  OAI22_X1  g0915(.A1(new_n835), .A2(new_n1048), .B1(new_n821), .B2(new_n806), .ZN(new_n1116));
  XNOR2_X1  g0916(.A(KEYINPUT114), .B(KEYINPUT52), .ZN(new_n1117));
  XNOR2_X1  g0917(.A(new_n1116), .B(new_n1117), .ZN(new_n1118));
  OAI221_X1 g0918(.A(new_n264), .B1(new_n210), .B2(new_n815), .C1(new_n818), .C2(new_n812), .ZN(new_n1119));
  AOI21_X1  g0919(.A(new_n1119), .B1(G116), .B2(new_n804), .ZN(new_n1120));
  NAND2_X1  g0920(.A1(new_n876), .A2(G294), .ZN(new_n1121));
  AOI22_X1  g0921(.A1(new_n828), .A2(G322), .B1(new_n830), .B2(G303), .ZN(new_n1122));
  NAND4_X1  g0922(.A1(new_n1118), .A2(new_n1120), .A3(new_n1121), .A4(new_n1122), .ZN(new_n1123));
  AOI21_X1  g0923(.A(new_n794), .B1(new_n1115), .B2(new_n1123), .ZN(new_n1124));
  NOR2_X1   g0924(.A1(new_n252), .A2(new_n1036), .ZN(new_n1125));
  AOI211_X1 g0925(.A(new_n1076), .B(new_n1125), .C1(G97), .C2(new_n227), .ZN(new_n1126));
  NOR3_X1   g0926(.A1(new_n1124), .A2(new_n789), .A3(new_n1126), .ZN(new_n1127));
  AOI22_X1  g0927(.A1(new_n1103), .A2(new_n785), .B1(new_n1107), .B2(new_n1127), .ZN(new_n1128));
  NAND2_X1  g0928(.A1(new_n1106), .A2(new_n1128), .ZN(G390));
  OAI21_X1  g0929(.A(new_n940), .B1(new_n946), .B2(new_n957), .ZN(new_n1130));
  NAND4_X1  g0930(.A1(new_n1130), .A2(new_n928), .A3(new_n931), .A4(new_n937), .ZN(new_n1131));
  AOI21_X1  g0931(.A(new_n941), .B1(new_n935), .B2(new_n921), .ZN(new_n1132));
  NAND3_X1  g0932(.A1(new_n746), .A2(new_n708), .A3(new_n870), .ZN(new_n1133));
  INV_X1    g0933(.A(new_n945), .ZN(new_n1134));
  AND2_X1   g0934(.A1(new_n1133), .A2(new_n1134), .ZN(new_n1135));
  NAND2_X1  g0935(.A1(new_n957), .A2(KEYINPUT115), .ZN(new_n1136));
  INV_X1    g0936(.A(KEYINPUT115), .ZN(new_n1137));
  NAND3_X1  g0937(.A1(new_n955), .A2(new_n1137), .A3(new_n956), .ZN(new_n1138));
  NAND2_X1  g0938(.A1(new_n1136), .A2(new_n1138), .ZN(new_n1139));
  OAI21_X1  g0939(.A(new_n1132), .B1(new_n1135), .B2(new_n1139), .ZN(new_n1140));
  AND2_X1   g0940(.A1(new_n955), .A2(new_n956), .ZN(new_n1141));
  NAND4_X1  g0941(.A1(new_n778), .A2(new_n714), .A3(new_n870), .A4(new_n1141), .ZN(new_n1142));
  AND3_X1   g0942(.A1(new_n1131), .A2(new_n1140), .A3(new_n1142), .ZN(new_n1143));
  NAND3_X1  g0943(.A1(new_n969), .A2(new_n974), .A3(G330), .ZN(new_n1144));
  AOI21_X1  g0944(.A(new_n1144), .B1(new_n1131), .B2(new_n1140), .ZN(new_n1145));
  NOR2_X1   g0945(.A1(new_n1143), .A2(new_n1145), .ZN(new_n1146));
  AND2_X1   g0946(.A1(new_n937), .A2(new_n931), .ZN(new_n1147));
  NAND3_X1  g0947(.A1(new_n1147), .A2(new_n848), .A3(new_n928), .ZN(new_n1148));
  INV_X1    g0948(.A(new_n874), .ZN(new_n1149));
  OAI21_X1  g0949(.A(new_n786), .B1(new_n1149), .B2(new_n292), .ZN(new_n1150));
  AOI211_X1 g0950(.A(new_n315), .B(new_n841), .C1(G68), .C2(new_n879), .ZN(new_n1151));
  AOI22_X1  g0951(.A1(G107), .A2(new_n830), .B1(new_n822), .B2(G116), .ZN(new_n1152));
  NAND3_X1  g0952(.A1(new_n1151), .A2(new_n1111), .A3(new_n1152), .ZN(new_n1153));
  AOI22_X1  g0953(.A1(new_n876), .A2(G97), .B1(new_n801), .B2(G283), .ZN(new_n1154));
  OAI21_X1  g0954(.A(new_n1154), .B1(new_n753), .B2(new_n827), .ZN(new_n1155));
  NAND2_X1  g0955(.A1(new_n801), .A2(G128), .ZN(new_n1156));
  INV_X1    g0956(.A(G132), .ZN(new_n1157));
  INV_X1    g0957(.A(G137), .ZN(new_n1158));
  OAI221_X1 g0958(.A(new_n1156), .B1(new_n821), .B2(new_n1157), .C1(new_n1158), .C2(new_n829), .ZN(new_n1159));
  NAND2_X1  g0959(.A1(new_n817), .A2(G150), .ZN(new_n1160));
  XOR2_X1   g0960(.A(new_n1160), .B(KEYINPUT53), .Z(new_n1161));
  NAND2_X1  g0961(.A1(new_n828), .A2(G125), .ZN(new_n1162));
  XOR2_X1   g0962(.A(KEYINPUT54), .B(G143), .Z(new_n1163));
  XNOR2_X1  g0963(.A(new_n1163), .B(KEYINPUT117), .ZN(new_n1164));
  NAND2_X1  g0964(.A1(new_n876), .A2(new_n1164), .ZN(new_n1165));
  OAI21_X1  g0965(.A(new_n315), .B1(new_n815), .B2(new_n201), .ZN(new_n1166));
  AOI21_X1  g0966(.A(new_n1166), .B1(G159), .B2(new_n804), .ZN(new_n1167));
  NAND4_X1  g0967(.A1(new_n1161), .A2(new_n1162), .A3(new_n1165), .A4(new_n1167), .ZN(new_n1168));
  OAI22_X1  g0968(.A1(new_n1153), .A2(new_n1155), .B1(new_n1159), .B2(new_n1168), .ZN(new_n1169));
  AOI21_X1  g0969(.A(new_n1150), .B1(new_n1169), .B2(new_n793), .ZN(new_n1170));
  AOI22_X1  g0970(.A1(new_n1146), .A2(new_n785), .B1(new_n1148), .B2(new_n1170), .ZN(new_n1171));
  NAND2_X1  g0971(.A1(new_n1131), .A2(new_n1140), .ZN(new_n1172));
  INV_X1    g0972(.A(new_n1144), .ZN(new_n1173));
  NAND2_X1  g0973(.A1(new_n1172), .A2(new_n1173), .ZN(new_n1174));
  NAND3_X1  g0974(.A1(new_n1131), .A2(new_n1140), .A3(new_n1142), .ZN(new_n1175));
  NAND2_X1  g0975(.A1(new_n1174), .A2(new_n1175), .ZN(new_n1176));
  NAND3_X1  g0976(.A1(new_n466), .A2(G330), .A3(new_n974), .ZN(new_n1177));
  AND3_X1   g0977(.A1(new_n965), .A2(new_n685), .A3(new_n1177), .ZN(new_n1178));
  NAND3_X1  g0978(.A1(new_n974), .A2(G330), .A3(new_n870), .ZN(new_n1179));
  AND2_X1   g0979(.A1(new_n1179), .A2(new_n1139), .ZN(new_n1180));
  NAND2_X1  g0980(.A1(new_n1135), .A2(new_n1142), .ZN(new_n1181));
  NOR2_X1   g0981(.A1(new_n1180), .A2(new_n1181), .ZN(new_n1182));
  NAND3_X1  g0982(.A1(new_n778), .A2(new_n714), .A3(new_n870), .ZN(new_n1183));
  NAND2_X1  g0983(.A1(new_n1183), .A2(new_n957), .ZN(new_n1184));
  AOI21_X1  g0984(.A(new_n946), .B1(new_n1184), .B2(new_n1144), .ZN(new_n1185));
  OAI21_X1  g0985(.A(new_n1178), .B1(new_n1182), .B2(new_n1185), .ZN(new_n1186));
  AOI21_X1  g0986(.A(new_n725), .B1(new_n1176), .B2(new_n1186), .ZN(new_n1187));
  NAND2_X1  g0987(.A1(new_n1179), .A2(new_n1139), .ZN(new_n1188));
  NAND3_X1  g0988(.A1(new_n1188), .A2(new_n1135), .A3(new_n1142), .ZN(new_n1189));
  NAND2_X1  g0989(.A1(new_n974), .A2(G330), .ZN(new_n1190));
  INV_X1    g0990(.A(new_n1190), .ZN(new_n1191));
  AOI22_X1  g0991(.A1(new_n1191), .A2(new_n969), .B1(new_n1183), .B2(new_n957), .ZN(new_n1192));
  OAI21_X1  g0992(.A(new_n1189), .B1(new_n1192), .B2(new_n946), .ZN(new_n1193));
  NAND4_X1  g0993(.A1(new_n1174), .A2(new_n1175), .A3(new_n1178), .A4(new_n1193), .ZN(new_n1194));
  AOI21_X1  g0994(.A(KEYINPUT116), .B1(new_n1187), .B2(new_n1194), .ZN(new_n1195));
  OAI21_X1  g0995(.A(new_n1186), .B1(new_n1143), .B2(new_n1145), .ZN(new_n1196));
  AND4_X1   g0996(.A1(KEYINPUT116), .A2(new_n1196), .A3(new_n1194), .A4(new_n724), .ZN(new_n1197));
  OAI21_X1  g0997(.A(new_n1171), .B1(new_n1195), .B2(new_n1197), .ZN(G378));
  NAND2_X1  g0998(.A1(new_n311), .A2(new_n344), .ZN(new_n1199));
  AND2_X1   g0999(.A1(new_n305), .A2(new_n914), .ZN(new_n1200));
  OR2_X1    g1000(.A1(new_n1199), .A2(new_n1200), .ZN(new_n1201));
  NAND2_X1  g1001(.A1(new_n1199), .A2(new_n1200), .ZN(new_n1202));
  NAND2_X1  g1002(.A1(new_n1201), .A2(new_n1202), .ZN(new_n1203));
  XNOR2_X1  g1003(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1204));
  INV_X1    g1004(.A(new_n1204), .ZN(new_n1205));
  NAND2_X1  g1005(.A1(new_n1203), .A2(new_n1205), .ZN(new_n1206));
  NAND3_X1  g1006(.A1(new_n1201), .A2(new_n1202), .A3(new_n1204), .ZN(new_n1207));
  AND2_X1   g1007(.A1(new_n1206), .A2(new_n1207), .ZN(new_n1208));
  AOI21_X1  g1008(.A(KEYINPUT40), .B1(new_n975), .B2(new_n960), .ZN(new_n1209));
  NAND2_X1  g1009(.A1(new_n976), .A2(KEYINPUT40), .ZN(new_n1210));
  OAI21_X1  g1010(.A(G330), .B1(new_n979), .B2(new_n1210), .ZN(new_n1211));
  OAI21_X1  g1011(.A(new_n1208), .B1(new_n1209), .B2(new_n1211), .ZN(new_n1212));
  NAND2_X1  g1012(.A1(new_n1206), .A2(new_n1207), .ZN(new_n1213));
  NAND4_X1  g1013(.A1(new_n977), .A2(new_n1213), .A3(new_n980), .A4(G330), .ZN(new_n1214));
  NAND2_X1  g1014(.A1(new_n1212), .A2(new_n1214), .ZN(new_n1215));
  OAI21_X1  g1015(.A(new_n1215), .B1(new_n962), .B2(new_n963), .ZN(new_n1216));
  AOI21_X1  g1016(.A(new_n940), .B1(new_n1147), .B2(new_n928), .ZN(new_n1217));
  INV_X1    g1017(.A(new_n961), .ZN(new_n1218));
  OAI21_X1  g1018(.A(KEYINPUT107), .B1(new_n1217), .B2(new_n1218), .ZN(new_n1219));
  NAND3_X1  g1019(.A1(new_n942), .A2(new_n943), .A3(new_n961), .ZN(new_n1220));
  NAND4_X1  g1020(.A1(new_n1219), .A2(new_n1220), .A3(new_n1214), .A4(new_n1212), .ZN(new_n1221));
  NAND3_X1  g1021(.A1(new_n1216), .A2(new_n1221), .A3(new_n785), .ZN(new_n1222));
  OAI21_X1  g1022(.A(new_n786), .B1(new_n1149), .B2(new_n902), .ZN(new_n1223));
  AOI22_X1  g1023(.A1(new_n830), .A2(G97), .B1(new_n801), .B2(G116), .ZN(new_n1224));
  OAI21_X1  g1024(.A(new_n1224), .B1(new_n812), .B2(new_n827), .ZN(new_n1225));
  NAND3_X1  g1025(.A1(new_n1080), .A2(new_n272), .A3(new_n350), .ZN(new_n1226));
  XNOR2_X1  g1026(.A(new_n1226), .B(KEYINPUT119), .ZN(new_n1227));
  NOR2_X1   g1027(.A1(new_n815), .A2(new_n836), .ZN(new_n1228));
  XNOR2_X1  g1028(.A(new_n1228), .B(KEYINPUT118), .ZN(new_n1229));
  OAI21_X1  g1029(.A(new_n1229), .B1(new_n1035), .B2(new_n809), .ZN(new_n1230));
  OAI22_X1  g1030(.A1(new_n821), .A2(new_n210), .B1(new_n425), .B2(new_n842), .ZN(new_n1231));
  NOR4_X1   g1031(.A1(new_n1225), .A2(new_n1227), .A3(new_n1230), .A4(new_n1231), .ZN(new_n1232));
  NAND2_X1  g1032(.A1(new_n350), .A2(new_n272), .ZN(new_n1233));
  AOI21_X1  g1033(.A(G50), .B1(new_n260), .B2(new_n272), .ZN(new_n1234));
  AOI22_X1  g1034(.A1(new_n1232), .A2(KEYINPUT58), .B1(new_n1233), .B2(new_n1234), .ZN(new_n1235));
  AOI22_X1  g1035(.A1(new_n822), .A2(G128), .B1(new_n1164), .B2(new_n817), .ZN(new_n1236));
  AOI22_X1  g1036(.A1(new_n876), .A2(G137), .B1(G150), .B2(new_n804), .ZN(new_n1237));
  AOI22_X1  g1037(.A1(new_n830), .A2(G132), .B1(new_n801), .B2(G125), .ZN(new_n1238));
  NAND3_X1  g1038(.A1(new_n1236), .A2(new_n1237), .A3(new_n1238), .ZN(new_n1239));
  NOR2_X1   g1039(.A1(new_n1239), .A2(KEYINPUT59), .ZN(new_n1240));
  NAND2_X1  g1040(.A1(new_n1239), .A2(KEYINPUT59), .ZN(new_n1241));
  AOI211_X1 g1041(.A(G33), .B(G41), .C1(new_n879), .C2(G159), .ZN(new_n1242));
  XNOR2_X1  g1042(.A(KEYINPUT120), .B(G124), .ZN(new_n1243));
  OAI211_X1 g1043(.A(new_n1241), .B(new_n1242), .C1(new_n827), .C2(new_n1243), .ZN(new_n1244));
  OAI221_X1 g1044(.A(new_n1235), .B1(KEYINPUT58), .B2(new_n1232), .C1(new_n1240), .C2(new_n1244), .ZN(new_n1245));
  AOI21_X1  g1045(.A(new_n1223), .B1(new_n1245), .B2(new_n793), .ZN(new_n1246));
  OAI21_X1  g1046(.A(new_n1246), .B1(new_n1213), .B2(new_n849), .ZN(new_n1247));
  AND3_X1   g1047(.A1(new_n1222), .A2(KEYINPUT121), .A3(new_n1247), .ZN(new_n1248));
  AOI21_X1  g1048(.A(KEYINPUT121), .B1(new_n1222), .B2(new_n1247), .ZN(new_n1249));
  OR2_X1    g1049(.A1(new_n1248), .A2(new_n1249), .ZN(new_n1250));
  INV_X1    g1050(.A(KEYINPUT57), .ZN(new_n1251));
  NAND2_X1  g1051(.A1(new_n1216), .A2(new_n1221), .ZN(new_n1252));
  NAND3_X1  g1052(.A1(new_n965), .A2(new_n685), .A3(new_n1177), .ZN(new_n1253));
  AOI21_X1  g1053(.A(new_n1253), .B1(new_n1146), .B2(new_n1193), .ZN(new_n1254));
  OAI21_X1  g1054(.A(new_n1251), .B1(new_n1252), .B2(new_n1254), .ZN(new_n1255));
  NAND2_X1  g1055(.A1(new_n1194), .A2(new_n1178), .ZN(new_n1256));
  NAND4_X1  g1056(.A1(new_n1256), .A2(KEYINPUT57), .A3(new_n1221), .A4(new_n1216), .ZN(new_n1257));
  NAND3_X1  g1057(.A1(new_n1255), .A2(new_n724), .A3(new_n1257), .ZN(new_n1258));
  NAND2_X1  g1058(.A1(new_n1250), .A2(new_n1258), .ZN(G375));
  INV_X1    g1059(.A(KEYINPUT122), .ZN(new_n1260));
  NAND2_X1  g1060(.A1(new_n1184), .A2(new_n1144), .ZN(new_n1261));
  INV_X1    g1061(.A(new_n946), .ZN(new_n1262));
  NAND2_X1  g1062(.A1(new_n1261), .A2(new_n1262), .ZN(new_n1263));
  AOI21_X1  g1063(.A(new_n784), .B1(new_n1263), .B2(new_n1189), .ZN(new_n1264));
  AOI21_X1  g1064(.A(new_n849), .B1(new_n1136), .B2(new_n1138), .ZN(new_n1265));
  OAI21_X1  g1065(.A(new_n357), .B1(new_n818), .B2(new_n361), .ZN(new_n1266));
  OAI21_X1  g1066(.A(new_n1229), .B1(new_n1157), .B2(new_n835), .ZN(new_n1267));
  AOI211_X1 g1067(.A(new_n1266), .B(new_n1267), .C1(G50), .C2(new_n804), .ZN(new_n1268));
  OAI22_X1  g1068(.A1(new_n1158), .A2(new_n821), .B1(new_n809), .B2(new_n1045), .ZN(new_n1269));
  AND2_X1   g1069(.A1(new_n830), .A2(new_n1164), .ZN(new_n1270));
  AOI211_X1 g1070(.A(new_n1269), .B(new_n1270), .C1(G128), .C2(new_n828), .ZN(new_n1271));
  OAI22_X1  g1071(.A1(new_n827), .A2(new_n819), .B1(new_n809), .B2(new_n210), .ZN(new_n1272));
  AOI21_X1  g1072(.A(new_n1272), .B1(G283), .B2(new_n822), .ZN(new_n1273));
  OAI22_X1  g1073(.A1(new_n835), .A2(new_n753), .B1(new_n829), .B2(new_n473), .ZN(new_n1274));
  AOI21_X1  g1074(.A(new_n315), .B1(new_n879), .B2(G77), .ZN(new_n1275));
  OAI211_X1 g1075(.A(new_n1275), .B(new_n1081), .C1(new_n216), .C2(new_n818), .ZN(new_n1276));
  NOR2_X1   g1076(.A1(new_n1274), .A2(new_n1276), .ZN(new_n1277));
  AOI22_X1  g1077(.A1(new_n1268), .A2(new_n1271), .B1(new_n1273), .B2(new_n1277), .ZN(new_n1278));
  OAI221_X1 g1078(.A(new_n786), .B1(G68), .B2(new_n1149), .C1(new_n1278), .C2(new_n794), .ZN(new_n1279));
  NOR2_X1   g1079(.A1(new_n1265), .A2(new_n1279), .ZN(new_n1280));
  OAI21_X1  g1080(.A(new_n1260), .B1(new_n1264), .B2(new_n1280), .ZN(new_n1281));
  NAND2_X1  g1081(.A1(new_n1193), .A2(new_n785), .ZN(new_n1282));
  INV_X1    g1082(.A(new_n1280), .ZN(new_n1283));
  NAND3_X1  g1083(.A1(new_n1282), .A2(KEYINPUT122), .A3(new_n1283), .ZN(new_n1284));
  NAND2_X1  g1084(.A1(new_n1281), .A2(new_n1284), .ZN(new_n1285));
  NAND3_X1  g1085(.A1(new_n1263), .A2(new_n1253), .A3(new_n1189), .ZN(new_n1286));
  NAND3_X1  g1086(.A1(new_n1186), .A2(new_n1286), .A3(new_n1013), .ZN(new_n1287));
  NAND2_X1  g1087(.A1(new_n1285), .A2(new_n1287), .ZN(G381));
  NOR2_X1   g1088(.A1(G390), .A2(G384), .ZN(new_n1289));
  NAND3_X1  g1089(.A1(new_n1289), .A2(new_n1034), .A3(new_n1062), .ZN(new_n1290));
  OR2_X1    g1090(.A1(G393), .A2(G396), .ZN(new_n1291));
  NOR3_X1   g1091(.A1(new_n1290), .A2(G381), .A3(new_n1291), .ZN(new_n1292));
  INV_X1    g1092(.A(G375), .ZN(new_n1293));
  NAND2_X1  g1093(.A1(new_n1187), .A2(new_n1194), .ZN(new_n1294));
  AND2_X1   g1094(.A1(new_n1294), .A2(new_n1171), .ZN(new_n1295));
  NAND3_X1  g1095(.A1(new_n1292), .A2(new_n1293), .A3(new_n1295), .ZN(new_n1296));
  AND2_X1   g1096(.A1(new_n1296), .A2(KEYINPUT123), .ZN(new_n1297));
  NOR2_X1   g1097(.A1(new_n1296), .A2(KEYINPUT123), .ZN(new_n1298));
  OR2_X1    g1098(.A1(new_n1297), .A2(new_n1298), .ZN(G407));
  AND2_X1   g1099(.A1(new_n1295), .A2(new_n706), .ZN(new_n1300));
  NAND2_X1  g1100(.A1(new_n1293), .A2(new_n1300), .ZN(new_n1301));
  OAI211_X1 g1101(.A(G213), .B(new_n1301), .C1(new_n1297), .C2(new_n1298), .ZN(G409));
  OAI211_X1 g1102(.A(new_n1258), .B(G378), .C1(new_n1249), .C2(new_n1248), .ZN(new_n1303));
  AND2_X1   g1103(.A1(new_n1216), .A2(new_n1221), .ZN(new_n1304));
  NAND4_X1  g1104(.A1(new_n1304), .A2(KEYINPUT124), .A3(new_n1013), .A4(new_n1256), .ZN(new_n1305));
  AND2_X1   g1105(.A1(new_n1222), .A2(new_n1247), .ZN(new_n1306));
  INV_X1    g1106(.A(KEYINPUT124), .ZN(new_n1307));
  NAND3_X1  g1107(.A1(new_n1216), .A2(new_n1221), .A3(new_n1013), .ZN(new_n1308));
  OAI21_X1  g1108(.A(new_n1307), .B1(new_n1308), .B2(new_n1254), .ZN(new_n1309));
  NAND3_X1  g1109(.A1(new_n1305), .A2(new_n1306), .A3(new_n1309), .ZN(new_n1310));
  NAND2_X1  g1110(.A1(new_n1310), .A2(new_n1295), .ZN(new_n1311));
  NAND2_X1  g1111(.A1(new_n1303), .A2(new_n1311), .ZN(new_n1312));
  NAND2_X1  g1112(.A1(new_n706), .A2(G213), .ZN(new_n1313));
  INV_X1    g1113(.A(KEYINPUT60), .ZN(new_n1314));
  NAND2_X1  g1114(.A1(new_n1286), .A2(new_n1314), .ZN(new_n1315));
  NAND4_X1  g1115(.A1(new_n1263), .A2(KEYINPUT60), .A3(new_n1253), .A4(new_n1189), .ZN(new_n1316));
  NAND4_X1  g1116(.A1(new_n1315), .A2(new_n1316), .A3(new_n724), .A4(new_n1186), .ZN(new_n1317));
  AOI21_X1  g1117(.A(G384), .B1(new_n1285), .B2(new_n1317), .ZN(new_n1318));
  INV_X1    g1118(.A(new_n1318), .ZN(new_n1319));
  NAND3_X1  g1119(.A1(new_n1285), .A2(G384), .A3(new_n1317), .ZN(new_n1320));
  NAND2_X1  g1120(.A1(new_n1319), .A2(new_n1320), .ZN(new_n1321));
  INV_X1    g1121(.A(new_n1321), .ZN(new_n1322));
  NAND3_X1  g1122(.A1(new_n1312), .A2(new_n1313), .A3(new_n1322), .ZN(new_n1323));
  NAND2_X1  g1123(.A1(new_n1323), .A2(KEYINPUT62), .ZN(new_n1324));
  NAND2_X1  g1124(.A1(new_n1312), .A2(new_n1313), .ZN(new_n1325));
  INV_X1    g1125(.A(KEYINPUT125), .ZN(new_n1326));
  AND3_X1   g1126(.A1(new_n706), .A2(G213), .A3(G2897), .ZN(new_n1327));
  INV_X1    g1127(.A(new_n1320), .ZN(new_n1328));
  OAI211_X1 g1128(.A(new_n1326), .B(new_n1327), .C1(new_n1328), .C2(new_n1318), .ZN(new_n1329));
  NAND3_X1  g1129(.A1(new_n1319), .A2(KEYINPUT125), .A3(new_n1320), .ZN(new_n1330));
  NAND2_X1  g1130(.A1(new_n1329), .A2(new_n1330), .ZN(new_n1331));
  AOI21_X1  g1131(.A(new_n1327), .B1(new_n1321), .B2(new_n1326), .ZN(new_n1332));
  NOR2_X1   g1132(.A1(new_n1331), .A2(new_n1332), .ZN(new_n1333));
  NAND2_X1  g1133(.A1(new_n1325), .A2(new_n1333), .ZN(new_n1334));
  INV_X1    g1134(.A(KEYINPUT61), .ZN(new_n1335));
  INV_X1    g1135(.A(KEYINPUT62), .ZN(new_n1336));
  NAND4_X1  g1136(.A1(new_n1312), .A2(new_n1336), .A3(new_n1313), .A4(new_n1322), .ZN(new_n1337));
  NAND4_X1  g1137(.A1(new_n1324), .A2(new_n1334), .A3(new_n1335), .A4(new_n1337), .ZN(new_n1338));
  NAND2_X1  g1138(.A1(new_n1338), .A2(KEYINPUT127), .ZN(new_n1339));
  XNOR2_X1  g1139(.A(G393), .B(new_n862), .ZN(new_n1340));
  INV_X1    g1140(.A(new_n1340), .ZN(new_n1341));
  NAND3_X1  g1141(.A1(new_n1034), .A2(new_n1062), .A3(G390), .ZN(new_n1342));
  INV_X1    g1142(.A(new_n1062), .ZN(new_n1343));
  OAI211_X1 g1143(.A(new_n1106), .B(new_n1128), .C1(new_n1033), .C2(new_n1343), .ZN(new_n1344));
  NAND2_X1  g1144(.A1(new_n1342), .A2(new_n1344), .ZN(new_n1345));
  AOI21_X1  g1145(.A(new_n1341), .B1(new_n1345), .B2(KEYINPUT126), .ZN(new_n1346));
  INV_X1    g1146(.A(new_n1346), .ZN(new_n1347));
  NAND3_X1  g1147(.A1(new_n1345), .A2(KEYINPUT126), .A3(new_n1341), .ZN(new_n1348));
  NAND2_X1  g1148(.A1(new_n1347), .A2(new_n1348), .ZN(new_n1349));
  AOI21_X1  g1149(.A(KEYINPUT61), .B1(new_n1325), .B2(new_n1333), .ZN(new_n1350));
  INV_X1    g1150(.A(KEYINPUT127), .ZN(new_n1351));
  NAND4_X1  g1151(.A1(new_n1350), .A2(new_n1324), .A3(new_n1351), .A4(new_n1337), .ZN(new_n1352));
  NAND3_X1  g1152(.A1(new_n1339), .A2(new_n1349), .A3(new_n1352), .ZN(new_n1353));
  AND3_X1   g1153(.A1(new_n1345), .A2(KEYINPUT126), .A3(new_n1341), .ZN(new_n1354));
  NOR2_X1   g1154(.A1(new_n1354), .A2(new_n1346), .ZN(new_n1355));
  INV_X1    g1155(.A(new_n1323), .ZN(new_n1356));
  OR2_X1    g1156(.A1(new_n1356), .A2(KEYINPUT63), .ZN(new_n1357));
  NAND2_X1  g1157(.A1(new_n1356), .A2(KEYINPUT63), .ZN(new_n1358));
  NAND4_X1  g1158(.A1(new_n1355), .A2(new_n1357), .A3(new_n1350), .A4(new_n1358), .ZN(new_n1359));
  NAND2_X1  g1159(.A1(new_n1353), .A2(new_n1359), .ZN(G405));
  NAND2_X1  g1160(.A1(G375), .A2(new_n1295), .ZN(new_n1361));
  AND2_X1   g1161(.A1(new_n1361), .A2(new_n1303), .ZN(new_n1362));
  AND2_X1   g1162(.A1(new_n1362), .A2(new_n1321), .ZN(new_n1363));
  NOR2_X1   g1163(.A1(new_n1362), .A2(new_n1321), .ZN(new_n1364));
  OAI21_X1  g1164(.A(new_n1349), .B1(new_n1363), .B2(new_n1364), .ZN(new_n1365));
  NOR2_X1   g1165(.A1(new_n1363), .A2(new_n1364), .ZN(new_n1366));
  NAND2_X1  g1166(.A1(new_n1366), .A2(new_n1355), .ZN(new_n1367));
  NAND2_X1  g1167(.A1(new_n1365), .A2(new_n1367), .ZN(G402));
endmodule


