//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 1 1 1 0 1 1 0 0 1 0 1 1 1 1 1 0 0 0 1 0 0 0 0 0 1 0 1 1 0 0 0 0 0 1 1 0 0 0 0 1 0 1 1 0 0 0 1 0 1 1 0 0 0 1 1 0 0 0 1 0 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:23:59 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n705, new_n706, new_n707, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n730, new_n731, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n744, new_n745, new_n746, new_n747, new_n748, new_n749,
    new_n750, new_n751, new_n752, new_n753, new_n754, new_n755, new_n756,
    new_n757, new_n759, new_n760, new_n761, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n790, new_n791, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n817,
    new_n818, new_n819, new_n820, new_n821, new_n822, new_n823, new_n824,
    new_n825, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n920, new_n921, new_n922, new_n923, new_n924,
    new_n925, new_n926, new_n927, new_n928, new_n929, new_n930, new_n931,
    new_n932, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n944, new_n945, new_n946, new_n948,
    new_n949, new_n950, new_n951, new_n952, new_n953, new_n954, new_n955,
    new_n957, new_n958, new_n959, new_n960, new_n961, new_n962, new_n963,
    new_n964, new_n965, new_n966, new_n967, new_n968, new_n969, new_n970,
    new_n971, new_n972, new_n973, new_n974, new_n975, new_n976, new_n977,
    new_n978, new_n980, new_n981, new_n982, new_n983, new_n984, new_n985,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1017, new_n1018, new_n1019,
    new_n1020, new_n1021, new_n1022, new_n1023, new_n1024, new_n1025;
  OAI21_X1  g000(.A(G214), .B1(G237), .B2(G902), .ZN(new_n187));
  INV_X1    g001(.A(G146), .ZN(new_n188));
  NAND2_X1  g002(.A1(new_n188), .A2(G143), .ZN(new_n189));
  INV_X1    g003(.A(G143), .ZN(new_n190));
  NAND2_X1  g004(.A1(new_n190), .A2(G146), .ZN(new_n191));
  NAND4_X1  g005(.A1(new_n189), .A2(new_n191), .A3(KEYINPUT0), .A4(G128), .ZN(new_n192));
  XNOR2_X1  g006(.A(G143), .B(G146), .ZN(new_n193));
  XNOR2_X1  g007(.A(KEYINPUT0), .B(G128), .ZN(new_n194));
  OAI21_X1  g008(.A(new_n192), .B1(new_n193), .B2(new_n194), .ZN(new_n195));
  INV_X1    g009(.A(new_n195), .ZN(new_n196));
  XNOR2_X1  g010(.A(KEYINPUT67), .B(G125), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n196), .A2(new_n197), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n189), .A2(new_n191), .ZN(new_n199));
  XNOR2_X1  g013(.A(KEYINPUT65), .B(G128), .ZN(new_n200));
  INV_X1    g014(.A(KEYINPUT1), .ZN(new_n201));
  AOI21_X1  g015(.A(new_n201), .B1(G143), .B2(new_n188), .ZN(new_n202));
  OAI21_X1  g016(.A(new_n199), .B1(new_n200), .B2(new_n202), .ZN(new_n203));
  NAND3_X1  g017(.A1(new_n193), .A2(new_n201), .A3(G128), .ZN(new_n204));
  AND2_X1   g018(.A1(new_n203), .A2(new_n204), .ZN(new_n205));
  OAI21_X1  g019(.A(new_n198), .B1(new_n197), .B2(new_n205), .ZN(new_n206));
  XNOR2_X1  g020(.A(KEYINPUT80), .B(G224), .ZN(new_n207));
  INV_X1    g021(.A(G953), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n209), .A2(KEYINPUT7), .ZN(new_n210));
  XNOR2_X1  g024(.A(new_n206), .B(new_n210), .ZN(new_n211));
  INV_X1    g025(.A(G104), .ZN(new_n212));
  OAI21_X1  g026(.A(KEYINPUT75), .B1(new_n212), .B2(G107), .ZN(new_n213));
  INV_X1    g027(.A(KEYINPUT75), .ZN(new_n214));
  INV_X1    g028(.A(G107), .ZN(new_n215));
  NAND3_X1  g029(.A1(new_n214), .A2(new_n215), .A3(G104), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n212), .A2(G107), .ZN(new_n217));
  NAND3_X1  g031(.A1(new_n213), .A2(new_n216), .A3(new_n217), .ZN(new_n218));
  NAND3_X1  g032(.A1(new_n218), .A2(KEYINPUT76), .A3(G101), .ZN(new_n219));
  INV_X1    g033(.A(KEYINPUT73), .ZN(new_n220));
  OAI21_X1  g034(.A(new_n220), .B1(new_n215), .B2(G104), .ZN(new_n221));
  NAND3_X1  g035(.A1(new_n212), .A2(KEYINPUT73), .A3(G107), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  INV_X1    g037(.A(KEYINPUT72), .ZN(new_n224));
  NAND3_X1  g038(.A1(new_n224), .A2(new_n215), .A3(G104), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n225), .A2(KEYINPUT3), .ZN(new_n226));
  INV_X1    g040(.A(G101), .ZN(new_n227));
  INV_X1    g041(.A(KEYINPUT3), .ZN(new_n228));
  NAND4_X1  g042(.A1(new_n224), .A2(new_n228), .A3(new_n215), .A4(G104), .ZN(new_n229));
  NAND4_X1  g043(.A1(new_n223), .A2(new_n226), .A3(new_n227), .A4(new_n229), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n219), .A2(new_n230), .ZN(new_n231));
  AOI21_X1  g045(.A(KEYINPUT76), .B1(new_n218), .B2(G101), .ZN(new_n232));
  NOR2_X1   g046(.A1(new_n231), .A2(new_n232), .ZN(new_n233));
  INV_X1    g047(.A(G116), .ZN(new_n234));
  OR2_X1    g048(.A1(new_n234), .A2(G119), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n234), .A2(G119), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n235), .A2(new_n236), .ZN(new_n237));
  INV_X1    g051(.A(new_n237), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n238), .A2(KEYINPUT5), .ZN(new_n239));
  NOR2_X1   g053(.A1(new_n235), .A2(KEYINPUT5), .ZN(new_n240));
  INV_X1    g054(.A(G113), .ZN(new_n241));
  NOR2_X1   g055(.A1(new_n240), .A2(new_n241), .ZN(new_n242));
  XNOR2_X1  g056(.A(KEYINPUT2), .B(G113), .ZN(new_n243));
  INV_X1    g057(.A(new_n243), .ZN(new_n244));
  AOI22_X1  g058(.A1(new_n239), .A2(new_n242), .B1(new_n238), .B2(new_n244), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n233), .A2(new_n245), .ZN(new_n246));
  XNOR2_X1  g060(.A(G110), .B(G122), .ZN(new_n247));
  NAND3_X1  g061(.A1(new_n223), .A2(new_n226), .A3(new_n229), .ZN(new_n248));
  INV_X1    g062(.A(KEYINPUT74), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n248), .A2(new_n249), .ZN(new_n250));
  INV_X1    g064(.A(KEYINPUT4), .ZN(new_n251));
  NAND4_X1  g065(.A1(new_n223), .A2(new_n226), .A3(KEYINPUT74), .A4(new_n229), .ZN(new_n252));
  NAND4_X1  g066(.A1(new_n250), .A2(new_n251), .A3(G101), .A4(new_n252), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n238), .A2(new_n244), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n237), .A2(new_n243), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n254), .A2(new_n255), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n253), .A2(new_n256), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n230), .A2(KEYINPUT4), .ZN(new_n258));
  AOI21_X1  g072(.A(new_n227), .B1(new_n248), .B2(new_n249), .ZN(new_n259));
  AOI21_X1  g073(.A(new_n258), .B1(new_n259), .B2(new_n252), .ZN(new_n260));
  OAI211_X1 g074(.A(new_n246), .B(new_n247), .C1(new_n257), .C2(new_n260), .ZN(new_n261));
  XOR2_X1   g075(.A(new_n233), .B(new_n245), .Z(new_n262));
  XOR2_X1   g076(.A(new_n247), .B(KEYINPUT8), .Z(new_n263));
  OAI211_X1 g077(.A(new_n211), .B(new_n261), .C1(new_n262), .C2(new_n263), .ZN(new_n264));
  INV_X1    g078(.A(G902), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n264), .A2(new_n265), .ZN(new_n266));
  OAI21_X1  g080(.A(G210), .B1(G237), .B2(G902), .ZN(new_n267));
  XNOR2_X1  g081(.A(new_n267), .B(KEYINPUT81), .ZN(new_n268));
  OAI21_X1  g082(.A(new_n246), .B1(new_n257), .B2(new_n260), .ZN(new_n269));
  INV_X1    g083(.A(KEYINPUT78), .ZN(new_n270));
  NAND2_X1  g084(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  OAI211_X1 g085(.A(new_n246), .B(KEYINPUT78), .C1(new_n257), .C2(new_n260), .ZN(new_n272));
  NOR2_X1   g086(.A1(new_n247), .A2(KEYINPUT6), .ZN(new_n273));
  NAND3_X1  g087(.A1(new_n271), .A2(new_n272), .A3(new_n273), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n274), .A2(KEYINPUT79), .ZN(new_n275));
  INV_X1    g089(.A(KEYINPUT79), .ZN(new_n276));
  NAND4_X1  g090(.A1(new_n271), .A2(new_n276), .A3(new_n272), .A4(new_n273), .ZN(new_n277));
  INV_X1    g091(.A(new_n247), .ZN(new_n278));
  NAND3_X1  g092(.A1(new_n271), .A2(new_n272), .A3(new_n278), .ZN(new_n279));
  AND2_X1   g093(.A1(new_n261), .A2(KEYINPUT6), .ZN(new_n280));
  AOI22_X1  g094(.A1(new_n275), .A2(new_n277), .B1(new_n279), .B2(new_n280), .ZN(new_n281));
  XNOR2_X1  g095(.A(new_n206), .B(new_n209), .ZN(new_n282));
  AOI211_X1 g096(.A(new_n266), .B(new_n268), .C1(new_n281), .C2(new_n282), .ZN(new_n283));
  INV_X1    g097(.A(new_n268), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n275), .A2(new_n277), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n279), .A2(new_n280), .ZN(new_n286));
  NAND3_X1  g100(.A1(new_n285), .A2(new_n282), .A3(new_n286), .ZN(new_n287));
  INV_X1    g101(.A(new_n266), .ZN(new_n288));
  AOI21_X1  g102(.A(new_n284), .B1(new_n287), .B2(new_n288), .ZN(new_n289));
  OAI21_X1  g103(.A(new_n187), .B1(new_n283), .B2(new_n289), .ZN(new_n290));
  XNOR2_X1  g104(.A(G110), .B(G140), .ZN(new_n291));
  AND2_X1   g105(.A1(new_n208), .A2(G227), .ZN(new_n292));
  XNOR2_X1  g106(.A(new_n291), .B(new_n292), .ZN(new_n293));
  INV_X1    g107(.A(KEYINPUT77), .ZN(new_n294));
  OAI21_X1  g108(.A(new_n205), .B1(new_n231), .B2(new_n232), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n218), .A2(G101), .ZN(new_n296));
  INV_X1    g110(.A(KEYINPUT76), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n296), .A2(new_n297), .ZN(new_n298));
  INV_X1    g112(.A(G128), .ZN(new_n299));
  OAI21_X1  g113(.A(new_n199), .B1(new_n202), .B2(new_n299), .ZN(new_n300));
  NAND2_X1  g114(.A1(new_n300), .A2(new_n204), .ZN(new_n301));
  NAND4_X1  g115(.A1(new_n298), .A2(new_n301), .A3(new_n230), .A4(new_n219), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n295), .A2(new_n302), .ZN(new_n303));
  INV_X1    g117(.A(KEYINPUT11), .ZN(new_n304));
  INV_X1    g118(.A(G134), .ZN(new_n305));
  OAI21_X1  g119(.A(new_n304), .B1(new_n305), .B2(G137), .ZN(new_n306));
  INV_X1    g120(.A(G137), .ZN(new_n307));
  NAND3_X1  g121(.A1(new_n307), .A2(KEYINPUT11), .A3(G134), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n305), .A2(G137), .ZN(new_n309));
  NAND3_X1  g123(.A1(new_n306), .A2(new_n308), .A3(new_n309), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n310), .A2(G131), .ZN(new_n311));
  INV_X1    g125(.A(G131), .ZN(new_n312));
  NAND4_X1  g126(.A1(new_n306), .A2(new_n308), .A3(new_n312), .A4(new_n309), .ZN(new_n313));
  NAND2_X1  g127(.A1(new_n311), .A2(new_n313), .ZN(new_n314));
  AOI21_X1  g128(.A(KEYINPUT12), .B1(new_n303), .B2(new_n314), .ZN(new_n315));
  INV_X1    g129(.A(KEYINPUT12), .ZN(new_n316));
  INV_X1    g130(.A(new_n314), .ZN(new_n317));
  AOI211_X1 g131(.A(new_n316), .B(new_n317), .C1(new_n295), .C2(new_n302), .ZN(new_n318));
  OR2_X1    g132(.A1(new_n315), .A2(new_n318), .ZN(new_n319));
  NAND3_X1  g133(.A1(new_n250), .A2(G101), .A3(new_n252), .ZN(new_n320));
  INV_X1    g134(.A(new_n258), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n320), .A2(new_n321), .ZN(new_n322));
  NAND3_X1  g136(.A1(new_n322), .A2(new_n196), .A3(new_n253), .ZN(new_n323));
  INV_X1    g137(.A(KEYINPUT10), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n302), .A2(new_n324), .ZN(new_n325));
  NOR2_X1   g139(.A1(new_n205), .A2(new_n324), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n233), .A2(new_n326), .ZN(new_n327));
  NAND4_X1  g141(.A1(new_n323), .A2(new_n317), .A3(new_n325), .A4(new_n327), .ZN(new_n328));
  AOI21_X1  g142(.A(new_n294), .B1(new_n319), .B2(new_n328), .ZN(new_n329));
  OAI211_X1 g143(.A(new_n328), .B(new_n294), .C1(new_n318), .C2(new_n315), .ZN(new_n330));
  INV_X1    g144(.A(new_n330), .ZN(new_n331));
  OAI21_X1  g145(.A(new_n293), .B1(new_n329), .B2(new_n331), .ZN(new_n332));
  INV_X1    g146(.A(new_n293), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n328), .A2(new_n333), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n253), .A2(new_n196), .ZN(new_n335));
  OAI211_X1 g149(.A(new_n327), .B(new_n325), .C1(new_n335), .C2(new_n260), .ZN(new_n336));
  AOI21_X1  g150(.A(new_n334), .B1(new_n314), .B2(new_n336), .ZN(new_n337));
  INV_X1    g151(.A(new_n337), .ZN(new_n338));
  NAND3_X1  g152(.A1(new_n332), .A2(G469), .A3(new_n338), .ZN(new_n339));
  INV_X1    g153(.A(G469), .ZN(new_n340));
  NOR2_X1   g154(.A1(new_n340), .A2(new_n265), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n336), .A2(new_n314), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n342), .A2(new_n328), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n343), .A2(new_n293), .ZN(new_n344));
  OAI211_X1 g158(.A(new_n328), .B(new_n333), .C1(new_n318), .C2(new_n315), .ZN(new_n345));
  AOI21_X1  g159(.A(G902), .B1(new_n344), .B2(new_n345), .ZN(new_n346));
  AOI21_X1  g160(.A(new_n341), .B1(new_n346), .B2(new_n340), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n339), .A2(new_n347), .ZN(new_n348));
  INV_X1    g162(.A(G221), .ZN(new_n349));
  XNOR2_X1  g163(.A(KEYINPUT9), .B(G234), .ZN(new_n350));
  INV_X1    g164(.A(new_n350), .ZN(new_n351));
  AOI21_X1  g165(.A(new_n349), .B1(new_n351), .B2(new_n265), .ZN(new_n352));
  INV_X1    g166(.A(new_n352), .ZN(new_n353));
  NOR2_X1   g167(.A1(new_n234), .A2(G122), .ZN(new_n354));
  INV_X1    g168(.A(KEYINPUT14), .ZN(new_n355));
  OAI21_X1  g169(.A(G107), .B1(new_n354), .B2(new_n355), .ZN(new_n356));
  XNOR2_X1  g170(.A(G116), .B(G122), .ZN(new_n357));
  XOR2_X1   g171(.A(new_n356), .B(new_n357), .Z(new_n358));
  NAND2_X1  g172(.A1(new_n190), .A2(G128), .ZN(new_n359));
  INV_X1    g173(.A(new_n359), .ZN(new_n360));
  AOI21_X1  g174(.A(new_n360), .B1(new_n200), .B2(G143), .ZN(new_n361));
  NOR2_X1   g175(.A1(new_n361), .A2(new_n305), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n299), .A2(KEYINPUT65), .ZN(new_n363));
  INV_X1    g177(.A(KEYINPUT65), .ZN(new_n364));
  NAND2_X1  g178(.A1(new_n364), .A2(G128), .ZN(new_n365));
  NAND3_X1  g179(.A1(new_n363), .A2(new_n365), .A3(G143), .ZN(new_n366));
  NAND3_X1  g180(.A1(new_n366), .A2(new_n305), .A3(new_n359), .ZN(new_n367));
  INV_X1    g181(.A(new_n367), .ZN(new_n368));
  OAI21_X1  g182(.A(new_n358), .B1(new_n362), .B2(new_n368), .ZN(new_n369));
  INV_X1    g183(.A(G217), .ZN(new_n370));
  NOR3_X1   g184(.A1(new_n350), .A2(new_n370), .A3(G953), .ZN(new_n371));
  INV_X1    g185(.A(KEYINPUT13), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n372), .A2(KEYINPUT85), .ZN(new_n373));
  INV_X1    g187(.A(KEYINPUT85), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n374), .A2(KEYINPUT13), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n373), .A2(new_n375), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n376), .A2(new_n360), .ZN(new_n377));
  NAND3_X1  g191(.A1(new_n359), .A2(new_n373), .A3(new_n375), .ZN(new_n378));
  NAND3_X1  g192(.A1(new_n377), .A2(new_n378), .A3(new_n366), .ZN(new_n379));
  NAND2_X1  g193(.A1(new_n379), .A2(G134), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n357), .A2(new_n215), .ZN(new_n381));
  INV_X1    g195(.A(G122), .ZN(new_n382));
  NOR2_X1   g196(.A1(new_n382), .A2(G116), .ZN(new_n383));
  OAI21_X1  g197(.A(G107), .B1(new_n354), .B2(new_n383), .ZN(new_n384));
  AOI22_X1  g198(.A1(new_n361), .A2(new_n305), .B1(new_n381), .B2(new_n384), .ZN(new_n385));
  AND3_X1   g199(.A1(new_n380), .A2(KEYINPUT86), .A3(new_n385), .ZN(new_n386));
  AOI21_X1  g200(.A(KEYINPUT86), .B1(new_n380), .B2(new_n385), .ZN(new_n387));
  OAI211_X1 g201(.A(new_n369), .B(new_n371), .C1(new_n386), .C2(new_n387), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n388), .A2(KEYINPUT87), .ZN(new_n389));
  INV_X1    g203(.A(KEYINPUT86), .ZN(new_n390));
  AOI22_X1  g204(.A1(new_n360), .A2(new_n376), .B1(new_n200), .B2(G143), .ZN(new_n391));
  AOI21_X1  g205(.A(new_n305), .B1(new_n391), .B2(new_n378), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n381), .A2(new_n384), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n393), .A2(new_n367), .ZN(new_n394));
  OAI21_X1  g208(.A(new_n390), .B1(new_n392), .B2(new_n394), .ZN(new_n395));
  NAND3_X1  g209(.A1(new_n380), .A2(new_n385), .A3(KEYINPUT86), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n395), .A2(new_n396), .ZN(new_n397));
  INV_X1    g211(.A(KEYINPUT87), .ZN(new_n398));
  NAND4_X1  g212(.A1(new_n397), .A2(new_n398), .A3(new_n369), .A4(new_n371), .ZN(new_n399));
  OAI21_X1  g213(.A(new_n369), .B1(new_n386), .B2(new_n387), .ZN(new_n400));
  INV_X1    g214(.A(new_n371), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n400), .A2(new_n401), .ZN(new_n402));
  NAND3_X1  g216(.A1(new_n389), .A2(new_n399), .A3(new_n402), .ZN(new_n403));
  INV_X1    g217(.A(KEYINPUT88), .ZN(new_n404));
  NAND3_X1  g218(.A1(new_n403), .A2(new_n404), .A3(new_n265), .ZN(new_n405));
  INV_X1    g219(.A(G478), .ZN(new_n406));
  NOR2_X1   g220(.A1(new_n406), .A2(KEYINPUT15), .ZN(new_n407));
  NAND2_X1  g221(.A1(new_n405), .A2(new_n407), .ZN(new_n408));
  INV_X1    g222(.A(new_n407), .ZN(new_n409));
  NAND4_X1  g223(.A1(new_n403), .A2(new_n404), .A3(new_n265), .A4(new_n409), .ZN(new_n410));
  INV_X1    g224(.A(G952), .ZN(new_n411));
  AOI211_X1 g225(.A(G953), .B(new_n411), .C1(G234), .C2(G237), .ZN(new_n412));
  INV_X1    g226(.A(G234), .ZN(new_n413));
  INV_X1    g227(.A(G237), .ZN(new_n414));
  OAI211_X1 g228(.A(G902), .B(G953), .C1(new_n413), .C2(new_n414), .ZN(new_n415));
  XOR2_X1   g229(.A(new_n415), .B(KEYINPUT89), .Z(new_n416));
  INV_X1    g230(.A(new_n416), .ZN(new_n417));
  XNOR2_X1  g231(.A(KEYINPUT21), .B(G898), .ZN(new_n418));
  AOI21_X1  g232(.A(new_n412), .B1(new_n417), .B2(new_n418), .ZN(new_n419));
  INV_X1    g233(.A(new_n419), .ZN(new_n420));
  NAND3_X1  g234(.A1(new_n408), .A2(new_n410), .A3(new_n420), .ZN(new_n421));
  INV_X1    g235(.A(KEYINPUT20), .ZN(new_n422));
  INV_X1    g236(.A(KEYINPUT18), .ZN(new_n423));
  NOR2_X1   g237(.A1(new_n423), .A2(new_n312), .ZN(new_n424));
  NAND3_X1  g238(.A1(new_n414), .A2(new_n208), .A3(G214), .ZN(new_n425));
  NOR2_X1   g239(.A1(new_n425), .A2(new_n190), .ZN(new_n426));
  NOR2_X1   g240(.A1(G237), .A2(G953), .ZN(new_n427));
  AOI21_X1  g241(.A(G143), .B1(new_n427), .B2(G214), .ZN(new_n428));
  OAI21_X1  g242(.A(new_n424), .B1(new_n426), .B2(new_n428), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n425), .A2(new_n190), .ZN(new_n430));
  NAND3_X1  g244(.A1(new_n427), .A2(G143), .A3(G214), .ZN(new_n431));
  OAI211_X1 g245(.A(new_n430), .B(new_n431), .C1(new_n423), .C2(new_n312), .ZN(new_n432));
  OR2_X1    g246(.A1(KEYINPUT67), .A2(G125), .ZN(new_n433));
  NAND2_X1  g247(.A1(KEYINPUT67), .A2(G125), .ZN(new_n434));
  NAND3_X1  g248(.A1(new_n433), .A2(G140), .A3(new_n434), .ZN(new_n435));
  INV_X1    g249(.A(G140), .ZN(new_n436));
  NAND2_X1  g250(.A1(new_n436), .A2(G125), .ZN(new_n437));
  AOI21_X1  g251(.A(new_n188), .B1(new_n435), .B2(new_n437), .ZN(new_n438));
  INV_X1    g252(.A(G125), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n439), .A2(G140), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n437), .A2(new_n440), .ZN(new_n441));
  NOR2_X1   g255(.A1(new_n441), .A2(G146), .ZN(new_n442));
  OAI211_X1 g256(.A(new_n429), .B(new_n432), .C1(new_n438), .C2(new_n442), .ZN(new_n443));
  INV_X1    g257(.A(KEYINPUT82), .ZN(new_n444));
  XNOR2_X1  g258(.A(new_n443), .B(new_n444), .ZN(new_n445));
  XNOR2_X1  g259(.A(G113), .B(G122), .ZN(new_n446));
  XNOR2_X1  g260(.A(new_n446), .B(new_n212), .ZN(new_n447));
  XOR2_X1   g261(.A(new_n447), .B(KEYINPUT83), .Z(new_n448));
  OAI21_X1  g262(.A(G131), .B1(new_n426), .B2(new_n428), .ZN(new_n449));
  INV_X1    g263(.A(KEYINPUT17), .ZN(new_n450));
  NAND3_X1  g264(.A1(new_n430), .A2(new_n312), .A3(new_n431), .ZN(new_n451));
  NAND3_X1  g265(.A1(new_n449), .A2(new_n450), .A3(new_n451), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n452), .A2(KEYINPUT84), .ZN(new_n453));
  INV_X1    g267(.A(KEYINPUT84), .ZN(new_n454));
  NAND4_X1  g268(.A1(new_n449), .A2(new_n454), .A3(new_n450), .A4(new_n451), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n453), .A2(new_n455), .ZN(new_n456));
  INV_X1    g270(.A(new_n449), .ZN(new_n457));
  NAND2_X1  g271(.A1(new_n457), .A2(KEYINPUT17), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n456), .A2(new_n458), .ZN(new_n459));
  NAND3_X1  g273(.A1(new_n435), .A2(KEYINPUT16), .A3(new_n437), .ZN(new_n460));
  NOR2_X1   g274(.A1(KEYINPUT16), .A2(G140), .ZN(new_n461));
  AOI21_X1  g275(.A(new_n188), .B1(new_n197), .B2(new_n461), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n460), .A2(new_n462), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n463), .A2(KEYINPUT68), .ZN(new_n464));
  INV_X1    g278(.A(KEYINPUT68), .ZN(new_n465));
  NAND3_X1  g279(.A1(new_n460), .A2(new_n462), .A3(new_n465), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n464), .A2(new_n466), .ZN(new_n467));
  NAND2_X1  g281(.A1(new_n197), .A2(new_n461), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n460), .A2(new_n468), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n469), .A2(new_n188), .ZN(new_n470));
  NAND2_X1  g284(.A1(new_n470), .A2(KEYINPUT69), .ZN(new_n471));
  AOI21_X1  g285(.A(G146), .B1(new_n460), .B2(new_n468), .ZN(new_n472));
  INV_X1    g286(.A(KEYINPUT69), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n472), .A2(new_n473), .ZN(new_n474));
  NAND3_X1  g288(.A1(new_n467), .A2(new_n471), .A3(new_n474), .ZN(new_n475));
  OAI211_X1 g289(.A(new_n445), .B(new_n448), .C1(new_n459), .C2(new_n475), .ZN(new_n476));
  NAND2_X1  g290(.A1(new_n449), .A2(new_n451), .ZN(new_n477));
  AOI21_X1  g291(.A(KEYINPUT19), .B1(new_n437), .B2(new_n440), .ZN(new_n478));
  AND2_X1   g292(.A1(new_n435), .A2(new_n437), .ZN(new_n479));
  AOI21_X1  g293(.A(new_n478), .B1(new_n479), .B2(KEYINPUT19), .ZN(new_n480));
  OAI211_X1 g294(.A(new_n463), .B(new_n477), .C1(new_n480), .C2(G146), .ZN(new_n481));
  AND2_X1   g295(.A1(new_n443), .A2(new_n444), .ZN(new_n482));
  NOR2_X1   g296(.A1(new_n443), .A2(new_n444), .ZN(new_n483));
  OAI21_X1  g297(.A(new_n481), .B1(new_n482), .B2(new_n483), .ZN(new_n484));
  INV_X1    g298(.A(new_n447), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n484), .A2(new_n485), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n476), .A2(new_n486), .ZN(new_n487));
  NOR2_X1   g301(.A1(G475), .A2(G902), .ZN(new_n488));
  AOI21_X1  g302(.A(new_n422), .B1(new_n487), .B2(new_n488), .ZN(new_n489));
  INV_X1    g303(.A(new_n488), .ZN(new_n490));
  AOI211_X1 g304(.A(KEYINPUT20), .B(new_n490), .C1(new_n476), .C2(new_n486), .ZN(new_n491));
  OAI21_X1  g305(.A(new_n445), .B1(new_n459), .B2(new_n475), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n492), .A2(new_n485), .ZN(new_n493));
  AOI21_X1  g307(.A(G902), .B1(new_n493), .B2(new_n476), .ZN(new_n494));
  INV_X1    g308(.A(G475), .ZN(new_n495));
  OAI22_X1  g309(.A1(new_n489), .A2(new_n491), .B1(new_n494), .B2(new_n495), .ZN(new_n496));
  NOR2_X1   g310(.A1(new_n421), .A2(new_n496), .ZN(new_n497));
  NAND3_X1  g311(.A1(new_n348), .A2(new_n353), .A3(new_n497), .ZN(new_n498));
  NOR2_X1   g312(.A1(new_n290), .A2(new_n498), .ZN(new_n499));
  INV_X1    g313(.A(G472), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n203), .A2(new_n204), .ZN(new_n501));
  OR3_X1    g315(.A1(new_n305), .A2(KEYINPUT64), .A3(G137), .ZN(new_n502));
  INV_X1    g316(.A(new_n309), .ZN(new_n503));
  OAI21_X1  g317(.A(KEYINPUT64), .B1(new_n305), .B2(G137), .ZN(new_n504));
  OAI211_X1 g318(.A(new_n502), .B(G131), .C1(new_n503), .C2(new_n504), .ZN(new_n505));
  AND3_X1   g319(.A1(new_n501), .A2(new_n313), .A3(new_n505), .ZN(new_n506));
  AOI21_X1  g320(.A(new_n195), .B1(new_n311), .B2(new_n313), .ZN(new_n507));
  NOR3_X1   g321(.A1(new_n506), .A2(new_n256), .A3(new_n507), .ZN(new_n508));
  AND2_X1   g322(.A1(new_n254), .A2(new_n255), .ZN(new_n509));
  NAND2_X1  g323(.A1(new_n196), .A2(new_n314), .ZN(new_n510));
  NAND3_X1  g324(.A1(new_n501), .A2(new_n313), .A3(new_n505), .ZN(new_n511));
  AOI21_X1  g325(.A(new_n509), .B1(new_n510), .B2(new_n511), .ZN(new_n512));
  OAI21_X1  g326(.A(KEYINPUT28), .B1(new_n508), .B2(new_n512), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n427), .A2(G210), .ZN(new_n514));
  XNOR2_X1  g328(.A(new_n514), .B(KEYINPUT27), .ZN(new_n515));
  XNOR2_X1  g329(.A(KEYINPUT26), .B(G101), .ZN(new_n516));
  XNOR2_X1  g330(.A(new_n515), .B(new_n516), .ZN(new_n517));
  NAND3_X1  g331(.A1(new_n509), .A2(new_n510), .A3(new_n511), .ZN(new_n518));
  INV_X1    g332(.A(KEYINPUT28), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  NAND3_X1  g334(.A1(new_n513), .A2(new_n517), .A3(new_n520), .ZN(new_n521));
  INV_X1    g335(.A(KEYINPUT29), .ZN(new_n522));
  NOR2_X1   g336(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  NOR2_X1   g337(.A1(new_n523), .A2(G902), .ZN(new_n524));
  INV_X1    g338(.A(KEYINPUT66), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n525), .A2(KEYINPUT30), .ZN(new_n526));
  NOR2_X1   g340(.A1(new_n525), .A2(KEYINPUT30), .ZN(new_n527));
  INV_X1    g341(.A(new_n527), .ZN(new_n528));
  OAI211_X1 g342(.A(new_n526), .B(new_n528), .C1(new_n506), .C2(new_n507), .ZN(new_n529));
  INV_X1    g343(.A(KEYINPUT30), .ZN(new_n530));
  NAND4_X1  g344(.A1(new_n510), .A2(new_n511), .A3(KEYINPUT66), .A4(new_n530), .ZN(new_n531));
  NAND2_X1  g345(.A1(new_n529), .A2(new_n531), .ZN(new_n532));
  AOI21_X1  g346(.A(new_n508), .B1(new_n532), .B2(new_n256), .ZN(new_n533));
  OAI211_X1 g347(.A(new_n521), .B(new_n522), .C1(new_n533), .C2(new_n517), .ZN(new_n534));
  AOI21_X1  g348(.A(new_n500), .B1(new_n524), .B2(new_n534), .ZN(new_n535));
  AOI21_X1  g349(.A(new_n509), .B1(new_n529), .B2(new_n531), .ZN(new_n536));
  INV_X1    g350(.A(new_n517), .ZN(new_n537));
  NOR4_X1   g351(.A1(new_n536), .A2(KEYINPUT31), .A3(new_n508), .A4(new_n537), .ZN(new_n538));
  OAI21_X1  g352(.A(new_n256), .B1(new_n506), .B2(new_n507), .ZN(new_n539));
  AOI21_X1  g353(.A(new_n519), .B1(new_n539), .B2(new_n518), .ZN(new_n540));
  INV_X1    g354(.A(new_n520), .ZN(new_n541));
  OAI21_X1  g355(.A(new_n537), .B1(new_n540), .B2(new_n541), .ZN(new_n542));
  INV_X1    g356(.A(KEYINPUT31), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  NAND2_X1  g358(.A1(new_n533), .A2(new_n517), .ZN(new_n545));
  AOI21_X1  g359(.A(new_n538), .B1(new_n544), .B2(new_n545), .ZN(new_n546));
  NOR2_X1   g360(.A1(G472), .A2(G902), .ZN(new_n547));
  INV_X1    g361(.A(new_n547), .ZN(new_n548));
  OAI21_X1  g362(.A(KEYINPUT32), .B1(new_n546), .B2(new_n548), .ZN(new_n549));
  NOR3_X1   g363(.A1(new_n536), .A2(new_n508), .A3(new_n537), .ZN(new_n550));
  NAND2_X1  g364(.A1(new_n550), .A2(new_n543), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n513), .A2(new_n520), .ZN(new_n552));
  AOI21_X1  g366(.A(KEYINPUT31), .B1(new_n552), .B2(new_n537), .ZN(new_n553));
  OAI21_X1  g367(.A(new_n551), .B1(new_n553), .B2(new_n550), .ZN(new_n554));
  INV_X1    g368(.A(KEYINPUT32), .ZN(new_n555));
  NAND3_X1  g369(.A1(new_n554), .A2(new_n555), .A3(new_n547), .ZN(new_n556));
  AOI21_X1  g370(.A(new_n535), .B1(new_n549), .B2(new_n556), .ZN(new_n557));
  AOI21_X1  g371(.A(new_n370), .B1(G234), .B2(new_n265), .ZN(new_n558));
  INV_X1    g372(.A(new_n558), .ZN(new_n559));
  NAND3_X1  g373(.A1(new_n200), .A2(KEYINPUT23), .A3(G119), .ZN(new_n560));
  AOI21_X1  g374(.A(KEYINPUT23), .B1(new_n299), .B2(G119), .ZN(new_n561));
  NOR2_X1   g375(.A1(new_n299), .A2(G119), .ZN(new_n562));
  NOR2_X1   g376(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n560), .A2(new_n563), .ZN(new_n564));
  AOI21_X1  g378(.A(new_n562), .B1(new_n200), .B2(G119), .ZN(new_n565));
  XOR2_X1   g379(.A(KEYINPUT24), .B(G110), .Z(new_n566));
  OAI22_X1  g380(.A1(new_n564), .A2(G110), .B1(new_n565), .B2(new_n566), .ZN(new_n567));
  INV_X1    g381(.A(new_n442), .ZN(new_n568));
  NAND3_X1  g382(.A1(new_n567), .A2(new_n463), .A3(new_n568), .ZN(new_n569));
  INV_X1    g383(.A(KEYINPUT70), .ZN(new_n570));
  AOI22_X1  g384(.A1(new_n564), .A2(G110), .B1(new_n565), .B2(new_n566), .ZN(new_n571));
  AND3_X1   g385(.A1(new_n460), .A2(new_n462), .A3(new_n465), .ZN(new_n572));
  AOI21_X1  g386(.A(new_n465), .B1(new_n460), .B2(new_n462), .ZN(new_n573));
  OAI22_X1  g387(.A1(new_n572), .A2(new_n573), .B1(new_n472), .B2(new_n473), .ZN(new_n574));
  INV_X1    g388(.A(new_n474), .ZN(new_n575));
  OAI211_X1 g389(.A(new_n570), .B(new_n571), .C1(new_n574), .C2(new_n575), .ZN(new_n576));
  INV_X1    g390(.A(new_n576), .ZN(new_n577));
  AOI21_X1  g391(.A(new_n570), .B1(new_n475), .B2(new_n571), .ZN(new_n578));
  OAI21_X1  g392(.A(new_n569), .B1(new_n577), .B2(new_n578), .ZN(new_n579));
  XNOR2_X1  g393(.A(KEYINPUT22), .B(G137), .ZN(new_n580));
  NOR3_X1   g394(.A1(new_n349), .A2(new_n413), .A3(G953), .ZN(new_n581));
  XOR2_X1   g395(.A(new_n580), .B(new_n581), .Z(new_n582));
  INV_X1    g396(.A(new_n582), .ZN(new_n583));
  NAND2_X1  g397(.A1(new_n579), .A2(new_n583), .ZN(new_n584));
  OAI21_X1  g398(.A(new_n571), .B1(new_n574), .B2(new_n575), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n585), .A2(KEYINPUT70), .ZN(new_n586));
  NAND2_X1  g400(.A1(new_n586), .A2(new_n576), .ZN(new_n587));
  NAND3_X1  g401(.A1(new_n587), .A2(new_n569), .A3(new_n582), .ZN(new_n588));
  NAND3_X1  g402(.A1(new_n584), .A2(new_n265), .A3(new_n588), .ZN(new_n589));
  INV_X1    g403(.A(KEYINPUT25), .ZN(new_n590));
  NAND2_X1  g404(.A1(new_n589), .A2(new_n590), .ZN(new_n591));
  NAND4_X1  g405(.A1(new_n584), .A2(KEYINPUT25), .A3(new_n265), .A4(new_n588), .ZN(new_n592));
  AOI21_X1  g406(.A(new_n559), .B1(new_n591), .B2(new_n592), .ZN(new_n593));
  AOI21_X1  g407(.A(new_n582), .B1(new_n587), .B2(new_n569), .ZN(new_n594));
  INV_X1    g408(.A(new_n569), .ZN(new_n595));
  AOI211_X1 g409(.A(new_n595), .B(new_n583), .C1(new_n586), .C2(new_n576), .ZN(new_n596));
  NOR2_X1   g410(.A1(new_n594), .A2(new_n596), .ZN(new_n597));
  INV_X1    g411(.A(new_n597), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n559), .A2(new_n265), .ZN(new_n599));
  XNOR2_X1  g413(.A(new_n599), .B(KEYINPUT71), .ZN(new_n600));
  NOR2_X1   g414(.A1(new_n598), .A2(new_n600), .ZN(new_n601));
  NOR3_X1   g415(.A1(new_n557), .A2(new_n593), .A3(new_n601), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n499), .A2(new_n602), .ZN(new_n603));
  XNOR2_X1  g417(.A(new_n603), .B(G101), .ZN(G3));
  AOI21_X1  g418(.A(KEYINPUT25), .B1(new_n597), .B2(new_n265), .ZN(new_n605));
  INV_X1    g419(.A(new_n592), .ZN(new_n606));
  OAI21_X1  g420(.A(new_n558), .B1(new_n605), .B2(new_n606), .ZN(new_n607));
  INV_X1    g421(.A(new_n601), .ZN(new_n608));
  AOI22_X1  g422(.A1(new_n542), .A2(new_n543), .B1(new_n533), .B2(new_n517), .ZN(new_n609));
  OAI21_X1  g423(.A(new_n265), .B1(new_n609), .B2(new_n538), .ZN(new_n610));
  AOI22_X1  g424(.A1(new_n610), .A2(G472), .B1(new_n554), .B2(new_n547), .ZN(new_n611));
  NAND3_X1  g425(.A1(new_n607), .A2(new_n608), .A3(new_n611), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n348), .A2(new_n353), .ZN(new_n613));
  OAI21_X1  g427(.A(KEYINPUT90), .B1(new_n612), .B2(new_n613), .ZN(new_n614));
  NOR2_X1   g428(.A1(new_n593), .A2(new_n601), .ZN(new_n615));
  INV_X1    g429(.A(KEYINPUT90), .ZN(new_n616));
  AOI21_X1  g430(.A(new_n352), .B1(new_n339), .B2(new_n347), .ZN(new_n617));
  NAND4_X1  g431(.A1(new_n615), .A2(new_n616), .A3(new_n617), .A4(new_n611), .ZN(new_n618));
  INV_X1    g432(.A(KEYINPUT33), .ZN(new_n619));
  NAND2_X1  g433(.A1(new_n403), .A2(new_n619), .ZN(new_n620));
  NAND3_X1  g434(.A1(new_n402), .A2(KEYINPUT33), .A3(new_n388), .ZN(new_n621));
  NOR2_X1   g435(.A1(new_n406), .A2(G902), .ZN(new_n622));
  NAND3_X1  g436(.A1(new_n620), .A2(new_n621), .A3(new_n622), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n403), .A2(new_n265), .ZN(new_n624));
  NAND2_X1  g438(.A1(new_n624), .A2(new_n406), .ZN(new_n625));
  NAND2_X1  g439(.A1(new_n623), .A2(new_n625), .ZN(new_n626));
  INV_X1    g440(.A(new_n626), .ZN(new_n627));
  NOR2_X1   g441(.A1(new_n574), .A2(new_n575), .ZN(new_n628));
  AOI22_X1  g442(.A1(new_n453), .A2(new_n455), .B1(KEYINPUT17), .B2(new_n457), .ZN(new_n629));
  INV_X1    g443(.A(new_n482), .ZN(new_n630));
  INV_X1    g444(.A(new_n483), .ZN(new_n631));
  AOI22_X1  g445(.A1(new_n628), .A2(new_n629), .B1(new_n630), .B2(new_n631), .ZN(new_n632));
  OAI21_X1  g446(.A(new_n476), .B1(new_n632), .B2(new_n447), .ZN(new_n633));
  AOI21_X1  g447(.A(new_n495), .B1(new_n633), .B2(new_n265), .ZN(new_n634));
  INV_X1    g448(.A(new_n489), .ZN(new_n635));
  NAND3_X1  g449(.A1(new_n487), .A2(new_n422), .A3(new_n488), .ZN(new_n636));
  AOI21_X1  g450(.A(new_n634), .B1(new_n635), .B2(new_n636), .ZN(new_n637));
  NOR2_X1   g451(.A1(new_n627), .A2(new_n637), .ZN(new_n638));
  OAI211_X1 g452(.A(new_n187), .B(new_n420), .C1(new_n283), .C2(new_n289), .ZN(new_n639));
  INV_X1    g453(.A(new_n639), .ZN(new_n640));
  NAND4_X1  g454(.A1(new_n614), .A2(new_n618), .A3(new_n638), .A4(new_n640), .ZN(new_n641));
  XOR2_X1   g455(.A(KEYINPUT34), .B(G104), .Z(new_n642));
  XNOR2_X1  g456(.A(new_n641), .B(new_n642), .ZN(G6));
  INV_X1    g457(.A(KEYINPUT91), .ZN(new_n644));
  NOR2_X1   g458(.A1(new_n636), .A2(new_n644), .ZN(new_n645));
  NOR2_X1   g459(.A1(new_n489), .A2(new_n491), .ZN(new_n646));
  AOI21_X1  g460(.A(new_n645), .B1(new_n646), .B2(new_n644), .ZN(new_n647));
  AOI21_X1  g461(.A(new_n634), .B1(new_n408), .B2(new_n410), .ZN(new_n648));
  AND2_X1   g462(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  AND2_X1   g463(.A1(new_n640), .A2(new_n649), .ZN(new_n650));
  NAND3_X1  g464(.A1(new_n650), .A2(new_n618), .A3(new_n614), .ZN(new_n651));
  XOR2_X1   g465(.A(KEYINPUT35), .B(G107), .Z(new_n652));
  XNOR2_X1  g466(.A(new_n651), .B(new_n652), .ZN(G9));
  OR2_X1    g467(.A1(new_n583), .A2(KEYINPUT36), .ZN(new_n654));
  XNOR2_X1  g468(.A(new_n579), .B(new_n654), .ZN(new_n655));
  NOR2_X1   g469(.A1(new_n655), .A2(new_n600), .ZN(new_n656));
  NOR2_X1   g470(.A1(new_n593), .A2(new_n656), .ZN(new_n657));
  INV_X1    g471(.A(new_n657), .ZN(new_n658));
  NAND3_X1  g472(.A1(new_n499), .A2(new_n611), .A3(new_n658), .ZN(new_n659));
  XOR2_X1   g473(.A(KEYINPUT37), .B(G110), .Z(new_n660));
  XNOR2_X1  g474(.A(new_n659), .B(new_n660), .ZN(G12));
  INV_X1    g475(.A(new_n187), .ZN(new_n662));
  NAND2_X1  g476(.A1(new_n287), .A2(new_n288), .ZN(new_n663));
  NAND2_X1  g477(.A1(new_n663), .A2(new_n268), .ZN(new_n664));
  NAND3_X1  g478(.A1(new_n287), .A2(new_n288), .A3(new_n284), .ZN(new_n665));
  AOI21_X1  g479(.A(new_n662), .B1(new_n664), .B2(new_n665), .ZN(new_n666));
  NAND2_X1  g480(.A1(new_n646), .A2(new_n644), .ZN(new_n667));
  INV_X1    g481(.A(new_n645), .ZN(new_n668));
  INV_X1    g482(.A(new_n412), .ZN(new_n669));
  OAI21_X1  g483(.A(new_n669), .B1(new_n416), .B2(G900), .ZN(new_n670));
  XNOR2_X1  g484(.A(new_n670), .B(KEYINPUT92), .ZN(new_n671));
  NAND4_X1  g485(.A1(new_n648), .A2(new_n667), .A3(new_n668), .A4(new_n671), .ZN(new_n672));
  NAND2_X1  g486(.A1(new_n672), .A2(KEYINPUT93), .ZN(new_n673));
  INV_X1    g487(.A(KEYINPUT93), .ZN(new_n674));
  NAND4_X1  g488(.A1(new_n647), .A2(new_n674), .A3(new_n648), .A4(new_n671), .ZN(new_n675));
  NAND3_X1  g489(.A1(new_n666), .A2(new_n673), .A3(new_n675), .ZN(new_n676));
  INV_X1    g490(.A(KEYINPUT94), .ZN(new_n677));
  NAND2_X1  g491(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  NOR3_X1   g492(.A1(new_n657), .A2(new_n613), .A3(new_n557), .ZN(new_n679));
  NAND4_X1  g493(.A1(new_n666), .A2(new_n673), .A3(KEYINPUT94), .A4(new_n675), .ZN(new_n680));
  NAND3_X1  g494(.A1(new_n678), .A2(new_n679), .A3(new_n680), .ZN(new_n681));
  XNOR2_X1  g495(.A(new_n681), .B(G128), .ZN(G30));
  NAND2_X1  g496(.A1(new_n408), .A2(new_n410), .ZN(new_n683));
  NAND4_X1  g497(.A1(new_n657), .A2(new_n187), .A3(new_n496), .A4(new_n683), .ZN(new_n684));
  XNOR2_X1  g498(.A(new_n684), .B(KEYINPUT97), .ZN(new_n685));
  XNOR2_X1  g499(.A(new_n671), .B(KEYINPUT39), .ZN(new_n686));
  NAND2_X1  g500(.A1(new_n617), .A2(new_n686), .ZN(new_n687));
  XOR2_X1   g501(.A(new_n687), .B(KEYINPUT40), .Z(new_n688));
  NAND2_X1  g502(.A1(new_n549), .A2(new_n556), .ZN(new_n689));
  NOR2_X1   g503(.A1(new_n508), .A2(new_n512), .ZN(new_n690));
  NOR2_X1   g504(.A1(new_n690), .A2(new_n517), .ZN(new_n691));
  OAI21_X1  g505(.A(KEYINPUT95), .B1(new_n550), .B2(new_n691), .ZN(new_n692));
  NAND2_X1  g506(.A1(new_n692), .A2(new_n265), .ZN(new_n693));
  NOR3_X1   g507(.A1(new_n550), .A2(KEYINPUT95), .A3(new_n691), .ZN(new_n694));
  OAI21_X1  g508(.A(G472), .B1(new_n693), .B2(new_n694), .ZN(new_n695));
  NAND2_X1  g509(.A1(new_n689), .A2(new_n695), .ZN(new_n696));
  INV_X1    g510(.A(KEYINPUT96), .ZN(new_n697));
  NAND2_X1  g511(.A1(new_n696), .A2(new_n697), .ZN(new_n698));
  NAND3_X1  g512(.A1(new_n689), .A2(KEYINPUT96), .A3(new_n695), .ZN(new_n699));
  NAND2_X1  g513(.A1(new_n698), .A2(new_n699), .ZN(new_n700));
  NAND2_X1  g514(.A1(new_n664), .A2(new_n665), .ZN(new_n701));
  XNOR2_X1  g515(.A(new_n701), .B(KEYINPUT38), .ZN(new_n702));
  NAND4_X1  g516(.A1(new_n685), .A2(new_n688), .A3(new_n700), .A4(new_n702), .ZN(new_n703));
  XNOR2_X1  g517(.A(new_n703), .B(G143), .ZN(G45));
  AND3_X1   g518(.A1(new_n626), .A2(new_n496), .A3(new_n671), .ZN(new_n705));
  AND2_X1   g519(.A1(new_n666), .A2(new_n705), .ZN(new_n706));
  NAND2_X1  g520(.A1(new_n706), .A2(new_n679), .ZN(new_n707));
  XNOR2_X1  g521(.A(new_n707), .B(G146), .ZN(G48));
  INV_X1    g522(.A(new_n535), .ZN(new_n709));
  NOR3_X1   g523(.A1(new_n546), .A2(KEYINPUT32), .A3(new_n548), .ZN(new_n710));
  AOI21_X1  g524(.A(new_n555), .B1(new_n554), .B2(new_n547), .ZN(new_n711));
  OAI21_X1  g525(.A(new_n709), .B1(new_n710), .B2(new_n711), .ZN(new_n712));
  NAND3_X1  g526(.A1(new_n712), .A2(new_n608), .A3(new_n607), .ZN(new_n713));
  NOR2_X1   g527(.A1(new_n315), .A2(new_n318), .ZN(new_n714));
  NOR2_X1   g528(.A1(new_n334), .A2(new_n714), .ZN(new_n715));
  AOI21_X1  g529(.A(new_n333), .B1(new_n342), .B2(new_n328), .ZN(new_n716));
  OAI211_X1 g530(.A(new_n340), .B(new_n265), .C1(new_n715), .C2(new_n716), .ZN(new_n717));
  INV_X1    g531(.A(KEYINPUT98), .ZN(new_n718));
  NAND2_X1  g532(.A1(new_n717), .A2(new_n718), .ZN(new_n719));
  NAND2_X1  g533(.A1(new_n344), .A2(new_n345), .ZN(new_n720));
  AOI21_X1  g534(.A(new_n340), .B1(new_n720), .B2(new_n265), .ZN(new_n721));
  NOR2_X1   g535(.A1(new_n719), .A2(new_n721), .ZN(new_n722));
  NOR3_X1   g536(.A1(new_n346), .A2(new_n718), .A3(new_n340), .ZN(new_n723));
  OAI21_X1  g537(.A(new_n353), .B1(new_n722), .B2(new_n723), .ZN(new_n724));
  NOR2_X1   g538(.A1(new_n713), .A2(new_n724), .ZN(new_n725));
  NAND3_X1  g539(.A1(new_n725), .A2(new_n638), .A3(new_n640), .ZN(new_n726));
  XNOR2_X1  g540(.A(KEYINPUT41), .B(G113), .ZN(new_n727));
  XNOR2_X1  g541(.A(new_n727), .B(KEYINPUT99), .ZN(new_n728));
  XNOR2_X1  g542(.A(new_n726), .B(new_n728), .ZN(G15));
  NAND2_X1  g543(.A1(new_n650), .A2(new_n725), .ZN(new_n730));
  XNOR2_X1  g544(.A(KEYINPUT100), .B(G116), .ZN(new_n731));
  XNOR2_X1  g545(.A(new_n730), .B(new_n731), .ZN(G18));
  NOR4_X1   g546(.A1(new_n657), .A2(new_n557), .A3(new_n496), .A4(new_n421), .ZN(new_n733));
  NOR3_X1   g547(.A1(new_n290), .A2(new_n724), .A3(KEYINPUT101), .ZN(new_n734));
  INV_X1    g548(.A(KEYINPUT101), .ZN(new_n735));
  INV_X1    g549(.A(new_n723), .ZN(new_n736));
  OAI21_X1  g550(.A(new_n265), .B1(new_n715), .B2(new_n716), .ZN(new_n737));
  NAND2_X1  g551(.A1(new_n737), .A2(G469), .ZN(new_n738));
  NAND3_X1  g552(.A1(new_n738), .A2(new_n718), .A3(new_n717), .ZN(new_n739));
  AOI21_X1  g553(.A(new_n352), .B1(new_n736), .B2(new_n739), .ZN(new_n740));
  AOI21_X1  g554(.A(new_n735), .B1(new_n666), .B2(new_n740), .ZN(new_n741));
  OAI21_X1  g555(.A(new_n733), .B1(new_n734), .B2(new_n741), .ZN(new_n742));
  XNOR2_X1  g556(.A(new_n742), .B(G119), .ZN(G21));
  OAI211_X1 g557(.A(new_n353), .B(new_n420), .C1(new_n722), .C2(new_n723), .ZN(new_n744));
  INV_X1    g558(.A(KEYINPUT102), .ZN(new_n745));
  NAND2_X1  g559(.A1(new_n546), .A2(new_n745), .ZN(new_n746));
  AOI21_X1  g560(.A(new_n548), .B1(new_n609), .B2(KEYINPUT102), .ZN(new_n747));
  AOI22_X1  g561(.A1(new_n746), .A2(new_n747), .B1(new_n610), .B2(G472), .ZN(new_n748));
  NAND3_X1  g562(.A1(new_n607), .A2(new_n608), .A3(new_n748), .ZN(new_n749));
  NOR2_X1   g563(.A1(new_n744), .A2(new_n749), .ZN(new_n750));
  INV_X1    g564(.A(KEYINPUT103), .ZN(new_n751));
  INV_X1    g565(.A(new_n683), .ZN(new_n752));
  OAI21_X1  g566(.A(new_n751), .B1(new_n752), .B2(new_n637), .ZN(new_n753));
  NAND3_X1  g567(.A1(new_n683), .A2(new_n496), .A3(KEYINPUT103), .ZN(new_n754));
  NAND2_X1  g568(.A1(new_n753), .A2(new_n754), .ZN(new_n755));
  NOR2_X1   g569(.A1(new_n755), .A2(new_n290), .ZN(new_n756));
  NAND2_X1  g570(.A1(new_n750), .A2(new_n756), .ZN(new_n757));
  XNOR2_X1  g571(.A(new_n757), .B(G122), .ZN(G24));
  OAI211_X1 g572(.A(new_n705), .B(new_n748), .C1(new_n593), .C2(new_n656), .ZN(new_n759));
  INV_X1    g573(.A(new_n759), .ZN(new_n760));
  OAI21_X1  g574(.A(new_n760), .B1(new_n734), .B2(new_n741), .ZN(new_n761));
  XNOR2_X1  g575(.A(new_n761), .B(G125), .ZN(G27));
  INV_X1    g576(.A(new_n341), .ZN(new_n763));
  NAND2_X1  g577(.A1(new_n717), .A2(new_n763), .ZN(new_n764));
  NOR2_X1   g578(.A1(new_n336), .A2(new_n314), .ZN(new_n765));
  OAI21_X1  g579(.A(KEYINPUT77), .B1(new_n714), .B2(new_n765), .ZN(new_n766));
  AOI21_X1  g580(.A(new_n333), .B1(new_n766), .B2(new_n330), .ZN(new_n767));
  NOR3_X1   g581(.A1(new_n767), .A2(new_n340), .A3(new_n337), .ZN(new_n768));
  INV_X1    g582(.A(KEYINPUT104), .ZN(new_n769));
  AOI21_X1  g583(.A(new_n764), .B1(new_n768), .B2(new_n769), .ZN(new_n770));
  NAND2_X1  g584(.A1(new_n339), .A2(KEYINPUT104), .ZN(new_n771));
  AOI21_X1  g585(.A(new_n352), .B1(new_n770), .B2(new_n771), .ZN(new_n772));
  NOR3_X1   g586(.A1(new_n283), .A2(new_n289), .A3(new_n662), .ZN(new_n773));
  NAND4_X1  g587(.A1(new_n772), .A2(new_n602), .A3(new_n705), .A4(new_n773), .ZN(new_n774));
  INV_X1    g588(.A(KEYINPUT42), .ZN(new_n775));
  AOI21_X1  g589(.A(KEYINPUT106), .B1(new_n775), .B2(KEYINPUT105), .ZN(new_n776));
  NAND2_X1  g590(.A1(new_n774), .A2(new_n776), .ZN(new_n777));
  NAND4_X1  g591(.A1(new_n332), .A2(new_n769), .A3(G469), .A4(new_n338), .ZN(new_n778));
  NAND2_X1  g592(.A1(new_n778), .A2(new_n347), .ZN(new_n779));
  NAND2_X1  g593(.A1(new_n766), .A2(new_n330), .ZN(new_n780));
  AOI21_X1  g594(.A(new_n337), .B1(new_n780), .B2(new_n293), .ZN(new_n781));
  AOI21_X1  g595(.A(new_n769), .B1(new_n781), .B2(G469), .ZN(new_n782));
  OAI21_X1  g596(.A(new_n353), .B1(new_n779), .B2(new_n782), .ZN(new_n783));
  NAND3_X1  g597(.A1(new_n664), .A2(new_n187), .A3(new_n665), .ZN(new_n784));
  NOR2_X1   g598(.A1(new_n783), .A2(new_n784), .ZN(new_n785));
  AOI21_X1  g599(.A(new_n776), .B1(KEYINPUT106), .B2(new_n775), .ZN(new_n786));
  NAND4_X1  g600(.A1(new_n785), .A2(new_n602), .A3(new_n705), .A4(new_n786), .ZN(new_n787));
  NAND2_X1  g601(.A1(new_n777), .A2(new_n787), .ZN(new_n788));
  XNOR2_X1  g602(.A(new_n788), .B(new_n312), .ZN(G33));
  AND2_X1   g603(.A1(new_n673), .A2(new_n675), .ZN(new_n790));
  NAND3_X1  g604(.A1(new_n785), .A2(new_n790), .A3(new_n602), .ZN(new_n791));
  XNOR2_X1  g605(.A(new_n791), .B(G134), .ZN(G36));
  NAND2_X1  g606(.A1(new_n637), .A2(new_n626), .ZN(new_n793));
  INV_X1    g607(.A(KEYINPUT43), .ZN(new_n794));
  XNOR2_X1  g608(.A(new_n793), .B(new_n794), .ZN(new_n795));
  INV_X1    g609(.A(new_n611), .ZN(new_n796));
  NAND3_X1  g610(.A1(new_n795), .A2(new_n796), .A3(new_n658), .ZN(new_n797));
  INV_X1    g611(.A(KEYINPUT44), .ZN(new_n798));
  OR2_X1    g612(.A1(new_n797), .A2(new_n798), .ZN(new_n799));
  XNOR2_X1  g613(.A(new_n773), .B(KEYINPUT107), .ZN(new_n800));
  NAND2_X1  g614(.A1(new_n797), .A2(new_n798), .ZN(new_n801));
  NAND3_X1  g615(.A1(new_n799), .A2(new_n800), .A3(new_n801), .ZN(new_n802));
  NAND2_X1  g616(.A1(new_n802), .A2(KEYINPUT108), .ZN(new_n803));
  INV_X1    g617(.A(KEYINPUT46), .ZN(new_n804));
  OR2_X1    g618(.A1(new_n781), .A2(KEYINPUT45), .ZN(new_n805));
  NAND2_X1  g619(.A1(new_n781), .A2(KEYINPUT45), .ZN(new_n806));
  NAND3_X1  g620(.A1(new_n805), .A2(G469), .A3(new_n806), .ZN(new_n807));
  INV_X1    g621(.A(new_n807), .ZN(new_n808));
  OAI21_X1  g622(.A(new_n804), .B1(new_n808), .B2(new_n341), .ZN(new_n809));
  NAND3_X1  g623(.A1(new_n807), .A2(KEYINPUT46), .A3(new_n763), .ZN(new_n810));
  NAND3_X1  g624(.A1(new_n809), .A2(new_n717), .A3(new_n810), .ZN(new_n811));
  AND3_X1   g625(.A1(new_n811), .A2(new_n353), .A3(new_n686), .ZN(new_n812));
  INV_X1    g626(.A(KEYINPUT108), .ZN(new_n813));
  NAND4_X1  g627(.A1(new_n799), .A2(new_n813), .A3(new_n800), .A4(new_n801), .ZN(new_n814));
  NAND3_X1  g628(.A1(new_n803), .A2(new_n812), .A3(new_n814), .ZN(new_n815));
  XNOR2_X1  g629(.A(new_n815), .B(G137), .ZN(G39));
  NAND2_X1  g630(.A1(new_n811), .A2(new_n353), .ZN(new_n817));
  INV_X1    g631(.A(KEYINPUT47), .ZN(new_n818));
  NAND2_X1  g632(.A1(new_n817), .A2(new_n818), .ZN(new_n819));
  NAND3_X1  g633(.A1(new_n811), .A2(KEYINPUT47), .A3(new_n353), .ZN(new_n820));
  NAND2_X1  g634(.A1(new_n819), .A2(new_n820), .ZN(new_n821));
  NAND2_X1  g635(.A1(new_n607), .A2(new_n608), .ZN(new_n822));
  NAND4_X1  g636(.A1(new_n773), .A2(new_n822), .A3(new_n557), .A4(new_n705), .ZN(new_n823));
  XNOR2_X1  g637(.A(new_n823), .B(KEYINPUT109), .ZN(new_n824));
  NAND2_X1  g638(.A1(new_n821), .A2(new_n824), .ZN(new_n825));
  XNOR2_X1  g639(.A(new_n825), .B(G140), .ZN(G42));
  INV_X1    g640(.A(KEYINPUT54), .ZN(new_n827));
  AND2_X1   g641(.A1(new_n657), .A2(new_n671), .ZN(new_n828));
  NAND4_X1  g642(.A1(new_n700), .A2(new_n756), .A3(new_n828), .A4(new_n772), .ZN(new_n829));
  NAND4_X1  g643(.A1(new_n681), .A2(new_n761), .A3(new_n707), .A4(new_n829), .ZN(new_n830));
  XNOR2_X1  g644(.A(new_n830), .B(KEYINPUT52), .ZN(new_n831));
  INV_X1    g645(.A(KEYINPUT53), .ZN(new_n832));
  INV_X1    g646(.A(new_n634), .ZN(new_n833));
  AND4_X1   g647(.A1(new_n833), .A2(new_n647), .A3(new_n752), .A4(new_n671), .ZN(new_n834));
  NAND3_X1  g648(.A1(new_n679), .A2(new_n773), .A3(new_n834), .ZN(new_n835));
  AOI21_X1  g649(.A(KEYINPUT111), .B1(new_n785), .B2(new_n760), .ZN(new_n836));
  INV_X1    g650(.A(KEYINPUT111), .ZN(new_n837));
  NOR4_X1   g651(.A1(new_n783), .A2(new_n759), .A3(new_n784), .A4(new_n837), .ZN(new_n838));
  OAI21_X1  g652(.A(new_n835), .B1(new_n836), .B2(new_n838), .ZN(new_n839));
  NAND3_X1  g653(.A1(new_n777), .A2(new_n787), .A3(new_n791), .ZN(new_n840));
  NOR2_X1   g654(.A1(new_n839), .A2(new_n840), .ZN(new_n841));
  NAND2_X1  g655(.A1(new_n637), .A2(new_n683), .ZN(new_n842));
  NOR2_X1   g656(.A1(new_n639), .A2(new_n842), .ZN(new_n843));
  NAND3_X1  g657(.A1(new_n614), .A2(new_n843), .A3(new_n618), .ZN(new_n844));
  NAND2_X1  g658(.A1(new_n844), .A2(new_n659), .ZN(new_n845));
  NAND2_X1  g659(.A1(new_n845), .A2(KEYINPUT110), .ZN(new_n846));
  INV_X1    g660(.A(KEYINPUT110), .ZN(new_n847));
  NAND3_X1  g661(.A1(new_n844), .A2(new_n847), .A3(new_n659), .ZN(new_n848));
  NAND2_X1  g662(.A1(new_n846), .A2(new_n848), .ZN(new_n849));
  OAI211_X1 g663(.A(new_n725), .B(new_n640), .C1(new_n638), .C2(new_n649), .ZN(new_n850));
  AOI22_X1  g664(.A1(new_n756), .A2(new_n750), .B1(new_n499), .B2(new_n602), .ZN(new_n851));
  AND4_X1   g665(.A1(new_n641), .A2(new_n742), .A3(new_n850), .A4(new_n851), .ZN(new_n852));
  NAND3_X1  g666(.A1(new_n841), .A2(new_n849), .A3(new_n852), .ZN(new_n853));
  NOR3_X1   g667(.A1(new_n831), .A2(new_n832), .A3(new_n853), .ZN(new_n854));
  AND3_X1   g668(.A1(new_n841), .A2(new_n849), .A3(new_n852), .ZN(new_n855));
  AND2_X1   g669(.A1(new_n680), .A2(new_n679), .ZN(new_n856));
  AOI22_X1  g670(.A1(new_n856), .A2(new_n678), .B1(new_n679), .B2(new_n706), .ZN(new_n857));
  NAND4_X1  g671(.A1(new_n857), .A2(KEYINPUT52), .A3(new_n761), .A4(new_n829), .ZN(new_n858));
  INV_X1    g672(.A(KEYINPUT52), .ZN(new_n859));
  NAND2_X1  g673(.A1(new_n830), .A2(new_n859), .ZN(new_n860));
  NAND2_X1  g674(.A1(new_n858), .A2(new_n860), .ZN(new_n861));
  AOI21_X1  g675(.A(KEYINPUT53), .B1(new_n855), .B2(new_n861), .ZN(new_n862));
  OAI21_X1  g676(.A(new_n827), .B1(new_n854), .B2(new_n862), .ZN(new_n863));
  OAI21_X1  g677(.A(new_n832), .B1(new_n831), .B2(new_n853), .ZN(new_n864));
  NAND3_X1  g678(.A1(new_n855), .A2(KEYINPUT53), .A3(new_n861), .ZN(new_n865));
  NAND3_X1  g679(.A1(new_n864), .A2(KEYINPUT54), .A3(new_n865), .ZN(new_n866));
  NAND2_X1  g680(.A1(new_n863), .A2(new_n866), .ZN(new_n867));
  INV_X1    g681(.A(new_n702), .ZN(new_n868));
  INV_X1    g682(.A(new_n749), .ZN(new_n869));
  AND3_X1   g683(.A1(new_n795), .A2(new_n869), .A3(new_n412), .ZN(new_n870));
  NOR2_X1   g684(.A1(new_n724), .A2(new_n187), .ZN(new_n871));
  NAND4_X1  g685(.A1(new_n868), .A2(new_n870), .A3(KEYINPUT50), .A4(new_n871), .ZN(new_n872));
  INV_X1    g686(.A(KEYINPUT50), .ZN(new_n873));
  NAND4_X1  g687(.A1(new_n871), .A2(new_n795), .A3(new_n869), .A4(new_n412), .ZN(new_n874));
  OAI21_X1  g688(.A(new_n873), .B1(new_n874), .B2(new_n702), .ZN(new_n875));
  NOR2_X1   g689(.A1(new_n724), .A2(new_n669), .ZN(new_n876));
  AND3_X1   g690(.A1(new_n876), .A2(new_n773), .A3(new_n795), .ZN(new_n877));
  AND2_X1   g691(.A1(new_n658), .A2(new_n748), .ZN(new_n878));
  AOI22_X1  g692(.A1(new_n872), .A2(new_n875), .B1(new_n877), .B2(new_n878), .ZN(new_n879));
  NAND2_X1  g693(.A1(new_n876), .A2(new_n773), .ZN(new_n880));
  NAND3_X1  g694(.A1(new_n698), .A2(new_n615), .A3(new_n699), .ZN(new_n881));
  NOR2_X1   g695(.A1(new_n880), .A2(new_n881), .ZN(new_n882));
  INV_X1    g696(.A(KEYINPUT112), .ZN(new_n883));
  NAND2_X1  g697(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  OAI21_X1  g698(.A(KEYINPUT112), .B1(new_n880), .B2(new_n881), .ZN(new_n885));
  NAND4_X1  g699(.A1(new_n884), .A2(new_n637), .A3(new_n627), .A4(new_n885), .ZN(new_n886));
  NAND2_X1  g700(.A1(new_n879), .A2(new_n886), .ZN(new_n887));
  NAND2_X1  g701(.A1(new_n736), .A2(new_n739), .ZN(new_n888));
  NAND2_X1  g702(.A1(new_n888), .A2(new_n352), .ZN(new_n889));
  NAND3_X1  g703(.A1(new_n819), .A2(new_n820), .A3(new_n889), .ZN(new_n890));
  AND2_X1   g704(.A1(new_n800), .A2(new_n870), .ZN(new_n891));
  AOI21_X1  g705(.A(new_n887), .B1(new_n890), .B2(new_n891), .ZN(new_n892));
  NOR2_X1   g706(.A1(new_n892), .A2(KEYINPUT51), .ZN(new_n893));
  NAND2_X1  g707(.A1(new_n877), .A2(new_n602), .ZN(new_n894));
  XNOR2_X1  g708(.A(new_n894), .B(KEYINPUT48), .ZN(new_n895));
  NAND3_X1  g709(.A1(new_n884), .A2(new_n638), .A3(new_n885), .ZN(new_n896));
  OR2_X1    g710(.A1(new_n734), .A2(new_n741), .ZN(new_n897));
  AOI211_X1 g711(.A(new_n411), .B(G953), .C1(new_n897), .C2(new_n870), .ZN(new_n898));
  NAND3_X1  g712(.A1(new_n895), .A2(new_n896), .A3(new_n898), .ZN(new_n899));
  NOR2_X1   g713(.A1(new_n893), .A2(new_n899), .ZN(new_n900));
  INV_X1    g714(.A(KEYINPUT114), .ZN(new_n901));
  OR2_X1    g715(.A1(new_n890), .A2(new_n901), .ZN(new_n902));
  NAND2_X1  g716(.A1(new_n890), .A2(new_n901), .ZN(new_n903));
  AND3_X1   g717(.A1(new_n902), .A2(new_n903), .A3(new_n891), .ZN(new_n904));
  NOR2_X1   g718(.A1(new_n887), .A2(KEYINPUT113), .ZN(new_n905));
  INV_X1    g719(.A(KEYINPUT113), .ZN(new_n906));
  AOI21_X1  g720(.A(new_n906), .B1(new_n879), .B2(new_n886), .ZN(new_n907));
  OAI21_X1  g721(.A(KEYINPUT51), .B1(new_n905), .B2(new_n907), .ZN(new_n908));
  NOR2_X1   g722(.A1(new_n904), .A2(new_n908), .ZN(new_n909));
  INV_X1    g723(.A(KEYINPUT115), .ZN(new_n910));
  NOR2_X1   g724(.A1(new_n909), .A2(new_n910), .ZN(new_n911));
  NOR3_X1   g725(.A1(new_n904), .A2(new_n908), .A3(KEYINPUT115), .ZN(new_n912));
  OAI211_X1 g726(.A(new_n867), .B(new_n900), .C1(new_n911), .C2(new_n912), .ZN(new_n913));
  NAND2_X1  g727(.A1(new_n411), .A2(new_n208), .ZN(new_n914));
  NAND2_X1  g728(.A1(new_n913), .A2(new_n914), .ZN(new_n915));
  XOR2_X1   g729(.A(new_n888), .B(KEYINPUT49), .Z(new_n916));
  OR4_X1    g730(.A1(new_n822), .A2(new_n662), .A3(new_n352), .A4(new_n793), .ZN(new_n917));
  OR4_X1    g731(.A1(new_n700), .A2(new_n916), .A3(new_n917), .A4(new_n702), .ZN(new_n918));
  NAND2_X1  g732(.A1(new_n915), .A2(new_n918), .ZN(G75));
  NOR2_X1   g733(.A1(new_n208), .A2(G952), .ZN(new_n920));
  INV_X1    g734(.A(new_n920), .ZN(new_n921));
  AOI21_X1  g735(.A(new_n265), .B1(new_n864), .B2(new_n865), .ZN(new_n922));
  NAND2_X1  g736(.A1(new_n922), .A2(new_n268), .ZN(new_n923));
  INV_X1    g737(.A(KEYINPUT56), .ZN(new_n924));
  NAND2_X1  g738(.A1(new_n923), .A2(new_n924), .ZN(new_n925));
  XNOR2_X1  g739(.A(new_n281), .B(new_n282), .ZN(new_n926));
  XNOR2_X1  g740(.A(new_n926), .B(KEYINPUT55), .ZN(new_n927));
  OAI21_X1  g741(.A(new_n921), .B1(new_n925), .B2(new_n927), .ZN(new_n928));
  NAND2_X1  g742(.A1(new_n925), .A2(new_n927), .ZN(new_n929));
  INV_X1    g743(.A(KEYINPUT116), .ZN(new_n930));
  NAND2_X1  g744(.A1(new_n929), .A2(new_n930), .ZN(new_n931));
  NAND3_X1  g745(.A1(new_n925), .A2(KEYINPUT116), .A3(new_n927), .ZN(new_n932));
  AOI21_X1  g746(.A(new_n928), .B1(new_n931), .B2(new_n932), .ZN(G51));
  XNOR2_X1  g747(.A(new_n341), .B(KEYINPUT117), .ZN(new_n934));
  XOR2_X1   g748(.A(new_n934), .B(KEYINPUT57), .Z(new_n935));
  NAND3_X1  g749(.A1(new_n863), .A2(new_n866), .A3(new_n935), .ZN(new_n936));
  INV_X1    g750(.A(KEYINPUT118), .ZN(new_n937));
  NAND3_X1  g751(.A1(new_n936), .A2(new_n937), .A3(new_n720), .ZN(new_n938));
  NAND2_X1  g752(.A1(new_n922), .A2(new_n808), .ZN(new_n939));
  AND2_X1   g753(.A1(new_n938), .A2(new_n939), .ZN(new_n940));
  NAND2_X1  g754(.A1(new_n936), .A2(new_n720), .ZN(new_n941));
  NAND2_X1  g755(.A1(new_n941), .A2(KEYINPUT118), .ZN(new_n942));
  AOI21_X1  g756(.A(new_n920), .B1(new_n940), .B2(new_n942), .ZN(G54));
  AND2_X1   g757(.A1(KEYINPUT58), .A2(G475), .ZN(new_n944));
  AND3_X1   g758(.A1(new_n922), .A2(new_n487), .A3(new_n944), .ZN(new_n945));
  AOI21_X1  g759(.A(new_n487), .B1(new_n922), .B2(new_n944), .ZN(new_n946));
  NOR3_X1   g760(.A1(new_n945), .A2(new_n946), .A3(new_n920), .ZN(G60));
  NAND2_X1  g761(.A1(G478), .A2(G902), .ZN(new_n948));
  XNOR2_X1  g762(.A(new_n948), .B(KEYINPUT119), .ZN(new_n949));
  XNOR2_X1  g763(.A(new_n949), .B(KEYINPUT59), .ZN(new_n950));
  NAND3_X1  g764(.A1(new_n863), .A2(new_n866), .A3(new_n950), .ZN(new_n951));
  AND2_X1   g765(.A1(new_n620), .A2(new_n621), .ZN(new_n952));
  INV_X1    g766(.A(new_n952), .ZN(new_n953));
  AND2_X1   g767(.A1(new_n951), .A2(new_n953), .ZN(new_n954));
  NOR2_X1   g768(.A1(new_n951), .A2(new_n953), .ZN(new_n955));
  NOR3_X1   g769(.A1(new_n954), .A2(new_n955), .A3(new_n920), .ZN(G63));
  NAND2_X1  g770(.A1(new_n864), .A2(new_n865), .ZN(new_n957));
  INV_X1    g771(.A(new_n655), .ZN(new_n958));
  XNOR2_X1  g772(.A(KEYINPUT120), .B(KEYINPUT60), .ZN(new_n959));
  NOR2_X1   g773(.A1(new_n370), .A2(new_n265), .ZN(new_n960));
  XNOR2_X1  g774(.A(new_n959), .B(new_n960), .ZN(new_n961));
  NAND3_X1  g775(.A1(new_n957), .A2(new_n958), .A3(new_n961), .ZN(new_n962));
  AOI21_X1  g776(.A(KEYINPUT61), .B1(new_n962), .B2(KEYINPUT121), .ZN(new_n963));
  INV_X1    g777(.A(new_n963), .ZN(new_n964));
  INV_X1    g778(.A(new_n961), .ZN(new_n965));
  AOI21_X1  g779(.A(new_n965), .B1(new_n864), .B2(new_n865), .ZN(new_n966));
  AOI21_X1  g780(.A(new_n920), .B1(new_n966), .B2(new_n958), .ZN(new_n967));
  INV_X1    g781(.A(KEYINPUT122), .ZN(new_n968));
  OAI21_X1  g782(.A(new_n961), .B1(new_n854), .B2(new_n862), .ZN(new_n969));
  NAND2_X1  g783(.A1(new_n969), .A2(new_n598), .ZN(new_n970));
  AND3_X1   g784(.A1(new_n967), .A2(new_n968), .A3(new_n970), .ZN(new_n971));
  AOI21_X1  g785(.A(new_n968), .B1(new_n967), .B2(new_n970), .ZN(new_n972));
  OAI21_X1  g786(.A(new_n964), .B1(new_n971), .B2(new_n972), .ZN(new_n973));
  NAND2_X1  g787(.A1(new_n962), .A2(new_n921), .ZN(new_n974));
  NOR2_X1   g788(.A1(new_n966), .A2(new_n597), .ZN(new_n975));
  OAI21_X1  g789(.A(KEYINPUT122), .B1(new_n974), .B2(new_n975), .ZN(new_n976));
  NAND3_X1  g790(.A1(new_n967), .A2(new_n968), .A3(new_n970), .ZN(new_n977));
  NAND3_X1  g791(.A1(new_n976), .A2(new_n963), .A3(new_n977), .ZN(new_n978));
  NAND2_X1  g792(.A1(new_n973), .A2(new_n978), .ZN(G66));
  INV_X1    g793(.A(new_n418), .ZN(new_n980));
  AOI21_X1  g794(.A(new_n208), .B1(new_n980), .B2(new_n207), .ZN(new_n981));
  NAND2_X1  g795(.A1(new_n849), .A2(new_n852), .ZN(new_n982));
  AOI21_X1  g796(.A(new_n981), .B1(new_n982), .B2(new_n208), .ZN(new_n983));
  INV_X1    g797(.A(G898), .ZN(new_n984));
  AOI21_X1  g798(.A(new_n281), .B1(new_n984), .B2(G953), .ZN(new_n985));
  XNOR2_X1  g799(.A(new_n983), .B(new_n985), .ZN(G69));
  XNOR2_X1  g800(.A(new_n480), .B(KEYINPUT123), .ZN(new_n987));
  XNOR2_X1  g801(.A(new_n532), .B(new_n987), .ZN(new_n988));
  XNOR2_X1  g802(.A(new_n988), .B(KEYINPUT124), .ZN(new_n989));
  AND2_X1   g803(.A1(new_n825), .A2(new_n815), .ZN(new_n990));
  AND3_X1   g804(.A1(new_n681), .A2(new_n707), .A3(new_n761), .ZN(new_n991));
  NAND2_X1  g805(.A1(new_n991), .A2(new_n703), .ZN(new_n992));
  OR2_X1    g806(.A1(new_n992), .A2(KEYINPUT62), .ZN(new_n993));
  NAND2_X1  g807(.A1(new_n992), .A2(KEYINPUT62), .ZN(new_n994));
  AOI21_X1  g808(.A(new_n638), .B1(new_n637), .B2(new_n683), .ZN(new_n995));
  OR4_X1    g809(.A1(new_n713), .A2(new_n995), .A3(new_n687), .A4(new_n784), .ZN(new_n996));
  NAND4_X1  g810(.A1(new_n990), .A2(new_n993), .A3(new_n994), .A4(new_n996), .ZN(new_n997));
  AOI21_X1  g811(.A(new_n989), .B1(new_n997), .B2(new_n208), .ZN(new_n998));
  NOR3_X1   g812(.A1(new_n713), .A2(new_n755), .A3(new_n290), .ZN(new_n999));
  AOI21_X1  g813(.A(new_n840), .B1(new_n812), .B2(new_n999), .ZN(new_n1000));
  NAND4_X1  g814(.A1(new_n825), .A2(new_n815), .A3(new_n991), .A4(new_n1000), .ZN(new_n1001));
  NOR2_X1   g815(.A1(new_n1001), .A2(G953), .ZN(new_n1002));
  INV_X1    g816(.A(G900), .ZN(new_n1003));
  OAI21_X1  g817(.A(new_n988), .B1(new_n1003), .B2(new_n208), .ZN(new_n1004));
  NOR2_X1   g818(.A1(new_n1002), .A2(new_n1004), .ZN(new_n1005));
  NOR2_X1   g819(.A1(new_n998), .A2(new_n1005), .ZN(new_n1006));
  AOI21_X1  g820(.A(new_n208), .B1(G227), .B2(G900), .ZN(new_n1007));
  XOR2_X1   g821(.A(new_n1006), .B(new_n1007), .Z(G72));
  NAND2_X1  g822(.A1(G472), .A2(G902), .ZN(new_n1009));
  XOR2_X1   g823(.A(new_n1009), .B(KEYINPUT63), .Z(new_n1010));
  XOR2_X1   g824(.A(new_n1010), .B(KEYINPUT125), .Z(new_n1011));
  OAI21_X1  g825(.A(new_n1011), .B1(new_n997), .B2(new_n982), .ZN(new_n1012));
  INV_X1    g826(.A(new_n533), .ZN(new_n1013));
  NAND3_X1  g827(.A1(new_n1012), .A2(new_n1013), .A3(new_n517), .ZN(new_n1014));
  NOR2_X1   g828(.A1(new_n533), .A2(new_n517), .ZN(new_n1015));
  OAI21_X1  g829(.A(new_n1010), .B1(new_n1015), .B2(new_n550), .ZN(new_n1016));
  XOR2_X1   g830(.A(new_n1016), .B(KEYINPUT126), .Z(new_n1017));
  NAND2_X1  g831(.A1(new_n957), .A2(new_n1017), .ZN(new_n1018));
  OAI21_X1  g832(.A(new_n1011), .B1(new_n1001), .B2(new_n982), .ZN(new_n1019));
  NOR2_X1   g833(.A1(new_n1013), .A2(new_n517), .ZN(new_n1020));
  AOI21_X1  g834(.A(new_n920), .B1(new_n1019), .B2(new_n1020), .ZN(new_n1021));
  NAND3_X1  g835(.A1(new_n1014), .A2(new_n1018), .A3(new_n1021), .ZN(new_n1022));
  INV_X1    g836(.A(KEYINPUT127), .ZN(new_n1023));
  NAND2_X1  g837(.A1(new_n1022), .A2(new_n1023), .ZN(new_n1024));
  NAND4_X1  g838(.A1(new_n1014), .A2(KEYINPUT127), .A3(new_n1018), .A4(new_n1021), .ZN(new_n1025));
  NAND2_X1  g839(.A1(new_n1024), .A2(new_n1025), .ZN(G57));
endmodule


