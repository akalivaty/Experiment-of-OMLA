//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 0 0 1 1 0 0 0 1 0 1 1 1 0 0 0 0 0 1 0 0 1 0 0 1 1 0 1 1 1 0 1 1 1 1 0 1 0 0 1 0 1 0 1 0 0 1 1 0 0 0 1 1 0 0 0 0 1 0 0 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:18:28 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n698, new_n699,
    new_n700, new_n701, new_n702, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n709, new_n710, new_n712, new_n713, new_n714, new_n715,
    new_n716, new_n717, new_n718, new_n719, new_n720, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n741, new_n742, new_n743, new_n744, new_n745,
    new_n746, new_n747, new_n748, new_n749, new_n750, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n764, new_n765, new_n766, new_n767, new_n769,
    new_n770, new_n771, new_n772, new_n774, new_n775, new_n776, new_n777,
    new_n779, new_n780, new_n781, new_n782, new_n783, new_n784, new_n785,
    new_n786, new_n787, new_n789, new_n791, new_n792, new_n793, new_n794,
    new_n795, new_n796, new_n797, new_n798, new_n799, new_n800, new_n801,
    new_n802, new_n803, new_n804, new_n805, new_n806, new_n807, new_n808,
    new_n809, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n819, new_n820, new_n821, new_n822, new_n823, new_n824,
    new_n825, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n882, new_n884,
    new_n885, new_n886, new_n888, new_n889, new_n890, new_n891, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n946, new_n947, new_n949, new_n950, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n963, new_n964, new_n966, new_n967, new_n968, new_n969,
    new_n970, new_n971, new_n972, new_n974, new_n975, new_n976, new_n977,
    new_n978, new_n980, new_n981, new_n982, new_n983, new_n984, new_n985,
    new_n986, new_n987, new_n988, new_n989, new_n990, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1006, new_n1007;
  AND2_X1   g000(.A1(G227gat), .A2(G233gat), .ZN(new_n202));
  INV_X1    g001(.A(new_n202), .ZN(new_n203));
  INV_X1    g002(.A(G190gat), .ZN(new_n204));
  AND2_X1   g003(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n205));
  NOR2_X1   g004(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n206));
  OAI21_X1  g005(.A(new_n204), .B1(new_n205), .B2(new_n206), .ZN(new_n207));
  NAND2_X1  g006(.A1(new_n207), .A2(KEYINPUT28), .ZN(new_n208));
  NOR2_X1   g007(.A1(G169gat), .A2(G176gat), .ZN(new_n209));
  INV_X1    g008(.A(KEYINPUT26), .ZN(new_n210));
  NAND2_X1  g009(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  OAI21_X1  g010(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n212));
  NAND3_X1  g011(.A1(KEYINPUT66), .A2(G169gat), .A3(G176gat), .ZN(new_n213));
  INV_X1    g012(.A(new_n213), .ZN(new_n214));
  AOI21_X1  g013(.A(KEYINPUT66), .B1(G169gat), .B2(G176gat), .ZN(new_n215));
  OAI211_X1 g014(.A(new_n211), .B(new_n212), .C1(new_n214), .C2(new_n215), .ZN(new_n216));
  INV_X1    g015(.A(G183gat), .ZN(new_n217));
  OAI21_X1  g016(.A(KEYINPUT27), .B1(new_n217), .B2(KEYINPUT67), .ZN(new_n218));
  INV_X1    g017(.A(KEYINPUT67), .ZN(new_n219));
  INV_X1    g018(.A(KEYINPUT27), .ZN(new_n220));
  NAND3_X1  g019(.A1(new_n219), .A2(new_n220), .A3(G183gat), .ZN(new_n221));
  INV_X1    g020(.A(KEYINPUT28), .ZN(new_n222));
  NAND4_X1  g021(.A1(new_n218), .A2(new_n221), .A3(new_n222), .A4(new_n204), .ZN(new_n223));
  NAND2_X1  g022(.A1(G183gat), .A2(G190gat), .ZN(new_n224));
  NAND4_X1  g023(.A1(new_n208), .A2(new_n216), .A3(new_n223), .A4(new_n224), .ZN(new_n225));
  INV_X1    g024(.A(G169gat), .ZN(new_n226));
  INV_X1    g025(.A(G176gat), .ZN(new_n227));
  NAND3_X1  g026(.A1(new_n226), .A2(new_n227), .A3(KEYINPUT23), .ZN(new_n228));
  INV_X1    g027(.A(KEYINPUT23), .ZN(new_n229));
  OAI21_X1  g028(.A(new_n229), .B1(G169gat), .B2(G176gat), .ZN(new_n230));
  OAI211_X1 g029(.A(new_n228), .B(new_n230), .C1(new_n214), .C2(new_n215), .ZN(new_n231));
  INV_X1    g030(.A(KEYINPUT24), .ZN(new_n232));
  NAND3_X1  g031(.A1(new_n232), .A2(G183gat), .A3(G190gat), .ZN(new_n233));
  NAND2_X1  g032(.A1(new_n224), .A2(KEYINPUT24), .ZN(new_n234));
  NOR2_X1   g033(.A1(G183gat), .A2(G190gat), .ZN(new_n235));
  OAI21_X1  g034(.A(new_n233), .B1(new_n234), .B2(new_n235), .ZN(new_n236));
  OAI21_X1  g035(.A(KEYINPUT25), .B1(new_n231), .B2(new_n236), .ZN(new_n237));
  AND2_X1   g036(.A1(new_n225), .A2(new_n237), .ZN(new_n238));
  INV_X1    g037(.A(G127gat), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n239), .A2(KEYINPUT68), .ZN(new_n240));
  INV_X1    g039(.A(KEYINPUT68), .ZN(new_n241));
  NAND2_X1  g040(.A1(new_n241), .A2(G127gat), .ZN(new_n242));
  NAND3_X1  g041(.A1(new_n240), .A2(new_n242), .A3(G134gat), .ZN(new_n243));
  OR2_X1    g042(.A1(G127gat), .A2(G134gat), .ZN(new_n244));
  XNOR2_X1  g043(.A(G113gat), .B(G120gat), .ZN(new_n245));
  OAI211_X1 g044(.A(new_n243), .B(new_n244), .C1(KEYINPUT1), .C2(new_n245), .ZN(new_n246));
  INV_X1    g045(.A(KEYINPUT69), .ZN(new_n247));
  INV_X1    g046(.A(G113gat), .ZN(new_n248));
  OAI21_X1  g047(.A(new_n247), .B1(new_n248), .B2(G120gat), .ZN(new_n249));
  NAND2_X1  g048(.A1(new_n248), .A2(G120gat), .ZN(new_n250));
  INV_X1    g049(.A(G120gat), .ZN(new_n251));
  NAND3_X1  g050(.A1(new_n251), .A2(KEYINPUT69), .A3(G113gat), .ZN(new_n252));
  NAND3_X1  g051(.A1(new_n249), .A2(new_n250), .A3(new_n252), .ZN(new_n253));
  INV_X1    g052(.A(KEYINPUT1), .ZN(new_n254));
  XNOR2_X1  g053(.A(G127gat), .B(G134gat), .ZN(new_n255));
  NAND3_X1  g054(.A1(new_n253), .A2(new_n254), .A3(new_n255), .ZN(new_n256));
  AND2_X1   g055(.A1(new_n246), .A2(new_n256), .ZN(new_n257));
  INV_X1    g056(.A(KEYINPUT64), .ZN(new_n258));
  AOI21_X1  g057(.A(KEYINPUT25), .B1(new_n236), .B2(new_n258), .ZN(new_n259));
  INV_X1    g058(.A(KEYINPUT65), .ZN(new_n260));
  NAND2_X1  g059(.A1(new_n228), .A2(new_n260), .ZN(new_n261));
  NAND3_X1  g060(.A1(new_n209), .A2(KEYINPUT65), .A3(KEYINPUT23), .ZN(new_n262));
  INV_X1    g061(.A(new_n215), .ZN(new_n263));
  AOI22_X1  g062(.A1(new_n261), .A2(new_n262), .B1(new_n263), .B2(new_n213), .ZN(new_n264));
  OAI211_X1 g063(.A(KEYINPUT64), .B(new_n233), .C1(new_n234), .C2(new_n235), .ZN(new_n265));
  NAND4_X1  g064(.A1(new_n259), .A2(new_n230), .A3(new_n264), .A4(new_n265), .ZN(new_n266));
  NAND3_X1  g065(.A1(new_n238), .A2(new_n257), .A3(new_n266), .ZN(new_n267));
  NAND2_X1  g066(.A1(new_n246), .A2(new_n256), .ZN(new_n268));
  NAND2_X1  g067(.A1(new_n261), .A2(new_n262), .ZN(new_n269));
  NAND2_X1  g068(.A1(new_n263), .A2(new_n213), .ZN(new_n270));
  NAND4_X1  g069(.A1(new_n269), .A2(new_n265), .A3(new_n230), .A4(new_n270), .ZN(new_n271));
  INV_X1    g070(.A(KEYINPUT25), .ZN(new_n272));
  NOR2_X1   g071(.A1(new_n224), .A2(KEYINPUT24), .ZN(new_n273));
  AOI21_X1  g072(.A(new_n232), .B1(G183gat), .B2(G190gat), .ZN(new_n274));
  INV_X1    g073(.A(new_n235), .ZN(new_n275));
  AOI21_X1  g074(.A(new_n273), .B1(new_n274), .B2(new_n275), .ZN(new_n276));
  OAI21_X1  g075(.A(new_n272), .B1(new_n276), .B2(KEYINPUT64), .ZN(new_n277));
  NOR2_X1   g076(.A1(new_n271), .A2(new_n277), .ZN(new_n278));
  NAND2_X1  g077(.A1(new_n225), .A2(new_n237), .ZN(new_n279));
  OAI21_X1  g078(.A(new_n268), .B1(new_n278), .B2(new_n279), .ZN(new_n280));
  AOI21_X1  g079(.A(new_n203), .B1(new_n267), .B2(new_n280), .ZN(new_n281));
  OR2_X1    g080(.A1(new_n281), .A2(KEYINPUT33), .ZN(new_n282));
  XOR2_X1   g081(.A(G15gat), .B(G43gat), .Z(new_n283));
  XNOR2_X1  g082(.A(G71gat), .B(G99gat), .ZN(new_n284));
  XNOR2_X1  g083(.A(new_n283), .B(new_n284), .ZN(new_n285));
  NAND2_X1  g084(.A1(new_n282), .A2(new_n285), .ZN(new_n286));
  INV_X1    g085(.A(KEYINPUT32), .ZN(new_n287));
  OAI21_X1  g086(.A(KEYINPUT34), .B1(new_n281), .B2(new_n287), .ZN(new_n288));
  INV_X1    g087(.A(new_n288), .ZN(new_n289));
  NOR3_X1   g088(.A1(new_n281), .A2(new_n287), .A3(KEYINPUT34), .ZN(new_n290));
  NAND3_X1  g089(.A1(new_n267), .A2(new_n280), .A3(new_n203), .ZN(new_n291));
  INV_X1    g090(.A(new_n291), .ZN(new_n292));
  NOR3_X1   g091(.A1(new_n289), .A2(new_n290), .A3(new_n292), .ZN(new_n293));
  OR3_X1    g092(.A1(new_n281), .A2(new_n287), .A3(KEYINPUT34), .ZN(new_n294));
  AOI21_X1  g093(.A(new_n291), .B1(new_n294), .B2(new_n288), .ZN(new_n295));
  OAI21_X1  g094(.A(new_n286), .B1(new_n293), .B2(new_n295), .ZN(new_n296));
  OAI21_X1  g095(.A(new_n292), .B1(new_n289), .B2(new_n290), .ZN(new_n297));
  NAND3_X1  g096(.A1(new_n294), .A2(new_n291), .A3(new_n288), .ZN(new_n298));
  NAND4_X1  g097(.A1(new_n297), .A2(new_n282), .A3(new_n298), .A4(new_n285), .ZN(new_n299));
  NAND2_X1  g098(.A1(new_n296), .A2(new_n299), .ZN(new_n300));
  INV_X1    g099(.A(KEYINPUT36), .ZN(new_n301));
  NAND2_X1  g100(.A1(new_n300), .A2(new_n301), .ZN(new_n302));
  NAND3_X1  g101(.A1(new_n296), .A2(new_n299), .A3(KEYINPUT36), .ZN(new_n303));
  NAND2_X1  g102(.A1(new_n302), .A2(new_n303), .ZN(new_n304));
  XNOR2_X1  g103(.A(G78gat), .B(G106gat), .ZN(new_n305));
  XNOR2_X1  g104(.A(KEYINPUT31), .B(G50gat), .ZN(new_n306));
  XNOR2_X1  g105(.A(new_n305), .B(new_n306), .ZN(new_n307));
  INV_X1    g106(.A(G228gat), .ZN(new_n308));
  INV_X1    g107(.A(G233gat), .ZN(new_n309));
  NOR2_X1   g108(.A1(new_n308), .A2(new_n309), .ZN(new_n310));
  INV_X1    g109(.A(new_n310), .ZN(new_n311));
  NAND2_X1  g110(.A1(G155gat), .A2(G162gat), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n312), .A2(KEYINPUT2), .ZN(new_n313));
  INV_X1    g112(.A(KEYINPUT75), .ZN(new_n314));
  NAND2_X1  g113(.A1(new_n313), .A2(new_n314), .ZN(new_n315));
  NAND3_X1  g114(.A1(new_n312), .A2(KEYINPUT75), .A3(KEYINPUT2), .ZN(new_n316));
  XNOR2_X1  g115(.A(G155gat), .B(G162gat), .ZN(new_n317));
  AND3_X1   g116(.A1(new_n315), .A2(new_n316), .A3(new_n317), .ZN(new_n318));
  INV_X1    g117(.A(G148gat), .ZN(new_n319));
  NAND2_X1  g118(.A1(new_n319), .A2(G141gat), .ZN(new_n320));
  INV_X1    g119(.A(G141gat), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n321), .A2(G148gat), .ZN(new_n322));
  NAND2_X1  g121(.A1(new_n320), .A2(new_n322), .ZN(new_n323));
  INV_X1    g122(.A(KEYINPUT2), .ZN(new_n324));
  AOI22_X1  g123(.A1(new_n323), .A2(new_n324), .B1(G155gat), .B2(G162gat), .ZN(new_n325));
  NOR2_X1   g124(.A1(G155gat), .A2(G162gat), .ZN(new_n326));
  XNOR2_X1  g125(.A(new_n326), .B(KEYINPUT74), .ZN(new_n327));
  AOI22_X1  g126(.A1(new_n318), .A2(new_n323), .B1(new_n325), .B2(new_n327), .ZN(new_n328));
  XNOR2_X1  g127(.A(G197gat), .B(G204gat), .ZN(new_n329));
  INV_X1    g128(.A(KEYINPUT22), .ZN(new_n330));
  INV_X1    g129(.A(G211gat), .ZN(new_n331));
  INV_X1    g130(.A(G218gat), .ZN(new_n332));
  OAI21_X1  g131(.A(new_n330), .B1(new_n331), .B2(new_n332), .ZN(new_n333));
  NAND2_X1  g132(.A1(new_n329), .A2(new_n333), .ZN(new_n334));
  XNOR2_X1  g133(.A(G211gat), .B(G218gat), .ZN(new_n335));
  INV_X1    g134(.A(new_n335), .ZN(new_n336));
  NAND2_X1  g135(.A1(new_n334), .A2(new_n336), .ZN(new_n337));
  NAND3_X1  g136(.A1(new_n335), .A2(new_n329), .A3(new_n333), .ZN(new_n338));
  NAND2_X1  g137(.A1(new_n337), .A2(new_n338), .ZN(new_n339));
  INV_X1    g138(.A(KEYINPUT29), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n339), .A2(new_n340), .ZN(new_n341));
  INV_X1    g140(.A(KEYINPUT3), .ZN(new_n342));
  AOI21_X1  g141(.A(new_n328), .B1(new_n341), .B2(new_n342), .ZN(new_n343));
  NAND2_X1  g142(.A1(new_n323), .A2(new_n324), .ZN(new_n344));
  NAND3_X1  g143(.A1(new_n327), .A2(new_n344), .A3(new_n312), .ZN(new_n345));
  NAND4_X1  g144(.A1(new_n315), .A2(new_n323), .A3(new_n317), .A4(new_n316), .ZN(new_n346));
  NAND3_X1  g145(.A1(new_n345), .A2(new_n342), .A3(new_n346), .ZN(new_n347));
  INV_X1    g146(.A(KEYINPUT70), .ZN(new_n348));
  NAND3_X1  g147(.A1(new_n337), .A2(new_n348), .A3(new_n338), .ZN(new_n349));
  NAND3_X1  g148(.A1(new_n334), .A2(KEYINPUT70), .A3(new_n336), .ZN(new_n350));
  AOI22_X1  g149(.A1(new_n347), .A2(new_n340), .B1(new_n349), .B2(new_n350), .ZN(new_n351));
  OAI21_X1  g150(.A(new_n311), .B1(new_n343), .B2(new_n351), .ZN(new_n352));
  INV_X1    g151(.A(new_n352), .ZN(new_n353));
  NAND3_X1  g152(.A1(new_n349), .A2(new_n340), .A3(new_n350), .ZN(new_n354));
  AOI21_X1  g153(.A(new_n328), .B1(new_n354), .B2(new_n342), .ZN(new_n355));
  NOR3_X1   g154(.A1(new_n355), .A2(new_n311), .A3(new_n351), .ZN(new_n356));
  NOR3_X1   g155(.A1(new_n353), .A2(new_n356), .A3(G22gat), .ZN(new_n357));
  INV_X1    g156(.A(G22gat), .ZN(new_n358));
  INV_X1    g157(.A(new_n351), .ZN(new_n359));
  AND2_X1   g158(.A1(new_n354), .A2(new_n342), .ZN(new_n360));
  OAI211_X1 g159(.A(new_n359), .B(new_n310), .C1(new_n360), .C2(new_n328), .ZN(new_n361));
  AOI21_X1  g160(.A(new_n358), .B1(new_n361), .B2(new_n352), .ZN(new_n362));
  OAI21_X1  g161(.A(new_n307), .B1(new_n357), .B2(new_n362), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n357), .A2(KEYINPUT78), .ZN(new_n364));
  OAI21_X1  g163(.A(G22gat), .B1(new_n353), .B2(new_n356), .ZN(new_n365));
  NAND3_X1  g164(.A1(new_n361), .A2(new_n352), .A3(new_n358), .ZN(new_n366));
  NOR2_X1   g165(.A1(new_n307), .A2(KEYINPUT78), .ZN(new_n367));
  NAND3_X1  g166(.A1(new_n365), .A2(new_n366), .A3(new_n367), .ZN(new_n368));
  NAND3_X1  g167(.A1(new_n363), .A2(new_n364), .A3(new_n368), .ZN(new_n369));
  NAND2_X1  g168(.A1(new_n369), .A2(KEYINPUT79), .ZN(new_n370));
  INV_X1    g169(.A(KEYINPUT79), .ZN(new_n371));
  NAND4_X1  g170(.A1(new_n363), .A2(new_n364), .A3(new_n371), .A4(new_n368), .ZN(new_n372));
  NAND2_X1  g171(.A1(new_n370), .A2(new_n372), .ZN(new_n373));
  INV_X1    g172(.A(KEYINPUT71), .ZN(new_n374));
  OAI21_X1  g173(.A(new_n374), .B1(new_n278), .B2(new_n279), .ZN(new_n375));
  NAND4_X1  g174(.A1(new_n266), .A2(KEYINPUT71), .A3(new_n237), .A4(new_n225), .ZN(new_n376));
  NAND2_X1  g175(.A1(new_n375), .A2(new_n376), .ZN(new_n377));
  INV_X1    g176(.A(G226gat), .ZN(new_n378));
  NOR2_X1   g177(.A1(new_n378), .A2(new_n309), .ZN(new_n379));
  NOR2_X1   g178(.A1(new_n379), .A2(KEYINPUT29), .ZN(new_n380));
  NAND2_X1  g179(.A1(new_n377), .A2(new_n380), .ZN(new_n381));
  NAND2_X1  g180(.A1(new_n349), .A2(new_n350), .ZN(new_n382));
  INV_X1    g181(.A(new_n379), .ZN(new_n383));
  NOR3_X1   g182(.A1(new_n278), .A2(new_n279), .A3(new_n383), .ZN(new_n384));
  INV_X1    g183(.A(new_n384), .ZN(new_n385));
  NAND3_X1  g184(.A1(new_n381), .A2(new_n382), .A3(new_n385), .ZN(new_n386));
  NAND2_X1  g185(.A1(new_n386), .A2(KEYINPUT72), .ZN(new_n387));
  NAND3_X1  g186(.A1(new_n375), .A2(new_n379), .A3(new_n376), .ZN(new_n388));
  OAI21_X1  g187(.A(new_n380), .B1(new_n278), .B2(new_n279), .ZN(new_n389));
  AOI21_X1  g188(.A(new_n382), .B1(new_n388), .B2(new_n389), .ZN(new_n390));
  INV_X1    g189(.A(new_n390), .ZN(new_n391));
  AOI21_X1  g190(.A(new_n384), .B1(new_n377), .B2(new_n380), .ZN(new_n392));
  INV_X1    g191(.A(KEYINPUT72), .ZN(new_n393));
  NAND3_X1  g192(.A1(new_n392), .A2(new_n393), .A3(new_n382), .ZN(new_n394));
  NAND3_X1  g193(.A1(new_n387), .A2(new_n391), .A3(new_n394), .ZN(new_n395));
  XNOR2_X1  g194(.A(G64gat), .B(G92gat), .ZN(new_n396));
  INV_X1    g195(.A(G36gat), .ZN(new_n397));
  XNOR2_X1  g196(.A(new_n396), .B(new_n397), .ZN(new_n398));
  XNOR2_X1  g197(.A(KEYINPUT73), .B(G8gat), .ZN(new_n399));
  XOR2_X1   g198(.A(new_n398), .B(new_n399), .Z(new_n400));
  NAND2_X1  g199(.A1(new_n395), .A2(new_n400), .ZN(new_n401));
  INV_X1    g200(.A(new_n400), .ZN(new_n402));
  NAND4_X1  g201(.A1(new_n387), .A2(new_n402), .A3(new_n391), .A4(new_n394), .ZN(new_n403));
  NAND3_X1  g202(.A1(new_n401), .A2(KEYINPUT30), .A3(new_n403), .ZN(new_n404));
  AOI21_X1  g203(.A(new_n393), .B1(new_n392), .B2(new_n382), .ZN(new_n405));
  INV_X1    g204(.A(new_n380), .ZN(new_n406));
  AOI21_X1  g205(.A(new_n406), .B1(new_n375), .B2(new_n376), .ZN(new_n407));
  INV_X1    g206(.A(new_n382), .ZN(new_n408));
  NOR4_X1   g207(.A1(new_n407), .A2(KEYINPUT72), .A3(new_n408), .A4(new_n384), .ZN(new_n409));
  NOR3_X1   g208(.A1(new_n405), .A2(new_n409), .A3(new_n390), .ZN(new_n410));
  INV_X1    g209(.A(KEYINPUT30), .ZN(new_n411));
  NAND3_X1  g210(.A1(new_n410), .A2(new_n411), .A3(new_n402), .ZN(new_n412));
  NAND2_X1  g211(.A1(G225gat), .A2(G233gat), .ZN(new_n413));
  INV_X1    g212(.A(new_n413), .ZN(new_n414));
  XNOR2_X1  g213(.A(G141gat), .B(G148gat), .ZN(new_n415));
  OAI21_X1  g214(.A(new_n312), .B1(new_n415), .B2(KEYINPUT2), .ZN(new_n416));
  INV_X1    g215(.A(KEYINPUT74), .ZN(new_n417));
  XNOR2_X1  g216(.A(new_n326), .B(new_n417), .ZN(new_n418));
  OAI21_X1  g217(.A(new_n346), .B1(new_n416), .B2(new_n418), .ZN(new_n419));
  NOR2_X1   g218(.A1(new_n419), .A2(new_n268), .ZN(new_n420));
  AOI22_X1  g219(.A1(new_n345), .A2(new_n346), .B1(new_n246), .B2(new_n256), .ZN(new_n421));
  OAI21_X1  g220(.A(new_n414), .B1(new_n420), .B2(new_n421), .ZN(new_n422));
  INV_X1    g221(.A(KEYINPUT76), .ZN(new_n423));
  NAND3_X1  g222(.A1(new_n422), .A2(new_n423), .A3(KEYINPUT5), .ZN(new_n424));
  NAND2_X1  g223(.A1(new_n419), .A2(new_n268), .ZN(new_n425));
  NAND4_X1  g224(.A1(new_n345), .A2(new_n256), .A3(new_n246), .A4(new_n346), .ZN(new_n426));
  AOI21_X1  g225(.A(new_n413), .B1(new_n425), .B2(new_n426), .ZN(new_n427));
  INV_X1    g226(.A(KEYINPUT5), .ZN(new_n428));
  OAI21_X1  g227(.A(KEYINPUT76), .B1(new_n427), .B2(new_n428), .ZN(new_n429));
  NAND2_X1  g228(.A1(new_n419), .A2(KEYINPUT3), .ZN(new_n430));
  NAND3_X1  g229(.A1(new_n430), .A2(new_n268), .A3(new_n347), .ZN(new_n431));
  NAND3_X1  g230(.A1(new_n328), .A2(new_n257), .A3(KEYINPUT4), .ZN(new_n432));
  INV_X1    g231(.A(KEYINPUT4), .ZN(new_n433));
  NAND2_X1  g232(.A1(new_n426), .A2(new_n433), .ZN(new_n434));
  NAND4_X1  g233(.A1(new_n431), .A2(new_n413), .A3(new_n432), .A4(new_n434), .ZN(new_n435));
  NAND3_X1  g234(.A1(new_n424), .A2(new_n429), .A3(new_n435), .ZN(new_n436));
  OAI21_X1  g235(.A(KEYINPUT77), .B1(new_n435), .B2(KEYINPUT5), .ZN(new_n437));
  NAND2_X1  g236(.A1(new_n436), .A2(new_n437), .ZN(new_n438));
  NAND4_X1  g237(.A1(new_n424), .A2(new_n429), .A3(KEYINPUT77), .A4(new_n435), .ZN(new_n439));
  NAND2_X1  g238(.A1(new_n438), .A2(new_n439), .ZN(new_n440));
  XNOR2_X1  g239(.A(G1gat), .B(G29gat), .ZN(new_n441));
  XNOR2_X1  g240(.A(new_n441), .B(G85gat), .ZN(new_n442));
  XNOR2_X1  g241(.A(KEYINPUT0), .B(G57gat), .ZN(new_n443));
  XOR2_X1   g242(.A(new_n442), .B(new_n443), .Z(new_n444));
  INV_X1    g243(.A(new_n444), .ZN(new_n445));
  NAND3_X1  g244(.A1(new_n440), .A2(KEYINPUT6), .A3(new_n445), .ZN(new_n446));
  NAND2_X1  g245(.A1(new_n440), .A2(new_n445), .ZN(new_n447));
  INV_X1    g246(.A(KEYINPUT6), .ZN(new_n448));
  NAND3_X1  g247(.A1(new_n438), .A2(new_n444), .A3(new_n439), .ZN(new_n449));
  NAND3_X1  g248(.A1(new_n447), .A2(new_n448), .A3(new_n449), .ZN(new_n450));
  AOI22_X1  g249(.A1(new_n404), .A2(new_n412), .B1(new_n446), .B2(new_n450), .ZN(new_n451));
  OAI21_X1  g250(.A(new_n304), .B1(new_n373), .B2(new_n451), .ZN(new_n452));
  NAND3_X1  g251(.A1(new_n440), .A2(KEYINPUT6), .A3(new_n445), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n449), .A2(new_n448), .ZN(new_n454));
  XOR2_X1   g253(.A(new_n444), .B(KEYINPUT80), .Z(new_n455));
  AOI21_X1  g254(.A(new_n455), .B1(new_n438), .B2(new_n439), .ZN(new_n456));
  OAI211_X1 g255(.A(new_n403), .B(new_n453), .C1(new_n454), .C2(new_n456), .ZN(new_n457));
  INV_X1    g256(.A(new_n457), .ZN(new_n458));
  INV_X1    g257(.A(KEYINPUT37), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n388), .A2(new_n389), .ZN(new_n460));
  AOI21_X1  g259(.A(new_n459), .B1(new_n460), .B2(new_n382), .ZN(new_n461));
  INV_X1    g260(.A(KEYINPUT82), .ZN(new_n462));
  NAND3_X1  g261(.A1(new_n381), .A2(new_n408), .A3(new_n385), .ZN(new_n463));
  AND3_X1   g262(.A1(new_n461), .A2(new_n462), .A3(new_n463), .ZN(new_n464));
  AOI21_X1  g263(.A(new_n462), .B1(new_n461), .B2(new_n463), .ZN(new_n465));
  NOR3_X1   g264(.A1(new_n464), .A2(new_n465), .A3(KEYINPUT38), .ZN(new_n466));
  AOI21_X1  g265(.A(new_n402), .B1(new_n410), .B2(new_n459), .ZN(new_n467));
  NAND3_X1  g266(.A1(new_n466), .A2(new_n467), .A3(KEYINPUT83), .ZN(new_n468));
  INV_X1    g267(.A(KEYINPUT83), .ZN(new_n469));
  NAND2_X1  g268(.A1(new_n460), .A2(new_n382), .ZN(new_n470));
  NAND3_X1  g269(.A1(new_n463), .A2(new_n470), .A3(KEYINPUT37), .ZN(new_n471));
  NAND2_X1  g270(.A1(new_n471), .A2(KEYINPUT82), .ZN(new_n472));
  INV_X1    g271(.A(KEYINPUT38), .ZN(new_n473));
  NAND3_X1  g272(.A1(new_n461), .A2(new_n462), .A3(new_n463), .ZN(new_n474));
  NAND3_X1  g273(.A1(new_n472), .A2(new_n473), .A3(new_n474), .ZN(new_n475));
  NAND4_X1  g274(.A1(new_n387), .A2(new_n459), .A3(new_n391), .A4(new_n394), .ZN(new_n476));
  NAND2_X1  g275(.A1(new_n476), .A2(new_n400), .ZN(new_n477));
  OAI21_X1  g276(.A(new_n469), .B1(new_n475), .B2(new_n477), .ZN(new_n478));
  NAND3_X1  g277(.A1(new_n458), .A2(new_n468), .A3(new_n478), .ZN(new_n479));
  INV_X1    g278(.A(KEYINPUT84), .ZN(new_n480));
  NAND2_X1  g279(.A1(new_n479), .A2(new_n480), .ZN(new_n481));
  NOR2_X1   g280(.A1(new_n410), .A2(new_n459), .ZN(new_n482));
  OAI21_X1  g281(.A(KEYINPUT38), .B1(new_n482), .B2(new_n477), .ZN(new_n483));
  NAND4_X1  g282(.A1(new_n458), .A2(new_n468), .A3(new_n478), .A4(KEYINPUT84), .ZN(new_n484));
  NAND3_X1  g283(.A1(new_n481), .A2(new_n483), .A3(new_n484), .ZN(new_n485));
  INV_X1    g284(.A(new_n373), .ZN(new_n486));
  NAND2_X1  g285(.A1(new_n404), .A2(new_n412), .ZN(new_n487));
  INV_X1    g286(.A(new_n487), .ZN(new_n488));
  NAND3_X1  g287(.A1(new_n431), .A2(new_n434), .A3(new_n432), .ZN(new_n489));
  NAND2_X1  g288(.A1(new_n489), .A2(new_n414), .ZN(new_n490));
  NAND3_X1  g289(.A1(new_n425), .A2(new_n413), .A3(new_n426), .ZN(new_n491));
  NAND3_X1  g290(.A1(new_n490), .A2(KEYINPUT39), .A3(new_n491), .ZN(new_n492));
  OAI211_X1 g291(.A(new_n492), .B(new_n455), .C1(KEYINPUT39), .C2(new_n490), .ZN(new_n493));
  INV_X1    g292(.A(KEYINPUT81), .ZN(new_n494));
  INV_X1    g293(.A(KEYINPUT40), .ZN(new_n495));
  NAND3_X1  g294(.A1(new_n493), .A2(new_n494), .A3(new_n495), .ZN(new_n496));
  OAI21_X1  g295(.A(new_n496), .B1(new_n495), .B2(new_n493), .ZN(new_n497));
  AOI21_X1  g296(.A(new_n494), .B1(new_n493), .B2(new_n495), .ZN(new_n498));
  NOR3_X1   g297(.A1(new_n497), .A2(new_n498), .A3(new_n456), .ZN(new_n499));
  AOI21_X1  g298(.A(new_n486), .B1(new_n488), .B2(new_n499), .ZN(new_n500));
  AOI21_X1  g299(.A(new_n452), .B1(new_n485), .B2(new_n500), .ZN(new_n501));
  INV_X1    g300(.A(new_n300), .ZN(new_n502));
  NAND3_X1  g301(.A1(new_n451), .A2(new_n502), .A3(new_n373), .ZN(new_n503));
  NAND2_X1  g302(.A1(new_n503), .A2(KEYINPUT35), .ZN(new_n504));
  AND2_X1   g303(.A1(new_n438), .A2(new_n439), .ZN(new_n505));
  OAI211_X1 g304(.A(new_n448), .B(new_n449), .C1(new_n505), .C2(new_n455), .ZN(new_n506));
  AOI21_X1  g305(.A(KEYINPUT35), .B1(new_n506), .B2(new_n453), .ZN(new_n507));
  NAND4_X1  g306(.A1(new_n487), .A2(new_n502), .A3(new_n373), .A4(new_n507), .ZN(new_n508));
  NAND2_X1  g307(.A1(new_n508), .A2(KEYINPUT85), .ZN(new_n509));
  AOI21_X1  g308(.A(new_n300), .B1(new_n372), .B2(new_n370), .ZN(new_n510));
  INV_X1    g309(.A(KEYINPUT85), .ZN(new_n511));
  NAND4_X1  g310(.A1(new_n510), .A2(new_n511), .A3(new_n487), .A4(new_n507), .ZN(new_n512));
  AND3_X1   g311(.A1(new_n504), .A2(new_n509), .A3(new_n512), .ZN(new_n513));
  OR2_X1    g312(.A1(new_n501), .A2(new_n513), .ZN(new_n514));
  INV_X1    g313(.A(KEYINPUT14), .ZN(new_n515));
  INV_X1    g314(.A(G29gat), .ZN(new_n516));
  NAND3_X1  g315(.A1(new_n515), .A2(new_n516), .A3(new_n397), .ZN(new_n517));
  INV_X1    g316(.A(KEYINPUT87), .ZN(new_n518));
  OAI21_X1  g317(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n519));
  NAND3_X1  g318(.A1(new_n517), .A2(new_n518), .A3(new_n519), .ZN(new_n520));
  OAI211_X1 g319(.A(KEYINPUT87), .B(KEYINPUT14), .C1(G29gat), .C2(G36gat), .ZN(new_n521));
  OAI211_X1 g320(.A(new_n520), .B(new_n521), .C1(new_n516), .C2(new_n397), .ZN(new_n522));
  XNOR2_X1  g321(.A(G43gat), .B(G50gat), .ZN(new_n523));
  NAND3_X1  g322(.A1(new_n522), .A2(KEYINPUT15), .A3(new_n523), .ZN(new_n524));
  INV_X1    g323(.A(G50gat), .ZN(new_n525));
  NAND2_X1  g324(.A1(new_n525), .A2(G43gat), .ZN(new_n526));
  INV_X1    g325(.A(G43gat), .ZN(new_n527));
  NAND2_X1  g326(.A1(new_n527), .A2(G50gat), .ZN(new_n528));
  NAND2_X1  g327(.A1(new_n526), .A2(new_n528), .ZN(new_n529));
  INV_X1    g328(.A(KEYINPUT15), .ZN(new_n530));
  AOI22_X1  g329(.A1(new_n529), .A2(new_n530), .B1(G29gat), .B2(G36gat), .ZN(new_n531));
  AOI22_X1  g330(.A1(new_n523), .A2(KEYINPUT15), .B1(new_n517), .B2(new_n519), .ZN(new_n532));
  AND3_X1   g331(.A1(new_n531), .A2(new_n532), .A3(KEYINPUT88), .ZN(new_n533));
  AOI21_X1  g332(.A(KEYINPUT88), .B1(new_n531), .B2(new_n532), .ZN(new_n534));
  OAI21_X1  g333(.A(new_n524), .B1(new_n533), .B2(new_n534), .ZN(new_n535));
  INV_X1    g334(.A(KEYINPUT17), .ZN(new_n536));
  NAND2_X1  g335(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  XOR2_X1   g336(.A(G15gat), .B(G22gat), .Z(new_n538));
  INV_X1    g337(.A(G1gat), .ZN(new_n539));
  NAND2_X1  g338(.A1(new_n538), .A2(new_n539), .ZN(new_n540));
  INV_X1    g339(.A(KEYINPUT89), .ZN(new_n541));
  XNOR2_X1  g340(.A(G15gat), .B(G22gat), .ZN(new_n542));
  NAND2_X1  g341(.A1(new_n539), .A2(KEYINPUT16), .ZN(new_n543));
  AOI21_X1  g342(.A(new_n541), .B1(new_n542), .B2(new_n543), .ZN(new_n544));
  NAND2_X1  g343(.A1(new_n540), .A2(new_n544), .ZN(new_n545));
  NAND2_X1  g344(.A1(new_n545), .A2(G8gat), .ZN(new_n546));
  INV_X1    g345(.A(KEYINPUT90), .ZN(new_n547));
  INV_X1    g346(.A(G8gat), .ZN(new_n548));
  NAND3_X1  g347(.A1(new_n540), .A2(new_n544), .A3(new_n548), .ZN(new_n549));
  NAND3_X1  g348(.A1(new_n546), .A2(new_n547), .A3(new_n549), .ZN(new_n550));
  OAI211_X1 g349(.A(new_n524), .B(KEYINPUT17), .C1(new_n533), .C2(new_n534), .ZN(new_n551));
  NAND2_X1  g350(.A1(new_n546), .A2(new_n549), .ZN(new_n552));
  NAND2_X1  g351(.A1(new_n552), .A2(KEYINPUT90), .ZN(new_n553));
  NAND4_X1  g352(.A1(new_n537), .A2(new_n550), .A3(new_n551), .A4(new_n553), .ZN(new_n554));
  NAND2_X1  g353(.A1(new_n535), .A2(new_n552), .ZN(new_n555));
  NAND2_X1  g354(.A1(G229gat), .A2(G233gat), .ZN(new_n556));
  NAND3_X1  g355(.A1(new_n554), .A2(new_n555), .A3(new_n556), .ZN(new_n557));
  NOR2_X1   g356(.A1(KEYINPUT91), .A2(KEYINPUT18), .ZN(new_n558));
  INV_X1    g357(.A(new_n558), .ZN(new_n559));
  NAND2_X1  g358(.A1(new_n557), .A2(new_n559), .ZN(new_n560));
  NAND4_X1  g359(.A1(new_n554), .A2(new_n555), .A3(new_n556), .A4(new_n558), .ZN(new_n561));
  NAND2_X1  g360(.A1(new_n560), .A2(new_n561), .ZN(new_n562));
  OR2_X1    g361(.A1(new_n535), .A2(new_n552), .ZN(new_n563));
  NAND2_X1  g362(.A1(new_n563), .A2(new_n555), .ZN(new_n564));
  XNOR2_X1  g363(.A(KEYINPUT92), .B(KEYINPUT13), .ZN(new_n565));
  XNOR2_X1  g364(.A(new_n565), .B(new_n556), .ZN(new_n566));
  INV_X1    g365(.A(new_n566), .ZN(new_n567));
  AOI21_X1  g366(.A(KEYINPUT93), .B1(new_n564), .B2(new_n567), .ZN(new_n568));
  INV_X1    g367(.A(KEYINPUT93), .ZN(new_n569));
  AOI211_X1 g368(.A(new_n569), .B(new_n566), .C1(new_n563), .C2(new_n555), .ZN(new_n570));
  NOR2_X1   g369(.A1(new_n568), .A2(new_n570), .ZN(new_n571));
  NAND2_X1  g370(.A1(new_n562), .A2(new_n571), .ZN(new_n572));
  XNOR2_X1  g371(.A(KEYINPUT86), .B(KEYINPUT11), .ZN(new_n573));
  XNOR2_X1  g372(.A(G169gat), .B(G197gat), .ZN(new_n574));
  XNOR2_X1  g373(.A(new_n573), .B(new_n574), .ZN(new_n575));
  XNOR2_X1  g374(.A(G113gat), .B(G141gat), .ZN(new_n576));
  XNOR2_X1  g375(.A(new_n575), .B(new_n576), .ZN(new_n577));
  XNOR2_X1  g376(.A(new_n577), .B(KEYINPUT12), .ZN(new_n578));
  NAND2_X1  g377(.A1(new_n572), .A2(new_n578), .ZN(new_n579));
  INV_X1    g378(.A(new_n578), .ZN(new_n580));
  NAND3_X1  g379(.A1(new_n562), .A2(new_n571), .A3(new_n580), .ZN(new_n581));
  NAND2_X1  g380(.A1(new_n579), .A2(new_n581), .ZN(new_n582));
  INV_X1    g381(.A(new_n582), .ZN(new_n583));
  XOR2_X1   g382(.A(G57gat), .B(G64gat), .Z(new_n584));
  AOI21_X1  g383(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n585));
  INV_X1    g384(.A(KEYINPUT94), .ZN(new_n586));
  AND2_X1   g385(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  NOR2_X1   g386(.A1(new_n585), .A2(new_n586), .ZN(new_n588));
  OAI21_X1  g387(.A(new_n584), .B1(new_n587), .B2(new_n588), .ZN(new_n589));
  INV_X1    g388(.A(KEYINPUT95), .ZN(new_n590));
  OR2_X1    g389(.A1(G71gat), .A2(G78gat), .ZN(new_n591));
  NAND2_X1  g390(.A1(G71gat), .A2(G78gat), .ZN(new_n592));
  NAND2_X1  g391(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  NAND3_X1  g392(.A1(new_n589), .A2(new_n590), .A3(new_n593), .ZN(new_n594));
  XNOR2_X1  g393(.A(new_n585), .B(new_n586), .ZN(new_n595));
  NAND2_X1  g394(.A1(new_n593), .A2(new_n590), .ZN(new_n596));
  NAND3_X1  g395(.A1(new_n591), .A2(KEYINPUT95), .A3(new_n592), .ZN(new_n597));
  NAND4_X1  g396(.A1(new_n595), .A2(new_n596), .A3(new_n597), .A4(new_n584), .ZN(new_n598));
  NAND2_X1  g397(.A1(new_n594), .A2(new_n598), .ZN(new_n599));
  OR2_X1    g398(.A1(G99gat), .A2(G106gat), .ZN(new_n600));
  INV_X1    g399(.A(KEYINPUT98), .ZN(new_n601));
  NAND2_X1  g400(.A1(G99gat), .A2(G106gat), .ZN(new_n602));
  NAND3_X1  g401(.A1(new_n600), .A2(new_n601), .A3(new_n602), .ZN(new_n603));
  AND2_X1   g402(.A1(G99gat), .A2(G106gat), .ZN(new_n604));
  NOR2_X1   g403(.A1(G99gat), .A2(G106gat), .ZN(new_n605));
  OAI21_X1  g404(.A(KEYINPUT98), .B1(new_n604), .B2(new_n605), .ZN(new_n606));
  NAND2_X1  g405(.A1(new_n603), .A2(new_n606), .ZN(new_n607));
  INV_X1    g406(.A(G85gat), .ZN(new_n608));
  INV_X1    g407(.A(G92gat), .ZN(new_n609));
  AOI22_X1  g408(.A1(KEYINPUT8), .A2(new_n602), .B1(new_n608), .B2(new_n609), .ZN(new_n610));
  INV_X1    g409(.A(KEYINPUT7), .ZN(new_n611));
  OAI211_X1 g410(.A(KEYINPUT97), .B(new_n611), .C1(new_n608), .C2(new_n609), .ZN(new_n612));
  OAI21_X1  g411(.A(KEYINPUT97), .B1(new_n608), .B2(new_n609), .ZN(new_n613));
  INV_X1    g412(.A(KEYINPUT97), .ZN(new_n614));
  NAND3_X1  g413(.A1(new_n614), .A2(G85gat), .A3(G92gat), .ZN(new_n615));
  NAND3_X1  g414(.A1(new_n613), .A2(new_n615), .A3(KEYINPUT7), .ZN(new_n616));
  NAND4_X1  g415(.A1(new_n607), .A2(new_n610), .A3(new_n612), .A4(new_n616), .ZN(new_n617));
  NAND3_X1  g416(.A1(new_n616), .A2(new_n610), .A3(new_n612), .ZN(new_n618));
  AND2_X1   g417(.A1(new_n603), .A2(new_n606), .ZN(new_n619));
  NAND2_X1  g418(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  NAND3_X1  g419(.A1(new_n599), .A2(new_n617), .A3(new_n620), .ZN(new_n621));
  INV_X1    g420(.A(KEYINPUT10), .ZN(new_n622));
  NAND3_X1  g421(.A1(new_n620), .A2(KEYINPUT99), .A3(new_n617), .ZN(new_n623));
  AND2_X1   g422(.A1(new_n616), .A2(new_n612), .ZN(new_n624));
  INV_X1    g423(.A(KEYINPUT99), .ZN(new_n625));
  NAND4_X1  g424(.A1(new_n624), .A2(new_n625), .A3(new_n607), .A4(new_n610), .ZN(new_n626));
  NAND2_X1  g425(.A1(new_n623), .A2(new_n626), .ZN(new_n627));
  OAI211_X1 g426(.A(new_n621), .B(new_n622), .C1(new_n627), .C2(new_n599), .ZN(new_n628));
  NAND3_X1  g427(.A1(new_n627), .A2(KEYINPUT10), .A3(new_n599), .ZN(new_n629));
  NAND2_X1  g428(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  NAND2_X1  g429(.A1(G230gat), .A2(G233gat), .ZN(new_n631));
  XOR2_X1   g430(.A(new_n631), .B(KEYINPUT101), .Z(new_n632));
  INV_X1    g431(.A(new_n632), .ZN(new_n633));
  NAND2_X1  g432(.A1(new_n630), .A2(new_n633), .ZN(new_n634));
  OAI21_X1  g433(.A(new_n621), .B1(new_n627), .B2(new_n599), .ZN(new_n635));
  NAND2_X1  g434(.A1(new_n635), .A2(new_n632), .ZN(new_n636));
  NAND2_X1  g435(.A1(new_n634), .A2(new_n636), .ZN(new_n637));
  XNOR2_X1  g436(.A(G120gat), .B(G148gat), .ZN(new_n638));
  XNOR2_X1  g437(.A(G176gat), .B(G204gat), .ZN(new_n639));
  XNOR2_X1  g438(.A(new_n638), .B(new_n639), .ZN(new_n640));
  NAND2_X1  g439(.A1(new_n637), .A2(new_n640), .ZN(new_n641));
  INV_X1    g440(.A(new_n640), .ZN(new_n642));
  NAND3_X1  g441(.A1(new_n634), .A2(new_n636), .A3(new_n642), .ZN(new_n643));
  NAND2_X1  g442(.A1(new_n641), .A2(new_n643), .ZN(new_n644));
  NOR2_X1   g443(.A1(new_n583), .A2(new_n644), .ZN(new_n645));
  AOI21_X1  g444(.A(new_n552), .B1(KEYINPUT21), .B2(new_n599), .ZN(new_n646));
  XNOR2_X1  g445(.A(new_n646), .B(KEYINPUT96), .ZN(new_n647));
  NOR2_X1   g446(.A1(new_n599), .A2(KEYINPUT21), .ZN(new_n648));
  INV_X1    g447(.A(new_n648), .ZN(new_n649));
  NOR2_X1   g448(.A1(new_n647), .A2(new_n649), .ZN(new_n650));
  INV_X1    g449(.A(new_n650), .ZN(new_n651));
  NAND2_X1  g450(.A1(new_n647), .A2(new_n649), .ZN(new_n652));
  NAND4_X1  g451(.A1(new_n651), .A2(G231gat), .A3(G233gat), .A4(new_n652), .ZN(new_n653));
  INV_X1    g452(.A(new_n652), .ZN(new_n654));
  INV_X1    g453(.A(G231gat), .ZN(new_n655));
  OAI22_X1  g454(.A1(new_n654), .A2(new_n650), .B1(new_n655), .B2(new_n309), .ZN(new_n656));
  NAND2_X1  g455(.A1(new_n653), .A2(new_n656), .ZN(new_n657));
  XNOR2_X1  g456(.A(G183gat), .B(G211gat), .ZN(new_n658));
  XNOR2_X1  g457(.A(new_n658), .B(new_n239), .ZN(new_n659));
  NAND2_X1  g458(.A1(new_n657), .A2(new_n659), .ZN(new_n660));
  INV_X1    g459(.A(new_n659), .ZN(new_n661));
  NAND3_X1  g460(.A1(new_n653), .A2(new_n656), .A3(new_n661), .ZN(new_n662));
  NAND2_X1  g461(.A1(new_n660), .A2(new_n662), .ZN(new_n663));
  XNOR2_X1  g462(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n664));
  XNOR2_X1  g463(.A(new_n664), .B(G155gat), .ZN(new_n665));
  INV_X1    g464(.A(new_n665), .ZN(new_n666));
  NAND2_X1  g465(.A1(new_n663), .A2(new_n666), .ZN(new_n667));
  NAND3_X1  g466(.A1(new_n660), .A2(new_n665), .A3(new_n662), .ZN(new_n668));
  AND2_X1   g467(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  AND2_X1   g468(.A1(new_n623), .A2(new_n626), .ZN(new_n670));
  NAND3_X1  g469(.A1(new_n537), .A2(new_n670), .A3(new_n551), .ZN(new_n671));
  NAND3_X1  g470(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n672));
  NAND2_X1  g471(.A1(new_n627), .A2(new_n535), .ZN(new_n673));
  XOR2_X1   g472(.A(G190gat), .B(G218gat), .Z(new_n674));
  INV_X1    g473(.A(KEYINPUT100), .ZN(new_n675));
  NOR2_X1   g474(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  INV_X1    g475(.A(new_n676), .ZN(new_n677));
  NAND4_X1  g476(.A1(new_n671), .A2(new_n672), .A3(new_n673), .A4(new_n677), .ZN(new_n678));
  XNOR2_X1  g477(.A(G134gat), .B(G162gat), .ZN(new_n679));
  NAND2_X1  g478(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  INV_X1    g479(.A(new_n680), .ZN(new_n681));
  NOR2_X1   g480(.A1(new_n678), .A2(new_n679), .ZN(new_n682));
  NAND2_X1  g481(.A1(new_n674), .A2(new_n675), .ZN(new_n683));
  AOI21_X1  g482(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n684));
  XOR2_X1   g483(.A(new_n683), .B(new_n684), .Z(new_n685));
  INV_X1    g484(.A(new_n685), .ZN(new_n686));
  NOR3_X1   g485(.A1(new_n681), .A2(new_n682), .A3(new_n686), .ZN(new_n687));
  OR2_X1    g486(.A1(new_n678), .A2(new_n679), .ZN(new_n688));
  AOI21_X1  g487(.A(new_n685), .B1(new_n688), .B2(new_n680), .ZN(new_n689));
  NOR2_X1   g488(.A1(new_n687), .A2(new_n689), .ZN(new_n690));
  NOR2_X1   g489(.A1(new_n669), .A2(new_n690), .ZN(new_n691));
  NAND3_X1  g490(.A1(new_n514), .A2(new_n645), .A3(new_n691), .ZN(new_n692));
  XNOR2_X1  g491(.A(new_n692), .B(KEYINPUT102), .ZN(new_n693));
  NAND2_X1  g492(.A1(new_n450), .A2(new_n446), .ZN(new_n694));
  INV_X1    g493(.A(new_n694), .ZN(new_n695));
  NAND2_X1  g494(.A1(new_n693), .A2(new_n695), .ZN(new_n696));
  XNOR2_X1  g495(.A(new_n696), .B(G1gat), .ZN(G1324gat));
  OR2_X1    g496(.A1(new_n692), .A2(KEYINPUT102), .ZN(new_n698));
  NAND2_X1  g497(.A1(new_n692), .A2(KEYINPUT102), .ZN(new_n699));
  AOI21_X1  g498(.A(new_n487), .B1(new_n698), .B2(new_n699), .ZN(new_n700));
  NAND2_X1  g499(.A1(KEYINPUT16), .A2(G8gat), .ZN(new_n701));
  OR2_X1    g500(.A1(KEYINPUT16), .A2(G8gat), .ZN(new_n702));
  NAND3_X1  g501(.A1(new_n700), .A2(new_n701), .A3(new_n702), .ZN(new_n703));
  INV_X1    g502(.A(KEYINPUT42), .ZN(new_n704));
  NAND2_X1  g503(.A1(new_n703), .A2(new_n704), .ZN(new_n705));
  OR2_X1    g504(.A1(new_n700), .A2(new_n548), .ZN(new_n706));
  NAND4_X1  g505(.A1(new_n700), .A2(KEYINPUT42), .A3(new_n701), .A4(new_n702), .ZN(new_n707));
  NAND3_X1  g506(.A1(new_n705), .A2(new_n706), .A3(new_n707), .ZN(G1325gat));
  AOI21_X1  g507(.A(G15gat), .B1(new_n693), .B2(new_n502), .ZN(new_n709));
  AOI21_X1  g508(.A(new_n304), .B1(new_n698), .B2(new_n699), .ZN(new_n710));
  AOI21_X1  g509(.A(new_n709), .B1(G15gat), .B2(new_n710), .ZN(G1326gat));
  NAND2_X1  g510(.A1(new_n693), .A2(new_n486), .ZN(new_n712));
  NAND2_X1  g511(.A1(new_n712), .A2(G22gat), .ZN(new_n713));
  XNOR2_X1  g512(.A(KEYINPUT103), .B(KEYINPUT43), .ZN(new_n714));
  NAND3_X1  g513(.A1(new_n693), .A2(new_n358), .A3(new_n486), .ZN(new_n715));
  NAND3_X1  g514(.A1(new_n713), .A2(new_n714), .A3(new_n715), .ZN(new_n716));
  INV_X1    g515(.A(new_n714), .ZN(new_n717));
  AOI211_X1 g516(.A(G22gat), .B(new_n373), .C1(new_n698), .C2(new_n699), .ZN(new_n718));
  AOI21_X1  g517(.A(new_n358), .B1(new_n693), .B2(new_n486), .ZN(new_n719));
  OAI21_X1  g518(.A(new_n717), .B1(new_n718), .B2(new_n719), .ZN(new_n720));
  NAND2_X1  g519(.A1(new_n716), .A2(new_n720), .ZN(G1327gat));
  OAI21_X1  g520(.A(new_n690), .B1(new_n501), .B2(new_n513), .ZN(new_n722));
  INV_X1    g521(.A(KEYINPUT44), .ZN(new_n723));
  NAND2_X1  g522(.A1(new_n722), .A2(new_n723), .ZN(new_n724));
  OAI211_X1 g523(.A(KEYINPUT44), .B(new_n690), .C1(new_n501), .C2(new_n513), .ZN(new_n725));
  AND2_X1   g524(.A1(new_n724), .A2(new_n725), .ZN(new_n726));
  NAND2_X1  g525(.A1(new_n669), .A2(new_n645), .ZN(new_n727));
  INV_X1    g526(.A(new_n727), .ZN(new_n728));
  NAND3_X1  g527(.A1(new_n726), .A2(new_n695), .A3(new_n728), .ZN(new_n729));
  NAND2_X1  g528(.A1(new_n729), .A2(G29gat), .ZN(new_n730));
  INV_X1    g529(.A(KEYINPUT45), .ZN(new_n731));
  NAND3_X1  g530(.A1(new_n514), .A2(new_n690), .A3(new_n728), .ZN(new_n732));
  NOR2_X1   g531(.A1(new_n732), .A2(G29gat), .ZN(new_n733));
  AOI21_X1  g532(.A(new_n731), .B1(new_n733), .B2(new_n695), .ZN(new_n734));
  NOR4_X1   g533(.A1(new_n732), .A2(KEYINPUT45), .A3(G29gat), .A4(new_n694), .ZN(new_n735));
  OAI21_X1  g534(.A(new_n730), .B1(new_n734), .B2(new_n735), .ZN(new_n736));
  NAND2_X1  g535(.A1(new_n736), .A2(KEYINPUT104), .ZN(new_n737));
  INV_X1    g536(.A(KEYINPUT104), .ZN(new_n738));
  OAI211_X1 g537(.A(new_n730), .B(new_n738), .C1(new_n734), .C2(new_n735), .ZN(new_n739));
  NAND2_X1  g538(.A1(new_n737), .A2(new_n739), .ZN(G1328gat));
  NOR3_X1   g539(.A1(new_n732), .A2(G36gat), .A3(new_n487), .ZN(new_n741));
  INV_X1    g540(.A(KEYINPUT46), .ZN(new_n742));
  OR2_X1    g541(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  NAND3_X1  g542(.A1(new_n726), .A2(new_n488), .A3(new_n728), .ZN(new_n744));
  NAND2_X1  g543(.A1(new_n744), .A2(G36gat), .ZN(new_n745));
  NAND2_X1  g544(.A1(new_n741), .A2(new_n742), .ZN(new_n746));
  NAND3_X1  g545(.A1(new_n743), .A2(new_n745), .A3(new_n746), .ZN(new_n747));
  INV_X1    g546(.A(KEYINPUT105), .ZN(new_n748));
  NAND2_X1  g547(.A1(new_n747), .A2(new_n748), .ZN(new_n749));
  NAND4_X1  g548(.A1(new_n743), .A2(new_n745), .A3(KEYINPUT105), .A4(new_n746), .ZN(new_n750));
  NAND2_X1  g549(.A1(new_n749), .A2(new_n750), .ZN(G1329gat));
  INV_X1    g550(.A(new_n304), .ZN(new_n752));
  NAND4_X1  g551(.A1(new_n724), .A2(new_n752), .A3(new_n725), .A4(new_n728), .ZN(new_n753));
  INV_X1    g552(.A(KEYINPUT106), .ZN(new_n754));
  OR2_X1    g553(.A1(new_n753), .A2(new_n754), .ZN(new_n755));
  NAND2_X1  g554(.A1(new_n753), .A2(new_n754), .ZN(new_n756));
  NAND3_X1  g555(.A1(new_n755), .A2(G43gat), .A3(new_n756), .ZN(new_n757));
  INV_X1    g556(.A(new_n732), .ZN(new_n758));
  NAND3_X1  g557(.A1(new_n758), .A2(new_n527), .A3(new_n502), .ZN(new_n759));
  NAND3_X1  g558(.A1(new_n757), .A2(KEYINPUT47), .A3(new_n759), .ZN(new_n760));
  NAND2_X1  g559(.A1(new_n753), .A2(G43gat), .ZN(new_n761));
  AND2_X1   g560(.A1(new_n759), .A2(new_n761), .ZN(new_n762));
  OAI21_X1  g561(.A(new_n760), .B1(KEYINPUT47), .B2(new_n762), .ZN(G1330gat));
  NAND3_X1  g562(.A1(new_n758), .A2(new_n525), .A3(new_n486), .ZN(new_n764));
  AND3_X1   g563(.A1(new_n726), .A2(new_n486), .A3(new_n728), .ZN(new_n765));
  OAI21_X1  g564(.A(new_n764), .B1(new_n765), .B2(new_n525), .ZN(new_n766));
  AOI21_X1  g565(.A(KEYINPUT48), .B1(new_n764), .B2(KEYINPUT107), .ZN(new_n767));
  XNOR2_X1  g566(.A(new_n766), .B(new_n767), .ZN(G1331gat));
  NOR3_X1   g567(.A1(new_n669), .A2(new_n582), .A3(new_n690), .ZN(new_n769));
  NAND3_X1  g568(.A1(new_n514), .A2(new_n644), .A3(new_n769), .ZN(new_n770));
  NOR2_X1   g569(.A1(new_n770), .A2(new_n694), .ZN(new_n771));
  XOR2_X1   g570(.A(KEYINPUT108), .B(G57gat), .Z(new_n772));
  XNOR2_X1  g571(.A(new_n771), .B(new_n772), .ZN(G1332gat));
  AOI21_X1  g572(.A(new_n487), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n774));
  XNOR2_X1  g573(.A(new_n774), .B(KEYINPUT109), .ZN(new_n775));
  NOR2_X1   g574(.A1(new_n770), .A2(new_n775), .ZN(new_n776));
  NOR2_X1   g575(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n777));
  XNOR2_X1  g576(.A(new_n776), .B(new_n777), .ZN(G1333gat));
  INV_X1    g577(.A(G71gat), .ZN(new_n779));
  OAI21_X1  g578(.A(new_n779), .B1(new_n770), .B2(new_n300), .ZN(new_n780));
  NOR2_X1   g579(.A1(new_n770), .A2(new_n779), .ZN(new_n781));
  AND3_X1   g580(.A1(new_n781), .A2(KEYINPUT110), .A3(new_n752), .ZN(new_n782));
  AOI21_X1  g581(.A(KEYINPUT110), .B1(new_n781), .B2(new_n752), .ZN(new_n783));
  OAI21_X1  g582(.A(new_n780), .B1(new_n782), .B2(new_n783), .ZN(new_n784));
  NAND2_X1  g583(.A1(new_n784), .A2(KEYINPUT50), .ZN(new_n785));
  INV_X1    g584(.A(KEYINPUT50), .ZN(new_n786));
  OAI211_X1 g585(.A(new_n786), .B(new_n780), .C1(new_n782), .C2(new_n783), .ZN(new_n787));
  NAND2_X1  g586(.A1(new_n785), .A2(new_n787), .ZN(G1334gat));
  NOR2_X1   g587(.A1(new_n770), .A2(new_n373), .ZN(new_n789));
  XOR2_X1   g588(.A(new_n789), .B(G78gat), .Z(G1335gat));
  NAND2_X1  g589(.A1(new_n667), .A2(new_n668), .ZN(new_n791));
  INV_X1    g590(.A(new_n644), .ZN(new_n792));
  NOR3_X1   g591(.A1(new_n791), .A2(new_n582), .A3(new_n792), .ZN(new_n793));
  NAND3_X1  g592(.A1(new_n724), .A2(new_n725), .A3(new_n793), .ZN(new_n794));
  INV_X1    g593(.A(KEYINPUT111), .ZN(new_n795));
  NAND2_X1  g594(.A1(new_n794), .A2(new_n795), .ZN(new_n796));
  NAND4_X1  g595(.A1(new_n724), .A2(KEYINPUT111), .A3(new_n725), .A4(new_n793), .ZN(new_n797));
  NAND2_X1  g596(.A1(new_n796), .A2(new_n797), .ZN(new_n798));
  NAND2_X1  g597(.A1(new_n798), .A2(new_n695), .ZN(new_n799));
  INV_X1    g598(.A(KEYINPUT112), .ZN(new_n800));
  NAND2_X1  g599(.A1(new_n799), .A2(new_n800), .ZN(new_n801));
  NAND3_X1  g600(.A1(new_n798), .A2(KEYINPUT112), .A3(new_n695), .ZN(new_n802));
  NAND3_X1  g601(.A1(new_n801), .A2(G85gat), .A3(new_n802), .ZN(new_n803));
  NOR2_X1   g602(.A1(new_n791), .A2(new_n582), .ZN(new_n804));
  OAI211_X1 g603(.A(new_n690), .B(new_n804), .C1(new_n501), .C2(new_n513), .ZN(new_n805));
  AND2_X1   g604(.A1(new_n805), .A2(KEYINPUT51), .ZN(new_n806));
  NOR2_X1   g605(.A1(new_n805), .A2(KEYINPUT51), .ZN(new_n807));
  NOR2_X1   g606(.A1(new_n806), .A2(new_n807), .ZN(new_n808));
  NAND4_X1  g607(.A1(new_n808), .A2(new_n608), .A3(new_n695), .A4(new_n644), .ZN(new_n809));
  NAND2_X1  g608(.A1(new_n803), .A2(new_n809), .ZN(G1336gat));
  AOI21_X1  g609(.A(new_n609), .B1(new_n798), .B2(new_n488), .ZN(new_n811));
  NAND3_X1  g610(.A1(new_n808), .A2(new_n644), .A3(new_n488), .ZN(new_n812));
  NOR2_X1   g611(.A1(new_n812), .A2(G92gat), .ZN(new_n813));
  OAI21_X1  g612(.A(KEYINPUT52), .B1(new_n811), .B2(new_n813), .ZN(new_n814));
  OAI21_X1  g613(.A(G92gat), .B1(new_n794), .B2(new_n487), .ZN(new_n815));
  INV_X1    g614(.A(KEYINPUT52), .ZN(new_n816));
  OAI211_X1 g615(.A(new_n815), .B(new_n816), .C1(new_n812), .C2(G92gat), .ZN(new_n817));
  NAND2_X1  g616(.A1(new_n814), .A2(new_n817), .ZN(G1337gat));
  INV_X1    g617(.A(G99gat), .ZN(new_n819));
  NAND4_X1  g618(.A1(new_n808), .A2(new_n819), .A3(new_n644), .A4(new_n502), .ZN(new_n820));
  AOI21_X1  g619(.A(new_n304), .B1(new_n796), .B2(new_n797), .ZN(new_n821));
  OAI21_X1  g620(.A(new_n820), .B1(new_n821), .B2(new_n819), .ZN(new_n822));
  INV_X1    g621(.A(KEYINPUT113), .ZN(new_n823));
  NAND2_X1  g622(.A1(new_n822), .A2(new_n823), .ZN(new_n824));
  OAI211_X1 g623(.A(KEYINPUT113), .B(new_n820), .C1(new_n821), .C2(new_n819), .ZN(new_n825));
  NAND2_X1  g624(.A1(new_n824), .A2(new_n825), .ZN(G1338gat));
  XOR2_X1   g625(.A(KEYINPUT114), .B(G106gat), .Z(new_n827));
  INV_X1    g626(.A(new_n827), .ZN(new_n828));
  AOI21_X1  g627(.A(new_n828), .B1(new_n798), .B2(new_n486), .ZN(new_n829));
  NAND3_X1  g628(.A1(new_n808), .A2(new_n644), .A3(new_n486), .ZN(new_n830));
  NOR2_X1   g629(.A1(new_n830), .A2(G106gat), .ZN(new_n831));
  OAI21_X1  g630(.A(KEYINPUT53), .B1(new_n829), .B2(new_n831), .ZN(new_n832));
  OAI21_X1  g631(.A(new_n827), .B1(new_n794), .B2(new_n373), .ZN(new_n833));
  INV_X1    g632(.A(KEYINPUT53), .ZN(new_n834));
  OAI211_X1 g633(.A(new_n833), .B(new_n834), .C1(new_n830), .C2(G106gat), .ZN(new_n835));
  NAND2_X1  g634(.A1(new_n832), .A2(new_n835), .ZN(G1339gat));
  NAND3_X1  g635(.A1(new_n628), .A2(new_n632), .A3(new_n629), .ZN(new_n837));
  NAND2_X1  g636(.A1(new_n837), .A2(KEYINPUT115), .ZN(new_n838));
  INV_X1    g637(.A(KEYINPUT115), .ZN(new_n839));
  NAND4_X1  g638(.A1(new_n628), .A2(new_n839), .A3(new_n632), .A4(new_n629), .ZN(new_n840));
  NAND4_X1  g639(.A1(new_n838), .A2(new_n634), .A3(KEYINPUT54), .A4(new_n840), .ZN(new_n841));
  AOI21_X1  g640(.A(new_n632), .B1(new_n628), .B2(new_n629), .ZN(new_n842));
  INV_X1    g641(.A(KEYINPUT54), .ZN(new_n843));
  AOI21_X1  g642(.A(new_n642), .B1(new_n842), .B2(new_n843), .ZN(new_n844));
  AOI21_X1  g643(.A(KEYINPUT55), .B1(new_n841), .B2(new_n844), .ZN(new_n845));
  INV_X1    g644(.A(new_n845), .ZN(new_n846));
  NAND3_X1  g645(.A1(new_n841), .A2(KEYINPUT55), .A3(new_n844), .ZN(new_n847));
  NAND3_X1  g646(.A1(new_n847), .A2(KEYINPUT116), .A3(new_n643), .ZN(new_n848));
  INV_X1    g647(.A(new_n848), .ZN(new_n849));
  AOI21_X1  g648(.A(KEYINPUT116), .B1(new_n847), .B2(new_n643), .ZN(new_n850));
  OAI211_X1 g649(.A(new_n582), .B(new_n846), .C1(new_n849), .C2(new_n850), .ZN(new_n851));
  NAND2_X1  g650(.A1(new_n554), .A2(new_n555), .ZN(new_n852));
  INV_X1    g651(.A(new_n556), .ZN(new_n853));
  AOI21_X1  g652(.A(KEYINPUT117), .B1(new_n852), .B2(new_n853), .ZN(new_n854));
  INV_X1    g653(.A(KEYINPUT117), .ZN(new_n855));
  AOI211_X1 g654(.A(new_n855), .B(new_n556), .C1(new_n554), .C2(new_n555), .ZN(new_n856));
  NOR2_X1   g655(.A1(new_n564), .A2(new_n567), .ZN(new_n857));
  NOR3_X1   g656(.A1(new_n854), .A2(new_n856), .A3(new_n857), .ZN(new_n858));
  OAI21_X1  g657(.A(KEYINPUT118), .B1(new_n858), .B2(new_n577), .ZN(new_n859));
  NAND2_X1  g658(.A1(new_n852), .A2(new_n853), .ZN(new_n860));
  NAND2_X1  g659(.A1(new_n860), .A2(new_n855), .ZN(new_n861));
  INV_X1    g660(.A(new_n857), .ZN(new_n862));
  NAND3_X1  g661(.A1(new_n852), .A2(KEYINPUT117), .A3(new_n853), .ZN(new_n863));
  NAND3_X1  g662(.A1(new_n861), .A2(new_n862), .A3(new_n863), .ZN(new_n864));
  INV_X1    g663(.A(KEYINPUT118), .ZN(new_n865));
  INV_X1    g664(.A(new_n577), .ZN(new_n866));
  NAND3_X1  g665(.A1(new_n864), .A2(new_n865), .A3(new_n866), .ZN(new_n867));
  NAND4_X1  g666(.A1(new_n859), .A2(new_n581), .A3(new_n644), .A4(new_n867), .ZN(new_n868));
  AOI21_X1  g667(.A(new_n690), .B1(new_n851), .B2(new_n868), .ZN(new_n869));
  NOR2_X1   g668(.A1(new_n849), .A2(new_n850), .ZN(new_n870));
  NAND4_X1  g669(.A1(new_n690), .A2(new_n859), .A3(new_n581), .A4(new_n867), .ZN(new_n871));
  NOR3_X1   g670(.A1(new_n870), .A2(new_n871), .A3(new_n845), .ZN(new_n872));
  OAI21_X1  g671(.A(new_n669), .B1(new_n869), .B2(new_n872), .ZN(new_n873));
  INV_X1    g672(.A(new_n690), .ZN(new_n874));
  NAND4_X1  g673(.A1(new_n791), .A2(new_n583), .A3(new_n792), .A4(new_n874), .ZN(new_n875));
  NAND2_X1  g674(.A1(new_n873), .A2(new_n875), .ZN(new_n876));
  AND2_X1   g675(.A1(new_n876), .A2(new_n510), .ZN(new_n877));
  NOR2_X1   g676(.A1(new_n488), .A2(new_n694), .ZN(new_n878));
  NAND2_X1  g677(.A1(new_n877), .A2(new_n878), .ZN(new_n879));
  NOR2_X1   g678(.A1(new_n879), .A2(new_n583), .ZN(new_n880));
  XNOR2_X1  g679(.A(new_n880), .B(new_n248), .ZN(G1340gat));
  NOR2_X1   g680(.A1(new_n879), .A2(new_n792), .ZN(new_n882));
  XNOR2_X1  g681(.A(new_n882), .B(new_n251), .ZN(G1341gat));
  NOR2_X1   g682(.A1(new_n879), .A2(new_n669), .ZN(new_n884));
  NAND2_X1  g683(.A1(new_n240), .A2(new_n242), .ZN(new_n885));
  XOR2_X1   g684(.A(new_n885), .B(KEYINPUT119), .Z(new_n886));
  XNOR2_X1  g685(.A(new_n884), .B(new_n886), .ZN(G1342gat));
  NOR2_X1   g686(.A1(new_n879), .A2(new_n874), .ZN(new_n888));
  NOR2_X1   g687(.A1(KEYINPUT56), .A2(G134gat), .ZN(new_n889));
  AND2_X1   g688(.A1(KEYINPUT56), .A2(G134gat), .ZN(new_n890));
  OAI21_X1  g689(.A(new_n888), .B1(new_n889), .B2(new_n890), .ZN(new_n891));
  OAI21_X1  g690(.A(new_n891), .B1(new_n888), .B2(new_n889), .ZN(G1343gat));
  NAND2_X1  g691(.A1(new_n876), .A2(new_n486), .ZN(new_n893));
  INV_X1    g692(.A(KEYINPUT120), .ZN(new_n894));
  INV_X1    g693(.A(KEYINPUT57), .ZN(new_n895));
  NAND3_X1  g694(.A1(new_n893), .A2(new_n894), .A3(new_n895), .ZN(new_n896));
  INV_X1    g695(.A(new_n875), .ZN(new_n897));
  AND3_X1   g696(.A1(new_n859), .A2(new_n581), .A3(new_n867), .ZN(new_n898));
  NAND2_X1  g697(.A1(new_n847), .A2(new_n643), .ZN(new_n899));
  INV_X1    g698(.A(KEYINPUT116), .ZN(new_n900));
  NAND2_X1  g699(.A1(new_n899), .A2(new_n900), .ZN(new_n901));
  NAND2_X1  g700(.A1(new_n901), .A2(new_n848), .ZN(new_n902));
  NAND4_X1  g701(.A1(new_n898), .A2(new_n902), .A3(new_n690), .A4(new_n846), .ZN(new_n903));
  AND2_X1   g702(.A1(new_n847), .A2(new_n643), .ZN(new_n904));
  NAND3_X1  g703(.A1(new_n582), .A2(new_n904), .A3(new_n846), .ZN(new_n905));
  NAND2_X1  g704(.A1(new_n905), .A2(new_n868), .ZN(new_n906));
  NAND2_X1  g705(.A1(new_n906), .A2(new_n874), .ZN(new_n907));
  AOI21_X1  g706(.A(new_n791), .B1(new_n903), .B2(new_n907), .ZN(new_n908));
  OAI211_X1 g707(.A(KEYINPUT57), .B(new_n486), .C1(new_n897), .C2(new_n908), .ZN(new_n909));
  AOI21_X1  g708(.A(new_n373), .B1(new_n873), .B2(new_n875), .ZN(new_n910));
  OAI21_X1  g709(.A(KEYINPUT120), .B1(new_n910), .B2(KEYINPUT57), .ZN(new_n911));
  NAND3_X1  g710(.A1(new_n896), .A2(new_n909), .A3(new_n911), .ZN(new_n912));
  NAND2_X1  g711(.A1(new_n878), .A2(new_n304), .ZN(new_n913));
  INV_X1    g712(.A(new_n913), .ZN(new_n914));
  NAND2_X1  g713(.A1(new_n912), .A2(new_n914), .ZN(new_n915));
  OAI21_X1  g714(.A(G141gat), .B1(new_n915), .B2(new_n583), .ZN(new_n916));
  NOR2_X1   g715(.A1(new_n893), .A2(new_n913), .ZN(new_n917));
  NAND2_X1  g716(.A1(new_n582), .A2(new_n321), .ZN(new_n918));
  XNOR2_X1  g717(.A(new_n918), .B(KEYINPUT121), .ZN(new_n919));
  NAND2_X1  g718(.A1(new_n917), .A2(new_n919), .ZN(new_n920));
  NAND2_X1  g719(.A1(new_n916), .A2(new_n920), .ZN(new_n921));
  NAND2_X1  g720(.A1(new_n921), .A2(KEYINPUT58), .ZN(new_n922));
  INV_X1    g721(.A(KEYINPUT58), .ZN(new_n923));
  NAND3_X1  g722(.A1(new_n916), .A2(new_n923), .A3(new_n920), .ZN(new_n924));
  NAND2_X1  g723(.A1(new_n922), .A2(new_n924), .ZN(G1344gat));
  NAND3_X1  g724(.A1(new_n917), .A2(new_n319), .A3(new_n644), .ZN(new_n926));
  INV_X1    g725(.A(new_n915), .ZN(new_n927));
  AOI211_X1 g726(.A(KEYINPUT59), .B(new_n319), .C1(new_n927), .C2(new_n644), .ZN(new_n928));
  INV_X1    g727(.A(KEYINPUT59), .ZN(new_n929));
  INV_X1    g728(.A(KEYINPUT122), .ZN(new_n930));
  AOI21_X1  g729(.A(new_n690), .B1(new_n905), .B2(new_n868), .ZN(new_n931));
  OAI21_X1  g730(.A(new_n930), .B1(new_n872), .B2(new_n931), .ZN(new_n932));
  NAND3_X1  g731(.A1(new_n907), .A2(KEYINPUT122), .A3(new_n903), .ZN(new_n933));
  NAND3_X1  g732(.A1(new_n932), .A2(new_n933), .A3(new_n669), .ZN(new_n934));
  NAND2_X1  g733(.A1(new_n934), .A2(new_n875), .ZN(new_n935));
  NAND2_X1  g734(.A1(new_n935), .A2(new_n486), .ZN(new_n936));
  INV_X1    g735(.A(KEYINPUT123), .ZN(new_n937));
  NAND3_X1  g736(.A1(new_n936), .A2(new_n937), .A3(new_n895), .ZN(new_n938));
  NAND2_X1  g737(.A1(new_n910), .A2(KEYINPUT57), .ZN(new_n939));
  AOI21_X1  g738(.A(new_n373), .B1(new_n934), .B2(new_n875), .ZN(new_n940));
  OAI21_X1  g739(.A(KEYINPUT123), .B1(new_n940), .B2(KEYINPUT57), .ZN(new_n941));
  NAND3_X1  g740(.A1(new_n938), .A2(new_n939), .A3(new_n941), .ZN(new_n942));
  NAND3_X1  g741(.A1(new_n942), .A2(new_n644), .A3(new_n914), .ZN(new_n943));
  AOI21_X1  g742(.A(new_n929), .B1(new_n943), .B2(G148gat), .ZN(new_n944));
  OAI21_X1  g743(.A(new_n926), .B1(new_n928), .B2(new_n944), .ZN(G1345gat));
  AOI21_X1  g744(.A(G155gat), .B1(new_n917), .B2(new_n791), .ZN(new_n946));
  AND2_X1   g745(.A1(new_n791), .A2(G155gat), .ZN(new_n947));
  AOI21_X1  g746(.A(new_n946), .B1(new_n927), .B2(new_n947), .ZN(G1346gat));
  AOI21_X1  g747(.A(G162gat), .B1(new_n917), .B2(new_n690), .ZN(new_n949));
  AND2_X1   g748(.A1(new_n690), .A2(G162gat), .ZN(new_n950));
  AOI21_X1  g749(.A(new_n949), .B1(new_n927), .B2(new_n950), .ZN(G1347gat));
  NOR2_X1   g750(.A1(new_n695), .A2(new_n487), .ZN(new_n952));
  AND2_X1   g751(.A1(new_n877), .A2(new_n952), .ZN(new_n953));
  NAND3_X1  g752(.A1(new_n953), .A2(new_n226), .A3(new_n582), .ZN(new_n954));
  XOR2_X1   g753(.A(new_n952), .B(KEYINPUT124), .Z(new_n955));
  NAND2_X1  g754(.A1(new_n877), .A2(new_n955), .ZN(new_n956));
  NAND2_X1  g755(.A1(new_n956), .A2(KEYINPUT125), .ZN(new_n957));
  INV_X1    g756(.A(KEYINPUT125), .ZN(new_n958));
  NAND3_X1  g757(.A1(new_n877), .A2(new_n958), .A3(new_n955), .ZN(new_n959));
  AND2_X1   g758(.A1(new_n957), .A2(new_n959), .ZN(new_n960));
  AND2_X1   g759(.A1(new_n960), .A2(new_n582), .ZN(new_n961));
  OAI21_X1  g760(.A(new_n954), .B1(new_n961), .B2(new_n226), .ZN(G1348gat));
  AOI21_X1  g761(.A(G176gat), .B1(new_n953), .B2(new_n644), .ZN(new_n963));
  NOR2_X1   g762(.A1(new_n792), .A2(new_n227), .ZN(new_n964));
  AOI21_X1  g763(.A(new_n963), .B1(new_n960), .B2(new_n964), .ZN(G1349gat));
  NAND3_X1  g764(.A1(new_n957), .A2(new_n791), .A3(new_n959), .ZN(new_n966));
  NAND2_X1  g765(.A1(new_n966), .A2(G183gat), .ZN(new_n967));
  OAI211_X1 g766(.A(new_n953), .B(new_n791), .C1(new_n206), .C2(new_n205), .ZN(new_n968));
  NAND2_X1  g767(.A1(new_n967), .A2(new_n968), .ZN(new_n969));
  NAND2_X1  g768(.A1(new_n969), .A2(KEYINPUT60), .ZN(new_n970));
  INV_X1    g769(.A(KEYINPUT60), .ZN(new_n971));
  NAND3_X1  g770(.A1(new_n967), .A2(new_n968), .A3(new_n971), .ZN(new_n972));
  NAND2_X1  g771(.A1(new_n970), .A2(new_n972), .ZN(G1350gat));
  NAND3_X1  g772(.A1(new_n953), .A2(new_n204), .A3(new_n690), .ZN(new_n974));
  NAND3_X1  g773(.A1(new_n957), .A2(new_n690), .A3(new_n959), .ZN(new_n975));
  INV_X1    g774(.A(KEYINPUT61), .ZN(new_n976));
  AND3_X1   g775(.A1(new_n975), .A2(new_n976), .A3(G190gat), .ZN(new_n977));
  AOI21_X1  g776(.A(new_n976), .B1(new_n975), .B2(G190gat), .ZN(new_n978));
  OAI21_X1  g777(.A(new_n974), .B1(new_n977), .B2(new_n978), .ZN(G1351gat));
  INV_X1    g778(.A(KEYINPUT126), .ZN(new_n980));
  AND2_X1   g779(.A1(new_n955), .A2(new_n304), .ZN(new_n981));
  NAND3_X1  g780(.A1(new_n942), .A2(new_n582), .A3(new_n981), .ZN(new_n982));
  NAND2_X1  g781(.A1(new_n982), .A2(G197gat), .ZN(new_n983));
  INV_X1    g782(.A(new_n952), .ZN(new_n984));
  NOR3_X1   g783(.A1(new_n893), .A2(new_n752), .A3(new_n984), .ZN(new_n985));
  INV_X1    g784(.A(G197gat), .ZN(new_n986));
  NAND3_X1  g785(.A1(new_n985), .A2(new_n986), .A3(new_n582), .ZN(new_n987));
  AOI21_X1  g786(.A(new_n980), .B1(new_n983), .B2(new_n987), .ZN(new_n988));
  INV_X1    g787(.A(new_n987), .ZN(new_n989));
  AOI211_X1 g788(.A(KEYINPUT126), .B(new_n989), .C1(new_n982), .C2(G197gat), .ZN(new_n990));
  NOR2_X1   g789(.A1(new_n988), .A2(new_n990), .ZN(G1352gat));
  INV_X1    g790(.A(new_n985), .ZN(new_n992));
  NOR3_X1   g791(.A1(new_n992), .A2(G204gat), .A3(new_n792), .ZN(new_n993));
  XNOR2_X1  g792(.A(new_n993), .B(KEYINPUT62), .ZN(new_n994));
  NAND3_X1  g793(.A1(new_n942), .A2(new_n644), .A3(new_n981), .ZN(new_n995));
  NAND2_X1  g794(.A1(new_n995), .A2(G204gat), .ZN(new_n996));
  NAND2_X1  g795(.A1(new_n994), .A2(new_n996), .ZN(G1353gat));
  NAND3_X1  g796(.A1(new_n942), .A2(new_n791), .A3(new_n981), .ZN(new_n998));
  NAND2_X1  g797(.A1(new_n998), .A2(G211gat), .ZN(new_n999));
  NAND2_X1  g798(.A1(new_n999), .A2(KEYINPUT63), .ZN(new_n1000));
  INV_X1    g799(.A(KEYINPUT63), .ZN(new_n1001));
  NAND3_X1  g800(.A1(new_n998), .A2(new_n1001), .A3(G211gat), .ZN(new_n1002));
  NAND3_X1  g801(.A1(new_n985), .A2(new_n331), .A3(new_n791), .ZN(new_n1003));
  XNOR2_X1  g802(.A(new_n1003), .B(KEYINPUT127), .ZN(new_n1004));
  NAND3_X1  g803(.A1(new_n1000), .A2(new_n1002), .A3(new_n1004), .ZN(G1354gat));
  NAND3_X1  g804(.A1(new_n985), .A2(new_n332), .A3(new_n690), .ZN(new_n1006));
  AND3_X1   g805(.A1(new_n942), .A2(new_n690), .A3(new_n981), .ZN(new_n1007));
  OAI21_X1  g806(.A(new_n1006), .B1(new_n1007), .B2(new_n332), .ZN(G1355gat));
endmodule


