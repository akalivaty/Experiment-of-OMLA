//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 1 1 0 1 0 0 1 1 0 0 0 1 0 1 1 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 0 0 0 0 0 0 1 0 0 1 0 0 1 1 0 0 1 1 1 1 0 1 0 0 0 1 1 0 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:16:19 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n650, new_n651, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n681, new_n682,
    new_n683, new_n684, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n725, new_n726, new_n727, new_n728,
    new_n730, new_n731, new_n732, new_n733, new_n735, new_n736, new_n738,
    new_n739, new_n740, new_n741, new_n742, new_n743, new_n744, new_n745,
    new_n746, new_n747, new_n748, new_n749, new_n750, new_n751, new_n752,
    new_n753, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n771, new_n772, new_n773, new_n774, new_n775,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n820,
    new_n821, new_n822, new_n824, new_n825, new_n826, new_n828, new_n829,
    new_n830, new_n831, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n863, new_n864, new_n866, new_n867, new_n868,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n878, new_n879, new_n880, new_n882, new_n883, new_n884, new_n885,
    new_n886, new_n887, new_n888, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n915, new_n916, new_n917,
    new_n918, new_n919, new_n920, new_n922, new_n923;
  NAND2_X1  g000(.A1(G29gat), .A2(G36gat), .ZN(new_n202));
  XOR2_X1   g001(.A(new_n202), .B(KEYINPUT93), .Z(new_n203));
  OAI21_X1  g002(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n204));
  INV_X1    g003(.A(new_n204), .ZN(new_n205));
  NOR3_X1   g004(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n206));
  OAI21_X1  g005(.A(new_n203), .B1(new_n205), .B2(new_n206), .ZN(new_n207));
  XNOR2_X1  g006(.A(G43gat), .B(G50gat), .ZN(new_n208));
  INV_X1    g007(.A(KEYINPUT92), .ZN(new_n209));
  XNOR2_X1  g008(.A(new_n208), .B(new_n209), .ZN(new_n210));
  NAND3_X1  g009(.A1(new_n207), .A2(KEYINPUT15), .A3(new_n210), .ZN(new_n211));
  NAND2_X1  g010(.A1(new_n210), .A2(KEYINPUT15), .ZN(new_n212));
  OAI211_X1 g011(.A(new_n212), .B(new_n203), .C1(KEYINPUT15), .C2(new_n208), .ZN(new_n213));
  XNOR2_X1  g012(.A(new_n206), .B(KEYINPUT95), .ZN(new_n214));
  NAND2_X1  g013(.A1(new_n204), .A2(KEYINPUT94), .ZN(new_n215));
  XNOR2_X1  g014(.A(new_n214), .B(new_n215), .ZN(new_n216));
  OAI21_X1  g015(.A(new_n211), .B1(new_n213), .B2(new_n216), .ZN(new_n217));
  XNOR2_X1  g016(.A(new_n217), .B(KEYINPUT17), .ZN(new_n218));
  XNOR2_X1  g017(.A(G15gat), .B(G22gat), .ZN(new_n219));
  INV_X1    g018(.A(G1gat), .ZN(new_n220));
  NAND3_X1  g019(.A1(new_n219), .A2(KEYINPUT16), .A3(new_n220), .ZN(new_n221));
  OAI21_X1  g020(.A(new_n221), .B1(new_n220), .B2(new_n219), .ZN(new_n222));
  INV_X1    g021(.A(G8gat), .ZN(new_n223));
  AOI21_X1  g022(.A(new_n222), .B1(KEYINPUT96), .B2(new_n223), .ZN(new_n224));
  NOR2_X1   g023(.A1(new_n223), .A2(KEYINPUT96), .ZN(new_n225));
  XNOR2_X1  g024(.A(new_n224), .B(new_n225), .ZN(new_n226));
  INV_X1    g025(.A(new_n226), .ZN(new_n227));
  MUX2_X1   g026(.A(new_n217), .B(new_n218), .S(new_n227), .Z(new_n228));
  NAND2_X1  g027(.A1(G229gat), .A2(G233gat), .ZN(new_n229));
  XNOR2_X1  g028(.A(new_n229), .B(KEYINPUT97), .ZN(new_n230));
  NOR2_X1   g029(.A1(new_n228), .A2(new_n230), .ZN(new_n231));
  XOR2_X1   g030(.A(new_n231), .B(KEYINPUT18), .Z(new_n232));
  XOR2_X1   g031(.A(new_n226), .B(new_n217), .Z(new_n233));
  XOR2_X1   g032(.A(new_n230), .B(KEYINPUT13), .Z(new_n234));
  OAI21_X1  g033(.A(new_n232), .B1(new_n233), .B2(new_n234), .ZN(new_n235));
  XNOR2_X1  g034(.A(G113gat), .B(G141gat), .ZN(new_n236));
  XNOR2_X1  g035(.A(new_n236), .B(G197gat), .ZN(new_n237));
  XNOR2_X1  g036(.A(new_n237), .B(KEYINPUT11), .ZN(new_n238));
  INV_X1    g037(.A(G169gat), .ZN(new_n239));
  XNOR2_X1  g038(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XOR2_X1   g039(.A(new_n240), .B(KEYINPUT12), .Z(new_n241));
  NOR2_X1   g040(.A1(new_n235), .A2(new_n241), .ZN(new_n242));
  XNOR2_X1  g041(.A(new_n242), .B(KEYINPUT98), .ZN(new_n243));
  XNOR2_X1  g042(.A(new_n241), .B(KEYINPUT91), .ZN(new_n244));
  NAND2_X1  g043(.A1(new_n235), .A2(new_n244), .ZN(new_n245));
  NAND2_X1  g044(.A1(new_n243), .A2(new_n245), .ZN(new_n246));
  INV_X1    g045(.A(new_n246), .ZN(new_n247));
  INV_X1    g046(.A(KEYINPUT78), .ZN(new_n248));
  NAND2_X1  g047(.A1(G183gat), .A2(G190gat), .ZN(new_n249));
  NAND2_X1  g048(.A1(G169gat), .A2(G176gat), .ZN(new_n250));
  NAND2_X1  g049(.A1(new_n250), .A2(KEYINPUT65), .ZN(new_n251));
  INV_X1    g050(.A(KEYINPUT65), .ZN(new_n252));
  NAND3_X1  g051(.A1(new_n252), .A2(G169gat), .A3(G176gat), .ZN(new_n253));
  NAND2_X1  g052(.A1(new_n251), .A2(new_n253), .ZN(new_n254));
  INV_X1    g053(.A(KEYINPUT26), .ZN(new_n255));
  NOR2_X1   g054(.A1(G169gat), .A2(G176gat), .ZN(new_n256));
  NOR4_X1   g055(.A1(KEYINPUT73), .A2(KEYINPUT26), .A3(G169gat), .A4(G176gat), .ZN(new_n257));
  INV_X1    g056(.A(KEYINPUT73), .ZN(new_n258));
  AOI21_X1  g057(.A(new_n258), .B1(new_n256), .B2(new_n255), .ZN(new_n259));
  OAI221_X1 g058(.A(new_n254), .B1(new_n255), .B2(new_n256), .C1(new_n257), .C2(new_n259), .ZN(new_n260));
  INV_X1    g059(.A(KEYINPUT28), .ZN(new_n261));
  INV_X1    g060(.A(G190gat), .ZN(new_n262));
  INV_X1    g061(.A(KEYINPUT27), .ZN(new_n263));
  NAND2_X1  g062(.A1(new_n263), .A2(G183gat), .ZN(new_n264));
  OAI21_X1  g063(.A(new_n262), .B1(new_n264), .B2(KEYINPUT70), .ZN(new_n265));
  INV_X1    g064(.A(KEYINPUT70), .ZN(new_n266));
  AOI21_X1  g065(.A(new_n263), .B1(new_n266), .B2(G183gat), .ZN(new_n267));
  OAI21_X1  g066(.A(new_n261), .B1(new_n265), .B2(new_n267), .ZN(new_n268));
  XNOR2_X1  g067(.A(new_n268), .B(KEYINPUT71), .ZN(new_n269));
  XNOR2_X1  g068(.A(KEYINPUT27), .B(G183gat), .ZN(new_n270));
  NAND3_X1  g069(.A1(new_n270), .A2(KEYINPUT28), .A3(new_n262), .ZN(new_n271));
  XOR2_X1   g070(.A(new_n271), .B(KEYINPUT72), .Z(new_n272));
  OAI211_X1 g071(.A(new_n249), .B(new_n260), .C1(new_n269), .C2(new_n272), .ZN(new_n273));
  OAI21_X1  g072(.A(KEYINPUT64), .B1(new_n256), .B2(KEYINPUT23), .ZN(new_n274));
  INV_X1    g073(.A(KEYINPUT64), .ZN(new_n275));
  INV_X1    g074(.A(KEYINPUT23), .ZN(new_n276));
  OAI211_X1 g075(.A(new_n275), .B(new_n276), .C1(G169gat), .C2(G176gat), .ZN(new_n277));
  NAND2_X1  g076(.A1(new_n274), .A2(new_n277), .ZN(new_n278));
  AOI22_X1  g077(.A1(new_n251), .A2(new_n253), .B1(KEYINPUT23), .B2(new_n256), .ZN(new_n279));
  NAND2_X1  g078(.A1(new_n278), .A2(new_n279), .ZN(new_n280));
  NAND2_X1  g079(.A1(new_n280), .A2(KEYINPUT66), .ZN(new_n281));
  NOR2_X1   g080(.A1(new_n249), .A2(KEYINPUT24), .ZN(new_n282));
  INV_X1    g081(.A(KEYINPUT24), .ZN(new_n283));
  AOI21_X1  g082(.A(new_n283), .B1(G183gat), .B2(G190gat), .ZN(new_n284));
  NOR2_X1   g083(.A1(G183gat), .A2(G190gat), .ZN(new_n285));
  INV_X1    g084(.A(new_n285), .ZN(new_n286));
  AOI21_X1  g085(.A(new_n282), .B1(new_n284), .B2(new_n286), .ZN(new_n287));
  INV_X1    g086(.A(KEYINPUT66), .ZN(new_n288));
  NAND3_X1  g087(.A1(new_n278), .A2(new_n279), .A3(new_n288), .ZN(new_n289));
  NAND3_X1  g088(.A1(new_n281), .A2(new_n287), .A3(new_n289), .ZN(new_n290));
  INV_X1    g089(.A(KEYINPUT25), .ZN(new_n291));
  NAND2_X1  g090(.A1(new_n290), .A2(new_n291), .ZN(new_n292));
  INV_X1    g091(.A(KEYINPUT69), .ZN(new_n293));
  INV_X1    g092(.A(KEYINPUT68), .ZN(new_n294));
  INV_X1    g093(.A(KEYINPUT67), .ZN(new_n295));
  NAND2_X1  g094(.A1(new_n254), .A2(new_n295), .ZN(new_n296));
  NAND3_X1  g095(.A1(new_n251), .A2(new_n253), .A3(KEYINPUT67), .ZN(new_n297));
  NAND3_X1  g096(.A1(new_n296), .A2(new_n278), .A3(new_n297), .ZN(new_n298));
  AOI21_X1  g097(.A(new_n291), .B1(new_n256), .B2(KEYINPUT23), .ZN(new_n299));
  NAND2_X1  g098(.A1(new_n287), .A2(new_n299), .ZN(new_n300));
  OAI21_X1  g099(.A(new_n294), .B1(new_n298), .B2(new_n300), .ZN(new_n301));
  AND3_X1   g100(.A1(new_n251), .A2(new_n253), .A3(KEYINPUT67), .ZN(new_n302));
  AOI21_X1  g101(.A(KEYINPUT67), .B1(new_n251), .B2(new_n253), .ZN(new_n303));
  NOR2_X1   g102(.A1(new_n302), .A2(new_n303), .ZN(new_n304));
  INV_X1    g103(.A(new_n299), .ZN(new_n305));
  NAND3_X1  g104(.A1(new_n283), .A2(G183gat), .A3(G190gat), .ZN(new_n306));
  NAND2_X1  g105(.A1(new_n249), .A2(KEYINPUT24), .ZN(new_n307));
  OAI21_X1  g106(.A(new_n306), .B1(new_n307), .B2(new_n285), .ZN(new_n308));
  NOR2_X1   g107(.A1(new_n305), .A2(new_n308), .ZN(new_n309));
  NAND4_X1  g108(.A1(new_n304), .A2(new_n309), .A3(KEYINPUT68), .A4(new_n278), .ZN(new_n310));
  NAND2_X1  g109(.A1(new_n301), .A2(new_n310), .ZN(new_n311));
  AND3_X1   g110(.A1(new_n292), .A2(new_n293), .A3(new_n311), .ZN(new_n312));
  AOI21_X1  g111(.A(new_n293), .B1(new_n292), .B2(new_n311), .ZN(new_n313));
  OAI21_X1  g112(.A(new_n273), .B1(new_n312), .B2(new_n313), .ZN(new_n314));
  INV_X1    g113(.A(KEYINPUT75), .ZN(new_n315));
  NAND2_X1  g114(.A1(new_n314), .A2(new_n315), .ZN(new_n316));
  OAI211_X1 g115(.A(KEYINPUT75), .B(new_n273), .C1(new_n312), .C2(new_n313), .ZN(new_n317));
  NAND2_X1  g116(.A1(new_n316), .A2(new_n317), .ZN(new_n318));
  NAND2_X1  g117(.A1(G226gat), .A2(G233gat), .ZN(new_n319));
  INV_X1    g118(.A(new_n319), .ZN(new_n320));
  AOI21_X1  g119(.A(new_n248), .B1(new_n318), .B2(new_n320), .ZN(new_n321));
  AOI211_X1 g120(.A(KEYINPUT78), .B(new_n319), .C1(new_n316), .C2(new_n317), .ZN(new_n322));
  NOR2_X1   g121(.A1(new_n321), .A2(new_n322), .ZN(new_n323));
  INV_X1    g122(.A(G211gat), .ZN(new_n324));
  INV_X1    g123(.A(G218gat), .ZN(new_n325));
  NOR2_X1   g124(.A1(new_n324), .A2(new_n325), .ZN(new_n326));
  INV_X1    g125(.A(new_n326), .ZN(new_n327));
  NAND2_X1  g126(.A1(new_n324), .A2(new_n325), .ZN(new_n328));
  INV_X1    g127(.A(KEYINPUT22), .ZN(new_n329));
  OAI21_X1  g128(.A(new_n327), .B1(new_n328), .B2(new_n329), .ZN(new_n330));
  XOR2_X1   g129(.A(G197gat), .B(G204gat), .Z(new_n331));
  INV_X1    g130(.A(new_n331), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n330), .A2(new_n332), .ZN(new_n333));
  OAI211_X1 g132(.A(new_n327), .B(new_n328), .C1(new_n331), .C2(new_n329), .ZN(new_n334));
  NAND2_X1  g133(.A1(new_n333), .A2(new_n334), .ZN(new_n335));
  NAND2_X1  g134(.A1(new_n292), .A2(new_n311), .ZN(new_n336));
  NAND2_X1  g135(.A1(new_n273), .A2(new_n336), .ZN(new_n337));
  INV_X1    g136(.A(KEYINPUT29), .ZN(new_n338));
  AOI21_X1  g137(.A(new_n320), .B1(new_n337), .B2(new_n338), .ZN(new_n339));
  INV_X1    g138(.A(KEYINPUT77), .ZN(new_n340));
  XNOR2_X1  g139(.A(new_n339), .B(new_n340), .ZN(new_n341));
  NAND4_X1  g140(.A1(new_n323), .A2(KEYINPUT79), .A3(new_n335), .A4(new_n341), .ZN(new_n342));
  NAND2_X1  g141(.A1(new_n336), .A2(KEYINPUT69), .ZN(new_n343));
  NAND3_X1  g142(.A1(new_n292), .A2(new_n293), .A3(new_n311), .ZN(new_n344));
  NAND2_X1  g143(.A1(new_n343), .A2(new_n344), .ZN(new_n345));
  AOI21_X1  g144(.A(KEYINPUT75), .B1(new_n345), .B2(new_n273), .ZN(new_n346));
  INV_X1    g145(.A(new_n317), .ZN(new_n347));
  OAI21_X1  g146(.A(new_n320), .B1(new_n346), .B2(new_n347), .ZN(new_n348));
  NAND2_X1  g147(.A1(new_n348), .A2(KEYINPUT78), .ZN(new_n349));
  NAND3_X1  g148(.A1(new_n318), .A2(new_n248), .A3(new_n320), .ZN(new_n350));
  NAND4_X1  g149(.A1(new_n349), .A2(new_n335), .A3(new_n350), .A4(new_n341), .ZN(new_n351));
  INV_X1    g150(.A(KEYINPUT79), .ZN(new_n352));
  NAND2_X1  g151(.A1(new_n351), .A2(new_n352), .ZN(new_n353));
  NOR2_X1   g152(.A1(new_n320), .A2(KEYINPUT29), .ZN(new_n354));
  OAI21_X1  g153(.A(new_n354), .B1(new_n346), .B2(new_n347), .ZN(new_n355));
  INV_X1    g154(.A(new_n335), .ZN(new_n356));
  NAND3_X1  g155(.A1(new_n273), .A2(new_n336), .A3(new_n320), .ZN(new_n357));
  NAND3_X1  g156(.A1(new_n355), .A2(new_n356), .A3(new_n357), .ZN(new_n358));
  INV_X1    g157(.A(KEYINPUT76), .ZN(new_n359));
  NAND2_X1  g158(.A1(new_n358), .A2(new_n359), .ZN(new_n360));
  NAND4_X1  g159(.A1(new_n355), .A2(KEYINPUT76), .A3(new_n356), .A4(new_n357), .ZN(new_n361));
  NAND2_X1  g160(.A1(new_n360), .A2(new_n361), .ZN(new_n362));
  NAND3_X1  g161(.A1(new_n342), .A2(new_n353), .A3(new_n362), .ZN(new_n363));
  XNOR2_X1  g162(.A(G8gat), .B(G36gat), .ZN(new_n364));
  INV_X1    g163(.A(G64gat), .ZN(new_n365));
  XNOR2_X1  g164(.A(new_n364), .B(new_n365), .ZN(new_n366));
  INV_X1    g165(.A(G92gat), .ZN(new_n367));
  XNOR2_X1  g166(.A(new_n366), .B(new_n367), .ZN(new_n368));
  XOR2_X1   g167(.A(new_n368), .B(KEYINPUT80), .Z(new_n369));
  INV_X1    g168(.A(new_n369), .ZN(new_n370));
  NAND2_X1  g169(.A1(new_n363), .A2(new_n370), .ZN(new_n371));
  INV_X1    g170(.A(new_n368), .ZN(new_n372));
  NAND4_X1  g171(.A1(new_n342), .A2(new_n353), .A3(new_n362), .A4(new_n372), .ZN(new_n373));
  NAND3_X1  g172(.A1(new_n371), .A2(KEYINPUT30), .A3(new_n373), .ZN(new_n374));
  OR2_X1    g173(.A1(new_n373), .A2(KEYINPUT30), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n374), .A2(new_n375), .ZN(new_n376));
  NAND2_X1  g175(.A1(new_n376), .A2(KEYINPUT89), .ZN(new_n377));
  INV_X1    g176(.A(KEYINPUT89), .ZN(new_n378));
  NAND3_X1  g177(.A1(new_n374), .A2(new_n378), .A3(new_n375), .ZN(new_n379));
  INV_X1    g178(.A(G155gat), .ZN(new_n380));
  INV_X1    g179(.A(G162gat), .ZN(new_n381));
  OAI21_X1  g180(.A(KEYINPUT2), .B1(new_n380), .B2(new_n381), .ZN(new_n382));
  XNOR2_X1  g181(.A(new_n382), .B(KEYINPUT82), .ZN(new_n383));
  INV_X1    g182(.A(G148gat), .ZN(new_n384));
  NAND2_X1  g183(.A1(new_n384), .A2(G141gat), .ZN(new_n385));
  XOR2_X1   g184(.A(KEYINPUT81), .B(G141gat), .Z(new_n386));
  OAI21_X1  g185(.A(new_n385), .B1(new_n386), .B2(new_n384), .ZN(new_n387));
  XNOR2_X1  g186(.A(G155gat), .B(G162gat), .ZN(new_n388));
  NAND3_X1  g187(.A1(new_n383), .A2(new_n387), .A3(new_n388), .ZN(new_n389));
  INV_X1    g188(.A(KEYINPUT83), .ZN(new_n390));
  XNOR2_X1  g189(.A(new_n389), .B(new_n390), .ZN(new_n391));
  INV_X1    g190(.A(new_n388), .ZN(new_n392));
  XNOR2_X1  g191(.A(G141gat), .B(G148gat), .ZN(new_n393));
  OAI21_X1  g192(.A(new_n392), .B1(KEYINPUT2), .B2(new_n393), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n391), .A2(new_n394), .ZN(new_n395));
  INV_X1    g194(.A(G120gat), .ZN(new_n396));
  NAND2_X1  g195(.A1(new_n396), .A2(G113gat), .ZN(new_n397));
  INV_X1    g196(.A(G113gat), .ZN(new_n398));
  NAND2_X1  g197(.A1(new_n398), .A2(G120gat), .ZN(new_n399));
  AOI21_X1  g198(.A(KEYINPUT1), .B1(new_n397), .B2(new_n399), .ZN(new_n400));
  XNOR2_X1  g199(.A(new_n400), .B(G127gat), .ZN(new_n401));
  INV_X1    g200(.A(G134gat), .ZN(new_n402));
  XNOR2_X1  g201(.A(new_n401), .B(new_n402), .ZN(new_n403));
  INV_X1    g202(.A(new_n403), .ZN(new_n404));
  OAI21_X1  g203(.A(KEYINPUT4), .B1(new_n395), .B2(new_n404), .ZN(new_n405));
  OR2_X1    g204(.A1(new_n405), .A2(KEYINPUT87), .ZN(new_n406));
  NOR2_X1   g205(.A1(new_n395), .A2(new_n404), .ZN(new_n407));
  INV_X1    g206(.A(KEYINPUT4), .ZN(new_n408));
  NAND2_X1  g207(.A1(new_n407), .A2(new_n408), .ZN(new_n409));
  NAND2_X1  g208(.A1(new_n409), .A2(KEYINPUT86), .ZN(new_n410));
  NAND2_X1  g209(.A1(new_n405), .A2(KEYINPUT87), .ZN(new_n411));
  INV_X1    g210(.A(KEYINPUT86), .ZN(new_n412));
  NAND3_X1  g211(.A1(new_n407), .A2(new_n412), .A3(new_n408), .ZN(new_n413));
  NAND4_X1  g212(.A1(new_n406), .A2(new_n410), .A3(new_n411), .A4(new_n413), .ZN(new_n414));
  OR2_X1    g213(.A1(new_n395), .A2(KEYINPUT3), .ZN(new_n415));
  XNOR2_X1  g214(.A(new_n403), .B(KEYINPUT84), .ZN(new_n416));
  NAND2_X1  g215(.A1(new_n395), .A2(KEYINPUT3), .ZN(new_n417));
  NAND3_X1  g216(.A1(new_n415), .A2(new_n416), .A3(new_n417), .ZN(new_n418));
  AND2_X1   g217(.A1(new_n414), .A2(new_n418), .ZN(new_n419));
  NAND2_X1  g218(.A1(G225gat), .A2(G233gat), .ZN(new_n420));
  NOR3_X1   g219(.A1(new_n419), .A2(KEYINPUT39), .A3(new_n420), .ZN(new_n421));
  XNOR2_X1  g220(.A(G1gat), .B(G29gat), .ZN(new_n422));
  XNOR2_X1  g221(.A(new_n422), .B(KEYINPUT0), .ZN(new_n423));
  XNOR2_X1  g222(.A(new_n423), .B(G57gat), .ZN(new_n424));
  INV_X1    g223(.A(G85gat), .ZN(new_n425));
  XNOR2_X1  g224(.A(new_n424), .B(new_n425), .ZN(new_n426));
  INV_X1    g225(.A(new_n426), .ZN(new_n427));
  NOR2_X1   g226(.A1(new_n421), .A2(new_n427), .ZN(new_n428));
  AOI21_X1  g227(.A(new_n407), .B1(new_n395), .B2(new_n416), .ZN(new_n429));
  NAND2_X1  g228(.A1(new_n429), .A2(new_n420), .ZN(new_n430));
  OAI211_X1 g229(.A(KEYINPUT39), .B(new_n430), .C1(new_n419), .C2(new_n420), .ZN(new_n431));
  AND3_X1   g230(.A1(new_n428), .A2(KEYINPUT40), .A3(new_n431), .ZN(new_n432));
  AOI21_X1  g231(.A(KEYINPUT40), .B1(new_n428), .B2(new_n431), .ZN(new_n433));
  OR2_X1    g232(.A1(new_n429), .A2(new_n420), .ZN(new_n434));
  NAND3_X1  g233(.A1(new_n409), .A2(KEYINPUT85), .A3(new_n405), .ZN(new_n435));
  NAND2_X1  g234(.A1(new_n435), .A2(new_n420), .ZN(new_n436));
  OR3_X1    g235(.A1(new_n407), .A2(KEYINPUT85), .A3(new_n408), .ZN(new_n437));
  NAND2_X1  g236(.A1(new_n437), .A2(new_n418), .ZN(new_n438));
  OAI211_X1 g237(.A(KEYINPUT5), .B(new_n434), .C1(new_n436), .C2(new_n438), .ZN(new_n439));
  INV_X1    g238(.A(KEYINPUT5), .ZN(new_n440));
  NAND4_X1  g239(.A1(new_n414), .A2(new_n440), .A3(new_n420), .A4(new_n418), .ZN(new_n441));
  AOI21_X1  g240(.A(new_n426), .B1(new_n439), .B2(new_n441), .ZN(new_n442));
  NOR3_X1   g241(.A1(new_n432), .A2(new_n433), .A3(new_n442), .ZN(new_n443));
  NAND3_X1  g242(.A1(new_n377), .A2(new_n379), .A3(new_n443), .ZN(new_n444));
  XNOR2_X1  g243(.A(G22gat), .B(G50gat), .ZN(new_n445));
  INV_X1    g244(.A(new_n445), .ZN(new_n446));
  NOR2_X1   g245(.A1(new_n395), .A2(KEYINPUT3), .ZN(new_n447));
  OAI21_X1  g246(.A(new_n356), .B1(new_n447), .B2(KEYINPUT29), .ZN(new_n448));
  AND2_X1   g247(.A1(new_n391), .A2(new_n394), .ZN(new_n449));
  AOI21_X1  g248(.A(KEYINPUT3), .B1(new_n335), .B2(new_n338), .ZN(new_n450));
  OAI21_X1  g249(.A(new_n448), .B1(new_n449), .B2(new_n450), .ZN(new_n451));
  NAND2_X1  g250(.A1(G228gat), .A2(G233gat), .ZN(new_n452));
  INV_X1    g251(.A(new_n452), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n451), .A2(new_n453), .ZN(new_n454));
  XNOR2_X1  g253(.A(new_n334), .B(KEYINPUT88), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n455), .A2(new_n333), .ZN(new_n456));
  AOI21_X1  g255(.A(KEYINPUT3), .B1(new_n456), .B2(new_n338), .ZN(new_n457));
  OAI211_X1 g256(.A(new_n448), .B(new_n452), .C1(new_n449), .C2(new_n457), .ZN(new_n458));
  INV_X1    g257(.A(KEYINPUT31), .ZN(new_n459));
  NAND3_X1  g258(.A1(new_n454), .A2(new_n458), .A3(new_n459), .ZN(new_n460));
  INV_X1    g259(.A(new_n460), .ZN(new_n461));
  AOI21_X1  g260(.A(new_n459), .B1(new_n454), .B2(new_n458), .ZN(new_n462));
  XOR2_X1   g261(.A(G78gat), .B(G106gat), .Z(new_n463));
  NOR3_X1   g262(.A1(new_n461), .A2(new_n462), .A3(new_n463), .ZN(new_n464));
  INV_X1    g263(.A(new_n463), .ZN(new_n465));
  NAND2_X1  g264(.A1(new_n454), .A2(new_n458), .ZN(new_n466));
  NAND2_X1  g265(.A1(new_n466), .A2(KEYINPUT31), .ZN(new_n467));
  AOI21_X1  g266(.A(new_n465), .B1(new_n467), .B2(new_n460), .ZN(new_n468));
  OAI21_X1  g267(.A(new_n446), .B1(new_n464), .B2(new_n468), .ZN(new_n469));
  OAI21_X1  g268(.A(new_n463), .B1(new_n461), .B2(new_n462), .ZN(new_n470));
  NAND3_X1  g269(.A1(new_n467), .A2(new_n460), .A3(new_n465), .ZN(new_n471));
  NAND3_X1  g270(.A1(new_n470), .A2(new_n471), .A3(new_n445), .ZN(new_n472));
  NAND2_X1  g271(.A1(new_n469), .A2(new_n472), .ZN(new_n473));
  INV_X1    g272(.A(new_n473), .ZN(new_n474));
  NAND2_X1  g273(.A1(new_n363), .A2(KEYINPUT37), .ZN(new_n475));
  INV_X1    g274(.A(KEYINPUT37), .ZN(new_n476));
  NAND4_X1  g275(.A1(new_n342), .A2(new_n353), .A3(new_n476), .A4(new_n362), .ZN(new_n477));
  NAND4_X1  g276(.A1(new_n475), .A2(KEYINPUT38), .A3(new_n368), .A4(new_n477), .ZN(new_n478));
  NAND4_X1  g277(.A1(new_n349), .A2(new_n356), .A3(new_n350), .A4(new_n341), .ZN(new_n479));
  NAND3_X1  g278(.A1(new_n355), .A2(new_n335), .A3(new_n357), .ZN(new_n480));
  NAND3_X1  g279(.A1(new_n479), .A2(KEYINPUT37), .A3(new_n480), .ZN(new_n481));
  INV_X1    g280(.A(KEYINPUT90), .ZN(new_n482));
  AOI21_X1  g281(.A(new_n369), .B1(new_n481), .B2(new_n482), .ZN(new_n483));
  NAND4_X1  g282(.A1(new_n479), .A2(KEYINPUT90), .A3(KEYINPUT37), .A4(new_n480), .ZN(new_n484));
  AND3_X1   g283(.A1(new_n483), .A2(new_n477), .A3(new_n484), .ZN(new_n485));
  INV_X1    g284(.A(KEYINPUT38), .ZN(new_n486));
  NAND2_X1  g285(.A1(new_n373), .A2(new_n486), .ZN(new_n487));
  OAI21_X1  g286(.A(new_n478), .B1(new_n485), .B2(new_n487), .ZN(new_n488));
  NAND3_X1  g287(.A1(new_n439), .A2(new_n441), .A3(new_n426), .ZN(new_n489));
  INV_X1    g288(.A(KEYINPUT6), .ZN(new_n490));
  NAND2_X1  g289(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  NOR2_X1   g290(.A1(new_n491), .A2(new_n442), .ZN(new_n492));
  AOI211_X1 g291(.A(new_n490), .B(new_n426), .C1(new_n439), .C2(new_n441), .ZN(new_n493));
  NOR2_X1   g292(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  AOI21_X1  g293(.A(new_n474), .B1(new_n488), .B2(new_n494), .ZN(new_n495));
  NAND2_X1  g294(.A1(new_n444), .A2(new_n495), .ZN(new_n496));
  AOI21_X1  g295(.A(new_n494), .B1(new_n374), .B2(new_n375), .ZN(new_n497));
  NAND2_X1  g296(.A1(new_n314), .A2(new_n404), .ZN(new_n498));
  OAI211_X1 g297(.A(new_n403), .B(new_n273), .C1(new_n312), .C2(new_n313), .ZN(new_n499));
  NAND2_X1  g298(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  INV_X1    g299(.A(G227gat), .ZN(new_n501));
  INV_X1    g300(.A(G233gat), .ZN(new_n502));
  NOR2_X1   g301(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  NOR2_X1   g302(.A1(new_n500), .A2(new_n503), .ZN(new_n504));
  INV_X1    g303(.A(new_n504), .ZN(new_n505));
  INV_X1    g304(.A(KEYINPUT34), .ZN(new_n506));
  NAND2_X1  g305(.A1(new_n500), .A2(new_n503), .ZN(new_n507));
  XNOR2_X1  g306(.A(G15gat), .B(G43gat), .ZN(new_n508));
  XNOR2_X1  g307(.A(new_n508), .B(G71gat), .ZN(new_n509));
  INV_X1    g308(.A(G99gat), .ZN(new_n510));
  XNOR2_X1  g309(.A(new_n509), .B(new_n510), .ZN(new_n511));
  NAND2_X1  g310(.A1(new_n511), .A2(KEYINPUT33), .ZN(new_n512));
  NAND3_X1  g311(.A1(new_n507), .A2(KEYINPUT32), .A3(new_n512), .ZN(new_n513));
  INV_X1    g312(.A(KEYINPUT74), .ZN(new_n514));
  NAND2_X1  g313(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  INV_X1    g314(.A(new_n503), .ZN(new_n516));
  AOI21_X1  g315(.A(new_n516), .B1(new_n498), .B2(new_n499), .ZN(new_n517));
  INV_X1    g316(.A(KEYINPUT32), .ZN(new_n518));
  NOR2_X1   g317(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  NAND3_X1  g318(.A1(new_n519), .A2(KEYINPUT74), .A3(new_n512), .ZN(new_n520));
  NAND2_X1  g319(.A1(new_n515), .A2(new_n520), .ZN(new_n521));
  INV_X1    g320(.A(new_n511), .ZN(new_n522));
  NAND2_X1  g321(.A1(new_n518), .A2(KEYINPUT33), .ZN(new_n523));
  AOI21_X1  g322(.A(new_n522), .B1(new_n507), .B2(new_n523), .ZN(new_n524));
  INV_X1    g323(.A(new_n524), .ZN(new_n525));
  AOI21_X1  g324(.A(new_n506), .B1(new_n521), .B2(new_n525), .ZN(new_n526));
  AOI211_X1 g325(.A(KEYINPUT34), .B(new_n524), .C1(new_n515), .C2(new_n520), .ZN(new_n527));
  OAI21_X1  g326(.A(new_n505), .B1(new_n526), .B2(new_n527), .ZN(new_n528));
  AOI21_X1  g327(.A(KEYINPUT74), .B1(new_n519), .B2(new_n512), .ZN(new_n529));
  INV_X1    g328(.A(new_n512), .ZN(new_n530));
  NOR4_X1   g329(.A1(new_n517), .A2(new_n514), .A3(new_n518), .A4(new_n530), .ZN(new_n531));
  OAI21_X1  g330(.A(new_n525), .B1(new_n529), .B2(new_n531), .ZN(new_n532));
  NAND2_X1  g331(.A1(new_n532), .A2(KEYINPUT34), .ZN(new_n533));
  NAND3_X1  g332(.A1(new_n521), .A2(new_n506), .A3(new_n525), .ZN(new_n534));
  NAND3_X1  g333(.A1(new_n533), .A2(new_n534), .A3(new_n504), .ZN(new_n535));
  AND3_X1   g334(.A1(new_n528), .A2(KEYINPUT36), .A3(new_n535), .ZN(new_n536));
  AOI21_X1  g335(.A(KEYINPUT36), .B1(new_n528), .B2(new_n535), .ZN(new_n537));
  OAI22_X1  g336(.A1(new_n497), .A2(new_n473), .B1(new_n536), .B2(new_n537), .ZN(new_n538));
  INV_X1    g337(.A(new_n538), .ZN(new_n539));
  NAND2_X1  g338(.A1(new_n496), .A2(new_n539), .ZN(new_n540));
  XNOR2_X1  g339(.A(new_n491), .B(new_n442), .ZN(new_n541));
  NAND2_X1  g340(.A1(new_n376), .A2(new_n541), .ZN(new_n542));
  NAND4_X1  g341(.A1(new_n473), .A2(KEYINPUT35), .A3(new_n535), .A4(new_n528), .ZN(new_n543));
  NOR2_X1   g342(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  AND4_X1   g343(.A1(new_n541), .A2(new_n473), .A3(new_n535), .A4(new_n528), .ZN(new_n545));
  INV_X1    g344(.A(new_n379), .ZN(new_n546));
  AOI21_X1  g345(.A(new_n378), .B1(new_n374), .B2(new_n375), .ZN(new_n547));
  OAI21_X1  g346(.A(new_n545), .B1(new_n546), .B2(new_n547), .ZN(new_n548));
  INV_X1    g347(.A(KEYINPUT35), .ZN(new_n549));
  AOI21_X1  g348(.A(new_n544), .B1(new_n548), .B2(new_n549), .ZN(new_n550));
  AOI21_X1  g349(.A(new_n247), .B1(new_n540), .B2(new_n550), .ZN(new_n551));
  NAND2_X1  g350(.A1(G85gat), .A2(G92gat), .ZN(new_n552));
  XNOR2_X1  g351(.A(new_n552), .B(KEYINPUT7), .ZN(new_n553));
  NAND2_X1  g352(.A1(G99gat), .A2(G106gat), .ZN(new_n554));
  AOI22_X1  g353(.A1(KEYINPUT8), .A2(new_n554), .B1(new_n425), .B2(new_n367), .ZN(new_n555));
  NAND2_X1  g354(.A1(new_n553), .A2(new_n555), .ZN(new_n556));
  XNOR2_X1  g355(.A(G99gat), .B(G106gat), .ZN(new_n557));
  XOR2_X1   g356(.A(new_n556), .B(new_n557), .Z(new_n558));
  NAND2_X1  g357(.A1(new_n218), .A2(new_n558), .ZN(new_n559));
  INV_X1    g358(.A(new_n558), .ZN(new_n560));
  NAND2_X1  g359(.A1(new_n217), .A2(new_n560), .ZN(new_n561));
  NAND3_X1  g360(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n562));
  NAND3_X1  g361(.A1(new_n559), .A2(new_n561), .A3(new_n562), .ZN(new_n563));
  XNOR2_X1  g362(.A(G190gat), .B(G218gat), .ZN(new_n564));
  OR2_X1    g363(.A1(new_n563), .A2(new_n564), .ZN(new_n565));
  XNOR2_X1  g364(.A(new_n565), .B(KEYINPUT103), .ZN(new_n566));
  NAND2_X1  g365(.A1(new_n563), .A2(new_n564), .ZN(new_n567));
  XOR2_X1   g366(.A(new_n567), .B(KEYINPUT104), .Z(new_n568));
  NAND2_X1  g367(.A1(new_n566), .A2(new_n568), .ZN(new_n569));
  INV_X1    g368(.A(KEYINPUT41), .ZN(new_n570));
  INV_X1    g369(.A(G232gat), .ZN(new_n571));
  OAI21_X1  g370(.A(new_n570), .B1(new_n571), .B2(new_n502), .ZN(new_n572));
  XNOR2_X1  g371(.A(new_n569), .B(new_n572), .ZN(new_n573));
  AND2_X1   g372(.A1(new_n573), .A2(new_n402), .ZN(new_n574));
  NOR2_X1   g373(.A1(new_n573), .A2(new_n402), .ZN(new_n575));
  OAI21_X1  g374(.A(new_n381), .B1(new_n574), .B2(new_n575), .ZN(new_n576));
  XOR2_X1   g375(.A(new_n569), .B(new_n572), .Z(new_n577));
  NAND2_X1  g376(.A1(new_n577), .A2(G134gat), .ZN(new_n578));
  NAND2_X1  g377(.A1(new_n573), .A2(new_n402), .ZN(new_n579));
  NAND3_X1  g378(.A1(new_n578), .A2(G162gat), .A3(new_n579), .ZN(new_n580));
  NAND2_X1  g379(.A1(new_n576), .A2(new_n580), .ZN(new_n581));
  INV_X1    g380(.A(G57gat), .ZN(new_n582));
  OR3_X1    g381(.A1(new_n582), .A2(KEYINPUT99), .A3(G64gat), .ZN(new_n583));
  OAI21_X1  g382(.A(KEYINPUT99), .B1(new_n582), .B2(G64gat), .ZN(new_n584));
  OAI211_X1 g383(.A(new_n583), .B(new_n584), .C1(G57gat), .C2(new_n365), .ZN(new_n585));
  XOR2_X1   g384(.A(G71gat), .B(G78gat), .Z(new_n586));
  INV_X1    g385(.A(new_n586), .ZN(new_n587));
  INV_X1    g386(.A(KEYINPUT9), .ZN(new_n588));
  INV_X1    g387(.A(G71gat), .ZN(new_n589));
  INV_X1    g388(.A(G78gat), .ZN(new_n590));
  OAI21_X1  g389(.A(new_n588), .B1(new_n589), .B2(new_n590), .ZN(new_n591));
  NAND2_X1  g390(.A1(new_n591), .A2(KEYINPUT100), .ZN(new_n592));
  OR2_X1    g391(.A1(new_n591), .A2(KEYINPUT100), .ZN(new_n593));
  NAND4_X1  g392(.A1(new_n585), .A2(new_n587), .A3(new_n592), .A4(new_n593), .ZN(new_n594));
  XNOR2_X1  g393(.A(G57gat), .B(G64gat), .ZN(new_n595));
  OAI21_X1  g394(.A(new_n586), .B1(new_n588), .B2(new_n595), .ZN(new_n596));
  NAND2_X1  g395(.A1(new_n594), .A2(new_n596), .ZN(new_n597));
  INV_X1    g396(.A(KEYINPUT21), .ZN(new_n598));
  NAND2_X1  g397(.A1(new_n597), .A2(new_n598), .ZN(new_n599));
  XNOR2_X1  g398(.A(G127gat), .B(G155gat), .ZN(new_n600));
  XNOR2_X1  g399(.A(new_n599), .B(new_n600), .ZN(new_n601));
  XNOR2_X1  g400(.A(G183gat), .B(G211gat), .ZN(new_n602));
  XOR2_X1   g401(.A(new_n601), .B(new_n602), .Z(new_n603));
  NAND2_X1  g402(.A1(G231gat), .A2(G233gat), .ZN(new_n604));
  XOR2_X1   g403(.A(new_n603), .B(new_n604), .Z(new_n605));
  OAI21_X1  g404(.A(new_n227), .B1(new_n598), .B2(new_n597), .ZN(new_n606));
  XNOR2_X1  g405(.A(KEYINPUT102), .B(KEYINPUT20), .ZN(new_n607));
  XNOR2_X1  g406(.A(new_n606), .B(new_n607), .ZN(new_n608));
  XOR2_X1   g407(.A(KEYINPUT101), .B(KEYINPUT19), .Z(new_n609));
  XNOR2_X1  g408(.A(new_n608), .B(new_n609), .ZN(new_n610));
  XNOR2_X1  g409(.A(new_n605), .B(new_n610), .ZN(new_n611));
  INV_X1    g410(.A(new_n611), .ZN(new_n612));
  INV_X1    g411(.A(KEYINPUT10), .ZN(new_n613));
  NOR3_X1   g412(.A1(new_n558), .A2(new_n613), .A3(new_n597), .ZN(new_n614));
  AOI22_X1  g413(.A1(new_n560), .A2(KEYINPUT105), .B1(new_n596), .B2(new_n594), .ZN(new_n615));
  NOR2_X1   g414(.A1(new_n560), .A2(KEYINPUT105), .ZN(new_n616));
  XOR2_X1   g415(.A(new_n615), .B(new_n616), .Z(new_n617));
  AOI21_X1  g416(.A(new_n614), .B1(new_n617), .B2(new_n613), .ZN(new_n618));
  NAND2_X1  g417(.A1(G230gat), .A2(G233gat), .ZN(new_n619));
  INV_X1    g418(.A(new_n619), .ZN(new_n620));
  OR2_X1    g419(.A1(new_n618), .A2(new_n620), .ZN(new_n621));
  OAI21_X1  g420(.A(new_n621), .B1(new_n619), .B2(new_n617), .ZN(new_n622));
  XNOR2_X1  g421(.A(G120gat), .B(G148gat), .ZN(new_n623));
  XNOR2_X1  g422(.A(new_n623), .B(G176gat), .ZN(new_n624));
  XNOR2_X1  g423(.A(new_n624), .B(G204gat), .ZN(new_n625));
  XNOR2_X1  g424(.A(new_n622), .B(new_n625), .ZN(new_n626));
  XOR2_X1   g425(.A(new_n626), .B(KEYINPUT106), .Z(new_n627));
  INV_X1    g426(.A(new_n627), .ZN(new_n628));
  NOR3_X1   g427(.A1(new_n581), .A2(new_n612), .A3(new_n628), .ZN(new_n629));
  NAND2_X1  g428(.A1(new_n551), .A2(new_n629), .ZN(new_n630));
  NOR2_X1   g429(.A1(new_n630), .A2(new_n541), .ZN(new_n631));
  XNOR2_X1  g430(.A(new_n631), .B(new_n220), .ZN(G1324gat));
  INV_X1    g431(.A(new_n630), .ZN(new_n633));
  NOR2_X1   g432(.A1(new_n546), .A2(new_n547), .ZN(new_n634));
  NAND2_X1  g433(.A1(KEYINPUT16), .A2(G8gat), .ZN(new_n635));
  NAND3_X1  g434(.A1(new_n633), .A2(new_n634), .A3(new_n635), .ZN(new_n636));
  INV_X1    g435(.A(new_n636), .ZN(new_n637));
  OAI21_X1  g436(.A(new_n637), .B1(KEYINPUT16), .B2(G8gat), .ZN(new_n638));
  INV_X1    g437(.A(new_n634), .ZN(new_n639));
  OAI21_X1  g438(.A(G8gat), .B1(new_n630), .B2(new_n639), .ZN(new_n640));
  NAND2_X1  g439(.A1(new_n638), .A2(new_n640), .ZN(new_n641));
  MUX2_X1   g440(.A(new_n638), .B(new_n641), .S(KEYINPUT42), .Z(G1325gat));
  NOR2_X1   g441(.A1(new_n536), .A2(new_n537), .ZN(new_n643));
  AND3_X1   g442(.A1(new_n633), .A2(G15gat), .A3(new_n643), .ZN(new_n644));
  INV_X1    g443(.A(new_n528), .ZN(new_n645));
  INV_X1    g444(.A(new_n535), .ZN(new_n646));
  NOR2_X1   g445(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  AOI21_X1  g446(.A(G15gat), .B1(new_n633), .B2(new_n647), .ZN(new_n648));
  NOR2_X1   g447(.A1(new_n644), .A2(new_n648), .ZN(G1326gat));
  NOR2_X1   g448(.A1(new_n630), .A2(new_n473), .ZN(new_n650));
  XOR2_X1   g449(.A(KEYINPUT43), .B(G22gat), .Z(new_n651));
  XNOR2_X1  g450(.A(new_n650), .B(new_n651), .ZN(G1327gat));
  NAND3_X1  g451(.A1(new_n581), .A2(new_n612), .A3(new_n627), .ZN(new_n653));
  INV_X1    g452(.A(KEYINPUT107), .ZN(new_n654));
  OR2_X1    g453(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  NAND2_X1  g454(.A1(new_n655), .A2(new_n551), .ZN(new_n656));
  AOI21_X1  g455(.A(new_n656), .B1(new_n654), .B2(new_n653), .ZN(new_n657));
  INV_X1    g456(.A(G29gat), .ZN(new_n658));
  NAND3_X1  g457(.A1(new_n657), .A2(new_n658), .A3(new_n494), .ZN(new_n659));
  XOR2_X1   g458(.A(KEYINPUT108), .B(KEYINPUT45), .Z(new_n660));
  XNOR2_X1  g459(.A(new_n659), .B(new_n660), .ZN(new_n661));
  NOR3_X1   g460(.A1(new_n247), .A2(new_n611), .A3(new_n628), .ZN(new_n662));
  INV_X1    g461(.A(KEYINPUT44), .ZN(new_n663));
  NAND2_X1  g462(.A1(new_n581), .A2(new_n663), .ZN(new_n664));
  NAND4_X1  g463(.A1(new_n541), .A2(new_n473), .A3(new_n535), .A4(new_n528), .ZN(new_n665));
  AOI21_X1  g464(.A(new_n665), .B1(new_n377), .B2(new_n379), .ZN(new_n666));
  OAI22_X1  g465(.A1(new_n666), .A2(KEYINPUT35), .B1(new_n542), .B2(new_n543), .ZN(new_n667));
  AOI21_X1  g466(.A(new_n538), .B1(new_n495), .B2(new_n444), .ZN(new_n668));
  OAI21_X1  g467(.A(KEYINPUT109), .B1(new_n667), .B2(new_n668), .ZN(new_n669));
  INV_X1    g468(.A(KEYINPUT109), .ZN(new_n670));
  NAND3_X1  g469(.A1(new_n540), .A2(new_n670), .A3(new_n550), .ZN(new_n671));
  AOI21_X1  g470(.A(new_n664), .B1(new_n669), .B2(new_n671), .ZN(new_n672));
  NAND2_X1  g471(.A1(new_n540), .A2(new_n550), .ZN(new_n673));
  AOI21_X1  g472(.A(new_n663), .B1(new_n673), .B2(new_n581), .ZN(new_n674));
  OAI21_X1  g473(.A(new_n662), .B1(new_n672), .B2(new_n674), .ZN(new_n675));
  INV_X1    g474(.A(KEYINPUT110), .ZN(new_n676));
  NAND2_X1  g475(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  OAI211_X1 g476(.A(KEYINPUT110), .B(new_n662), .C1(new_n672), .C2(new_n674), .ZN(new_n678));
  AOI21_X1  g477(.A(new_n541), .B1(new_n677), .B2(new_n678), .ZN(new_n679));
  OAI21_X1  g478(.A(new_n661), .B1(new_n658), .B2(new_n679), .ZN(G1328gat));
  INV_X1    g479(.A(G36gat), .ZN(new_n681));
  NAND3_X1  g480(.A1(new_n657), .A2(new_n681), .A3(new_n634), .ZN(new_n682));
  XOR2_X1   g481(.A(new_n682), .B(KEYINPUT46), .Z(new_n683));
  AOI21_X1  g482(.A(new_n639), .B1(new_n677), .B2(new_n678), .ZN(new_n684));
  OAI21_X1  g483(.A(new_n683), .B1(new_n681), .B2(new_n684), .ZN(G1329gat));
  INV_X1    g484(.A(new_n664), .ZN(new_n686));
  NOR3_X1   g485(.A1(new_n667), .A2(new_n668), .A3(KEYINPUT109), .ZN(new_n687));
  AOI21_X1  g486(.A(new_n670), .B1(new_n540), .B2(new_n550), .ZN(new_n688));
  OAI21_X1  g487(.A(new_n686), .B1(new_n687), .B2(new_n688), .ZN(new_n689));
  NAND2_X1  g488(.A1(new_n673), .A2(new_n581), .ZN(new_n690));
  NAND2_X1  g489(.A1(new_n690), .A2(KEYINPUT44), .ZN(new_n691));
  NAND2_X1  g490(.A1(new_n689), .A2(new_n691), .ZN(new_n692));
  AOI21_X1  g491(.A(KEYINPUT110), .B1(new_n692), .B2(new_n662), .ZN(new_n693));
  INV_X1    g492(.A(new_n678), .ZN(new_n694));
  OAI21_X1  g493(.A(new_n643), .B1(new_n693), .B2(new_n694), .ZN(new_n695));
  INV_X1    g494(.A(KEYINPUT112), .ZN(new_n696));
  NAND3_X1  g495(.A1(new_n695), .A2(new_n696), .A3(G43gat), .ZN(new_n697));
  INV_X1    g496(.A(new_n643), .ZN(new_n698));
  AOI21_X1  g497(.A(new_n698), .B1(new_n677), .B2(new_n678), .ZN(new_n699));
  INV_X1    g498(.A(G43gat), .ZN(new_n700));
  OAI21_X1  g499(.A(KEYINPUT112), .B1(new_n699), .B2(new_n700), .ZN(new_n701));
  NAND3_X1  g500(.A1(new_n657), .A2(new_n700), .A3(new_n647), .ZN(new_n702));
  NAND3_X1  g501(.A1(new_n697), .A2(new_n701), .A3(new_n702), .ZN(new_n703));
  XNOR2_X1  g502(.A(KEYINPUT111), .B(KEYINPUT47), .ZN(new_n704));
  NAND2_X1  g503(.A1(new_n703), .A2(new_n704), .ZN(new_n705));
  OAI21_X1  g504(.A(G43gat), .B1(new_n675), .B2(new_n698), .ZN(new_n706));
  NAND3_X1  g505(.A1(new_n702), .A2(KEYINPUT47), .A3(new_n706), .ZN(new_n707));
  NAND2_X1  g506(.A1(new_n705), .A2(new_n707), .ZN(G1330gat));
  INV_X1    g507(.A(G50gat), .ZN(new_n709));
  NAND3_X1  g508(.A1(new_n657), .A2(new_n709), .A3(new_n474), .ZN(new_n710));
  OAI21_X1  g509(.A(G50gat), .B1(new_n675), .B2(new_n473), .ZN(new_n711));
  NAND3_X1  g510(.A1(new_n710), .A2(KEYINPUT48), .A3(new_n711), .ZN(new_n712));
  OAI21_X1  g511(.A(new_n474), .B1(new_n693), .B2(new_n694), .ZN(new_n713));
  NAND2_X1  g512(.A1(new_n713), .A2(G50gat), .ZN(new_n714));
  AND2_X1   g513(.A1(new_n714), .A2(new_n710), .ZN(new_n715));
  OAI21_X1  g514(.A(new_n712), .B1(new_n715), .B2(KEYINPUT48), .ZN(G1331gat));
  NOR2_X1   g515(.A1(new_n581), .A2(new_n612), .ZN(new_n717));
  NOR2_X1   g516(.A1(new_n246), .A2(new_n627), .ZN(new_n718));
  OAI211_X1 g517(.A(new_n717), .B(new_n718), .C1(new_n687), .C2(new_n688), .ZN(new_n719));
  OR2_X1    g518(.A1(new_n719), .A2(KEYINPUT113), .ZN(new_n720));
  NAND2_X1  g519(.A1(new_n719), .A2(KEYINPUT113), .ZN(new_n721));
  NAND2_X1  g520(.A1(new_n720), .A2(new_n721), .ZN(new_n722));
  NOR2_X1   g521(.A1(new_n722), .A2(new_n541), .ZN(new_n723));
  XNOR2_X1  g522(.A(new_n723), .B(new_n582), .ZN(G1332gat));
  NOR2_X1   g523(.A1(new_n722), .A2(new_n639), .ZN(new_n725));
  NOR2_X1   g524(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n726));
  AND2_X1   g525(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n727));
  OAI21_X1  g526(.A(new_n725), .B1(new_n726), .B2(new_n727), .ZN(new_n728));
  OAI21_X1  g527(.A(new_n728), .B1(new_n725), .B2(new_n726), .ZN(G1333gat));
  INV_X1    g528(.A(new_n647), .ZN(new_n730));
  OAI21_X1  g529(.A(new_n589), .B1(new_n722), .B2(new_n730), .ZN(new_n731));
  NAND4_X1  g530(.A1(new_n720), .A2(G71gat), .A3(new_n643), .A4(new_n721), .ZN(new_n732));
  NAND2_X1  g531(.A1(new_n731), .A2(new_n732), .ZN(new_n733));
  XNOR2_X1  g532(.A(new_n733), .B(KEYINPUT50), .ZN(G1334gat));
  NOR2_X1   g533(.A1(new_n722), .A2(new_n473), .ZN(new_n735));
  XOR2_X1   g534(.A(KEYINPUT114), .B(G78gat), .Z(new_n736));
  XNOR2_X1  g535(.A(new_n735), .B(new_n736), .ZN(G1335gat));
  NAND2_X1  g536(.A1(new_n247), .A2(new_n612), .ZN(new_n738));
  AOI21_X1  g537(.A(new_n738), .B1(new_n689), .B2(new_n691), .ZN(new_n739));
  NOR2_X1   g538(.A1(new_n627), .A2(new_n541), .ZN(new_n740));
  NAND2_X1  g539(.A1(new_n739), .A2(new_n740), .ZN(new_n741));
  NAND2_X1  g540(.A1(new_n741), .A2(G85gat), .ZN(new_n742));
  INV_X1    g541(.A(new_n738), .ZN(new_n743));
  NAND3_X1  g542(.A1(new_n673), .A2(new_n743), .A3(new_n581), .ZN(new_n744));
  INV_X1    g543(.A(KEYINPUT51), .ZN(new_n745));
  OR2_X1    g544(.A1(new_n744), .A2(new_n745), .ZN(new_n746));
  OR2_X1    g545(.A1(new_n746), .A2(KEYINPUT115), .ZN(new_n747));
  NAND2_X1  g546(.A1(new_n744), .A2(new_n745), .ZN(new_n748));
  NAND3_X1  g547(.A1(new_n746), .A2(KEYINPUT115), .A3(new_n748), .ZN(new_n749));
  AND3_X1   g548(.A1(new_n747), .A2(KEYINPUT116), .A3(new_n749), .ZN(new_n750));
  AOI21_X1  g549(.A(KEYINPUT116), .B1(new_n747), .B2(new_n749), .ZN(new_n751));
  NOR2_X1   g550(.A1(new_n750), .A2(new_n751), .ZN(new_n752));
  NAND2_X1  g551(.A1(new_n740), .A2(new_n425), .ZN(new_n753));
  OAI21_X1  g552(.A(new_n742), .B1(new_n752), .B2(new_n753), .ZN(G1336gat));
  NOR2_X1   g553(.A1(new_n639), .A2(new_n627), .ZN(new_n755));
  NAND2_X1  g554(.A1(new_n739), .A2(new_n755), .ZN(new_n756));
  OR2_X1    g555(.A1(new_n756), .A2(KEYINPUT119), .ZN(new_n757));
  NAND2_X1  g556(.A1(new_n756), .A2(KEYINPUT119), .ZN(new_n758));
  NAND3_X1  g557(.A1(new_n757), .A2(G92gat), .A3(new_n758), .ZN(new_n759));
  INV_X1    g558(.A(KEYINPUT52), .ZN(new_n760));
  NAND2_X1  g559(.A1(new_n747), .A2(new_n749), .ZN(new_n761));
  NAND2_X1  g560(.A1(new_n755), .A2(new_n367), .ZN(new_n762));
  OAI211_X1 g561(.A(new_n759), .B(new_n760), .C1(new_n761), .C2(new_n762), .ZN(new_n763));
  AOI211_X1 g562(.A(KEYINPUT117), .B(new_n367), .C1(new_n739), .C2(new_n755), .ZN(new_n764));
  INV_X1    g563(.A(KEYINPUT117), .ZN(new_n765));
  AOI21_X1  g564(.A(new_n765), .B1(new_n756), .B2(G92gat), .ZN(new_n766));
  NAND2_X1  g565(.A1(new_n746), .A2(new_n748), .ZN(new_n767));
  XOR2_X1   g566(.A(new_n762), .B(KEYINPUT118), .Z(new_n768));
  AOI211_X1 g567(.A(new_n764), .B(new_n766), .C1(new_n767), .C2(new_n768), .ZN(new_n769));
  OAI21_X1  g568(.A(new_n763), .B1(new_n769), .B2(new_n760), .ZN(G1337gat));
  OAI211_X1 g569(.A(new_n628), .B(new_n743), .C1(new_n672), .C2(new_n674), .ZN(new_n771));
  OR3_X1    g570(.A1(new_n771), .A2(KEYINPUT120), .A3(new_n698), .ZN(new_n772));
  OAI21_X1  g571(.A(KEYINPUT120), .B1(new_n771), .B2(new_n698), .ZN(new_n773));
  NAND3_X1  g572(.A1(new_n772), .A2(G99gat), .A3(new_n773), .ZN(new_n774));
  OAI211_X1 g573(.A(new_n510), .B(new_n647), .C1(new_n750), .C2(new_n751), .ZN(new_n775));
  OAI21_X1  g574(.A(new_n774), .B1(new_n775), .B2(new_n627), .ZN(G1338gat));
  OAI21_X1  g575(.A(G106gat), .B1(new_n771), .B2(new_n473), .ZN(new_n777));
  OR2_X1    g576(.A1(new_n777), .A2(KEYINPUT121), .ZN(new_n778));
  NOR3_X1   g577(.A1(new_n627), .A2(G106gat), .A3(new_n473), .ZN(new_n779));
  NAND2_X1  g578(.A1(new_n767), .A2(new_n779), .ZN(new_n780));
  NAND2_X1  g579(.A1(new_n777), .A2(KEYINPUT121), .ZN(new_n781));
  AND3_X1   g580(.A1(new_n778), .A2(new_n780), .A3(new_n781), .ZN(new_n782));
  INV_X1    g581(.A(KEYINPUT53), .ZN(new_n783));
  INV_X1    g582(.A(new_n777), .ZN(new_n784));
  INV_X1    g583(.A(new_n779), .ZN(new_n785));
  OAI21_X1  g584(.A(new_n783), .B1(new_n761), .B2(new_n785), .ZN(new_n786));
  OAI22_X1  g585(.A1(new_n782), .A2(new_n783), .B1(new_n784), .B2(new_n786), .ZN(G1339gat));
  NAND2_X1  g586(.A1(new_n618), .A2(new_n620), .ZN(new_n788));
  NAND3_X1  g587(.A1(new_n621), .A2(KEYINPUT54), .A3(new_n788), .ZN(new_n789));
  OAI211_X1 g588(.A(new_n789), .B(new_n625), .C1(KEYINPUT54), .C2(new_n621), .ZN(new_n790));
  XOR2_X1   g589(.A(new_n790), .B(KEYINPUT55), .Z(new_n791));
  NOR2_X1   g590(.A1(new_n622), .A2(new_n625), .ZN(new_n792));
  NOR2_X1   g591(.A1(new_n791), .A2(new_n792), .ZN(new_n793));
  INV_X1    g592(.A(new_n793), .ZN(new_n794));
  NOR3_X1   g593(.A1(new_n574), .A2(new_n575), .A3(new_n381), .ZN(new_n795));
  AOI21_X1  g594(.A(G162gat), .B1(new_n578), .B2(new_n579), .ZN(new_n796));
  OAI21_X1  g595(.A(new_n794), .B1(new_n795), .B2(new_n796), .ZN(new_n797));
  NAND3_X1  g596(.A1(new_n576), .A2(new_n580), .A3(new_n627), .ZN(new_n798));
  INV_X1    g597(.A(new_n240), .ZN(new_n799));
  NAND2_X1  g598(.A1(new_n228), .A2(new_n230), .ZN(new_n800));
  NAND2_X1  g599(.A1(new_n233), .A2(new_n234), .ZN(new_n801));
  AOI21_X1  g600(.A(new_n799), .B1(new_n800), .B2(new_n801), .ZN(new_n802));
  INV_X1    g601(.A(new_n802), .ZN(new_n803));
  NAND2_X1  g602(.A1(new_n243), .A2(new_n803), .ZN(new_n804));
  INV_X1    g603(.A(new_n804), .ZN(new_n805));
  NAND3_X1  g604(.A1(new_n797), .A2(new_n798), .A3(new_n805), .ZN(new_n806));
  NOR2_X1   g605(.A1(new_n795), .A2(new_n796), .ZN(new_n807));
  NAND3_X1  g606(.A1(new_n807), .A2(new_n246), .A3(new_n793), .ZN(new_n808));
  AOI21_X1  g607(.A(new_n611), .B1(new_n806), .B2(new_n808), .ZN(new_n809));
  AND2_X1   g608(.A1(new_n629), .A2(new_n247), .ZN(new_n810));
  NOR2_X1   g609(.A1(new_n809), .A2(new_n810), .ZN(new_n811));
  NOR2_X1   g610(.A1(new_n811), .A2(new_n474), .ZN(new_n812));
  NOR2_X1   g611(.A1(new_n634), .A2(new_n541), .ZN(new_n813));
  AND2_X1   g612(.A1(new_n812), .A2(new_n813), .ZN(new_n814));
  NAND2_X1  g613(.A1(new_n814), .A2(new_n647), .ZN(new_n815));
  XNOR2_X1  g614(.A(KEYINPUT122), .B(G113gat), .ZN(new_n816));
  OR3_X1    g615(.A1(new_n815), .A2(new_n247), .A3(new_n816), .ZN(new_n817));
  OAI21_X1  g616(.A(new_n816), .B1(new_n815), .B2(new_n247), .ZN(new_n818));
  NAND2_X1  g617(.A1(new_n817), .A2(new_n818), .ZN(G1340gat));
  INV_X1    g618(.A(new_n815), .ZN(new_n820));
  NAND3_X1  g619(.A1(new_n820), .A2(new_n396), .A3(new_n628), .ZN(new_n821));
  OAI21_X1  g620(.A(G120gat), .B1(new_n815), .B2(new_n627), .ZN(new_n822));
  NAND2_X1  g621(.A1(new_n821), .A2(new_n822), .ZN(G1341gat));
  AOI21_X1  g622(.A(G127gat), .B1(new_n820), .B2(new_n611), .ZN(new_n824));
  INV_X1    g623(.A(G127gat), .ZN(new_n825));
  NOR3_X1   g624(.A1(new_n815), .A2(new_n825), .A3(new_n612), .ZN(new_n826));
  NOR2_X1   g625(.A1(new_n824), .A2(new_n826), .ZN(G1342gat));
  XOR2_X1   g626(.A(KEYINPUT56), .B(G134gat), .Z(new_n828));
  NAND3_X1  g627(.A1(new_n820), .A2(new_n581), .A3(new_n828), .ZN(new_n829));
  NOR2_X1   g628(.A1(KEYINPUT56), .A2(G134gat), .ZN(new_n830));
  OAI21_X1  g629(.A(new_n830), .B1(new_n815), .B2(new_n807), .ZN(new_n831));
  AND2_X1   g630(.A1(new_n829), .A2(new_n831), .ZN(G1343gat));
  OAI21_X1  g631(.A(new_n474), .B1(new_n809), .B2(new_n810), .ZN(new_n833));
  NAND2_X1  g632(.A1(new_n833), .A2(KEYINPUT57), .ZN(new_n834));
  INV_X1    g633(.A(KEYINPUT57), .ZN(new_n835));
  OAI211_X1 g634(.A(new_n835), .B(new_n474), .C1(new_n809), .C2(new_n810), .ZN(new_n836));
  NAND4_X1  g635(.A1(new_n834), .A2(new_n698), .A3(new_n813), .A4(new_n836), .ZN(new_n837));
  OAI21_X1  g636(.A(new_n386), .B1(new_n837), .B2(new_n247), .ZN(new_n838));
  NAND2_X1  g637(.A1(new_n629), .A2(new_n247), .ZN(new_n839));
  AOI21_X1  g638(.A(new_n804), .B1(new_n581), .B2(new_n794), .ZN(new_n840));
  NOR2_X1   g639(.A1(new_n581), .A2(new_n247), .ZN(new_n841));
  AOI22_X1  g640(.A1(new_n840), .A2(new_n798), .B1(new_n841), .B2(new_n793), .ZN(new_n842));
  OAI21_X1  g641(.A(new_n839), .B1(new_n842), .B2(new_n611), .ZN(new_n843));
  NAND3_X1  g642(.A1(new_n843), .A2(new_n474), .A3(new_n698), .ZN(new_n844));
  INV_X1    g643(.A(new_n844), .ZN(new_n845));
  INV_X1    g644(.A(G141gat), .ZN(new_n846));
  NAND4_X1  g645(.A1(new_n845), .A2(new_n846), .A3(new_n246), .A4(new_n813), .ZN(new_n847));
  NAND2_X1  g646(.A1(new_n838), .A2(new_n847), .ZN(new_n848));
  INV_X1    g647(.A(KEYINPUT58), .ZN(new_n849));
  INV_X1    g648(.A(KEYINPUT123), .ZN(new_n850));
  AOI21_X1  g649(.A(new_n849), .B1(new_n847), .B2(new_n850), .ZN(new_n851));
  NAND2_X1  g650(.A1(new_n848), .A2(new_n851), .ZN(new_n852));
  OAI211_X1 g651(.A(new_n838), .B(new_n847), .C1(new_n850), .C2(new_n849), .ZN(new_n853));
  NAND2_X1  g652(.A1(new_n852), .A2(new_n853), .ZN(G1344gat));
  NOR3_X1   g653(.A1(new_n844), .A2(new_n541), .A3(new_n634), .ZN(new_n855));
  NAND3_X1  g654(.A1(new_n855), .A2(new_n384), .A3(new_n628), .ZN(new_n856));
  OAI21_X1  g655(.A(G148gat), .B1(new_n837), .B2(new_n627), .ZN(new_n857));
  AND2_X1   g656(.A1(new_n857), .A2(KEYINPUT59), .ZN(new_n858));
  INV_X1    g657(.A(KEYINPUT59), .ZN(new_n859));
  OAI211_X1 g658(.A(new_n859), .B(G148gat), .C1(new_n837), .C2(new_n627), .ZN(new_n860));
  INV_X1    g659(.A(new_n860), .ZN(new_n861));
  OAI21_X1  g660(.A(new_n856), .B1(new_n858), .B2(new_n861), .ZN(G1345gat));
  OAI21_X1  g661(.A(G155gat), .B1(new_n837), .B2(new_n612), .ZN(new_n863));
  NAND3_X1  g662(.A1(new_n855), .A2(new_n380), .A3(new_n611), .ZN(new_n864));
  NAND2_X1  g663(.A1(new_n863), .A2(new_n864), .ZN(G1346gat));
  NOR2_X1   g664(.A1(new_n855), .A2(G162gat), .ZN(new_n866));
  NOR2_X1   g665(.A1(new_n574), .A2(new_n575), .ZN(new_n867));
  NAND2_X1  g666(.A1(new_n837), .A2(G162gat), .ZN(new_n868));
  AOI21_X1  g667(.A(new_n866), .B1(new_n867), .B2(new_n868), .ZN(G1347gat));
  NOR3_X1   g668(.A1(new_n639), .A2(new_n494), .A3(new_n730), .ZN(new_n870));
  OR2_X1    g669(.A1(new_n870), .A2(KEYINPUT124), .ZN(new_n871));
  NAND2_X1  g670(.A1(new_n870), .A2(KEYINPUT124), .ZN(new_n872));
  NAND3_X1  g671(.A1(new_n812), .A2(new_n871), .A3(new_n872), .ZN(new_n873));
  OAI21_X1  g672(.A(G169gat), .B1(new_n873), .B2(new_n247), .ZN(new_n874));
  NOR3_X1   g673(.A1(new_n811), .A2(new_n639), .A3(new_n665), .ZN(new_n875));
  NAND3_X1  g674(.A1(new_n875), .A2(new_n239), .A3(new_n246), .ZN(new_n876));
  NAND2_X1  g675(.A1(new_n874), .A2(new_n876), .ZN(G1348gat));
  OAI21_X1  g676(.A(G176gat), .B1(new_n873), .B2(new_n627), .ZN(new_n878));
  INV_X1    g677(.A(G176gat), .ZN(new_n879));
  NAND4_X1  g678(.A1(new_n843), .A2(new_n879), .A3(new_n545), .A4(new_n755), .ZN(new_n880));
  NAND2_X1  g679(.A1(new_n878), .A2(new_n880), .ZN(G1349gat));
  OAI21_X1  g680(.A(G183gat), .B1(new_n873), .B2(new_n612), .ZN(new_n882));
  AND2_X1   g681(.A1(new_n611), .A2(new_n270), .ZN(new_n883));
  AOI21_X1  g682(.A(KEYINPUT125), .B1(new_n875), .B2(new_n883), .ZN(new_n884));
  NAND2_X1  g683(.A1(new_n882), .A2(new_n884), .ZN(new_n885));
  NAND2_X1  g684(.A1(new_n885), .A2(KEYINPUT60), .ZN(new_n886));
  INV_X1    g685(.A(KEYINPUT60), .ZN(new_n887));
  NAND3_X1  g686(.A1(new_n882), .A2(new_n887), .A3(new_n884), .ZN(new_n888));
  NAND2_X1  g687(.A1(new_n886), .A2(new_n888), .ZN(G1350gat));
  NAND3_X1  g688(.A1(new_n875), .A2(new_n262), .A3(new_n581), .ZN(new_n890));
  NAND4_X1  g689(.A1(new_n812), .A2(new_n581), .A3(new_n871), .A4(new_n872), .ZN(new_n891));
  INV_X1    g690(.A(KEYINPUT61), .ZN(new_n892));
  AND3_X1   g691(.A1(new_n891), .A2(new_n892), .A3(G190gat), .ZN(new_n893));
  AOI21_X1  g692(.A(new_n892), .B1(new_n891), .B2(G190gat), .ZN(new_n894));
  OAI21_X1  g693(.A(new_n890), .B1(new_n893), .B2(new_n894), .ZN(G1351gat));
  NOR2_X1   g694(.A1(new_n639), .A2(new_n494), .ZN(new_n896));
  NAND4_X1  g695(.A1(new_n834), .A2(new_n698), .A3(new_n836), .A4(new_n896), .ZN(new_n897));
  OAI21_X1  g696(.A(G197gat), .B1(new_n897), .B2(new_n247), .ZN(new_n898));
  NOR3_X1   g697(.A1(new_n844), .A2(new_n494), .A3(new_n639), .ZN(new_n899));
  INV_X1    g698(.A(G197gat), .ZN(new_n900));
  NAND3_X1  g699(.A1(new_n899), .A2(new_n900), .A3(new_n246), .ZN(new_n901));
  NAND2_X1  g700(.A1(new_n898), .A2(new_n901), .ZN(G1352gat));
  INV_X1    g701(.A(new_n897), .ZN(new_n903));
  NAND3_X1  g702(.A1(new_n903), .A2(KEYINPUT127), .A3(new_n628), .ZN(new_n904));
  XNOR2_X1  g703(.A(KEYINPUT126), .B(G204gat), .ZN(new_n905));
  INV_X1    g704(.A(KEYINPUT127), .ZN(new_n906));
  OAI21_X1  g705(.A(new_n906), .B1(new_n897), .B2(new_n627), .ZN(new_n907));
  NAND3_X1  g706(.A1(new_n904), .A2(new_n905), .A3(new_n907), .ZN(new_n908));
  NAND3_X1  g707(.A1(new_n845), .A2(new_n628), .A3(new_n896), .ZN(new_n909));
  NOR2_X1   g708(.A1(new_n909), .A2(new_n905), .ZN(new_n910));
  NOR2_X1   g709(.A1(new_n910), .A2(KEYINPUT62), .ZN(new_n911));
  INV_X1    g710(.A(KEYINPUT62), .ZN(new_n912));
  NOR3_X1   g711(.A1(new_n909), .A2(new_n912), .A3(new_n905), .ZN(new_n913));
  OAI21_X1  g712(.A(new_n908), .B1(new_n911), .B2(new_n913), .ZN(G1353gat));
  NAND3_X1  g713(.A1(new_n899), .A2(new_n324), .A3(new_n611), .ZN(new_n915));
  OAI21_X1  g714(.A(G211gat), .B1(new_n897), .B2(new_n612), .ZN(new_n916));
  INV_X1    g715(.A(KEYINPUT63), .ZN(new_n917));
  AND2_X1   g716(.A1(new_n916), .A2(new_n917), .ZN(new_n918));
  OAI211_X1 g717(.A(KEYINPUT63), .B(G211gat), .C1(new_n897), .C2(new_n612), .ZN(new_n919));
  INV_X1    g718(.A(new_n919), .ZN(new_n920));
  OAI21_X1  g719(.A(new_n915), .B1(new_n918), .B2(new_n920), .ZN(G1354gat));
  AOI21_X1  g720(.A(G218gat), .B1(new_n899), .B2(new_n581), .ZN(new_n922));
  NOR3_X1   g721(.A1(new_n897), .A2(new_n325), .A3(new_n807), .ZN(new_n923));
  NOR2_X1   g722(.A1(new_n922), .A2(new_n923), .ZN(G1355gat));
endmodule


