

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365,
         n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376,
         n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387,
         n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398,
         n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409,
         n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420,
         n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431,
         n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442,
         n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453,
         n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464,
         n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475,
         n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486,
         n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497,
         n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508,
         n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585,
         n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596,
         n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607,
         n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618,
         n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629,
         n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640,
         n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651,
         n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662,
         n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673,
         n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684,
         n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695,
         n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706,
         n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717,
         n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728,
         n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739,
         n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750,
         n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, n761,
         n762, n763, n764, n765;

  XNOR2_X1 U376 ( .A(n420), .B(KEYINPUT1), .ZN(n560) );
  INV_X1 U377 ( .A(G953), .ZN(n753) );
  AND2_X1 U378 ( .A1(n375), .A2(n374), .ZN(n355) );
  NAND2_X2 U379 ( .A1(n405), .A2(n355), .ZN(n398) );
  AND2_X2 U380 ( .A1(n422), .A2(n421), .ZN(n405) );
  XNOR2_X2 U381 ( .A(n398), .B(n569), .ZN(n629) );
  NAND2_X2 U382 ( .A1(n473), .A2(n472), .ZN(n503) );
  OR2_X2 U383 ( .A1(n721), .A2(n360), .ZN(n413) );
  XNOR2_X2 U384 ( .A(n737), .B(n514), .ZN(n721) );
  XNOR2_X2 U385 ( .A(n406), .B(KEYINPUT33), .ZN(n681) );
  NAND2_X2 U386 ( .A1(n434), .A2(n435), .ZN(n406) );
  INV_X1 U387 ( .A(n630), .ZN(n751) );
  NAND2_X1 U388 ( .A1(n659), .A2(n686), .ZN(n581) );
  AND2_X1 U389 ( .A1(n452), .A2(n765), .ZN(n422) );
  OR2_X1 U390 ( .A1(n763), .A2(n566), .ZN(n374) );
  XNOR2_X1 U391 ( .A(n562), .B(KEYINPUT32), .ZN(n763) );
  XNOR2_X1 U392 ( .A(KEYINPUT106), .B(n568), .ZN(n765) );
  XNOR2_X1 U393 ( .A(n558), .B(n559), .ZN(n563) );
  NOR2_X1 U394 ( .A1(n685), .A2(n687), .ZN(n605) );
  INV_X1 U395 ( .A(n549), .ZN(n356) );
  XNOR2_X1 U396 ( .A(n501), .B(n482), .ZN(n635) );
  XNOR2_X1 U397 ( .A(n456), .B(n455), .ZN(n512) );
  XNOR2_X1 U398 ( .A(G119), .B(KEYINPUT90), .ZN(n479) );
  XNOR2_X1 U399 ( .A(G137), .B(KEYINPUT5), .ZN(n480) );
  XOR2_X1 U400 ( .A(G902), .B(KEYINPUT15), .Z(n626) );
  INV_X1 U401 ( .A(KEYINPUT113), .ZN(n603) );
  XNOR2_X1 U402 ( .A(G116), .B(KEYINPUT70), .ZN(n477) );
  BUF_X1 U403 ( .A(n503), .Z(n357) );
  NOR2_X2 U404 ( .A1(n631), .A2(n630), .ZN(n632) );
  BUF_X1 U405 ( .A(n629), .Z(n744) );
  BUF_X1 U406 ( .A(n728), .Z(n733) );
  NOR2_X1 U407 ( .A1(n764), .A2(n760), .ZN(n615) );
  OR2_X1 U408 ( .A1(G237), .A2(G902), .ZN(n517) );
  NAND2_X1 U409 ( .A1(n416), .A2(n626), .ZN(n415) );
  INV_X1 U410 ( .A(KEYINPUT4), .ZN(n474) );
  XNOR2_X1 U411 ( .A(KEYINPUT102), .B(n546), .ZN(n591) );
  XNOR2_X1 U412 ( .A(n533), .B(n407), .ZN(n535) );
  XNOR2_X1 U413 ( .A(n534), .B(n408), .ZN(n407) );
  XNOR2_X1 U414 ( .A(n493), .B(n492), .ZN(n564) );
  XNOR2_X1 U415 ( .A(n491), .B(n490), .ZN(n492) );
  XNOR2_X1 U416 ( .A(n376), .B(n423), .ZN(n375) );
  INV_X1 U417 ( .A(KEYINPUT105), .ZN(n423) );
  INV_X1 U418 ( .A(G143), .ZN(n471) );
  AND2_X1 U419 ( .A1(n616), .A2(n367), .ZN(n464) );
  INV_X1 U420 ( .A(KEYINPUT48), .ZN(n462) );
  NAND2_X1 U421 ( .A1(n502), .A2(n393), .ZN(n392) );
  INV_X1 U422 ( .A(G902), .ZN(n393) );
  NOR2_X1 U423 ( .A1(G953), .A2(G237), .ZN(n530) );
  XNOR2_X1 U424 ( .A(n478), .B(G113), .ZN(n455) );
  XNOR2_X1 U425 ( .A(n477), .B(n479), .ZN(n456) );
  INV_X1 U426 ( .A(KEYINPUT3), .ZN(n478) );
  NAND2_X1 U427 ( .A1(G234), .A2(G237), .ZN(n518) );
  NAND2_X1 U428 ( .A1(n721), .A2(n682), .ZN(n381) );
  NAND2_X1 U429 ( .A1(n360), .A2(n682), .ZN(n380) );
  NOR2_X1 U430 ( .A1(n359), .A2(n417), .ZN(n411) );
  AND2_X1 U431 ( .A1(n382), .A2(n415), .ZN(n414) );
  AND2_X1 U432 ( .A1(n384), .A2(n359), .ZN(n383) );
  OR2_X1 U433 ( .A1(n721), .A2(n385), .ZN(n378) );
  NAND2_X1 U434 ( .A1(n415), .A2(n516), .ZN(n384) );
  XNOR2_X1 U435 ( .A(n460), .B(n497), .ZN(n499) );
  XNOR2_X1 U436 ( .A(n498), .B(n461), .ZN(n460) );
  NOR2_X1 U437 ( .A1(n610), .A2(n609), .ZN(n611) );
  XNOR2_X1 U438 ( .A(n538), .B(n537), .ZN(n556) );
  INV_X1 U439 ( .A(KEYINPUT6), .ZN(n429) );
  INV_X1 U440 ( .A(n564), .ZN(n694) );
  XNOR2_X1 U441 ( .A(n467), .B(n465), .ZN(n487) );
  XNOR2_X1 U442 ( .A(n485), .B(n486), .ZN(n467) );
  XNOR2_X1 U443 ( .A(n544), .B(n447), .ZN(n446) );
  XNOR2_X1 U444 ( .A(n515), .B(KEYINPUT77), .ZN(n516) );
  INV_X1 U445 ( .A(G128), .ZN(n470) );
  XNOR2_X1 U446 ( .A(G143), .B(G131), .ZN(n534) );
  INV_X1 U447 ( .A(KEYINPUT98), .ZN(n408) );
  XNOR2_X1 U448 ( .A(G113), .B(G104), .ZN(n526) );
  XOR2_X1 U449 ( .A(G140), .B(G122), .Z(n527) );
  XOR2_X1 U450 ( .A(KEYINPUT11), .B(KEYINPUT12), .Z(n532) );
  INV_X1 U451 ( .A(KEYINPUT75), .ZN(n461) );
  XNOR2_X1 U452 ( .A(n459), .B(G140), .ZN(n497) );
  INV_X1 U453 ( .A(G137), .ZN(n459) );
  XNOR2_X1 U454 ( .A(n432), .B(n431), .ZN(n511) );
  XNOR2_X1 U455 ( .A(KEYINPUT89), .B(G110), .ZN(n431) );
  XNOR2_X1 U456 ( .A(n433), .B(G107), .ZN(n432) );
  INV_X1 U457 ( .A(G104), .ZN(n433) );
  XNOR2_X1 U458 ( .A(KEYINPUT4), .B(KEYINPUT91), .ZN(n504) );
  XOR2_X1 U459 ( .A(KEYINPUT18), .B(KEYINPUT17), .Z(n505) );
  XOR2_X1 U460 ( .A(G146), .B(G125), .Z(n508) );
  XOR2_X1 U461 ( .A(G101), .B(KEYINPUT69), .Z(n509) );
  AND2_X1 U462 ( .A1(n672), .A2(n618), .ZN(n442) );
  INV_X1 U463 ( .A(n670), .ZN(n618) );
  XNOR2_X1 U464 ( .A(KEYINPUT38), .B(n622), .ZN(n683) );
  AND2_X1 U465 ( .A1(n590), .A2(n436), .ZN(n608) );
  XNOR2_X1 U466 ( .A(n589), .B(KEYINPUT109), .ZN(n590) );
  NAND2_X2 U467 ( .A1(n394), .A2(n391), .ZN(n420) );
  AND2_X1 U468 ( .A1(n396), .A2(n395), .ZN(n394) );
  NAND2_X1 U469 ( .A1(G469), .A2(G902), .ZN(n395) );
  AND2_X1 U470 ( .A1(n564), .A2(n468), .ZN(n696) );
  INV_X1 U471 ( .A(n693), .ZN(n468) );
  XNOR2_X1 U472 ( .A(n437), .B(n512), .ZN(n482) );
  XNOR2_X1 U473 ( .A(n469), .B(n481), .ZN(n437) );
  XNOR2_X1 U474 ( .A(n457), .B(n512), .ZN(n737) );
  XNOR2_X1 U475 ( .A(n511), .B(n513), .ZN(n457) );
  XOR2_X1 U476 ( .A(G122), .B(KEYINPUT16), .Z(n513) );
  XNOR2_X1 U477 ( .A(n439), .B(KEYINPUT24), .ZN(n485) );
  XNOR2_X1 U478 ( .A(G110), .B(KEYINPUT23), .ZN(n439) );
  XNOR2_X1 U479 ( .A(G128), .B(G119), .ZN(n486) );
  XNOR2_X1 U480 ( .A(n484), .B(n466), .ZN(n543) );
  INV_X1 U481 ( .A(KEYINPUT8), .ZN(n466) );
  XNOR2_X1 U482 ( .A(n540), .B(n542), .ZN(n447) );
  NAND2_X1 U483 ( .A1(n448), .A2(n661), .ZN(n619) );
  NOR2_X1 U484 ( .A1(n450), .A2(n449), .ZN(n448) );
  NAND2_X1 U485 ( .A1(n694), .A2(n368), .ZN(n449) );
  INV_X1 U486 ( .A(n591), .ZN(n440) );
  XNOR2_X1 U487 ( .A(n388), .B(n387), .ZN(n451) );
  INV_X1 U488 ( .A(n523), .ZN(n387) );
  OR2_X1 U489 ( .A1(n753), .A2(n571), .ZN(n572) );
  AND2_X1 U490 ( .A1(n386), .A2(n379), .ZN(n412) );
  NAND2_X1 U491 ( .A1(n381), .A2(n369), .ZN(n386) );
  XNOR2_X1 U492 ( .A(n547), .B(KEYINPUT103), .ZN(n651) );
  XNOR2_X1 U493 ( .A(n388), .B(n365), .ZN(n551) );
  XNOR2_X1 U494 ( .A(n640), .B(n639), .ZN(n641) );
  XNOR2_X1 U495 ( .A(n607), .B(n404), .ZN(n760) );
  XNOR2_X1 U496 ( .A(KEYINPUT42), .B(KEYINPUT114), .ZN(n404) );
  XNOR2_X1 U497 ( .A(n613), .B(KEYINPUT40), .ZN(n764) );
  NAND2_X1 U498 ( .A1(n425), .A2(n424), .ZN(n562) );
  AND2_X1 U499 ( .A1(n561), .A2(n450), .ZN(n424) );
  NOR2_X1 U500 ( .A1(n697), .A2(n356), .ZN(n438) );
  XNOR2_X1 U501 ( .A(n612), .B(KEYINPUT107), .ZN(n661) );
  AND2_X1 U502 ( .A1(n551), .A2(n397), .ZN(n652) );
  NOR2_X1 U503 ( .A1(n356), .A2(n589), .ZN(n397) );
  XNOR2_X1 U504 ( .A(n734), .B(n735), .ZN(n400) );
  XNOR2_X1 U505 ( .A(n731), .B(n732), .ZN(n401) );
  XNOR2_X1 U506 ( .A(n729), .B(n730), .ZN(n399) );
  INV_X1 U507 ( .A(KEYINPUT56), .ZN(n402) );
  NAND2_X1 U508 ( .A1(G214), .A2(n517), .ZN(n682) );
  XNOR2_X1 U509 ( .A(n549), .B(n429), .ZN(n554) );
  AND2_X1 U510 ( .A1(n454), .A2(n566), .ZN(n358) );
  XNOR2_X1 U511 ( .A(KEYINPUT19), .B(KEYINPUT67), .ZN(n359) );
  OR2_X1 U512 ( .A1(n416), .A2(n626), .ZN(n360) );
  XOR2_X1 U513 ( .A(n539), .B(n541), .Z(n361) );
  XOR2_X1 U514 ( .A(n509), .B(n508), .Z(n362) );
  AND2_X1 U515 ( .A1(G224), .A2(n753), .ZN(n363) );
  OR2_X1 U516 ( .A1(n574), .A2(n521), .ZN(n364) );
  XOR2_X1 U517 ( .A(n523), .B(KEYINPUT94), .Z(n365) );
  AND2_X1 U518 ( .A1(n556), .A2(n440), .ZN(n366) );
  AND2_X1 U519 ( .A1(n586), .A2(n585), .ZN(n367) );
  INV_X1 U520 ( .A(n435), .ZN(n450) );
  AND2_X1 U521 ( .A1(n598), .A2(n682), .ZN(n368) );
  BUF_X1 U522 ( .A(n560), .Z(n697) );
  AND2_X1 U523 ( .A1(n380), .A2(n359), .ZN(n369) );
  INV_X1 U524 ( .A(G469), .ZN(n502) );
  XNOR2_X1 U525 ( .A(KEYINPUT71), .B(KEYINPUT34), .ZN(n370) );
  XOR2_X1 U526 ( .A(n635), .B(KEYINPUT62), .Z(n371) );
  XNOR2_X1 U527 ( .A(n723), .B(n722), .ZN(n372) );
  INV_X1 U528 ( .A(n736), .ZN(n643) );
  XOR2_X1 U529 ( .A(n638), .B(n637), .Z(n373) );
  NAND2_X1 U530 ( .A1(n377), .A2(n686), .ZN(n376) );
  XNOR2_X1 U531 ( .A(n524), .B(KEYINPUT97), .ZN(n377) );
  NAND2_X1 U532 ( .A1(n378), .A2(n383), .ZN(n379) );
  NAND2_X1 U533 ( .A1(n721), .A2(n416), .ZN(n382) );
  INV_X1 U534 ( .A(n415), .ZN(n385) );
  NAND2_X2 U535 ( .A1(n389), .A2(n364), .ZN(n388) );
  INV_X1 U536 ( .A(n579), .ZN(n389) );
  AND2_X1 U537 ( .A1(n358), .A2(n390), .ZN(n453) );
  NAND2_X1 U538 ( .A1(n390), .A2(n454), .ZN(n419) );
  XNOR2_X1 U539 ( .A(n390), .B(G122), .ZN(G24) );
  XNOR2_X2 U540 ( .A(n553), .B(n552), .ZN(n390) );
  NAND2_X1 U541 ( .A1(n725), .A2(G469), .ZN(n396) );
  XNOR2_X2 U542 ( .A(n501), .B(n500), .ZN(n725) );
  OR2_X1 U543 ( .A1(n725), .A2(n392), .ZN(n391) );
  NOR2_X1 U544 ( .A1(n399), .A2(n736), .ZN(G54) );
  NOR2_X1 U545 ( .A1(n400), .A2(n736), .ZN(G66) );
  NOR2_X1 U546 ( .A1(n401), .A2(n736), .ZN(G63) );
  NAND2_X1 U547 ( .A1(n412), .A2(n409), .ZN(n579) );
  XNOR2_X1 U548 ( .A(n403), .B(n402), .ZN(G51) );
  NAND2_X1 U549 ( .A1(n428), .A2(n643), .ZN(n403) );
  NOR2_X1 U550 ( .A1(n563), .A2(n564), .ZN(n565) );
  NAND2_X1 U551 ( .A1(n414), .A2(n413), .ZN(n622) );
  INV_X1 U552 ( .A(n550), .ZN(n434) );
  NAND2_X1 U553 ( .A1(n463), .A2(n464), .ZN(n444) );
  XNOR2_X1 U554 ( .A(n446), .B(n445), .ZN(n732) );
  NOR2_X2 U555 ( .A1(n665), .A2(n652), .ZN(n524) );
  XNOR2_X2 U556 ( .A(n522), .B(KEYINPUT31), .ZN(n665) );
  NAND2_X1 U557 ( .A1(n565), .A2(n438), .ZN(n454) );
  NAND2_X1 U558 ( .A1(n414), .A2(n410), .ZN(n409) );
  AND2_X1 U559 ( .A1(n413), .A2(n411), .ZN(n410) );
  INV_X1 U560 ( .A(n516), .ZN(n416) );
  INV_X1 U561 ( .A(n682), .ZN(n417) );
  XNOR2_X2 U562 ( .A(n418), .B(n475), .ZN(n749) );
  XNOR2_X1 U563 ( .A(n418), .B(n361), .ZN(n445) );
  XNOR2_X2 U564 ( .A(n503), .B(G134), .ZN(n418) );
  NAND2_X1 U565 ( .A1(n419), .A2(KEYINPUT44), .ZN(n452) );
  NAND2_X1 U566 ( .A1(n696), .A2(n420), .ZN(n589) );
  NAND2_X1 U567 ( .A1(n577), .A2(n420), .ZN(n578) );
  NAND2_X1 U568 ( .A1(n453), .A2(n763), .ZN(n421) );
  NOR2_X1 U569 ( .A1(n563), .A2(n435), .ZN(n426) );
  INV_X1 U570 ( .A(n563), .ZN(n425) );
  NAND2_X1 U571 ( .A1(n426), .A2(n567), .ZN(n568) );
  XNOR2_X1 U572 ( .A(n427), .B(n373), .ZN(G57) );
  NAND2_X1 U573 ( .A1(n430), .A2(n643), .ZN(n427) );
  XNOR2_X1 U574 ( .A(n724), .B(n372), .ZN(n428) );
  XNOR2_X2 U575 ( .A(n483), .B(G472), .ZN(n549) );
  XNOR2_X1 U576 ( .A(n636), .B(n371), .ZN(n430) );
  NAND2_X1 U577 ( .A1(n543), .A2(G221), .ZN(n465) );
  INV_X1 U578 ( .A(n554), .ZN(n435) );
  XNOR2_X1 U579 ( .A(n458), .B(n370), .ZN(n441) );
  NAND2_X1 U580 ( .A1(n441), .A2(n366), .ZN(n553) );
  XNOR2_X1 U581 ( .A(n615), .B(n614), .ZN(n463) );
  XNOR2_X1 U582 ( .A(n588), .B(n587), .ZN(n436) );
  XNOR2_X1 U583 ( .A(n444), .B(n462), .ZN(n443) );
  NOR2_X1 U584 ( .A1(G902), .A2(n735), .ZN(n493) );
  NOR2_X2 U585 ( .A1(n606), .A2(n580), .ZN(n659) );
  INV_X1 U586 ( .A(n454), .ZN(n655) );
  NAND2_X1 U587 ( .A1(n443), .A2(n442), .ZN(n630) );
  NOR2_X2 U588 ( .A1(G902), .A2(n635), .ZN(n483) );
  NAND2_X1 U589 ( .A1(n451), .A2(n557), .ZN(n558) );
  NAND2_X1 U590 ( .A1(n451), .A2(n704), .ZN(n522) );
  NAND2_X1 U591 ( .A1(n681), .A2(n551), .ZN(n458) );
  NAND2_X1 U592 ( .A1(n644), .A2(n643), .ZN(n646) );
  XNOR2_X1 U593 ( .A(n642), .B(n641), .ZN(n644) );
  NOR2_X1 U594 ( .A1(G952), .A2(n753), .ZN(n736) );
  XOR2_X1 U595 ( .A(n480), .B(KEYINPUT96), .Z(n469) );
  INV_X1 U596 ( .A(KEYINPUT44), .ZN(n566) );
  XNOR2_X1 U597 ( .A(n474), .B(G131), .ZN(n475) );
  XNOR2_X1 U598 ( .A(n509), .B(G146), .ZN(n476) );
  XNOR2_X1 U599 ( .A(n510), .B(n362), .ZN(n514) );
  XNOR2_X1 U600 ( .A(n603), .B(KEYINPUT41), .ZN(n604) );
  XNOR2_X1 U601 ( .A(n511), .B(n499), .ZN(n500) );
  INV_X1 U602 ( .A(KEYINPUT60), .ZN(n645) );
  NAND2_X1 U603 ( .A1(G143), .A2(n470), .ZN(n473) );
  NAND2_X1 U604 ( .A1(n471), .A2(G128), .ZN(n472) );
  XNOR2_X2 U605 ( .A(n749), .B(n476), .ZN(n501) );
  NAND2_X1 U606 ( .A1(n530), .A2(G210), .ZN(n481) );
  XNOR2_X1 U607 ( .A(n508), .B(KEYINPUT10), .ZN(n525) );
  XNOR2_X1 U608 ( .A(n497), .B(n525), .ZN(n750) );
  NAND2_X1 U609 ( .A1(G234), .A2(n753), .ZN(n484) );
  XNOR2_X1 U610 ( .A(n750), .B(n487), .ZN(n735) );
  INV_X1 U611 ( .A(n626), .ZN(n488) );
  NAND2_X1 U612 ( .A1(n488), .A2(G234), .ZN(n489) );
  XNOR2_X1 U613 ( .A(n489), .B(KEYINPUT20), .ZN(n494) );
  NAND2_X1 U614 ( .A1(G217), .A2(n494), .ZN(n491) );
  XNOR2_X1 U615 ( .A(KEYINPUT25), .B(KEYINPUT74), .ZN(n490) );
  XOR2_X1 U616 ( .A(KEYINPUT95), .B(KEYINPUT21), .Z(n496) );
  NAND2_X1 U617 ( .A1(n494), .A2(G221), .ZN(n495) );
  XNOR2_X1 U618 ( .A(n496), .B(n495), .ZN(n693) );
  NAND2_X1 U619 ( .A1(G227), .A2(n753), .ZN(n498) );
  NAND2_X1 U620 ( .A1(n696), .A2(n560), .ZN(n550) );
  NOR2_X1 U621 ( .A1(n549), .A2(n550), .ZN(n704) );
  XNOR2_X1 U622 ( .A(n357), .B(n363), .ZN(n507) );
  XNOR2_X1 U623 ( .A(n505), .B(n504), .ZN(n506) );
  XNOR2_X1 U624 ( .A(n507), .B(n506), .ZN(n510) );
  NAND2_X1 U625 ( .A1(G210), .A2(n517), .ZN(n515) );
  XNOR2_X1 U626 ( .A(n518), .B(KEYINPUT92), .ZN(n519) );
  XNOR2_X1 U627 ( .A(KEYINPUT14), .B(n519), .ZN(n520) );
  NAND2_X1 U628 ( .A1(G952), .A2(n520), .ZN(n712) );
  NOR2_X1 U629 ( .A1(G953), .A2(n712), .ZN(n574) );
  NAND2_X1 U630 ( .A1(n520), .A2(G902), .ZN(n571) );
  XNOR2_X1 U631 ( .A(G898), .B(KEYINPUT93), .ZN(n743) );
  NAND2_X1 U632 ( .A1(G953), .A2(n743), .ZN(n739) );
  NOR2_X1 U633 ( .A1(n571), .A2(n739), .ZN(n521) );
  XNOR2_X1 U634 ( .A(KEYINPUT68), .B(KEYINPUT0), .ZN(n523) );
  XNOR2_X1 U635 ( .A(KEYINPUT13), .B(G475), .ZN(n538) );
  INV_X1 U636 ( .A(n525), .ZN(n529) );
  XNOR2_X1 U637 ( .A(n527), .B(n526), .ZN(n528) );
  XNOR2_X1 U638 ( .A(n529), .B(n528), .ZN(n536) );
  NAND2_X1 U639 ( .A1(G214), .A2(n530), .ZN(n531) );
  XNOR2_X1 U640 ( .A(n532), .B(n531), .ZN(n533) );
  XNOR2_X1 U641 ( .A(n536), .B(n535), .ZN(n640) );
  NOR2_X1 U642 ( .A1(G902), .A2(n640), .ZN(n537) );
  XOR2_X1 U643 ( .A(KEYINPUT9), .B(G122), .Z(n540) );
  XNOR2_X1 U644 ( .A(G116), .B(G107), .ZN(n539) );
  XOR2_X1 U645 ( .A(KEYINPUT100), .B(KEYINPUT99), .Z(n542) );
  XNOR2_X1 U646 ( .A(KEYINPUT7), .B(KEYINPUT101), .ZN(n541) );
  NAND2_X1 U647 ( .A1(G217), .A2(n543), .ZN(n544) );
  NOR2_X1 U648 ( .A1(n732), .A2(G902), .ZN(n545) );
  XNOR2_X1 U649 ( .A(n545), .B(G478), .ZN(n546) );
  NAND2_X1 U650 ( .A1(n556), .A2(n591), .ZN(n612) );
  NOR2_X1 U651 ( .A1(n591), .A2(n556), .ZN(n547) );
  NAND2_X1 U652 ( .A1(n612), .A2(n651), .ZN(n548) );
  XNOR2_X1 U653 ( .A(KEYINPUT104), .B(n548), .ZN(n686) );
  XOR2_X1 U654 ( .A(KEYINPUT76), .B(KEYINPUT35), .Z(n552) );
  XNOR2_X1 U655 ( .A(KEYINPUT22), .B(KEYINPUT72), .ZN(n555) );
  XNOR2_X1 U656 ( .A(n555), .B(KEYINPUT66), .ZN(n559) );
  INV_X1 U657 ( .A(n556), .ZN(n594) );
  NAND2_X1 U658 ( .A1(n591), .A2(n594), .ZN(n685) );
  NOR2_X1 U659 ( .A1(n685), .A2(n693), .ZN(n557) );
  AND2_X1 U660 ( .A1(n697), .A2(n694), .ZN(n561) );
  NOR2_X1 U661 ( .A1(n697), .A2(n694), .ZN(n567) );
  XOR2_X1 U662 ( .A(KEYINPUT85), .B(KEYINPUT45), .Z(n569) );
  NAND2_X1 U663 ( .A1(n629), .A2(n626), .ZN(n570) );
  XNOR2_X1 U664 ( .A(n570), .B(KEYINPUT83), .ZN(n624) );
  NOR2_X1 U665 ( .A1(G900), .A2(n572), .ZN(n573) );
  NOR2_X1 U666 ( .A1(n574), .A2(n573), .ZN(n609) );
  NOR2_X1 U667 ( .A1(n693), .A2(n609), .ZN(n598) );
  NAND2_X1 U668 ( .A1(n598), .A2(n694), .ZN(n575) );
  NOR2_X1 U669 ( .A1(n549), .A2(n575), .ZN(n576) );
  XNOR2_X1 U670 ( .A(KEYINPUT28), .B(n576), .ZN(n577) );
  XNOR2_X1 U671 ( .A(n578), .B(KEYINPUT112), .ZN(n606) );
  BUF_X1 U672 ( .A(n579), .Z(n580) );
  XNOR2_X1 U673 ( .A(n581), .B(KEYINPUT47), .ZN(n583) );
  INV_X1 U674 ( .A(KEYINPUT79), .ZN(n582) );
  NAND2_X1 U675 ( .A1(n583), .A2(n582), .ZN(n586) );
  NAND2_X1 U676 ( .A1(KEYINPUT47), .A2(n686), .ZN(n584) );
  NAND2_X1 U677 ( .A1(n584), .A2(KEYINPUT79), .ZN(n585) );
  NAND2_X1 U678 ( .A1(n356), .A2(n682), .ZN(n588) );
  XOR2_X1 U679 ( .A(KEYINPUT30), .B(KEYINPUT110), .Z(n587) );
  INV_X1 U680 ( .A(n608), .ZN(n593) );
  OR2_X1 U681 ( .A1(n622), .A2(n591), .ZN(n592) );
  NOR2_X1 U682 ( .A1(n593), .A2(n592), .ZN(n596) );
  NOR2_X1 U683 ( .A1(n594), .A2(n609), .ZN(n595) );
  NAND2_X1 U684 ( .A1(n596), .A2(n595), .ZN(n597) );
  XNOR2_X1 U685 ( .A(KEYINPUT111), .B(n597), .ZN(n762) );
  NAND2_X1 U686 ( .A1(n659), .A2(KEYINPUT79), .ZN(n601) );
  NOR2_X1 U687 ( .A1(n622), .A2(n619), .ZN(n599) );
  XNOR2_X1 U688 ( .A(n599), .B(KEYINPUT36), .ZN(n600) );
  NAND2_X1 U689 ( .A1(n600), .A2(n697), .ZN(n669) );
  NAND2_X1 U690 ( .A1(n601), .A2(n669), .ZN(n602) );
  NOR2_X1 U691 ( .A1(n762), .A2(n602), .ZN(n616) );
  NAND2_X1 U692 ( .A1(n683), .A2(n682), .ZN(n687) );
  XNOR2_X1 U693 ( .A(n605), .B(n604), .ZN(n713) );
  NOR2_X1 U694 ( .A1(n606), .A2(n713), .ZN(n607) );
  NAND2_X1 U695 ( .A1(n608), .A2(n683), .ZN(n610) );
  XNOR2_X1 U696 ( .A(n611), .B(KEYINPUT39), .ZN(n617) );
  NOR2_X1 U697 ( .A1(n617), .A2(n612), .ZN(n613) );
  XNOR2_X1 U698 ( .A(KEYINPUT64), .B(KEYINPUT46), .ZN(n614) );
  NOR2_X1 U699 ( .A1(n617), .A2(n651), .ZN(n670) );
  OR2_X1 U700 ( .A1(n619), .A2(n697), .ZN(n621) );
  XNOR2_X1 U701 ( .A(KEYINPUT108), .B(KEYINPUT43), .ZN(n620) );
  XNOR2_X1 U702 ( .A(n621), .B(n620), .ZN(n623) );
  NAND2_X1 U703 ( .A1(n623), .A2(n622), .ZN(n672) );
  NAND2_X1 U704 ( .A1(n624), .A2(n751), .ZN(n625) );
  XNOR2_X1 U705 ( .A(n625), .B(KEYINPUT82), .ZN(n628) );
  NAND2_X1 U706 ( .A1(KEYINPUT2), .A2(n626), .ZN(n627) );
  NAND2_X1 U707 ( .A1(n628), .A2(n627), .ZN(n633) );
  NAND2_X1 U708 ( .A1(n744), .A2(KEYINPUT2), .ZN(n631) );
  XNOR2_X1 U709 ( .A(n632), .B(KEYINPUT73), .ZN(n679) );
  NAND2_X1 U710 ( .A1(n633), .A2(n679), .ZN(n634) );
  XNOR2_X2 U711 ( .A(n634), .B(KEYINPUT65), .ZN(n728) );
  NAND2_X1 U712 ( .A1(n728), .A2(G472), .ZN(n636) );
  XNOR2_X1 U713 ( .A(KEYINPUT86), .B(KEYINPUT88), .ZN(n638) );
  INV_X1 U714 ( .A(KEYINPUT63), .ZN(n637) );
  NAND2_X1 U715 ( .A1(n728), .A2(G475), .ZN(n642) );
  XOR2_X1 U716 ( .A(KEYINPUT59), .B(KEYINPUT125), .Z(n639) );
  XNOR2_X1 U717 ( .A(n646), .B(n645), .ZN(G60) );
  NAND2_X1 U718 ( .A1(n652), .A2(n661), .ZN(n647) );
  XNOR2_X1 U719 ( .A(n647), .B(G104), .ZN(G6) );
  XOR2_X1 U720 ( .A(KEYINPUT27), .B(KEYINPUT116), .Z(n649) );
  XNOR2_X1 U721 ( .A(G107), .B(KEYINPUT26), .ZN(n648) );
  XNOR2_X1 U722 ( .A(n649), .B(n648), .ZN(n650) );
  XOR2_X1 U723 ( .A(KEYINPUT115), .B(n650), .Z(n654) );
  INV_X1 U724 ( .A(n651), .ZN(n664) );
  NAND2_X1 U725 ( .A1(n652), .A2(n664), .ZN(n653) );
  XNOR2_X1 U726 ( .A(n654), .B(n653), .ZN(G9) );
  XOR2_X1 U727 ( .A(G110), .B(n655), .Z(G12) );
  XOR2_X1 U728 ( .A(KEYINPUT117), .B(KEYINPUT29), .Z(n657) );
  NAND2_X1 U729 ( .A1(n659), .A2(n664), .ZN(n656) );
  XNOR2_X1 U730 ( .A(n657), .B(n656), .ZN(n658) );
  XOR2_X1 U731 ( .A(G128), .B(n658), .Z(G30) );
  NAND2_X1 U732 ( .A1(n659), .A2(n661), .ZN(n660) );
  XNOR2_X1 U733 ( .A(n660), .B(G146), .ZN(G48) );
  NAND2_X1 U734 ( .A1(n665), .A2(n661), .ZN(n662) );
  XNOR2_X1 U735 ( .A(n662), .B(KEYINPUT118), .ZN(n663) );
  XNOR2_X1 U736 ( .A(G113), .B(n663), .ZN(G15) );
  XOR2_X1 U737 ( .A(G116), .B(KEYINPUT119), .Z(n667) );
  NAND2_X1 U738 ( .A1(n665), .A2(n664), .ZN(n666) );
  XNOR2_X1 U739 ( .A(n667), .B(n666), .ZN(G18) );
  XOR2_X1 U740 ( .A(G125), .B(KEYINPUT37), .Z(n668) );
  XNOR2_X1 U741 ( .A(n669), .B(n668), .ZN(G27) );
  XOR2_X1 U742 ( .A(G134), .B(n670), .Z(n671) );
  XNOR2_X1 U743 ( .A(KEYINPUT120), .B(n671), .ZN(G36) );
  XNOR2_X1 U744 ( .A(G140), .B(n672), .ZN(G42) );
  XNOR2_X1 U745 ( .A(KEYINPUT2), .B(KEYINPUT78), .ZN(n674) );
  OR2_X1 U746 ( .A1(n751), .A2(n674), .ZN(n673) );
  XNOR2_X1 U747 ( .A(n673), .B(KEYINPUT81), .ZN(n677) );
  NOR2_X1 U748 ( .A1(n744), .A2(n674), .ZN(n675) );
  XNOR2_X1 U749 ( .A(n675), .B(KEYINPUT80), .ZN(n676) );
  NOR2_X1 U750 ( .A1(n677), .A2(n676), .ZN(n678) );
  NAND2_X1 U751 ( .A1(n679), .A2(n678), .ZN(n680) );
  XNOR2_X1 U752 ( .A(n680), .B(KEYINPUT84), .ZN(n718) );
  INV_X1 U753 ( .A(n681), .ZN(n714) );
  NOR2_X1 U754 ( .A1(n683), .A2(n682), .ZN(n684) );
  NOR2_X1 U755 ( .A1(n685), .A2(n684), .ZN(n690) );
  INV_X1 U756 ( .A(n686), .ZN(n688) );
  NOR2_X1 U757 ( .A1(n688), .A2(n687), .ZN(n689) );
  NOR2_X1 U758 ( .A1(n690), .A2(n689), .ZN(n691) );
  XOR2_X1 U759 ( .A(KEYINPUT123), .B(n691), .Z(n692) );
  NOR2_X1 U760 ( .A1(n714), .A2(n692), .ZN(n709) );
  AND2_X1 U761 ( .A1(n694), .A2(n693), .ZN(n695) );
  XNOR2_X1 U762 ( .A(KEYINPUT49), .B(n695), .ZN(n701) );
  XOR2_X1 U763 ( .A(KEYINPUT121), .B(KEYINPUT50), .Z(n699) );
  OR2_X1 U764 ( .A1(n697), .A2(n696), .ZN(n698) );
  XNOR2_X1 U765 ( .A(n699), .B(n698), .ZN(n700) );
  NAND2_X1 U766 ( .A1(n701), .A2(n700), .ZN(n702) );
  NOR2_X1 U767 ( .A1(n356), .A2(n702), .ZN(n703) );
  NOR2_X1 U768 ( .A1(n704), .A2(n703), .ZN(n705) );
  XOR2_X1 U769 ( .A(n705), .B(KEYINPUT122), .Z(n706) );
  XNOR2_X1 U770 ( .A(KEYINPUT51), .B(n706), .ZN(n707) );
  NOR2_X1 U771 ( .A1(n713), .A2(n707), .ZN(n708) );
  NOR2_X1 U772 ( .A1(n709), .A2(n708), .ZN(n710) );
  XNOR2_X1 U773 ( .A(n710), .B(KEYINPUT52), .ZN(n711) );
  NOR2_X1 U774 ( .A1(n712), .A2(n711), .ZN(n716) );
  NOR2_X1 U775 ( .A1(n714), .A2(n713), .ZN(n715) );
  NOR2_X1 U776 ( .A1(n716), .A2(n715), .ZN(n717) );
  NAND2_X1 U777 ( .A1(n718), .A2(n717), .ZN(n719) );
  NOR2_X1 U778 ( .A1(n719), .A2(G953), .ZN(n720) );
  XNOR2_X1 U779 ( .A(n720), .B(KEYINPUT53), .ZN(G75) );
  NAND2_X1 U780 ( .A1(n728), .A2(G210), .ZN(n724) );
  XOR2_X1 U781 ( .A(KEYINPUT54), .B(KEYINPUT55), .Z(n723) );
  XNOR2_X1 U782 ( .A(n721), .B(KEYINPUT87), .ZN(n722) );
  XOR2_X1 U783 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n727) );
  XNOR2_X1 U784 ( .A(n725), .B(KEYINPUT124), .ZN(n726) );
  XNOR2_X1 U785 ( .A(n727), .B(n726), .ZN(n730) );
  NAND2_X1 U786 ( .A1(n733), .A2(G469), .ZN(n729) );
  NAND2_X1 U787 ( .A1(G478), .A2(n733), .ZN(n731) );
  NAND2_X1 U788 ( .A1(n733), .A2(G217), .ZN(n734) );
  XOR2_X1 U789 ( .A(n737), .B(G101), .Z(n738) );
  XNOR2_X1 U790 ( .A(KEYINPUT126), .B(n738), .ZN(n740) );
  NAND2_X1 U791 ( .A1(n740), .A2(n739), .ZN(n748) );
  NAND2_X1 U792 ( .A1(G953), .A2(G224), .ZN(n741) );
  XOR2_X1 U793 ( .A(KEYINPUT61), .B(n741), .Z(n742) );
  NOR2_X1 U794 ( .A1(n743), .A2(n742), .ZN(n746) );
  AND2_X1 U795 ( .A1(n744), .A2(n753), .ZN(n745) );
  NOR2_X1 U796 ( .A1(n746), .A2(n745), .ZN(n747) );
  XNOR2_X1 U797 ( .A(n748), .B(n747), .ZN(G69) );
  XOR2_X1 U798 ( .A(n749), .B(n750), .Z(n755) );
  INV_X1 U799 ( .A(n755), .ZN(n752) );
  XNOR2_X1 U800 ( .A(n752), .B(n751), .ZN(n754) );
  NAND2_X1 U801 ( .A1(n754), .A2(n753), .ZN(n759) );
  XNOR2_X1 U802 ( .A(G227), .B(n755), .ZN(n756) );
  NAND2_X1 U803 ( .A1(n756), .A2(G900), .ZN(n757) );
  NAND2_X1 U804 ( .A1(n757), .A2(G953), .ZN(n758) );
  NAND2_X1 U805 ( .A1(n759), .A2(n758), .ZN(G72) );
  XNOR2_X1 U806 ( .A(n760), .B(G137), .ZN(n761) );
  XNOR2_X1 U807 ( .A(n761), .B(KEYINPUT127), .ZN(G39) );
  XOR2_X1 U808 ( .A(G143), .B(n762), .Z(G45) );
  XNOR2_X1 U809 ( .A(n763), .B(G119), .ZN(G21) );
  XOR2_X1 U810 ( .A(n764), .B(G131), .Z(G33) );
  XNOR2_X1 U811 ( .A(G101), .B(n765), .ZN(G3) );
endmodule

