//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 1 1 1 1 1 0 0 1 1 1 0 1 1 0 0 1 1 0 0 1 0 0 0 1 1 1 0 0 1 0 0 0 0 0 1 0 0 0 1 0 1 0 0 0 0 0 1 1 0 1 0 1 0 0 0 0 0 0 0 1 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:37:14 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n205, new_n206, new_n207, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n241, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n251, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1108, new_n1109, new_n1110, new_n1111, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1249, new_n1250, new_n1251, new_n1252, new_n1253,
    new_n1254, new_n1255, new_n1256, new_n1257, new_n1258, new_n1259,
    new_n1260, new_n1261, new_n1262, new_n1263, new_n1264, new_n1265,
    new_n1266, new_n1267, new_n1268, new_n1269, new_n1270, new_n1271,
    new_n1272, new_n1274, new_n1275, new_n1276, new_n1277, new_n1278,
    new_n1280, new_n1281, new_n1282, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1346,
    new_n1347, new_n1348, new_n1349, new_n1351, new_n1352, new_n1353,
    new_n1354, new_n1355, new_n1356, new_n1357, new_n1358, new_n1359,
    new_n1360;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  INV_X1    g0004(.A(G97), .ZN(new_n205));
  INV_X1    g0005(.A(G107), .ZN(new_n206));
  NAND2_X1  g0006(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  NAND2_X1  g0007(.A1(new_n207), .A2(G87), .ZN(G355));
  INV_X1    g0008(.A(G1), .ZN(new_n209));
  INV_X1    g0009(.A(G20), .ZN(new_n210));
  NOR2_X1   g0010(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  INV_X1    g0011(.A(new_n211), .ZN(new_n212));
  NOR2_X1   g0012(.A1(new_n212), .A2(G13), .ZN(new_n213));
  OAI211_X1 g0013(.A(new_n213), .B(G250), .C1(G257), .C2(G264), .ZN(new_n214));
  XOR2_X1   g0014(.A(new_n214), .B(KEYINPUT64), .Z(new_n215));
  XNOR2_X1  g0015(.A(new_n215), .B(KEYINPUT0), .ZN(new_n216));
  AOI22_X1  g0016(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n217));
  XNOR2_X1  g0017(.A(new_n217), .B(KEYINPUT65), .ZN(new_n218));
  AOI22_X1  g0018(.A1(G58), .A2(G232), .B1(G116), .B2(G270), .ZN(new_n219));
  AOI22_X1  g0019(.A1(G50), .A2(G226), .B1(G68), .B2(G238), .ZN(new_n220));
  AOI22_X1  g0020(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n221));
  NAND3_X1  g0021(.A1(new_n219), .A2(new_n220), .A3(new_n221), .ZN(new_n222));
  OAI21_X1  g0022(.A(new_n212), .B1(new_n218), .B2(new_n222), .ZN(new_n223));
  XOR2_X1   g0023(.A(new_n223), .B(KEYINPUT66), .Z(new_n224));
  INV_X1    g0024(.A(KEYINPUT1), .ZN(new_n225));
  AND2_X1   g0025(.A1(new_n224), .A2(new_n225), .ZN(new_n226));
  NOR2_X1   g0026(.A1(new_n224), .A2(new_n225), .ZN(new_n227));
  INV_X1    g0027(.A(new_n201), .ZN(new_n228));
  NAND2_X1  g0028(.A1(new_n228), .A2(G50), .ZN(new_n229));
  NAND2_X1  g0029(.A1(G1), .A2(G13), .ZN(new_n230));
  NOR3_X1   g0030(.A1(new_n229), .A2(new_n210), .A3(new_n230), .ZN(new_n231));
  NOR4_X1   g0031(.A1(new_n216), .A2(new_n226), .A3(new_n227), .A4(new_n231), .ZN(G361));
  XNOR2_X1  g0032(.A(G238), .B(G244), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n233), .B(G232), .ZN(new_n234));
  XNOR2_X1  g0034(.A(KEYINPUT2), .B(G226), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XOR2_X1   g0036(.A(G264), .B(G270), .Z(new_n237));
  XNOR2_X1  g0037(.A(G250), .B(G257), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n236), .B(new_n239), .ZN(G358));
  XNOR2_X1  g0040(.A(G87), .B(G97), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n241), .B(KEYINPUT67), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n242), .B(KEYINPUT68), .ZN(new_n243));
  XOR2_X1   g0043(.A(G107), .B(G116), .Z(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  NAND2_X1  g0045(.A1(new_n202), .A2(G68), .ZN(new_n246));
  INV_X1    g0046(.A(G68), .ZN(new_n247));
  NAND2_X1  g0047(.A1(new_n247), .A2(G50), .ZN(new_n248));
  NAND2_X1  g0048(.A1(new_n246), .A2(new_n248), .ZN(new_n249));
  XNOR2_X1  g0049(.A(G58), .B(G77), .ZN(new_n250));
  XNOR2_X1  g0050(.A(new_n249), .B(new_n250), .ZN(new_n251));
  XNOR2_X1  g0051(.A(new_n245), .B(new_n251), .ZN(G351));
  INV_X1    g0052(.A(G169), .ZN(new_n253));
  NAND3_X1  g0053(.A1(new_n209), .A2(G13), .A3(G20), .ZN(new_n254));
  NOR2_X1   g0054(.A1(new_n254), .A2(G116), .ZN(new_n255));
  INV_X1    g0055(.A(new_n254), .ZN(new_n256));
  NAND3_X1  g0056(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n257));
  NAND2_X1  g0057(.A1(new_n257), .A2(new_n230), .ZN(new_n258));
  NOR2_X1   g0058(.A1(new_n256), .A2(new_n258), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n209), .A2(G33), .ZN(new_n260));
  NAND2_X1  g0060(.A1(new_n259), .A2(new_n260), .ZN(new_n261));
  INV_X1    g0061(.A(new_n261), .ZN(new_n262));
  AOI21_X1  g0062(.A(new_n255), .B1(new_n262), .B2(G116), .ZN(new_n263));
  NAND2_X1  g0063(.A1(G33), .A2(G283), .ZN(new_n264));
  OAI211_X1 g0064(.A(new_n264), .B(new_n210), .C1(G33), .C2(new_n205), .ZN(new_n265));
  OAI211_X1 g0065(.A(new_n265), .B(new_n258), .C1(new_n210), .C2(G116), .ZN(new_n266));
  INV_X1    g0066(.A(KEYINPUT20), .ZN(new_n267));
  XNOR2_X1  g0067(.A(new_n266), .B(new_n267), .ZN(new_n268));
  AOI21_X1  g0068(.A(new_n253), .B1(new_n263), .B2(new_n268), .ZN(new_n269));
  AOI21_X1  g0069(.A(new_n230), .B1(G33), .B2(G41), .ZN(new_n270));
  INV_X1    g0070(.A(new_n270), .ZN(new_n271));
  INV_X1    g0071(.A(G1698), .ZN(new_n272));
  INV_X1    g0072(.A(KEYINPUT3), .ZN(new_n273));
  INV_X1    g0073(.A(KEYINPUT70), .ZN(new_n274));
  INV_X1    g0074(.A(G33), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n274), .A2(new_n275), .ZN(new_n276));
  NAND2_X1  g0076(.A1(KEYINPUT70), .A2(G33), .ZN(new_n277));
  AOI21_X1  g0077(.A(new_n273), .B1(new_n276), .B2(new_n277), .ZN(new_n278));
  NOR2_X1   g0078(.A1(KEYINPUT3), .A2(G33), .ZN(new_n279));
  OAI211_X1 g0079(.A(G257), .B(new_n272), .C1(new_n278), .C2(new_n279), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n280), .A2(KEYINPUT81), .ZN(new_n281));
  AND2_X1   g0081(.A1(KEYINPUT70), .A2(G33), .ZN(new_n282));
  NOR2_X1   g0082(.A1(KEYINPUT70), .A2(G33), .ZN(new_n283));
  OAI21_X1  g0083(.A(KEYINPUT3), .B1(new_n282), .B2(new_n283), .ZN(new_n284));
  INV_X1    g0084(.A(new_n279), .ZN(new_n285));
  AOI21_X1  g0085(.A(G1698), .B1(new_n284), .B2(new_n285), .ZN(new_n286));
  INV_X1    g0086(.A(KEYINPUT81), .ZN(new_n287));
  NAND3_X1  g0087(.A1(new_n286), .A2(new_n287), .A3(G257), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n281), .A2(new_n288), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n284), .A2(new_n285), .ZN(new_n290));
  NAND3_X1  g0090(.A1(new_n290), .A2(G264), .A3(G1698), .ZN(new_n291));
  NAND2_X1  g0091(.A1(KEYINPUT3), .A2(G33), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n285), .A2(new_n292), .ZN(new_n293));
  INV_X1    g0093(.A(new_n293), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n294), .A2(G303), .ZN(new_n295));
  AND2_X1   g0095(.A1(new_n291), .A2(new_n295), .ZN(new_n296));
  AOI21_X1  g0096(.A(new_n271), .B1(new_n289), .B2(new_n296), .ZN(new_n297));
  INV_X1    g0097(.A(G41), .ZN(new_n298));
  AND3_X1   g0098(.A1(new_n298), .A2(KEYINPUT75), .A3(KEYINPUT5), .ZN(new_n299));
  AOI21_X1  g0099(.A(KEYINPUT75), .B1(new_n298), .B2(KEYINPUT5), .ZN(new_n300));
  NOR2_X1   g0100(.A1(new_n299), .A2(new_n300), .ZN(new_n301));
  INV_X1    g0101(.A(G45), .ZN(new_n302));
  NOR2_X1   g0102(.A1(new_n302), .A2(G1), .ZN(new_n303));
  INV_X1    g0103(.A(KEYINPUT74), .ZN(new_n304));
  INV_X1    g0104(.A(KEYINPUT5), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n305), .A2(G41), .ZN(new_n306));
  NAND3_X1  g0106(.A1(new_n303), .A2(new_n304), .A3(new_n306), .ZN(new_n307));
  OAI211_X1 g0107(.A(new_n209), .B(G45), .C1(new_n298), .C2(KEYINPUT5), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n308), .A2(KEYINPUT74), .ZN(new_n309));
  INV_X1    g0109(.A(G274), .ZN(new_n310));
  INV_X1    g0110(.A(new_n230), .ZN(new_n311));
  NAND2_X1  g0111(.A1(G33), .A2(G41), .ZN(new_n312));
  AOI21_X1  g0112(.A(new_n310), .B1(new_n311), .B2(new_n312), .ZN(new_n313));
  NAND4_X1  g0113(.A1(new_n301), .A2(new_n307), .A3(new_n309), .A4(new_n313), .ZN(new_n314));
  INV_X1    g0114(.A(KEYINPUT75), .ZN(new_n315));
  OAI21_X1  g0115(.A(new_n315), .B1(new_n305), .B2(G41), .ZN(new_n316));
  NAND3_X1  g0116(.A1(new_n298), .A2(KEYINPUT75), .A3(KEYINPUT5), .ZN(new_n317));
  NAND4_X1  g0117(.A1(new_n316), .A2(new_n317), .A3(new_n303), .A4(new_n306), .ZN(new_n318));
  NAND3_X1  g0118(.A1(new_n318), .A2(new_n271), .A3(G270), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n314), .A2(new_n319), .ZN(new_n320));
  OAI211_X1 g0120(.A(new_n269), .B(KEYINPUT21), .C1(new_n297), .C2(new_n320), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n321), .A2(KEYINPUT82), .ZN(new_n322));
  INV_X1    g0122(.A(new_n320), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n291), .A2(new_n295), .ZN(new_n324));
  AOI21_X1  g0124(.A(new_n324), .B1(new_n288), .B2(new_n281), .ZN(new_n325));
  OAI21_X1  g0125(.A(new_n323), .B1(new_n325), .B2(new_n271), .ZN(new_n326));
  INV_X1    g0126(.A(KEYINPUT82), .ZN(new_n327));
  NAND4_X1  g0127(.A1(new_n326), .A2(new_n327), .A3(KEYINPUT21), .A4(new_n269), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n322), .A2(new_n328), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n326), .A2(G200), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n263), .A2(new_n268), .ZN(new_n331));
  INV_X1    g0131(.A(new_n331), .ZN(new_n332));
  INV_X1    g0132(.A(G190), .ZN(new_n333));
  OAI211_X1 g0133(.A(new_n330), .B(new_n332), .C1(new_n333), .C2(new_n326), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n326), .A2(new_n269), .ZN(new_n335));
  XNOR2_X1  g0135(.A(KEYINPUT83), .B(KEYINPUT21), .ZN(new_n336));
  INV_X1    g0136(.A(G179), .ZN(new_n337));
  NOR2_X1   g0137(.A1(new_n320), .A2(new_n337), .ZN(new_n338));
  INV_X1    g0138(.A(new_n338), .ZN(new_n339));
  NOR2_X1   g0139(.A1(new_n297), .A2(new_n339), .ZN(new_n340));
  AOI22_X1  g0140(.A1(new_n335), .A2(new_n336), .B1(new_n331), .B2(new_n340), .ZN(new_n341));
  AND3_X1   g0141(.A1(new_n329), .A2(new_n334), .A3(new_n341), .ZN(new_n342));
  XNOR2_X1  g0142(.A(KEYINPUT8), .B(G58), .ZN(new_n343));
  NOR2_X1   g0143(.A1(new_n275), .A2(G20), .ZN(new_n344));
  INV_X1    g0144(.A(new_n344), .ZN(new_n345));
  INV_X1    g0145(.A(G150), .ZN(new_n346));
  NOR2_X1   g0146(.A1(G20), .A2(G33), .ZN(new_n347));
  INV_X1    g0147(.A(new_n347), .ZN(new_n348));
  OAI22_X1  g0148(.A1(new_n343), .A2(new_n345), .B1(new_n346), .B2(new_n348), .ZN(new_n349));
  AOI21_X1  g0149(.A(new_n349), .B1(G20), .B2(new_n203), .ZN(new_n350));
  INV_X1    g0150(.A(new_n258), .ZN(new_n351));
  NOR2_X1   g0151(.A1(new_n350), .A2(new_n351), .ZN(new_n352));
  INV_X1    g0152(.A(KEYINPUT9), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n351), .A2(new_n254), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n209), .A2(G20), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n355), .A2(G50), .ZN(new_n356));
  OAI22_X1  g0156(.A1(new_n354), .A2(new_n356), .B1(G50), .B2(new_n254), .ZN(new_n357));
  NOR3_X1   g0157(.A1(new_n352), .A2(new_n353), .A3(new_n357), .ZN(new_n358));
  INV_X1    g0158(.A(new_n358), .ZN(new_n359));
  AOI21_X1  g0159(.A(G1), .B1(new_n298), .B2(new_n302), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n313), .A2(new_n360), .ZN(new_n361));
  NOR2_X1   g0161(.A1(new_n270), .A2(new_n360), .ZN(new_n362));
  INV_X1    g0162(.A(new_n362), .ZN(new_n363));
  INV_X1    g0163(.A(G226), .ZN(new_n364));
  OAI21_X1  g0164(.A(new_n361), .B1(new_n363), .B2(new_n364), .ZN(new_n365));
  NAND3_X1  g0165(.A1(new_n293), .A2(G222), .A3(new_n272), .ZN(new_n366));
  INV_X1    g0166(.A(G77), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n293), .A2(G1698), .ZN(new_n368));
  INV_X1    g0168(.A(G223), .ZN(new_n369));
  OAI221_X1 g0169(.A(new_n366), .B1(new_n367), .B2(new_n293), .C1(new_n368), .C2(new_n369), .ZN(new_n370));
  AOI21_X1  g0170(.A(new_n365), .B1(new_n370), .B2(new_n270), .ZN(new_n371));
  INV_X1    g0171(.A(G200), .ZN(new_n372));
  OR2_X1    g0172(.A1(new_n371), .A2(new_n372), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n371), .A2(G190), .ZN(new_n374));
  OAI21_X1  g0174(.A(new_n353), .B1(new_n352), .B2(new_n357), .ZN(new_n375));
  NAND4_X1  g0175(.A1(new_n359), .A2(new_n373), .A3(new_n374), .A4(new_n375), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n376), .A2(KEYINPUT10), .ZN(new_n377));
  INV_X1    g0177(.A(new_n375), .ZN(new_n378));
  NOR2_X1   g0178(.A1(new_n378), .A2(new_n358), .ZN(new_n379));
  INV_X1    g0179(.A(KEYINPUT10), .ZN(new_n380));
  NAND4_X1  g0180(.A1(new_n379), .A2(new_n380), .A3(new_n374), .A4(new_n373), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n377), .A2(new_n381), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n256), .A2(new_n247), .ZN(new_n383));
  XNOR2_X1  g0183(.A(new_n383), .B(KEYINPUT12), .ZN(new_n384));
  AOI22_X1  g0184(.A1(new_n347), .A2(G50), .B1(G20), .B2(new_n247), .ZN(new_n385));
  OAI21_X1  g0185(.A(new_n385), .B1(new_n345), .B2(new_n367), .ZN(new_n386));
  NAND3_X1  g0186(.A1(new_n386), .A2(KEYINPUT11), .A3(new_n258), .ZN(new_n387));
  NAND3_X1  g0187(.A1(new_n259), .A2(G68), .A3(new_n355), .ZN(new_n388));
  NAND3_X1  g0188(.A1(new_n384), .A2(new_n387), .A3(new_n388), .ZN(new_n389));
  AOI21_X1  g0189(.A(KEYINPUT11), .B1(new_n386), .B2(new_n258), .ZN(new_n390));
  NOR2_X1   g0190(.A1(new_n389), .A2(new_n390), .ZN(new_n391));
  INV_X1    g0191(.A(new_n391), .ZN(new_n392));
  INV_X1    g0192(.A(KEYINPUT13), .ZN(new_n393));
  AND2_X1   g0193(.A1(KEYINPUT3), .A2(G33), .ZN(new_n394));
  OAI211_X1 g0194(.A(G232), .B(G1698), .C1(new_n394), .C2(new_n279), .ZN(new_n395));
  OAI211_X1 g0195(.A(G226), .B(new_n272), .C1(new_n394), .C2(new_n279), .ZN(new_n396));
  NAND2_X1  g0196(.A1(G33), .A2(G97), .ZN(new_n397));
  NAND3_X1  g0197(.A1(new_n395), .A2(new_n396), .A3(new_n397), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n398), .A2(new_n270), .ZN(new_n399));
  AOI22_X1  g0199(.A1(new_n362), .A2(G238), .B1(new_n313), .B2(new_n360), .ZN(new_n400));
  AOI21_X1  g0200(.A(new_n393), .B1(new_n399), .B2(new_n400), .ZN(new_n401));
  INV_X1    g0201(.A(new_n401), .ZN(new_n402));
  NAND3_X1  g0202(.A1(new_n399), .A2(new_n400), .A3(new_n393), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n402), .A2(new_n403), .ZN(new_n404));
  INV_X1    g0204(.A(new_n404), .ZN(new_n405));
  AOI21_X1  g0205(.A(new_n392), .B1(new_n405), .B2(G190), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n404), .A2(G200), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n406), .A2(new_n407), .ZN(new_n408));
  OAI21_X1  g0208(.A(KEYINPUT69), .B1(new_n371), .B2(G169), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n371), .A2(new_n337), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n409), .A2(new_n410), .ZN(new_n411));
  INV_X1    g0211(.A(KEYINPUT69), .ZN(new_n412));
  OAI221_X1 g0212(.A(new_n411), .B1(new_n412), .B2(new_n410), .C1(new_n352), .C2(new_n357), .ZN(new_n413));
  NAND3_X1  g0213(.A1(new_n259), .A2(G77), .A3(new_n355), .ZN(new_n414));
  OAI21_X1  g0214(.A(new_n414), .B1(G77), .B2(new_n254), .ZN(new_n415));
  INV_X1    g0215(.A(G58), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n416), .A2(KEYINPUT8), .ZN(new_n417));
  INV_X1    g0217(.A(KEYINPUT8), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n418), .A2(G58), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n417), .A2(new_n419), .ZN(new_n420));
  AOI22_X1  g0220(.A1(new_n420), .A2(new_n347), .B1(G20), .B2(G77), .ZN(new_n421));
  XNOR2_X1  g0221(.A(KEYINPUT15), .B(G87), .ZN(new_n422));
  INV_X1    g0222(.A(new_n422), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n423), .A2(new_n344), .ZN(new_n424));
  AOI21_X1  g0224(.A(new_n351), .B1(new_n421), .B2(new_n424), .ZN(new_n425));
  NOR2_X1   g0225(.A1(new_n415), .A2(new_n425), .ZN(new_n426));
  INV_X1    g0226(.A(new_n426), .ZN(new_n427));
  INV_X1    g0227(.A(G244), .ZN(new_n428));
  OAI21_X1  g0228(.A(new_n361), .B1(new_n363), .B2(new_n428), .ZN(new_n429));
  NAND3_X1  g0229(.A1(new_n293), .A2(G232), .A3(new_n272), .ZN(new_n430));
  INV_X1    g0230(.A(G238), .ZN(new_n431));
  OAI221_X1 g0231(.A(new_n430), .B1(new_n206), .B2(new_n293), .C1(new_n368), .C2(new_n431), .ZN(new_n432));
  AOI21_X1  g0232(.A(new_n429), .B1(new_n432), .B2(new_n270), .ZN(new_n433));
  OAI21_X1  g0233(.A(new_n427), .B1(new_n433), .B2(G169), .ZN(new_n434));
  AND2_X1   g0234(.A1(new_n433), .A2(new_n337), .ZN(new_n435));
  OR2_X1    g0235(.A1(new_n434), .A2(new_n435), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n433), .A2(G190), .ZN(new_n437));
  OAI211_X1 g0237(.A(new_n437), .B(new_n426), .C1(new_n372), .C2(new_n433), .ZN(new_n438));
  AND2_X1   g0238(.A1(new_n436), .A2(new_n438), .ZN(new_n439));
  NAND4_X1  g0239(.A1(new_n382), .A2(new_n408), .A3(new_n413), .A4(new_n439), .ZN(new_n440));
  NAND3_X1  g0240(.A1(new_n284), .A2(new_n210), .A3(new_n285), .ZN(new_n441));
  NAND2_X1  g0241(.A1(new_n441), .A2(KEYINPUT7), .ZN(new_n442));
  INV_X1    g0242(.A(KEYINPUT7), .ZN(new_n443));
  NAND4_X1  g0243(.A1(new_n284), .A2(new_n443), .A3(new_n210), .A4(new_n285), .ZN(new_n444));
  NAND3_X1  g0244(.A1(new_n442), .A2(G68), .A3(new_n444), .ZN(new_n445));
  INV_X1    g0245(.A(KEYINPUT71), .ZN(new_n446));
  INV_X1    g0246(.A(G159), .ZN(new_n447));
  OAI21_X1  g0247(.A(new_n446), .B1(new_n348), .B2(new_n447), .ZN(new_n448));
  NAND3_X1  g0248(.A1(new_n347), .A2(KEYINPUT71), .A3(G159), .ZN(new_n449));
  NAND2_X1  g0249(.A1(new_n448), .A2(new_n449), .ZN(new_n450));
  NOR2_X1   g0250(.A1(new_n416), .A2(new_n247), .ZN(new_n451));
  OAI21_X1  g0251(.A(G20), .B1(new_n451), .B2(new_n201), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n450), .A2(new_n452), .ZN(new_n453));
  INV_X1    g0253(.A(new_n453), .ZN(new_n454));
  NAND3_X1  g0254(.A1(new_n445), .A2(KEYINPUT16), .A3(new_n454), .ZN(new_n455));
  INV_X1    g0255(.A(KEYINPUT16), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n292), .A2(new_n210), .ZN(new_n457));
  NOR2_X1   g0257(.A1(new_n457), .A2(new_n443), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n276), .A2(new_n277), .ZN(new_n459));
  OAI21_X1  g0259(.A(new_n458), .B1(KEYINPUT3), .B2(new_n459), .ZN(new_n460));
  OAI21_X1  g0260(.A(new_n443), .B1(new_n457), .B2(new_n279), .ZN(new_n461));
  AOI21_X1  g0261(.A(new_n247), .B1(new_n460), .B2(new_n461), .ZN(new_n462));
  OAI21_X1  g0262(.A(new_n456), .B1(new_n462), .B2(new_n453), .ZN(new_n463));
  NAND3_X1  g0263(.A1(new_n455), .A2(new_n258), .A3(new_n463), .ZN(new_n464));
  NAND2_X1  g0264(.A1(new_n420), .A2(new_n355), .ZN(new_n465));
  OAI22_X1  g0265(.A1(new_n354), .A2(new_n465), .B1(new_n254), .B2(new_n420), .ZN(new_n466));
  INV_X1    g0266(.A(KEYINPUT72), .ZN(new_n467));
  XNOR2_X1  g0267(.A(new_n466), .B(new_n467), .ZN(new_n468));
  INV_X1    g0268(.A(new_n468), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n464), .A2(new_n469), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n364), .A2(G1698), .ZN(new_n471));
  OAI21_X1  g0271(.A(new_n471), .B1(G223), .B2(G1698), .ZN(new_n472));
  INV_X1    g0272(.A(new_n472), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n290), .A2(new_n473), .ZN(new_n474));
  NAND2_X1  g0274(.A1(G33), .A2(G87), .ZN(new_n475));
  AOI21_X1  g0275(.A(new_n271), .B1(new_n474), .B2(new_n475), .ZN(new_n476));
  AOI22_X1  g0276(.A1(new_n362), .A2(G232), .B1(new_n313), .B2(new_n360), .ZN(new_n477));
  INV_X1    g0277(.A(new_n477), .ZN(new_n478));
  OAI21_X1  g0278(.A(new_n253), .B1(new_n476), .B2(new_n478), .ZN(new_n479));
  AOI21_X1  g0279(.A(new_n472), .B1(new_n285), .B2(new_n284), .ZN(new_n480));
  INV_X1    g0280(.A(new_n475), .ZN(new_n481));
  OAI21_X1  g0281(.A(new_n270), .B1(new_n480), .B2(new_n481), .ZN(new_n482));
  NAND3_X1  g0282(.A1(new_n482), .A2(new_n337), .A3(new_n477), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n479), .A2(new_n483), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n484), .A2(KEYINPUT73), .ZN(new_n485));
  INV_X1    g0285(.A(KEYINPUT73), .ZN(new_n486));
  NAND3_X1  g0286(.A1(new_n479), .A2(new_n486), .A3(new_n483), .ZN(new_n487));
  NAND3_X1  g0287(.A1(new_n470), .A2(new_n485), .A3(new_n487), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n488), .A2(KEYINPUT18), .ZN(new_n489));
  AOI21_X1  g0289(.A(new_n247), .B1(new_n441), .B2(KEYINPUT7), .ZN(new_n490));
  AOI21_X1  g0290(.A(new_n453), .B1(new_n490), .B2(new_n444), .ZN(new_n491));
  AOI21_X1  g0291(.A(new_n351), .B1(new_n491), .B2(KEYINPUT16), .ZN(new_n492));
  AOI21_X1  g0292(.A(new_n468), .B1(new_n492), .B2(new_n463), .ZN(new_n493));
  OAI21_X1  g0293(.A(new_n372), .B1(new_n476), .B2(new_n478), .ZN(new_n494));
  NAND3_X1  g0294(.A1(new_n482), .A2(new_n333), .A3(new_n477), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n493), .A2(new_n496), .ZN(new_n497));
  INV_X1    g0297(.A(KEYINPUT17), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  INV_X1    g0299(.A(KEYINPUT18), .ZN(new_n500));
  NAND4_X1  g0300(.A1(new_n470), .A2(new_n485), .A3(new_n500), .A4(new_n487), .ZN(new_n501));
  AND3_X1   g0301(.A1(new_n496), .A2(new_n464), .A3(new_n469), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n502), .A2(KEYINPUT17), .ZN(new_n503));
  NAND4_X1  g0303(.A1(new_n489), .A2(new_n499), .A3(new_n501), .A4(new_n503), .ZN(new_n504));
  INV_X1    g0304(.A(KEYINPUT14), .ZN(new_n505));
  AND3_X1   g0305(.A1(new_n399), .A2(new_n400), .A3(new_n393), .ZN(new_n506));
  OAI211_X1 g0306(.A(new_n505), .B(G169), .C1(new_n506), .C2(new_n401), .ZN(new_n507));
  OAI21_X1  g0307(.A(new_n507), .B1(new_n404), .B2(new_n337), .ZN(new_n508));
  AOI21_X1  g0308(.A(new_n505), .B1(new_n404), .B2(G169), .ZN(new_n509));
  OAI21_X1  g0309(.A(new_n392), .B1(new_n508), .B2(new_n509), .ZN(new_n510));
  INV_X1    g0310(.A(new_n510), .ZN(new_n511));
  OR3_X1    g0311(.A1(new_n440), .A2(new_n504), .A3(new_n511), .ZN(new_n512));
  INV_X1    g0312(.A(new_n512), .ZN(new_n513));
  NAND3_X1  g0313(.A1(new_n318), .A2(new_n271), .A3(G257), .ZN(new_n514));
  AND2_X1   g0314(.A1(new_n314), .A2(new_n514), .ZN(new_n515));
  AND2_X1   g0315(.A1(KEYINPUT4), .A2(G244), .ZN(new_n516));
  OAI211_X1 g0316(.A(new_n272), .B(new_n516), .C1(new_n394), .C2(new_n279), .ZN(new_n517));
  OAI211_X1 g0317(.A(G250), .B(G1698), .C1(new_n394), .C2(new_n279), .ZN(new_n518));
  NAND3_X1  g0318(.A1(new_n517), .A2(new_n518), .A3(new_n264), .ZN(new_n519));
  OAI211_X1 g0319(.A(G244), .B(new_n272), .C1(new_n278), .C2(new_n279), .ZN(new_n520));
  INV_X1    g0320(.A(KEYINPUT4), .ZN(new_n521));
  AOI21_X1  g0321(.A(new_n519), .B1(new_n520), .B2(new_n521), .ZN(new_n522));
  OAI211_X1 g0322(.A(new_n515), .B(new_n337), .C1(new_n522), .C2(new_n271), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n523), .A2(KEYINPUT76), .ZN(new_n524));
  NOR2_X1   g0324(.A1(new_n522), .A2(new_n271), .ZN(new_n525));
  INV_X1    g0325(.A(new_n515), .ZN(new_n526));
  OAI21_X1  g0326(.A(new_n253), .B1(new_n525), .B2(new_n526), .ZN(new_n527));
  AOI21_X1  g0327(.A(new_n428), .B1(new_n284), .B2(new_n285), .ZN(new_n528));
  AOI21_X1  g0328(.A(KEYINPUT4), .B1(new_n528), .B2(new_n272), .ZN(new_n529));
  OAI21_X1  g0329(.A(new_n270), .B1(new_n529), .B2(new_n519), .ZN(new_n530));
  INV_X1    g0330(.A(KEYINPUT76), .ZN(new_n531));
  NAND4_X1  g0331(.A1(new_n530), .A2(new_n531), .A3(new_n337), .A4(new_n515), .ZN(new_n532));
  AOI21_X1  g0332(.A(new_n206), .B1(new_n460), .B2(new_n461), .ZN(new_n533));
  INV_X1    g0333(.A(KEYINPUT6), .ZN(new_n534));
  NOR3_X1   g0334(.A1(new_n534), .A2(new_n205), .A3(G107), .ZN(new_n535));
  XNOR2_X1  g0335(.A(G97), .B(G107), .ZN(new_n536));
  AOI21_X1  g0336(.A(new_n535), .B1(new_n534), .B2(new_n536), .ZN(new_n537));
  OAI22_X1  g0337(.A1(new_n537), .A2(new_n210), .B1(new_n367), .B2(new_n348), .ZN(new_n538));
  OAI21_X1  g0338(.A(new_n258), .B1(new_n533), .B2(new_n538), .ZN(new_n539));
  NOR2_X1   g0339(.A1(new_n254), .A2(G97), .ZN(new_n540));
  AOI21_X1  g0340(.A(new_n540), .B1(new_n262), .B2(G97), .ZN(new_n541));
  NAND2_X1  g0341(.A1(new_n539), .A2(new_n541), .ZN(new_n542));
  NAND4_X1  g0342(.A1(new_n524), .A2(new_n527), .A3(new_n532), .A4(new_n542), .ZN(new_n543));
  OAI21_X1  g0343(.A(G200), .B1(new_n525), .B2(new_n526), .ZN(new_n544));
  NAND3_X1  g0344(.A1(new_n530), .A2(G190), .A3(new_n515), .ZN(new_n545));
  NAND4_X1  g0345(.A1(new_n544), .A2(new_n539), .A3(new_n541), .A4(new_n545), .ZN(new_n546));
  AND2_X1   g0346(.A1(new_n543), .A2(new_n546), .ZN(new_n547));
  NAND4_X1  g0347(.A1(new_n290), .A2(KEYINPUT22), .A3(new_n210), .A4(G87), .ZN(new_n548));
  INV_X1    g0348(.A(KEYINPUT22), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n210), .A2(G87), .ZN(new_n550));
  OAI21_X1  g0350(.A(new_n549), .B1(new_n294), .B2(new_n550), .ZN(new_n551));
  INV_X1    g0351(.A(G116), .ZN(new_n552));
  AOI21_X1  g0352(.A(new_n552), .B1(new_n276), .B2(new_n277), .ZN(new_n553));
  INV_X1    g0353(.A(KEYINPUT23), .ZN(new_n554));
  OAI21_X1  g0354(.A(new_n554), .B1(new_n210), .B2(G107), .ZN(new_n555));
  NAND3_X1  g0355(.A1(new_n206), .A2(KEYINPUT23), .A3(G20), .ZN(new_n556));
  AOI22_X1  g0356(.A1(new_n553), .A2(new_n210), .B1(new_n555), .B2(new_n556), .ZN(new_n557));
  NAND3_X1  g0357(.A1(new_n548), .A2(new_n551), .A3(new_n557), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n558), .A2(KEYINPUT24), .ZN(new_n559));
  INV_X1    g0359(.A(KEYINPUT24), .ZN(new_n560));
  NAND4_X1  g0360(.A1(new_n548), .A2(new_n551), .A3(new_n560), .A4(new_n557), .ZN(new_n561));
  AOI21_X1  g0361(.A(new_n351), .B1(new_n559), .B2(new_n561), .ZN(new_n562));
  AND3_X1   g0362(.A1(new_n256), .A2(KEYINPUT25), .A3(new_n206), .ZN(new_n563));
  AOI21_X1  g0363(.A(KEYINPUT25), .B1(new_n256), .B2(new_n206), .ZN(new_n564));
  OAI22_X1  g0364(.A1(new_n261), .A2(new_n206), .B1(new_n563), .B2(new_n564), .ZN(new_n565));
  NOR2_X1   g0365(.A1(new_n562), .A2(new_n565), .ZN(new_n566));
  NAND3_X1  g0366(.A1(new_n290), .A2(G250), .A3(new_n272), .ZN(new_n567));
  OAI211_X1 g0367(.A(G257), .B(G1698), .C1(new_n278), .C2(new_n279), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n459), .A2(G294), .ZN(new_n569));
  NAND3_X1  g0369(.A1(new_n567), .A2(new_n568), .A3(new_n569), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n570), .A2(new_n270), .ZN(new_n571));
  NAND3_X1  g0371(.A1(new_n318), .A2(new_n271), .A3(G264), .ZN(new_n572));
  INV_X1    g0372(.A(KEYINPUT84), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n572), .A2(new_n573), .ZN(new_n574));
  NAND4_X1  g0374(.A1(new_n318), .A2(new_n271), .A3(KEYINPUT84), .A4(G264), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  NAND3_X1  g0376(.A1(new_n571), .A2(new_n314), .A3(new_n576), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n577), .A2(G200), .ZN(new_n578));
  OAI211_X1 g0378(.A(new_n566), .B(new_n578), .C1(new_n333), .C2(new_n577), .ZN(new_n579));
  AND2_X1   g0379(.A1(new_n547), .A2(new_n579), .ZN(new_n580));
  NAND3_X1  g0380(.A1(new_n577), .A2(KEYINPUT85), .A3(G169), .ZN(new_n581));
  AOI22_X1  g0381(.A1(new_n570), .A2(new_n270), .B1(new_n574), .B2(new_n575), .ZN(new_n582));
  NAND3_X1  g0382(.A1(new_n582), .A2(G179), .A3(new_n314), .ZN(new_n583));
  AND2_X1   g0383(.A1(new_n581), .A2(new_n583), .ZN(new_n584));
  AOI21_X1  g0384(.A(new_n253), .B1(new_n582), .B2(new_n314), .ZN(new_n585));
  OR2_X1    g0385(.A1(new_n585), .A2(KEYINPUT85), .ZN(new_n586));
  AOI21_X1  g0386(.A(new_n566), .B1(new_n584), .B2(new_n586), .ZN(new_n587));
  OAI211_X1 g0387(.A(G244), .B(G1698), .C1(new_n278), .C2(new_n279), .ZN(new_n588));
  OAI211_X1 g0388(.A(G238), .B(new_n272), .C1(new_n278), .C2(new_n279), .ZN(new_n589));
  INV_X1    g0389(.A(new_n553), .ZN(new_n590));
  NAND3_X1  g0390(.A1(new_n588), .A2(new_n589), .A3(new_n590), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n591), .A2(new_n270), .ZN(new_n592));
  OR2_X1    g0392(.A1(new_n303), .A2(G250), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n303), .A2(new_n310), .ZN(new_n594));
  NAND3_X1  g0394(.A1(new_n593), .A2(new_n271), .A3(new_n594), .ZN(new_n595));
  AOI21_X1  g0395(.A(G169), .B1(new_n592), .B2(new_n595), .ZN(new_n596));
  INV_X1    g0396(.A(new_n595), .ZN(new_n597));
  AOI211_X1 g0397(.A(G179), .B(new_n597), .C1(new_n591), .C2(new_n270), .ZN(new_n598));
  OAI21_X1  g0398(.A(KEYINPUT77), .B1(new_n596), .B2(new_n598), .ZN(new_n599));
  AOI211_X1 g0399(.A(G20), .B(new_n247), .C1(new_n284), .C2(new_n285), .ZN(new_n600));
  OR2_X1    g0400(.A1(KEYINPUT78), .A2(G87), .ZN(new_n601));
  NOR2_X1   g0401(.A1(G97), .A2(G107), .ZN(new_n602));
  NAND2_X1  g0402(.A1(KEYINPUT78), .A2(G87), .ZN(new_n603));
  NAND3_X1  g0403(.A1(new_n601), .A2(new_n602), .A3(new_n603), .ZN(new_n604));
  INV_X1    g0404(.A(KEYINPUT19), .ZN(new_n605));
  AOI21_X1  g0405(.A(new_n605), .B1(new_n397), .B2(new_n210), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n604), .A2(new_n606), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n344), .A2(G97), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n608), .A2(new_n605), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n607), .A2(new_n609), .ZN(new_n610));
  OAI21_X1  g0410(.A(new_n258), .B1(new_n600), .B2(new_n610), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n422), .A2(new_n256), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n262), .A2(new_n423), .ZN(new_n613));
  NAND3_X1  g0413(.A1(new_n611), .A2(new_n612), .A3(new_n613), .ZN(new_n614));
  INV_X1    g0414(.A(KEYINPUT79), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  NAND4_X1  g0416(.A1(new_n611), .A2(new_n613), .A3(KEYINPUT79), .A4(new_n612), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  AOI21_X1  g0418(.A(new_n553), .B1(new_n286), .B2(G238), .ZN(new_n619));
  AOI21_X1  g0419(.A(new_n271), .B1(new_n619), .B2(new_n588), .ZN(new_n620));
  OAI21_X1  g0420(.A(new_n253), .B1(new_n620), .B2(new_n597), .ZN(new_n621));
  INV_X1    g0421(.A(KEYINPUT77), .ZN(new_n622));
  NAND3_X1  g0422(.A1(new_n592), .A2(new_n337), .A3(new_n595), .ZN(new_n623));
  NAND3_X1  g0423(.A1(new_n621), .A2(new_n622), .A3(new_n623), .ZN(new_n624));
  NAND3_X1  g0424(.A1(new_n599), .A2(new_n618), .A3(new_n624), .ZN(new_n625));
  OAI21_X1  g0425(.A(G200), .B1(new_n620), .B2(new_n597), .ZN(new_n626));
  NAND3_X1  g0426(.A1(new_n290), .A2(new_n210), .A3(G68), .ZN(new_n627));
  AOI22_X1  g0427(.A1(new_n604), .A2(new_n606), .B1(new_n608), .B2(new_n605), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  AOI22_X1  g0429(.A1(new_n629), .A2(new_n258), .B1(new_n256), .B2(new_n422), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n262), .A2(G87), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n630), .A2(new_n631), .ZN(new_n632));
  INV_X1    g0432(.A(new_n632), .ZN(new_n633));
  AND4_X1   g0433(.A1(KEYINPUT80), .A2(new_n592), .A3(G190), .A4(new_n595), .ZN(new_n634));
  AOI21_X1  g0434(.A(new_n597), .B1(new_n591), .B2(new_n270), .ZN(new_n635));
  AOI21_X1  g0435(.A(KEYINPUT80), .B1(new_n635), .B2(G190), .ZN(new_n636));
  OAI211_X1 g0436(.A(new_n626), .B(new_n633), .C1(new_n634), .C2(new_n636), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n625), .A2(new_n637), .ZN(new_n638));
  NOR2_X1   g0438(.A1(new_n587), .A2(new_n638), .ZN(new_n639));
  AND4_X1   g0439(.A1(new_n342), .A2(new_n513), .A3(new_n580), .A4(new_n639), .ZN(G372));
  INV_X1    g0440(.A(KEYINPUT88), .ZN(new_n641));
  NOR2_X1   g0441(.A1(new_n382), .A2(new_n641), .ZN(new_n642));
  AOI21_X1  g0442(.A(KEYINPUT88), .B1(new_n377), .B2(new_n381), .ZN(new_n643));
  OR2_X1    g0443(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  INV_X1    g0444(.A(new_n436), .ZN(new_n645));
  AOI21_X1  g0445(.A(new_n511), .B1(new_n408), .B2(new_n645), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n499), .A2(new_n503), .ZN(new_n647));
  NOR2_X1   g0447(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n489), .A2(new_n501), .ZN(new_n649));
  OAI21_X1  g0449(.A(new_n644), .B1(new_n648), .B2(new_n649), .ZN(new_n650));
  AND2_X1   g0450(.A1(new_n650), .A2(new_n413), .ZN(new_n651));
  AND3_X1   g0451(.A1(new_n591), .A2(KEYINPUT86), .A3(new_n270), .ZN(new_n652));
  AOI21_X1  g0452(.A(KEYINPUT86), .B1(new_n591), .B2(new_n270), .ZN(new_n653));
  OAI21_X1  g0453(.A(new_n595), .B1(new_n652), .B2(new_n653), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n654), .A2(new_n253), .ZN(new_n655));
  AOI21_X1  g0455(.A(new_n598), .B1(new_n616), .B2(new_n617), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n329), .A2(new_n341), .ZN(new_n658));
  NOR2_X1   g0458(.A1(new_n658), .A2(new_n587), .ZN(new_n659));
  NAND3_X1  g0459(.A1(new_n592), .A2(G190), .A3(new_n595), .ZN(new_n660));
  INV_X1    g0460(.A(KEYINPUT80), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  NAND3_X1  g0462(.A1(new_n635), .A2(KEYINPUT80), .A3(G190), .ZN(new_n663));
  AOI21_X1  g0463(.A(new_n632), .B1(new_n662), .B2(new_n663), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n654), .A2(G200), .ZN(new_n665));
  AOI22_X1  g0465(.A1(new_n664), .A2(new_n665), .B1(new_n655), .B2(new_n656), .ZN(new_n666));
  NAND3_X1  g0466(.A1(new_n666), .A2(new_n579), .A3(new_n547), .ZN(new_n667));
  OAI21_X1  g0467(.A(new_n657), .B1(new_n659), .B2(new_n667), .ZN(new_n668));
  AND4_X1   g0468(.A1(new_n524), .A2(new_n527), .A3(new_n532), .A4(new_n542), .ZN(new_n669));
  AND4_X1   g0469(.A1(KEYINPUT26), .A2(new_n625), .A3(new_n669), .A4(new_n637), .ZN(new_n670));
  NAND3_X1  g0470(.A1(new_n524), .A2(new_n527), .A3(new_n532), .ZN(new_n671));
  INV_X1    g0471(.A(KEYINPUT87), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  NAND4_X1  g0473(.A1(new_n524), .A2(new_n527), .A3(KEYINPUT87), .A4(new_n532), .ZN(new_n674));
  NAND4_X1  g0474(.A1(new_n666), .A2(new_n542), .A3(new_n673), .A4(new_n674), .ZN(new_n675));
  INV_X1    g0475(.A(KEYINPUT26), .ZN(new_n676));
  AOI21_X1  g0476(.A(new_n670), .B1(new_n675), .B2(new_n676), .ZN(new_n677));
  OAI21_X1  g0477(.A(new_n513), .B1(new_n668), .B2(new_n677), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n651), .A2(new_n678), .ZN(G369));
  NAND3_X1  g0479(.A1(new_n209), .A2(new_n210), .A3(G13), .ZN(new_n680));
  OR2_X1    g0480(.A1(new_n680), .A2(KEYINPUT27), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n680), .A2(KEYINPUT27), .ZN(new_n682));
  NAND3_X1  g0482(.A1(new_n681), .A2(G213), .A3(new_n682), .ZN(new_n683));
  INV_X1    g0483(.A(G343), .ZN(new_n684));
  NOR2_X1   g0484(.A1(new_n683), .A2(new_n684), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n331), .A2(new_n685), .ZN(new_n686));
  MUX2_X1   g0486(.A(new_n658), .B(new_n342), .S(new_n686), .Z(new_n687));
  NAND2_X1  g0487(.A1(new_n687), .A2(G330), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n584), .A2(new_n586), .ZN(new_n689));
  INV_X1    g0489(.A(new_n566), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  INV_X1    g0491(.A(new_n685), .ZN(new_n692));
  OAI21_X1  g0492(.A(new_n579), .B1(new_n566), .B2(new_n692), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n691), .A2(new_n693), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n587), .A2(new_n692), .ZN(new_n695));
  AND2_X1   g0495(.A1(new_n694), .A2(new_n695), .ZN(new_n696));
  INV_X1    g0496(.A(new_n696), .ZN(new_n697));
  NOR2_X1   g0497(.A1(new_n688), .A2(new_n697), .ZN(new_n698));
  AOI21_X1  g0498(.A(new_n685), .B1(new_n329), .B2(new_n341), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n696), .A2(new_n699), .ZN(new_n700));
  NAND2_X1  g0500(.A1(new_n700), .A2(new_n695), .ZN(new_n701));
  OR2_X1    g0501(.A1(new_n698), .A2(new_n701), .ZN(G399));
  INV_X1    g0502(.A(new_n213), .ZN(new_n703));
  NOR2_X1   g0503(.A1(new_n703), .A2(G41), .ZN(new_n704));
  INV_X1    g0504(.A(new_n704), .ZN(new_n705));
  NAND2_X1  g0505(.A1(new_n705), .A2(G1), .ZN(new_n706));
  OR2_X1    g0506(.A1(new_n604), .A2(G116), .ZN(new_n707));
  OAI22_X1  g0507(.A1(new_n706), .A2(new_n707), .B1(new_n229), .B2(new_n705), .ZN(new_n708));
  XNOR2_X1  g0508(.A(new_n708), .B(KEYINPUT28), .ZN(new_n709));
  INV_X1    g0509(.A(G330), .ZN(new_n710));
  NAND4_X1  g0510(.A1(new_n582), .A2(new_n635), .A3(new_n530), .A4(new_n515), .ZN(new_n711));
  OAI21_X1  g0511(.A(new_n338), .B1(new_n325), .B2(new_n271), .ZN(new_n712));
  OAI21_X1  g0512(.A(KEYINPUT89), .B1(new_n711), .B2(new_n712), .ZN(new_n713));
  NAND2_X1  g0513(.A1(new_n713), .A2(KEYINPUT30), .ZN(new_n714));
  INV_X1    g0514(.A(KEYINPUT90), .ZN(new_n715));
  NAND2_X1  g0515(.A1(new_n654), .A2(new_n715), .ZN(new_n716));
  AOI21_X1  g0516(.A(G179), .B1(new_n530), .B2(new_n515), .ZN(new_n717));
  AND2_X1   g0517(.A1(new_n717), .A2(new_n577), .ZN(new_n718));
  OAI211_X1 g0518(.A(KEYINPUT90), .B(new_n595), .C1(new_n652), .C2(new_n653), .ZN(new_n719));
  NAND4_X1  g0519(.A1(new_n716), .A2(new_n718), .A3(new_n326), .A4(new_n719), .ZN(new_n720));
  INV_X1    g0520(.A(KEYINPUT30), .ZN(new_n721));
  OAI211_X1 g0521(.A(KEYINPUT89), .B(new_n721), .C1(new_n711), .C2(new_n712), .ZN(new_n722));
  NAND3_X1  g0522(.A1(new_n714), .A2(new_n720), .A3(new_n722), .ZN(new_n723));
  AND3_X1   g0523(.A1(new_n723), .A2(KEYINPUT31), .A3(new_n685), .ZN(new_n724));
  AOI21_X1  g0524(.A(KEYINPUT31), .B1(new_n723), .B2(new_n685), .ZN(new_n725));
  NOR2_X1   g0525(.A1(new_n724), .A2(new_n725), .ZN(new_n726));
  NAND4_X1  g0526(.A1(new_n639), .A2(new_n342), .A3(new_n580), .A4(new_n692), .ZN(new_n727));
  AOI21_X1  g0527(.A(new_n710), .B1(new_n726), .B2(new_n727), .ZN(new_n728));
  NAND3_X1  g0528(.A1(new_n691), .A2(new_n329), .A3(new_n341), .ZN(new_n729));
  INV_X1    g0529(.A(new_n667), .ZN(new_n730));
  NAND2_X1  g0530(.A1(new_n729), .A2(new_n730), .ZN(new_n731));
  NAND4_X1  g0531(.A1(new_n625), .A2(new_n676), .A3(new_n669), .A4(new_n637), .ZN(new_n732));
  NAND2_X1  g0532(.A1(new_n732), .A2(new_n657), .ZN(new_n733));
  AOI21_X1  g0533(.A(new_n733), .B1(KEYINPUT26), .B2(new_n675), .ZN(new_n734));
  INV_X1    g0534(.A(KEYINPUT91), .ZN(new_n735));
  OAI21_X1  g0535(.A(new_n731), .B1(new_n734), .B2(new_n735), .ZN(new_n736));
  NAND2_X1  g0536(.A1(new_n664), .A2(new_n665), .ZN(new_n737));
  NAND3_X1  g0537(.A1(new_n737), .A2(new_n657), .A3(new_n542), .ZN(new_n738));
  NAND2_X1  g0538(.A1(new_n673), .A2(new_n674), .ZN(new_n739));
  OAI21_X1  g0539(.A(KEYINPUT26), .B1(new_n738), .B2(new_n739), .ZN(new_n740));
  AND2_X1   g0540(.A1(new_n732), .A2(new_n657), .ZN(new_n741));
  NAND2_X1  g0541(.A1(new_n740), .A2(new_n741), .ZN(new_n742));
  NOR2_X1   g0542(.A1(new_n742), .A2(KEYINPUT91), .ZN(new_n743));
  OAI211_X1 g0543(.A(KEYINPUT29), .B(new_n692), .C1(new_n736), .C2(new_n743), .ZN(new_n744));
  OAI21_X1  g0544(.A(new_n692), .B1(new_n668), .B2(new_n677), .ZN(new_n745));
  INV_X1    g0545(.A(KEYINPUT29), .ZN(new_n746));
  NAND2_X1  g0546(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  AOI21_X1  g0547(.A(new_n728), .B1(new_n744), .B2(new_n747), .ZN(new_n748));
  OAI21_X1  g0548(.A(new_n709), .B1(new_n748), .B2(G1), .ZN(G364));
  AOI21_X1  g0549(.A(new_n230), .B1(G20), .B2(new_n253), .ZN(new_n750));
  INV_X1    g0550(.A(new_n750), .ZN(new_n751));
  NOR2_X1   g0551(.A1(new_n210), .A2(G179), .ZN(new_n752));
  NAND3_X1  g0552(.A1(new_n752), .A2(new_n333), .A3(new_n372), .ZN(new_n753));
  OAI21_X1  g0553(.A(KEYINPUT32), .B1(new_n753), .B2(new_n447), .ZN(new_n754));
  NAND2_X1  g0554(.A1(new_n601), .A2(new_n603), .ZN(new_n755));
  INV_X1    g0555(.A(new_n755), .ZN(new_n756));
  NAND3_X1  g0556(.A1(new_n752), .A2(G190), .A3(G200), .ZN(new_n757));
  OAI21_X1  g0557(.A(new_n754), .B1(new_n756), .B2(new_n757), .ZN(new_n758));
  NAND2_X1  g0558(.A1(G20), .A2(G179), .ZN(new_n759));
  NOR3_X1   g0559(.A1(new_n759), .A2(new_n372), .A3(G190), .ZN(new_n760));
  AOI21_X1  g0560(.A(new_n758), .B1(G68), .B2(new_n760), .ZN(new_n761));
  NOR3_X1   g0561(.A1(new_n753), .A2(KEYINPUT32), .A3(new_n447), .ZN(new_n762));
  NOR3_X1   g0562(.A1(new_n333), .A2(G179), .A3(G200), .ZN(new_n763));
  NOR2_X1   g0563(.A1(new_n763), .A2(new_n210), .ZN(new_n764));
  NOR2_X1   g0564(.A1(new_n764), .A2(new_n205), .ZN(new_n765));
  NAND3_X1  g0565(.A1(new_n752), .A2(new_n333), .A3(G200), .ZN(new_n766));
  NOR2_X1   g0566(.A1(new_n766), .A2(new_n206), .ZN(new_n767));
  NOR4_X1   g0567(.A1(new_n762), .A2(new_n765), .A3(new_n767), .A4(new_n294), .ZN(new_n768));
  AOI21_X1  g0568(.A(G200), .B1(new_n759), .B2(KEYINPUT94), .ZN(new_n769));
  OAI21_X1  g0569(.A(new_n769), .B1(KEYINPUT94), .B2(new_n759), .ZN(new_n770));
  NOR2_X1   g0570(.A1(new_n770), .A2(G190), .ZN(new_n771));
  NAND2_X1  g0571(.A1(new_n771), .A2(G77), .ZN(new_n772));
  NAND4_X1  g0572(.A1(G20), .A2(G179), .A3(G190), .A4(G200), .ZN(new_n773));
  NAND2_X1  g0573(.A1(new_n773), .A2(KEYINPUT95), .ZN(new_n774));
  INV_X1    g0574(.A(new_n774), .ZN(new_n775));
  NOR2_X1   g0575(.A1(new_n773), .A2(KEYINPUT95), .ZN(new_n776));
  NOR2_X1   g0576(.A1(new_n775), .A2(new_n776), .ZN(new_n777));
  INV_X1    g0577(.A(new_n777), .ZN(new_n778));
  NOR2_X1   g0578(.A1(new_n770), .A2(new_n333), .ZN(new_n779));
  AOI22_X1  g0579(.A1(new_n778), .A2(G50), .B1(new_n779), .B2(G58), .ZN(new_n780));
  NAND4_X1  g0580(.A1(new_n761), .A2(new_n768), .A3(new_n772), .A4(new_n780), .ZN(new_n781));
  INV_X1    g0581(.A(G303), .ZN(new_n782));
  NOR2_X1   g0582(.A1(new_n757), .A2(new_n782), .ZN(new_n783));
  INV_X1    g0583(.A(new_n753), .ZN(new_n784));
  AOI211_X1 g0584(.A(new_n293), .B(new_n783), .C1(G329), .C2(new_n784), .ZN(new_n785));
  AOI22_X1  g0585(.A1(new_n778), .A2(G326), .B1(new_n771), .B2(G311), .ZN(new_n786));
  INV_X1    g0586(.A(new_n760), .ZN(new_n787));
  XOR2_X1   g0587(.A(KEYINPUT33), .B(G317), .Z(new_n788));
  INV_X1    g0588(.A(G283), .ZN(new_n789));
  OAI22_X1  g0589(.A1(new_n787), .A2(new_n788), .B1(new_n766), .B2(new_n789), .ZN(new_n790));
  INV_X1    g0590(.A(new_n764), .ZN(new_n791));
  AOI21_X1  g0591(.A(new_n790), .B1(G294), .B2(new_n791), .ZN(new_n792));
  NAND2_X1  g0592(.A1(new_n779), .A2(G322), .ZN(new_n793));
  NAND4_X1  g0593(.A1(new_n785), .A2(new_n786), .A3(new_n792), .A4(new_n793), .ZN(new_n794));
  AOI21_X1  g0594(.A(new_n751), .B1(new_n781), .B2(new_n794), .ZN(new_n795));
  AND2_X1   g0595(.A1(new_n210), .A2(G13), .ZN(new_n796));
  AOI21_X1  g0596(.A(new_n209), .B1(new_n796), .B2(G45), .ZN(new_n797));
  INV_X1    g0597(.A(new_n797), .ZN(new_n798));
  NOR2_X1   g0598(.A1(new_n704), .A2(new_n798), .ZN(new_n799));
  INV_X1    g0599(.A(new_n799), .ZN(new_n800));
  NOR2_X1   g0600(.A1(new_n251), .A2(new_n302), .ZN(new_n801));
  NOR2_X1   g0601(.A1(new_n703), .A2(new_n290), .ZN(new_n802));
  INV_X1    g0602(.A(new_n802), .ZN(new_n803));
  INV_X1    g0603(.A(new_n229), .ZN(new_n804));
  AOI21_X1  g0604(.A(new_n803), .B1(new_n302), .B2(new_n804), .ZN(new_n805));
  AOI21_X1  g0605(.A(new_n801), .B1(new_n805), .B2(KEYINPUT92), .ZN(new_n806));
  OAI21_X1  g0606(.A(new_n806), .B1(KEYINPUT92), .B2(new_n805), .ZN(new_n807));
  NOR2_X1   g0607(.A1(new_n703), .A2(new_n294), .ZN(new_n808));
  AOI22_X1  g0608(.A1(new_n808), .A2(G355), .B1(new_n552), .B2(new_n703), .ZN(new_n809));
  NAND2_X1  g0609(.A1(new_n807), .A2(new_n809), .ZN(new_n810));
  NOR2_X1   g0610(.A1(G13), .A2(G33), .ZN(new_n811));
  INV_X1    g0611(.A(new_n811), .ZN(new_n812));
  OR3_X1    g0612(.A1(new_n812), .A2(KEYINPUT93), .A3(G20), .ZN(new_n813));
  OAI21_X1  g0613(.A(KEYINPUT93), .B1(new_n812), .B2(G20), .ZN(new_n814));
  NAND2_X1  g0614(.A1(new_n813), .A2(new_n814), .ZN(new_n815));
  NOR2_X1   g0615(.A1(new_n815), .A2(new_n750), .ZN(new_n816));
  AOI211_X1 g0616(.A(new_n795), .B(new_n800), .C1(new_n810), .C2(new_n816), .ZN(new_n817));
  INV_X1    g0617(.A(new_n815), .ZN(new_n818));
  OAI21_X1  g0618(.A(new_n817), .B1(new_n687), .B2(new_n818), .ZN(new_n819));
  NAND2_X1  g0619(.A1(new_n688), .A2(new_n800), .ZN(new_n820));
  NOR2_X1   g0620(.A1(new_n687), .A2(G330), .ZN(new_n821));
  OAI21_X1  g0621(.A(new_n819), .B1(new_n820), .B2(new_n821), .ZN(new_n822));
  XOR2_X1   g0622(.A(new_n822), .B(KEYINPUT96), .Z(G396));
  NAND2_X1  g0623(.A1(new_n645), .A2(new_n692), .ZN(new_n824));
  OAI21_X1  g0624(.A(new_n438), .B1(new_n426), .B2(new_n692), .ZN(new_n825));
  NAND2_X1  g0625(.A1(new_n825), .A2(new_n436), .ZN(new_n826));
  NAND2_X1  g0626(.A1(new_n824), .A2(new_n826), .ZN(new_n827));
  NAND2_X1  g0627(.A1(new_n745), .A2(new_n827), .ZN(new_n828));
  INV_X1    g0628(.A(new_n827), .ZN(new_n829));
  OAI211_X1 g0629(.A(new_n692), .B(new_n829), .C1(new_n668), .C2(new_n677), .ZN(new_n830));
  AOI21_X1  g0630(.A(new_n728), .B1(new_n828), .B2(new_n830), .ZN(new_n831));
  AOI21_X1  g0631(.A(new_n831), .B1(new_n705), .B2(new_n797), .ZN(new_n832));
  NAND3_X1  g0632(.A1(new_n828), .A2(new_n728), .A3(new_n830), .ZN(new_n833));
  NAND2_X1  g0633(.A1(new_n832), .A2(new_n833), .ZN(new_n834));
  AOI211_X1 g0634(.A(new_n293), .B(new_n765), .C1(G311), .C2(new_n784), .ZN(new_n835));
  OAI22_X1  g0635(.A1(new_n787), .A2(new_n789), .B1(new_n757), .B2(new_n206), .ZN(new_n836));
  INV_X1    g0636(.A(G87), .ZN(new_n837));
  NOR2_X1   g0637(.A1(new_n766), .A2(new_n837), .ZN(new_n838));
  NOR2_X1   g0638(.A1(new_n836), .A2(new_n838), .ZN(new_n839));
  NAND2_X1  g0639(.A1(new_n778), .A2(G303), .ZN(new_n840));
  AOI22_X1  g0640(.A1(G116), .A2(new_n771), .B1(new_n779), .B2(G294), .ZN(new_n841));
  NAND4_X1  g0641(.A1(new_n835), .A2(new_n839), .A3(new_n840), .A4(new_n841), .ZN(new_n842));
  AOI22_X1  g0642(.A1(new_n778), .A2(G137), .B1(new_n771), .B2(G159), .ZN(new_n843));
  AOI22_X1  g0643(.A1(new_n779), .A2(G143), .B1(G150), .B2(new_n760), .ZN(new_n844));
  NAND3_X1  g0644(.A1(new_n843), .A2(KEYINPUT34), .A3(new_n844), .ZN(new_n845));
  INV_X1    g0645(.A(new_n290), .ZN(new_n846));
  AOI21_X1  g0646(.A(new_n846), .B1(G132), .B2(new_n784), .ZN(new_n847));
  INV_X1    g0647(.A(new_n757), .ZN(new_n848));
  NAND2_X1  g0648(.A1(new_n848), .A2(G50), .ZN(new_n849));
  NOR2_X1   g0649(.A1(new_n766), .A2(new_n247), .ZN(new_n850));
  AOI21_X1  g0650(.A(new_n850), .B1(G58), .B2(new_n791), .ZN(new_n851));
  NAND4_X1  g0651(.A1(new_n845), .A2(new_n847), .A3(new_n849), .A4(new_n851), .ZN(new_n852));
  AOI21_X1  g0652(.A(KEYINPUT34), .B1(new_n843), .B2(new_n844), .ZN(new_n853));
  OAI21_X1  g0653(.A(new_n842), .B1(new_n852), .B2(new_n853), .ZN(new_n854));
  AOI21_X1  g0654(.A(new_n751), .B1(new_n854), .B2(KEYINPUT97), .ZN(new_n855));
  OAI21_X1  g0655(.A(new_n855), .B1(KEYINPUT97), .B2(new_n854), .ZN(new_n856));
  NOR2_X1   g0656(.A1(new_n750), .A2(new_n811), .ZN(new_n857));
  AOI21_X1  g0657(.A(new_n800), .B1(new_n367), .B2(new_n857), .ZN(new_n858));
  OAI211_X1 g0658(.A(new_n856), .B(new_n858), .C1(new_n812), .C2(new_n829), .ZN(new_n859));
  AND2_X1   g0659(.A1(new_n834), .A2(new_n859), .ZN(new_n860));
  INV_X1    g0660(.A(new_n860), .ZN(G384));
  INV_X1    g0661(.A(new_n537), .ZN(new_n862));
  OR2_X1    g0662(.A1(new_n862), .A2(KEYINPUT35), .ZN(new_n863));
  NAND2_X1  g0663(.A1(new_n862), .A2(KEYINPUT35), .ZN(new_n864));
  NOR3_X1   g0664(.A1(new_n230), .A2(new_n210), .A3(new_n552), .ZN(new_n865));
  NAND3_X1  g0665(.A1(new_n863), .A2(new_n864), .A3(new_n865), .ZN(new_n866));
  XOR2_X1   g0666(.A(new_n866), .B(KEYINPUT36), .Z(new_n867));
  OR3_X1    g0667(.A1(new_n229), .A2(new_n367), .A3(new_n451), .ZN(new_n868));
  AOI211_X1 g0668(.A(new_n209), .B(G13), .C1(new_n868), .C2(new_n246), .ZN(new_n869));
  NOR2_X1   g0669(.A1(new_n867), .A2(new_n869), .ZN(new_n870));
  INV_X1    g0670(.A(KEYINPUT38), .ZN(new_n871));
  INV_X1    g0671(.A(new_n487), .ZN(new_n872));
  AOI21_X1  g0672(.A(new_n486), .B1(new_n479), .B2(new_n483), .ZN(new_n873));
  NOR2_X1   g0673(.A1(new_n872), .A2(new_n873), .ZN(new_n874));
  AOI21_X1  g0674(.A(new_n502), .B1(new_n874), .B2(new_n470), .ZN(new_n875));
  INV_X1    g0675(.A(KEYINPUT37), .ZN(new_n876));
  INV_X1    g0676(.A(new_n683), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n470), .A2(new_n877), .ZN(new_n878));
  NAND4_X1  g0678(.A1(new_n875), .A2(KEYINPUT99), .A3(new_n876), .A4(new_n878), .ZN(new_n879));
  NAND4_X1  g0679(.A1(new_n488), .A2(new_n497), .A3(new_n878), .A4(new_n876), .ZN(new_n880));
  INV_X1    g0680(.A(KEYINPUT99), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n880), .A2(new_n881), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n875), .A2(new_n878), .ZN(new_n883));
  AOI22_X1  g0683(.A1(new_n879), .A2(new_n882), .B1(new_n883), .B2(KEYINPUT37), .ZN(new_n884));
  INV_X1    g0684(.A(new_n878), .ZN(new_n885));
  AND2_X1   g0685(.A1(new_n504), .A2(new_n885), .ZN(new_n886));
  OAI21_X1  g0686(.A(new_n871), .B1(new_n884), .B2(new_n886), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n445), .A2(new_n454), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n888), .A2(new_n456), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n492), .A2(new_n889), .ZN(new_n890));
  AOI21_X1  g0690(.A(new_n683), .B1(new_n890), .B2(new_n469), .ZN(new_n891));
  NOR2_X1   g0691(.A1(new_n891), .A2(new_n502), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n890), .A2(new_n469), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n874), .A2(new_n893), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n892), .A2(new_n894), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n895), .A2(KEYINPUT37), .ZN(new_n896));
  AND2_X1   g0696(.A1(new_n880), .A2(new_n881), .ZN(new_n897));
  NOR2_X1   g0697(.A1(new_n880), .A2(new_n881), .ZN(new_n898));
  OAI21_X1  g0698(.A(new_n896), .B1(new_n897), .B2(new_n898), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n504), .A2(new_n891), .ZN(new_n900));
  NAND3_X1  g0700(.A1(new_n899), .A2(KEYINPUT38), .A3(new_n900), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n887), .A2(new_n901), .ZN(new_n902));
  INV_X1    g0702(.A(KEYINPUT39), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n902), .A2(new_n903), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n510), .A2(KEYINPUT98), .ZN(new_n905));
  INV_X1    g0705(.A(KEYINPUT98), .ZN(new_n906));
  OAI211_X1 g0706(.A(new_n906), .B(new_n392), .C1(new_n508), .C2(new_n509), .ZN(new_n907));
  AND2_X1   g0707(.A1(new_n905), .A2(new_n907), .ZN(new_n908));
  NOR2_X1   g0708(.A1(new_n908), .A2(new_n685), .ZN(new_n909));
  AOI21_X1  g0709(.A(new_n876), .B1(new_n892), .B2(new_n894), .ZN(new_n910));
  AOI21_X1  g0710(.A(new_n910), .B1(new_n879), .B2(new_n882), .ZN(new_n911));
  AND2_X1   g0711(.A1(new_n504), .A2(new_n891), .ZN(new_n912));
  OAI21_X1  g0712(.A(new_n871), .B1(new_n911), .B2(new_n912), .ZN(new_n913));
  NAND3_X1  g0713(.A1(new_n901), .A2(new_n913), .A3(KEYINPUT39), .ZN(new_n914));
  NAND3_X1  g0714(.A1(new_n904), .A2(new_n909), .A3(new_n914), .ZN(new_n915));
  NOR2_X1   g0715(.A1(new_n391), .A2(new_n692), .ZN(new_n916));
  AOI21_X1  g0716(.A(new_n916), .B1(new_n406), .B2(new_n407), .ZN(new_n917));
  NAND3_X1  g0717(.A1(new_n905), .A2(new_n907), .A3(new_n917), .ZN(new_n918));
  NOR2_X1   g0718(.A1(new_n508), .A2(new_n509), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n408), .A2(new_n919), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n920), .A2(new_n916), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n918), .A2(new_n921), .ZN(new_n922));
  INV_X1    g0722(.A(new_n922), .ZN(new_n923));
  AOI21_X1  g0723(.A(new_n923), .B1(new_n830), .B2(new_n824), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n901), .A2(new_n913), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n924), .A2(new_n925), .ZN(new_n926));
  NAND2_X1  g0726(.A1(new_n649), .A2(new_n683), .ZN(new_n927));
  NAND3_X1  g0727(.A1(new_n915), .A2(new_n926), .A3(new_n927), .ZN(new_n928));
  XOR2_X1   g0728(.A(new_n928), .B(KEYINPUT101), .Z(new_n929));
  INV_X1    g0729(.A(KEYINPUT100), .ZN(new_n930));
  AOI21_X1  g0730(.A(new_n512), .B1(new_n745), .B2(new_n746), .ZN(new_n931));
  AOI21_X1  g0731(.A(new_n930), .B1(new_n744), .B2(new_n931), .ZN(new_n932));
  INV_X1    g0732(.A(new_n932), .ZN(new_n933));
  NAND3_X1  g0733(.A1(new_n744), .A2(new_n931), .A3(new_n930), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n933), .A2(new_n934), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n935), .A2(new_n651), .ZN(new_n936));
  XNOR2_X1  g0736(.A(new_n929), .B(new_n936), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n922), .A2(new_n829), .ZN(new_n938));
  AOI21_X1  g0738(.A(new_n938), .B1(new_n726), .B2(new_n727), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n925), .A2(new_n939), .ZN(new_n940));
  INV_X1    g0740(.A(KEYINPUT40), .ZN(new_n941));
  NAND2_X1  g0741(.A1(new_n940), .A2(new_n941), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n723), .A2(new_n685), .ZN(new_n943));
  INV_X1    g0743(.A(KEYINPUT31), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n943), .A2(new_n944), .ZN(new_n945));
  NAND3_X1  g0745(.A1(new_n723), .A2(KEYINPUT31), .A3(new_n685), .ZN(new_n946));
  NAND3_X1  g0746(.A1(new_n727), .A2(new_n945), .A3(new_n946), .ZN(new_n947));
  AOI21_X1  g0747(.A(new_n827), .B1(new_n918), .B2(new_n921), .ZN(new_n948));
  AND3_X1   g0748(.A1(new_n947), .A2(new_n948), .A3(KEYINPUT40), .ZN(new_n949));
  NAND2_X1  g0749(.A1(new_n949), .A2(new_n902), .ZN(new_n950));
  NAND2_X1  g0750(.A1(new_n942), .A2(new_n950), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n513), .A2(new_n947), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n951), .A2(new_n952), .ZN(new_n953));
  AOI22_X1  g0753(.A1(new_n940), .A2(new_n941), .B1(new_n949), .B2(new_n902), .ZN(new_n954));
  NAND3_X1  g0754(.A1(new_n954), .A2(new_n513), .A3(new_n947), .ZN(new_n955));
  NAND3_X1  g0755(.A1(new_n953), .A2(new_n955), .A3(G330), .ZN(new_n956));
  NAND2_X1  g0756(.A1(new_n937), .A2(new_n956), .ZN(new_n957));
  OAI21_X1  g0757(.A(new_n957), .B1(new_n209), .B2(new_n796), .ZN(new_n958));
  NOR2_X1   g0758(.A1(new_n937), .A2(new_n956), .ZN(new_n959));
  OAI21_X1  g0759(.A(new_n870), .B1(new_n958), .B2(new_n959), .ZN(G367));
  OAI21_X1  g0760(.A(new_n666), .B1(new_n633), .B2(new_n692), .ZN(new_n961));
  NAND2_X1  g0761(.A1(new_n632), .A2(new_n685), .ZN(new_n962));
  OAI21_X1  g0762(.A(new_n961), .B1(new_n657), .B2(new_n962), .ZN(new_n963));
  NAND2_X1  g0763(.A1(new_n963), .A2(KEYINPUT43), .ZN(new_n964));
  INV_X1    g0764(.A(KEYINPUT103), .ZN(new_n965));
  NAND2_X1  g0765(.A1(new_n542), .A2(new_n685), .ZN(new_n966));
  NAND2_X1  g0766(.A1(new_n547), .A2(new_n966), .ZN(new_n967));
  INV_X1    g0767(.A(KEYINPUT102), .ZN(new_n968));
  OAI211_X1 g0768(.A(new_n967), .B(new_n968), .C1(new_n739), .C2(new_n966), .ZN(new_n969));
  OR3_X1    g0769(.A1(new_n739), .A2(new_n968), .A3(new_n966), .ZN(new_n970));
  NAND2_X1  g0770(.A1(new_n969), .A2(new_n970), .ZN(new_n971));
  INV_X1    g0771(.A(new_n971), .ZN(new_n972));
  NAND2_X1  g0772(.A1(new_n972), .A2(new_n587), .ZN(new_n973));
  AOI21_X1  g0773(.A(new_n965), .B1(new_n973), .B2(new_n543), .ZN(new_n974));
  INV_X1    g0774(.A(new_n974), .ZN(new_n975));
  NAND3_X1  g0775(.A1(new_n973), .A2(new_n965), .A3(new_n543), .ZN(new_n976));
  NAND3_X1  g0776(.A1(new_n975), .A2(new_n692), .A3(new_n976), .ZN(new_n977));
  INV_X1    g0777(.A(KEYINPUT104), .ZN(new_n978));
  OAI21_X1  g0778(.A(KEYINPUT42), .B1(new_n700), .B2(new_n971), .ZN(new_n979));
  NAND3_X1  g0779(.A1(new_n977), .A2(new_n978), .A3(new_n979), .ZN(new_n980));
  OR3_X1    g0780(.A1(new_n700), .A2(KEYINPUT42), .A3(new_n971), .ZN(new_n981));
  NAND2_X1  g0781(.A1(new_n980), .A2(new_n981), .ZN(new_n982));
  AOI21_X1  g0782(.A(new_n978), .B1(new_n977), .B2(new_n979), .ZN(new_n983));
  OAI21_X1  g0783(.A(new_n964), .B1(new_n982), .B2(new_n983), .ZN(new_n984));
  NOR2_X1   g0784(.A1(new_n963), .A2(KEYINPUT43), .ZN(new_n985));
  OR2_X1    g0785(.A1(new_n984), .A2(new_n985), .ZN(new_n986));
  NAND2_X1  g0786(.A1(new_n984), .A2(new_n985), .ZN(new_n987));
  NAND2_X1  g0787(.A1(new_n986), .A2(new_n987), .ZN(new_n988));
  INV_X1    g0788(.A(new_n698), .ZN(new_n989));
  NOR2_X1   g0789(.A1(new_n989), .A2(new_n971), .ZN(new_n990));
  XNOR2_X1  g0790(.A(new_n990), .B(KEYINPUT105), .ZN(new_n991));
  OR2_X1    g0791(.A1(new_n988), .A2(new_n991), .ZN(new_n992));
  XOR2_X1   g0792(.A(new_n797), .B(KEYINPUT107), .Z(new_n993));
  INV_X1    g0793(.A(new_n748), .ZN(new_n994));
  NAND2_X1  g0794(.A1(new_n701), .A2(new_n971), .ZN(new_n995));
  XOR2_X1   g0795(.A(new_n995), .B(KEYINPUT44), .Z(new_n996));
  NOR2_X1   g0796(.A1(new_n701), .A2(new_n971), .ZN(new_n997));
  XNOR2_X1  g0797(.A(new_n997), .B(KEYINPUT45), .ZN(new_n998));
  AND3_X1   g0798(.A1(new_n996), .A2(new_n989), .A3(new_n998), .ZN(new_n999));
  AOI21_X1  g0799(.A(new_n989), .B1(new_n996), .B2(new_n998), .ZN(new_n1000));
  NOR2_X1   g0800(.A1(new_n999), .A2(new_n1000), .ZN(new_n1001));
  XOR2_X1   g0801(.A(new_n696), .B(new_n699), .Z(new_n1002));
  XNOR2_X1  g0802(.A(new_n1002), .B(new_n688), .ZN(new_n1003));
  AOI21_X1  g0803(.A(new_n994), .B1(new_n1001), .B2(new_n1003), .ZN(new_n1004));
  XOR2_X1   g0804(.A(KEYINPUT106), .B(KEYINPUT41), .Z(new_n1005));
  XNOR2_X1  g0805(.A(new_n704), .B(new_n1005), .ZN(new_n1006));
  OAI21_X1  g0806(.A(new_n993), .B1(new_n1004), .B2(new_n1006), .ZN(new_n1007));
  NAND2_X1  g0807(.A1(new_n988), .A2(new_n991), .ZN(new_n1008));
  NAND3_X1  g0808(.A1(new_n992), .A2(new_n1007), .A3(new_n1008), .ZN(new_n1009));
  NOR2_X1   g0809(.A1(new_n803), .A2(new_n239), .ZN(new_n1010));
  OAI21_X1  g0810(.A(new_n816), .B1(new_n213), .B2(new_n422), .ZN(new_n1011));
  OAI21_X1  g0811(.A(new_n799), .B1(new_n1010), .B2(new_n1011), .ZN(new_n1012));
  AOI22_X1  g0812(.A1(new_n791), .A2(G107), .B1(G294), .B2(new_n760), .ZN(new_n1013));
  INV_X1    g0813(.A(new_n766), .ZN(new_n1014));
  NAND2_X1  g0814(.A1(new_n1014), .A2(G97), .ZN(new_n1015));
  INV_X1    g0815(.A(new_n779), .ZN(new_n1016));
  OAI211_X1 g0816(.A(new_n1013), .B(new_n1015), .C1(new_n1016), .C2(new_n782), .ZN(new_n1017));
  INV_X1    g0817(.A(new_n771), .ZN(new_n1018));
  INV_X1    g0818(.A(G311), .ZN(new_n1019));
  OAI22_X1  g0819(.A1(new_n1018), .A2(new_n789), .B1(new_n1019), .B2(new_n777), .ZN(new_n1020));
  NOR2_X1   g0820(.A1(new_n1017), .A2(new_n1020), .ZN(new_n1021));
  NAND3_X1  g0821(.A1(new_n848), .A2(KEYINPUT46), .A3(G116), .ZN(new_n1022));
  INV_X1    g0822(.A(KEYINPUT46), .ZN(new_n1023));
  OAI21_X1  g0823(.A(new_n1023), .B1(new_n757), .B2(new_n552), .ZN(new_n1024));
  AOI21_X1  g0824(.A(new_n290), .B1(G317), .B2(new_n784), .ZN(new_n1025));
  NAND4_X1  g0825(.A1(new_n1021), .A2(new_n1022), .A3(new_n1024), .A4(new_n1025), .ZN(new_n1026));
  NAND2_X1  g0826(.A1(new_n778), .A2(G143), .ZN(new_n1027));
  NAND2_X1  g0827(.A1(new_n1014), .A2(G77), .ZN(new_n1028));
  AOI22_X1  g0828(.A1(new_n791), .A2(G68), .B1(G159), .B2(new_n760), .ZN(new_n1029));
  NAND4_X1  g0829(.A1(new_n1027), .A2(new_n293), .A3(new_n1028), .A4(new_n1029), .ZN(new_n1030));
  XNOR2_X1  g0830(.A(KEYINPUT108), .B(G137), .ZN(new_n1031));
  OAI22_X1  g0831(.A1(new_n416), .A2(new_n757), .B1(new_n753), .B2(new_n1031), .ZN(new_n1032));
  INV_X1    g0832(.A(KEYINPUT109), .ZN(new_n1033));
  AOI22_X1  g0833(.A1(G50), .A2(new_n771), .B1(new_n1032), .B2(new_n1033), .ZN(new_n1034));
  OAI221_X1 g0834(.A(new_n1034), .B1(new_n1033), .B2(new_n1032), .C1(new_n346), .C2(new_n1016), .ZN(new_n1035));
  OAI21_X1  g0835(.A(new_n1026), .B1(new_n1030), .B2(new_n1035), .ZN(new_n1036));
  XNOR2_X1  g0836(.A(new_n1036), .B(KEYINPUT47), .ZN(new_n1037));
  AOI21_X1  g0837(.A(new_n1012), .B1(new_n1037), .B2(new_n750), .ZN(new_n1038));
  OAI21_X1  g0838(.A(new_n1038), .B1(new_n963), .B2(new_n818), .ZN(new_n1039));
  NAND2_X1  g0839(.A1(new_n1009), .A2(new_n1039), .ZN(G387));
  INV_X1    g0840(.A(new_n993), .ZN(new_n1041));
  NAND2_X1  g0841(.A1(new_n1003), .A2(new_n1041), .ZN(new_n1042));
  AOI22_X1  g0842(.A1(new_n808), .A2(new_n707), .B1(new_n206), .B2(new_n703), .ZN(new_n1043));
  XOR2_X1   g0843(.A(new_n707), .B(KEYINPUT110), .Z(new_n1044));
  OR3_X1    g0844(.A1(new_n343), .A2(KEYINPUT50), .A3(G50), .ZN(new_n1045));
  OAI21_X1  g0845(.A(KEYINPUT50), .B1(new_n343), .B2(G50), .ZN(new_n1046));
  AOI21_X1  g0846(.A(G45), .B1(G68), .B2(G77), .ZN(new_n1047));
  NAND3_X1  g0847(.A1(new_n1045), .A2(new_n1046), .A3(new_n1047), .ZN(new_n1048));
  OAI21_X1  g0848(.A(new_n802), .B1(new_n1044), .B2(new_n1048), .ZN(new_n1049));
  INV_X1    g0849(.A(KEYINPUT111), .ZN(new_n1050));
  OAI22_X1  g0850(.A1(new_n1049), .A2(new_n1050), .B1(new_n302), .B2(new_n236), .ZN(new_n1051));
  AND2_X1   g0851(.A1(new_n1049), .A2(new_n1050), .ZN(new_n1052));
  OAI21_X1  g0852(.A(new_n1043), .B1(new_n1051), .B2(new_n1052), .ZN(new_n1053));
  AOI21_X1  g0853(.A(new_n800), .B1(new_n1053), .B2(new_n816), .ZN(new_n1054));
  OAI22_X1  g0854(.A1(new_n1018), .A2(new_n247), .B1(new_n447), .B2(new_n777), .ZN(new_n1055));
  AOI21_X1  g0855(.A(new_n846), .B1(G150), .B2(new_n784), .ZN(new_n1056));
  AOI22_X1  g0856(.A1(new_n791), .A2(new_n423), .B1(new_n420), .B2(new_n760), .ZN(new_n1057));
  NAND2_X1  g0857(.A1(new_n848), .A2(G77), .ZN(new_n1058));
  NAND4_X1  g0858(.A1(new_n1056), .A2(new_n1015), .A3(new_n1057), .A4(new_n1058), .ZN(new_n1059));
  AOI211_X1 g0859(.A(new_n1055), .B(new_n1059), .C1(G50), .C2(new_n779), .ZN(new_n1060));
  AOI22_X1  g0860(.A1(new_n791), .A2(G283), .B1(new_n848), .B2(G294), .ZN(new_n1061));
  AOI22_X1  g0861(.A1(new_n771), .A2(G303), .B1(G311), .B2(new_n760), .ZN(new_n1062));
  INV_X1    g0862(.A(G317), .ZN(new_n1063));
  INV_X1    g0863(.A(G322), .ZN(new_n1064));
  OAI221_X1 g0864(.A(new_n1062), .B1(new_n1063), .B2(new_n1016), .C1(new_n1064), .C2(new_n777), .ZN(new_n1065));
  INV_X1    g0865(.A(KEYINPUT48), .ZN(new_n1066));
  OAI21_X1  g0866(.A(new_n1061), .B1(new_n1065), .B2(new_n1066), .ZN(new_n1067));
  XOR2_X1   g0867(.A(new_n1067), .B(KEYINPUT112), .Z(new_n1068));
  NAND2_X1  g0868(.A1(new_n1065), .A2(new_n1066), .ZN(new_n1069));
  NAND2_X1  g0869(.A1(new_n1068), .A2(new_n1069), .ZN(new_n1070));
  XNOR2_X1  g0870(.A(new_n1070), .B(KEYINPUT49), .ZN(new_n1071));
  NOR2_X1   g0871(.A1(new_n766), .A2(new_n552), .ZN(new_n1072));
  AOI211_X1 g0872(.A(new_n290), .B(new_n1072), .C1(G326), .C2(new_n784), .ZN(new_n1073));
  AOI21_X1  g0873(.A(new_n1060), .B1(new_n1071), .B2(new_n1073), .ZN(new_n1074));
  OAI221_X1 g0874(.A(new_n1054), .B1(new_n696), .B2(new_n818), .C1(new_n1074), .C2(new_n751), .ZN(new_n1075));
  NAND2_X1  g0875(.A1(new_n1003), .A2(new_n748), .ZN(new_n1076));
  NAND2_X1  g0876(.A1(new_n1076), .A2(new_n704), .ZN(new_n1077));
  NOR2_X1   g0877(.A1(new_n1003), .A2(new_n748), .ZN(new_n1078));
  OAI211_X1 g0878(.A(new_n1042), .B(new_n1075), .C1(new_n1077), .C2(new_n1078), .ZN(G393));
  INV_X1    g0879(.A(new_n1001), .ZN(new_n1080));
  NAND2_X1  g0880(.A1(new_n1080), .A2(new_n1076), .ZN(new_n1081));
  INV_X1    g0881(.A(new_n1076), .ZN(new_n1082));
  AOI21_X1  g0882(.A(new_n705), .B1(new_n1001), .B2(new_n1082), .ZN(new_n1083));
  AND2_X1   g0883(.A1(new_n1081), .A2(new_n1083), .ZN(new_n1084));
  OAI221_X1 g0884(.A(new_n816), .B1(new_n205), .B2(new_n213), .C1(new_n245), .C2(new_n803), .ZN(new_n1085));
  INV_X1    g0885(.A(KEYINPUT113), .ZN(new_n1086));
  AOI21_X1  g0886(.A(new_n800), .B1(new_n1085), .B2(new_n1086), .ZN(new_n1087));
  OAI21_X1  g0887(.A(new_n1087), .B1(new_n1086), .B2(new_n1085), .ZN(new_n1088));
  NOR2_X1   g0888(.A1(new_n764), .A2(new_n367), .ZN(new_n1089));
  AOI211_X1 g0889(.A(new_n838), .B(new_n1089), .C1(G68), .C2(new_n848), .ZN(new_n1090));
  AOI21_X1  g0890(.A(new_n846), .B1(G143), .B2(new_n784), .ZN(new_n1091));
  NAND2_X1  g0891(.A1(new_n1090), .A2(new_n1091), .ZN(new_n1092));
  AOI22_X1  g0892(.A1(new_n771), .A2(new_n420), .B1(G50), .B2(new_n760), .ZN(new_n1093));
  AOI21_X1  g0893(.A(new_n1092), .B1(KEYINPUT114), .B2(new_n1093), .ZN(new_n1094));
  OAI21_X1  g0894(.A(new_n1094), .B1(KEYINPUT114), .B2(new_n1093), .ZN(new_n1095));
  AOI22_X1  g0895(.A1(new_n778), .A2(G150), .B1(new_n779), .B2(G159), .ZN(new_n1096));
  XNOR2_X1  g0896(.A(new_n1096), .B(KEYINPUT51), .ZN(new_n1097));
  NOR2_X1   g0897(.A1(new_n1095), .A2(new_n1097), .ZN(new_n1098));
  OR2_X1    g0898(.A1(new_n1098), .A2(KEYINPUT115), .ZN(new_n1099));
  NAND2_X1  g0899(.A1(new_n1098), .A2(KEYINPUT115), .ZN(new_n1100));
  OAI22_X1  g0900(.A1(new_n1016), .A2(new_n1019), .B1(new_n1063), .B2(new_n777), .ZN(new_n1101));
  XNOR2_X1  g0901(.A(new_n1101), .B(KEYINPUT52), .ZN(new_n1102));
  OAI221_X1 g0902(.A(new_n294), .B1(new_n753), .B2(new_n1064), .C1(new_n206), .C2(new_n766), .ZN(new_n1103));
  AOI22_X1  g0903(.A1(new_n848), .A2(G283), .B1(G303), .B2(new_n760), .ZN(new_n1104));
  OAI21_X1  g0904(.A(new_n1104), .B1(new_n552), .B2(new_n764), .ZN(new_n1105));
  AOI211_X1 g0905(.A(new_n1103), .B(new_n1105), .C1(G294), .C2(new_n771), .ZN(new_n1106));
  NAND2_X1  g0906(.A1(new_n1102), .A2(new_n1106), .ZN(new_n1107));
  NAND3_X1  g0907(.A1(new_n1099), .A2(new_n1100), .A3(new_n1107), .ZN(new_n1108));
  AOI21_X1  g0908(.A(new_n1088), .B1(new_n750), .B2(new_n1108), .ZN(new_n1109));
  OAI21_X1  g0909(.A(new_n1109), .B1(new_n972), .B2(new_n818), .ZN(new_n1110));
  OAI21_X1  g0910(.A(new_n1110), .B1(new_n1080), .B2(new_n993), .ZN(new_n1111));
  OR2_X1    g0911(.A1(new_n1084), .A2(new_n1111), .ZN(G390));
  INV_X1    g0912(.A(new_n914), .ZN(new_n1113));
  AOI21_X1  g0913(.A(KEYINPUT39), .B1(new_n887), .B2(new_n901), .ZN(new_n1114));
  OAI21_X1  g0914(.A(new_n811), .B1(new_n1113), .B2(new_n1114), .ZN(new_n1115));
  INV_X1    g0915(.A(new_n857), .ZN(new_n1116));
  OAI21_X1  g0916(.A(new_n799), .B1(new_n420), .B2(new_n1116), .ZN(new_n1117));
  NOR2_X1   g0917(.A1(new_n757), .A2(new_n837), .ZN(new_n1118));
  AOI211_X1 g0918(.A(new_n1118), .B(new_n1089), .C1(G107), .C2(new_n760), .ZN(new_n1119));
  AOI211_X1 g0919(.A(new_n293), .B(new_n850), .C1(G294), .C2(new_n784), .ZN(new_n1120));
  NAND2_X1  g0920(.A1(new_n778), .A2(G283), .ZN(new_n1121));
  AOI22_X1  g0921(.A1(G97), .A2(new_n771), .B1(new_n779), .B2(G116), .ZN(new_n1122));
  NAND4_X1  g0922(.A1(new_n1119), .A2(new_n1120), .A3(new_n1121), .A4(new_n1122), .ZN(new_n1123));
  XNOR2_X1  g0923(.A(KEYINPUT54), .B(G143), .ZN(new_n1124));
  INV_X1    g0924(.A(new_n1124), .ZN(new_n1125));
  INV_X1    g0925(.A(new_n1031), .ZN(new_n1126));
  AOI22_X1  g0926(.A1(new_n771), .A2(new_n1125), .B1(new_n760), .B2(new_n1126), .ZN(new_n1127));
  XOR2_X1   g0927(.A(new_n1127), .B(KEYINPUT117), .Z(new_n1128));
  INV_X1    g0928(.A(G125), .ZN(new_n1129));
  OAI221_X1 g0929(.A(new_n293), .B1(new_n753), .B2(new_n1129), .C1(new_n202), .C2(new_n766), .ZN(new_n1130));
  AOI21_X1  g0930(.A(new_n1130), .B1(G159), .B2(new_n791), .ZN(new_n1131));
  NOR2_X1   g0931(.A1(new_n757), .A2(new_n346), .ZN(new_n1132));
  XNOR2_X1  g0932(.A(new_n1132), .B(KEYINPUT53), .ZN(new_n1133));
  AOI22_X1  g0933(.A1(new_n778), .A2(G128), .B1(new_n779), .B2(G132), .ZN(new_n1134));
  NAND3_X1  g0934(.A1(new_n1131), .A2(new_n1133), .A3(new_n1134), .ZN(new_n1135));
  OAI21_X1  g0935(.A(new_n1123), .B1(new_n1128), .B2(new_n1135), .ZN(new_n1136));
  AOI21_X1  g0936(.A(new_n1117), .B1(new_n1136), .B2(new_n750), .ZN(new_n1137));
  NAND2_X1  g0937(.A1(new_n1115), .A2(new_n1137), .ZN(new_n1138));
  NAND4_X1  g0938(.A1(new_n947), .A2(G330), .A3(new_n829), .A4(new_n922), .ZN(new_n1139));
  INV_X1    g0939(.A(new_n1139), .ZN(new_n1140));
  INV_X1    g0940(.A(new_n909), .ZN(new_n1141));
  NAND2_X1  g0941(.A1(new_n902), .A2(new_n1141), .ZN(new_n1142));
  OAI211_X1 g0942(.A(new_n692), .B(new_n826), .C1(new_n736), .C2(new_n743), .ZN(new_n1143));
  NAND2_X1  g0943(.A1(new_n1143), .A2(new_n824), .ZN(new_n1144));
  AOI21_X1  g0944(.A(new_n1142), .B1(new_n1144), .B2(new_n922), .ZN(new_n1145));
  NAND2_X1  g0945(.A1(new_n830), .A2(new_n824), .ZN(new_n1146));
  NAND2_X1  g0946(.A1(new_n1146), .A2(new_n922), .ZN(new_n1147));
  AOI22_X1  g0947(.A1(new_n1147), .A2(new_n1141), .B1(new_n904), .B2(new_n914), .ZN(new_n1148));
  OAI21_X1  g0948(.A(new_n1140), .B1(new_n1145), .B2(new_n1148), .ZN(new_n1149));
  OAI22_X1  g0949(.A1(new_n1113), .A2(new_n1114), .B1(new_n924), .B2(new_n909), .ZN(new_n1150));
  AOI21_X1  g0950(.A(new_n923), .B1(new_n1143), .B2(new_n824), .ZN(new_n1151));
  OAI211_X1 g0951(.A(new_n1150), .B(new_n1139), .C1(new_n1151), .C2(new_n1142), .ZN(new_n1152));
  NAND2_X1  g0952(.A1(new_n1149), .A2(new_n1152), .ZN(new_n1153));
  OAI21_X1  g0953(.A(new_n1138), .B1(new_n1153), .B2(new_n993), .ZN(new_n1154));
  AOI21_X1  g0954(.A(new_n922), .B1(new_n728), .B2(new_n829), .ZN(new_n1155));
  OAI21_X1  g0955(.A(new_n1146), .B1(new_n1155), .B2(new_n1140), .ZN(new_n1156));
  NAND3_X1  g0956(.A1(new_n947), .A2(G330), .A3(new_n829), .ZN(new_n1157));
  NAND2_X1  g0957(.A1(new_n1157), .A2(new_n923), .ZN(new_n1158));
  NAND2_X1  g0958(.A1(new_n1158), .A2(new_n1139), .ZN(new_n1159));
  OAI21_X1  g0959(.A(new_n1156), .B1(new_n1144), .B2(new_n1159), .ZN(new_n1160));
  NAND2_X1  g0960(.A1(new_n728), .A2(new_n513), .ZN(new_n1161));
  NAND4_X1  g0961(.A1(new_n1160), .A2(new_n935), .A3(new_n651), .A4(new_n1161), .ZN(new_n1162));
  NAND2_X1  g0962(.A1(new_n1153), .A2(new_n1162), .ZN(new_n1163));
  AND3_X1   g0963(.A1(new_n744), .A2(new_n930), .A3(new_n931), .ZN(new_n1164));
  OAI211_X1 g0964(.A(new_n651), .B(new_n1161), .C1(new_n1164), .C2(new_n932), .ZN(new_n1165));
  INV_X1    g0965(.A(new_n1165), .ZN(new_n1166));
  NAND4_X1  g0966(.A1(new_n1166), .A2(new_n1149), .A3(new_n1152), .A4(new_n1160), .ZN(new_n1167));
  NAND3_X1  g0967(.A1(new_n1163), .A2(new_n1167), .A3(new_n704), .ZN(new_n1168));
  INV_X1    g0968(.A(KEYINPUT116), .ZN(new_n1169));
  NAND2_X1  g0969(.A1(new_n1168), .A2(new_n1169), .ZN(new_n1170));
  AOI21_X1  g0970(.A(new_n705), .B1(new_n1153), .B2(new_n1162), .ZN(new_n1171));
  NAND3_X1  g0971(.A1(new_n1171), .A2(KEYINPUT116), .A3(new_n1167), .ZN(new_n1172));
  AOI21_X1  g0972(.A(new_n1154), .B1(new_n1170), .B2(new_n1172), .ZN(new_n1173));
  INV_X1    g0973(.A(new_n1173), .ZN(G378));
  AOI22_X1  g0974(.A1(new_n1158), .A2(new_n1139), .B1(new_n824), .B2(new_n830), .ZN(new_n1175));
  INV_X1    g0975(.A(new_n1144), .ZN(new_n1176));
  NOR2_X1   g0976(.A1(new_n1155), .A2(new_n1140), .ZN(new_n1177));
  AOI21_X1  g0977(.A(new_n1175), .B1(new_n1176), .B2(new_n1177), .ZN(new_n1178));
  OAI21_X1  g0978(.A(new_n1166), .B1(new_n1153), .B2(new_n1178), .ZN(new_n1179));
  NAND2_X1  g0979(.A1(new_n644), .A2(new_n413), .ZN(new_n1180));
  NOR2_X1   g0980(.A1(new_n352), .A2(new_n357), .ZN(new_n1181));
  NOR2_X1   g0981(.A1(new_n1181), .A2(new_n683), .ZN(new_n1182));
  NAND2_X1  g0982(.A1(new_n1180), .A2(new_n1182), .ZN(new_n1183));
  INV_X1    g0983(.A(new_n1182), .ZN(new_n1184));
  OAI211_X1 g0984(.A(new_n413), .B(new_n1184), .C1(new_n642), .C2(new_n643), .ZN(new_n1185));
  XNOR2_X1  g0985(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1186));
  NAND3_X1  g0986(.A1(new_n1183), .A2(new_n1185), .A3(new_n1186), .ZN(new_n1187));
  INV_X1    g0987(.A(new_n1186), .ZN(new_n1188));
  AOI21_X1  g0988(.A(new_n1184), .B1(new_n644), .B2(new_n413), .ZN(new_n1189));
  INV_X1    g0989(.A(new_n1185), .ZN(new_n1190));
  OAI21_X1  g0990(.A(new_n1188), .B1(new_n1189), .B2(new_n1190), .ZN(new_n1191));
  NAND2_X1  g0991(.A1(new_n1187), .A2(new_n1191), .ZN(new_n1192));
  AND3_X1   g0992(.A1(new_n954), .A2(G330), .A3(new_n1192), .ZN(new_n1193));
  AOI21_X1  g0993(.A(new_n1192), .B1(new_n954), .B2(G330), .ZN(new_n1194));
  OAI21_X1  g0994(.A(new_n928), .B1(new_n1193), .B2(new_n1194), .ZN(new_n1195));
  INV_X1    g0995(.A(new_n1192), .ZN(new_n1196));
  OAI21_X1  g0996(.A(new_n1196), .B1(new_n951), .B2(new_n710), .ZN(new_n1197));
  INV_X1    g0997(.A(new_n928), .ZN(new_n1198));
  NAND3_X1  g0998(.A1(new_n954), .A2(G330), .A3(new_n1192), .ZN(new_n1199));
  NAND3_X1  g0999(.A1(new_n1197), .A2(new_n1198), .A3(new_n1199), .ZN(new_n1200));
  INV_X1    g1000(.A(KEYINPUT119), .ZN(new_n1201));
  NAND3_X1  g1001(.A1(new_n1195), .A2(new_n1200), .A3(new_n1201), .ZN(new_n1202));
  NAND4_X1  g1002(.A1(new_n1197), .A2(new_n1198), .A3(KEYINPUT119), .A4(new_n1199), .ZN(new_n1203));
  NAND3_X1  g1003(.A1(new_n1179), .A2(new_n1202), .A3(new_n1203), .ZN(new_n1204));
  INV_X1    g1004(.A(KEYINPUT57), .ZN(new_n1205));
  NAND2_X1  g1005(.A1(new_n1204), .A2(new_n1205), .ZN(new_n1206));
  NAND2_X1  g1006(.A1(new_n1206), .A2(KEYINPUT120), .ZN(new_n1207));
  INV_X1    g1007(.A(KEYINPUT120), .ZN(new_n1208));
  NAND3_X1  g1008(.A1(new_n1204), .A2(new_n1208), .A3(new_n1205), .ZN(new_n1209));
  AOI21_X1  g1009(.A(new_n1205), .B1(new_n1195), .B2(new_n1200), .ZN(new_n1210));
  NAND2_X1  g1010(.A1(new_n1210), .A2(new_n1179), .ZN(new_n1211));
  NAND2_X1  g1011(.A1(new_n1211), .A2(new_n704), .ZN(new_n1212));
  INV_X1    g1012(.A(new_n1212), .ZN(new_n1213));
  NAND3_X1  g1013(.A1(new_n1207), .A2(new_n1209), .A3(new_n1213), .ZN(new_n1214));
  NAND3_X1  g1014(.A1(new_n1202), .A2(new_n1041), .A3(new_n1203), .ZN(new_n1215));
  NAND2_X1  g1015(.A1(new_n1196), .A2(new_n811), .ZN(new_n1216));
  AOI22_X1  g1016(.A1(new_n778), .A2(G116), .B1(new_n779), .B2(G107), .ZN(new_n1217));
  OAI21_X1  g1017(.A(new_n1217), .B1(new_n422), .B2(new_n1018), .ZN(new_n1218));
  OAI211_X1 g1018(.A(new_n846), .B(new_n298), .C1(new_n789), .C2(new_n753), .ZN(new_n1219));
  AOI22_X1  g1019(.A1(new_n1014), .A2(G58), .B1(new_n760), .B2(G97), .ZN(new_n1220));
  OAI211_X1 g1020(.A(new_n1220), .B(new_n1058), .C1(new_n247), .C2(new_n764), .ZN(new_n1221));
  NOR3_X1   g1021(.A1(new_n1218), .A2(new_n1219), .A3(new_n1221), .ZN(new_n1222));
  XNOR2_X1  g1022(.A(KEYINPUT118), .B(KEYINPUT58), .ZN(new_n1223));
  INV_X1    g1023(.A(new_n1223), .ZN(new_n1224));
  NAND2_X1  g1024(.A1(new_n1222), .A2(new_n1224), .ZN(new_n1225));
  OAI21_X1  g1025(.A(new_n298), .B1(new_n284), .B2(new_n275), .ZN(new_n1226));
  NAND2_X1  g1026(.A1(new_n1226), .A2(new_n202), .ZN(new_n1227));
  AND2_X1   g1027(.A1(new_n1225), .A2(new_n1227), .ZN(new_n1228));
  INV_X1    g1028(.A(G128), .ZN(new_n1229));
  OAI22_X1  g1029(.A1(new_n1016), .A2(new_n1229), .B1(new_n1129), .B2(new_n777), .ZN(new_n1230));
  NAND2_X1  g1030(.A1(new_n791), .A2(G150), .ZN(new_n1231));
  NAND2_X1  g1031(.A1(new_n848), .A2(new_n1125), .ZN(new_n1232));
  NAND2_X1  g1032(.A1(new_n760), .A2(G132), .ZN(new_n1233));
  NAND3_X1  g1033(.A1(new_n1231), .A2(new_n1232), .A3(new_n1233), .ZN(new_n1234));
  AOI211_X1 g1034(.A(new_n1230), .B(new_n1234), .C1(G137), .C2(new_n771), .ZN(new_n1235));
  INV_X1    g1035(.A(new_n1235), .ZN(new_n1236));
  NAND2_X1  g1036(.A1(new_n1236), .A2(KEYINPUT59), .ZN(new_n1237));
  NAND2_X1  g1037(.A1(new_n1014), .A2(G159), .ZN(new_n1238));
  AOI211_X1 g1038(.A(G33), .B(G41), .C1(new_n784), .C2(G124), .ZN(new_n1239));
  NAND3_X1  g1039(.A1(new_n1237), .A2(new_n1238), .A3(new_n1239), .ZN(new_n1240));
  NOR2_X1   g1040(.A1(new_n1236), .A2(KEYINPUT59), .ZN(new_n1241));
  OAI221_X1 g1041(.A(new_n1228), .B1(new_n1224), .B2(new_n1222), .C1(new_n1240), .C2(new_n1241), .ZN(new_n1242));
  NAND2_X1  g1042(.A1(new_n1242), .A2(new_n750), .ZN(new_n1243));
  AOI21_X1  g1043(.A(new_n800), .B1(new_n202), .B2(new_n857), .ZN(new_n1244));
  NAND3_X1  g1044(.A1(new_n1216), .A2(new_n1243), .A3(new_n1244), .ZN(new_n1245));
  NAND2_X1  g1045(.A1(new_n1215), .A2(new_n1245), .ZN(new_n1246));
  INV_X1    g1046(.A(new_n1246), .ZN(new_n1247));
  NAND2_X1  g1047(.A1(new_n1214), .A2(new_n1247), .ZN(G375));
  INV_X1    g1048(.A(new_n1162), .ZN(new_n1249));
  NOR2_X1   g1049(.A1(new_n1249), .A2(new_n1006), .ZN(new_n1250));
  NAND2_X1  g1050(.A1(new_n1165), .A2(new_n1178), .ZN(new_n1251));
  NAND2_X1  g1051(.A1(new_n1250), .A2(new_n1251), .ZN(new_n1252));
  NAND2_X1  g1052(.A1(new_n923), .A2(new_n811), .ZN(new_n1253));
  OAI21_X1  g1053(.A(new_n799), .B1(G68), .B2(new_n1116), .ZN(new_n1254));
  OAI21_X1  g1054(.A(new_n290), .B1(new_n416), .B2(new_n766), .ZN(new_n1255));
  INV_X1    g1055(.A(KEYINPUT121), .ZN(new_n1256));
  AOI22_X1  g1056(.A1(new_n1255), .A2(new_n1256), .B1(new_n779), .B2(new_n1126), .ZN(new_n1257));
  INV_X1    g1057(.A(KEYINPUT122), .ZN(new_n1258));
  OAI22_X1  g1058(.A1(new_n753), .A2(new_n1229), .B1(new_n757), .B2(new_n447), .ZN(new_n1259));
  OAI221_X1 g1059(.A(new_n1257), .B1(new_n1258), .B2(new_n1259), .C1(new_n346), .C2(new_n1018), .ZN(new_n1260));
  AOI22_X1  g1060(.A1(new_n778), .A2(G132), .B1(new_n1259), .B2(new_n1258), .ZN(new_n1261));
  AOI22_X1  g1061(.A1(new_n791), .A2(G50), .B1(new_n760), .B2(new_n1125), .ZN(new_n1262));
  OAI211_X1 g1062(.A(new_n1261), .B(new_n1262), .C1(new_n1256), .C2(new_n1255), .ZN(new_n1263));
  AOI22_X1  g1063(.A1(new_n791), .A2(new_n423), .B1(G116), .B2(new_n760), .ZN(new_n1264));
  AOI21_X1  g1064(.A(new_n293), .B1(new_n784), .B2(G303), .ZN(new_n1265));
  NAND2_X1  g1065(.A1(new_n848), .A2(G97), .ZN(new_n1266));
  NAND4_X1  g1066(.A1(new_n1264), .A2(new_n1028), .A3(new_n1265), .A4(new_n1266), .ZN(new_n1267));
  AOI22_X1  g1067(.A1(new_n778), .A2(G294), .B1(new_n771), .B2(G107), .ZN(new_n1268));
  OAI21_X1  g1068(.A(new_n1268), .B1(new_n789), .B2(new_n1016), .ZN(new_n1269));
  OAI22_X1  g1069(.A1(new_n1260), .A2(new_n1263), .B1(new_n1267), .B2(new_n1269), .ZN(new_n1270));
  AOI21_X1  g1070(.A(new_n1254), .B1(new_n1270), .B2(new_n750), .ZN(new_n1271));
  AOI22_X1  g1071(.A1(new_n1160), .A2(new_n1041), .B1(new_n1253), .B2(new_n1271), .ZN(new_n1272));
  NAND2_X1  g1072(.A1(new_n1252), .A2(new_n1272), .ZN(G381));
  NOR2_X1   g1073(.A1(new_n1084), .A2(new_n1111), .ZN(new_n1274));
  NAND2_X1  g1074(.A1(new_n1274), .A2(new_n860), .ZN(new_n1275));
  OR4_X1    g1075(.A1(G396), .A2(new_n1275), .A3(G393), .A4(G381), .ZN(new_n1276));
  AOI21_X1  g1076(.A(new_n1154), .B1(new_n1167), .B2(new_n1171), .ZN(new_n1277));
  INV_X1    g1077(.A(new_n1277), .ZN(new_n1278));
  OR4_X1    g1078(.A1(G387), .A2(new_n1276), .A3(G375), .A4(new_n1278), .ZN(G407));
  INV_X1    g1079(.A(G213), .ZN(new_n1280));
  NOR2_X1   g1080(.A1(new_n1280), .A2(G343), .ZN(new_n1281));
  NAND4_X1  g1081(.A1(new_n1214), .A2(new_n1247), .A3(new_n1277), .A4(new_n1281), .ZN(new_n1282));
  NAND3_X1  g1082(.A1(G407), .A2(G213), .A3(new_n1282), .ZN(G409));
  XOR2_X1   g1083(.A(G393), .B(G396), .Z(new_n1284));
  NAND2_X1  g1084(.A1(G390), .A2(new_n1284), .ZN(new_n1285));
  INV_X1    g1085(.A(new_n1284), .ZN(new_n1286));
  NAND2_X1  g1086(.A1(new_n1274), .A2(new_n1286), .ZN(new_n1287));
  NAND2_X1  g1087(.A1(new_n1285), .A2(new_n1287), .ZN(new_n1288));
  NAND2_X1  g1088(.A1(new_n1288), .A2(G387), .ZN(new_n1289));
  NAND4_X1  g1089(.A1(new_n1285), .A2(new_n1039), .A3(new_n1009), .A4(new_n1287), .ZN(new_n1290));
  NAND2_X1  g1090(.A1(new_n1289), .A2(new_n1290), .ZN(new_n1291));
  INV_X1    g1091(.A(KEYINPUT126), .ZN(new_n1292));
  INV_X1    g1092(.A(KEYINPUT61), .ZN(new_n1293));
  NAND3_X1  g1093(.A1(new_n1214), .A2(G378), .A3(new_n1247), .ZN(new_n1294));
  OR2_X1    g1094(.A1(new_n1204), .A2(new_n1006), .ZN(new_n1295));
  INV_X1    g1095(.A(new_n1245), .ZN(new_n1296));
  NAND2_X1  g1096(.A1(new_n1195), .A2(new_n1200), .ZN(new_n1297));
  AOI21_X1  g1097(.A(new_n1296), .B1(new_n1297), .B2(new_n1041), .ZN(new_n1298));
  AOI21_X1  g1098(.A(new_n1278), .B1(new_n1295), .B2(new_n1298), .ZN(new_n1299));
  INV_X1    g1099(.A(new_n1299), .ZN(new_n1300));
  AOI21_X1  g1100(.A(new_n1281), .B1(new_n1294), .B2(new_n1300), .ZN(new_n1301));
  NAND2_X1  g1101(.A1(new_n1281), .A2(G2897), .ZN(new_n1302));
  NAND3_X1  g1102(.A1(new_n1165), .A2(new_n1178), .A3(KEYINPUT60), .ZN(new_n1303));
  NAND2_X1  g1103(.A1(new_n1303), .A2(KEYINPUT123), .ZN(new_n1304));
  AOI21_X1  g1104(.A(new_n705), .B1(new_n1166), .B2(new_n1160), .ZN(new_n1305));
  INV_X1    g1105(.A(KEYINPUT123), .ZN(new_n1306));
  NAND4_X1  g1106(.A1(new_n1165), .A2(new_n1178), .A3(new_n1306), .A4(KEYINPUT60), .ZN(new_n1307));
  INV_X1    g1107(.A(KEYINPUT60), .ZN(new_n1308));
  NAND2_X1  g1108(.A1(new_n1251), .A2(new_n1308), .ZN(new_n1309));
  NAND4_X1  g1109(.A1(new_n1304), .A2(new_n1305), .A3(new_n1307), .A4(new_n1309), .ZN(new_n1310));
  NAND3_X1  g1110(.A1(new_n1310), .A2(G384), .A3(new_n1272), .ZN(new_n1311));
  INV_X1    g1111(.A(new_n1311), .ZN(new_n1312));
  AOI21_X1  g1112(.A(G384), .B1(new_n1310), .B2(new_n1272), .ZN(new_n1313));
  INV_X1    g1113(.A(KEYINPUT125), .ZN(new_n1314));
  NOR3_X1   g1114(.A1(new_n1312), .A2(new_n1313), .A3(new_n1314), .ZN(new_n1315));
  NAND2_X1  g1115(.A1(new_n1310), .A2(new_n1272), .ZN(new_n1316));
  NAND2_X1  g1116(.A1(new_n1316), .A2(new_n860), .ZN(new_n1317));
  AOI21_X1  g1117(.A(KEYINPUT125), .B1(new_n1317), .B2(new_n1311), .ZN(new_n1318));
  OAI21_X1  g1118(.A(new_n1302), .B1(new_n1315), .B2(new_n1318), .ZN(new_n1319));
  NAND3_X1  g1119(.A1(new_n1317), .A2(KEYINPUT125), .A3(new_n1311), .ZN(new_n1320));
  NAND3_X1  g1120(.A1(new_n1320), .A2(G2897), .A3(new_n1281), .ZN(new_n1321));
  NAND2_X1  g1121(.A1(new_n1319), .A2(new_n1321), .ZN(new_n1322));
  OAI211_X1 g1122(.A(new_n1292), .B(new_n1293), .C1(new_n1301), .C2(new_n1322), .ZN(new_n1323));
  INV_X1    g1123(.A(new_n1281), .ZN(new_n1324));
  NOR2_X1   g1124(.A1(new_n1312), .A2(new_n1313), .ZN(new_n1325));
  AOI21_X1  g1125(.A(new_n1212), .B1(new_n1206), .B2(KEYINPUT120), .ZN(new_n1326));
  AOI211_X1 g1126(.A(new_n1246), .B(new_n1173), .C1(new_n1326), .C2(new_n1209), .ZN(new_n1327));
  OAI211_X1 g1127(.A(new_n1324), .B(new_n1325), .C1(new_n1327), .C2(new_n1299), .ZN(new_n1328));
  NAND2_X1  g1128(.A1(new_n1328), .A2(KEYINPUT62), .ZN(new_n1329));
  INV_X1    g1129(.A(KEYINPUT62), .ZN(new_n1330));
  NAND3_X1  g1130(.A1(new_n1301), .A2(new_n1330), .A3(new_n1325), .ZN(new_n1331));
  NAND3_X1  g1131(.A1(new_n1323), .A2(new_n1329), .A3(new_n1331), .ZN(new_n1332));
  OAI21_X1  g1132(.A(new_n1324), .B1(new_n1327), .B2(new_n1299), .ZN(new_n1333));
  OAI21_X1  g1133(.A(new_n1314), .B1(new_n1312), .B2(new_n1313), .ZN(new_n1334));
  AOI22_X1  g1134(.A1(new_n1334), .A2(new_n1320), .B1(G2897), .B2(new_n1281), .ZN(new_n1335));
  NOR2_X1   g1135(.A1(new_n1315), .A2(new_n1302), .ZN(new_n1336));
  NOR2_X1   g1136(.A1(new_n1335), .A2(new_n1336), .ZN(new_n1337));
  NAND2_X1  g1137(.A1(new_n1333), .A2(new_n1337), .ZN(new_n1338));
  AOI21_X1  g1138(.A(new_n1292), .B1(new_n1338), .B2(new_n1293), .ZN(new_n1339));
  OAI21_X1  g1139(.A(new_n1291), .B1(new_n1332), .B2(new_n1339), .ZN(new_n1340));
  NAND2_X1  g1140(.A1(new_n1333), .A2(KEYINPUT124), .ZN(new_n1341));
  INV_X1    g1141(.A(KEYINPUT124), .ZN(new_n1342));
  NAND2_X1  g1142(.A1(new_n1301), .A2(new_n1342), .ZN(new_n1343));
  NAND3_X1  g1143(.A1(new_n1341), .A2(new_n1343), .A3(new_n1337), .ZN(new_n1344));
  NOR2_X1   g1144(.A1(new_n1291), .A2(KEYINPUT61), .ZN(new_n1345));
  INV_X1    g1145(.A(KEYINPUT63), .ZN(new_n1346));
  NAND2_X1  g1146(.A1(new_n1328), .A2(new_n1346), .ZN(new_n1347));
  NAND3_X1  g1147(.A1(new_n1301), .A2(KEYINPUT63), .A3(new_n1325), .ZN(new_n1348));
  NAND4_X1  g1148(.A1(new_n1344), .A2(new_n1345), .A3(new_n1347), .A4(new_n1348), .ZN(new_n1349));
  NAND2_X1  g1149(.A1(new_n1340), .A2(new_n1349), .ZN(G405));
  NAND2_X1  g1150(.A1(G375), .A2(new_n1277), .ZN(new_n1351));
  NAND2_X1  g1151(.A1(new_n1325), .A2(KEYINPUT127), .ZN(new_n1352));
  NAND3_X1  g1152(.A1(new_n1351), .A2(new_n1294), .A3(new_n1352), .ZN(new_n1353));
  INV_X1    g1153(.A(KEYINPUT127), .ZN(new_n1354));
  INV_X1    g1154(.A(new_n1325), .ZN(new_n1355));
  NAND3_X1  g1155(.A1(new_n1353), .A2(new_n1354), .A3(new_n1355), .ZN(new_n1356));
  NAND2_X1  g1156(.A1(new_n1355), .A2(new_n1354), .ZN(new_n1357));
  NAND4_X1  g1157(.A1(new_n1351), .A2(new_n1294), .A3(new_n1357), .A4(new_n1352), .ZN(new_n1358));
  NAND2_X1  g1158(.A1(new_n1356), .A2(new_n1358), .ZN(new_n1359));
  INV_X1    g1159(.A(new_n1291), .ZN(new_n1360));
  XNOR2_X1  g1160(.A(new_n1359), .B(new_n1360), .ZN(G402));
endmodule


