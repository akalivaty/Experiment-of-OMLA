//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 0 1 1 1 0 0 0 0 1 0 1 1 0 0 1 1 1 0 0 1 0 1 1 1 1 0 1 0 1 0 1 0 1 0 1 0 0 0 1 1 0 0 0 1 0 0 1 1 1 1 1 0 0 1 1 1 1 1 1 0 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:31:20 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n454, new_n458,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n488, new_n489,
    new_n490, new_n491, new_n492, new_n493, new_n494, new_n495, new_n496,
    new_n497, new_n498, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n514, new_n515, new_n516, new_n517, new_n518,
    new_n519, new_n520, new_n522, new_n523, new_n524, new_n525, new_n526,
    new_n527, new_n528, new_n529, new_n530, new_n531, new_n532, new_n533,
    new_n534, new_n535, new_n536, new_n537, new_n538, new_n539, new_n540,
    new_n541, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n557,
    new_n558, new_n559, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n576, new_n577, new_n578, new_n579, new_n580,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n591,
    new_n592, new_n593, new_n594, new_n595, new_n596, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n619, new_n622, new_n623, new_n625, new_n626,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n918, new_n919, new_n920, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1176, new_n1177, new_n1178;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n450));
  XNOR2_X1  g025(.A(KEYINPUT64), .B(KEYINPUT2), .ZN(new_n451));
  XNOR2_X1  g026(.A(new_n450), .B(new_n451), .ZN(new_n452));
  NOR4_X1   g027(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n453));
  INV_X1    g028(.A(new_n453), .ZN(new_n454));
  NOR2_X1   g029(.A1(new_n452), .A2(new_n454), .ZN(G325));
  INV_X1    g030(.A(G325), .ZN(G261));
  AOI22_X1  g031(.A1(new_n452), .A2(G2106), .B1(G567), .B2(new_n454), .ZN(G319));
  XNOR2_X1  g032(.A(KEYINPUT3), .B(G2104), .ZN(new_n458));
  AND2_X1   g033(.A1(new_n458), .A2(G125), .ZN(new_n459));
  AND2_X1   g034(.A1(G113), .A2(G2104), .ZN(new_n460));
  OAI21_X1  g035(.A(G2105), .B1(new_n459), .B2(new_n460), .ZN(new_n461));
  OR2_X1    g036(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n462));
  NAND2_X1  g037(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n463));
  AOI21_X1  g038(.A(G2105), .B1(new_n462), .B2(new_n463), .ZN(new_n464));
  INV_X1    g039(.A(G2105), .ZN(new_n465));
  AND2_X1   g040(.A1(new_n465), .A2(G2104), .ZN(new_n466));
  AOI22_X1  g041(.A1(new_n464), .A2(G137), .B1(G101), .B2(new_n466), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n461), .A2(new_n467), .ZN(new_n468));
  INV_X1    g043(.A(new_n468), .ZN(G160));
  OR2_X1    g044(.A1(G100), .A2(G2105), .ZN(new_n470));
  OAI211_X1 g045(.A(new_n470), .B(G2104), .C1(G112), .C2(new_n465), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n458), .A2(G2105), .ZN(new_n472));
  INV_X1    g047(.A(G124), .ZN(new_n473));
  OAI21_X1  g048(.A(new_n471), .B1(new_n472), .B2(new_n473), .ZN(new_n474));
  AOI21_X1  g049(.A(new_n474), .B1(G136), .B2(new_n464), .ZN(G162));
  NAND3_X1  g050(.A1(new_n458), .A2(G126), .A3(G2105), .ZN(new_n476));
  OR2_X1    g051(.A1(G102), .A2(G2105), .ZN(new_n477));
  OAI211_X1 g052(.A(new_n477), .B(G2104), .C1(G114), .C2(new_n465), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n476), .A2(new_n478), .ZN(new_n479));
  INV_X1    g054(.A(KEYINPUT65), .ZN(new_n480));
  INV_X1    g055(.A(KEYINPUT4), .ZN(new_n481));
  NOR2_X1   g056(.A1(new_n480), .A2(new_n481), .ZN(new_n482));
  NAND2_X1  g057(.A1(new_n458), .A2(new_n465), .ZN(new_n483));
  INV_X1    g058(.A(G138), .ZN(new_n484));
  OAI21_X1  g059(.A(new_n482), .B1(new_n483), .B2(new_n484), .ZN(new_n485));
  OAI211_X1 g060(.A(new_n464), .B(G138), .C1(new_n480), .C2(new_n481), .ZN(new_n486));
  AOI21_X1  g061(.A(new_n479), .B1(new_n485), .B2(new_n486), .ZN(G164));
  INV_X1    g062(.A(KEYINPUT5), .ZN(new_n488));
  NOR2_X1   g063(.A1(new_n488), .A2(G543), .ZN(new_n489));
  INV_X1    g064(.A(KEYINPUT66), .ZN(new_n490));
  INV_X1    g065(.A(G543), .ZN(new_n491));
  OAI21_X1  g066(.A(new_n490), .B1(new_n491), .B2(KEYINPUT5), .ZN(new_n492));
  NAND3_X1  g067(.A1(new_n488), .A2(KEYINPUT66), .A3(G543), .ZN(new_n493));
  AOI21_X1  g068(.A(new_n489), .B1(new_n492), .B2(new_n493), .ZN(new_n494));
  XNOR2_X1  g069(.A(KEYINPUT6), .B(G651), .ZN(new_n495));
  NAND2_X1  g070(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  INV_X1    g071(.A(G88), .ZN(new_n497));
  INV_X1    g072(.A(G50), .ZN(new_n498));
  NAND2_X1  g073(.A1(new_n495), .A2(G543), .ZN(new_n499));
  OAI22_X1  g074(.A1(new_n496), .A2(new_n497), .B1(new_n498), .B2(new_n499), .ZN(new_n500));
  NAND2_X1  g075(.A1(G75), .A2(G543), .ZN(new_n501));
  INV_X1    g076(.A(new_n489), .ZN(new_n502));
  AND3_X1   g077(.A1(new_n488), .A2(KEYINPUT66), .A3(G543), .ZN(new_n503));
  AOI21_X1  g078(.A(KEYINPUT66), .B1(new_n488), .B2(G543), .ZN(new_n504));
  OAI21_X1  g079(.A(new_n502), .B1(new_n503), .B2(new_n504), .ZN(new_n505));
  INV_X1    g080(.A(G62), .ZN(new_n506));
  OAI21_X1  g081(.A(new_n501), .B1(new_n505), .B2(new_n506), .ZN(new_n507));
  AOI21_X1  g082(.A(new_n500), .B1(G651), .B2(new_n507), .ZN(new_n508));
  NAND2_X1  g083(.A1(new_n508), .A2(KEYINPUT67), .ZN(new_n509));
  INV_X1    g084(.A(KEYINPUT67), .ZN(new_n510));
  AND2_X1   g085(.A1(new_n507), .A2(G651), .ZN(new_n511));
  OAI21_X1  g086(.A(new_n510), .B1(new_n511), .B2(new_n500), .ZN(new_n512));
  NAND2_X1  g087(.A1(new_n509), .A2(new_n512), .ZN(G166));
  AND2_X1   g088(.A1(new_n494), .A2(new_n495), .ZN(new_n514));
  AND2_X1   g089(.A1(new_n514), .A2(G89), .ZN(new_n515));
  NAND3_X1  g090(.A1(new_n494), .A2(G63), .A3(G651), .ZN(new_n516));
  NAND3_X1  g091(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n517));
  XNOR2_X1  g092(.A(new_n517), .B(KEYINPUT7), .ZN(new_n518));
  INV_X1    g093(.A(G51), .ZN(new_n519));
  OAI211_X1 g094(.A(new_n516), .B(new_n518), .C1(new_n519), .C2(new_n499), .ZN(new_n520));
  NOR2_X1   g095(.A1(new_n515), .A2(new_n520), .ZN(G168));
  INV_X1    g096(.A(KEYINPUT69), .ZN(new_n522));
  NAND2_X1  g097(.A1(G77), .A2(G543), .ZN(new_n523));
  INV_X1    g098(.A(new_n523), .ZN(new_n524));
  AOI21_X1  g099(.A(new_n524), .B1(new_n494), .B2(G64), .ZN(new_n525));
  OAI21_X1  g100(.A(G651), .B1(new_n525), .B2(KEYINPUT68), .ZN(new_n526));
  INV_X1    g101(.A(KEYINPUT68), .ZN(new_n527));
  AOI211_X1 g102(.A(new_n527), .B(new_n524), .C1(new_n494), .C2(G64), .ZN(new_n528));
  OAI21_X1  g103(.A(new_n522), .B1(new_n526), .B2(new_n528), .ZN(new_n529));
  XOR2_X1   g104(.A(KEYINPUT70), .B(G90), .Z(new_n530));
  NAND2_X1  g105(.A1(new_n514), .A2(new_n530), .ZN(new_n531));
  INV_X1    g106(.A(new_n499), .ZN(new_n532));
  NAND2_X1  g107(.A1(new_n532), .A2(G52), .ZN(new_n533));
  NAND2_X1  g108(.A1(new_n531), .A2(new_n533), .ZN(new_n534));
  INV_X1    g109(.A(new_n534), .ZN(new_n535));
  OAI211_X1 g110(.A(new_n502), .B(G64), .C1(new_n503), .C2(new_n504), .ZN(new_n536));
  NAND2_X1  g111(.A1(new_n536), .A2(new_n523), .ZN(new_n537));
  NAND2_X1  g112(.A1(new_n537), .A2(new_n527), .ZN(new_n538));
  NAND2_X1  g113(.A1(new_n525), .A2(KEYINPUT68), .ZN(new_n539));
  NAND4_X1  g114(.A1(new_n538), .A2(new_n539), .A3(KEYINPUT69), .A4(G651), .ZN(new_n540));
  NAND3_X1  g115(.A1(new_n529), .A2(new_n535), .A3(new_n540), .ZN(new_n541));
  INV_X1    g116(.A(new_n541), .ZN(G171));
  NAND3_X1  g117(.A1(new_n495), .A2(G43), .A3(G543), .ZN(new_n543));
  INV_X1    g118(.A(new_n543), .ZN(new_n544));
  AOI21_X1  g119(.A(new_n544), .B1(new_n514), .B2(G81), .ZN(new_n545));
  NAND2_X1  g120(.A1(G68), .A2(G543), .ZN(new_n546));
  INV_X1    g121(.A(new_n546), .ZN(new_n547));
  AOI21_X1  g122(.A(new_n547), .B1(new_n494), .B2(G56), .ZN(new_n548));
  INV_X1    g123(.A(KEYINPUT71), .ZN(new_n549));
  OAI21_X1  g124(.A(G651), .B1(new_n548), .B2(new_n549), .ZN(new_n550));
  AOI211_X1 g125(.A(KEYINPUT71), .B(new_n547), .C1(new_n494), .C2(G56), .ZN(new_n551));
  OAI21_X1  g126(.A(new_n545), .B1(new_n550), .B2(new_n551), .ZN(new_n552));
  INV_X1    g127(.A(G860), .ZN(new_n553));
  NOR2_X1   g128(.A1(new_n552), .A2(new_n553), .ZN(new_n554));
  XNOR2_X1  g129(.A(new_n554), .B(KEYINPUT72), .ZN(G153));
  NAND4_X1  g130(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  XOR2_X1   g131(.A(KEYINPUT73), .B(KEYINPUT8), .Z(new_n557));
  NAND2_X1  g132(.A1(G1), .A2(G3), .ZN(new_n558));
  XNOR2_X1  g133(.A(new_n557), .B(new_n558), .ZN(new_n559));
  NAND4_X1  g134(.A1(G319), .A2(G483), .A3(G661), .A4(new_n559), .ZN(G188));
  INV_X1    g135(.A(KEYINPUT74), .ZN(new_n561));
  NAND3_X1  g136(.A1(new_n494), .A2(G91), .A3(new_n495), .ZN(new_n562));
  NAND3_X1  g137(.A1(new_n495), .A2(G53), .A3(G543), .ZN(new_n563));
  NAND2_X1  g138(.A1(new_n563), .A2(KEYINPUT9), .ZN(new_n564));
  INV_X1    g139(.A(new_n564), .ZN(new_n565));
  NOR2_X1   g140(.A1(new_n563), .A2(KEYINPUT9), .ZN(new_n566));
  OAI21_X1  g141(.A(new_n562), .B1(new_n565), .B2(new_n566), .ZN(new_n567));
  INV_X1    g142(.A(G651), .ZN(new_n568));
  NAND2_X1  g143(.A1(new_n494), .A2(G65), .ZN(new_n569));
  NAND2_X1  g144(.A1(G78), .A2(G543), .ZN(new_n570));
  AOI21_X1  g145(.A(new_n568), .B1(new_n569), .B2(new_n570), .ZN(new_n571));
  OAI21_X1  g146(.A(new_n561), .B1(new_n567), .B2(new_n571), .ZN(new_n572));
  INV_X1    g147(.A(new_n572), .ZN(new_n573));
  NOR3_X1   g148(.A1(new_n567), .A2(new_n561), .A3(new_n571), .ZN(new_n574));
  NOR2_X1   g149(.A1(new_n573), .A2(new_n574), .ZN(G299));
  INV_X1    g150(.A(KEYINPUT75), .ZN(new_n576));
  NAND3_X1  g151(.A1(new_n538), .A2(new_n539), .A3(G651), .ZN(new_n577));
  AOI21_X1  g152(.A(new_n534), .B1(new_n577), .B2(new_n522), .ZN(new_n578));
  AOI21_X1  g153(.A(new_n576), .B1(new_n578), .B2(new_n540), .ZN(new_n579));
  AND4_X1   g154(.A1(new_n576), .A2(new_n529), .A3(new_n540), .A4(new_n535), .ZN(new_n580));
  NOR2_X1   g155(.A1(new_n579), .A2(new_n580), .ZN(G301));
  INV_X1    g156(.A(G168), .ZN(G286));
  INV_X1    g157(.A(G166), .ZN(G303));
  INV_X1    g158(.A(G87), .ZN(new_n584));
  INV_X1    g159(.A(G49), .ZN(new_n585));
  OAI22_X1  g160(.A1(new_n496), .A2(new_n584), .B1(new_n585), .B2(new_n499), .ZN(new_n586));
  INV_X1    g161(.A(G74), .ZN(new_n587));
  AOI21_X1  g162(.A(new_n568), .B1(new_n505), .B2(new_n587), .ZN(new_n588));
  NOR2_X1   g163(.A1(new_n586), .A2(new_n588), .ZN(new_n589));
  INV_X1    g164(.A(new_n589), .ZN(G288));
  AOI22_X1  g165(.A1(new_n514), .A2(G86), .B1(G48), .B2(new_n532), .ZN(new_n591));
  NAND2_X1  g166(.A1(G73), .A2(G543), .ZN(new_n592));
  XNOR2_X1  g167(.A(new_n592), .B(KEYINPUT76), .ZN(new_n593));
  INV_X1    g168(.A(G61), .ZN(new_n594));
  OAI21_X1  g169(.A(new_n593), .B1(new_n505), .B2(new_n594), .ZN(new_n595));
  NAND2_X1  g170(.A1(new_n595), .A2(G651), .ZN(new_n596));
  NAND2_X1  g171(.A1(new_n591), .A2(new_n596), .ZN(G305));
  AOI22_X1  g172(.A1(new_n494), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n598));
  NOR2_X1   g173(.A1(new_n598), .A2(new_n568), .ZN(new_n599));
  INV_X1    g174(.A(G85), .ZN(new_n600));
  XOR2_X1   g175(.A(KEYINPUT77), .B(G47), .Z(new_n601));
  OAI22_X1  g176(.A1(new_n496), .A2(new_n600), .B1(new_n499), .B2(new_n601), .ZN(new_n602));
  NOR2_X1   g177(.A1(new_n599), .A2(new_n602), .ZN(new_n603));
  INV_X1    g178(.A(new_n603), .ZN(G290));
  NAND2_X1  g179(.A1(G301), .A2(G868), .ZN(new_n605));
  INV_X1    g180(.A(KEYINPUT78), .ZN(new_n606));
  NOR2_X1   g181(.A1(new_n605), .A2(new_n606), .ZN(new_n607));
  AND3_X1   g182(.A1(new_n494), .A2(G92), .A3(new_n495), .ZN(new_n608));
  XNOR2_X1  g183(.A(new_n608), .B(KEYINPUT10), .ZN(new_n609));
  NAND2_X1  g184(.A1(G79), .A2(G543), .ZN(new_n610));
  INV_X1    g185(.A(G66), .ZN(new_n611));
  OAI21_X1  g186(.A(new_n610), .B1(new_n505), .B2(new_n611), .ZN(new_n612));
  AOI22_X1  g187(.A1(new_n612), .A2(G651), .B1(G54), .B2(new_n532), .ZN(new_n613));
  NAND2_X1  g188(.A1(new_n609), .A2(new_n613), .ZN(new_n614));
  INV_X1    g189(.A(G868), .ZN(new_n615));
  AOI21_X1  g190(.A(KEYINPUT78), .B1(new_n614), .B2(new_n615), .ZN(new_n616));
  AOI21_X1  g191(.A(new_n607), .B1(new_n605), .B2(new_n616), .ZN(G284));
  AOI21_X1  g192(.A(new_n607), .B1(new_n605), .B2(new_n616), .ZN(G321));
  NAND2_X1  g193(.A1(G299), .A2(new_n615), .ZN(new_n619));
  OAI21_X1  g194(.A(new_n619), .B1(new_n615), .B2(G168), .ZN(G297));
  OAI21_X1  g195(.A(new_n619), .B1(new_n615), .B2(G168), .ZN(G280));
  INV_X1    g196(.A(new_n614), .ZN(new_n622));
  INV_X1    g197(.A(G559), .ZN(new_n623));
  OAI21_X1  g198(.A(new_n622), .B1(new_n623), .B2(G860), .ZN(G148));
  NAND2_X1  g199(.A1(new_n552), .A2(new_n615), .ZN(new_n625));
  NOR2_X1   g200(.A1(new_n614), .A2(G559), .ZN(new_n626));
  OAI21_X1  g201(.A(new_n625), .B1(new_n626), .B2(new_n615), .ZN(G323));
  XNOR2_X1  g202(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g203(.A1(new_n464), .A2(G135), .ZN(new_n629));
  NOR2_X1   g204(.A1(new_n465), .A2(G111), .ZN(new_n630));
  OAI21_X1  g205(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n631));
  INV_X1    g206(.A(G123), .ZN(new_n632));
  OAI221_X1 g207(.A(new_n629), .B1(new_n630), .B2(new_n631), .C1(new_n632), .C2(new_n472), .ZN(new_n633));
  OR2_X1    g208(.A1(new_n633), .A2(KEYINPUT80), .ZN(new_n634));
  NAND2_X1  g209(.A1(new_n633), .A2(KEYINPUT80), .ZN(new_n635));
  NAND2_X1  g210(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  XOR2_X1   g211(.A(new_n636), .B(G2096), .Z(new_n637));
  NAND2_X1  g212(.A1(new_n458), .A2(new_n466), .ZN(new_n638));
  XOR2_X1   g213(.A(KEYINPUT79), .B(KEYINPUT12), .Z(new_n639));
  XNOR2_X1  g214(.A(new_n638), .B(new_n639), .ZN(new_n640));
  XNOR2_X1  g215(.A(KEYINPUT13), .B(G2100), .ZN(new_n641));
  XNOR2_X1  g216(.A(new_n640), .B(new_n641), .ZN(new_n642));
  NAND2_X1  g217(.A1(new_n637), .A2(new_n642), .ZN(G156));
  XNOR2_X1  g218(.A(G2443), .B(G2446), .ZN(new_n644));
  XNOR2_X1  g219(.A(new_n644), .B(KEYINPUT82), .ZN(new_n645));
  XNOR2_X1  g220(.A(new_n645), .B(G2451), .ZN(new_n646));
  XOR2_X1   g221(.A(G1341), .B(G1348), .Z(new_n647));
  XNOR2_X1  g222(.A(new_n646), .B(new_n647), .ZN(new_n648));
  XOR2_X1   g223(.A(KEYINPUT15), .B(G2435), .Z(new_n649));
  XNOR2_X1  g224(.A(new_n649), .B(G2438), .ZN(new_n650));
  XNOR2_X1  g225(.A(G2427), .B(G2430), .ZN(new_n651));
  XNOR2_X1  g226(.A(new_n651), .B(KEYINPUT83), .ZN(new_n652));
  OR2_X1    g227(.A1(new_n650), .A2(new_n652), .ZN(new_n653));
  NAND2_X1  g228(.A1(new_n650), .A2(new_n652), .ZN(new_n654));
  NAND3_X1  g229(.A1(new_n653), .A2(new_n654), .A3(KEYINPUT14), .ZN(new_n655));
  XNOR2_X1  g230(.A(new_n648), .B(new_n655), .ZN(new_n656));
  INV_X1    g231(.A(new_n656), .ZN(new_n657));
  XOR2_X1   g232(.A(KEYINPUT81), .B(KEYINPUT16), .Z(new_n658));
  XNOR2_X1  g233(.A(new_n658), .B(G2454), .ZN(new_n659));
  INV_X1    g234(.A(new_n659), .ZN(new_n660));
  OAI21_X1  g235(.A(G14), .B1(new_n657), .B2(new_n660), .ZN(new_n661));
  AOI21_X1  g236(.A(new_n661), .B1(new_n660), .B2(new_n657), .ZN(G401));
  XOR2_X1   g237(.A(G2084), .B(G2090), .Z(new_n663));
  XNOR2_X1  g238(.A(G2072), .B(G2078), .ZN(new_n664));
  XNOR2_X1  g239(.A(G2067), .B(G2678), .ZN(new_n665));
  NAND3_X1  g240(.A1(new_n663), .A2(new_n664), .A3(new_n665), .ZN(new_n666));
  XNOR2_X1  g241(.A(new_n666), .B(KEYINPUT84), .ZN(new_n667));
  XNOR2_X1  g242(.A(new_n667), .B(KEYINPUT18), .ZN(new_n668));
  INV_X1    g243(.A(new_n663), .ZN(new_n669));
  OAI21_X1  g244(.A(new_n669), .B1(new_n664), .B2(new_n665), .ZN(new_n670));
  XOR2_X1   g245(.A(new_n670), .B(KEYINPUT85), .Z(new_n671));
  XOR2_X1   g246(.A(new_n664), .B(KEYINPUT17), .Z(new_n672));
  NAND2_X1  g247(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  AOI21_X1  g248(.A(new_n671), .B1(new_n663), .B2(new_n672), .ZN(new_n674));
  OAI211_X1 g249(.A(new_n668), .B(new_n673), .C1(new_n674), .C2(new_n665), .ZN(new_n675));
  XOR2_X1   g250(.A(G2096), .B(G2100), .Z(new_n676));
  XNOR2_X1  g251(.A(new_n675), .B(new_n676), .ZN(G227));
  XNOR2_X1  g252(.A(G1971), .B(G1976), .ZN(new_n678));
  XNOR2_X1  g253(.A(new_n678), .B(KEYINPUT19), .ZN(new_n679));
  INV_X1    g254(.A(KEYINPUT86), .ZN(new_n680));
  XNOR2_X1  g255(.A(G1956), .B(G2474), .ZN(new_n681));
  INV_X1    g256(.A(new_n681), .ZN(new_n682));
  XNOR2_X1  g257(.A(G1961), .B(G1966), .ZN(new_n683));
  INV_X1    g258(.A(new_n683), .ZN(new_n684));
  NAND2_X1  g259(.A1(new_n682), .A2(new_n684), .ZN(new_n685));
  AOI21_X1  g260(.A(new_n679), .B1(new_n680), .B2(new_n685), .ZN(new_n686));
  OAI21_X1  g261(.A(new_n686), .B1(new_n680), .B2(new_n685), .ZN(new_n687));
  XNOR2_X1  g262(.A(new_n687), .B(KEYINPUT20), .ZN(new_n688));
  NOR2_X1   g263(.A1(new_n682), .A2(new_n684), .ZN(new_n689));
  INV_X1    g264(.A(new_n689), .ZN(new_n690));
  NAND3_X1  g265(.A1(new_n690), .A2(new_n685), .A3(new_n679), .ZN(new_n691));
  OAI211_X1 g266(.A(new_n688), .B(new_n691), .C1(new_n679), .C2(new_n690), .ZN(new_n692));
  XNOR2_X1  g267(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n693));
  XNOR2_X1  g268(.A(new_n692), .B(new_n693), .ZN(new_n694));
  XNOR2_X1  g269(.A(G1991), .B(G1996), .ZN(new_n695));
  XNOR2_X1  g270(.A(new_n695), .B(KEYINPUT87), .ZN(new_n696));
  XNOR2_X1  g271(.A(new_n694), .B(new_n696), .ZN(new_n697));
  XNOR2_X1  g272(.A(G1981), .B(G1986), .ZN(new_n698));
  OR2_X1    g273(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  NAND2_X1  g274(.A1(new_n697), .A2(new_n698), .ZN(new_n700));
  NAND2_X1  g275(.A1(new_n699), .A2(new_n700), .ZN(G229));
  NAND2_X1  g276(.A1(G299), .A2(G16), .ZN(new_n702));
  INV_X1    g277(.A(G16), .ZN(new_n703));
  NAND2_X1  g278(.A1(new_n703), .A2(G20), .ZN(new_n704));
  XNOR2_X1  g279(.A(new_n704), .B(KEYINPUT23), .ZN(new_n705));
  NAND2_X1  g280(.A1(new_n702), .A2(new_n705), .ZN(new_n706));
  XNOR2_X1  g281(.A(new_n706), .B(KEYINPUT99), .ZN(new_n707));
  XNOR2_X1  g282(.A(KEYINPUT98), .B(G1956), .ZN(new_n708));
  XNOR2_X1  g283(.A(new_n707), .B(new_n708), .ZN(new_n709));
  MUX2_X1   g284(.A(G19), .B(new_n552), .S(G16), .Z(new_n710));
  XOR2_X1   g285(.A(new_n710), .B(G1341), .Z(new_n711));
  NAND2_X1  g286(.A1(new_n622), .A2(G16), .ZN(new_n712));
  OAI21_X1  g287(.A(new_n712), .B1(G4), .B2(G16), .ZN(new_n713));
  INV_X1    g288(.A(G1348), .ZN(new_n714));
  AND2_X1   g289(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  NOR2_X1   g290(.A1(new_n713), .A2(new_n714), .ZN(new_n716));
  XOR2_X1   g291(.A(KEYINPUT88), .B(G29), .Z(new_n717));
  INV_X1    g292(.A(new_n717), .ZN(new_n718));
  NOR2_X1   g293(.A1(new_n718), .A2(G27), .ZN(new_n719));
  AOI21_X1  g294(.A(new_n719), .B1(G164), .B2(new_n718), .ZN(new_n720));
  XNOR2_X1  g295(.A(new_n720), .B(G2078), .ZN(new_n721));
  NOR2_X1   g296(.A1(new_n721), .A2(KEYINPUT96), .ZN(new_n722));
  NOR3_X1   g297(.A1(new_n715), .A2(new_n716), .A3(new_n722), .ZN(new_n723));
  NAND2_X1  g298(.A1(G162), .A2(new_n718), .ZN(new_n724));
  OAI21_X1  g299(.A(new_n724), .B1(G35), .B2(new_n718), .ZN(new_n725));
  XNOR2_X1  g300(.A(KEYINPUT97), .B(KEYINPUT29), .ZN(new_n726));
  XNOR2_X1  g301(.A(new_n726), .B(G2090), .ZN(new_n727));
  OR2_X1    g302(.A1(new_n725), .A2(new_n727), .ZN(new_n728));
  NAND2_X1  g303(.A1(new_n725), .A2(new_n727), .ZN(new_n729));
  OAI211_X1 g304(.A(new_n728), .B(new_n729), .C1(new_n636), .C2(new_n717), .ZN(new_n730));
  INV_X1    g305(.A(KEYINPUT24), .ZN(new_n731));
  OR2_X1    g306(.A1(new_n731), .A2(G34), .ZN(new_n732));
  NAND2_X1  g307(.A1(new_n731), .A2(G34), .ZN(new_n733));
  NAND3_X1  g308(.A1(new_n717), .A2(new_n732), .A3(new_n733), .ZN(new_n734));
  INV_X1    g309(.A(G29), .ZN(new_n735));
  OAI21_X1  g310(.A(new_n734), .B1(new_n468), .B2(new_n735), .ZN(new_n736));
  INV_X1    g311(.A(G2084), .ZN(new_n737));
  NOR2_X1   g312(.A1(new_n736), .A2(new_n737), .ZN(new_n738));
  XOR2_X1   g313(.A(new_n738), .B(KEYINPUT93), .Z(new_n739));
  AND3_X1   g314(.A1(new_n717), .A2(KEYINPUT28), .A3(G26), .ZN(new_n740));
  AOI21_X1  g315(.A(KEYINPUT28), .B1(new_n717), .B2(G26), .ZN(new_n741));
  NAND2_X1  g316(.A1(new_n464), .A2(G140), .ZN(new_n742));
  OR2_X1    g317(.A1(G104), .A2(G2105), .ZN(new_n743));
  OAI211_X1 g318(.A(new_n743), .B(G2104), .C1(G116), .C2(new_n465), .ZN(new_n744));
  INV_X1    g319(.A(G128), .ZN(new_n745));
  OAI211_X1 g320(.A(new_n742), .B(new_n744), .C1(new_n745), .C2(new_n472), .ZN(new_n746));
  AOI211_X1 g321(.A(new_n740), .B(new_n741), .C1(new_n746), .C2(G29), .ZN(new_n747));
  INV_X1    g322(.A(new_n747), .ZN(new_n748));
  AND2_X1   g323(.A1(new_n735), .A2(G32), .ZN(new_n749));
  AOI22_X1  g324(.A1(new_n464), .A2(G141), .B1(G105), .B2(new_n466), .ZN(new_n750));
  NAND3_X1  g325(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n751));
  XOR2_X1   g326(.A(new_n751), .B(KEYINPUT26), .Z(new_n752));
  INV_X1    g327(.A(G129), .ZN(new_n753));
  OAI211_X1 g328(.A(new_n750), .B(new_n752), .C1(new_n753), .C2(new_n472), .ZN(new_n754));
  AOI21_X1  g329(.A(new_n749), .B1(new_n754), .B2(G29), .ZN(new_n755));
  XNOR2_X1  g330(.A(KEYINPUT27), .B(G1996), .ZN(new_n756));
  OAI22_X1  g331(.A1(new_n748), .A2(G2067), .B1(new_n755), .B2(new_n756), .ZN(new_n757));
  NAND2_X1  g332(.A1(new_n755), .A2(new_n756), .ZN(new_n758));
  AND2_X1   g333(.A1(new_n458), .A2(G127), .ZN(new_n759));
  AND2_X1   g334(.A1(G115), .A2(G2104), .ZN(new_n760));
  OAI21_X1  g335(.A(G2105), .B1(new_n759), .B2(new_n760), .ZN(new_n761));
  NAND3_X1  g336(.A1(new_n465), .A2(G103), .A3(G2104), .ZN(new_n762));
  INV_X1    g337(.A(KEYINPUT25), .ZN(new_n763));
  OR2_X1    g338(.A1(new_n762), .A2(new_n763), .ZN(new_n764));
  NAND2_X1  g339(.A1(new_n762), .A2(new_n763), .ZN(new_n765));
  AOI22_X1  g340(.A1(new_n764), .A2(new_n765), .B1(new_n464), .B2(G139), .ZN(new_n766));
  NAND2_X1  g341(.A1(new_n761), .A2(new_n766), .ZN(new_n767));
  MUX2_X1   g342(.A(G33), .B(new_n767), .S(G29), .Z(new_n768));
  INV_X1    g343(.A(new_n768), .ZN(new_n769));
  INV_X1    g344(.A(G2072), .ZN(new_n770));
  OAI21_X1  g345(.A(new_n758), .B1(new_n769), .B2(new_n770), .ZN(new_n771));
  NOR4_X1   g346(.A1(new_n730), .A2(new_n739), .A3(new_n757), .A4(new_n771), .ZN(new_n772));
  NAND2_X1  g347(.A1(new_n703), .A2(G21), .ZN(new_n773));
  OAI21_X1  g348(.A(new_n773), .B1(G168), .B2(new_n703), .ZN(new_n774));
  INV_X1    g349(.A(G1966), .ZN(new_n775));
  XNOR2_X1  g350(.A(new_n774), .B(new_n775), .ZN(new_n776));
  XNOR2_X1  g351(.A(KEYINPUT94), .B(G28), .ZN(new_n777));
  INV_X1    g352(.A(KEYINPUT30), .ZN(new_n778));
  AOI21_X1  g353(.A(G29), .B1(new_n777), .B2(new_n778), .ZN(new_n779));
  OAI21_X1  g354(.A(new_n779), .B1(new_n778), .B2(new_n777), .ZN(new_n780));
  XNOR2_X1  g355(.A(KEYINPUT31), .B(G11), .ZN(new_n781));
  NAND2_X1  g356(.A1(new_n780), .A2(new_n781), .ZN(new_n782));
  AOI21_X1  g357(.A(new_n782), .B1(new_n769), .B2(new_n770), .ZN(new_n783));
  AOI22_X1  g358(.A1(new_n748), .A2(G2067), .B1(new_n736), .B2(new_n737), .ZN(new_n784));
  NAND3_X1  g359(.A1(new_n776), .A2(new_n783), .A3(new_n784), .ZN(new_n785));
  AOI21_X1  g360(.A(new_n785), .B1(KEYINPUT96), .B2(new_n721), .ZN(new_n786));
  AND4_X1   g361(.A1(new_n711), .A2(new_n723), .A3(new_n772), .A4(new_n786), .ZN(new_n787));
  NAND2_X1  g362(.A1(new_n703), .A2(G5), .ZN(new_n788));
  OAI21_X1  g363(.A(new_n788), .B1(G171), .B2(new_n703), .ZN(new_n789));
  XOR2_X1   g364(.A(new_n789), .B(KEYINPUT95), .Z(new_n790));
  OR2_X1    g365(.A1(new_n790), .A2(G1961), .ZN(new_n791));
  NAND2_X1  g366(.A1(new_n790), .A2(G1961), .ZN(new_n792));
  NAND4_X1  g367(.A1(new_n709), .A2(new_n787), .A3(new_n791), .A4(new_n792), .ZN(new_n793));
  NAND2_X1  g368(.A1(G166), .A2(G16), .ZN(new_n794));
  OAI21_X1  g369(.A(new_n794), .B1(G16), .B2(G22), .ZN(new_n795));
  OR2_X1    g370(.A1(new_n795), .A2(KEYINPUT92), .ZN(new_n796));
  NAND2_X1  g371(.A1(new_n795), .A2(KEYINPUT92), .ZN(new_n797));
  NAND2_X1  g372(.A1(new_n796), .A2(new_n797), .ZN(new_n798));
  INV_X1    g373(.A(G1971), .ZN(new_n799));
  NAND2_X1  g374(.A1(new_n798), .A2(new_n799), .ZN(new_n800));
  NAND3_X1  g375(.A1(new_n796), .A2(G1971), .A3(new_n797), .ZN(new_n801));
  AND2_X1   g376(.A1(new_n703), .A2(G6), .ZN(new_n802));
  AOI21_X1  g377(.A(new_n802), .B1(G305), .B2(G16), .ZN(new_n803));
  XNOR2_X1  g378(.A(new_n803), .B(KEYINPUT91), .ZN(new_n804));
  XOR2_X1   g379(.A(KEYINPUT32), .B(G1981), .Z(new_n805));
  XNOR2_X1  g380(.A(new_n804), .B(new_n805), .ZN(new_n806));
  NAND2_X1  g381(.A1(new_n703), .A2(G23), .ZN(new_n807));
  OAI21_X1  g382(.A(new_n807), .B1(new_n589), .B2(new_n703), .ZN(new_n808));
  XNOR2_X1  g383(.A(KEYINPUT33), .B(G1976), .ZN(new_n809));
  XNOR2_X1  g384(.A(new_n808), .B(new_n809), .ZN(new_n810));
  NAND4_X1  g385(.A1(new_n800), .A2(new_n801), .A3(new_n806), .A4(new_n810), .ZN(new_n811));
  XNOR2_X1  g386(.A(KEYINPUT90), .B(KEYINPUT34), .ZN(new_n812));
  OR2_X1    g387(.A1(new_n811), .A2(new_n812), .ZN(new_n813));
  NAND2_X1  g388(.A1(new_n811), .A2(new_n812), .ZN(new_n814));
  NAND2_X1  g389(.A1(new_n464), .A2(G131), .ZN(new_n815));
  NOR2_X1   g390(.A1(new_n465), .A2(G107), .ZN(new_n816));
  OAI21_X1  g391(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n817));
  INV_X1    g392(.A(G119), .ZN(new_n818));
  OAI221_X1 g393(.A(new_n815), .B1(new_n816), .B2(new_n817), .C1(new_n818), .C2(new_n472), .ZN(new_n819));
  MUX2_X1   g394(.A(G25), .B(new_n819), .S(new_n718), .Z(new_n820));
  XNOR2_X1  g395(.A(KEYINPUT35), .B(G1991), .ZN(new_n821));
  XOR2_X1   g396(.A(new_n820), .B(new_n821), .Z(new_n822));
  NAND2_X1  g397(.A1(new_n703), .A2(G24), .ZN(new_n823));
  XNOR2_X1  g398(.A(new_n823), .B(KEYINPUT89), .ZN(new_n824));
  OAI21_X1  g399(.A(new_n824), .B1(new_n603), .B2(new_n703), .ZN(new_n825));
  OAI21_X1  g400(.A(new_n822), .B1(G1986), .B2(new_n825), .ZN(new_n826));
  AOI21_X1  g401(.A(new_n826), .B1(G1986), .B2(new_n825), .ZN(new_n827));
  NAND3_X1  g402(.A1(new_n813), .A2(new_n814), .A3(new_n827), .ZN(new_n828));
  OR2_X1    g403(.A1(new_n828), .A2(KEYINPUT36), .ZN(new_n829));
  NAND2_X1  g404(.A1(new_n828), .A2(KEYINPUT36), .ZN(new_n830));
  AOI21_X1  g405(.A(new_n793), .B1(new_n829), .B2(new_n830), .ZN(G311));
  INV_X1    g406(.A(G311), .ZN(G150));
  NAND2_X1  g407(.A1(new_n622), .A2(G559), .ZN(new_n833));
  XNOR2_X1  g408(.A(new_n833), .B(KEYINPUT38), .ZN(new_n834));
  NAND2_X1  g409(.A1(new_n494), .A2(G67), .ZN(new_n835));
  NAND2_X1  g410(.A1(G80), .A2(G543), .ZN(new_n836));
  AOI21_X1  g411(.A(new_n568), .B1(new_n835), .B2(new_n836), .ZN(new_n837));
  NAND3_X1  g412(.A1(new_n494), .A2(G93), .A3(new_n495), .ZN(new_n838));
  NAND3_X1  g413(.A1(new_n495), .A2(G55), .A3(G543), .ZN(new_n839));
  NAND2_X1  g414(.A1(new_n838), .A2(new_n839), .ZN(new_n840));
  OR2_X1    g415(.A1(new_n837), .A2(new_n840), .ZN(new_n841));
  NAND2_X1  g416(.A1(new_n552), .A2(new_n841), .ZN(new_n842));
  OAI211_X1 g417(.A(new_n502), .B(G56), .C1(new_n503), .C2(new_n504), .ZN(new_n843));
  NAND2_X1  g418(.A1(new_n843), .A2(new_n546), .ZN(new_n844));
  NAND2_X1  g419(.A1(new_n844), .A2(KEYINPUT71), .ZN(new_n845));
  NAND2_X1  g420(.A1(new_n548), .A2(new_n549), .ZN(new_n846));
  NAND3_X1  g421(.A1(new_n845), .A2(new_n846), .A3(G651), .ZN(new_n847));
  NOR2_X1   g422(.A1(new_n837), .A2(new_n840), .ZN(new_n848));
  NAND3_X1  g423(.A1(new_n847), .A2(new_n848), .A3(new_n545), .ZN(new_n849));
  NAND2_X1  g424(.A1(new_n842), .A2(new_n849), .ZN(new_n850));
  INV_X1    g425(.A(new_n850), .ZN(new_n851));
  XNOR2_X1  g426(.A(new_n834), .B(new_n851), .ZN(new_n852));
  OR2_X1    g427(.A1(new_n852), .A2(KEYINPUT39), .ZN(new_n853));
  NAND2_X1  g428(.A1(new_n852), .A2(KEYINPUT39), .ZN(new_n854));
  NAND3_X1  g429(.A1(new_n853), .A2(new_n553), .A3(new_n854), .ZN(new_n855));
  NOR2_X1   g430(.A1(new_n848), .A2(new_n553), .ZN(new_n856));
  XNOR2_X1  g431(.A(new_n856), .B(KEYINPUT37), .ZN(new_n857));
  NAND2_X1  g432(.A1(new_n855), .A2(new_n857), .ZN(G145));
  AND3_X1   g433(.A1(new_n476), .A2(KEYINPUT101), .A3(new_n478), .ZN(new_n859));
  AOI21_X1  g434(.A(KEYINPUT101), .B1(new_n476), .B2(new_n478), .ZN(new_n860));
  NOR2_X1   g435(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  INV_X1    g436(.A(KEYINPUT100), .ZN(new_n862));
  AND3_X1   g437(.A1(new_n485), .A2(new_n862), .A3(new_n486), .ZN(new_n863));
  AOI21_X1  g438(.A(new_n862), .B1(new_n485), .B2(new_n486), .ZN(new_n864));
  OAI21_X1  g439(.A(new_n861), .B1(new_n863), .B2(new_n864), .ZN(new_n865));
  XNOR2_X1  g440(.A(new_n865), .B(new_n746), .ZN(new_n866));
  INV_X1    g441(.A(G130), .ZN(new_n867));
  NOR2_X1   g442(.A1(new_n465), .A2(G118), .ZN(new_n868));
  OAI21_X1  g443(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n869));
  OAI22_X1  g444(.A1(new_n472), .A2(new_n867), .B1(new_n868), .B2(new_n869), .ZN(new_n870));
  AOI21_X1  g445(.A(new_n870), .B1(G142), .B2(new_n464), .ZN(new_n871));
  XOR2_X1   g446(.A(new_n866), .B(new_n871), .Z(new_n872));
  XNOR2_X1  g447(.A(new_n767), .B(new_n754), .ZN(new_n873));
  XNOR2_X1  g448(.A(new_n819), .B(new_n640), .ZN(new_n874));
  XNOR2_X1  g449(.A(new_n873), .B(new_n874), .ZN(new_n875));
  XNOR2_X1  g450(.A(new_n872), .B(new_n875), .ZN(new_n876));
  XNOR2_X1  g451(.A(new_n636), .B(G160), .ZN(new_n877));
  XNOR2_X1  g452(.A(new_n877), .B(G162), .ZN(new_n878));
  AOI21_X1  g453(.A(G37), .B1(new_n876), .B2(new_n878), .ZN(new_n879));
  OAI21_X1  g454(.A(new_n879), .B1(new_n878), .B2(new_n876), .ZN(new_n880));
  XNOR2_X1  g455(.A(new_n880), .B(KEYINPUT40), .ZN(G395));
  XNOR2_X1  g456(.A(new_n626), .B(new_n850), .ZN(new_n882));
  OR2_X1    g457(.A1(new_n563), .A2(KEYINPUT9), .ZN(new_n883));
  AOI22_X1  g458(.A1(new_n883), .A2(new_n564), .B1(new_n514), .B2(G91), .ZN(new_n884));
  INV_X1    g459(.A(new_n571), .ZN(new_n885));
  NAND3_X1  g460(.A1(new_n884), .A2(KEYINPUT74), .A3(new_n885), .ZN(new_n886));
  AND4_X1   g461(.A1(new_n572), .A2(new_n886), .A3(new_n609), .A4(new_n613), .ZN(new_n887));
  AOI22_X1  g462(.A1(new_n572), .A2(new_n886), .B1(new_n609), .B2(new_n613), .ZN(new_n888));
  NOR2_X1   g463(.A1(new_n887), .A2(new_n888), .ZN(new_n889));
  OR3_X1    g464(.A1(new_n882), .A2(KEYINPUT102), .A3(new_n889), .ZN(new_n890));
  OAI21_X1  g465(.A(KEYINPUT102), .B1(new_n882), .B2(new_n889), .ZN(new_n891));
  INV_X1    g466(.A(KEYINPUT41), .ZN(new_n892));
  OAI21_X1  g467(.A(new_n892), .B1(new_n887), .B2(new_n888), .ZN(new_n893));
  OAI21_X1  g468(.A(new_n614), .B1(new_n573), .B2(new_n574), .ZN(new_n894));
  NAND4_X1  g469(.A1(new_n572), .A2(new_n886), .A3(new_n609), .A4(new_n613), .ZN(new_n895));
  NAND3_X1  g470(.A1(new_n894), .A2(KEYINPUT41), .A3(new_n895), .ZN(new_n896));
  NAND2_X1  g471(.A1(new_n893), .A2(new_n896), .ZN(new_n897));
  NAND2_X1  g472(.A1(new_n897), .A2(new_n882), .ZN(new_n898));
  NAND3_X1  g473(.A1(new_n890), .A2(new_n891), .A3(new_n898), .ZN(new_n899));
  OR2_X1    g474(.A1(new_n899), .A2(KEYINPUT42), .ZN(new_n900));
  XNOR2_X1  g475(.A(G305), .B(new_n603), .ZN(new_n901));
  NOR2_X1   g476(.A1(new_n508), .A2(KEYINPUT67), .ZN(new_n902));
  NOR3_X1   g477(.A1(new_n511), .A2(new_n510), .A3(new_n500), .ZN(new_n903));
  NOR3_X1   g478(.A1(new_n902), .A2(new_n903), .A3(new_n589), .ZN(new_n904));
  AOI21_X1  g479(.A(G288), .B1(new_n509), .B2(new_n512), .ZN(new_n905));
  OAI21_X1  g480(.A(new_n901), .B1(new_n904), .B2(new_n905), .ZN(new_n906));
  XOR2_X1   g481(.A(G305), .B(new_n603), .Z(new_n907));
  OAI21_X1  g482(.A(new_n589), .B1(new_n902), .B2(new_n903), .ZN(new_n908));
  NAND3_X1  g483(.A1(new_n509), .A2(new_n512), .A3(G288), .ZN(new_n909));
  NAND3_X1  g484(.A1(new_n907), .A2(new_n908), .A3(new_n909), .ZN(new_n910));
  AND2_X1   g485(.A1(new_n906), .A2(new_n910), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n899), .A2(KEYINPUT42), .ZN(new_n912));
  AND3_X1   g487(.A1(new_n900), .A2(new_n911), .A3(new_n912), .ZN(new_n913));
  AOI21_X1  g488(.A(new_n911), .B1(new_n900), .B2(new_n912), .ZN(new_n914));
  OAI21_X1  g489(.A(G868), .B1(new_n913), .B2(new_n914), .ZN(new_n915));
  NAND2_X1  g490(.A1(new_n841), .A2(new_n615), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n915), .A2(new_n916), .ZN(G295));
  INV_X1    g492(.A(KEYINPUT103), .ZN(new_n918));
  AND3_X1   g493(.A1(new_n915), .A2(new_n918), .A3(new_n916), .ZN(new_n919));
  AOI21_X1  g494(.A(new_n918), .B1(new_n915), .B2(new_n916), .ZN(new_n920));
  NOR2_X1   g495(.A1(new_n919), .A2(new_n920), .ZN(G331));
  AND3_X1   g496(.A1(new_n906), .A2(new_n910), .A3(KEYINPUT105), .ZN(new_n922));
  AOI21_X1  g497(.A(KEYINPUT105), .B1(new_n906), .B2(new_n910), .ZN(new_n923));
  NOR2_X1   g498(.A1(new_n922), .A2(new_n923), .ZN(new_n924));
  INV_X1    g499(.A(KEYINPUT104), .ZN(new_n925));
  AND3_X1   g500(.A1(new_n842), .A2(new_n925), .A3(new_n849), .ZN(new_n926));
  AOI21_X1  g501(.A(new_n925), .B1(new_n842), .B2(new_n849), .ZN(new_n927));
  NOR2_X1   g502(.A1(new_n926), .A2(new_n927), .ZN(new_n928));
  NAND2_X1  g503(.A1(new_n541), .A2(KEYINPUT75), .ZN(new_n929));
  NAND3_X1  g504(.A1(new_n578), .A2(new_n576), .A3(new_n540), .ZN(new_n930));
  AOI21_X1  g505(.A(G286), .B1(new_n929), .B2(new_n930), .ZN(new_n931));
  NAND2_X1  g506(.A1(new_n541), .A2(G286), .ZN(new_n932));
  INV_X1    g507(.A(new_n932), .ZN(new_n933));
  OAI21_X1  g508(.A(new_n928), .B1(new_n931), .B2(new_n933), .ZN(new_n934));
  OAI21_X1  g509(.A(G168), .B1(new_n579), .B2(new_n580), .ZN(new_n935));
  NOR2_X1   g510(.A1(new_n552), .A2(new_n841), .ZN(new_n936));
  AOI21_X1  g511(.A(new_n848), .B1(new_n847), .B2(new_n545), .ZN(new_n937));
  OAI21_X1  g512(.A(KEYINPUT104), .B1(new_n936), .B2(new_n937), .ZN(new_n938));
  NAND3_X1  g513(.A1(new_n842), .A2(new_n925), .A3(new_n849), .ZN(new_n939));
  NAND2_X1  g514(.A1(new_n938), .A2(new_n939), .ZN(new_n940));
  NAND3_X1  g515(.A1(new_n935), .A2(new_n940), .A3(new_n932), .ZN(new_n941));
  AND3_X1   g516(.A1(new_n934), .A2(new_n941), .A3(new_n897), .ZN(new_n942));
  AOI21_X1  g517(.A(new_n889), .B1(new_n934), .B2(new_n941), .ZN(new_n943));
  OAI21_X1  g518(.A(new_n924), .B1(new_n942), .B2(new_n943), .ZN(new_n944));
  INV_X1    g519(.A(new_n889), .ZN(new_n945));
  AND3_X1   g520(.A1(new_n935), .A2(new_n940), .A3(new_n932), .ZN(new_n946));
  AOI21_X1  g521(.A(new_n940), .B1(new_n935), .B2(new_n932), .ZN(new_n947));
  OAI21_X1  g522(.A(new_n945), .B1(new_n946), .B2(new_n947), .ZN(new_n948));
  NAND3_X1  g523(.A1(new_n934), .A2(new_n941), .A3(new_n897), .ZN(new_n949));
  NAND3_X1  g524(.A1(new_n948), .A2(new_n911), .A3(new_n949), .ZN(new_n950));
  INV_X1    g525(.A(G37), .ZN(new_n951));
  NAND3_X1  g526(.A1(new_n944), .A2(new_n950), .A3(new_n951), .ZN(new_n952));
  INV_X1    g527(.A(KEYINPUT107), .ZN(new_n953));
  OR2_X1    g528(.A1(new_n893), .A2(new_n953), .ZN(new_n954));
  NAND3_X1  g529(.A1(new_n893), .A2(new_n896), .A3(new_n953), .ZN(new_n955));
  AND4_X1   g530(.A1(new_n934), .A2(new_n954), .A3(new_n941), .A4(new_n955), .ZN(new_n956));
  OAI21_X1  g531(.A(new_n924), .B1(new_n956), .B2(new_n943), .ZN(new_n957));
  NAND3_X1  g532(.A1(new_n957), .A2(new_n951), .A3(new_n950), .ZN(new_n958));
  INV_X1    g533(.A(KEYINPUT109), .ZN(new_n959));
  AND3_X1   g534(.A1(new_n958), .A2(new_n959), .A3(KEYINPUT43), .ZN(new_n960));
  AOI21_X1  g535(.A(new_n959), .B1(new_n958), .B2(KEYINPUT43), .ZN(new_n961));
  OAI221_X1 g536(.A(KEYINPUT44), .B1(KEYINPUT43), .B2(new_n952), .C1(new_n960), .C2(new_n961), .ZN(new_n962));
  NAND2_X1  g537(.A1(new_n952), .A2(KEYINPUT43), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n963), .A2(KEYINPUT106), .ZN(new_n964));
  INV_X1    g539(.A(KEYINPUT106), .ZN(new_n965));
  NAND3_X1  g540(.A1(new_n952), .A2(new_n965), .A3(KEYINPUT43), .ZN(new_n966));
  INV_X1    g541(.A(KEYINPUT43), .ZN(new_n967));
  NAND4_X1  g542(.A1(new_n957), .A2(new_n967), .A3(new_n951), .A4(new_n950), .ZN(new_n968));
  NAND3_X1  g543(.A1(new_n964), .A2(new_n966), .A3(new_n968), .ZN(new_n969));
  INV_X1    g544(.A(KEYINPUT44), .ZN(new_n970));
  AND3_X1   g545(.A1(new_n969), .A2(KEYINPUT108), .A3(new_n970), .ZN(new_n971));
  AOI21_X1  g546(.A(KEYINPUT108), .B1(new_n969), .B2(new_n970), .ZN(new_n972));
  OAI21_X1  g547(.A(new_n962), .B1(new_n971), .B2(new_n972), .ZN(G397));
  NOR2_X1   g548(.A1(new_n746), .A2(G2067), .ZN(new_n974));
  NAND2_X1  g549(.A1(new_n485), .A2(new_n486), .ZN(new_n975));
  NAND2_X1  g550(.A1(new_n975), .A2(KEYINPUT100), .ZN(new_n976));
  NAND3_X1  g551(.A1(new_n485), .A2(new_n862), .A3(new_n486), .ZN(new_n977));
  NAND2_X1  g552(.A1(new_n976), .A2(new_n977), .ZN(new_n978));
  AOI21_X1  g553(.A(G1384), .B1(new_n978), .B2(new_n861), .ZN(new_n979));
  NAND3_X1  g554(.A1(new_n461), .A2(G40), .A3(new_n467), .ZN(new_n980));
  NOR3_X1   g555(.A1(new_n979), .A2(KEYINPUT45), .A3(new_n980), .ZN(new_n981));
  NAND3_X1  g556(.A1(new_n981), .A2(G1996), .A3(new_n754), .ZN(new_n982));
  XNOR2_X1  g557(.A(new_n982), .B(KEYINPUT110), .ZN(new_n983));
  XNOR2_X1  g558(.A(new_n746), .B(G2067), .ZN(new_n984));
  NOR2_X1   g559(.A1(new_n754), .A2(G1996), .ZN(new_n985));
  OR2_X1    g560(.A1(new_n984), .A2(new_n985), .ZN(new_n986));
  AOI21_X1  g561(.A(new_n983), .B1(new_n981), .B2(new_n986), .ZN(new_n987));
  NOR2_X1   g562(.A1(new_n819), .A2(new_n821), .ZN(new_n988));
  AOI21_X1  g563(.A(new_n974), .B1(new_n987), .B2(new_n988), .ZN(new_n989));
  INV_X1    g564(.A(new_n981), .ZN(new_n990));
  NOR2_X1   g565(.A1(new_n989), .A2(new_n990), .ZN(new_n991));
  INV_X1    g566(.A(G1996), .ZN(new_n992));
  NAND3_X1  g567(.A1(new_n981), .A2(KEYINPUT46), .A3(new_n992), .ZN(new_n993));
  XOR2_X1   g568(.A(new_n993), .B(KEYINPUT127), .Z(new_n994));
  AOI21_X1  g569(.A(KEYINPUT46), .B1(new_n981), .B2(new_n992), .ZN(new_n995));
  XNOR2_X1  g570(.A(new_n995), .B(KEYINPUT126), .ZN(new_n996));
  OAI21_X1  g571(.A(new_n981), .B1(new_n754), .B2(new_n984), .ZN(new_n997));
  NAND3_X1  g572(.A1(new_n994), .A2(new_n996), .A3(new_n997), .ZN(new_n998));
  XOR2_X1   g573(.A(new_n998), .B(KEYINPUT47), .Z(new_n999));
  AND2_X1   g574(.A1(new_n819), .A2(new_n821), .ZN(new_n1000));
  OAI21_X1  g575(.A(new_n981), .B1(new_n1000), .B2(new_n988), .ZN(new_n1001));
  AND2_X1   g576(.A1(new_n987), .A2(new_n1001), .ZN(new_n1002));
  NOR3_X1   g577(.A1(new_n990), .A2(G1986), .A3(G290), .ZN(new_n1003));
  XOR2_X1   g578(.A(new_n1003), .B(KEYINPUT48), .Z(new_n1004));
  AOI211_X1 g579(.A(new_n991), .B(new_n999), .C1(new_n1002), .C2(new_n1004), .ZN(new_n1005));
  INV_X1    g580(.A(G1981), .ZN(new_n1006));
  INV_X1    g581(.A(KEYINPUT114), .ZN(new_n1007));
  AOI21_X1  g582(.A(new_n1006), .B1(new_n596), .B2(new_n1007), .ZN(new_n1008));
  XNOR2_X1  g583(.A(new_n1008), .B(G305), .ZN(new_n1009));
  XNOR2_X1  g584(.A(new_n1009), .B(KEYINPUT115), .ZN(new_n1010));
  XOR2_X1   g585(.A(KEYINPUT116), .B(KEYINPUT49), .Z(new_n1011));
  NAND2_X1  g586(.A1(new_n1010), .A2(new_n1011), .ZN(new_n1012));
  INV_X1    g587(.A(KEYINPUT117), .ZN(new_n1013));
  NAND2_X1  g588(.A1(new_n1012), .A2(new_n1013), .ZN(new_n1014));
  NAND3_X1  g589(.A1(new_n1010), .A2(KEYINPUT117), .A3(new_n1011), .ZN(new_n1015));
  NAND2_X1  g590(.A1(new_n1014), .A2(new_n1015), .ZN(new_n1016));
  INV_X1    g591(.A(G1384), .ZN(new_n1017));
  INV_X1    g592(.A(new_n980), .ZN(new_n1018));
  NAND3_X1  g593(.A1(new_n865), .A2(new_n1017), .A3(new_n1018), .ZN(new_n1019));
  XOR2_X1   g594(.A(KEYINPUT113), .B(G8), .Z(new_n1020));
  INV_X1    g595(.A(new_n1020), .ZN(new_n1021));
  NAND2_X1  g596(.A1(new_n1019), .A2(new_n1021), .ZN(new_n1022));
  INV_X1    g597(.A(new_n1009), .ZN(new_n1023));
  AOI21_X1  g598(.A(new_n1022), .B1(new_n1023), .B2(KEYINPUT49), .ZN(new_n1024));
  NAND2_X1  g599(.A1(new_n1016), .A2(new_n1024), .ZN(new_n1025));
  INV_X1    g600(.A(G1976), .ZN(new_n1026));
  OAI211_X1 g601(.A(new_n1019), .B(new_n1021), .C1(new_n1026), .C2(G288), .ZN(new_n1027));
  AOI21_X1  g602(.A(KEYINPUT52), .B1(G288), .B2(new_n1026), .ZN(new_n1028));
  INV_X1    g603(.A(new_n1028), .ZN(new_n1029));
  NOR2_X1   g604(.A1(new_n1027), .A2(new_n1029), .ZN(new_n1030));
  AOI21_X1  g605(.A(new_n1030), .B1(KEYINPUT52), .B2(new_n1027), .ZN(new_n1031));
  INV_X1    g606(.A(G8), .ZN(new_n1032));
  INV_X1    g607(.A(KEYINPUT111), .ZN(new_n1033));
  INV_X1    g608(.A(new_n479), .ZN(new_n1034));
  AOI21_X1  g609(.A(G1384), .B1(new_n975), .B2(new_n1034), .ZN(new_n1035));
  INV_X1    g610(.A(KEYINPUT50), .ZN(new_n1036));
  OAI21_X1  g611(.A(new_n1033), .B1(new_n1035), .B2(new_n1036), .ZN(new_n1037));
  OAI211_X1 g612(.A(KEYINPUT111), .B(KEYINPUT50), .C1(G164), .C2(G1384), .ZN(new_n1038));
  NAND2_X1  g613(.A1(new_n1037), .A2(new_n1038), .ZN(new_n1039));
  NAND3_X1  g614(.A1(new_n865), .A2(new_n1036), .A3(new_n1017), .ZN(new_n1040));
  NAND3_X1  g615(.A1(new_n1039), .A2(new_n1018), .A3(new_n1040), .ZN(new_n1041));
  XNOR2_X1  g616(.A(KEYINPUT112), .B(G2090), .ZN(new_n1042));
  OR2_X1    g617(.A1(new_n1041), .A2(new_n1042), .ZN(new_n1043));
  NAND2_X1  g618(.A1(new_n975), .A2(new_n1034), .ZN(new_n1044));
  NAND2_X1  g619(.A1(new_n1044), .A2(new_n1017), .ZN(new_n1045));
  INV_X1    g620(.A(KEYINPUT45), .ZN(new_n1046));
  AOI21_X1  g621(.A(new_n980), .B1(new_n1045), .B2(new_n1046), .ZN(new_n1047));
  NAND2_X1  g622(.A1(new_n865), .A2(new_n1017), .ZN(new_n1048));
  OAI21_X1  g623(.A(new_n1047), .B1(new_n1048), .B2(new_n1046), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n1049), .A2(new_n799), .ZN(new_n1050));
  AOI21_X1  g625(.A(new_n1032), .B1(new_n1043), .B2(new_n1050), .ZN(new_n1051));
  INV_X1    g626(.A(new_n1051), .ZN(new_n1052));
  NAND2_X1  g627(.A1(G303), .A2(G8), .ZN(new_n1053));
  XNOR2_X1  g628(.A(new_n1053), .B(KEYINPUT55), .ZN(new_n1054));
  NAND2_X1  g629(.A1(new_n1052), .A2(new_n1054), .ZN(new_n1055));
  INV_X1    g630(.A(KEYINPUT63), .ZN(new_n1056));
  INV_X1    g631(.A(new_n1054), .ZN(new_n1057));
  AOI21_X1  g632(.A(new_n1056), .B1(new_n1057), .B2(new_n1051), .ZN(new_n1058));
  NAND4_X1  g633(.A1(new_n1025), .A2(new_n1031), .A3(new_n1055), .A4(new_n1058), .ZN(new_n1059));
  NOR2_X1   g634(.A1(new_n1045), .A2(new_n1046), .ZN(new_n1060));
  AOI21_X1  g635(.A(new_n980), .B1(new_n1048), .B2(new_n1046), .ZN(new_n1061));
  INV_X1    g636(.A(KEYINPUT120), .ZN(new_n1062));
  AOI21_X1  g637(.A(new_n1060), .B1(new_n1061), .B2(new_n1062), .ZN(new_n1063));
  AOI21_X1  g638(.A(KEYINPUT45), .B1(new_n865), .B2(new_n1017), .ZN(new_n1064));
  OAI21_X1  g639(.A(KEYINPUT120), .B1(new_n1064), .B2(new_n980), .ZN(new_n1065));
  AOI21_X1  g640(.A(G1966), .B1(new_n1063), .B2(new_n1065), .ZN(new_n1066));
  AND4_X1   g641(.A1(new_n737), .A2(new_n1039), .A3(new_n1018), .A4(new_n1040), .ZN(new_n1067));
  OAI21_X1  g642(.A(new_n1021), .B1(new_n1066), .B2(new_n1067), .ZN(new_n1068));
  NOR2_X1   g643(.A1(new_n1068), .A2(G286), .ZN(new_n1069));
  INV_X1    g644(.A(new_n1069), .ZN(new_n1070));
  OAI21_X1  g645(.A(KEYINPUT63), .B1(new_n1059), .B2(new_n1070), .ZN(new_n1071));
  INV_X1    g646(.A(new_n1024), .ZN(new_n1072));
  AOI21_X1  g647(.A(new_n1072), .B1(new_n1014), .B2(new_n1015), .ZN(new_n1073));
  NAND2_X1  g648(.A1(new_n589), .A2(new_n1026), .ZN(new_n1074));
  OAI22_X1  g649(.A1(new_n1073), .A2(new_n1074), .B1(G1981), .B2(G305), .ZN(new_n1075));
  XNOR2_X1  g650(.A(new_n1022), .B(KEYINPUT118), .ZN(new_n1076));
  INV_X1    g651(.A(new_n1031), .ZN(new_n1077));
  NOR2_X1   g652(.A1(new_n1073), .A2(new_n1077), .ZN(new_n1078));
  NOR2_X1   g653(.A1(new_n1052), .A2(new_n1054), .ZN(new_n1079));
  AOI22_X1  g654(.A1(new_n1075), .A2(new_n1076), .B1(new_n1078), .B2(new_n1079), .ZN(new_n1080));
  NAND2_X1  g655(.A1(new_n1071), .A2(new_n1080), .ZN(new_n1081));
  NAND2_X1  g656(.A1(G286), .A2(new_n1021), .ZN(new_n1082));
  OAI211_X1 g657(.A(new_n1062), .B(new_n1018), .C1(new_n979), .C2(KEYINPUT45), .ZN(new_n1083));
  INV_X1    g658(.A(new_n1060), .ZN(new_n1084));
  NAND3_X1  g659(.A1(new_n1065), .A2(new_n1083), .A3(new_n1084), .ZN(new_n1085));
  AOI21_X1  g660(.A(new_n1067), .B1(new_n1085), .B2(new_n775), .ZN(new_n1086));
  OAI21_X1  g661(.A(new_n1082), .B1(new_n1086), .B2(new_n1032), .ZN(new_n1087));
  OAI211_X1 g662(.A(G286), .B(new_n1021), .C1(new_n1066), .C2(new_n1067), .ZN(new_n1088));
  XNOR2_X1  g663(.A(KEYINPUT124), .B(KEYINPUT51), .ZN(new_n1089));
  NAND3_X1  g664(.A1(new_n1087), .A2(new_n1088), .A3(new_n1089), .ZN(new_n1090));
  INV_X1    g665(.A(KEYINPUT51), .ZN(new_n1091));
  NAND3_X1  g666(.A1(new_n1068), .A2(new_n1091), .A3(new_n1082), .ZN(new_n1092));
  NAND2_X1  g667(.A1(new_n1090), .A2(new_n1092), .ZN(new_n1093));
  INV_X1    g668(.A(KEYINPUT62), .ZN(new_n1094));
  NAND2_X1  g669(.A1(new_n1093), .A2(new_n1094), .ZN(new_n1095));
  NAND3_X1  g670(.A1(new_n1090), .A2(KEYINPUT62), .A3(new_n1092), .ZN(new_n1096));
  INV_X1    g671(.A(KEYINPUT53), .ZN(new_n1097));
  NOR2_X1   g672(.A1(new_n1097), .A2(G2078), .ZN(new_n1098));
  INV_X1    g673(.A(new_n1098), .ZN(new_n1099));
  NOR2_X1   g674(.A1(new_n1085), .A2(new_n1099), .ZN(new_n1100));
  OAI21_X1  g675(.A(new_n1097), .B1(new_n1049), .B2(G2078), .ZN(new_n1101));
  INV_X1    g676(.A(G1961), .ZN(new_n1102));
  NAND2_X1  g677(.A1(new_n1041), .A2(new_n1102), .ZN(new_n1103));
  NAND2_X1  g678(.A1(new_n1101), .A2(new_n1103), .ZN(new_n1104));
  OAI22_X1  g679(.A1(new_n1100), .A2(new_n1104), .B1(new_n579), .B2(new_n580), .ZN(new_n1105));
  INV_X1    g680(.A(new_n1105), .ZN(new_n1106));
  NAND3_X1  g681(.A1(new_n1095), .A2(new_n1096), .A3(new_n1106), .ZN(new_n1107));
  NAND2_X1  g682(.A1(new_n1059), .A2(new_n1069), .ZN(new_n1108));
  INV_X1    g683(.A(G1956), .ZN(new_n1109));
  AOI21_X1  g684(.A(new_n1036), .B1(new_n865), .B2(new_n1017), .ZN(new_n1110));
  OAI21_X1  g685(.A(new_n1018), .B1(new_n1045), .B2(KEYINPUT50), .ZN(new_n1111));
  OAI21_X1  g686(.A(new_n1109), .B1(new_n1110), .B2(new_n1111), .ZN(new_n1112));
  XNOR2_X1  g687(.A(KEYINPUT56), .B(G2072), .ZN(new_n1113));
  XNOR2_X1  g688(.A(new_n1113), .B(KEYINPUT121), .ZN(new_n1114));
  OAI211_X1 g689(.A(new_n1047), .B(new_n1114), .C1(new_n1048), .C2(new_n1046), .ZN(new_n1115));
  NAND2_X1  g690(.A1(new_n884), .A2(new_n885), .ZN(new_n1116));
  INV_X1    g691(.A(KEYINPUT57), .ZN(new_n1117));
  XNOR2_X1  g692(.A(new_n1116), .B(new_n1117), .ZN(new_n1118));
  NAND3_X1  g693(.A1(new_n1112), .A2(new_n1115), .A3(new_n1118), .ZN(new_n1119));
  XNOR2_X1  g694(.A(new_n1119), .B(KEYINPUT122), .ZN(new_n1120));
  NAND2_X1  g695(.A1(new_n1041), .A2(new_n714), .ZN(new_n1121));
  NOR2_X1   g696(.A1(new_n1019), .A2(G2067), .ZN(new_n1122));
  INV_X1    g697(.A(new_n1122), .ZN(new_n1123));
  AOI21_X1  g698(.A(new_n614), .B1(new_n1121), .B2(new_n1123), .ZN(new_n1124));
  NAND2_X1  g699(.A1(new_n1112), .A2(new_n1115), .ZN(new_n1125));
  INV_X1    g700(.A(new_n1118), .ZN(new_n1126));
  NAND2_X1  g701(.A1(new_n1125), .A2(new_n1126), .ZN(new_n1127));
  INV_X1    g702(.A(new_n1127), .ZN(new_n1128));
  OAI21_X1  g703(.A(new_n1120), .B1(new_n1124), .B2(new_n1128), .ZN(new_n1129));
  AOI211_X1 g704(.A(new_n622), .B(new_n1122), .C1(new_n1041), .C2(new_n714), .ZN(new_n1130));
  OAI21_X1  g705(.A(KEYINPUT60), .B1(new_n1130), .B2(new_n1124), .ZN(new_n1131));
  OAI211_X1 g706(.A(new_n1047), .B(new_n992), .C1(new_n1048), .C2(new_n1046), .ZN(new_n1132));
  XOR2_X1   g707(.A(KEYINPUT58), .B(G1341), .Z(new_n1133));
  NAND2_X1  g708(.A1(new_n1019), .A2(new_n1133), .ZN(new_n1134));
  AOI21_X1  g709(.A(new_n552), .B1(new_n1132), .B2(new_n1134), .ZN(new_n1135));
  INV_X1    g710(.A(KEYINPUT59), .ZN(new_n1136));
  XNOR2_X1  g711(.A(new_n1135), .B(new_n1136), .ZN(new_n1137));
  NAND3_X1  g712(.A1(new_n1127), .A2(KEYINPUT61), .A3(new_n1119), .ZN(new_n1138));
  NOR2_X1   g713(.A1(new_n614), .A2(KEYINPUT60), .ZN(new_n1139));
  NAND3_X1  g714(.A1(new_n1121), .A2(new_n1123), .A3(new_n1139), .ZN(new_n1140));
  NAND4_X1  g715(.A1(new_n1131), .A2(new_n1137), .A3(new_n1138), .A4(new_n1140), .ZN(new_n1141));
  AOI21_X1  g716(.A(KEYINPUT123), .B1(new_n1125), .B2(new_n1126), .ZN(new_n1142));
  INV_X1    g717(.A(KEYINPUT123), .ZN(new_n1143));
  AOI211_X1 g718(.A(new_n1143), .B(new_n1118), .C1(new_n1112), .C2(new_n1115), .ZN(new_n1144));
  NOR2_X1   g719(.A1(new_n1142), .A2(new_n1144), .ZN(new_n1145));
  AOI21_X1  g720(.A(KEYINPUT61), .B1(new_n1145), .B2(new_n1120), .ZN(new_n1146));
  OAI21_X1  g721(.A(new_n1129), .B1(new_n1141), .B2(new_n1146), .ZN(new_n1147));
  AND2_X1   g722(.A1(new_n1090), .A2(new_n1092), .ZN(new_n1148));
  AND2_X1   g723(.A1(new_n1101), .A2(new_n1103), .ZN(new_n1149));
  INV_X1    g724(.A(KEYINPUT125), .ZN(new_n1150));
  OAI211_X1 g725(.A(new_n1061), .B(new_n1098), .C1(new_n1046), .C2(new_n1048), .ZN(new_n1151));
  NAND4_X1  g726(.A1(new_n1149), .A2(new_n1150), .A3(G301), .A4(new_n1151), .ZN(new_n1152));
  NAND4_X1  g727(.A1(new_n1151), .A2(new_n1101), .A3(new_n1103), .A4(G301), .ZN(new_n1153));
  NAND2_X1  g728(.A1(new_n1153), .A2(KEYINPUT125), .ZN(new_n1154));
  NAND3_X1  g729(.A1(new_n1105), .A2(new_n1152), .A3(new_n1154), .ZN(new_n1155));
  INV_X1    g730(.A(KEYINPUT54), .ZN(new_n1156));
  NAND2_X1  g731(.A1(new_n1149), .A2(new_n1151), .ZN(new_n1157));
  AOI21_X1  g732(.A(new_n1156), .B1(new_n1157), .B2(G171), .ZN(new_n1158));
  OAI211_X1 g733(.A(new_n1149), .B(G301), .C1(new_n1085), .C2(new_n1099), .ZN(new_n1159));
  AOI22_X1  g734(.A1(new_n1155), .A2(new_n1156), .B1(new_n1158), .B2(new_n1159), .ZN(new_n1160));
  NAND3_X1  g735(.A1(new_n1147), .A2(new_n1148), .A3(new_n1160), .ZN(new_n1161));
  NAND3_X1  g736(.A1(new_n1107), .A2(new_n1108), .A3(new_n1161), .ZN(new_n1162));
  INV_X1    g737(.A(new_n1050), .ZN(new_n1163));
  NOR3_X1   g738(.A1(new_n1110), .A2(new_n1111), .A3(new_n1042), .ZN(new_n1164));
  OAI21_X1  g739(.A(new_n1021), .B1(new_n1163), .B2(new_n1164), .ZN(new_n1165));
  NAND2_X1  g740(.A1(new_n1054), .A2(new_n1165), .ZN(new_n1166));
  OAI21_X1  g741(.A(new_n1166), .B1(new_n1052), .B2(new_n1054), .ZN(new_n1167));
  OR2_X1    g742(.A1(new_n1078), .A2(KEYINPUT119), .ZN(new_n1168));
  NAND2_X1  g743(.A1(new_n1078), .A2(KEYINPUT119), .ZN(new_n1169));
  AOI21_X1  g744(.A(new_n1167), .B1(new_n1168), .B2(new_n1169), .ZN(new_n1170));
  AOI21_X1  g745(.A(new_n1081), .B1(new_n1162), .B2(new_n1170), .ZN(new_n1171));
  XNOR2_X1  g746(.A(new_n603), .B(G1986), .ZN(new_n1172));
  OAI21_X1  g747(.A(new_n1002), .B1(new_n990), .B2(new_n1172), .ZN(new_n1173));
  OAI21_X1  g748(.A(new_n1005), .B1(new_n1171), .B2(new_n1173), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g749(.A(G319), .ZN(new_n1176));
  NOR3_X1   g750(.A1(G401), .A2(new_n1176), .A3(G227), .ZN(new_n1177));
  AND4_X1   g751(.A1(new_n700), .A2(new_n699), .A3(new_n880), .A4(new_n1177), .ZN(new_n1178));
  NAND2_X1  g752(.A1(new_n1178), .A2(new_n969), .ZN(G225));
  INV_X1    g753(.A(G225), .ZN(G308));
endmodule


