//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 0 0 1 0 0 0 1 0 0 1 0 0 0 1 0 1 1 0 1 1 1 1 0 0 1 0 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 0 0 0 0 0 0 0 1 1 1 0 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:19:48 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n674, new_n675, new_n676, new_n677, new_n678,
    new_n679, new_n680, new_n681, new_n682, new_n683, new_n685, new_n686,
    new_n687, new_n688, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n724,
    new_n725, new_n726, new_n727, new_n728, new_n729, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n751, new_n752, new_n753, new_n754, new_n756,
    new_n757, new_n758, new_n759, new_n761, new_n762, new_n763, new_n764,
    new_n765, new_n767, new_n769, new_n770, new_n771, new_n772, new_n773,
    new_n774, new_n775, new_n776, new_n777, new_n778, new_n779, new_n780,
    new_n781, new_n782, new_n783, new_n784, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n796,
    new_n797, new_n798, new_n799, new_n800, new_n801, new_n802, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n844, new_n845, new_n846, new_n848, new_n849,
    new_n850, new_n851, new_n853, new_n854, new_n855, new_n856, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n895,
    new_n896, new_n897, new_n899, new_n900, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n912,
    new_n913, new_n915, new_n916, new_n917, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n940, new_n941, new_n942, new_n943, new_n945, new_n946;
  XNOR2_X1  g000(.A(G78gat), .B(G106gat), .ZN(new_n202));
  XNOR2_X1  g001(.A(new_n202), .B(G22gat), .ZN(new_n203));
  INV_X1    g002(.A(new_n203), .ZN(new_n204));
  INV_X1    g003(.A(G228gat), .ZN(new_n205));
  INV_X1    g004(.A(G233gat), .ZN(new_n206));
  NOR2_X1   g005(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  XNOR2_X1  g006(.A(G197gat), .B(G204gat), .ZN(new_n208));
  INV_X1    g007(.A(KEYINPUT22), .ZN(new_n209));
  INV_X1    g008(.A(G211gat), .ZN(new_n210));
  INV_X1    g009(.A(G218gat), .ZN(new_n211));
  OAI21_X1  g010(.A(new_n209), .B1(new_n210), .B2(new_n211), .ZN(new_n212));
  NAND2_X1  g011(.A1(new_n208), .A2(new_n212), .ZN(new_n213));
  XNOR2_X1  g012(.A(G211gat), .B(G218gat), .ZN(new_n214));
  INV_X1    g013(.A(new_n214), .ZN(new_n215));
  NAND2_X1  g014(.A1(new_n213), .A2(new_n215), .ZN(new_n216));
  NAND3_X1  g015(.A1(new_n214), .A2(new_n208), .A3(new_n212), .ZN(new_n217));
  NAND2_X1  g016(.A1(new_n216), .A2(new_n217), .ZN(new_n218));
  INV_X1    g017(.A(G141gat), .ZN(new_n219));
  NAND2_X1  g018(.A1(new_n219), .A2(G148gat), .ZN(new_n220));
  INV_X1    g019(.A(G148gat), .ZN(new_n221));
  NAND2_X1  g020(.A1(new_n221), .A2(G141gat), .ZN(new_n222));
  NAND2_X1  g021(.A1(new_n220), .A2(new_n222), .ZN(new_n223));
  XNOR2_X1  g022(.A(KEYINPUT73), .B(KEYINPUT2), .ZN(new_n224));
  INV_X1    g023(.A(G162gat), .ZN(new_n225));
  NAND2_X1  g024(.A1(new_n225), .A2(G155gat), .ZN(new_n226));
  INV_X1    g025(.A(G155gat), .ZN(new_n227));
  NAND2_X1  g026(.A1(new_n227), .A2(G162gat), .ZN(new_n228));
  AOI22_X1  g027(.A1(new_n223), .A2(new_n224), .B1(new_n226), .B2(new_n228), .ZN(new_n229));
  INV_X1    g028(.A(new_n229), .ZN(new_n230));
  INV_X1    g029(.A(KEYINPUT2), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n227), .A2(KEYINPUT76), .ZN(new_n232));
  INV_X1    g031(.A(KEYINPUT76), .ZN(new_n233));
  NAND2_X1  g032(.A1(new_n233), .A2(G155gat), .ZN(new_n234));
  NAND2_X1  g033(.A1(new_n232), .A2(new_n234), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n225), .A2(KEYINPUT77), .ZN(new_n236));
  INV_X1    g035(.A(KEYINPUT77), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n237), .A2(G162gat), .ZN(new_n238));
  NAND2_X1  g037(.A1(new_n236), .A2(new_n238), .ZN(new_n239));
  AOI21_X1  g038(.A(new_n231), .B1(new_n235), .B2(new_n239), .ZN(new_n240));
  OAI21_X1  g039(.A(KEYINPUT74), .B1(new_n221), .B2(G141gat), .ZN(new_n241));
  INV_X1    g040(.A(KEYINPUT74), .ZN(new_n242));
  NAND3_X1  g041(.A1(new_n242), .A2(new_n219), .A3(G148gat), .ZN(new_n243));
  NAND3_X1  g042(.A1(new_n241), .A2(new_n243), .A3(new_n222), .ZN(new_n244));
  INV_X1    g043(.A(new_n244), .ZN(new_n245));
  NOR2_X1   g044(.A1(new_n240), .A2(new_n245), .ZN(new_n246));
  INV_X1    g045(.A(KEYINPUT75), .ZN(new_n247));
  NOR2_X1   g046(.A1(new_n227), .A2(G162gat), .ZN(new_n248));
  NOR2_X1   g047(.A1(new_n225), .A2(G155gat), .ZN(new_n249));
  OAI21_X1  g048(.A(new_n247), .B1(new_n248), .B2(new_n249), .ZN(new_n250));
  NAND3_X1  g049(.A1(new_n226), .A2(new_n228), .A3(KEYINPUT75), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n250), .A2(new_n251), .ZN(new_n252));
  AOI21_X1  g051(.A(KEYINPUT78), .B1(new_n246), .B2(new_n252), .ZN(new_n253));
  XNOR2_X1  g052(.A(KEYINPUT76), .B(G155gat), .ZN(new_n254));
  XNOR2_X1  g053(.A(KEYINPUT77), .B(G162gat), .ZN(new_n255));
  OAI21_X1  g054(.A(KEYINPUT2), .B1(new_n254), .B2(new_n255), .ZN(new_n256));
  NAND4_X1  g055(.A1(new_n252), .A2(new_n256), .A3(KEYINPUT78), .A4(new_n244), .ZN(new_n257));
  INV_X1    g056(.A(new_n257), .ZN(new_n258));
  OAI21_X1  g057(.A(new_n230), .B1(new_n253), .B2(new_n258), .ZN(new_n259));
  OAI21_X1  g058(.A(KEYINPUT79), .B1(new_n259), .B2(KEYINPUT3), .ZN(new_n260));
  NAND3_X1  g059(.A1(new_n252), .A2(new_n256), .A3(new_n244), .ZN(new_n261));
  INV_X1    g060(.A(KEYINPUT78), .ZN(new_n262));
  NAND2_X1  g061(.A1(new_n261), .A2(new_n262), .ZN(new_n263));
  AOI21_X1  g062(.A(new_n229), .B1(new_n263), .B2(new_n257), .ZN(new_n264));
  INV_X1    g063(.A(KEYINPUT79), .ZN(new_n265));
  INV_X1    g064(.A(KEYINPUT3), .ZN(new_n266));
  NAND3_X1  g065(.A1(new_n264), .A2(new_n265), .A3(new_n266), .ZN(new_n267));
  NAND2_X1  g066(.A1(new_n260), .A2(new_n267), .ZN(new_n268));
  INV_X1    g067(.A(KEYINPUT29), .ZN(new_n269));
  AOI21_X1  g068(.A(new_n218), .B1(new_n268), .B2(new_n269), .ZN(new_n270));
  INV_X1    g069(.A(new_n218), .ZN(new_n271));
  OAI21_X1  g070(.A(new_n266), .B1(new_n271), .B2(KEYINPUT29), .ZN(new_n272));
  NAND2_X1  g071(.A1(new_n259), .A2(new_n272), .ZN(new_n273));
  INV_X1    g072(.A(new_n273), .ZN(new_n274));
  OAI21_X1  g073(.A(new_n207), .B1(new_n270), .B2(new_n274), .ZN(new_n275));
  NAND2_X1  g074(.A1(new_n263), .A2(new_n257), .ZN(new_n276));
  AND4_X1   g075(.A1(new_n265), .A2(new_n276), .A3(new_n266), .A4(new_n230), .ZN(new_n277));
  AOI21_X1  g076(.A(new_n265), .B1(new_n264), .B2(new_n266), .ZN(new_n278));
  OAI21_X1  g077(.A(new_n269), .B1(new_n277), .B2(new_n278), .ZN(new_n279));
  NAND2_X1  g078(.A1(new_n279), .A2(new_n271), .ZN(new_n280));
  NAND3_X1  g079(.A1(new_n216), .A2(KEYINPUT84), .A3(new_n217), .ZN(new_n281));
  INV_X1    g080(.A(KEYINPUT84), .ZN(new_n282));
  NAND3_X1  g081(.A1(new_n213), .A2(new_n282), .A3(new_n215), .ZN(new_n283));
  NAND3_X1  g082(.A1(new_n281), .A2(new_n269), .A3(new_n283), .ZN(new_n284));
  INV_X1    g083(.A(KEYINPUT85), .ZN(new_n285));
  NAND2_X1  g084(.A1(new_n284), .A2(new_n285), .ZN(new_n286));
  NAND4_X1  g085(.A1(new_n281), .A2(KEYINPUT85), .A3(new_n269), .A4(new_n283), .ZN(new_n287));
  NAND3_X1  g086(.A1(new_n286), .A2(new_n266), .A3(new_n287), .ZN(new_n288));
  NAND2_X1  g087(.A1(new_n288), .A2(new_n259), .ZN(new_n289));
  NAND2_X1  g088(.A1(new_n289), .A2(KEYINPUT86), .ZN(new_n290));
  INV_X1    g089(.A(KEYINPUT86), .ZN(new_n291));
  NAND3_X1  g090(.A1(new_n288), .A2(new_n291), .A3(new_n259), .ZN(new_n292));
  NAND2_X1  g091(.A1(new_n290), .A2(new_n292), .ZN(new_n293));
  INV_X1    g092(.A(new_n207), .ZN(new_n294));
  NAND3_X1  g093(.A1(new_n280), .A2(new_n293), .A3(new_n294), .ZN(new_n295));
  XNOR2_X1  g094(.A(KEYINPUT31), .B(G50gat), .ZN(new_n296));
  INV_X1    g095(.A(new_n296), .ZN(new_n297));
  AND3_X1   g096(.A1(new_n275), .A2(new_n295), .A3(new_n297), .ZN(new_n298));
  AOI21_X1  g097(.A(new_n297), .B1(new_n275), .B2(new_n295), .ZN(new_n299));
  OAI21_X1  g098(.A(new_n204), .B1(new_n298), .B2(new_n299), .ZN(new_n300));
  INV_X1    g099(.A(new_n292), .ZN(new_n301));
  AOI21_X1  g100(.A(new_n291), .B1(new_n288), .B2(new_n259), .ZN(new_n302));
  OAI21_X1  g101(.A(new_n294), .B1(new_n301), .B2(new_n302), .ZN(new_n303));
  NOR2_X1   g102(.A1(new_n303), .A2(new_n270), .ZN(new_n304));
  AOI21_X1  g103(.A(new_n294), .B1(new_n280), .B2(new_n273), .ZN(new_n305));
  OAI21_X1  g104(.A(new_n296), .B1(new_n304), .B2(new_n305), .ZN(new_n306));
  NAND3_X1  g105(.A1(new_n275), .A2(new_n295), .A3(new_n297), .ZN(new_n307));
  NAND3_X1  g106(.A1(new_n306), .A2(new_n203), .A3(new_n307), .ZN(new_n308));
  NAND2_X1  g107(.A1(new_n300), .A2(new_n308), .ZN(new_n309));
  INV_X1    g108(.A(new_n309), .ZN(new_n310));
  INV_X1    g109(.A(G113gat), .ZN(new_n311));
  INV_X1    g110(.A(G120gat), .ZN(new_n312));
  AOI21_X1  g111(.A(KEYINPUT1), .B1(new_n311), .B2(new_n312), .ZN(new_n313));
  XNOR2_X1  g112(.A(G127gat), .B(G134gat), .ZN(new_n314));
  XOR2_X1   g113(.A(KEYINPUT68), .B(G120gat), .Z(new_n315));
  OAI211_X1 g114(.A(new_n313), .B(new_n314), .C1(new_n315), .C2(new_n311), .ZN(new_n316));
  OAI21_X1  g115(.A(new_n313), .B1(new_n311), .B2(new_n312), .ZN(new_n317));
  INV_X1    g116(.A(new_n314), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n317), .A2(new_n318), .ZN(new_n319));
  NAND2_X1  g118(.A1(new_n316), .A2(new_n319), .ZN(new_n320));
  INV_X1    g119(.A(new_n320), .ZN(new_n321));
  OAI211_X1 g120(.A(new_n230), .B(new_n321), .C1(new_n253), .C2(new_n258), .ZN(new_n322));
  INV_X1    g121(.A(KEYINPUT4), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n322), .A2(new_n323), .ZN(new_n324));
  INV_X1    g123(.A(new_n324), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n322), .A2(KEYINPUT80), .ZN(new_n326));
  INV_X1    g125(.A(KEYINPUT80), .ZN(new_n327));
  NAND3_X1  g126(.A1(new_n264), .A2(new_n327), .A3(new_n321), .ZN(new_n328));
  NAND2_X1  g127(.A1(new_n326), .A2(new_n328), .ZN(new_n329));
  AOI21_X1  g128(.A(new_n325), .B1(new_n329), .B2(KEYINPUT4), .ZN(new_n330));
  INV_X1    g129(.A(new_n330), .ZN(new_n331));
  AOI21_X1  g130(.A(new_n321), .B1(new_n259), .B2(KEYINPUT3), .ZN(new_n332));
  OAI21_X1  g131(.A(new_n332), .B1(new_n277), .B2(new_n278), .ZN(new_n333));
  NAND2_X1  g132(.A1(G225gat), .A2(G233gat), .ZN(new_n334));
  XOR2_X1   g133(.A(KEYINPUT81), .B(KEYINPUT5), .Z(new_n335));
  NAND3_X1  g134(.A1(new_n333), .A2(new_n334), .A3(new_n335), .ZN(new_n336));
  OR2_X1    g135(.A1(new_n331), .A2(new_n336), .ZN(new_n337));
  NAND3_X1  g136(.A1(new_n264), .A2(KEYINPUT4), .A3(new_n321), .ZN(new_n338));
  NAND3_X1  g137(.A1(new_n326), .A2(new_n323), .A3(new_n328), .ZN(new_n339));
  NAND4_X1  g138(.A1(new_n333), .A2(new_n334), .A3(new_n338), .A4(new_n339), .ZN(new_n340));
  INV_X1    g139(.A(KEYINPUT82), .ZN(new_n341));
  NAND2_X1  g140(.A1(new_n259), .A2(new_n320), .ZN(new_n342));
  NAND3_X1  g141(.A1(new_n326), .A2(new_n328), .A3(new_n342), .ZN(new_n343));
  INV_X1    g142(.A(new_n334), .ZN(new_n344));
  AOI21_X1  g143(.A(new_n335), .B1(new_n343), .B2(new_n344), .ZN(new_n345));
  AND3_X1   g144(.A1(new_n340), .A2(new_n341), .A3(new_n345), .ZN(new_n346));
  AOI21_X1  g145(.A(new_n341), .B1(new_n340), .B2(new_n345), .ZN(new_n347));
  OAI21_X1  g146(.A(new_n337), .B1(new_n346), .B2(new_n347), .ZN(new_n348));
  XNOR2_X1  g147(.A(G1gat), .B(G29gat), .ZN(new_n349));
  XNOR2_X1  g148(.A(new_n349), .B(KEYINPUT0), .ZN(new_n350));
  XNOR2_X1  g149(.A(G57gat), .B(G85gat), .ZN(new_n351));
  XOR2_X1   g150(.A(new_n350), .B(new_n351), .Z(new_n352));
  INV_X1    g151(.A(new_n352), .ZN(new_n353));
  XNOR2_X1  g152(.A(KEYINPUT83), .B(KEYINPUT6), .ZN(new_n354));
  INV_X1    g153(.A(new_n354), .ZN(new_n355));
  NAND3_X1  g154(.A1(new_n348), .A2(new_n353), .A3(new_n355), .ZN(new_n356));
  NOR2_X1   g155(.A1(new_n331), .A2(new_n336), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n340), .A2(new_n345), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n358), .A2(KEYINPUT82), .ZN(new_n359));
  NAND3_X1  g158(.A1(new_n340), .A2(new_n341), .A3(new_n345), .ZN(new_n360));
  AOI21_X1  g159(.A(new_n357), .B1(new_n359), .B2(new_n360), .ZN(new_n361));
  OAI21_X1  g160(.A(new_n354), .B1(new_n361), .B2(new_n352), .ZN(new_n362));
  OAI211_X1 g161(.A(new_n352), .B(new_n337), .C1(new_n346), .C2(new_n347), .ZN(new_n363));
  INV_X1    g162(.A(new_n363), .ZN(new_n364));
  OAI21_X1  g163(.A(new_n356), .B1(new_n362), .B2(new_n364), .ZN(new_n365));
  XOR2_X1   g164(.A(G8gat), .B(G36gat), .Z(new_n366));
  XNOR2_X1  g165(.A(new_n366), .B(KEYINPUT72), .ZN(new_n367));
  XNOR2_X1  g166(.A(G64gat), .B(G92gat), .ZN(new_n368));
  XOR2_X1   g167(.A(new_n367), .B(new_n368), .Z(new_n369));
  NAND2_X1  g168(.A1(G183gat), .A2(G190gat), .ZN(new_n370));
  INV_X1    g169(.A(KEYINPUT24), .ZN(new_n371));
  NAND2_X1  g170(.A1(new_n370), .A2(new_n371), .ZN(new_n372));
  OR2_X1    g171(.A1(G183gat), .A2(G190gat), .ZN(new_n373));
  NAND3_X1  g172(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n374));
  NAND3_X1  g173(.A1(new_n372), .A2(new_n373), .A3(new_n374), .ZN(new_n375));
  NOR2_X1   g174(.A1(G169gat), .A2(G176gat), .ZN(new_n376));
  INV_X1    g175(.A(new_n376), .ZN(new_n377));
  NAND2_X1  g176(.A1(G169gat), .A2(G176gat), .ZN(new_n378));
  NAND2_X1  g177(.A1(new_n378), .A2(KEYINPUT23), .ZN(new_n379));
  NAND2_X1  g178(.A1(new_n377), .A2(new_n379), .ZN(new_n380));
  AND3_X1   g179(.A1(new_n376), .A2(KEYINPUT64), .A3(KEYINPUT23), .ZN(new_n381));
  AOI21_X1  g180(.A(KEYINPUT64), .B1(new_n376), .B2(KEYINPUT23), .ZN(new_n382));
  OAI211_X1 g181(.A(new_n375), .B(new_n380), .C1(new_n381), .C2(new_n382), .ZN(new_n383));
  INV_X1    g182(.A(KEYINPUT65), .ZN(new_n384));
  INV_X1    g183(.A(KEYINPUT25), .ZN(new_n385));
  AND3_X1   g184(.A1(new_n383), .A2(new_n384), .A3(new_n385), .ZN(new_n386));
  AOI21_X1  g185(.A(new_n384), .B1(new_n383), .B2(new_n385), .ZN(new_n387));
  NAND2_X1  g186(.A1(new_n373), .A2(new_n374), .ZN(new_n388));
  OR2_X1    g187(.A1(new_n371), .A2(KEYINPUT66), .ZN(new_n389));
  AOI22_X1  g188(.A1(new_n371), .A2(KEYINPUT66), .B1(G183gat), .B2(G190gat), .ZN(new_n390));
  AOI21_X1  g189(.A(new_n388), .B1(new_n389), .B2(new_n390), .ZN(new_n391));
  AOI21_X1  g190(.A(new_n385), .B1(new_n376), .B2(KEYINPUT23), .ZN(new_n392));
  NAND2_X1  g191(.A1(new_n380), .A2(new_n392), .ZN(new_n393));
  NOR2_X1   g192(.A1(new_n391), .A2(new_n393), .ZN(new_n394));
  NOR3_X1   g193(.A1(new_n386), .A2(new_n387), .A3(new_n394), .ZN(new_n395));
  XNOR2_X1  g194(.A(KEYINPUT27), .B(G183gat), .ZN(new_n396));
  INV_X1    g195(.A(G190gat), .ZN(new_n397));
  NAND2_X1  g196(.A1(new_n396), .A2(new_n397), .ZN(new_n398));
  INV_X1    g197(.A(KEYINPUT67), .ZN(new_n399));
  NAND3_X1  g198(.A1(new_n398), .A2(new_n399), .A3(KEYINPUT28), .ZN(new_n400));
  NAND2_X1  g199(.A1(new_n400), .A2(new_n370), .ZN(new_n401));
  XOR2_X1   g200(.A(KEYINPUT67), .B(KEYINPUT28), .Z(new_n402));
  NOR2_X1   g201(.A1(new_n377), .A2(KEYINPUT26), .ZN(new_n403));
  INV_X1    g202(.A(KEYINPUT26), .ZN(new_n404));
  AOI21_X1  g203(.A(new_n376), .B1(new_n404), .B2(new_n378), .ZN(new_n405));
  OAI22_X1  g204(.A1(new_n398), .A2(new_n402), .B1(new_n403), .B2(new_n405), .ZN(new_n406));
  NOR2_X1   g205(.A1(new_n401), .A2(new_n406), .ZN(new_n407));
  OAI21_X1  g206(.A(new_n269), .B1(new_n395), .B2(new_n407), .ZN(new_n408));
  NAND2_X1  g207(.A1(G226gat), .A2(G233gat), .ZN(new_n409));
  NAND2_X1  g208(.A1(new_n408), .A2(new_n409), .ZN(new_n410));
  OAI211_X1 g209(.A(G226gat), .B(G233gat), .C1(new_n395), .C2(new_n407), .ZN(new_n411));
  NAND3_X1  g210(.A1(new_n410), .A2(new_n218), .A3(new_n411), .ZN(new_n412));
  INV_X1    g211(.A(new_n412), .ZN(new_n413));
  AOI21_X1  g212(.A(new_n218), .B1(new_n410), .B2(new_n411), .ZN(new_n414));
  OAI21_X1  g213(.A(new_n369), .B1(new_n413), .B2(new_n414), .ZN(new_n415));
  NAND2_X1  g214(.A1(new_n410), .A2(new_n411), .ZN(new_n416));
  NAND2_X1  g215(.A1(new_n416), .A2(new_n271), .ZN(new_n417));
  INV_X1    g216(.A(new_n369), .ZN(new_n418));
  NAND3_X1  g217(.A1(new_n417), .A2(new_n412), .A3(new_n418), .ZN(new_n419));
  NAND3_X1  g218(.A1(new_n415), .A2(new_n419), .A3(KEYINPUT30), .ZN(new_n420));
  NOR2_X1   g219(.A1(new_n413), .A2(new_n414), .ZN(new_n421));
  INV_X1    g220(.A(KEYINPUT30), .ZN(new_n422));
  NAND3_X1  g221(.A1(new_n421), .A2(new_n422), .A3(new_n418), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n420), .A2(new_n423), .ZN(new_n424));
  AOI21_X1  g223(.A(new_n310), .B1(new_n365), .B2(new_n424), .ZN(new_n425));
  INV_X1    g224(.A(KEYINPUT71), .ZN(new_n426));
  INV_X1    g225(.A(KEYINPUT69), .ZN(new_n427));
  NAND2_X1  g226(.A1(new_n320), .A2(new_n427), .ZN(new_n428));
  NAND2_X1  g227(.A1(new_n321), .A2(KEYINPUT69), .ZN(new_n429));
  OAI211_X1 g228(.A(new_n428), .B(new_n429), .C1(new_n395), .C2(new_n407), .ZN(new_n430));
  INV_X1    g229(.A(G227gat), .ZN(new_n431));
  NOR2_X1   g230(.A1(new_n431), .A2(new_n206), .ZN(new_n432));
  INV_X1    g231(.A(new_n387), .ZN(new_n433));
  NAND3_X1  g232(.A1(new_n383), .A2(new_n384), .A3(new_n385), .ZN(new_n434));
  INV_X1    g233(.A(new_n394), .ZN(new_n435));
  NAND3_X1  g234(.A1(new_n433), .A2(new_n434), .A3(new_n435), .ZN(new_n436));
  INV_X1    g235(.A(new_n407), .ZN(new_n437));
  NAND4_X1  g236(.A1(new_n436), .A2(new_n427), .A3(new_n437), .A4(new_n320), .ZN(new_n438));
  NAND3_X1  g237(.A1(new_n430), .A2(new_n432), .A3(new_n438), .ZN(new_n439));
  INV_X1    g238(.A(KEYINPUT70), .ZN(new_n440));
  NAND2_X1  g239(.A1(new_n439), .A2(new_n440), .ZN(new_n441));
  NAND4_X1  g240(.A1(new_n430), .A2(new_n438), .A3(KEYINPUT70), .A4(new_n432), .ZN(new_n442));
  NAND2_X1  g241(.A1(new_n441), .A2(new_n442), .ZN(new_n443));
  INV_X1    g242(.A(KEYINPUT33), .ZN(new_n444));
  NAND2_X1  g243(.A1(new_n443), .A2(new_n444), .ZN(new_n445));
  AOI21_X1  g244(.A(new_n432), .B1(new_n430), .B2(new_n438), .ZN(new_n446));
  INV_X1    g245(.A(KEYINPUT34), .ZN(new_n447));
  XNOR2_X1  g246(.A(new_n446), .B(new_n447), .ZN(new_n448));
  XOR2_X1   g247(.A(G15gat), .B(G43gat), .Z(new_n449));
  XNOR2_X1  g248(.A(G71gat), .B(G99gat), .ZN(new_n450));
  XNOR2_X1  g249(.A(new_n449), .B(new_n450), .ZN(new_n451));
  NAND3_X1  g250(.A1(new_n445), .A2(new_n448), .A3(new_n451), .ZN(new_n452));
  AND2_X1   g251(.A1(new_n443), .A2(KEYINPUT32), .ZN(new_n453));
  NOR2_X1   g252(.A1(new_n446), .A2(new_n447), .ZN(new_n454));
  AOI211_X1 g253(.A(KEYINPUT34), .B(new_n432), .C1(new_n430), .C2(new_n438), .ZN(new_n455));
  NOR2_X1   g254(.A1(new_n454), .A2(new_n455), .ZN(new_n456));
  AOI21_X1  g255(.A(KEYINPUT33), .B1(new_n441), .B2(new_n442), .ZN(new_n457));
  INV_X1    g256(.A(new_n451), .ZN(new_n458));
  OAI21_X1  g257(.A(new_n456), .B1(new_n457), .B2(new_n458), .ZN(new_n459));
  AND3_X1   g258(.A1(new_n452), .A2(new_n453), .A3(new_n459), .ZN(new_n460));
  AOI21_X1  g259(.A(new_n453), .B1(new_n452), .B2(new_n459), .ZN(new_n461));
  OAI21_X1  g260(.A(new_n426), .B1(new_n460), .B2(new_n461), .ZN(new_n462));
  INV_X1    g261(.A(KEYINPUT36), .ZN(new_n463));
  NAND2_X1  g262(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  OAI211_X1 g263(.A(new_n426), .B(KEYINPUT36), .C1(new_n460), .C2(new_n461), .ZN(new_n465));
  NAND2_X1  g264(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  NOR2_X1   g265(.A1(new_n425), .A2(new_n466), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n330), .A2(new_n333), .ZN(new_n468));
  NAND2_X1  g267(.A1(new_n468), .A2(new_n344), .ZN(new_n469));
  NAND4_X1  g268(.A1(new_n326), .A2(new_n342), .A3(new_n328), .A4(new_n334), .ZN(new_n470));
  XNOR2_X1  g269(.A(new_n470), .B(KEYINPUT87), .ZN(new_n471));
  NAND3_X1  g270(.A1(new_n469), .A2(KEYINPUT39), .A3(new_n471), .ZN(new_n472));
  AOI21_X1  g271(.A(new_n334), .B1(new_n330), .B2(new_n333), .ZN(new_n473));
  INV_X1    g272(.A(KEYINPUT39), .ZN(new_n474));
  AOI21_X1  g273(.A(new_n353), .B1(new_n473), .B2(new_n474), .ZN(new_n475));
  AND3_X1   g274(.A1(new_n472), .A2(new_n475), .A3(KEYINPUT40), .ZN(new_n476));
  AOI21_X1  g275(.A(KEYINPUT40), .B1(new_n472), .B2(new_n475), .ZN(new_n477));
  NOR2_X1   g276(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  AOI21_X1  g277(.A(new_n424), .B1(new_n353), .B2(new_n348), .ZN(new_n479));
  AOI21_X1  g278(.A(new_n309), .B1(new_n478), .B2(new_n479), .ZN(new_n480));
  NAND2_X1  g279(.A1(new_n348), .A2(new_n353), .ZN(new_n481));
  NAND3_X1  g280(.A1(new_n481), .A2(new_n354), .A3(new_n363), .ZN(new_n482));
  INV_X1    g281(.A(KEYINPUT89), .ZN(new_n483));
  OAI21_X1  g282(.A(KEYINPUT37), .B1(new_n413), .B2(new_n414), .ZN(new_n484));
  INV_X1    g283(.A(KEYINPUT88), .ZN(new_n485));
  INV_X1    g284(.A(KEYINPUT37), .ZN(new_n486));
  NAND4_X1  g285(.A1(new_n417), .A2(new_n412), .A3(new_n485), .A4(new_n486), .ZN(new_n487));
  NAND3_X1  g286(.A1(new_n484), .A2(new_n487), .A3(new_n369), .ZN(new_n488));
  AOI21_X1  g287(.A(new_n485), .B1(new_n421), .B2(new_n486), .ZN(new_n489));
  OAI211_X1 g288(.A(new_n483), .B(KEYINPUT38), .C1(new_n488), .C2(new_n489), .ZN(new_n490));
  OAI21_X1  g289(.A(KEYINPUT38), .B1(new_n488), .B2(new_n489), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n491), .A2(KEYINPUT89), .ZN(new_n492));
  NAND3_X1  g291(.A1(new_n482), .A2(new_n490), .A3(new_n492), .ZN(new_n493));
  OR2_X1    g292(.A1(new_n488), .A2(new_n489), .ZN(new_n494));
  OAI211_X1 g293(.A(new_n356), .B(new_n419), .C1(new_n494), .C2(KEYINPUT38), .ZN(new_n495));
  OAI21_X1  g294(.A(new_n480), .B1(new_n493), .B2(new_n495), .ZN(new_n496));
  NOR2_X1   g295(.A1(new_n460), .A2(new_n461), .ZN(new_n497));
  NAND4_X1  g296(.A1(new_n365), .A2(new_n310), .A3(new_n424), .A4(new_n497), .ZN(new_n498));
  NAND2_X1  g297(.A1(new_n498), .A2(KEYINPUT35), .ZN(new_n499));
  INV_X1    g298(.A(new_n424), .ZN(new_n500));
  AOI21_X1  g299(.A(new_n500), .B1(new_n482), .B2(new_n356), .ZN(new_n501));
  NOR3_X1   g300(.A1(new_n309), .A2(new_n460), .A3(new_n461), .ZN(new_n502));
  INV_X1    g301(.A(KEYINPUT35), .ZN(new_n503));
  NAND3_X1  g302(.A1(new_n501), .A2(new_n502), .A3(new_n503), .ZN(new_n504));
  AOI22_X1  g303(.A1(new_n467), .A2(new_n496), .B1(new_n499), .B2(new_n504), .ZN(new_n505));
  INV_X1    g304(.A(KEYINPUT98), .ZN(new_n506));
  XNOR2_X1  g305(.A(G15gat), .B(G22gat), .ZN(new_n507));
  INV_X1    g306(.A(G1gat), .ZN(new_n508));
  NAND2_X1  g307(.A1(new_n508), .A2(KEYINPUT16), .ZN(new_n509));
  AND2_X1   g308(.A1(new_n507), .A2(new_n509), .ZN(new_n510));
  NOR2_X1   g309(.A1(new_n507), .A2(G1gat), .ZN(new_n511));
  OAI21_X1  g310(.A(G8gat), .B1(new_n510), .B2(new_n511), .ZN(new_n512));
  NAND2_X1  g311(.A1(new_n507), .A2(new_n509), .ZN(new_n513));
  INV_X1    g312(.A(G8gat), .ZN(new_n514));
  OAI211_X1 g313(.A(new_n513), .B(new_n514), .C1(G1gat), .C2(new_n507), .ZN(new_n515));
  AND2_X1   g314(.A1(new_n512), .A2(new_n515), .ZN(new_n516));
  XNOR2_X1  g315(.A(G43gat), .B(G50gat), .ZN(new_n517));
  NAND2_X1  g316(.A1(new_n517), .A2(KEYINPUT15), .ZN(new_n518));
  NAND2_X1  g317(.A1(G29gat), .A2(G36gat), .ZN(new_n519));
  INV_X1    g318(.A(KEYINPUT92), .ZN(new_n520));
  XNOR2_X1  g319(.A(new_n519), .B(new_n520), .ZN(new_n521));
  AND2_X1   g320(.A1(new_n518), .A2(new_n521), .ZN(new_n522));
  INV_X1    g321(.A(new_n517), .ZN(new_n523));
  INV_X1    g322(.A(KEYINPUT15), .ZN(new_n524));
  INV_X1    g323(.A(KEYINPUT14), .ZN(new_n525));
  INV_X1    g324(.A(G29gat), .ZN(new_n526));
  INV_X1    g325(.A(G36gat), .ZN(new_n527));
  NAND3_X1  g326(.A1(new_n525), .A2(new_n526), .A3(new_n527), .ZN(new_n528));
  OAI21_X1  g327(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n529));
  AOI22_X1  g328(.A1(new_n523), .A2(new_n524), .B1(new_n528), .B2(new_n529), .ZN(new_n530));
  NOR3_X1   g329(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n531));
  INV_X1    g330(.A(KEYINPUT91), .ZN(new_n532));
  OAI21_X1  g331(.A(new_n529), .B1(new_n531), .B2(new_n532), .ZN(new_n533));
  NOR2_X1   g332(.A1(new_n528), .A2(KEYINPUT91), .ZN(new_n534));
  OAI21_X1  g333(.A(new_n521), .B1(new_n533), .B2(new_n534), .ZN(new_n535));
  INV_X1    g334(.A(new_n518), .ZN(new_n536));
  AOI22_X1  g335(.A1(new_n522), .A2(new_n530), .B1(new_n535), .B2(new_n536), .ZN(new_n537));
  OAI21_X1  g336(.A(KEYINPUT94), .B1(new_n516), .B2(new_n537), .ZN(new_n538));
  NAND2_X1  g337(.A1(new_n522), .A2(new_n530), .ZN(new_n539));
  NAND2_X1  g338(.A1(new_n535), .A2(new_n536), .ZN(new_n540));
  NAND2_X1  g339(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  INV_X1    g340(.A(KEYINPUT94), .ZN(new_n542));
  NAND2_X1  g341(.A1(new_n512), .A2(new_n515), .ZN(new_n543));
  NAND3_X1  g342(.A1(new_n541), .A2(new_n542), .A3(new_n543), .ZN(new_n544));
  NAND2_X1  g343(.A1(new_n538), .A2(new_n544), .ZN(new_n545));
  INV_X1    g344(.A(KEYINPUT17), .ZN(new_n546));
  AND3_X1   g345(.A1(new_n539), .A2(new_n540), .A3(new_n546), .ZN(new_n547));
  AOI21_X1  g346(.A(new_n546), .B1(new_n539), .B2(new_n540), .ZN(new_n548));
  OAI21_X1  g347(.A(new_n516), .B1(new_n547), .B2(new_n548), .ZN(new_n549));
  NAND2_X1  g348(.A1(G229gat), .A2(G233gat), .ZN(new_n550));
  XOR2_X1   g349(.A(new_n550), .B(KEYINPUT93), .Z(new_n551));
  INV_X1    g350(.A(new_n551), .ZN(new_n552));
  NAND3_X1  g351(.A1(new_n545), .A2(new_n549), .A3(new_n552), .ZN(new_n553));
  INV_X1    g352(.A(KEYINPUT97), .ZN(new_n554));
  INV_X1    g353(.A(KEYINPUT18), .ZN(new_n555));
  AND3_X1   g354(.A1(new_n553), .A2(new_n554), .A3(new_n555), .ZN(new_n556));
  AOI21_X1  g355(.A(new_n554), .B1(new_n553), .B2(new_n555), .ZN(new_n557));
  NOR2_X1   g356(.A1(new_n556), .A2(new_n557), .ZN(new_n558));
  INV_X1    g357(.A(KEYINPUT95), .ZN(new_n559));
  OAI21_X1  g358(.A(new_n559), .B1(new_n541), .B2(new_n543), .ZN(new_n560));
  NAND3_X1  g359(.A1(new_n516), .A2(new_n537), .A3(KEYINPUT95), .ZN(new_n561));
  NAND3_X1  g360(.A1(new_n545), .A2(new_n560), .A3(new_n561), .ZN(new_n562));
  XNOR2_X1  g361(.A(new_n551), .B(KEYINPUT13), .ZN(new_n563));
  NAND2_X1  g362(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  NAND4_X1  g363(.A1(new_n545), .A2(new_n549), .A3(KEYINPUT18), .A4(new_n552), .ZN(new_n565));
  XNOR2_X1  g364(.A(G113gat), .B(G141gat), .ZN(new_n566));
  XNOR2_X1  g365(.A(KEYINPUT90), .B(KEYINPUT11), .ZN(new_n567));
  XNOR2_X1  g366(.A(new_n566), .B(new_n567), .ZN(new_n568));
  XNOR2_X1  g367(.A(G169gat), .B(G197gat), .ZN(new_n569));
  XNOR2_X1  g368(.A(new_n568), .B(new_n569), .ZN(new_n570));
  XOR2_X1   g369(.A(new_n570), .B(KEYINPUT12), .Z(new_n571));
  NAND3_X1  g370(.A1(new_n564), .A2(new_n565), .A3(new_n571), .ZN(new_n572));
  INV_X1    g371(.A(new_n572), .ZN(new_n573));
  AOI21_X1  g372(.A(new_n506), .B1(new_n558), .B2(new_n573), .ZN(new_n574));
  NOR4_X1   g373(.A1(new_n572), .A2(new_n556), .A3(new_n557), .A4(KEYINPUT98), .ZN(new_n575));
  NAND2_X1  g374(.A1(new_n553), .A2(new_n555), .ZN(new_n576));
  NAND3_X1  g375(.A1(new_n576), .A2(new_n564), .A3(new_n565), .ZN(new_n577));
  INV_X1    g376(.A(new_n571), .ZN(new_n578));
  NAND3_X1  g377(.A1(new_n577), .A2(KEYINPUT96), .A3(new_n578), .ZN(new_n579));
  INV_X1    g378(.A(new_n579), .ZN(new_n580));
  AOI21_X1  g379(.A(KEYINPUT96), .B1(new_n577), .B2(new_n578), .ZN(new_n581));
  OAI22_X1  g380(.A1(new_n574), .A2(new_n575), .B1(new_n580), .B2(new_n581), .ZN(new_n582));
  INV_X1    g381(.A(new_n582), .ZN(new_n583));
  AOI21_X1  g382(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n584));
  XNOR2_X1  g383(.A(new_n584), .B(KEYINPUT99), .ZN(new_n585));
  XNOR2_X1  g384(.A(G71gat), .B(G78gat), .ZN(new_n586));
  INV_X1    g385(.A(G64gat), .ZN(new_n587));
  NAND2_X1  g386(.A1(new_n587), .A2(G57gat), .ZN(new_n588));
  NAND2_X1  g387(.A1(new_n588), .A2(KEYINPUT100), .ZN(new_n589));
  INV_X1    g388(.A(KEYINPUT100), .ZN(new_n590));
  NAND3_X1  g389(.A1(new_n590), .A2(new_n587), .A3(G57gat), .ZN(new_n591));
  INV_X1    g390(.A(G57gat), .ZN(new_n592));
  NAND2_X1  g391(.A1(new_n592), .A2(G64gat), .ZN(new_n593));
  NAND3_X1  g392(.A1(new_n589), .A2(new_n591), .A3(new_n593), .ZN(new_n594));
  AND3_X1   g393(.A1(new_n585), .A2(new_n586), .A3(new_n594), .ZN(new_n595));
  NAND2_X1  g394(.A1(new_n593), .A2(new_n588), .ZN(new_n596));
  AOI21_X1  g395(.A(new_n586), .B1(new_n585), .B2(new_n596), .ZN(new_n597));
  OR2_X1    g396(.A1(new_n595), .A2(new_n597), .ZN(new_n598));
  INV_X1    g397(.A(KEYINPUT21), .ZN(new_n599));
  NAND2_X1  g398(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  NAND2_X1  g399(.A1(G231gat), .A2(G233gat), .ZN(new_n601));
  XNOR2_X1  g400(.A(new_n600), .B(new_n601), .ZN(new_n602));
  XOR2_X1   g401(.A(G127gat), .B(G155gat), .Z(new_n603));
  XNOR2_X1  g402(.A(new_n603), .B(KEYINPUT20), .ZN(new_n604));
  XNOR2_X1  g403(.A(new_n602), .B(new_n604), .ZN(new_n605));
  XNOR2_X1  g404(.A(G183gat), .B(G211gat), .ZN(new_n606));
  XNOR2_X1  g405(.A(new_n605), .B(new_n606), .ZN(new_n607));
  OAI21_X1  g406(.A(new_n516), .B1(new_n598), .B2(new_n599), .ZN(new_n608));
  XOR2_X1   g407(.A(KEYINPUT101), .B(KEYINPUT19), .Z(new_n609));
  XNOR2_X1  g408(.A(new_n608), .B(new_n609), .ZN(new_n610));
  INV_X1    g409(.A(new_n610), .ZN(new_n611));
  OR2_X1    g410(.A1(new_n607), .A2(new_n611), .ZN(new_n612));
  NAND2_X1  g411(.A1(new_n607), .A2(new_n611), .ZN(new_n613));
  NAND2_X1  g412(.A1(new_n612), .A2(new_n613), .ZN(new_n614));
  INV_X1    g413(.A(KEYINPUT102), .ZN(new_n615));
  NAND3_X1  g414(.A1(new_n615), .A2(G85gat), .A3(G92gat), .ZN(new_n616));
  INV_X1    g415(.A(KEYINPUT7), .ZN(new_n617));
  NAND2_X1  g416(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  NAND2_X1  g417(.A1(G99gat), .A2(G106gat), .ZN(new_n619));
  INV_X1    g418(.A(G85gat), .ZN(new_n620));
  INV_X1    g419(.A(G92gat), .ZN(new_n621));
  AOI22_X1  g420(.A1(KEYINPUT8), .A2(new_n619), .B1(new_n620), .B2(new_n621), .ZN(new_n622));
  NAND4_X1  g421(.A1(new_n615), .A2(KEYINPUT7), .A3(G85gat), .A4(G92gat), .ZN(new_n623));
  NAND3_X1  g422(.A1(new_n618), .A2(new_n622), .A3(new_n623), .ZN(new_n624));
  XNOR2_X1  g423(.A(G99gat), .B(G106gat), .ZN(new_n625));
  XNOR2_X1  g424(.A(new_n624), .B(new_n625), .ZN(new_n626));
  XNOR2_X1  g425(.A(new_n626), .B(KEYINPUT103), .ZN(new_n627));
  OAI21_X1  g426(.A(new_n627), .B1(new_n548), .B2(new_n547), .ZN(new_n628));
  XNOR2_X1  g427(.A(new_n628), .B(KEYINPUT104), .ZN(new_n629));
  INV_X1    g428(.A(new_n627), .ZN(new_n630));
  AND2_X1   g429(.A1(G232gat), .A2(G233gat), .ZN(new_n631));
  AOI22_X1  g430(.A1(new_n630), .A2(new_n541), .B1(KEYINPUT41), .B2(new_n631), .ZN(new_n632));
  NAND2_X1  g431(.A1(new_n629), .A2(new_n632), .ZN(new_n633));
  XOR2_X1   g432(.A(G190gat), .B(G218gat), .Z(new_n634));
  NAND2_X1  g433(.A1(new_n633), .A2(new_n634), .ZN(new_n635));
  NOR2_X1   g434(.A1(new_n631), .A2(KEYINPUT41), .ZN(new_n636));
  XNOR2_X1  g435(.A(G134gat), .B(G162gat), .ZN(new_n637));
  XNOR2_X1  g436(.A(new_n636), .B(new_n637), .ZN(new_n638));
  INV_X1    g437(.A(new_n634), .ZN(new_n639));
  NAND3_X1  g438(.A1(new_n629), .A2(new_n639), .A3(new_n632), .ZN(new_n640));
  AND3_X1   g439(.A1(new_n635), .A2(new_n638), .A3(new_n640), .ZN(new_n641));
  AOI21_X1  g440(.A(new_n638), .B1(new_n635), .B2(new_n640), .ZN(new_n642));
  NOR2_X1   g441(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  INV_X1    g442(.A(new_n643), .ZN(new_n644));
  NOR2_X1   g443(.A1(new_n595), .A2(new_n597), .ZN(new_n645));
  INV_X1    g444(.A(KEYINPUT105), .ZN(new_n646));
  OR2_X1    g445(.A1(new_n625), .A2(new_n646), .ZN(new_n647));
  XNOR2_X1  g446(.A(new_n647), .B(new_n624), .ZN(new_n648));
  NAND2_X1  g447(.A1(new_n645), .A2(new_n648), .ZN(new_n649));
  OAI211_X1 g448(.A(new_n649), .B(KEYINPUT106), .C1(new_n645), .C2(new_n626), .ZN(new_n650));
  INV_X1    g449(.A(KEYINPUT106), .ZN(new_n651));
  NAND3_X1  g450(.A1(new_n645), .A2(new_n648), .A3(new_n651), .ZN(new_n652));
  AOI21_X1  g451(.A(KEYINPUT10), .B1(new_n650), .B2(new_n652), .ZN(new_n653));
  INV_X1    g452(.A(KEYINPUT10), .ZN(new_n654));
  NOR3_X1   g453(.A1(new_n627), .A2(new_n654), .A3(new_n598), .ZN(new_n655));
  INV_X1    g454(.A(G230gat), .ZN(new_n656));
  OAI22_X1  g455(.A1(new_n653), .A2(new_n655), .B1(new_n656), .B2(new_n206), .ZN(new_n657));
  AND2_X1   g456(.A1(new_n650), .A2(new_n652), .ZN(new_n658));
  NOR2_X1   g457(.A1(new_n656), .A2(new_n206), .ZN(new_n659));
  NAND2_X1  g458(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  NAND2_X1  g459(.A1(new_n657), .A2(new_n660), .ZN(new_n661));
  XNOR2_X1  g460(.A(G120gat), .B(G148gat), .ZN(new_n662));
  XNOR2_X1  g461(.A(G176gat), .B(G204gat), .ZN(new_n663));
  XNOR2_X1  g462(.A(new_n662), .B(new_n663), .ZN(new_n664));
  OR2_X1    g463(.A1(new_n661), .A2(new_n664), .ZN(new_n665));
  NAND2_X1  g464(.A1(new_n661), .A2(new_n664), .ZN(new_n666));
  NAND2_X1  g465(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  INV_X1    g466(.A(new_n667), .ZN(new_n668));
  NAND3_X1  g467(.A1(new_n614), .A2(new_n644), .A3(new_n668), .ZN(new_n669));
  NOR3_X1   g468(.A1(new_n505), .A2(new_n583), .A3(new_n669), .ZN(new_n670));
  INV_X1    g469(.A(new_n365), .ZN(new_n671));
  NAND2_X1  g470(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  XNOR2_X1  g471(.A(new_n672), .B(G1gat), .ZN(G1324gat));
  NAND2_X1  g472(.A1(new_n670), .A2(new_n500), .ZN(new_n674));
  INV_X1    g473(.A(KEYINPUT42), .ZN(new_n675));
  XOR2_X1   g474(.A(KEYINPUT16), .B(G8gat), .Z(new_n676));
  INV_X1    g475(.A(new_n676), .ZN(new_n677));
  NOR4_X1   g476(.A1(new_n674), .A2(KEYINPUT107), .A3(new_n675), .A4(new_n677), .ZN(new_n678));
  INV_X1    g477(.A(KEYINPUT107), .ZN(new_n679));
  NOR2_X1   g478(.A1(new_n674), .A2(new_n677), .ZN(new_n680));
  AOI21_X1  g479(.A(new_n679), .B1(new_n680), .B2(KEYINPUT42), .ZN(new_n681));
  AOI21_X1  g480(.A(new_n514), .B1(new_n670), .B2(new_n500), .ZN(new_n682));
  OAI22_X1  g481(.A1(new_n682), .A2(new_n675), .B1(new_n674), .B2(new_n677), .ZN(new_n683));
  AOI21_X1  g482(.A(new_n678), .B1(new_n681), .B2(new_n683), .ZN(G1325gat));
  AND3_X1   g483(.A1(new_n670), .A2(G15gat), .A3(new_n466), .ZN(new_n685));
  AOI21_X1  g484(.A(G15gat), .B1(new_n670), .B2(new_n497), .ZN(new_n686));
  OR2_X1    g485(.A1(new_n686), .A2(KEYINPUT108), .ZN(new_n687));
  NAND2_X1  g486(.A1(new_n686), .A2(KEYINPUT108), .ZN(new_n688));
  AOI21_X1  g487(.A(new_n685), .B1(new_n687), .B2(new_n688), .ZN(G1326gat));
  NAND2_X1  g488(.A1(new_n670), .A2(new_n309), .ZN(new_n690));
  XNOR2_X1  g489(.A(new_n690), .B(KEYINPUT109), .ZN(new_n691));
  XNOR2_X1  g490(.A(KEYINPUT43), .B(G22gat), .ZN(new_n692));
  INV_X1    g491(.A(new_n692), .ZN(new_n693));
  NAND2_X1  g492(.A1(new_n691), .A2(new_n693), .ZN(new_n694));
  OR2_X1    g493(.A1(new_n690), .A2(KEYINPUT109), .ZN(new_n695));
  NAND2_X1  g494(.A1(new_n690), .A2(KEYINPUT109), .ZN(new_n696));
  NAND3_X1  g495(.A1(new_n695), .A2(new_n696), .A3(new_n692), .ZN(new_n697));
  NAND2_X1  g496(.A1(new_n694), .A2(new_n697), .ZN(G1327gat));
  INV_X1    g497(.A(KEYINPUT44), .ZN(new_n699));
  OAI21_X1  g498(.A(new_n699), .B1(new_n505), .B2(new_n644), .ZN(new_n700));
  INV_X1    g499(.A(new_n496), .ZN(new_n701));
  OAI211_X1 g500(.A(new_n464), .B(new_n465), .C1(new_n501), .C2(new_n310), .ZN(new_n702));
  AND3_X1   g501(.A1(new_n501), .A2(new_n502), .A3(new_n503), .ZN(new_n703));
  AOI21_X1  g502(.A(new_n503), .B1(new_n501), .B2(new_n502), .ZN(new_n704));
  OAI22_X1  g503(.A1(new_n701), .A2(new_n702), .B1(new_n703), .B2(new_n704), .ZN(new_n705));
  NAND3_X1  g504(.A1(new_n705), .A2(KEYINPUT44), .A3(new_n643), .ZN(new_n706));
  INV_X1    g505(.A(new_n614), .ZN(new_n707));
  NAND2_X1  g506(.A1(new_n707), .A2(new_n668), .ZN(new_n708));
  INV_X1    g507(.A(KEYINPUT110), .ZN(new_n709));
  NAND2_X1  g508(.A1(new_n582), .A2(new_n709), .ZN(new_n710));
  INV_X1    g509(.A(new_n710), .ZN(new_n711));
  OAI221_X1 g510(.A(KEYINPUT110), .B1(new_n580), .B2(new_n581), .C1(new_n574), .C2(new_n575), .ZN(new_n712));
  INV_X1    g511(.A(new_n712), .ZN(new_n713));
  NOR3_X1   g512(.A1(new_n708), .A2(new_n711), .A3(new_n713), .ZN(new_n714));
  NAND4_X1  g513(.A1(new_n700), .A2(new_n671), .A3(new_n706), .A4(new_n714), .ZN(new_n715));
  INV_X1    g514(.A(KEYINPUT111), .ZN(new_n716));
  AOI21_X1  g515(.A(new_n526), .B1(new_n715), .B2(new_n716), .ZN(new_n717));
  OAI21_X1  g516(.A(new_n717), .B1(new_n716), .B2(new_n715), .ZN(new_n718));
  NOR2_X1   g517(.A1(new_n505), .A2(new_n583), .ZN(new_n719));
  NOR2_X1   g518(.A1(new_n708), .A2(new_n644), .ZN(new_n720));
  NAND4_X1  g519(.A1(new_n719), .A2(new_n526), .A3(new_n671), .A4(new_n720), .ZN(new_n721));
  XNOR2_X1  g520(.A(new_n721), .B(KEYINPUT45), .ZN(new_n722));
  NAND2_X1  g521(.A1(new_n718), .A2(new_n722), .ZN(G1328gat));
  NAND4_X1  g522(.A1(new_n719), .A2(new_n527), .A3(new_n500), .A4(new_n720), .ZN(new_n724));
  INV_X1    g523(.A(KEYINPUT46), .ZN(new_n725));
  NOR2_X1   g524(.A1(new_n725), .A2(KEYINPUT112), .ZN(new_n726));
  AND2_X1   g525(.A1(new_n725), .A2(KEYINPUT112), .ZN(new_n727));
  OAI21_X1  g526(.A(new_n724), .B1(new_n726), .B2(new_n727), .ZN(new_n728));
  AND4_X1   g527(.A1(new_n500), .A2(new_n700), .A3(new_n706), .A4(new_n714), .ZN(new_n729));
  OAI221_X1 g528(.A(new_n728), .B1(new_n726), .B2(new_n724), .C1(new_n729), .C2(new_n527), .ZN(G1329gat));
  NAND4_X1  g529(.A1(new_n700), .A2(new_n466), .A3(new_n706), .A4(new_n714), .ZN(new_n731));
  NAND2_X1  g530(.A1(new_n731), .A2(G43gat), .ZN(new_n732));
  INV_X1    g531(.A(KEYINPUT47), .ZN(new_n733));
  INV_X1    g532(.A(G43gat), .ZN(new_n734));
  NAND4_X1  g533(.A1(new_n719), .A2(new_n734), .A3(new_n497), .A4(new_n720), .ZN(new_n735));
  AND3_X1   g534(.A1(new_n732), .A2(new_n733), .A3(new_n735), .ZN(new_n736));
  AOI21_X1  g535(.A(new_n733), .B1(new_n732), .B2(new_n735), .ZN(new_n737));
  NOR2_X1   g536(.A1(new_n736), .A2(new_n737), .ZN(G1330gat));
  NOR2_X1   g537(.A1(new_n310), .A2(G50gat), .ZN(new_n739));
  NAND4_X1  g538(.A1(new_n705), .A2(new_n582), .A3(new_n720), .A4(new_n739), .ZN(new_n740));
  NAND2_X1  g539(.A1(new_n740), .A2(KEYINPUT48), .ZN(new_n741));
  NAND4_X1  g540(.A1(new_n700), .A2(new_n309), .A3(new_n706), .A4(new_n714), .ZN(new_n742));
  AOI21_X1  g541(.A(new_n741), .B1(new_n742), .B2(G50gat), .ZN(new_n743));
  NOR2_X1   g542(.A1(new_n743), .A2(KEYINPUT114), .ZN(new_n744));
  INV_X1    g543(.A(KEYINPUT114), .ZN(new_n745));
  AOI211_X1 g544(.A(new_n745), .B(new_n741), .C1(new_n742), .C2(G50gat), .ZN(new_n746));
  INV_X1    g545(.A(new_n740), .ZN(new_n747));
  AOI21_X1  g546(.A(new_n747), .B1(new_n742), .B2(G50gat), .ZN(new_n748));
  XOR2_X1   g547(.A(KEYINPUT113), .B(KEYINPUT48), .Z(new_n749));
  OAI22_X1  g548(.A1(new_n744), .A2(new_n746), .B1(new_n748), .B2(new_n749), .ZN(G1331gat));
  NOR2_X1   g549(.A1(new_n711), .A2(new_n713), .ZN(new_n751));
  NOR4_X1   g550(.A1(new_n751), .A2(new_n707), .A3(new_n643), .A4(new_n668), .ZN(new_n752));
  NAND2_X1  g551(.A1(new_n705), .A2(new_n752), .ZN(new_n753));
  NOR2_X1   g552(.A1(new_n753), .A2(new_n365), .ZN(new_n754));
  XNOR2_X1  g553(.A(new_n754), .B(new_n592), .ZN(G1332gat));
  NOR2_X1   g554(.A1(new_n753), .A2(new_n424), .ZN(new_n756));
  NOR2_X1   g555(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n757));
  AND2_X1   g556(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n758));
  OAI21_X1  g557(.A(new_n756), .B1(new_n757), .B2(new_n758), .ZN(new_n759));
  OAI21_X1  g558(.A(new_n759), .B1(new_n756), .B2(new_n757), .ZN(G1333gat));
  AND2_X1   g559(.A1(new_n464), .A2(new_n465), .ZN(new_n761));
  OAI21_X1  g560(.A(G71gat), .B1(new_n753), .B2(new_n761), .ZN(new_n762));
  INV_X1    g561(.A(G71gat), .ZN(new_n763));
  NAND2_X1  g562(.A1(new_n497), .A2(new_n763), .ZN(new_n764));
  OAI21_X1  g563(.A(new_n762), .B1(new_n753), .B2(new_n764), .ZN(new_n765));
  XOR2_X1   g564(.A(new_n765), .B(KEYINPUT50), .Z(G1334gat));
  NOR2_X1   g565(.A1(new_n753), .A2(new_n310), .ZN(new_n767));
  XOR2_X1   g566(.A(new_n767), .B(G78gat), .Z(G1335gat));
  NOR3_X1   g567(.A1(new_n751), .A2(new_n614), .A3(new_n668), .ZN(new_n769));
  NAND3_X1  g568(.A1(new_n700), .A2(new_n706), .A3(new_n769), .ZN(new_n770));
  OAI21_X1  g569(.A(G85gat), .B1(new_n770), .B2(new_n365), .ZN(new_n771));
  NOR3_X1   g570(.A1(new_n365), .A2(G85gat), .A3(new_n668), .ZN(new_n772));
  NOR2_X1   g571(.A1(new_n751), .A2(new_n614), .ZN(new_n773));
  AND4_X1   g572(.A1(KEYINPUT51), .A2(new_n705), .A3(new_n643), .A4(new_n773), .ZN(new_n774));
  INV_X1    g573(.A(new_n425), .ZN(new_n775));
  NAND3_X1  g574(.A1(new_n775), .A2(new_n761), .A3(new_n496), .ZN(new_n776));
  NAND2_X1  g575(.A1(new_n499), .A2(new_n504), .ZN(new_n777));
  AOI21_X1  g576(.A(new_n644), .B1(new_n776), .B2(new_n777), .ZN(new_n778));
  AOI21_X1  g577(.A(KEYINPUT51), .B1(new_n778), .B2(new_n773), .ZN(new_n779));
  OAI21_X1  g578(.A(new_n772), .B1(new_n774), .B2(new_n779), .ZN(new_n780));
  NAND2_X1  g579(.A1(new_n771), .A2(new_n780), .ZN(new_n781));
  INV_X1    g580(.A(KEYINPUT115), .ZN(new_n782));
  NAND2_X1  g581(.A1(new_n781), .A2(new_n782), .ZN(new_n783));
  NAND3_X1  g582(.A1(new_n771), .A2(new_n780), .A3(KEYINPUT115), .ZN(new_n784));
  NAND2_X1  g583(.A1(new_n783), .A2(new_n784), .ZN(G1336gat));
  NAND4_X1  g584(.A1(new_n700), .A2(new_n500), .A3(new_n706), .A4(new_n769), .ZN(new_n786));
  NAND2_X1  g585(.A1(new_n786), .A2(G92gat), .ZN(new_n787));
  NAND2_X1  g586(.A1(new_n787), .A2(KEYINPUT116), .ZN(new_n788));
  NOR3_X1   g587(.A1(new_n668), .A2(G92gat), .A3(new_n424), .ZN(new_n789));
  OAI21_X1  g588(.A(new_n789), .B1(new_n774), .B2(new_n779), .ZN(new_n790));
  NAND2_X1  g589(.A1(new_n787), .A2(new_n790), .ZN(new_n791));
  NAND3_X1  g590(.A1(new_n788), .A2(new_n791), .A3(KEYINPUT52), .ZN(new_n792));
  INV_X1    g591(.A(KEYINPUT52), .ZN(new_n793));
  OAI211_X1 g592(.A(new_n787), .B(new_n790), .C1(KEYINPUT116), .C2(new_n793), .ZN(new_n794));
  NAND2_X1  g593(.A1(new_n792), .A2(new_n794), .ZN(G1337gat));
  OAI21_X1  g594(.A(G99gat), .B1(new_n770), .B2(new_n761), .ZN(new_n796));
  NOR2_X1   g595(.A1(new_n668), .A2(G99gat), .ZN(new_n797));
  OAI211_X1 g596(.A(new_n497), .B(new_n797), .C1(new_n774), .C2(new_n779), .ZN(new_n798));
  NAND2_X1  g597(.A1(new_n796), .A2(new_n798), .ZN(new_n799));
  INV_X1    g598(.A(KEYINPUT117), .ZN(new_n800));
  NAND2_X1  g599(.A1(new_n799), .A2(new_n800), .ZN(new_n801));
  NAND3_X1  g600(.A1(new_n796), .A2(new_n798), .A3(KEYINPUT117), .ZN(new_n802));
  NAND2_X1  g601(.A1(new_n801), .A2(new_n802), .ZN(G1338gat));
  NAND4_X1  g602(.A1(new_n700), .A2(new_n309), .A3(new_n706), .A4(new_n769), .ZN(new_n804));
  NAND2_X1  g603(.A1(new_n804), .A2(G106gat), .ZN(new_n805));
  NAND2_X1  g604(.A1(new_n805), .A2(KEYINPUT118), .ZN(new_n806));
  NOR3_X1   g605(.A1(new_n310), .A2(G106gat), .A3(new_n668), .ZN(new_n807));
  OAI21_X1  g606(.A(new_n807), .B1(new_n774), .B2(new_n779), .ZN(new_n808));
  NAND2_X1  g607(.A1(new_n805), .A2(new_n808), .ZN(new_n809));
  NAND3_X1  g608(.A1(new_n806), .A2(new_n809), .A3(KEYINPUT53), .ZN(new_n810));
  INV_X1    g609(.A(KEYINPUT53), .ZN(new_n811));
  OAI211_X1 g610(.A(new_n805), .B(new_n808), .C1(KEYINPUT118), .C2(new_n811), .ZN(new_n812));
  NAND2_X1  g611(.A1(new_n810), .A2(new_n812), .ZN(G1339gat));
  NAND3_X1  g612(.A1(new_n630), .A2(KEYINPUT10), .A3(new_n645), .ZN(new_n814));
  OAI211_X1 g613(.A(new_n659), .B(new_n814), .C1(new_n658), .C2(KEYINPUT10), .ZN(new_n815));
  NAND3_X1  g614(.A1(new_n815), .A2(new_n657), .A3(KEYINPUT54), .ZN(new_n816));
  INV_X1    g615(.A(KEYINPUT54), .ZN(new_n817));
  OAI221_X1 g616(.A(new_n817), .B1(new_n656), .B2(new_n206), .C1(new_n653), .C2(new_n655), .ZN(new_n818));
  NAND4_X1  g617(.A1(new_n816), .A2(KEYINPUT55), .A3(new_n664), .A4(new_n818), .ZN(new_n819));
  NAND2_X1  g618(.A1(new_n819), .A2(new_n665), .ZN(new_n820));
  AND2_X1   g619(.A1(new_n818), .A2(new_n664), .ZN(new_n821));
  AOI21_X1  g620(.A(KEYINPUT55), .B1(new_n821), .B2(new_n816), .ZN(new_n822));
  NOR2_X1   g621(.A1(new_n820), .A2(new_n822), .ZN(new_n823));
  NAND3_X1  g622(.A1(new_n710), .A2(new_n712), .A3(new_n823), .ZN(new_n824));
  OR2_X1    g623(.A1(new_n574), .A2(new_n575), .ZN(new_n825));
  INV_X1    g624(.A(new_n570), .ZN(new_n826));
  NOR2_X1   g625(.A1(new_n562), .A2(new_n563), .ZN(new_n827));
  AOI21_X1  g626(.A(new_n552), .B1(new_n545), .B2(new_n549), .ZN(new_n828));
  OAI21_X1  g627(.A(new_n826), .B1(new_n827), .B2(new_n828), .ZN(new_n829));
  NAND3_X1  g628(.A1(new_n825), .A2(new_n667), .A3(new_n829), .ZN(new_n830));
  AOI21_X1  g629(.A(new_n643), .B1(new_n824), .B2(new_n830), .ZN(new_n831));
  AND4_X1   g630(.A1(new_n825), .A2(new_n643), .A3(new_n823), .A4(new_n829), .ZN(new_n832));
  OAI21_X1  g631(.A(new_n707), .B1(new_n831), .B2(new_n832), .ZN(new_n833));
  OR2_X1    g632(.A1(new_n751), .A2(new_n669), .ZN(new_n834));
  AOI21_X1  g633(.A(new_n365), .B1(new_n833), .B2(new_n834), .ZN(new_n835));
  AND2_X1   g634(.A1(new_n835), .A2(new_n502), .ZN(new_n836));
  AND2_X1   g635(.A1(new_n836), .A2(new_n424), .ZN(new_n837));
  AOI21_X1  g636(.A(G113gat), .B1(new_n837), .B2(new_n751), .ZN(new_n838));
  AOI21_X1  g637(.A(new_n309), .B1(new_n833), .B2(new_n834), .ZN(new_n839));
  NAND4_X1  g638(.A1(new_n839), .A2(new_n671), .A3(new_n424), .A4(new_n497), .ZN(new_n840));
  XNOR2_X1  g639(.A(new_n840), .B(KEYINPUT119), .ZN(new_n841));
  NOR2_X1   g640(.A1(new_n583), .A2(new_n311), .ZN(new_n842));
  AOI21_X1  g641(.A(new_n838), .B1(new_n841), .B2(new_n842), .ZN(G1340gat));
  XOR2_X1   g642(.A(new_n840), .B(KEYINPUT119), .Z(new_n844));
  OAI21_X1  g643(.A(G120gat), .B1(new_n844), .B2(new_n668), .ZN(new_n845));
  NAND3_X1  g644(.A1(new_n837), .A2(new_n315), .A3(new_n667), .ZN(new_n846));
  NAND2_X1  g645(.A1(new_n845), .A2(new_n846), .ZN(G1341gat));
  AND3_X1   g646(.A1(new_n836), .A2(new_n424), .A3(new_n614), .ZN(new_n848));
  OR2_X1    g647(.A1(new_n848), .A2(KEYINPUT120), .ZN(new_n849));
  AOI21_X1  g648(.A(G127gat), .B1(new_n848), .B2(KEYINPUT120), .ZN(new_n850));
  AND2_X1   g649(.A1(new_n614), .A2(G127gat), .ZN(new_n851));
  AOI22_X1  g650(.A1(new_n849), .A2(new_n850), .B1(new_n841), .B2(new_n851), .ZN(G1342gat));
  OAI21_X1  g651(.A(G134gat), .B1(new_n844), .B2(new_n644), .ZN(new_n853));
  NOR3_X1   g652(.A1(new_n644), .A2(G134gat), .A3(new_n500), .ZN(new_n854));
  NAND2_X1  g653(.A1(new_n836), .A2(new_n854), .ZN(new_n855));
  XOR2_X1   g654(.A(new_n855), .B(KEYINPUT56), .Z(new_n856));
  NAND2_X1  g655(.A1(new_n853), .A2(new_n856), .ZN(G1343gat));
  NOR3_X1   g656(.A1(new_n466), .A2(new_n365), .A3(new_n500), .ZN(new_n858));
  NAND2_X1  g657(.A1(new_n833), .A2(new_n834), .ZN(new_n859));
  AOI21_X1  g658(.A(KEYINPUT57), .B1(new_n859), .B2(new_n309), .ZN(new_n860));
  NAND2_X1  g659(.A1(new_n309), .A2(KEYINPUT57), .ZN(new_n861));
  NAND2_X1  g660(.A1(new_n823), .A2(new_n582), .ZN(new_n862));
  AOI21_X1  g661(.A(new_n643), .B1(new_n862), .B2(new_n830), .ZN(new_n863));
  OAI21_X1  g662(.A(new_n707), .B1(new_n863), .B2(new_n832), .ZN(new_n864));
  AOI21_X1  g663(.A(new_n861), .B1(new_n834), .B2(new_n864), .ZN(new_n865));
  OAI211_X1 g664(.A(new_n751), .B(new_n858), .C1(new_n860), .C2(new_n865), .ZN(new_n866));
  NAND2_X1  g665(.A1(new_n866), .A2(G141gat), .ZN(new_n867));
  NOR3_X1   g666(.A1(new_n466), .A2(new_n310), .A3(new_n500), .ZN(new_n868));
  NOR2_X1   g667(.A1(new_n583), .A2(G141gat), .ZN(new_n869));
  NAND3_X1  g668(.A1(new_n835), .A2(new_n868), .A3(new_n869), .ZN(new_n870));
  NAND2_X1  g669(.A1(new_n867), .A2(new_n870), .ZN(new_n871));
  NAND2_X1  g670(.A1(new_n871), .A2(KEYINPUT58), .ZN(new_n872));
  XNOR2_X1  g671(.A(KEYINPUT122), .B(KEYINPUT58), .ZN(new_n873));
  NAND2_X1  g672(.A1(new_n870), .A2(KEYINPUT121), .ZN(new_n874));
  INV_X1    g673(.A(KEYINPUT121), .ZN(new_n875));
  NAND4_X1  g674(.A1(new_n835), .A2(new_n875), .A3(new_n868), .A4(new_n869), .ZN(new_n876));
  AOI21_X1  g675(.A(new_n873), .B1(new_n874), .B2(new_n876), .ZN(new_n877));
  OAI211_X1 g676(.A(new_n582), .B(new_n858), .C1(new_n860), .C2(new_n865), .ZN(new_n878));
  NAND2_X1  g677(.A1(new_n878), .A2(G141gat), .ZN(new_n879));
  AND3_X1   g678(.A1(new_n877), .A2(new_n879), .A3(KEYINPUT123), .ZN(new_n880));
  AOI21_X1  g679(.A(KEYINPUT123), .B1(new_n877), .B2(new_n879), .ZN(new_n881));
  OAI21_X1  g680(.A(new_n872), .B1(new_n880), .B2(new_n881), .ZN(G1344gat));
  OAI21_X1  g681(.A(new_n864), .B1(new_n582), .B2(new_n669), .ZN(new_n883));
  AOI21_X1  g682(.A(KEYINPUT57), .B1(new_n883), .B2(new_n309), .ZN(new_n884));
  AOI21_X1  g683(.A(new_n861), .B1(new_n833), .B2(new_n834), .ZN(new_n885));
  OR2_X1    g684(.A1(new_n884), .A2(new_n885), .ZN(new_n886));
  NAND3_X1  g685(.A1(new_n886), .A2(new_n667), .A3(new_n858), .ZN(new_n887));
  NAND3_X1  g686(.A1(new_n887), .A2(KEYINPUT59), .A3(G148gat), .ZN(new_n888));
  OAI21_X1  g687(.A(new_n858), .B1(new_n860), .B2(new_n865), .ZN(new_n889));
  OR3_X1    g688(.A1(new_n889), .A2(KEYINPUT59), .A3(new_n668), .ZN(new_n890));
  NAND2_X1  g689(.A1(new_n835), .A2(new_n868), .ZN(new_n891));
  OAI21_X1  g690(.A(KEYINPUT59), .B1(new_n891), .B2(new_n668), .ZN(new_n892));
  NAND2_X1  g691(.A1(new_n892), .A2(new_n221), .ZN(new_n893));
  NAND3_X1  g692(.A1(new_n888), .A2(new_n890), .A3(new_n893), .ZN(G1345gat));
  OAI21_X1  g693(.A(new_n235), .B1(new_n889), .B2(new_n707), .ZN(new_n895));
  INV_X1    g694(.A(new_n891), .ZN(new_n896));
  NAND3_X1  g695(.A1(new_n896), .A2(new_n254), .A3(new_n614), .ZN(new_n897));
  NAND2_X1  g696(.A1(new_n895), .A2(new_n897), .ZN(G1346gat));
  OAI21_X1  g697(.A(new_n239), .B1(new_n889), .B2(new_n644), .ZN(new_n899));
  NAND3_X1  g698(.A1(new_n896), .A2(new_n255), .A3(new_n643), .ZN(new_n900));
  NAND2_X1  g699(.A1(new_n899), .A2(new_n900), .ZN(G1347gat));
  AND3_X1   g700(.A1(new_n365), .A2(new_n500), .A3(new_n497), .ZN(new_n902));
  NAND2_X1  g701(.A1(new_n839), .A2(new_n902), .ZN(new_n903));
  INV_X1    g702(.A(G169gat), .ZN(new_n904));
  NOR3_X1   g703(.A1(new_n903), .A2(new_n904), .A3(new_n583), .ZN(new_n905));
  AOI21_X1  g704(.A(new_n671), .B1(new_n833), .B2(new_n834), .ZN(new_n906));
  AND2_X1   g705(.A1(new_n502), .A2(new_n500), .ZN(new_n907));
  NAND2_X1  g706(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  INV_X1    g707(.A(new_n908), .ZN(new_n909));
  NAND2_X1  g708(.A1(new_n909), .A2(new_n751), .ZN(new_n910));
  AOI21_X1  g709(.A(new_n905), .B1(new_n904), .B2(new_n910), .ZN(G1348gat));
  OR3_X1    g710(.A1(new_n908), .A2(G176gat), .A3(new_n668), .ZN(new_n912));
  OAI21_X1  g711(.A(G176gat), .B1(new_n903), .B2(new_n668), .ZN(new_n913));
  NAND2_X1  g712(.A1(new_n912), .A2(new_n913), .ZN(G1349gat));
  NAND3_X1  g713(.A1(new_n909), .A2(new_n396), .A3(new_n614), .ZN(new_n915));
  OAI21_X1  g714(.A(G183gat), .B1(new_n903), .B2(new_n707), .ZN(new_n916));
  NAND3_X1  g715(.A1(new_n915), .A2(KEYINPUT124), .A3(new_n916), .ZN(new_n917));
  XNOR2_X1  g716(.A(new_n917), .B(KEYINPUT60), .ZN(G1350gat));
  NAND3_X1  g717(.A1(new_n909), .A2(new_n397), .A3(new_n643), .ZN(new_n919));
  XNOR2_X1  g718(.A(new_n919), .B(KEYINPUT125), .ZN(new_n920));
  NAND3_X1  g719(.A1(new_n839), .A2(new_n643), .A3(new_n902), .ZN(new_n921));
  AND2_X1   g720(.A1(new_n921), .A2(G190gat), .ZN(new_n922));
  OR2_X1    g721(.A1(new_n922), .A2(KEYINPUT61), .ZN(new_n923));
  NAND2_X1  g722(.A1(new_n922), .A2(KEYINPUT61), .ZN(new_n924));
  NAND3_X1  g723(.A1(new_n920), .A2(new_n923), .A3(new_n924), .ZN(G1351gat));
  AND4_X1   g724(.A1(new_n309), .A2(new_n906), .A3(new_n500), .A4(new_n761), .ZN(new_n926));
  AOI21_X1  g725(.A(G197gat), .B1(new_n926), .B2(new_n751), .ZN(new_n927));
  NOR3_X1   g726(.A1(new_n466), .A2(new_n671), .A3(new_n424), .ZN(new_n928));
  NAND2_X1  g727(.A1(new_n886), .A2(new_n928), .ZN(new_n929));
  INV_X1    g728(.A(new_n929), .ZN(new_n930));
  AND2_X1   g729(.A1(new_n582), .A2(G197gat), .ZN(new_n931));
  AOI21_X1  g730(.A(new_n927), .B1(new_n930), .B2(new_n931), .ZN(G1352gat));
  XNOR2_X1  g731(.A(KEYINPUT126), .B(G204gat), .ZN(new_n933));
  OAI21_X1  g732(.A(new_n933), .B1(new_n929), .B2(new_n668), .ZN(new_n934));
  NOR2_X1   g733(.A1(new_n668), .A2(new_n933), .ZN(new_n935));
  NAND2_X1  g734(.A1(new_n926), .A2(new_n935), .ZN(new_n936));
  OR2_X1    g735(.A1(new_n936), .A2(KEYINPUT62), .ZN(new_n937));
  NAND2_X1  g736(.A1(new_n936), .A2(KEYINPUT62), .ZN(new_n938));
  NAND3_X1  g737(.A1(new_n934), .A2(new_n937), .A3(new_n938), .ZN(G1353gat));
  NAND3_X1  g738(.A1(new_n926), .A2(new_n210), .A3(new_n614), .ZN(new_n940));
  OAI211_X1 g739(.A(new_n614), .B(new_n928), .C1(new_n884), .C2(new_n885), .ZN(new_n941));
  AND3_X1   g740(.A1(new_n941), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n942));
  AOI21_X1  g741(.A(KEYINPUT63), .B1(new_n941), .B2(G211gat), .ZN(new_n943));
  OAI21_X1  g742(.A(new_n940), .B1(new_n942), .B2(new_n943), .ZN(G1354gat));
  OAI21_X1  g743(.A(G218gat), .B1(new_n929), .B2(new_n644), .ZN(new_n945));
  NAND3_X1  g744(.A1(new_n926), .A2(new_n211), .A3(new_n643), .ZN(new_n946));
  NAND2_X1  g745(.A1(new_n945), .A2(new_n946), .ZN(G1355gat));
endmodule


