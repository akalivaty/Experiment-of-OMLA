//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 0 0 1 0 1 0 1 0 1 1 1 0 0 1 1 1 1 1 1 1 1 1 1 0 0 0 1 1 1 0 1 0 0 1 0 1 1 0 1 0 1 1 0 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 1 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:20:20 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n622,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n633, new_n634, new_n635, new_n636, new_n637,
    new_n638, new_n639, new_n640, new_n641, new_n642, new_n644, new_n645,
    new_n646, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n701, new_n702, new_n703,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n730, new_n731, new_n732, new_n734, new_n735, new_n736,
    new_n738, new_n740, new_n741, new_n742, new_n743, new_n744, new_n745,
    new_n746, new_n747, new_n748, new_n749, new_n750, new_n751, new_n752,
    new_n753, new_n754, new_n755, new_n756, new_n757, new_n758, new_n759,
    new_n760, new_n761, new_n762, new_n763, new_n764, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n776, new_n777, new_n778, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n837, new_n838, new_n839, new_n841, new_n842,
    new_n843, new_n845, new_n846, new_n847, new_n848, new_n849, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n918, new_n919, new_n921, new_n922, new_n923, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n939, new_n940, new_n941,
    new_n942, new_n943, new_n944, new_n945, new_n947, new_n948, new_n949,
    new_n950, new_n951, new_n952, new_n953, new_n955, new_n956, new_n957,
    new_n958, new_n959, new_n960, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n968, new_n969, new_n970, new_n971, new_n972, new_n974,
    new_n975;
  NAND3_X1  g000(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n202));
  NAND2_X1  g001(.A1(new_n202), .A2(KEYINPUT64), .ZN(new_n203));
  INV_X1    g002(.A(KEYINPUT64), .ZN(new_n204));
  NAND4_X1  g003(.A1(new_n204), .A2(KEYINPUT24), .A3(G183gat), .A4(G190gat), .ZN(new_n205));
  NAND2_X1  g004(.A1(G183gat), .A2(G190gat), .ZN(new_n206));
  INV_X1    g005(.A(KEYINPUT24), .ZN(new_n207));
  NAND2_X1  g006(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  INV_X1    g007(.A(G183gat), .ZN(new_n209));
  INV_X1    g008(.A(G190gat), .ZN(new_n210));
  NAND2_X1  g009(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  NAND4_X1  g010(.A1(new_n203), .A2(new_n205), .A3(new_n208), .A4(new_n211), .ZN(new_n212));
  NAND2_X1  g011(.A1(G169gat), .A2(G176gat), .ZN(new_n213));
  INV_X1    g012(.A(new_n213), .ZN(new_n214));
  NOR2_X1   g013(.A1(G169gat), .A2(G176gat), .ZN(new_n215));
  AOI21_X1  g014(.A(new_n214), .B1(KEYINPUT23), .B2(new_n215), .ZN(new_n216));
  INV_X1    g015(.A(KEYINPUT23), .ZN(new_n217));
  OAI21_X1  g016(.A(new_n217), .B1(G169gat), .B2(G176gat), .ZN(new_n218));
  NAND4_X1  g017(.A1(new_n212), .A2(KEYINPUT25), .A3(new_n216), .A4(new_n218), .ZN(new_n219));
  INV_X1    g018(.A(KEYINPUT25), .ZN(new_n220));
  AND3_X1   g019(.A1(new_n208), .A2(new_n202), .A3(new_n211), .ZN(new_n221));
  NAND2_X1  g020(.A1(new_n215), .A2(KEYINPUT23), .ZN(new_n222));
  NAND3_X1  g021(.A1(new_n222), .A2(new_n218), .A3(new_n213), .ZN(new_n223));
  OAI21_X1  g022(.A(new_n220), .B1(new_n221), .B2(new_n223), .ZN(new_n224));
  NAND2_X1  g023(.A1(new_n219), .A2(new_n224), .ZN(new_n225));
  INV_X1    g024(.A(KEYINPUT28), .ZN(new_n226));
  NOR2_X1   g025(.A1(new_n226), .A2(G190gat), .ZN(new_n227));
  NAND2_X1  g026(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n228));
  INV_X1    g027(.A(new_n228), .ZN(new_n229));
  NOR2_X1   g028(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n230));
  INV_X1    g029(.A(KEYINPUT66), .ZN(new_n231));
  NOR3_X1   g030(.A1(new_n229), .A2(new_n230), .A3(new_n231), .ZN(new_n232));
  INV_X1    g031(.A(KEYINPUT27), .ZN(new_n233));
  NAND2_X1  g032(.A1(new_n233), .A2(new_n209), .ZN(new_n234));
  AOI21_X1  g033(.A(KEYINPUT66), .B1(new_n234), .B2(new_n228), .ZN(new_n235));
  OAI21_X1  g034(.A(new_n227), .B1(new_n232), .B2(new_n235), .ZN(new_n236));
  INV_X1    g035(.A(KEYINPUT65), .ZN(new_n237));
  AOI21_X1  g036(.A(G190gat), .B1(new_n234), .B2(new_n228), .ZN(new_n238));
  OAI21_X1  g037(.A(new_n237), .B1(new_n238), .B2(KEYINPUT28), .ZN(new_n239));
  OAI21_X1  g038(.A(new_n210), .B1(new_n229), .B2(new_n230), .ZN(new_n240));
  NAND3_X1  g039(.A1(new_n240), .A2(KEYINPUT65), .A3(new_n226), .ZN(new_n241));
  NAND3_X1  g040(.A1(new_n236), .A2(new_n239), .A3(new_n241), .ZN(new_n242));
  INV_X1    g041(.A(new_n215), .ZN(new_n243));
  OR2_X1    g042(.A1(new_n243), .A2(KEYINPUT26), .ZN(new_n244));
  AOI21_X1  g043(.A(new_n214), .B1(new_n243), .B2(KEYINPUT26), .ZN(new_n245));
  AOI22_X1  g044(.A1(new_n244), .A2(new_n245), .B1(G183gat), .B2(G190gat), .ZN(new_n246));
  AND3_X1   g045(.A1(new_n242), .A2(KEYINPUT67), .A3(new_n246), .ZN(new_n247));
  AOI21_X1  g046(.A(KEYINPUT67), .B1(new_n242), .B2(new_n246), .ZN(new_n248));
  OAI21_X1  g047(.A(new_n225), .B1(new_n247), .B2(new_n248), .ZN(new_n249));
  XOR2_X1   g048(.A(G127gat), .B(G134gat), .Z(new_n250));
  XNOR2_X1  g049(.A(G113gat), .B(G120gat), .ZN(new_n251));
  OAI21_X1  g050(.A(new_n250), .B1(KEYINPUT1), .B2(new_n251), .ZN(new_n252));
  XOR2_X1   g051(.A(G113gat), .B(G120gat), .Z(new_n253));
  INV_X1    g052(.A(KEYINPUT1), .ZN(new_n254));
  XNOR2_X1  g053(.A(G127gat), .B(G134gat), .ZN(new_n255));
  NAND3_X1  g054(.A1(new_n253), .A2(new_n254), .A3(new_n255), .ZN(new_n256));
  NAND2_X1  g055(.A1(new_n252), .A2(new_n256), .ZN(new_n257));
  NAND2_X1  g056(.A1(new_n249), .A2(new_n257), .ZN(new_n258));
  NAND2_X1  g057(.A1(G227gat), .A2(G233gat), .ZN(new_n259));
  AND2_X1   g058(.A1(new_n252), .A2(new_n256), .ZN(new_n260));
  OAI211_X1 g059(.A(new_n260), .B(new_n225), .C1(new_n247), .C2(new_n248), .ZN(new_n261));
  NAND3_X1  g060(.A1(new_n258), .A2(new_n259), .A3(new_n261), .ZN(new_n262));
  INV_X1    g061(.A(KEYINPUT71), .ZN(new_n263));
  AND3_X1   g062(.A1(new_n262), .A2(new_n263), .A3(KEYINPUT34), .ZN(new_n264));
  AOI21_X1  g063(.A(KEYINPUT34), .B1(new_n262), .B2(new_n263), .ZN(new_n265));
  NOR2_X1   g064(.A1(new_n264), .A2(new_n265), .ZN(new_n266));
  INV_X1    g065(.A(KEYINPUT69), .ZN(new_n267));
  XOR2_X1   g066(.A(G71gat), .B(G99gat), .Z(new_n268));
  XNOR2_X1  g067(.A(new_n268), .B(KEYINPUT70), .ZN(new_n269));
  XNOR2_X1  g068(.A(G15gat), .B(G43gat), .ZN(new_n270));
  XNOR2_X1  g069(.A(new_n269), .B(new_n270), .ZN(new_n271));
  AOI21_X1  g070(.A(new_n259), .B1(new_n258), .B2(new_n261), .ZN(new_n272));
  XNOR2_X1  g071(.A(KEYINPUT68), .B(KEYINPUT33), .ZN(new_n273));
  OAI211_X1 g072(.A(new_n267), .B(new_n271), .C1(new_n272), .C2(new_n273), .ZN(new_n274));
  AND2_X1   g073(.A1(new_n258), .A2(new_n261), .ZN(new_n275));
  OAI21_X1  g074(.A(KEYINPUT32), .B1(new_n275), .B2(new_n259), .ZN(new_n276));
  NAND2_X1  g075(.A1(new_n274), .A2(new_n276), .ZN(new_n277));
  OAI211_X1 g076(.A(KEYINPUT69), .B(new_n271), .C1(new_n272), .C2(new_n273), .ZN(new_n278));
  INV_X1    g077(.A(KEYINPUT32), .ZN(new_n279));
  NAND2_X1  g078(.A1(new_n271), .A2(new_n273), .ZN(new_n280));
  NOR3_X1   g079(.A1(new_n272), .A2(new_n279), .A3(new_n280), .ZN(new_n281));
  NAND2_X1  g080(.A1(new_n278), .A2(new_n281), .ZN(new_n282));
  AOI21_X1  g081(.A(new_n266), .B1(new_n277), .B2(new_n282), .ZN(new_n283));
  INV_X1    g082(.A(new_n283), .ZN(new_n284));
  NAND3_X1  g083(.A1(new_n266), .A2(new_n282), .A3(new_n277), .ZN(new_n285));
  NAND3_X1  g084(.A1(new_n284), .A2(KEYINPUT82), .A3(new_n285), .ZN(new_n286));
  XNOR2_X1  g085(.A(G197gat), .B(G204gat), .ZN(new_n287));
  INV_X1    g086(.A(G211gat), .ZN(new_n288));
  INV_X1    g087(.A(G218gat), .ZN(new_n289));
  NOR2_X1   g088(.A1(new_n288), .A2(new_n289), .ZN(new_n290));
  OAI21_X1  g089(.A(new_n287), .B1(KEYINPUT22), .B2(new_n290), .ZN(new_n291));
  XOR2_X1   g090(.A(G211gat), .B(G218gat), .Z(new_n292));
  XOR2_X1   g091(.A(new_n291), .B(new_n292), .Z(new_n293));
  INV_X1    g092(.A(KEYINPUT73), .ZN(new_n294));
  NAND2_X1  g093(.A1(new_n293), .A2(new_n294), .ZN(new_n295));
  NAND3_X1  g094(.A1(new_n291), .A2(KEYINPUT73), .A3(new_n292), .ZN(new_n296));
  INV_X1    g095(.A(KEYINPUT29), .ZN(new_n297));
  INV_X1    g096(.A(KEYINPUT3), .ZN(new_n298));
  NAND2_X1  g097(.A1(G155gat), .A2(G162gat), .ZN(new_n299));
  NAND2_X1  g098(.A1(new_n299), .A2(KEYINPUT2), .ZN(new_n300));
  INV_X1    g099(.A(G141gat), .ZN(new_n301));
  INV_X1    g100(.A(G148gat), .ZN(new_n302));
  NAND2_X1  g101(.A1(new_n301), .A2(new_n302), .ZN(new_n303));
  NAND2_X1  g102(.A1(G141gat), .A2(G148gat), .ZN(new_n304));
  NAND3_X1  g103(.A1(new_n300), .A2(new_n303), .A3(new_n304), .ZN(new_n305));
  XNOR2_X1  g104(.A(G155gat), .B(G162gat), .ZN(new_n306));
  INV_X1    g105(.A(KEYINPUT76), .ZN(new_n307));
  OAI21_X1  g106(.A(new_n307), .B1(G155gat), .B2(G162gat), .ZN(new_n308));
  AND3_X1   g107(.A1(new_n305), .A2(new_n306), .A3(new_n308), .ZN(new_n309));
  AOI21_X1  g108(.A(new_n306), .B1(new_n305), .B2(new_n308), .ZN(new_n310));
  OAI21_X1  g109(.A(new_n298), .B1(new_n309), .B2(new_n310), .ZN(new_n311));
  AOI22_X1  g110(.A1(new_n295), .A2(new_n296), .B1(new_n297), .B2(new_n311), .ZN(new_n312));
  INV_X1    g111(.A(G228gat), .ZN(new_n313));
  INV_X1    g112(.A(G233gat), .ZN(new_n314));
  NOR3_X1   g113(.A1(new_n312), .A2(new_n313), .A3(new_n314), .ZN(new_n315));
  NAND2_X1  g114(.A1(new_n295), .A2(new_n296), .ZN(new_n316));
  INV_X1    g115(.A(new_n316), .ZN(new_n317));
  AOI21_X1  g116(.A(KEYINPUT3), .B1(new_n317), .B2(new_n297), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n305), .A2(new_n308), .ZN(new_n319));
  INV_X1    g118(.A(new_n306), .ZN(new_n320));
  NAND2_X1  g119(.A1(new_n319), .A2(new_n320), .ZN(new_n321));
  NAND3_X1  g120(.A1(new_n305), .A2(new_n306), .A3(new_n308), .ZN(new_n322));
  NAND2_X1  g121(.A1(new_n321), .A2(new_n322), .ZN(new_n323));
  OAI21_X1  g122(.A(new_n315), .B1(new_n318), .B2(new_n323), .ZN(new_n324));
  OR2_X1    g123(.A1(new_n293), .A2(KEYINPUT29), .ZN(new_n325));
  AOI21_X1  g124(.A(new_n323), .B1(new_n325), .B2(new_n298), .ZN(new_n326));
  OAI22_X1  g125(.A1(new_n326), .A2(new_n312), .B1(new_n313), .B2(new_n314), .ZN(new_n327));
  AND2_X1   g126(.A1(new_n327), .A2(KEYINPUT79), .ZN(new_n328));
  NOR2_X1   g127(.A1(new_n327), .A2(KEYINPUT79), .ZN(new_n329));
  OAI21_X1  g128(.A(new_n324), .B1(new_n328), .B2(new_n329), .ZN(new_n330));
  XOR2_X1   g129(.A(G78gat), .B(G106gat), .Z(new_n331));
  XNOR2_X1  g130(.A(new_n331), .B(G22gat), .ZN(new_n332));
  XNOR2_X1  g131(.A(KEYINPUT31), .B(G50gat), .ZN(new_n333));
  XOR2_X1   g132(.A(new_n332), .B(new_n333), .Z(new_n334));
  INV_X1    g133(.A(new_n334), .ZN(new_n335));
  NAND2_X1  g134(.A1(new_n330), .A2(new_n335), .ZN(new_n336));
  OAI211_X1 g135(.A(new_n324), .B(new_n334), .C1(new_n328), .C2(new_n329), .ZN(new_n337));
  NAND2_X1  g136(.A1(new_n336), .A2(new_n337), .ZN(new_n338));
  INV_X1    g137(.A(KEYINPUT82), .ZN(new_n339));
  AND3_X1   g138(.A1(new_n266), .A2(new_n282), .A3(new_n277), .ZN(new_n340));
  OAI21_X1  g139(.A(new_n339), .B1(new_n340), .B2(new_n283), .ZN(new_n341));
  AND3_X1   g140(.A1(new_n286), .A2(new_n338), .A3(new_n341), .ZN(new_n342));
  XOR2_X1   g141(.A(G8gat), .B(G36gat), .Z(new_n343));
  XNOR2_X1  g142(.A(G64gat), .B(G92gat), .ZN(new_n344));
  XNOR2_X1  g143(.A(new_n343), .B(new_n344), .ZN(new_n345));
  XOR2_X1   g144(.A(new_n345), .B(KEYINPUT75), .Z(new_n346));
  NAND2_X1  g145(.A1(G226gat), .A2(G233gat), .ZN(new_n347));
  INV_X1    g146(.A(new_n347), .ZN(new_n348));
  NOR2_X1   g147(.A1(new_n348), .A2(KEYINPUT29), .ZN(new_n349));
  NAND2_X1  g148(.A1(new_n249), .A2(new_n349), .ZN(new_n350));
  INV_X1    g149(.A(KEYINPUT74), .ZN(new_n351));
  AOI221_X4 g150(.A(new_n351), .B1(new_n219), .B2(new_n224), .C1(new_n242), .C2(new_n246), .ZN(new_n352));
  NAND2_X1  g151(.A1(new_n242), .A2(new_n246), .ZN(new_n353));
  AOI21_X1  g152(.A(KEYINPUT74), .B1(new_n353), .B2(new_n225), .ZN(new_n354));
  OAI21_X1  g153(.A(new_n348), .B1(new_n352), .B2(new_n354), .ZN(new_n355));
  AND3_X1   g154(.A1(new_n350), .A2(new_n355), .A3(new_n316), .ZN(new_n356));
  INV_X1    g155(.A(new_n354), .ZN(new_n357));
  NAND3_X1  g156(.A1(new_n353), .A2(KEYINPUT74), .A3(new_n225), .ZN(new_n358));
  NAND3_X1  g157(.A1(new_n357), .A2(new_n358), .A3(new_n349), .ZN(new_n359));
  OAI211_X1 g158(.A(new_n348), .B(new_n225), .C1(new_n247), .C2(new_n248), .ZN(new_n360));
  AOI21_X1  g159(.A(new_n316), .B1(new_n359), .B2(new_n360), .ZN(new_n361));
  OAI21_X1  g160(.A(new_n346), .B1(new_n356), .B2(new_n361), .ZN(new_n362));
  NAND3_X1  g161(.A1(new_n350), .A2(new_n355), .A3(new_n316), .ZN(new_n363));
  NOR2_X1   g162(.A1(new_n352), .A2(new_n354), .ZN(new_n364));
  INV_X1    g163(.A(new_n225), .ZN(new_n365));
  INV_X1    g164(.A(KEYINPUT67), .ZN(new_n366));
  NAND2_X1  g165(.A1(new_n353), .A2(new_n366), .ZN(new_n367));
  NAND3_X1  g166(.A1(new_n242), .A2(KEYINPUT67), .A3(new_n246), .ZN(new_n368));
  AOI21_X1  g167(.A(new_n365), .B1(new_n367), .B2(new_n368), .ZN(new_n369));
  AOI22_X1  g168(.A1(new_n364), .A2(new_n349), .B1(new_n369), .B2(new_n348), .ZN(new_n370));
  OAI211_X1 g169(.A(new_n363), .B(new_n345), .C1(new_n370), .C2(new_n316), .ZN(new_n371));
  NAND3_X1  g170(.A1(new_n362), .A2(KEYINPUT30), .A3(new_n371), .ZN(new_n372));
  NAND2_X1  g171(.A1(new_n359), .A2(new_n360), .ZN(new_n373));
  NAND2_X1  g172(.A1(new_n373), .A2(new_n317), .ZN(new_n374));
  INV_X1    g173(.A(KEYINPUT30), .ZN(new_n375));
  NAND4_X1  g174(.A1(new_n374), .A2(new_n375), .A3(new_n363), .A4(new_n345), .ZN(new_n376));
  NAND2_X1  g175(.A1(new_n372), .A2(new_n376), .ZN(new_n377));
  XNOR2_X1  g176(.A(KEYINPUT77), .B(KEYINPUT6), .ZN(new_n378));
  INV_X1    g177(.A(new_n378), .ZN(new_n379));
  XNOR2_X1  g178(.A(G1gat), .B(G29gat), .ZN(new_n380));
  INV_X1    g179(.A(G85gat), .ZN(new_n381));
  XNOR2_X1  g180(.A(new_n380), .B(new_n381), .ZN(new_n382));
  XNOR2_X1  g181(.A(KEYINPUT0), .B(G57gat), .ZN(new_n383));
  XNOR2_X1  g182(.A(new_n382), .B(new_n383), .ZN(new_n384));
  INV_X1    g183(.A(new_n384), .ZN(new_n385));
  NAND2_X1  g184(.A1(G225gat), .A2(G233gat), .ZN(new_n386));
  NAND3_X1  g185(.A1(new_n321), .A2(KEYINPUT3), .A3(new_n322), .ZN(new_n387));
  NAND3_X1  g186(.A1(new_n311), .A2(new_n387), .A3(new_n257), .ZN(new_n388));
  NOR2_X1   g187(.A1(new_n309), .A2(new_n310), .ZN(new_n389));
  NOR3_X1   g188(.A1(new_n389), .A2(KEYINPUT4), .A3(new_n257), .ZN(new_n390));
  INV_X1    g189(.A(KEYINPUT4), .ZN(new_n391));
  AOI21_X1  g190(.A(new_n391), .B1(new_n323), .B2(new_n260), .ZN(new_n392));
  OAI211_X1 g191(.A(new_n386), .B(new_n388), .C1(new_n390), .C2(new_n392), .ZN(new_n393));
  INV_X1    g192(.A(KEYINPUT5), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n393), .A2(new_n394), .ZN(new_n395));
  NAND2_X1  g194(.A1(new_n389), .A2(new_n257), .ZN(new_n396));
  NAND2_X1  g195(.A1(new_n323), .A2(new_n260), .ZN(new_n397));
  NAND2_X1  g196(.A1(new_n396), .A2(new_n397), .ZN(new_n398));
  INV_X1    g197(.A(new_n386), .ZN(new_n399));
  NAND2_X1  g198(.A1(new_n398), .A2(new_n399), .ZN(new_n400));
  AND2_X1   g199(.A1(new_n393), .A2(new_n400), .ZN(new_n401));
  OAI211_X1 g200(.A(new_n385), .B(new_n395), .C1(new_n401), .C2(new_n394), .ZN(new_n402));
  INV_X1    g201(.A(new_n395), .ZN(new_n403));
  AOI21_X1  g202(.A(new_n394), .B1(new_n393), .B2(new_n400), .ZN(new_n404));
  OAI21_X1  g203(.A(new_n384), .B1(new_n403), .B2(new_n404), .ZN(new_n405));
  AOI21_X1  g204(.A(new_n379), .B1(new_n402), .B2(new_n405), .ZN(new_n406));
  AND2_X1   g205(.A1(new_n402), .A2(new_n379), .ZN(new_n407));
  NOR2_X1   g206(.A1(new_n406), .A2(new_n407), .ZN(new_n408));
  NAND2_X1  g207(.A1(new_n377), .A2(new_n408), .ZN(new_n409));
  NOR2_X1   g208(.A1(new_n409), .A2(KEYINPUT35), .ZN(new_n410));
  INV_X1    g209(.A(KEYINPUT78), .ZN(new_n411));
  NAND2_X1  g210(.A1(new_n409), .A2(new_n411), .ZN(new_n412));
  NAND3_X1  g211(.A1(new_n282), .A2(new_n277), .A3(KEYINPUT72), .ZN(new_n413));
  INV_X1    g212(.A(new_n266), .ZN(new_n414));
  NAND2_X1  g213(.A1(new_n413), .A2(new_n414), .ZN(new_n415));
  NAND4_X1  g214(.A1(new_n266), .A2(new_n282), .A3(new_n277), .A4(KEYINPUT72), .ZN(new_n416));
  NAND2_X1  g215(.A1(new_n415), .A2(new_n416), .ZN(new_n417));
  NAND3_X1  g216(.A1(new_n377), .A2(new_n408), .A3(KEYINPUT78), .ZN(new_n418));
  NAND4_X1  g217(.A1(new_n412), .A2(new_n417), .A3(new_n338), .A4(new_n418), .ZN(new_n419));
  AOI22_X1  g218(.A1(new_n342), .A2(new_n410), .B1(new_n419), .B2(KEYINPUT35), .ZN(new_n420));
  INV_X1    g219(.A(new_n338), .ZN(new_n421));
  NAND3_X1  g220(.A1(new_n412), .A2(new_n421), .A3(new_n418), .ZN(new_n422));
  OAI21_X1  g221(.A(new_n388), .B1(new_n390), .B2(new_n392), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n423), .A2(new_n399), .ZN(new_n424));
  NAND3_X1  g223(.A1(new_n396), .A2(new_n397), .A3(new_n386), .ZN(new_n425));
  NAND3_X1  g224(.A1(new_n424), .A2(KEYINPUT39), .A3(new_n425), .ZN(new_n426));
  INV_X1    g225(.A(KEYINPUT39), .ZN(new_n427));
  NAND3_X1  g226(.A1(new_n423), .A2(new_n427), .A3(new_n399), .ZN(new_n428));
  NAND4_X1  g227(.A1(new_n426), .A2(KEYINPUT40), .A3(new_n384), .A4(new_n428), .ZN(new_n429));
  NAND2_X1  g228(.A1(new_n429), .A2(new_n402), .ZN(new_n430));
  AND2_X1   g229(.A1(new_n428), .A2(new_n384), .ZN(new_n431));
  AOI21_X1  g230(.A(KEYINPUT40), .B1(new_n431), .B2(new_n426), .ZN(new_n432));
  NOR2_X1   g231(.A1(new_n430), .A2(new_n432), .ZN(new_n433));
  AND3_X1   g232(.A1(new_n433), .A2(new_n372), .A3(new_n376), .ZN(new_n434));
  NAND3_X1  g233(.A1(new_n350), .A2(new_n355), .A3(new_n317), .ZN(new_n435));
  OAI211_X1 g234(.A(new_n435), .B(KEYINPUT37), .C1(new_n370), .C2(new_n317), .ZN(new_n436));
  NAND2_X1  g235(.A1(new_n436), .A2(new_n346), .ZN(new_n437));
  INV_X1    g236(.A(KEYINPUT37), .ZN(new_n438));
  OAI211_X1 g237(.A(new_n363), .B(new_n438), .C1(new_n370), .C2(new_n316), .ZN(new_n439));
  NAND2_X1  g238(.A1(new_n439), .A2(KEYINPUT81), .ZN(new_n440));
  INV_X1    g239(.A(KEYINPUT81), .ZN(new_n441));
  NAND4_X1  g240(.A1(new_n374), .A2(new_n441), .A3(new_n438), .A4(new_n363), .ZN(new_n442));
  AOI21_X1  g241(.A(new_n437), .B1(new_n440), .B2(new_n442), .ZN(new_n443));
  XNOR2_X1  g242(.A(KEYINPUT80), .B(KEYINPUT38), .ZN(new_n444));
  INV_X1    g243(.A(new_n444), .ZN(new_n445));
  NAND2_X1  g244(.A1(new_n371), .A2(new_n445), .ZN(new_n446));
  AND2_X1   g245(.A1(new_n440), .A2(new_n442), .ZN(new_n447));
  OAI21_X1  g246(.A(KEYINPUT37), .B1(new_n356), .B2(new_n361), .ZN(new_n448));
  NOR2_X1   g247(.A1(new_n345), .A2(new_n445), .ZN(new_n449));
  NAND2_X1  g248(.A1(new_n448), .A2(new_n449), .ZN(new_n450));
  OAI22_X1  g249(.A1(new_n443), .A2(new_n446), .B1(new_n447), .B2(new_n450), .ZN(new_n451));
  INV_X1    g250(.A(new_n408), .ZN(new_n452));
  AOI21_X1  g251(.A(new_n434), .B1(new_n451), .B2(new_n452), .ZN(new_n453));
  OAI21_X1  g252(.A(new_n422), .B1(new_n453), .B2(new_n421), .ZN(new_n454));
  NAND3_X1  g253(.A1(new_n415), .A2(KEYINPUT36), .A3(new_n416), .ZN(new_n455));
  INV_X1    g254(.A(KEYINPUT36), .ZN(new_n456));
  OAI21_X1  g255(.A(new_n456), .B1(new_n340), .B2(new_n283), .ZN(new_n457));
  NAND2_X1  g256(.A1(new_n455), .A2(new_n457), .ZN(new_n458));
  INV_X1    g257(.A(new_n458), .ZN(new_n459));
  AOI21_X1  g258(.A(new_n420), .B1(new_n454), .B2(new_n459), .ZN(new_n460));
  INV_X1    g259(.A(G29gat), .ZN(new_n461));
  INV_X1    g260(.A(G36gat), .ZN(new_n462));
  AOI21_X1  g261(.A(KEYINPUT14), .B1(new_n461), .B2(new_n462), .ZN(new_n463));
  XNOR2_X1  g262(.A(KEYINPUT84), .B(G29gat), .ZN(new_n464));
  NAND2_X1  g263(.A1(new_n464), .A2(G36gat), .ZN(new_n465));
  NAND2_X1  g264(.A1(new_n461), .A2(new_n462), .ZN(new_n466));
  NAND2_X1  g265(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  AOI21_X1  g266(.A(new_n463), .B1(new_n467), .B2(KEYINPUT14), .ZN(new_n468));
  XNOR2_X1  g267(.A(G43gat), .B(G50gat), .ZN(new_n469));
  INV_X1    g268(.A(KEYINPUT83), .ZN(new_n470));
  AND2_X1   g269(.A1(new_n469), .A2(new_n470), .ZN(new_n471));
  OAI21_X1  g270(.A(KEYINPUT15), .B1(new_n469), .B2(new_n470), .ZN(new_n472));
  OAI22_X1  g271(.A1(new_n471), .A2(new_n472), .B1(KEYINPUT15), .B2(new_n469), .ZN(new_n473));
  NAND2_X1  g272(.A1(new_n468), .A2(new_n473), .ZN(new_n474));
  INV_X1    g273(.A(KEYINPUT14), .ZN(new_n475));
  AOI21_X1  g274(.A(new_n475), .B1(new_n465), .B2(new_n466), .ZN(new_n476));
  OAI22_X1  g275(.A1(new_n476), .A2(new_n463), .B1(new_n471), .B2(new_n472), .ZN(new_n477));
  NAND2_X1  g276(.A1(new_n474), .A2(new_n477), .ZN(new_n478));
  NAND2_X1  g277(.A1(new_n478), .A2(KEYINPUT85), .ZN(new_n479));
  INV_X1    g278(.A(KEYINPUT86), .ZN(new_n480));
  INV_X1    g279(.A(KEYINPUT17), .ZN(new_n481));
  INV_X1    g280(.A(KEYINPUT85), .ZN(new_n482));
  NAND3_X1  g281(.A1(new_n474), .A2(new_n482), .A3(new_n477), .ZN(new_n483));
  NAND4_X1  g282(.A1(new_n479), .A2(new_n480), .A3(new_n481), .A4(new_n483), .ZN(new_n484));
  AND3_X1   g283(.A1(new_n474), .A2(new_n482), .A3(new_n477), .ZN(new_n485));
  AOI21_X1  g284(.A(new_n482), .B1(new_n474), .B2(new_n477), .ZN(new_n486));
  NOR3_X1   g285(.A1(new_n485), .A2(new_n486), .A3(KEYINPUT17), .ZN(new_n487));
  AOI21_X1  g286(.A(new_n480), .B1(new_n478), .B2(KEYINPUT17), .ZN(new_n488));
  INV_X1    g287(.A(new_n488), .ZN(new_n489));
  OAI21_X1  g288(.A(new_n484), .B1(new_n487), .B2(new_n489), .ZN(new_n490));
  XNOR2_X1  g289(.A(G15gat), .B(G22gat), .ZN(new_n491));
  AND2_X1   g290(.A1(new_n491), .A2(KEYINPUT87), .ZN(new_n492));
  OR2_X1    g291(.A1(new_n492), .A2(G1gat), .ZN(new_n493));
  NAND2_X1  g292(.A1(new_n492), .A2(G1gat), .ZN(new_n494));
  INV_X1    g293(.A(KEYINPUT16), .ZN(new_n495));
  NAND2_X1  g294(.A1(new_n491), .A2(new_n495), .ZN(new_n496));
  NAND3_X1  g295(.A1(new_n493), .A2(new_n494), .A3(new_n496), .ZN(new_n497));
  XNOR2_X1  g296(.A(new_n497), .B(G8gat), .ZN(new_n498));
  INV_X1    g297(.A(new_n498), .ZN(new_n499));
  NAND2_X1  g298(.A1(new_n490), .A2(new_n499), .ZN(new_n500));
  INV_X1    g299(.A(KEYINPUT88), .ZN(new_n501));
  INV_X1    g300(.A(KEYINPUT18), .ZN(new_n502));
  NAND2_X1  g301(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  NAND2_X1  g302(.A1(G229gat), .A2(G233gat), .ZN(new_n504));
  NAND2_X1  g303(.A1(new_n479), .A2(new_n483), .ZN(new_n505));
  NOR2_X1   g304(.A1(new_n499), .A2(new_n505), .ZN(new_n506));
  INV_X1    g305(.A(new_n506), .ZN(new_n507));
  NAND4_X1  g306(.A1(new_n500), .A2(new_n503), .A3(new_n504), .A4(new_n507), .ZN(new_n508));
  NOR2_X1   g307(.A1(new_n501), .A2(new_n502), .ZN(new_n509));
  INV_X1    g308(.A(new_n509), .ZN(new_n510));
  NAND2_X1  g309(.A1(new_n508), .A2(new_n510), .ZN(new_n511));
  NAND2_X1  g310(.A1(new_n499), .A2(new_n505), .ZN(new_n512));
  NAND2_X1  g311(.A1(new_n507), .A2(new_n512), .ZN(new_n513));
  XOR2_X1   g312(.A(new_n504), .B(KEYINPUT13), .Z(new_n514));
  NAND2_X1  g313(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  NAND4_X1  g314(.A1(new_n500), .A2(new_n509), .A3(new_n504), .A4(new_n507), .ZN(new_n516));
  XNOR2_X1  g315(.A(G113gat), .B(G141gat), .ZN(new_n517));
  INV_X1    g316(.A(G197gat), .ZN(new_n518));
  XNOR2_X1  g317(.A(new_n517), .B(new_n518), .ZN(new_n519));
  XNOR2_X1  g318(.A(KEYINPUT11), .B(G169gat), .ZN(new_n520));
  XNOR2_X1  g319(.A(new_n519), .B(new_n520), .ZN(new_n521));
  XNOR2_X1  g320(.A(new_n521), .B(KEYINPUT12), .ZN(new_n522));
  NAND4_X1  g321(.A1(new_n511), .A2(new_n515), .A3(new_n516), .A4(new_n522), .ZN(new_n523));
  INV_X1    g322(.A(new_n523), .ZN(new_n524));
  AND2_X1   g323(.A1(new_n516), .A2(new_n515), .ZN(new_n525));
  AOI21_X1  g324(.A(new_n522), .B1(new_n525), .B2(new_n511), .ZN(new_n526));
  NOR2_X1   g325(.A1(new_n524), .A2(new_n526), .ZN(new_n527));
  NOR3_X1   g326(.A1(new_n460), .A2(KEYINPUT89), .A3(new_n527), .ZN(new_n528));
  INV_X1    g327(.A(KEYINPUT89), .ZN(new_n529));
  INV_X1    g328(.A(new_n420), .ZN(new_n530));
  NAND2_X1  g329(.A1(new_n454), .A2(new_n459), .ZN(new_n531));
  NAND2_X1  g330(.A1(new_n530), .A2(new_n531), .ZN(new_n532));
  INV_X1    g331(.A(new_n527), .ZN(new_n533));
  AOI21_X1  g332(.A(new_n529), .B1(new_n532), .B2(new_n533), .ZN(new_n534));
  NOR2_X1   g333(.A1(new_n528), .A2(new_n534), .ZN(new_n535));
  XNOR2_X1  g334(.A(G71gat), .B(G78gat), .ZN(new_n536));
  AOI21_X1  g335(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n537));
  XNOR2_X1  g336(.A(KEYINPUT90), .B(G57gat), .ZN(new_n538));
  NAND2_X1  g337(.A1(new_n538), .A2(G64gat), .ZN(new_n539));
  INV_X1    g338(.A(G64gat), .ZN(new_n540));
  NAND2_X1  g339(.A1(new_n540), .A2(G57gat), .ZN(new_n541));
  AOI21_X1  g340(.A(new_n537), .B1(new_n539), .B2(new_n541), .ZN(new_n542));
  INV_X1    g341(.A(KEYINPUT91), .ZN(new_n543));
  NAND2_X1  g342(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  NAND2_X1  g343(.A1(new_n542), .A2(KEYINPUT91), .ZN(new_n545));
  INV_X1    g344(.A(KEYINPUT9), .ZN(new_n546));
  OR2_X1    g345(.A1(new_n540), .A2(G57gat), .ZN(new_n547));
  AOI211_X1 g346(.A(new_n546), .B(new_n536), .C1(new_n541), .C2(new_n547), .ZN(new_n548));
  AOI22_X1  g347(.A1(new_n536), .A2(new_n544), .B1(new_n545), .B2(new_n548), .ZN(new_n549));
  XOR2_X1   g348(.A(KEYINPUT92), .B(KEYINPUT21), .Z(new_n550));
  NAND2_X1  g349(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  INV_X1    g350(.A(G127gat), .ZN(new_n552));
  XNOR2_X1  g351(.A(new_n551), .B(new_n552), .ZN(new_n553));
  INV_X1    g352(.A(G155gat), .ZN(new_n554));
  XNOR2_X1  g353(.A(new_n553), .B(new_n554), .ZN(new_n555));
  XNOR2_X1  g354(.A(G183gat), .B(G211gat), .ZN(new_n556));
  XNOR2_X1  g355(.A(new_n556), .B(KEYINPUT93), .ZN(new_n557));
  NAND2_X1  g356(.A1(G231gat), .A2(G233gat), .ZN(new_n558));
  XOR2_X1   g357(.A(new_n557), .B(new_n558), .Z(new_n559));
  XNOR2_X1  g358(.A(new_n555), .B(new_n559), .ZN(new_n560));
  INV_X1    g359(.A(KEYINPUT21), .ZN(new_n561));
  OAI21_X1  g360(.A(new_n499), .B1(new_n549), .B2(new_n561), .ZN(new_n562));
  XNOR2_X1  g361(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n563));
  XNOR2_X1  g362(.A(new_n562), .B(new_n563), .ZN(new_n564));
  XNOR2_X1  g363(.A(new_n560), .B(new_n564), .ZN(new_n565));
  XNOR2_X1  g364(.A(KEYINPUT95), .B(KEYINPUT7), .ZN(new_n566));
  INV_X1    g365(.A(G92gat), .ZN(new_n567));
  OR3_X1    g366(.A1(new_n566), .A2(new_n381), .A3(new_n567), .ZN(new_n568));
  OAI21_X1  g367(.A(new_n566), .B1(new_n381), .B2(new_n567), .ZN(new_n569));
  NAND2_X1  g368(.A1(G99gat), .A2(G106gat), .ZN(new_n570));
  AOI22_X1  g369(.A1(KEYINPUT8), .A2(new_n570), .B1(new_n381), .B2(new_n567), .ZN(new_n571));
  NAND3_X1  g370(.A1(new_n568), .A2(new_n569), .A3(new_n571), .ZN(new_n572));
  XOR2_X1   g371(.A(G99gat), .B(G106gat), .Z(new_n573));
  XNOR2_X1  g372(.A(new_n572), .B(new_n573), .ZN(new_n574));
  INV_X1    g373(.A(new_n574), .ZN(new_n575));
  NAND3_X1  g374(.A1(new_n479), .A2(new_n481), .A3(new_n483), .ZN(new_n576));
  NAND2_X1  g375(.A1(new_n576), .A2(new_n488), .ZN(new_n577));
  AOI21_X1  g376(.A(new_n575), .B1(new_n577), .B2(new_n484), .ZN(new_n578));
  XOR2_X1   g377(.A(G190gat), .B(G218gat), .Z(new_n579));
  NAND2_X1  g378(.A1(G232gat), .A2(G233gat), .ZN(new_n580));
  INV_X1    g379(.A(new_n580), .ZN(new_n581));
  NAND2_X1  g380(.A1(new_n581), .A2(KEYINPUT41), .ZN(new_n582));
  OAI21_X1  g381(.A(new_n582), .B1(new_n505), .B2(new_n574), .ZN(new_n583));
  OR3_X1    g382(.A1(new_n578), .A2(new_n579), .A3(new_n583), .ZN(new_n584));
  NOR2_X1   g383(.A1(new_n581), .A2(KEYINPUT41), .ZN(new_n585));
  XNOR2_X1  g384(.A(new_n585), .B(KEYINPUT94), .ZN(new_n586));
  XNOR2_X1  g385(.A(G134gat), .B(G162gat), .ZN(new_n587));
  XNOR2_X1  g386(.A(new_n586), .B(new_n587), .ZN(new_n588));
  OAI21_X1  g387(.A(new_n579), .B1(new_n578), .B2(new_n583), .ZN(new_n589));
  NAND3_X1  g388(.A1(new_n584), .A2(new_n588), .A3(new_n589), .ZN(new_n590));
  INV_X1    g389(.A(new_n590), .ZN(new_n591));
  AOI21_X1  g390(.A(new_n588), .B1(new_n584), .B2(new_n589), .ZN(new_n592));
  NOR2_X1   g391(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  INV_X1    g392(.A(new_n593), .ZN(new_n594));
  NAND2_X1  g393(.A1(new_n565), .A2(new_n594), .ZN(new_n595));
  XNOR2_X1  g394(.A(G120gat), .B(G148gat), .ZN(new_n596));
  XNOR2_X1  g395(.A(G176gat), .B(G204gat), .ZN(new_n597));
  XNOR2_X1  g396(.A(new_n596), .B(new_n597), .ZN(new_n598));
  NOR2_X1   g397(.A1(new_n574), .A2(new_n549), .ZN(new_n599));
  INV_X1    g398(.A(new_n599), .ZN(new_n600));
  NAND3_X1  g399(.A1(new_n600), .A2(KEYINPUT96), .A3(KEYINPUT10), .ZN(new_n601));
  INV_X1    g400(.A(new_n601), .ZN(new_n602));
  INV_X1    g401(.A(KEYINPUT10), .ZN(new_n603));
  INV_X1    g402(.A(KEYINPUT96), .ZN(new_n604));
  OAI21_X1  g403(.A(new_n603), .B1(new_n599), .B2(new_n604), .ZN(new_n605));
  NAND2_X1  g404(.A1(new_n574), .A2(new_n549), .ZN(new_n606));
  NAND2_X1  g405(.A1(new_n605), .A2(new_n606), .ZN(new_n607));
  NAND2_X1  g406(.A1(G230gat), .A2(G233gat), .ZN(new_n608));
  XOR2_X1   g407(.A(new_n608), .B(KEYINPUT97), .Z(new_n609));
  INV_X1    g408(.A(new_n609), .ZN(new_n610));
  NOR3_X1   g409(.A1(new_n602), .A2(new_n607), .A3(new_n610), .ZN(new_n611));
  AOI21_X1  g410(.A(new_n608), .B1(new_n600), .B2(new_n606), .ZN(new_n612));
  OAI21_X1  g411(.A(new_n598), .B1(new_n611), .B2(new_n612), .ZN(new_n613));
  NAND4_X1  g412(.A1(new_n601), .A2(new_n605), .A3(new_n606), .A4(new_n608), .ZN(new_n614));
  NOR2_X1   g413(.A1(new_n612), .A2(new_n598), .ZN(new_n615));
  NAND2_X1  g414(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  NAND2_X1  g415(.A1(new_n613), .A2(new_n616), .ZN(new_n617));
  NOR3_X1   g416(.A1(new_n535), .A2(new_n595), .A3(new_n617), .ZN(new_n618));
  NAND2_X1  g417(.A1(new_n618), .A2(new_n452), .ZN(new_n619));
  XOR2_X1   g418(.A(KEYINPUT98), .B(G1gat), .Z(new_n620));
  XNOR2_X1  g419(.A(new_n619), .B(new_n620), .ZN(G1324gat));
  INV_X1    g420(.A(new_n377), .ZN(new_n622));
  NAND2_X1  g421(.A1(new_n618), .A2(new_n622), .ZN(new_n623));
  INV_X1    g422(.A(KEYINPUT42), .ZN(new_n624));
  XNOR2_X1  g423(.A(KEYINPUT16), .B(G8gat), .ZN(new_n625));
  NOR3_X1   g424(.A1(new_n623), .A2(new_n624), .A3(new_n625), .ZN(new_n626));
  AOI21_X1  g425(.A(new_n626), .B1(G8gat), .B2(new_n623), .ZN(new_n627));
  OAI21_X1  g426(.A(new_n624), .B1(new_n623), .B2(new_n625), .ZN(new_n628));
  INV_X1    g427(.A(KEYINPUT99), .ZN(new_n629));
  OR2_X1    g428(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  NAND2_X1  g429(.A1(new_n628), .A2(new_n629), .ZN(new_n631));
  NAND3_X1  g430(.A1(new_n627), .A2(new_n630), .A3(new_n631), .ZN(G1325gat));
  AND2_X1   g431(.A1(new_n286), .A2(new_n341), .ZN(new_n633));
  AOI21_X1  g432(.A(G15gat), .B1(new_n618), .B2(new_n633), .ZN(new_n634));
  INV_X1    g433(.A(KEYINPUT100), .ZN(new_n635));
  AND3_X1   g434(.A1(new_n455), .A2(new_n457), .A3(new_n635), .ZN(new_n636));
  INV_X1    g435(.A(new_n636), .ZN(new_n637));
  AOI21_X1  g436(.A(new_n635), .B1(new_n455), .B2(new_n457), .ZN(new_n638));
  INV_X1    g437(.A(new_n638), .ZN(new_n639));
  NAND2_X1  g438(.A1(new_n637), .A2(new_n639), .ZN(new_n640));
  INV_X1    g439(.A(new_n640), .ZN(new_n641));
  AND2_X1   g440(.A1(new_n641), .A2(G15gat), .ZN(new_n642));
  AOI21_X1  g441(.A(new_n634), .B1(new_n618), .B2(new_n642), .ZN(G1326gat));
  NAND2_X1  g442(.A1(new_n618), .A2(new_n421), .ZN(new_n644));
  XNOR2_X1  g443(.A(new_n644), .B(KEYINPUT101), .ZN(new_n645));
  XNOR2_X1  g444(.A(KEYINPUT43), .B(G22gat), .ZN(new_n646));
  XNOR2_X1  g445(.A(new_n645), .B(new_n646), .ZN(G1327gat));
  NOR2_X1   g446(.A1(new_n565), .A2(new_n617), .ZN(new_n648));
  INV_X1    g447(.A(new_n648), .ZN(new_n649));
  NOR3_X1   g448(.A1(new_n535), .A2(new_n594), .A3(new_n649), .ZN(new_n650));
  NOR2_X1   g449(.A1(new_n408), .A2(new_n464), .ZN(new_n651));
  NAND2_X1  g450(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  NAND2_X1  g451(.A1(new_n652), .A2(KEYINPUT45), .ZN(new_n653));
  OR2_X1    g452(.A1(new_n652), .A2(KEYINPUT45), .ZN(new_n654));
  OAI21_X1  g453(.A(KEYINPUT44), .B1(new_n460), .B2(new_n594), .ZN(new_n655));
  INV_X1    g454(.A(new_n655), .ZN(new_n656));
  NAND2_X1  g455(.A1(new_n440), .A2(new_n442), .ZN(new_n657));
  INV_X1    g456(.A(new_n437), .ZN(new_n658));
  AOI21_X1  g457(.A(new_n446), .B1(new_n657), .B2(new_n658), .ZN(new_n659));
  AOI21_X1  g458(.A(new_n450), .B1(new_n440), .B2(new_n442), .ZN(new_n660));
  OAI21_X1  g459(.A(new_n452), .B1(new_n659), .B2(new_n660), .ZN(new_n661));
  INV_X1    g460(.A(new_n434), .ZN(new_n662));
  AOI21_X1  g461(.A(new_n421), .B1(new_n661), .B2(new_n662), .ZN(new_n663));
  AND3_X1   g462(.A1(new_n377), .A2(new_n408), .A3(KEYINPUT78), .ZN(new_n664));
  AOI21_X1  g463(.A(KEYINPUT78), .B1(new_n377), .B2(new_n408), .ZN(new_n665));
  NOR3_X1   g464(.A1(new_n664), .A2(new_n665), .A3(new_n338), .ZN(new_n666));
  OAI22_X1  g465(.A1(new_n636), .A2(new_n638), .B1(new_n663), .B2(new_n666), .ZN(new_n667));
  INV_X1    g466(.A(KEYINPUT103), .ZN(new_n668));
  NAND2_X1  g467(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  OAI211_X1 g468(.A(new_n454), .B(KEYINPUT103), .C1(new_n636), .C2(new_n638), .ZN(new_n670));
  NAND2_X1  g469(.A1(new_n669), .A2(new_n670), .ZN(new_n671));
  NAND2_X1  g470(.A1(new_n671), .A2(new_n530), .ZN(new_n672));
  NAND2_X1  g471(.A1(new_n672), .A2(KEYINPUT104), .ZN(new_n673));
  AOI21_X1  g472(.A(new_n420), .B1(new_n669), .B2(new_n670), .ZN(new_n674));
  INV_X1    g473(.A(KEYINPUT104), .ZN(new_n675));
  NAND2_X1  g474(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  NAND2_X1  g475(.A1(new_n673), .A2(new_n676), .ZN(new_n677));
  NOR2_X1   g476(.A1(new_n593), .A2(KEYINPUT105), .ZN(new_n678));
  INV_X1    g477(.A(KEYINPUT105), .ZN(new_n679));
  NOR3_X1   g478(.A1(new_n591), .A2(new_n592), .A3(new_n679), .ZN(new_n680));
  NOR2_X1   g479(.A1(new_n678), .A2(new_n680), .ZN(new_n681));
  INV_X1    g480(.A(new_n681), .ZN(new_n682));
  NOR2_X1   g481(.A1(new_n682), .A2(KEYINPUT44), .ZN(new_n683));
  AOI21_X1  g482(.A(new_n656), .B1(new_n677), .B2(new_n683), .ZN(new_n684));
  INV_X1    g483(.A(new_n522), .ZN(new_n685));
  AOI21_X1  g484(.A(new_n498), .B1(new_n577), .B2(new_n484), .ZN(new_n686));
  INV_X1    g485(.A(new_n504), .ZN(new_n687));
  NOR3_X1   g486(.A1(new_n686), .A2(new_n687), .A3(new_n506), .ZN(new_n688));
  AOI21_X1  g487(.A(new_n509), .B1(new_n688), .B2(new_n503), .ZN(new_n689));
  NAND2_X1  g488(.A1(new_n516), .A2(new_n515), .ZN(new_n690));
  OAI21_X1  g489(.A(new_n685), .B1(new_n689), .B2(new_n690), .ZN(new_n691));
  INV_X1    g490(.A(KEYINPUT102), .ZN(new_n692));
  AND3_X1   g491(.A1(new_n691), .A2(new_n692), .A3(new_n523), .ZN(new_n693));
  AOI21_X1  g492(.A(new_n692), .B1(new_n691), .B2(new_n523), .ZN(new_n694));
  NOR2_X1   g493(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  NOR3_X1   g494(.A1(new_n684), .A2(new_n649), .A3(new_n695), .ZN(new_n696));
  NAND2_X1  g495(.A1(new_n696), .A2(new_n452), .ZN(new_n697));
  AOI22_X1  g496(.A1(new_n653), .A2(new_n654), .B1(new_n697), .B2(new_n464), .ZN(new_n698));
  INV_X1    g497(.A(KEYINPUT106), .ZN(new_n699));
  XNOR2_X1  g498(.A(new_n698), .B(new_n699), .ZN(G1328gat));
  NAND3_X1  g499(.A1(new_n650), .A2(new_n462), .A3(new_n622), .ZN(new_n701));
  XOR2_X1   g500(.A(new_n701), .B(KEYINPUT46), .Z(new_n702));
  AND2_X1   g501(.A1(new_n696), .A2(new_n622), .ZN(new_n703));
  OAI21_X1  g502(.A(new_n702), .B1(new_n462), .B2(new_n703), .ZN(G1329gat));
  NOR2_X1   g503(.A1(KEYINPUT107), .A2(KEYINPUT47), .ZN(new_n705));
  INV_X1    g504(.A(G43gat), .ZN(new_n706));
  AND2_X1   g505(.A1(new_n633), .A2(new_n706), .ZN(new_n707));
  AOI21_X1  g506(.A(new_n705), .B1(new_n650), .B2(new_n707), .ZN(new_n708));
  AND2_X1   g507(.A1(new_n696), .A2(new_n641), .ZN(new_n709));
  OAI21_X1  g508(.A(new_n708), .B1(new_n709), .B2(new_n706), .ZN(new_n710));
  NAND2_X1  g509(.A1(KEYINPUT107), .A2(KEYINPUT47), .ZN(new_n711));
  XNOR2_X1  g510(.A(new_n710), .B(new_n711), .ZN(G1330gat));
  INV_X1    g511(.A(G50gat), .ZN(new_n713));
  NAND3_X1  g512(.A1(new_n650), .A2(new_n713), .A3(new_n421), .ZN(new_n714));
  NAND2_X1  g513(.A1(new_n696), .A2(new_n421), .ZN(new_n715));
  AND2_X1   g514(.A1(new_n715), .A2(KEYINPUT108), .ZN(new_n716));
  OAI21_X1  g515(.A(G50gat), .B1(new_n715), .B2(KEYINPUT108), .ZN(new_n717));
  OAI211_X1 g516(.A(KEYINPUT48), .B(new_n714), .C1(new_n716), .C2(new_n717), .ZN(new_n718));
  INV_X1    g517(.A(new_n714), .ZN(new_n719));
  AOI21_X1  g518(.A(new_n719), .B1(new_n715), .B2(G50gat), .ZN(new_n720));
  OAI21_X1  g519(.A(new_n718), .B1(KEYINPUT48), .B2(new_n720), .ZN(G1331gat));
  INV_X1    g520(.A(new_n695), .ZN(new_n722));
  INV_X1    g521(.A(new_n617), .ZN(new_n723));
  NOR3_X1   g522(.A1(new_n722), .A2(new_n595), .A3(new_n723), .ZN(new_n724));
  XNOR2_X1  g523(.A(new_n724), .B(KEYINPUT109), .ZN(new_n725));
  AOI21_X1  g524(.A(new_n725), .B1(new_n673), .B2(new_n676), .ZN(new_n726));
  NAND2_X1  g525(.A1(new_n726), .A2(new_n452), .ZN(new_n727));
  XNOR2_X1  g526(.A(new_n727), .B(KEYINPUT110), .ZN(new_n728));
  XOR2_X1   g527(.A(new_n728), .B(new_n538), .Z(G1332gat));
  NAND2_X1  g528(.A1(new_n726), .A2(new_n622), .ZN(new_n730));
  OAI21_X1  g529(.A(new_n730), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n731));
  XOR2_X1   g530(.A(KEYINPUT49), .B(G64gat), .Z(new_n732));
  OAI21_X1  g531(.A(new_n731), .B1(new_n730), .B2(new_n732), .ZN(G1333gat));
  AOI21_X1  g532(.A(G71gat), .B1(new_n726), .B2(new_n633), .ZN(new_n734));
  AND2_X1   g533(.A1(new_n641), .A2(G71gat), .ZN(new_n735));
  AOI21_X1  g534(.A(new_n734), .B1(new_n726), .B2(new_n735), .ZN(new_n736));
  XOR2_X1   g535(.A(new_n736), .B(KEYINPUT50), .Z(G1334gat));
  NAND2_X1  g536(.A1(new_n726), .A2(new_n421), .ZN(new_n738));
  XNOR2_X1  g537(.A(new_n738), .B(G78gat), .ZN(G1335gat));
  INV_X1    g538(.A(KEYINPUT111), .ZN(new_n740));
  AOI21_X1  g539(.A(new_n675), .B1(new_n671), .B2(new_n530), .ZN(new_n741));
  AOI211_X1 g540(.A(KEYINPUT104), .B(new_n420), .C1(new_n669), .C2(new_n670), .ZN(new_n742));
  OAI21_X1  g541(.A(new_n683), .B1(new_n741), .B2(new_n742), .ZN(new_n743));
  NAND2_X1  g542(.A1(new_n743), .A2(new_n655), .ZN(new_n744));
  NOR2_X1   g543(.A1(new_n722), .A2(new_n565), .ZN(new_n745));
  NAND2_X1  g544(.A1(new_n745), .A2(new_n617), .ZN(new_n746));
  INV_X1    g545(.A(new_n746), .ZN(new_n747));
  AOI21_X1  g546(.A(new_n740), .B1(new_n744), .B2(new_n747), .ZN(new_n748));
  INV_X1    g547(.A(new_n748), .ZN(new_n749));
  AOI211_X1 g548(.A(KEYINPUT111), .B(new_n746), .C1(new_n743), .C2(new_n655), .ZN(new_n750));
  INV_X1    g549(.A(new_n750), .ZN(new_n751));
  AOI21_X1  g550(.A(new_n408), .B1(new_n749), .B2(new_n751), .ZN(new_n752));
  NAND3_X1  g551(.A1(new_n672), .A2(KEYINPUT112), .A3(new_n593), .ZN(new_n753));
  INV_X1    g552(.A(KEYINPUT112), .ZN(new_n754));
  OAI21_X1  g553(.A(new_n754), .B1(new_n674), .B2(new_n594), .ZN(new_n755));
  NAND3_X1  g554(.A1(new_n753), .A2(new_n755), .A3(new_n745), .ZN(new_n756));
  INV_X1    g555(.A(KEYINPUT51), .ZN(new_n757));
  NAND2_X1  g556(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  INV_X1    g557(.A(new_n758), .ZN(new_n759));
  NAND4_X1  g558(.A1(new_n753), .A2(new_n755), .A3(KEYINPUT51), .A4(new_n745), .ZN(new_n760));
  INV_X1    g559(.A(new_n760), .ZN(new_n761));
  NOR2_X1   g560(.A1(new_n759), .A2(new_n761), .ZN(new_n762));
  NAND3_X1  g561(.A1(new_n617), .A2(new_n452), .A3(new_n381), .ZN(new_n763));
  XNOR2_X1  g562(.A(new_n763), .B(KEYINPUT113), .ZN(new_n764));
  OAI22_X1  g563(.A1(new_n752), .A2(new_n381), .B1(new_n762), .B2(new_n764), .ZN(G1336gat));
  INV_X1    g564(.A(KEYINPUT52), .ZN(new_n766));
  NOR3_X1   g565(.A1(new_n684), .A2(new_n377), .A3(new_n746), .ZN(new_n767));
  OAI21_X1  g566(.A(new_n617), .B1(new_n759), .B2(new_n761), .ZN(new_n768));
  NOR2_X1   g567(.A1(new_n377), .A2(G92gat), .ZN(new_n769));
  INV_X1    g568(.A(new_n769), .ZN(new_n770));
  OAI221_X1 g569(.A(new_n766), .B1(new_n767), .B2(new_n567), .C1(new_n768), .C2(new_n770), .ZN(new_n771));
  INV_X1    g570(.A(new_n768), .ZN(new_n772));
  OAI21_X1  g571(.A(new_n622), .B1(new_n748), .B2(new_n750), .ZN(new_n773));
  AOI22_X1  g572(.A1(new_n772), .A2(new_n769), .B1(new_n773), .B2(G92gat), .ZN(new_n774));
  OAI21_X1  g573(.A(new_n771), .B1(new_n774), .B2(new_n766), .ZN(G1337gat));
  INV_X1    g574(.A(G99gat), .ZN(new_n776));
  NAND3_X1  g575(.A1(new_n772), .A2(new_n776), .A3(new_n633), .ZN(new_n777));
  AOI21_X1  g576(.A(new_n640), .B1(new_n749), .B2(new_n751), .ZN(new_n778));
  OAI21_X1  g577(.A(new_n777), .B1(new_n778), .B2(new_n776), .ZN(G1338gat));
  NAND3_X1  g578(.A1(new_n744), .A2(new_n421), .A3(new_n747), .ZN(new_n780));
  AOI21_X1  g579(.A(KEYINPUT53), .B1(new_n780), .B2(G106gat), .ZN(new_n781));
  NOR2_X1   g580(.A1(new_n338), .A2(G106gat), .ZN(new_n782));
  INV_X1    g581(.A(new_n782), .ZN(new_n783));
  OAI21_X1  g582(.A(new_n781), .B1(new_n768), .B2(new_n783), .ZN(new_n784));
  AOI211_X1 g583(.A(new_n723), .B(new_n783), .C1(new_n758), .C2(new_n760), .ZN(new_n785));
  OAI21_X1  g584(.A(new_n421), .B1(new_n748), .B2(new_n750), .ZN(new_n786));
  AOI21_X1  g585(.A(new_n785), .B1(new_n786), .B2(G106gat), .ZN(new_n787));
  INV_X1    g586(.A(KEYINPUT53), .ZN(new_n788));
  OAI21_X1  g587(.A(new_n784), .B1(new_n787), .B2(new_n788), .ZN(new_n789));
  NAND2_X1  g588(.A1(new_n789), .A2(KEYINPUT114), .ZN(new_n790));
  INV_X1    g589(.A(KEYINPUT114), .ZN(new_n791));
  OAI211_X1 g590(.A(new_n791), .B(new_n784), .C1(new_n787), .C2(new_n788), .ZN(new_n792));
  NAND2_X1  g591(.A1(new_n790), .A2(new_n792), .ZN(G1339gat));
  OAI21_X1  g592(.A(new_n610), .B1(new_n602), .B2(new_n607), .ZN(new_n794));
  NAND3_X1  g593(.A1(new_n794), .A2(KEYINPUT54), .A3(new_n614), .ZN(new_n795));
  INV_X1    g594(.A(new_n607), .ZN(new_n796));
  INV_X1    g595(.A(KEYINPUT54), .ZN(new_n797));
  NAND4_X1  g596(.A1(new_n796), .A2(new_n797), .A3(new_n609), .A4(new_n601), .ZN(new_n798));
  NAND3_X1  g597(.A1(new_n795), .A2(new_n598), .A3(new_n798), .ZN(new_n799));
  INV_X1    g598(.A(KEYINPUT55), .ZN(new_n800));
  NAND2_X1  g599(.A1(new_n799), .A2(new_n800), .ZN(new_n801));
  NAND4_X1  g600(.A1(new_n795), .A2(KEYINPUT55), .A3(new_n598), .A4(new_n798), .ZN(new_n802));
  NAND3_X1  g601(.A1(new_n801), .A2(new_n616), .A3(new_n802), .ZN(new_n803));
  OAI21_X1  g602(.A(KEYINPUT102), .B1(new_n524), .B2(new_n526), .ZN(new_n804));
  NAND3_X1  g603(.A1(new_n691), .A2(new_n692), .A3(new_n523), .ZN(new_n805));
  AOI21_X1  g604(.A(new_n803), .B1(new_n804), .B2(new_n805), .ZN(new_n806));
  NOR2_X1   g605(.A1(new_n513), .A2(new_n514), .ZN(new_n807));
  AOI21_X1  g606(.A(new_n504), .B1(new_n500), .B2(new_n507), .ZN(new_n808));
  OAI21_X1  g607(.A(new_n521), .B1(new_n807), .B2(new_n808), .ZN(new_n809));
  NAND2_X1  g608(.A1(new_n523), .A2(new_n809), .ZN(new_n810));
  NOR2_X1   g609(.A1(new_n810), .A2(new_n723), .ZN(new_n811));
  OAI21_X1  g610(.A(KEYINPUT116), .B1(new_n806), .B2(new_n811), .ZN(new_n812));
  AND3_X1   g611(.A1(new_n801), .A2(new_n616), .A3(new_n802), .ZN(new_n813));
  OAI21_X1  g612(.A(new_n813), .B1(new_n693), .B2(new_n694), .ZN(new_n814));
  INV_X1    g613(.A(KEYINPUT116), .ZN(new_n815));
  INV_X1    g614(.A(new_n811), .ZN(new_n816));
  NAND3_X1  g615(.A1(new_n814), .A2(new_n815), .A3(new_n816), .ZN(new_n817));
  NAND3_X1  g616(.A1(new_n812), .A2(new_n682), .A3(new_n817), .ZN(new_n818));
  OR2_X1    g617(.A1(new_n810), .A2(KEYINPUT115), .ZN(new_n819));
  NAND2_X1  g618(.A1(new_n810), .A2(KEYINPUT115), .ZN(new_n820));
  AND3_X1   g619(.A1(new_n819), .A2(new_n813), .A3(new_n820), .ZN(new_n821));
  NAND2_X1  g620(.A1(new_n821), .A2(new_n681), .ZN(new_n822));
  AOI21_X1  g621(.A(new_n565), .B1(new_n818), .B2(new_n822), .ZN(new_n823));
  NOR3_X1   g622(.A1(new_n722), .A2(new_n595), .A3(new_n617), .ZN(new_n824));
  NOR2_X1   g623(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  NAND2_X1  g624(.A1(new_n452), .A2(new_n377), .ZN(new_n826));
  NOR2_X1   g625(.A1(new_n825), .A2(new_n826), .ZN(new_n827));
  NAND2_X1  g626(.A1(new_n417), .A2(new_n338), .ZN(new_n828));
  INV_X1    g627(.A(new_n828), .ZN(new_n829));
  NAND2_X1  g628(.A1(new_n827), .A2(new_n829), .ZN(new_n830));
  XOR2_X1   g629(.A(new_n830), .B(KEYINPUT117), .Z(new_n831));
  INV_X1    g630(.A(G113gat), .ZN(new_n832));
  NAND3_X1  g631(.A1(new_n831), .A2(new_n832), .A3(new_n722), .ZN(new_n833));
  NAND2_X1  g632(.A1(new_n827), .A2(new_n342), .ZN(new_n834));
  OAI21_X1  g633(.A(G113gat), .B1(new_n834), .B2(new_n527), .ZN(new_n835));
  NAND2_X1  g634(.A1(new_n833), .A2(new_n835), .ZN(G1340gat));
  INV_X1    g635(.A(G120gat), .ZN(new_n837));
  NAND3_X1  g636(.A1(new_n831), .A2(new_n837), .A3(new_n617), .ZN(new_n838));
  OAI21_X1  g637(.A(G120gat), .B1(new_n834), .B2(new_n723), .ZN(new_n839));
  NAND2_X1  g638(.A1(new_n838), .A2(new_n839), .ZN(G1341gat));
  INV_X1    g639(.A(new_n565), .ZN(new_n841));
  NOR3_X1   g640(.A1(new_n834), .A2(new_n552), .A3(new_n841), .ZN(new_n842));
  NAND3_X1  g641(.A1(new_n827), .A2(new_n829), .A3(new_n565), .ZN(new_n843));
  AOI21_X1  g642(.A(new_n842), .B1(new_n552), .B2(new_n843), .ZN(G1342gat));
  NOR3_X1   g643(.A1(new_n830), .A2(G134gat), .A3(new_n594), .ZN(new_n845));
  INV_X1    g644(.A(new_n845), .ZN(new_n846));
  OR2_X1    g645(.A1(new_n846), .A2(KEYINPUT56), .ZN(new_n847));
  OAI21_X1  g646(.A(G134gat), .B1(new_n834), .B2(new_n594), .ZN(new_n848));
  NAND2_X1  g647(.A1(new_n846), .A2(KEYINPUT56), .ZN(new_n849));
  NAND3_X1  g648(.A1(new_n847), .A2(new_n848), .A3(new_n849), .ZN(G1343gat));
  INV_X1    g649(.A(KEYINPUT121), .ZN(new_n851));
  INV_X1    g650(.A(KEYINPUT58), .ZN(new_n852));
  NOR2_X1   g651(.A1(new_n641), .A2(new_n826), .ZN(new_n853));
  INV_X1    g652(.A(new_n824), .ZN(new_n854));
  NOR2_X1   g653(.A1(new_n527), .A2(new_n803), .ZN(new_n855));
  OAI21_X1  g654(.A(new_n594), .B1(new_n855), .B2(new_n811), .ZN(new_n856));
  AND2_X1   g655(.A1(new_n822), .A2(new_n856), .ZN(new_n857));
  OAI21_X1  g656(.A(new_n854), .B1(new_n857), .B2(new_n565), .ZN(new_n858));
  INV_X1    g657(.A(KEYINPUT57), .ZN(new_n859));
  NOR2_X1   g658(.A1(new_n338), .A2(new_n859), .ZN(new_n860));
  NAND2_X1  g659(.A1(new_n858), .A2(new_n860), .ZN(new_n861));
  AND4_X1   g660(.A1(new_n681), .A2(new_n819), .A3(new_n813), .A4(new_n820), .ZN(new_n862));
  NAND2_X1  g661(.A1(new_n814), .A2(new_n816), .ZN(new_n863));
  AOI21_X1  g662(.A(new_n681), .B1(new_n863), .B2(KEYINPUT116), .ZN(new_n864));
  AOI21_X1  g663(.A(new_n862), .B1(new_n864), .B2(new_n817), .ZN(new_n865));
  OAI21_X1  g664(.A(new_n854), .B1(new_n865), .B2(new_n565), .ZN(new_n866));
  AOI21_X1  g665(.A(KEYINPUT57), .B1(new_n866), .B2(new_n421), .ZN(new_n867));
  INV_X1    g666(.A(KEYINPUT118), .ZN(new_n868));
  OAI21_X1  g667(.A(new_n861), .B1(new_n867), .B2(new_n868), .ZN(new_n869));
  OAI21_X1  g668(.A(new_n421), .B1(new_n823), .B2(new_n824), .ZN(new_n870));
  NAND2_X1  g669(.A1(new_n870), .A2(new_n859), .ZN(new_n871));
  NOR2_X1   g670(.A1(new_n871), .A2(KEYINPUT118), .ZN(new_n872));
  OAI211_X1 g671(.A(new_n722), .B(new_n853), .C1(new_n869), .C2(new_n872), .ZN(new_n873));
  NAND2_X1  g672(.A1(new_n873), .A2(G141gat), .ZN(new_n874));
  NAND2_X1  g673(.A1(new_n640), .A2(new_n421), .ZN(new_n875));
  OAI21_X1  g674(.A(new_n452), .B1(new_n875), .B2(KEYINPUT119), .ZN(new_n876));
  AOI21_X1  g675(.A(new_n876), .B1(KEYINPUT119), .B2(new_n875), .ZN(new_n877));
  NAND2_X1  g676(.A1(new_n866), .A2(new_n877), .ZN(new_n878));
  INV_X1    g677(.A(new_n878), .ZN(new_n879));
  NOR3_X1   g678(.A1(new_n527), .A2(G141gat), .A3(new_n622), .ZN(new_n880));
  NAND2_X1  g679(.A1(new_n879), .A2(new_n880), .ZN(new_n881));
  AOI21_X1  g680(.A(new_n852), .B1(new_n874), .B2(new_n881), .ZN(new_n882));
  NAND2_X1  g681(.A1(new_n878), .A2(KEYINPUT120), .ZN(new_n883));
  NOR2_X1   g682(.A1(new_n527), .A2(G141gat), .ZN(new_n884));
  INV_X1    g683(.A(KEYINPUT120), .ZN(new_n885));
  NAND3_X1  g684(.A1(new_n866), .A2(new_n877), .A3(new_n885), .ZN(new_n886));
  NAND4_X1  g685(.A1(new_n883), .A2(new_n377), .A3(new_n884), .A4(new_n886), .ZN(new_n887));
  NAND2_X1  g686(.A1(new_n887), .A2(new_n852), .ZN(new_n888));
  INV_X1    g687(.A(new_n853), .ZN(new_n889));
  AOI22_X1  g688(.A1(new_n871), .A2(KEYINPUT118), .B1(new_n858), .B2(new_n860), .ZN(new_n890));
  NAND2_X1  g689(.A1(new_n867), .A2(new_n868), .ZN(new_n891));
  AOI21_X1  g690(.A(new_n889), .B1(new_n890), .B2(new_n891), .ZN(new_n892));
  NAND2_X1  g691(.A1(new_n892), .A2(new_n533), .ZN(new_n893));
  AOI21_X1  g692(.A(new_n888), .B1(new_n893), .B2(G141gat), .ZN(new_n894));
  OAI21_X1  g693(.A(new_n851), .B1(new_n882), .B2(new_n894), .ZN(new_n895));
  INV_X1    g694(.A(new_n888), .ZN(new_n896));
  AOI211_X1 g695(.A(new_n527), .B(new_n889), .C1(new_n890), .C2(new_n891), .ZN(new_n897));
  OAI21_X1  g696(.A(new_n896), .B1(new_n897), .B2(new_n301), .ZN(new_n898));
  AOI22_X1  g697(.A1(new_n873), .A2(G141gat), .B1(new_n879), .B2(new_n880), .ZN(new_n899));
  OAI211_X1 g698(.A(new_n898), .B(KEYINPUT121), .C1(new_n852), .C2(new_n899), .ZN(new_n900));
  NAND2_X1  g699(.A1(new_n895), .A2(new_n900), .ZN(G1344gat));
  AND3_X1   g700(.A1(new_n883), .A2(new_n377), .A3(new_n886), .ZN(new_n902));
  NAND3_X1  g701(.A1(new_n902), .A2(new_n302), .A3(new_n617), .ZN(new_n903));
  AOI211_X1 g702(.A(KEYINPUT59), .B(new_n302), .C1(new_n892), .C2(new_n617), .ZN(new_n904));
  INV_X1    g703(.A(KEYINPUT59), .ZN(new_n905));
  NAND2_X1  g704(.A1(new_n821), .A2(new_n593), .ZN(new_n906));
  AOI21_X1  g705(.A(new_n565), .B1(new_n906), .B2(new_n856), .ZN(new_n907));
  NOR3_X1   g706(.A1(new_n595), .A2(new_n533), .A3(new_n617), .ZN(new_n908));
  OAI21_X1  g707(.A(new_n421), .B1(new_n907), .B2(new_n908), .ZN(new_n909));
  NAND2_X1  g708(.A1(new_n909), .A2(new_n859), .ZN(new_n910));
  XNOR2_X1  g709(.A(new_n910), .B(KEYINPUT122), .ZN(new_n911));
  INV_X1    g710(.A(new_n870), .ZN(new_n912));
  NAND2_X1  g711(.A1(new_n912), .A2(KEYINPUT57), .ZN(new_n913));
  NAND2_X1  g712(.A1(new_n911), .A2(new_n913), .ZN(new_n914));
  NAND3_X1  g713(.A1(new_n914), .A2(new_n617), .A3(new_n853), .ZN(new_n915));
  AOI21_X1  g714(.A(new_n905), .B1(new_n915), .B2(G148gat), .ZN(new_n916));
  OAI21_X1  g715(.A(new_n903), .B1(new_n904), .B2(new_n916), .ZN(G1345gat));
  AOI21_X1  g716(.A(G155gat), .B1(new_n902), .B2(new_n565), .ZN(new_n918));
  NOR2_X1   g717(.A1(new_n841), .A2(new_n554), .ZN(new_n919));
  AOI21_X1  g718(.A(new_n918), .B1(new_n892), .B2(new_n919), .ZN(G1346gat));
  INV_X1    g719(.A(G162gat), .ZN(new_n921));
  NAND3_X1  g720(.A1(new_n902), .A2(new_n921), .A3(new_n593), .ZN(new_n922));
  AND2_X1   g721(.A1(new_n892), .A2(new_n681), .ZN(new_n923));
  OAI21_X1  g722(.A(new_n922), .B1(new_n923), .B2(new_n921), .ZN(G1347gat));
  NAND2_X1  g723(.A1(new_n622), .A2(new_n408), .ZN(new_n925));
  NOR2_X1   g724(.A1(new_n825), .A2(new_n925), .ZN(new_n926));
  NAND2_X1  g725(.A1(new_n926), .A2(new_n342), .ZN(new_n927));
  OAI21_X1  g726(.A(G169gat), .B1(new_n927), .B2(new_n527), .ZN(new_n928));
  NAND2_X1  g727(.A1(new_n926), .A2(new_n829), .ZN(new_n929));
  OR2_X1    g728(.A1(new_n695), .A2(G169gat), .ZN(new_n930));
  OAI21_X1  g729(.A(new_n928), .B1(new_n929), .B2(new_n930), .ZN(G1348gat));
  INV_X1    g730(.A(new_n929), .ZN(new_n932));
  AOI21_X1  g731(.A(G176gat), .B1(new_n932), .B2(new_n617), .ZN(new_n933));
  NAND4_X1  g732(.A1(new_n926), .A2(G176gat), .A3(new_n342), .A4(new_n617), .ZN(new_n934));
  INV_X1    g733(.A(KEYINPUT123), .ZN(new_n935));
  AND2_X1   g734(.A1(new_n934), .A2(new_n935), .ZN(new_n936));
  NOR2_X1   g735(.A1(new_n934), .A2(new_n935), .ZN(new_n937));
  NOR3_X1   g736(.A1(new_n933), .A2(new_n936), .A3(new_n937), .ZN(G1349gat));
  INV_X1    g737(.A(KEYINPUT124), .ZN(new_n939));
  OAI21_X1  g738(.A(new_n939), .B1(new_n927), .B2(new_n841), .ZN(new_n940));
  NAND4_X1  g739(.A1(new_n926), .A2(KEYINPUT124), .A3(new_n342), .A4(new_n565), .ZN(new_n941));
  NAND3_X1  g740(.A1(new_n940), .A2(G183gat), .A3(new_n941), .ZN(new_n942));
  INV_X1    g741(.A(KEYINPUT125), .ZN(new_n943));
  OAI21_X1  g742(.A(new_n565), .B1(new_n235), .B2(new_n232), .ZN(new_n944));
  OAI211_X1 g743(.A(new_n942), .B(new_n943), .C1(new_n929), .C2(new_n944), .ZN(new_n945));
  XNOR2_X1  g744(.A(new_n945), .B(KEYINPUT60), .ZN(G1350gat));
  NAND3_X1  g745(.A1(new_n932), .A2(new_n210), .A3(new_n681), .ZN(new_n947));
  OAI21_X1  g746(.A(G190gat), .B1(new_n927), .B2(new_n594), .ZN(new_n948));
  AND2_X1   g747(.A1(new_n948), .A2(KEYINPUT61), .ZN(new_n949));
  INV_X1    g748(.A(KEYINPUT126), .ZN(new_n950));
  NAND2_X1  g749(.A1(new_n949), .A2(new_n950), .ZN(new_n951));
  OAI21_X1  g750(.A(new_n951), .B1(KEYINPUT61), .B2(new_n948), .ZN(new_n952));
  NOR2_X1   g751(.A1(new_n949), .A2(new_n950), .ZN(new_n953));
  OAI21_X1  g752(.A(new_n947), .B1(new_n952), .B2(new_n953), .ZN(G1351gat));
  NOR2_X1   g753(.A1(new_n641), .A2(new_n925), .ZN(new_n955));
  INV_X1    g754(.A(new_n955), .ZN(new_n956));
  AOI21_X1  g755(.A(new_n956), .B1(new_n911), .B2(new_n913), .ZN(new_n957));
  AOI21_X1  g756(.A(new_n518), .B1(new_n957), .B2(new_n533), .ZN(new_n958));
  NAND2_X1  g757(.A1(new_n912), .A2(new_n955), .ZN(new_n959));
  NOR3_X1   g758(.A1(new_n959), .A2(G197gat), .A3(new_n695), .ZN(new_n960));
  OR2_X1    g759(.A1(new_n958), .A2(new_n960), .ZN(G1352gat));
  OR3_X1    g760(.A1(new_n959), .A2(G204gat), .A3(new_n723), .ZN(new_n962));
  NAND2_X1  g761(.A1(new_n962), .A2(KEYINPUT62), .ZN(new_n963));
  XNOR2_X1  g762(.A(new_n963), .B(KEYINPUT127), .ZN(new_n964));
  NAND3_X1  g763(.A1(new_n914), .A2(new_n617), .A3(new_n955), .ZN(new_n965));
  NAND2_X1  g764(.A1(new_n965), .A2(G204gat), .ZN(new_n966));
  OAI211_X1 g765(.A(new_n964), .B(new_n966), .C1(KEYINPUT62), .C2(new_n962), .ZN(G1353gat));
  INV_X1    g766(.A(new_n959), .ZN(new_n968));
  NAND3_X1  g767(.A1(new_n968), .A2(new_n288), .A3(new_n565), .ZN(new_n969));
  AOI21_X1  g768(.A(new_n288), .B1(new_n957), .B2(new_n565), .ZN(new_n970));
  AND2_X1   g769(.A1(new_n970), .A2(KEYINPUT63), .ZN(new_n971));
  NOR2_X1   g770(.A1(new_n970), .A2(KEYINPUT63), .ZN(new_n972));
  OAI21_X1  g771(.A(new_n969), .B1(new_n971), .B2(new_n972), .ZN(G1354gat));
  AOI21_X1  g772(.A(G218gat), .B1(new_n968), .B2(new_n681), .ZN(new_n974));
  NOR2_X1   g773(.A1(new_n594), .A2(new_n289), .ZN(new_n975));
  AOI21_X1  g774(.A(new_n974), .B1(new_n957), .B2(new_n975), .ZN(G1355gat));
endmodule


