//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 1 0 1 0 1 1 0 1 1 0 1 1 1 1 0 1 1 1 1 0 1 1 1 1 1 0 1 0 0 1 1 1 1 0 1 0 0 0 0 1 0 1 0 1 0 0 1 0 0 0 0 1 1 1 1 1 0 0 0 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:20:13 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n677, new_n678,
    new_n679, new_n680, new_n681, new_n682, new_n683, new_n684, new_n685,
    new_n686, new_n687, new_n688, new_n689, new_n691, new_n692, new_n693,
    new_n694, new_n695, new_n696, new_n697, new_n699, new_n700, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n748, new_n749, new_n750, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n772, new_n773, new_n774, new_n775,
    new_n776, new_n777, new_n778, new_n780, new_n781, new_n782, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n790, new_n791, new_n792,
    new_n793, new_n795, new_n797, new_n798, new_n799, new_n800, new_n801,
    new_n802, new_n803, new_n804, new_n805, new_n806, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n816, new_n817,
    new_n818, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n870, new_n871, new_n872, new_n874, new_n875, new_n876, new_n877,
    new_n878, new_n880, new_n881, new_n882, new_n883, new_n884, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n941, new_n942, new_n943, new_n944,
    new_n946, new_n947, new_n948, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n959, new_n960, new_n961,
    new_n962, new_n964, new_n965, new_n966, new_n967, new_n968, new_n970,
    new_n971, new_n972, new_n973, new_n975, new_n976, new_n977, new_n978,
    new_n979, new_n980, new_n981, new_n982, new_n983, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n994,
    new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1009, new_n1010;
  XNOR2_X1  g000(.A(G78gat), .B(G106gat), .ZN(new_n202));
  XNOR2_X1  g001(.A(KEYINPUT31), .B(G50gat), .ZN(new_n203));
  XOR2_X1   g002(.A(new_n202), .B(new_n203), .Z(new_n204));
  XOR2_X1   g003(.A(new_n204), .B(KEYINPUT81), .Z(new_n205));
  XNOR2_X1  g004(.A(G211gat), .B(G218gat), .ZN(new_n206));
  INV_X1    g005(.A(KEYINPUT73), .ZN(new_n207));
  NOR2_X1   g006(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  INV_X1    g007(.A(G197gat), .ZN(new_n209));
  INV_X1    g008(.A(G204gat), .ZN(new_n210));
  NAND2_X1  g009(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  NAND2_X1  g010(.A1(G197gat), .A2(G204gat), .ZN(new_n212));
  NAND2_X1  g011(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  NAND2_X1  g012(.A1(G211gat), .A2(G218gat), .ZN(new_n214));
  INV_X1    g013(.A(KEYINPUT22), .ZN(new_n215));
  NAND2_X1  g014(.A1(new_n214), .A2(new_n215), .ZN(new_n216));
  NAND2_X1  g015(.A1(new_n213), .A2(new_n216), .ZN(new_n217));
  NOR2_X1   g016(.A1(new_n208), .A2(new_n217), .ZN(new_n218));
  AOI22_X1  g017(.A1(new_n211), .A2(new_n212), .B1(new_n215), .B2(new_n214), .ZN(new_n219));
  NOR3_X1   g018(.A1(new_n219), .A2(new_n207), .A3(new_n206), .ZN(new_n220));
  NOR2_X1   g019(.A1(new_n218), .A2(new_n220), .ZN(new_n221));
  NAND2_X1  g020(.A1(G155gat), .A2(G162gat), .ZN(new_n222));
  NAND2_X1  g021(.A1(new_n222), .A2(KEYINPUT2), .ZN(new_n223));
  INV_X1    g022(.A(KEYINPUT76), .ZN(new_n224));
  NAND2_X1  g023(.A1(new_n223), .A2(new_n224), .ZN(new_n225));
  XNOR2_X1  g024(.A(G155gat), .B(G162gat), .ZN(new_n226));
  XNOR2_X1  g025(.A(G141gat), .B(G148gat), .ZN(new_n227));
  AND2_X1   g026(.A1(new_n222), .A2(KEYINPUT2), .ZN(new_n228));
  OAI211_X1 g027(.A(new_n225), .B(new_n226), .C1(new_n227), .C2(new_n228), .ZN(new_n229));
  INV_X1    g028(.A(G141gat), .ZN(new_n230));
  NAND2_X1  g029(.A1(new_n230), .A2(G148gat), .ZN(new_n231));
  INV_X1    g030(.A(G148gat), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n232), .A2(G141gat), .ZN(new_n233));
  NAND2_X1  g032(.A1(new_n231), .A2(new_n233), .ZN(new_n234));
  AND2_X1   g033(.A1(G155gat), .A2(G162gat), .ZN(new_n235));
  NOR2_X1   g034(.A1(G155gat), .A2(G162gat), .ZN(new_n236));
  NOR2_X1   g035(.A1(new_n235), .A2(new_n236), .ZN(new_n237));
  OAI211_X1 g036(.A(new_n223), .B(new_n234), .C1(new_n237), .C2(new_n224), .ZN(new_n238));
  AOI21_X1  g037(.A(KEYINPUT3), .B1(new_n229), .B2(new_n238), .ZN(new_n239));
  OAI21_X1  g038(.A(new_n221), .B1(new_n239), .B2(KEYINPUT29), .ZN(new_n240));
  AND3_X1   g039(.A1(new_n240), .A2(G228gat), .A3(G233gat), .ZN(new_n241));
  NAND2_X1  g040(.A1(new_n229), .A2(new_n238), .ZN(new_n242));
  INV_X1    g041(.A(new_n242), .ZN(new_n243));
  INV_X1    g042(.A(KEYINPUT3), .ZN(new_n244));
  NAND2_X1  g043(.A1(new_n208), .A2(new_n217), .ZN(new_n245));
  OAI21_X1  g044(.A(new_n219), .B1(new_n207), .B2(new_n206), .ZN(new_n246));
  AOI21_X1  g045(.A(KEYINPUT29), .B1(new_n245), .B2(new_n246), .ZN(new_n247));
  OAI21_X1  g046(.A(new_n244), .B1(new_n247), .B2(KEYINPUT82), .ZN(new_n248));
  INV_X1    g047(.A(KEYINPUT82), .ZN(new_n249));
  AOI211_X1 g048(.A(new_n249), .B(KEYINPUT29), .C1(new_n245), .C2(new_n246), .ZN(new_n250));
  OAI21_X1  g049(.A(new_n243), .B1(new_n248), .B2(new_n250), .ZN(new_n251));
  NAND2_X1  g050(.A1(G228gat), .A2(G233gat), .ZN(new_n252));
  INV_X1    g051(.A(KEYINPUT29), .ZN(new_n253));
  INV_X1    g052(.A(new_n206), .ZN(new_n254));
  OAI21_X1  g053(.A(new_n253), .B1(new_n254), .B2(new_n219), .ZN(new_n255));
  NOR2_X1   g054(.A1(new_n217), .A2(new_n206), .ZN(new_n256));
  OAI21_X1  g055(.A(new_n244), .B1(new_n255), .B2(new_n256), .ZN(new_n257));
  NAND2_X1  g056(.A1(new_n257), .A2(new_n243), .ZN(new_n258));
  NAND2_X1  g057(.A1(new_n240), .A2(new_n258), .ZN(new_n259));
  AOI22_X1  g058(.A1(new_n241), .A2(new_n251), .B1(new_n252), .B2(new_n259), .ZN(new_n260));
  XOR2_X1   g059(.A(KEYINPUT83), .B(G22gat), .Z(new_n261));
  OAI21_X1  g060(.A(KEYINPUT84), .B1(new_n260), .B2(new_n261), .ZN(new_n262));
  NAND2_X1  g061(.A1(new_n259), .A2(new_n252), .ZN(new_n263));
  OAI21_X1  g062(.A(new_n253), .B1(new_n218), .B2(new_n220), .ZN(new_n264));
  AOI21_X1  g063(.A(KEYINPUT3), .B1(new_n264), .B2(new_n249), .ZN(new_n265));
  INV_X1    g064(.A(new_n250), .ZN(new_n266));
  AOI21_X1  g065(.A(new_n242), .B1(new_n265), .B2(new_n266), .ZN(new_n267));
  NAND3_X1  g066(.A1(new_n240), .A2(G228gat), .A3(G233gat), .ZN(new_n268));
  OAI21_X1  g067(.A(new_n263), .B1(new_n267), .B2(new_n268), .ZN(new_n269));
  INV_X1    g068(.A(KEYINPUT84), .ZN(new_n270));
  INV_X1    g069(.A(new_n261), .ZN(new_n271));
  NAND3_X1  g070(.A1(new_n269), .A2(new_n270), .A3(new_n271), .ZN(new_n272));
  NAND2_X1  g071(.A1(new_n262), .A2(new_n272), .ZN(new_n273));
  NAND2_X1  g072(.A1(new_n260), .A2(new_n261), .ZN(new_n274));
  AOI21_X1  g073(.A(new_n205), .B1(new_n273), .B2(new_n274), .ZN(new_n275));
  INV_X1    g074(.A(new_n204), .ZN(new_n276));
  NAND2_X1  g075(.A1(new_n274), .A2(new_n276), .ZN(new_n277));
  OR2_X1    g076(.A1(new_n269), .A2(KEYINPUT85), .ZN(new_n278));
  INV_X1    g077(.A(G22gat), .ZN(new_n279));
  AOI21_X1  g078(.A(new_n279), .B1(new_n269), .B2(KEYINPUT85), .ZN(new_n280));
  AOI21_X1  g079(.A(new_n277), .B1(new_n278), .B2(new_n280), .ZN(new_n281));
  OR2_X1    g080(.A1(new_n275), .A2(new_n281), .ZN(new_n282));
  NOR2_X1   g081(.A1(G169gat), .A2(G176gat), .ZN(new_n283));
  NAND2_X1  g082(.A1(new_n283), .A2(KEYINPUT23), .ZN(new_n284));
  NAND2_X1  g083(.A1(G169gat), .A2(G176gat), .ZN(new_n285));
  INV_X1    g084(.A(KEYINPUT23), .ZN(new_n286));
  OAI21_X1  g085(.A(new_n286), .B1(G169gat), .B2(G176gat), .ZN(new_n287));
  AND4_X1   g086(.A1(KEYINPUT25), .A2(new_n284), .A3(new_n285), .A4(new_n287), .ZN(new_n288));
  NAND2_X1  g087(.A1(G183gat), .A2(G190gat), .ZN(new_n289));
  INV_X1    g088(.A(KEYINPUT65), .ZN(new_n290));
  NAND2_X1  g089(.A1(new_n289), .A2(new_n290), .ZN(new_n291));
  INV_X1    g090(.A(KEYINPUT24), .ZN(new_n292));
  NAND3_X1  g091(.A1(KEYINPUT65), .A2(G183gat), .A3(G190gat), .ZN(new_n293));
  NAND3_X1  g092(.A1(new_n291), .A2(new_n292), .A3(new_n293), .ZN(new_n294));
  OAI21_X1  g093(.A(KEYINPUT66), .B1(G183gat), .B2(G190gat), .ZN(new_n295));
  NAND3_X1  g094(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n296));
  NAND2_X1  g095(.A1(new_n295), .A2(new_n296), .ZN(new_n297));
  AND2_X1   g096(.A1(KEYINPUT24), .A2(G183gat), .ZN(new_n298));
  NAND3_X1  g097(.A1(new_n298), .A2(KEYINPUT66), .A3(G190gat), .ZN(new_n299));
  NAND3_X1  g098(.A1(new_n294), .A2(new_n297), .A3(new_n299), .ZN(new_n300));
  NAND2_X1  g099(.A1(new_n288), .A2(new_n300), .ZN(new_n301));
  INV_X1    g100(.A(KEYINPUT25), .ZN(new_n302));
  NAND3_X1  g101(.A1(new_n284), .A2(new_n285), .A3(new_n287), .ZN(new_n303));
  OAI21_X1  g102(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n304));
  AOI22_X1  g103(.A1(new_n289), .A2(new_n304), .B1(new_n298), .B2(G190gat), .ZN(new_n305));
  OAI21_X1  g104(.A(new_n302), .B1(new_n303), .B2(new_n305), .ZN(new_n306));
  NAND2_X1  g105(.A1(new_n301), .A2(new_n306), .ZN(new_n307));
  INV_X1    g106(.A(KEYINPUT68), .ZN(new_n308));
  INV_X1    g107(.A(KEYINPUT67), .ZN(new_n309));
  INV_X1    g108(.A(KEYINPUT27), .ZN(new_n310));
  NOR2_X1   g109(.A1(new_n310), .A2(G183gat), .ZN(new_n311));
  INV_X1    g110(.A(G183gat), .ZN(new_n312));
  NOR2_X1   g111(.A1(new_n312), .A2(KEYINPUT27), .ZN(new_n313));
  OAI21_X1  g112(.A(new_n309), .B1(new_n311), .B2(new_n313), .ZN(new_n314));
  NAND2_X1  g113(.A1(new_n312), .A2(KEYINPUT27), .ZN(new_n315));
  NAND2_X1  g114(.A1(new_n310), .A2(G183gat), .ZN(new_n316));
  NAND3_X1  g115(.A1(new_n315), .A2(new_n316), .A3(KEYINPUT67), .ZN(new_n317));
  INV_X1    g116(.A(KEYINPUT28), .ZN(new_n318));
  NOR2_X1   g117(.A1(new_n318), .A2(G190gat), .ZN(new_n319));
  NAND3_X1  g118(.A1(new_n314), .A2(new_n317), .A3(new_n319), .ZN(new_n320));
  INV_X1    g119(.A(G190gat), .ZN(new_n321));
  NAND3_X1  g120(.A1(new_n315), .A2(new_n316), .A3(new_n321), .ZN(new_n322));
  NAND2_X1  g121(.A1(new_n322), .A2(new_n318), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n320), .A2(new_n323), .ZN(new_n324));
  NAND2_X1  g123(.A1(new_n283), .A2(KEYINPUT26), .ZN(new_n325));
  INV_X1    g124(.A(KEYINPUT26), .ZN(new_n326));
  NAND2_X1  g125(.A1(new_n285), .A2(new_n326), .ZN(new_n327));
  OAI211_X1 g126(.A(new_n325), .B(new_n289), .C1(new_n327), .C2(new_n283), .ZN(new_n328));
  INV_X1    g127(.A(new_n328), .ZN(new_n329));
  AOI21_X1  g128(.A(new_n308), .B1(new_n324), .B2(new_n329), .ZN(new_n330));
  AOI211_X1 g129(.A(KEYINPUT68), .B(new_n328), .C1(new_n320), .C2(new_n323), .ZN(new_n331));
  OAI21_X1  g130(.A(new_n307), .B1(new_n330), .B2(new_n331), .ZN(new_n332));
  INV_X1    g131(.A(G120gat), .ZN(new_n333));
  NAND2_X1  g132(.A1(new_n333), .A2(G113gat), .ZN(new_n334));
  INV_X1    g133(.A(G113gat), .ZN(new_n335));
  NAND2_X1  g134(.A1(new_n335), .A2(G120gat), .ZN(new_n336));
  NAND2_X1  g135(.A1(new_n334), .A2(new_n336), .ZN(new_n337));
  XNOR2_X1  g136(.A(G127gat), .B(G134gat), .ZN(new_n338));
  INV_X1    g137(.A(KEYINPUT1), .ZN(new_n339));
  NAND3_X1  g138(.A1(new_n337), .A2(new_n338), .A3(new_n339), .ZN(new_n340));
  INV_X1    g139(.A(new_n340), .ZN(new_n341));
  NOR2_X1   g140(.A1(G127gat), .A2(G134gat), .ZN(new_n342));
  INV_X1    g141(.A(new_n342), .ZN(new_n343));
  XNOR2_X1  g142(.A(G113gat), .B(G120gat), .ZN(new_n344));
  OAI21_X1  g143(.A(new_n343), .B1(new_n344), .B2(KEYINPUT1), .ZN(new_n345));
  INV_X1    g144(.A(G127gat), .ZN(new_n346));
  INV_X1    g145(.A(G134gat), .ZN(new_n347));
  NAND2_X1  g146(.A1(new_n347), .A2(KEYINPUT69), .ZN(new_n348));
  INV_X1    g147(.A(KEYINPUT69), .ZN(new_n349));
  NAND2_X1  g148(.A1(new_n349), .A2(G134gat), .ZN(new_n350));
  AOI21_X1  g149(.A(new_n346), .B1(new_n348), .B2(new_n350), .ZN(new_n351));
  OAI21_X1  g150(.A(KEYINPUT70), .B1(new_n345), .B2(new_n351), .ZN(new_n352));
  AOI21_X1  g151(.A(new_n342), .B1(new_n337), .B2(new_n339), .ZN(new_n353));
  INV_X1    g152(.A(new_n351), .ZN(new_n354));
  INV_X1    g153(.A(KEYINPUT70), .ZN(new_n355));
  NAND3_X1  g154(.A1(new_n353), .A2(new_n354), .A3(new_n355), .ZN(new_n356));
  AOI21_X1  g155(.A(new_n341), .B1(new_n352), .B2(new_n356), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n332), .A2(new_n357), .ZN(new_n358));
  NOR3_X1   g157(.A1(new_n345), .A2(KEYINPUT70), .A3(new_n351), .ZN(new_n359));
  AOI21_X1  g158(.A(new_n355), .B1(new_n353), .B2(new_n354), .ZN(new_n360));
  OAI21_X1  g159(.A(new_n340), .B1(new_n359), .B2(new_n360), .ZN(new_n361));
  OAI211_X1 g160(.A(new_n361), .B(new_n307), .C1(new_n330), .C2(new_n331), .ZN(new_n362));
  NAND2_X1  g161(.A1(G227gat), .A2(G233gat), .ZN(new_n363));
  XNOR2_X1  g162(.A(new_n363), .B(KEYINPUT64), .ZN(new_n364));
  NAND3_X1  g163(.A1(new_n358), .A2(new_n362), .A3(new_n364), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n365), .A2(KEYINPUT32), .ZN(new_n366));
  INV_X1    g165(.A(KEYINPUT33), .ZN(new_n367));
  NAND2_X1  g166(.A1(new_n365), .A2(new_n367), .ZN(new_n368));
  XOR2_X1   g167(.A(G15gat), .B(G43gat), .Z(new_n369));
  XNOR2_X1  g168(.A(G71gat), .B(G99gat), .ZN(new_n370));
  XNOR2_X1  g169(.A(new_n369), .B(new_n370), .ZN(new_n371));
  NAND3_X1  g170(.A1(new_n366), .A2(new_n368), .A3(new_n371), .ZN(new_n372));
  INV_X1    g171(.A(new_n371), .ZN(new_n373));
  OAI211_X1 g172(.A(new_n365), .B(KEYINPUT32), .C1(new_n367), .C2(new_n373), .ZN(new_n374));
  NAND2_X1  g173(.A1(new_n372), .A2(new_n374), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n358), .A2(new_n362), .ZN(new_n376));
  NAND2_X1  g175(.A1(new_n376), .A2(new_n363), .ZN(new_n377));
  NOR2_X1   g176(.A1(new_n364), .A2(KEYINPUT34), .ZN(new_n378));
  AOI22_X1  g177(.A1(new_n377), .A2(KEYINPUT34), .B1(new_n376), .B2(new_n378), .ZN(new_n379));
  INV_X1    g178(.A(new_n379), .ZN(new_n380));
  NAND2_X1  g179(.A1(new_n375), .A2(new_n380), .ZN(new_n381));
  INV_X1    g180(.A(KEYINPUT71), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n381), .A2(new_n382), .ZN(new_n383));
  AOI21_X1  g182(.A(new_n379), .B1(new_n372), .B2(new_n374), .ZN(new_n384));
  NAND2_X1  g183(.A1(new_n384), .A2(KEYINPUT71), .ZN(new_n385));
  NAND3_X1  g184(.A1(new_n372), .A2(new_n379), .A3(new_n374), .ZN(new_n386));
  NAND4_X1  g185(.A1(new_n282), .A2(new_n383), .A3(new_n385), .A4(new_n386), .ZN(new_n387));
  XNOR2_X1  g186(.A(G8gat), .B(G36gat), .ZN(new_n388));
  XNOR2_X1  g187(.A(G64gat), .B(G92gat), .ZN(new_n389));
  XOR2_X1   g188(.A(new_n388), .B(new_n389), .Z(new_n390));
  NAND2_X1  g189(.A1(G226gat), .A2(G233gat), .ZN(new_n391));
  INV_X1    g190(.A(new_n391), .ZN(new_n392));
  AOI21_X1  g191(.A(new_n392), .B1(new_n332), .B2(new_n253), .ZN(new_n393));
  INV_X1    g192(.A(KEYINPUT74), .ZN(new_n394));
  AOI22_X1  g193(.A1(new_n324), .A2(new_n329), .B1(new_n301), .B2(new_n306), .ZN(new_n395));
  OAI21_X1  g194(.A(new_n394), .B1(new_n395), .B2(new_n391), .ZN(new_n396));
  NAND2_X1  g195(.A1(new_n304), .A2(new_n289), .ZN(new_n397));
  NAND2_X1  g196(.A1(new_n397), .A2(new_n296), .ZN(new_n398));
  NAND4_X1  g197(.A1(new_n398), .A2(new_n284), .A3(new_n285), .A4(new_n287), .ZN(new_n399));
  AOI22_X1  g198(.A1(new_n399), .A2(new_n302), .B1(new_n288), .B2(new_n300), .ZN(new_n400));
  AOI21_X1  g199(.A(new_n328), .B1(new_n320), .B2(new_n323), .ZN(new_n401));
  OAI211_X1 g200(.A(KEYINPUT74), .B(new_n392), .C1(new_n400), .C2(new_n401), .ZN(new_n402));
  NAND2_X1  g201(.A1(new_n396), .A2(new_n402), .ZN(new_n403));
  OAI21_X1  g202(.A(new_n221), .B1(new_n393), .B2(new_n403), .ZN(new_n404));
  NAND2_X1  g203(.A1(new_n332), .A2(new_n392), .ZN(new_n405));
  NAND2_X1  g204(.A1(new_n324), .A2(new_n329), .ZN(new_n406));
  AOI21_X1  g205(.A(KEYINPUT29), .B1(new_n406), .B2(new_n307), .ZN(new_n407));
  OAI21_X1  g206(.A(KEYINPUT75), .B1(new_n407), .B2(new_n392), .ZN(new_n408));
  INV_X1    g207(.A(new_n221), .ZN(new_n409));
  INV_X1    g208(.A(KEYINPUT75), .ZN(new_n410));
  OAI211_X1 g209(.A(new_n410), .B(new_n391), .C1(new_n395), .C2(KEYINPUT29), .ZN(new_n411));
  NAND4_X1  g210(.A1(new_n405), .A2(new_n408), .A3(new_n409), .A4(new_n411), .ZN(new_n412));
  AOI21_X1  g211(.A(new_n390), .B1(new_n404), .B2(new_n412), .ZN(new_n413));
  INV_X1    g212(.A(KEYINPUT30), .ZN(new_n414));
  NOR2_X1   g213(.A1(new_n413), .A2(new_n414), .ZN(new_n415));
  AND3_X1   g214(.A1(new_n404), .A2(new_n390), .A3(new_n412), .ZN(new_n416));
  INV_X1    g215(.A(new_n416), .ZN(new_n417));
  NAND2_X1  g216(.A1(new_n415), .A2(new_n417), .ZN(new_n418));
  AND4_X1   g217(.A1(new_n414), .A2(new_n404), .A3(new_n390), .A4(new_n412), .ZN(new_n419));
  INV_X1    g218(.A(new_n419), .ZN(new_n420));
  NAND2_X1  g219(.A1(new_n418), .A2(new_n420), .ZN(new_n421));
  NAND2_X1  g220(.A1(G225gat), .A2(G233gat), .ZN(new_n422));
  XOR2_X1   g221(.A(new_n422), .B(KEYINPUT77), .Z(new_n423));
  INV_X1    g222(.A(new_n423), .ZN(new_n424));
  NAND2_X1  g223(.A1(new_n361), .A2(new_n243), .ZN(new_n425));
  OAI211_X1 g224(.A(new_n340), .B(new_n242), .C1(new_n359), .C2(new_n360), .ZN(new_n426));
  AOI21_X1  g225(.A(new_n424), .B1(new_n425), .B2(new_n426), .ZN(new_n427));
  INV_X1    g226(.A(KEYINPUT5), .ZN(new_n428));
  OAI21_X1  g227(.A(KEYINPUT78), .B1(new_n427), .B2(new_n428), .ZN(new_n429));
  NAND2_X1  g228(.A1(new_n242), .A2(new_n244), .ZN(new_n430));
  NAND3_X1  g229(.A1(new_n229), .A2(new_n238), .A3(KEYINPUT3), .ZN(new_n431));
  NAND2_X1  g230(.A1(new_n430), .A2(new_n431), .ZN(new_n432));
  OAI211_X1 g231(.A(new_n426), .B(KEYINPUT4), .C1(new_n432), .C2(new_n357), .ZN(new_n433));
  INV_X1    g232(.A(KEYINPUT4), .ZN(new_n434));
  NAND3_X1  g233(.A1(new_n357), .A2(new_n434), .A3(new_n242), .ZN(new_n435));
  NAND2_X1  g234(.A1(new_n433), .A2(new_n435), .ZN(new_n436));
  NAND2_X1  g235(.A1(new_n436), .A2(new_n424), .ZN(new_n437));
  INV_X1    g236(.A(new_n426), .ZN(new_n438));
  NAND2_X1  g237(.A1(new_n352), .A2(new_n356), .ZN(new_n439));
  AOI21_X1  g238(.A(new_n242), .B1(new_n439), .B2(new_n340), .ZN(new_n440));
  OAI21_X1  g239(.A(new_n423), .B1(new_n438), .B2(new_n440), .ZN(new_n441));
  INV_X1    g240(.A(KEYINPUT78), .ZN(new_n442));
  NAND3_X1  g241(.A1(new_n441), .A2(new_n442), .A3(KEYINPUT5), .ZN(new_n443));
  NAND3_X1  g242(.A1(new_n429), .A2(new_n437), .A3(new_n443), .ZN(new_n444));
  NAND3_X1  g243(.A1(new_n436), .A2(new_n428), .A3(new_n424), .ZN(new_n445));
  NAND2_X1  g244(.A1(new_n444), .A2(new_n445), .ZN(new_n446));
  XOR2_X1   g245(.A(KEYINPUT79), .B(KEYINPUT0), .Z(new_n447));
  XNOR2_X1  g246(.A(new_n447), .B(KEYINPUT80), .ZN(new_n448));
  XNOR2_X1  g247(.A(G1gat), .B(G29gat), .ZN(new_n449));
  XNOR2_X1  g248(.A(new_n448), .B(new_n449), .ZN(new_n450));
  XNOR2_X1  g249(.A(G57gat), .B(G85gat), .ZN(new_n451));
  XOR2_X1   g250(.A(new_n450), .B(new_n451), .Z(new_n452));
  NAND2_X1  g251(.A1(new_n452), .A2(KEYINPUT6), .ZN(new_n453));
  INV_X1    g252(.A(new_n452), .ZN(new_n454));
  INV_X1    g253(.A(KEYINPUT6), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n454), .A2(new_n455), .ZN(new_n456));
  NAND3_X1  g255(.A1(new_n446), .A2(new_n453), .A3(new_n456), .ZN(new_n457));
  NAND4_X1  g256(.A1(new_n444), .A2(new_n455), .A3(new_n445), .A4(new_n454), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n421), .A2(new_n459), .ZN(new_n460));
  OAI21_X1  g259(.A(KEYINPUT35), .B1(new_n387), .B2(new_n460), .ZN(new_n461));
  INV_X1    g260(.A(new_n386), .ZN(new_n462));
  NOR2_X1   g261(.A1(new_n462), .A2(new_n384), .ZN(new_n463));
  NAND2_X1  g262(.A1(new_n282), .A2(new_n463), .ZN(new_n464));
  INV_X1    g263(.A(KEYINPUT35), .ZN(new_n465));
  NAND3_X1  g264(.A1(new_n421), .A2(new_n465), .A3(new_n459), .ZN(new_n466));
  OR2_X1    g265(.A1(new_n464), .A2(new_n466), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n461), .A2(new_n467), .ZN(new_n468));
  AND3_X1   g267(.A1(new_n457), .A2(new_n458), .A3(new_n417), .ZN(new_n469));
  INV_X1    g268(.A(new_n390), .ZN(new_n470));
  INV_X1    g269(.A(KEYINPUT37), .ZN(new_n471));
  NAND2_X1  g270(.A1(new_n412), .A2(new_n471), .ZN(new_n472));
  NAND2_X1  g271(.A1(new_n406), .A2(KEYINPUT68), .ZN(new_n473));
  NAND2_X1  g272(.A1(new_n401), .A2(new_n308), .ZN(new_n474));
  AOI21_X1  g273(.A(new_n400), .B1(new_n473), .B2(new_n474), .ZN(new_n475));
  OAI21_X1  g274(.A(new_n391), .B1(new_n475), .B2(KEYINPUT29), .ZN(new_n476));
  NAND2_X1  g275(.A1(new_n406), .A2(new_n307), .ZN(new_n477));
  AOI21_X1  g276(.A(KEYINPUT74), .B1(new_n477), .B2(new_n392), .ZN(new_n478));
  INV_X1    g277(.A(new_n402), .ZN(new_n479));
  NOR2_X1   g278(.A1(new_n478), .A2(new_n479), .ZN(new_n480));
  AOI21_X1  g279(.A(new_n409), .B1(new_n476), .B2(new_n480), .ZN(new_n481));
  OAI21_X1  g280(.A(new_n470), .B1(new_n472), .B2(new_n481), .ZN(new_n482));
  NOR2_X1   g281(.A1(new_n482), .A2(KEYINPUT38), .ZN(new_n483));
  OAI21_X1  g282(.A(new_n409), .B1(new_n393), .B2(new_n403), .ZN(new_n484));
  NAND4_X1  g283(.A1(new_n405), .A2(new_n408), .A3(new_n221), .A4(new_n411), .ZN(new_n485));
  NAND3_X1  g284(.A1(new_n484), .A2(KEYINPUT37), .A3(new_n485), .ZN(new_n486));
  INV_X1    g285(.A(KEYINPUT87), .ZN(new_n487));
  OR2_X1    g286(.A1(new_n486), .A2(new_n487), .ZN(new_n488));
  NAND2_X1  g287(.A1(new_n486), .A2(new_n487), .ZN(new_n489));
  NAND3_X1  g288(.A1(new_n483), .A2(new_n488), .A3(new_n489), .ZN(new_n490));
  AOI21_X1  g289(.A(new_n471), .B1(new_n404), .B2(new_n412), .ZN(new_n491));
  OAI21_X1  g290(.A(KEYINPUT38), .B1(new_n482), .B2(new_n491), .ZN(new_n492));
  INV_X1    g291(.A(KEYINPUT88), .ZN(new_n493));
  NAND2_X1  g292(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  OAI211_X1 g293(.A(KEYINPUT88), .B(KEYINPUT38), .C1(new_n482), .C2(new_n491), .ZN(new_n495));
  NAND4_X1  g294(.A1(new_n469), .A2(new_n490), .A3(new_n494), .A4(new_n495), .ZN(new_n496));
  INV_X1    g295(.A(KEYINPUT89), .ZN(new_n497));
  NAND2_X1  g296(.A1(new_n273), .A2(new_n274), .ZN(new_n498));
  INV_X1    g297(.A(new_n205), .ZN(new_n499));
  NAND2_X1  g298(.A1(new_n278), .A2(new_n280), .ZN(new_n500));
  INV_X1    g299(.A(new_n277), .ZN(new_n501));
  AOI22_X1  g300(.A1(new_n498), .A2(new_n499), .B1(new_n500), .B2(new_n501), .ZN(new_n502));
  NOR3_X1   g301(.A1(new_n416), .A2(new_n413), .A3(new_n414), .ZN(new_n503));
  NOR2_X1   g302(.A1(new_n503), .A2(new_n419), .ZN(new_n504));
  XOR2_X1   g303(.A(KEYINPUT86), .B(KEYINPUT39), .Z(new_n505));
  NAND4_X1  g304(.A1(new_n433), .A2(new_n423), .A3(new_n435), .A4(new_n505), .ZN(new_n506));
  AND2_X1   g305(.A1(new_n452), .A2(new_n506), .ZN(new_n507));
  INV_X1    g306(.A(KEYINPUT40), .ZN(new_n508));
  NOR2_X1   g307(.A1(new_n436), .A2(new_n424), .ZN(new_n509));
  NAND3_X1  g308(.A1(new_n425), .A2(new_n424), .A3(new_n426), .ZN(new_n510));
  NAND2_X1  g309(.A1(new_n510), .A2(KEYINPUT39), .ZN(new_n511));
  OAI211_X1 g310(.A(new_n507), .B(new_n508), .C1(new_n509), .C2(new_n511), .ZN(new_n512));
  NOR2_X1   g311(.A1(new_n509), .A2(new_n511), .ZN(new_n513));
  NAND2_X1  g312(.A1(new_n452), .A2(new_n506), .ZN(new_n514));
  OAI21_X1  g313(.A(KEYINPUT40), .B1(new_n513), .B2(new_n514), .ZN(new_n515));
  AOI22_X1  g314(.A1(new_n512), .A2(new_n515), .B1(new_n446), .B2(new_n454), .ZN(new_n516));
  AOI21_X1  g315(.A(new_n502), .B1(new_n504), .B2(new_n516), .ZN(new_n517));
  AND3_X1   g316(.A1(new_n496), .A2(new_n497), .A3(new_n517), .ZN(new_n518));
  AOI21_X1  g317(.A(new_n497), .B1(new_n496), .B2(new_n517), .ZN(new_n519));
  NOR2_X1   g318(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  NAND2_X1  g319(.A1(new_n460), .A2(new_n502), .ZN(new_n521));
  AND2_X1   g320(.A1(new_n386), .A2(KEYINPUT36), .ZN(new_n522));
  INV_X1    g321(.A(KEYINPUT72), .ZN(new_n523));
  NAND4_X1  g322(.A1(new_n383), .A2(new_n522), .A3(new_n523), .A4(new_n385), .ZN(new_n524));
  OAI21_X1  g323(.A(new_n524), .B1(KEYINPUT36), .B2(new_n463), .ZN(new_n525));
  AND3_X1   g324(.A1(new_n375), .A2(KEYINPUT71), .A3(new_n380), .ZN(new_n526));
  AOI21_X1  g325(.A(KEYINPUT71), .B1(new_n375), .B2(new_n380), .ZN(new_n527));
  NOR2_X1   g326(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  AOI21_X1  g327(.A(new_n523), .B1(new_n528), .B2(new_n522), .ZN(new_n529));
  OAI21_X1  g328(.A(new_n521), .B1(new_n525), .B2(new_n529), .ZN(new_n530));
  OAI21_X1  g329(.A(new_n468), .B1(new_n520), .B2(new_n530), .ZN(new_n531));
  XNOR2_X1  g330(.A(G113gat), .B(G141gat), .ZN(new_n532));
  XNOR2_X1  g331(.A(new_n532), .B(G197gat), .ZN(new_n533));
  XOR2_X1   g332(.A(KEYINPUT11), .B(G169gat), .Z(new_n534));
  XNOR2_X1  g333(.A(new_n533), .B(new_n534), .ZN(new_n535));
  XOR2_X1   g334(.A(new_n535), .B(KEYINPUT12), .Z(new_n536));
  XNOR2_X1  g335(.A(G15gat), .B(G22gat), .ZN(new_n537));
  XNOR2_X1  g336(.A(new_n537), .B(KEYINPUT90), .ZN(new_n538));
  INV_X1    g337(.A(KEYINPUT16), .ZN(new_n539));
  OAI21_X1  g338(.A(new_n538), .B1(new_n539), .B2(G1gat), .ZN(new_n540));
  OR2_X1    g339(.A1(new_n537), .A2(KEYINPUT90), .ZN(new_n541));
  INV_X1    g340(.A(G1gat), .ZN(new_n542));
  NAND2_X1  g341(.A1(new_n537), .A2(KEYINPUT90), .ZN(new_n543));
  NAND3_X1  g342(.A1(new_n541), .A2(new_n542), .A3(new_n543), .ZN(new_n544));
  INV_X1    g343(.A(G8gat), .ZN(new_n545));
  OAI211_X1 g344(.A(new_n540), .B(new_n544), .C1(KEYINPUT91), .C2(new_n545), .ZN(new_n546));
  NAND2_X1  g345(.A1(new_n540), .A2(new_n544), .ZN(new_n547));
  AOI21_X1  g346(.A(new_n545), .B1(new_n544), .B2(KEYINPUT91), .ZN(new_n548));
  NAND2_X1  g347(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  INV_X1    g348(.A(G36gat), .ZN(new_n550));
  AND2_X1   g349(.A1(KEYINPUT14), .A2(G29gat), .ZN(new_n551));
  NOR2_X1   g350(.A1(KEYINPUT14), .A2(G29gat), .ZN(new_n552));
  OAI21_X1  g351(.A(new_n550), .B1(new_n551), .B2(new_n552), .ZN(new_n553));
  INV_X1    g352(.A(G29gat), .ZN(new_n554));
  NAND3_X1  g353(.A1(new_n554), .A2(KEYINPUT14), .A3(G36gat), .ZN(new_n555));
  NAND2_X1  g354(.A1(new_n553), .A2(new_n555), .ZN(new_n556));
  OR2_X1    g355(.A1(new_n556), .A2(KEYINPUT15), .ZN(new_n557));
  NAND2_X1  g356(.A1(new_n556), .A2(KEYINPUT15), .ZN(new_n558));
  XNOR2_X1  g357(.A(G43gat), .B(G50gat), .ZN(new_n559));
  NAND3_X1  g358(.A1(new_n557), .A2(new_n558), .A3(new_n559), .ZN(new_n560));
  OR2_X1    g359(.A1(new_n558), .A2(new_n559), .ZN(new_n561));
  NAND2_X1  g360(.A1(new_n560), .A2(new_n561), .ZN(new_n562));
  NOR2_X1   g361(.A1(new_n562), .A2(KEYINPUT17), .ZN(new_n563));
  INV_X1    g362(.A(KEYINPUT17), .ZN(new_n564));
  AOI21_X1  g363(.A(new_n564), .B1(new_n560), .B2(new_n561), .ZN(new_n565));
  OAI211_X1 g364(.A(new_n546), .B(new_n549), .C1(new_n563), .C2(new_n565), .ZN(new_n566));
  NAND2_X1  g365(.A1(new_n549), .A2(new_n546), .ZN(new_n567));
  NAND2_X1  g366(.A1(new_n567), .A2(new_n562), .ZN(new_n568));
  NAND2_X1  g367(.A1(G229gat), .A2(G233gat), .ZN(new_n569));
  XOR2_X1   g368(.A(new_n569), .B(KEYINPUT92), .Z(new_n570));
  INV_X1    g369(.A(new_n570), .ZN(new_n571));
  NAND4_X1  g370(.A1(new_n566), .A2(new_n568), .A3(KEYINPUT18), .A4(new_n571), .ZN(new_n572));
  XNOR2_X1  g371(.A(new_n572), .B(KEYINPUT93), .ZN(new_n573));
  AND2_X1   g372(.A1(new_n549), .A2(new_n546), .ZN(new_n574));
  INV_X1    g373(.A(KEYINPUT94), .ZN(new_n575));
  NAND4_X1  g374(.A1(new_n574), .A2(new_n575), .A3(new_n560), .A4(new_n561), .ZN(new_n576));
  OAI21_X1  g375(.A(KEYINPUT94), .B1(new_n567), .B2(new_n562), .ZN(new_n577));
  NAND3_X1  g376(.A1(new_n576), .A2(new_n568), .A3(new_n577), .ZN(new_n578));
  XNOR2_X1  g377(.A(new_n570), .B(KEYINPUT13), .ZN(new_n579));
  NAND2_X1  g378(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  NAND3_X1  g379(.A1(new_n566), .A2(new_n571), .A3(new_n568), .ZN(new_n581));
  INV_X1    g380(.A(KEYINPUT18), .ZN(new_n582));
  NAND2_X1  g381(.A1(new_n581), .A2(new_n582), .ZN(new_n583));
  NAND2_X1  g382(.A1(new_n580), .A2(new_n583), .ZN(new_n584));
  OAI21_X1  g383(.A(new_n536), .B1(new_n573), .B2(new_n584), .ZN(new_n585));
  INV_X1    g384(.A(KEYINPUT93), .ZN(new_n586));
  XNOR2_X1  g385(.A(new_n572), .B(new_n586), .ZN(new_n587));
  INV_X1    g386(.A(new_n536), .ZN(new_n588));
  AOI22_X1  g387(.A1(new_n578), .A2(new_n579), .B1(new_n581), .B2(new_n582), .ZN(new_n589));
  NAND3_X1  g388(.A1(new_n587), .A2(new_n588), .A3(new_n589), .ZN(new_n590));
  NAND3_X1  g389(.A1(new_n585), .A2(KEYINPUT95), .A3(new_n590), .ZN(new_n591));
  INV_X1    g390(.A(KEYINPUT95), .ZN(new_n592));
  OAI211_X1 g391(.A(new_n592), .B(new_n536), .C1(new_n573), .C2(new_n584), .ZN(new_n593));
  NAND2_X1  g392(.A1(new_n591), .A2(new_n593), .ZN(new_n594));
  INV_X1    g393(.A(new_n594), .ZN(new_n595));
  XNOR2_X1  g394(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n596));
  INV_X1    g395(.A(G155gat), .ZN(new_n597));
  XNOR2_X1  g396(.A(new_n596), .B(new_n597), .ZN(new_n598));
  XNOR2_X1  g397(.A(G183gat), .B(G211gat), .ZN(new_n599));
  XOR2_X1   g398(.A(new_n598), .B(new_n599), .Z(new_n600));
  INV_X1    g399(.A(new_n600), .ZN(new_n601));
  XOR2_X1   g400(.A(G57gat), .B(G64gat), .Z(new_n602));
  NAND2_X1  g401(.A1(G71gat), .A2(G78gat), .ZN(new_n603));
  INV_X1    g402(.A(KEYINPUT9), .ZN(new_n604));
  NAND2_X1  g403(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  NAND2_X1  g404(.A1(new_n602), .A2(new_n605), .ZN(new_n606));
  XOR2_X1   g405(.A(G71gat), .B(G78gat), .Z(new_n607));
  XNOR2_X1  g406(.A(new_n606), .B(new_n607), .ZN(new_n608));
  INV_X1    g407(.A(KEYINPUT21), .ZN(new_n609));
  NAND2_X1  g408(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  NAND2_X1  g409(.A1(G231gat), .A2(G233gat), .ZN(new_n611));
  XNOR2_X1  g410(.A(new_n610), .B(new_n611), .ZN(new_n612));
  XNOR2_X1  g411(.A(new_n612), .B(new_n346), .ZN(new_n613));
  INV_X1    g412(.A(KEYINPUT96), .ZN(new_n614));
  XNOR2_X1  g413(.A(new_n608), .B(new_n614), .ZN(new_n615));
  AOI21_X1  g414(.A(new_n567), .B1(KEYINPUT21), .B2(new_n615), .ZN(new_n616));
  AND2_X1   g415(.A1(new_n613), .A2(new_n616), .ZN(new_n617));
  NOR2_X1   g416(.A1(new_n613), .A2(new_n616), .ZN(new_n618));
  OAI21_X1  g417(.A(new_n601), .B1(new_n617), .B2(new_n618), .ZN(new_n619));
  OR2_X1    g418(.A1(new_n613), .A2(new_n616), .ZN(new_n620));
  NAND2_X1  g419(.A1(new_n613), .A2(new_n616), .ZN(new_n621));
  NAND3_X1  g420(.A1(new_n620), .A2(new_n621), .A3(new_n600), .ZN(new_n622));
  NAND2_X1  g421(.A1(new_n619), .A2(new_n622), .ZN(new_n623));
  NAND2_X1  g422(.A1(G85gat), .A2(G92gat), .ZN(new_n624));
  XNOR2_X1  g423(.A(new_n624), .B(KEYINPUT7), .ZN(new_n625));
  NAND2_X1  g424(.A1(G99gat), .A2(G106gat), .ZN(new_n626));
  INV_X1    g425(.A(G85gat), .ZN(new_n627));
  INV_X1    g426(.A(G92gat), .ZN(new_n628));
  AOI22_X1  g427(.A1(KEYINPUT8), .A2(new_n626), .B1(new_n627), .B2(new_n628), .ZN(new_n629));
  NAND2_X1  g428(.A1(new_n625), .A2(new_n629), .ZN(new_n630));
  XNOR2_X1  g429(.A(G99gat), .B(G106gat), .ZN(new_n631));
  XNOR2_X1  g430(.A(new_n630), .B(new_n631), .ZN(new_n632));
  INV_X1    g431(.A(new_n632), .ZN(new_n633));
  OAI21_X1  g432(.A(new_n633), .B1(new_n563), .B2(new_n565), .ZN(new_n634));
  AND2_X1   g433(.A1(G232gat), .A2(G233gat), .ZN(new_n635));
  AOI22_X1  g434(.A1(new_n562), .A2(new_n632), .B1(KEYINPUT41), .B2(new_n635), .ZN(new_n636));
  NAND2_X1  g435(.A1(new_n634), .A2(new_n636), .ZN(new_n637));
  XOR2_X1   g436(.A(G190gat), .B(G218gat), .Z(new_n638));
  INV_X1    g437(.A(new_n638), .ZN(new_n639));
  XNOR2_X1  g438(.A(new_n637), .B(new_n639), .ZN(new_n640));
  NOR2_X1   g439(.A1(new_n635), .A2(KEYINPUT41), .ZN(new_n641));
  XNOR2_X1  g440(.A(G134gat), .B(G162gat), .ZN(new_n642));
  XNOR2_X1  g441(.A(new_n641), .B(new_n642), .ZN(new_n643));
  XNOR2_X1  g442(.A(new_n640), .B(new_n643), .ZN(new_n644));
  INV_X1    g443(.A(KEYINPUT97), .ZN(new_n645));
  XNOR2_X1  g444(.A(new_n608), .B(KEYINPUT96), .ZN(new_n646));
  NAND2_X1  g445(.A1(new_n632), .A2(KEYINPUT10), .ZN(new_n647));
  NOR2_X1   g446(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  OR2_X1    g447(.A1(new_n632), .A2(new_n608), .ZN(new_n649));
  NAND2_X1  g448(.A1(new_n632), .A2(new_n608), .ZN(new_n650));
  AOI21_X1  g449(.A(KEYINPUT10), .B1(new_n649), .B2(new_n650), .ZN(new_n651));
  OAI21_X1  g450(.A(new_n645), .B1(new_n648), .B2(new_n651), .ZN(new_n652));
  XNOR2_X1  g451(.A(new_n632), .B(new_n608), .ZN(new_n653));
  INV_X1    g452(.A(KEYINPUT10), .ZN(new_n654));
  NAND2_X1  g453(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  NAND3_X1  g454(.A1(new_n615), .A2(KEYINPUT10), .A3(new_n632), .ZN(new_n656));
  NAND3_X1  g455(.A1(new_n655), .A2(new_n656), .A3(KEYINPUT97), .ZN(new_n657));
  NAND2_X1  g456(.A1(G230gat), .A2(G233gat), .ZN(new_n658));
  NAND3_X1  g457(.A1(new_n652), .A2(new_n657), .A3(new_n658), .ZN(new_n659));
  XNOR2_X1  g458(.A(G120gat), .B(G148gat), .ZN(new_n660));
  XNOR2_X1  g459(.A(G176gat), .B(G204gat), .ZN(new_n661));
  XOR2_X1   g460(.A(new_n660), .B(new_n661), .Z(new_n662));
  OAI211_X1 g461(.A(new_n659), .B(new_n662), .C1(new_n653), .C2(new_n658), .ZN(new_n663));
  XOR2_X1   g462(.A(new_n662), .B(KEYINPUT98), .Z(new_n664));
  NOR2_X1   g463(.A1(new_n648), .A2(new_n651), .ZN(new_n665));
  INV_X1    g464(.A(new_n658), .ZN(new_n666));
  NOR2_X1   g465(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  NOR2_X1   g466(.A1(new_n653), .A2(new_n658), .ZN(new_n668));
  OAI21_X1  g467(.A(new_n664), .B1(new_n667), .B2(new_n668), .ZN(new_n669));
  NAND2_X1  g468(.A1(new_n663), .A2(new_n669), .ZN(new_n670));
  INV_X1    g469(.A(new_n670), .ZN(new_n671));
  AND3_X1   g470(.A1(new_n623), .A2(new_n644), .A3(new_n671), .ZN(new_n672));
  NAND3_X1  g471(.A1(new_n531), .A2(new_n595), .A3(new_n672), .ZN(new_n673));
  NOR2_X1   g472(.A1(new_n673), .A2(new_n459), .ZN(new_n674));
  XNOR2_X1  g473(.A(KEYINPUT99), .B(G1gat), .ZN(new_n675));
  XNOR2_X1  g474(.A(new_n674), .B(new_n675), .ZN(G1324gat));
  NOR2_X1   g475(.A1(new_n673), .A2(new_n421), .ZN(new_n677));
  NOR2_X1   g476(.A1(new_n677), .A2(KEYINPUT100), .ZN(new_n678));
  INV_X1    g477(.A(new_n678), .ZN(new_n679));
  NAND2_X1  g478(.A1(new_n677), .A2(KEYINPUT100), .ZN(new_n680));
  AND3_X1   g479(.A1(new_n679), .A2(G8gat), .A3(new_n680), .ZN(new_n681));
  XOR2_X1   g480(.A(KEYINPUT16), .B(G8gat), .Z(new_n682));
  AND2_X1   g481(.A1(new_n682), .A2(KEYINPUT42), .ZN(new_n683));
  AOI21_X1  g482(.A(new_n681), .B1(new_n677), .B2(new_n683), .ZN(new_n684));
  INV_X1    g483(.A(new_n682), .ZN(new_n685));
  AOI21_X1  g484(.A(new_n685), .B1(new_n679), .B2(new_n680), .ZN(new_n686));
  NOR2_X1   g485(.A1(new_n686), .A2(KEYINPUT42), .ZN(new_n687));
  AND2_X1   g486(.A1(new_n687), .A2(KEYINPUT101), .ZN(new_n688));
  NOR2_X1   g487(.A1(new_n687), .A2(KEYINPUT101), .ZN(new_n689));
  OAI21_X1  g488(.A(new_n684), .B1(new_n688), .B2(new_n689), .ZN(G1325gat));
  NAND3_X1  g489(.A1(new_n383), .A2(new_n522), .A3(new_n385), .ZN(new_n691));
  NAND2_X1  g490(.A1(new_n691), .A2(KEYINPUT72), .ZN(new_n692));
  OR2_X1    g491(.A1(new_n463), .A2(KEYINPUT36), .ZN(new_n693));
  NAND3_X1  g492(.A1(new_n692), .A2(new_n693), .A3(new_n524), .ZN(new_n694));
  OAI21_X1  g493(.A(G15gat), .B1(new_n673), .B2(new_n694), .ZN(new_n695));
  INV_X1    g494(.A(G15gat), .ZN(new_n696));
  NAND2_X1  g495(.A1(new_n463), .A2(new_n696), .ZN(new_n697));
  OAI21_X1  g496(.A(new_n695), .B1(new_n673), .B2(new_n697), .ZN(G1326gat));
  NOR2_X1   g497(.A1(new_n673), .A2(new_n282), .ZN(new_n699));
  XOR2_X1   g498(.A(KEYINPUT43), .B(G22gat), .Z(new_n700));
  XNOR2_X1  g499(.A(new_n699), .B(new_n700), .ZN(G1327gat));
  INV_X1    g500(.A(KEYINPUT106), .ZN(new_n702));
  OAI211_X1 g501(.A(new_n521), .B(new_n694), .C1(new_n518), .C2(new_n519), .ZN(new_n703));
  NAND2_X1  g502(.A1(new_n703), .A2(KEYINPUT104), .ZN(new_n704));
  NAND2_X1  g503(.A1(new_n496), .A2(new_n517), .ZN(new_n705));
  NAND2_X1  g504(.A1(new_n705), .A2(KEYINPUT89), .ZN(new_n706));
  NAND3_X1  g505(.A1(new_n496), .A2(new_n517), .A3(new_n497), .ZN(new_n707));
  NAND2_X1  g506(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  INV_X1    g507(.A(KEYINPUT104), .ZN(new_n709));
  NAND4_X1  g508(.A1(new_n708), .A2(new_n709), .A3(new_n521), .A4(new_n694), .ZN(new_n710));
  OAI21_X1  g509(.A(new_n386), .B1(new_n275), .B2(new_n281), .ZN(new_n711));
  NOR3_X1   g510(.A1(new_n711), .A2(new_n526), .A3(new_n527), .ZN(new_n712));
  INV_X1    g511(.A(new_n460), .ZN(new_n713));
  AOI21_X1  g512(.A(new_n465), .B1(new_n712), .B2(new_n713), .ZN(new_n714));
  NOR2_X1   g513(.A1(new_n464), .A2(new_n466), .ZN(new_n715));
  OAI21_X1  g514(.A(KEYINPUT105), .B1(new_n714), .B2(new_n715), .ZN(new_n716));
  INV_X1    g515(.A(KEYINPUT105), .ZN(new_n717));
  NAND3_X1  g516(.A1(new_n461), .A2(new_n467), .A3(new_n717), .ZN(new_n718));
  NAND2_X1  g517(.A1(new_n716), .A2(new_n718), .ZN(new_n719));
  NAND3_X1  g518(.A1(new_n704), .A2(new_n710), .A3(new_n719), .ZN(new_n720));
  NOR2_X1   g519(.A1(new_n644), .A2(KEYINPUT44), .ZN(new_n721));
  INV_X1    g520(.A(new_n644), .ZN(new_n722));
  NAND2_X1  g521(.A1(new_n531), .A2(new_n722), .ZN(new_n723));
  AOI22_X1  g522(.A1(new_n720), .A2(new_n721), .B1(new_n723), .B2(KEYINPUT44), .ZN(new_n724));
  AND3_X1   g523(.A1(new_n591), .A2(KEYINPUT103), .A3(new_n593), .ZN(new_n725));
  AOI21_X1  g524(.A(KEYINPUT103), .B1(new_n591), .B2(new_n593), .ZN(new_n726));
  NOR2_X1   g525(.A1(new_n725), .A2(new_n726), .ZN(new_n727));
  INV_X1    g526(.A(new_n727), .ZN(new_n728));
  NOR2_X1   g527(.A1(new_n623), .A2(new_n670), .ZN(new_n729));
  INV_X1    g528(.A(new_n729), .ZN(new_n730));
  NOR2_X1   g529(.A1(new_n728), .A2(new_n730), .ZN(new_n731));
  INV_X1    g530(.A(new_n731), .ZN(new_n732));
  OAI21_X1  g531(.A(new_n702), .B1(new_n724), .B2(new_n732), .ZN(new_n733));
  INV_X1    g532(.A(new_n721), .ZN(new_n734));
  AOI22_X1  g533(.A1(new_n703), .A2(KEYINPUT104), .B1(new_n716), .B2(new_n718), .ZN(new_n735));
  AOI21_X1  g534(.A(new_n734), .B1(new_n735), .B2(new_n710), .ZN(new_n736));
  INV_X1    g535(.A(KEYINPUT44), .ZN(new_n737));
  AOI21_X1  g536(.A(new_n737), .B1(new_n531), .B2(new_n722), .ZN(new_n738));
  OAI211_X1 g537(.A(KEYINPUT106), .B(new_n731), .C1(new_n736), .C2(new_n738), .ZN(new_n739));
  NAND2_X1  g538(.A1(new_n733), .A2(new_n739), .ZN(new_n740));
  OAI21_X1  g539(.A(G29gat), .B1(new_n740), .B2(new_n459), .ZN(new_n741));
  AND4_X1   g540(.A1(new_n531), .A2(new_n595), .A3(new_n722), .A4(new_n729), .ZN(new_n742));
  INV_X1    g541(.A(new_n459), .ZN(new_n743));
  NAND3_X1  g542(.A1(new_n742), .A2(new_n554), .A3(new_n743), .ZN(new_n744));
  XOR2_X1   g543(.A(KEYINPUT102), .B(KEYINPUT45), .Z(new_n745));
  XNOR2_X1  g544(.A(new_n744), .B(new_n745), .ZN(new_n746));
  NAND2_X1  g545(.A1(new_n741), .A2(new_n746), .ZN(G1328gat));
  OAI21_X1  g546(.A(G36gat), .B1(new_n740), .B2(new_n421), .ZN(new_n748));
  NAND3_X1  g547(.A1(new_n742), .A2(new_n550), .A3(new_n504), .ZN(new_n749));
  XOR2_X1   g548(.A(new_n749), .B(KEYINPUT46), .Z(new_n750));
  NAND2_X1  g549(.A1(new_n748), .A2(new_n750), .ZN(G1329gat));
  INV_X1    g550(.A(G43gat), .ZN(new_n752));
  AND3_X1   g551(.A1(new_n742), .A2(new_n752), .A3(new_n463), .ZN(new_n753));
  INV_X1    g552(.A(new_n694), .ZN(new_n754));
  NAND3_X1  g553(.A1(new_n733), .A2(new_n754), .A3(new_n739), .ZN(new_n755));
  AOI21_X1  g554(.A(new_n753), .B1(new_n755), .B2(G43gat), .ZN(new_n756));
  NOR2_X1   g555(.A1(new_n724), .A2(new_n732), .ZN(new_n757));
  AOI21_X1  g556(.A(new_n752), .B1(new_n757), .B2(new_n754), .ZN(new_n758));
  INV_X1    g557(.A(KEYINPUT47), .ZN(new_n759));
  OR2_X1    g558(.A1(new_n753), .A2(new_n759), .ZN(new_n760));
  OAI22_X1  g559(.A1(new_n756), .A2(KEYINPUT47), .B1(new_n758), .B2(new_n760), .ZN(G1330gat));
  INV_X1    g560(.A(KEYINPUT107), .ZN(new_n762));
  NAND3_X1  g561(.A1(new_n733), .A2(new_n502), .A3(new_n739), .ZN(new_n763));
  NAND2_X1  g562(.A1(new_n763), .A2(G50gat), .ZN(new_n764));
  OR2_X1    g563(.A1(new_n282), .A2(G50gat), .ZN(new_n765));
  INV_X1    g564(.A(new_n765), .ZN(new_n766));
  NAND2_X1  g565(.A1(new_n742), .A2(new_n766), .ZN(new_n767));
  INV_X1    g566(.A(KEYINPUT48), .ZN(new_n768));
  NAND2_X1  g567(.A1(new_n767), .A2(new_n768), .ZN(new_n769));
  INV_X1    g568(.A(new_n769), .ZN(new_n770));
  NAND2_X1  g569(.A1(new_n764), .A2(new_n770), .ZN(new_n771));
  OAI211_X1 g570(.A(new_n502), .B(new_n731), .C1(new_n736), .C2(new_n738), .ZN(new_n772));
  NAND2_X1  g571(.A1(new_n772), .A2(G50gat), .ZN(new_n773));
  AOI21_X1  g572(.A(new_n768), .B1(new_n773), .B2(new_n767), .ZN(new_n774));
  INV_X1    g573(.A(new_n774), .ZN(new_n775));
  AOI21_X1  g574(.A(new_n762), .B1(new_n771), .B2(new_n775), .ZN(new_n776));
  AOI21_X1  g575(.A(new_n769), .B1(new_n763), .B2(G50gat), .ZN(new_n777));
  NOR3_X1   g576(.A1(new_n777), .A2(KEYINPUT107), .A3(new_n774), .ZN(new_n778));
  NOR2_X1   g577(.A1(new_n776), .A2(new_n778), .ZN(G1331gat));
  NAND4_X1  g578(.A1(new_n728), .A2(new_n623), .A3(new_n644), .A4(new_n670), .ZN(new_n780));
  AOI21_X1  g579(.A(new_n780), .B1(new_n735), .B2(new_n710), .ZN(new_n781));
  NAND2_X1  g580(.A1(new_n781), .A2(new_n743), .ZN(new_n782));
  XNOR2_X1  g581(.A(new_n782), .B(G57gat), .ZN(G1332gat));
  XOR2_X1   g582(.A(new_n781), .B(KEYINPUT108), .Z(new_n784));
  XNOR2_X1  g583(.A(new_n421), .B(KEYINPUT109), .ZN(new_n785));
  AOI21_X1  g584(.A(new_n785), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n786));
  NAND2_X1  g585(.A1(new_n784), .A2(new_n786), .ZN(new_n787));
  NOR2_X1   g586(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n788));
  XOR2_X1   g587(.A(new_n787), .B(new_n788), .Z(G1333gat));
  AOI21_X1  g588(.A(G71gat), .B1(new_n781), .B2(new_n463), .ZN(new_n790));
  AND2_X1   g589(.A1(new_n754), .A2(G71gat), .ZN(new_n791));
  AOI21_X1  g590(.A(new_n790), .B1(new_n784), .B2(new_n791), .ZN(new_n792));
  XNOR2_X1  g591(.A(KEYINPUT110), .B(KEYINPUT50), .ZN(new_n793));
  XNOR2_X1  g592(.A(new_n792), .B(new_n793), .ZN(G1334gat));
  NAND2_X1  g593(.A1(new_n784), .A2(new_n502), .ZN(new_n795));
  XNOR2_X1  g594(.A(new_n795), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g595(.A1(new_n727), .A2(new_n623), .ZN(new_n797));
  NAND3_X1  g596(.A1(new_n720), .A2(new_n722), .A3(new_n797), .ZN(new_n798));
  NAND2_X1  g597(.A1(new_n798), .A2(KEYINPUT51), .ZN(new_n799));
  INV_X1    g598(.A(KEYINPUT51), .ZN(new_n800));
  NAND4_X1  g599(.A1(new_n720), .A2(new_n800), .A3(new_n722), .A4(new_n797), .ZN(new_n801));
  AND3_X1   g600(.A1(new_n799), .A2(new_n670), .A3(new_n801), .ZN(new_n802));
  NAND3_X1  g601(.A1(new_n802), .A2(new_n627), .A3(new_n743), .ZN(new_n803));
  NOR3_X1   g602(.A1(new_n727), .A2(new_n623), .A3(new_n671), .ZN(new_n804));
  OAI21_X1  g603(.A(new_n804), .B1(new_n736), .B2(new_n738), .ZN(new_n805));
  OAI21_X1  g604(.A(G85gat), .B1(new_n805), .B2(new_n459), .ZN(new_n806));
  NAND2_X1  g605(.A1(new_n803), .A2(new_n806), .ZN(G1336gat));
  INV_X1    g606(.A(new_n785), .ZN(new_n808));
  NAND3_X1  g607(.A1(new_n802), .A2(new_n628), .A3(new_n808), .ZN(new_n809));
  INV_X1    g608(.A(KEYINPUT52), .ZN(new_n810));
  OAI21_X1  g609(.A(G92gat), .B1(new_n805), .B2(new_n785), .ZN(new_n811));
  NAND3_X1  g610(.A1(new_n809), .A2(new_n810), .A3(new_n811), .ZN(new_n812));
  OAI21_X1  g611(.A(G92gat), .B1(new_n805), .B2(new_n421), .ZN(new_n813));
  AND2_X1   g612(.A1(new_n809), .A2(new_n813), .ZN(new_n814));
  OAI21_X1  g613(.A(new_n812), .B1(new_n814), .B2(new_n810), .ZN(G1337gat));
  INV_X1    g614(.A(G99gat), .ZN(new_n816));
  NOR3_X1   g615(.A1(new_n805), .A2(new_n816), .A3(new_n694), .ZN(new_n817));
  NAND2_X1  g616(.A1(new_n802), .A2(new_n463), .ZN(new_n818));
  AOI21_X1  g617(.A(new_n817), .B1(new_n818), .B2(new_n816), .ZN(G1338gat));
  OR2_X1    g618(.A1(new_n282), .A2(G106gat), .ZN(new_n820));
  INV_X1    g619(.A(new_n820), .ZN(new_n821));
  NAND4_X1  g620(.A1(new_n799), .A2(new_n670), .A3(new_n801), .A4(new_n821), .ZN(new_n822));
  OAI211_X1 g621(.A(new_n502), .B(new_n804), .C1(new_n736), .C2(new_n738), .ZN(new_n823));
  NAND2_X1  g622(.A1(new_n823), .A2(G106gat), .ZN(new_n824));
  INV_X1    g623(.A(KEYINPUT53), .ZN(new_n825));
  NAND3_X1  g624(.A1(new_n822), .A2(new_n824), .A3(new_n825), .ZN(new_n826));
  NAND2_X1  g625(.A1(new_n824), .A2(KEYINPUT111), .ZN(new_n827));
  INV_X1    g626(.A(KEYINPUT111), .ZN(new_n828));
  NAND3_X1  g627(.A1(new_n823), .A2(new_n828), .A3(G106gat), .ZN(new_n829));
  NAND3_X1  g628(.A1(new_n827), .A2(new_n829), .A3(new_n822), .ZN(new_n830));
  INV_X1    g629(.A(KEYINPUT112), .ZN(new_n831));
  AND3_X1   g630(.A1(new_n830), .A2(new_n831), .A3(KEYINPUT53), .ZN(new_n832));
  AOI21_X1  g631(.A(new_n831), .B1(new_n830), .B2(KEYINPUT53), .ZN(new_n833));
  OAI21_X1  g632(.A(new_n826), .B1(new_n832), .B2(new_n833), .ZN(G1339gat));
  INV_X1    g633(.A(new_n623), .ZN(new_n835));
  INV_X1    g634(.A(KEYINPUT103), .ZN(new_n836));
  NAND2_X1  g635(.A1(new_n594), .A2(new_n836), .ZN(new_n837));
  NAND3_X1  g636(.A1(new_n591), .A2(KEYINPUT103), .A3(new_n593), .ZN(new_n838));
  INV_X1    g637(.A(KEYINPUT54), .ZN(new_n839));
  OAI211_X1 g638(.A(new_n839), .B(new_n658), .C1(new_n648), .C2(new_n651), .ZN(new_n840));
  INV_X1    g639(.A(new_n662), .ZN(new_n841));
  NAND2_X1  g640(.A1(new_n840), .A2(new_n841), .ZN(new_n842));
  AOI21_X1  g641(.A(new_n839), .B1(new_n665), .B2(new_n666), .ZN(new_n843));
  AOI21_X1  g642(.A(new_n842), .B1(new_n843), .B2(new_n659), .ZN(new_n844));
  AND2_X1   g643(.A1(new_n844), .A2(KEYINPUT55), .ZN(new_n845));
  OAI21_X1  g644(.A(new_n663), .B1(new_n844), .B2(KEYINPUT55), .ZN(new_n846));
  NOR2_X1   g645(.A1(new_n845), .A2(new_n846), .ZN(new_n847));
  NAND3_X1  g646(.A1(new_n837), .A2(new_n838), .A3(new_n847), .ZN(new_n848));
  NOR2_X1   g647(.A1(new_n578), .A2(new_n579), .ZN(new_n849));
  AOI21_X1  g648(.A(new_n571), .B1(new_n566), .B2(new_n568), .ZN(new_n850));
  OAI21_X1  g649(.A(new_n535), .B1(new_n849), .B2(new_n850), .ZN(new_n851));
  NAND3_X1  g650(.A1(new_n590), .A2(new_n670), .A3(new_n851), .ZN(new_n852));
  XNOR2_X1  g651(.A(new_n852), .B(KEYINPUT113), .ZN(new_n853));
  INV_X1    g652(.A(new_n853), .ZN(new_n854));
  AOI21_X1  g653(.A(new_n722), .B1(new_n848), .B2(new_n854), .ZN(new_n855));
  NAND4_X1  g654(.A1(new_n847), .A2(new_n590), .A3(new_n722), .A4(new_n851), .ZN(new_n856));
  INV_X1    g655(.A(new_n856), .ZN(new_n857));
  OAI21_X1  g656(.A(new_n835), .B1(new_n855), .B2(new_n857), .ZN(new_n858));
  INV_X1    g657(.A(new_n672), .ZN(new_n859));
  NOR2_X1   g658(.A1(new_n727), .A2(new_n859), .ZN(new_n860));
  INV_X1    g659(.A(new_n860), .ZN(new_n861));
  AOI21_X1  g660(.A(new_n459), .B1(new_n858), .B2(new_n861), .ZN(new_n862));
  AND2_X1   g661(.A1(new_n862), .A2(new_n712), .ZN(new_n863));
  NAND3_X1  g662(.A1(new_n863), .A2(new_n727), .A3(new_n785), .ZN(new_n864));
  AOI21_X1  g663(.A(new_n464), .B1(new_n858), .B2(new_n861), .ZN(new_n865));
  NOR2_X1   g664(.A1(new_n808), .A2(new_n459), .ZN(new_n866));
  AND2_X1   g665(.A1(new_n865), .A2(new_n866), .ZN(new_n867));
  NOR2_X1   g666(.A1(new_n594), .A2(new_n335), .ZN(new_n868));
  AOI22_X1  g667(.A1(new_n864), .A2(new_n335), .B1(new_n867), .B2(new_n868), .ZN(G1340gat));
  NAND3_X1  g668(.A1(new_n867), .A2(G120gat), .A3(new_n670), .ZN(new_n870));
  AND3_X1   g669(.A1(new_n863), .A2(new_n670), .A3(new_n785), .ZN(new_n871));
  OAI21_X1  g670(.A(new_n870), .B1(new_n871), .B2(G120gat), .ZN(new_n872));
  XNOR2_X1  g671(.A(new_n872), .B(KEYINPUT114), .ZN(G1341gat));
  NAND3_X1  g672(.A1(new_n867), .A2(G127gat), .A3(new_n623), .ZN(new_n874));
  NAND4_X1  g673(.A1(new_n862), .A2(new_n712), .A3(new_n623), .A4(new_n785), .ZN(new_n875));
  AND2_X1   g674(.A1(new_n875), .A2(KEYINPUT115), .ZN(new_n876));
  OAI21_X1  g675(.A(new_n346), .B1(new_n875), .B2(KEYINPUT115), .ZN(new_n877));
  OAI21_X1  g676(.A(new_n874), .B1(new_n876), .B2(new_n877), .ZN(new_n878));
  XNOR2_X1  g677(.A(new_n878), .B(KEYINPUT116), .ZN(G1342gat));
  NOR2_X1   g678(.A1(new_n644), .A2(new_n504), .ZN(new_n880));
  NAND4_X1  g679(.A1(new_n863), .A2(new_n348), .A3(new_n350), .A4(new_n880), .ZN(new_n881));
  AND2_X1   g680(.A1(new_n881), .A2(KEYINPUT56), .ZN(new_n882));
  AOI21_X1  g681(.A(new_n347), .B1(new_n867), .B2(new_n722), .ZN(new_n883));
  NOR2_X1   g682(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  OAI21_X1  g683(.A(new_n884), .B1(KEYINPUT56), .B2(new_n881), .ZN(G1343gat));
  NOR2_X1   g684(.A1(new_n754), .A2(new_n282), .ZN(new_n886));
  NAND3_X1  g685(.A1(new_n862), .A2(new_n785), .A3(new_n886), .ZN(new_n887));
  NOR3_X1   g686(.A1(new_n887), .A2(G141gat), .A3(new_n594), .ZN(new_n888));
  NOR2_X1   g687(.A1(new_n888), .A2(KEYINPUT58), .ZN(new_n889));
  NAND3_X1  g688(.A1(new_n847), .A2(new_n591), .A3(new_n593), .ZN(new_n890));
  AOI21_X1  g689(.A(new_n722), .B1(new_n890), .B2(new_n852), .ZN(new_n891));
  OAI21_X1  g690(.A(new_n835), .B1(new_n891), .B2(new_n857), .ZN(new_n892));
  INV_X1    g691(.A(KEYINPUT117), .ZN(new_n893));
  AOI21_X1  g692(.A(new_n860), .B1(new_n892), .B2(new_n893), .ZN(new_n894));
  OAI211_X1 g693(.A(KEYINPUT117), .B(new_n835), .C1(new_n891), .C2(new_n857), .ZN(new_n895));
  NAND2_X1  g694(.A1(new_n894), .A2(new_n895), .ZN(new_n896));
  NAND2_X1  g695(.A1(new_n502), .A2(KEYINPUT57), .ZN(new_n897));
  INV_X1    g696(.A(new_n897), .ZN(new_n898));
  NAND2_X1  g697(.A1(new_n896), .A2(new_n898), .ZN(new_n899));
  AOI21_X1  g698(.A(new_n282), .B1(new_n858), .B2(new_n861), .ZN(new_n900));
  OAI21_X1  g699(.A(new_n899), .B1(new_n900), .B2(KEYINPUT57), .ZN(new_n901));
  NAND2_X1  g700(.A1(new_n866), .A2(new_n694), .ZN(new_n902));
  INV_X1    g701(.A(new_n902), .ZN(new_n903));
  NAND3_X1  g702(.A1(new_n901), .A2(new_n595), .A3(new_n903), .ZN(new_n904));
  INV_X1    g703(.A(KEYINPUT119), .ZN(new_n905));
  NAND2_X1  g704(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  NAND2_X1  g705(.A1(new_n906), .A2(G141gat), .ZN(new_n907));
  NOR2_X1   g706(.A1(new_n904), .A2(new_n905), .ZN(new_n908));
  OAI21_X1  g707(.A(new_n889), .B1(new_n907), .B2(new_n908), .ZN(new_n909));
  AOI21_X1  g708(.A(new_n897), .B1(new_n894), .B2(new_n895), .ZN(new_n910));
  INV_X1    g709(.A(new_n847), .ZN(new_n911));
  NOR3_X1   g710(.A1(new_n725), .A2(new_n726), .A3(new_n911), .ZN(new_n912));
  OAI21_X1  g711(.A(new_n644), .B1(new_n912), .B2(new_n853), .ZN(new_n913));
  AOI21_X1  g712(.A(new_n623), .B1(new_n913), .B2(new_n856), .ZN(new_n914));
  OAI21_X1  g713(.A(new_n502), .B1(new_n914), .B2(new_n860), .ZN(new_n915));
  INV_X1    g714(.A(KEYINPUT57), .ZN(new_n916));
  AOI21_X1  g715(.A(new_n910), .B1(new_n915), .B2(new_n916), .ZN(new_n917));
  OAI21_X1  g716(.A(KEYINPUT118), .B1(new_n917), .B2(new_n902), .ZN(new_n918));
  INV_X1    g717(.A(KEYINPUT118), .ZN(new_n919));
  NAND3_X1  g718(.A1(new_n901), .A2(new_n919), .A3(new_n903), .ZN(new_n920));
  NAND3_X1  g719(.A1(new_n918), .A2(new_n727), .A3(new_n920), .ZN(new_n921));
  AOI21_X1  g720(.A(new_n888), .B1(new_n921), .B2(G141gat), .ZN(new_n922));
  INV_X1    g721(.A(KEYINPUT58), .ZN(new_n923));
  OAI21_X1  g722(.A(new_n909), .B1(new_n922), .B2(new_n923), .ZN(G1344gat));
  NAND2_X1  g723(.A1(new_n594), .A2(new_n672), .ZN(new_n925));
  XNOR2_X1  g724(.A(new_n925), .B(KEYINPUT120), .ZN(new_n926));
  NAND2_X1  g725(.A1(new_n926), .A2(new_n892), .ZN(new_n927));
  INV_X1    g726(.A(KEYINPUT121), .ZN(new_n928));
  AOI21_X1  g727(.A(new_n282), .B1(new_n927), .B2(new_n928), .ZN(new_n929));
  NAND3_X1  g728(.A1(new_n926), .A2(KEYINPUT121), .A3(new_n892), .ZN(new_n930));
  AOI21_X1  g729(.A(KEYINPUT57), .B1(new_n929), .B2(new_n930), .ZN(new_n931));
  AOI21_X1  g730(.A(new_n897), .B1(new_n858), .B2(new_n861), .ZN(new_n932));
  OAI211_X1 g731(.A(new_n670), .B(new_n903), .C1(new_n931), .C2(new_n932), .ZN(new_n933));
  INV_X1    g732(.A(new_n933), .ZN(new_n934));
  OAI21_X1  g733(.A(KEYINPUT59), .B1(new_n934), .B2(new_n232), .ZN(new_n935));
  AND3_X1   g734(.A1(new_n918), .A2(new_n670), .A3(new_n920), .ZN(new_n936));
  OR2_X1    g735(.A1(new_n232), .A2(KEYINPUT59), .ZN(new_n937));
  OAI21_X1  g736(.A(new_n935), .B1(new_n936), .B2(new_n937), .ZN(new_n938));
  OR3_X1    g737(.A1(new_n887), .A2(G148gat), .A3(new_n671), .ZN(new_n939));
  NAND2_X1  g738(.A1(new_n938), .A2(new_n939), .ZN(G1345gat));
  NAND4_X1  g739(.A1(new_n918), .A2(G155gat), .A3(new_n623), .A4(new_n920), .ZN(new_n941));
  OAI21_X1  g740(.A(new_n597), .B1(new_n887), .B2(new_n835), .ZN(new_n942));
  AND3_X1   g741(.A1(new_n941), .A2(KEYINPUT122), .A3(new_n942), .ZN(new_n943));
  AOI21_X1  g742(.A(KEYINPUT122), .B1(new_n941), .B2(new_n942), .ZN(new_n944));
  NOR2_X1   g743(.A1(new_n943), .A2(new_n944), .ZN(G1346gat));
  INV_X1    g744(.A(G162gat), .ZN(new_n946));
  NAND4_X1  g745(.A1(new_n862), .A2(new_n946), .A3(new_n880), .A4(new_n886), .ZN(new_n947));
  AND3_X1   g746(.A1(new_n918), .A2(new_n722), .A3(new_n920), .ZN(new_n948));
  OAI21_X1  g747(.A(new_n947), .B1(new_n948), .B2(new_n946), .ZN(G1347gat));
  AOI21_X1  g748(.A(new_n743), .B1(new_n858), .B2(new_n861), .ZN(new_n950));
  NOR2_X1   g749(.A1(new_n785), .A2(new_n387), .ZN(new_n951));
  NAND2_X1  g750(.A1(new_n950), .A2(new_n951), .ZN(new_n952));
  INV_X1    g751(.A(new_n952), .ZN(new_n953));
  AOI21_X1  g752(.A(G169gat), .B1(new_n953), .B2(new_n727), .ZN(new_n954));
  NOR2_X1   g753(.A1(new_n743), .A2(new_n421), .ZN(new_n955));
  AND2_X1   g754(.A1(new_n865), .A2(new_n955), .ZN(new_n956));
  AND2_X1   g755(.A1(new_n595), .A2(G169gat), .ZN(new_n957));
  AOI21_X1  g756(.A(new_n954), .B1(new_n956), .B2(new_n957), .ZN(G1348gat));
  INV_X1    g757(.A(new_n956), .ZN(new_n959));
  OAI21_X1  g758(.A(G176gat), .B1(new_n959), .B2(new_n671), .ZN(new_n960));
  INV_X1    g759(.A(G176gat), .ZN(new_n961));
  NAND3_X1  g760(.A1(new_n953), .A2(new_n961), .A3(new_n670), .ZN(new_n962));
  NAND2_X1  g761(.A1(new_n960), .A2(new_n962), .ZN(G1349gat));
  NAND3_X1  g762(.A1(new_n865), .A2(new_n623), .A3(new_n955), .ZN(new_n964));
  AOI21_X1  g763(.A(new_n312), .B1(new_n964), .B2(KEYINPUT123), .ZN(new_n965));
  OAI21_X1  g764(.A(new_n965), .B1(KEYINPUT123), .B2(new_n964), .ZN(new_n966));
  NAND4_X1  g765(.A1(new_n953), .A2(new_n314), .A3(new_n317), .A4(new_n623), .ZN(new_n967));
  NAND2_X1  g766(.A1(new_n966), .A2(new_n967), .ZN(new_n968));
  XNOR2_X1  g767(.A(new_n968), .B(KEYINPUT60), .ZN(G1350gat));
  NAND3_X1  g768(.A1(new_n953), .A2(new_n321), .A3(new_n722), .ZN(new_n970));
  OAI21_X1  g769(.A(G190gat), .B1(new_n959), .B2(new_n644), .ZN(new_n971));
  AND2_X1   g770(.A1(new_n971), .A2(KEYINPUT61), .ZN(new_n972));
  NOR2_X1   g771(.A1(new_n971), .A2(KEYINPUT61), .ZN(new_n973));
  OAI21_X1  g772(.A(new_n970), .B1(new_n972), .B2(new_n973), .ZN(G1351gat));
  NAND2_X1  g773(.A1(new_n886), .A2(new_n808), .ZN(new_n975));
  XNOR2_X1  g774(.A(new_n975), .B(KEYINPUT124), .ZN(new_n976));
  AND2_X1   g775(.A1(new_n976), .A2(new_n950), .ZN(new_n977));
  AOI21_X1  g776(.A(G197gat), .B1(new_n977), .B2(new_n727), .ZN(new_n978));
  NOR2_X1   g777(.A1(new_n931), .A2(new_n932), .ZN(new_n979));
  NAND2_X1  g778(.A1(new_n694), .A2(new_n955), .ZN(new_n980));
  XNOR2_X1  g779(.A(new_n980), .B(KEYINPUT125), .ZN(new_n981));
  NOR2_X1   g780(.A1(new_n979), .A2(new_n981), .ZN(new_n982));
  NOR2_X1   g781(.A1(new_n594), .A2(new_n209), .ZN(new_n983));
  AOI21_X1  g782(.A(new_n978), .B1(new_n982), .B2(new_n983), .ZN(G1352gat));
  NAND3_X1  g783(.A1(new_n977), .A2(new_n210), .A3(new_n670), .ZN(new_n985));
  OAI21_X1  g784(.A(new_n985), .B1(KEYINPUT126), .B2(KEYINPUT62), .ZN(new_n986));
  NAND2_X1  g785(.A1(KEYINPUT126), .A2(KEYINPUT62), .ZN(new_n987));
  NAND2_X1  g786(.A1(new_n986), .A2(new_n987), .ZN(new_n988));
  OR2_X1    g787(.A1(new_n931), .A2(new_n932), .ZN(new_n989));
  NAND2_X1  g788(.A1(new_n989), .A2(new_n670), .ZN(new_n990));
  OAI21_X1  g789(.A(G204gat), .B1(new_n990), .B2(new_n981), .ZN(new_n991));
  NAND3_X1  g790(.A1(new_n985), .A2(KEYINPUT126), .A3(KEYINPUT62), .ZN(new_n992));
  NAND3_X1  g791(.A1(new_n988), .A2(new_n991), .A3(new_n992), .ZN(G1353gat));
  INV_X1    g792(.A(KEYINPUT63), .ZN(new_n994));
  INV_X1    g793(.A(KEYINPUT127), .ZN(new_n995));
  INV_X1    g794(.A(new_n980), .ZN(new_n996));
  NAND2_X1  g795(.A1(new_n996), .A2(new_n623), .ZN(new_n997));
  INV_X1    g796(.A(new_n997), .ZN(new_n998));
  AOI21_X1  g797(.A(new_n995), .B1(new_n989), .B2(new_n998), .ZN(new_n999));
  OAI211_X1 g798(.A(new_n995), .B(new_n998), .C1(new_n931), .C2(new_n932), .ZN(new_n1000));
  NAND2_X1  g799(.A1(new_n1000), .A2(G211gat), .ZN(new_n1001));
  OAI21_X1  g800(.A(new_n994), .B1(new_n999), .B2(new_n1001), .ZN(new_n1002));
  OAI21_X1  g801(.A(KEYINPUT127), .B1(new_n979), .B2(new_n997), .ZN(new_n1003));
  NAND4_X1  g802(.A1(new_n1003), .A2(KEYINPUT63), .A3(G211gat), .A4(new_n1000), .ZN(new_n1004));
  NAND2_X1  g803(.A1(new_n1002), .A2(new_n1004), .ZN(new_n1005));
  INV_X1    g804(.A(G211gat), .ZN(new_n1006));
  NAND3_X1  g805(.A1(new_n977), .A2(new_n1006), .A3(new_n623), .ZN(new_n1007));
  NAND2_X1  g806(.A1(new_n1005), .A2(new_n1007), .ZN(G1354gat));
  AOI21_X1  g807(.A(G218gat), .B1(new_n977), .B2(new_n722), .ZN(new_n1009));
  AND2_X1   g808(.A1(new_n722), .A2(G218gat), .ZN(new_n1010));
  AOI21_X1  g809(.A(new_n1009), .B1(new_n982), .B2(new_n1010), .ZN(G1355gat));
endmodule


