//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 0 0 1 1 1 1 1 0 0 0 0 0 1 1 0 0 1 1 1 1 0 0 0 1 0 1 0 1 1 1 0 0 0 1 1 1 0 0 1 0 0 0 0 0 0 0 0 0 1 1 1 0 0 1 0 1 0 1 1 1 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:41:01 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n205, new_n206, new_n207, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n692, new_n693, new_n694, new_n695, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1087,
    new_n1088, new_n1089, new_n1090, new_n1091, new_n1092, new_n1093,
    new_n1094, new_n1095, new_n1096, new_n1097, new_n1098, new_n1099,
    new_n1100, new_n1101, new_n1102, new_n1103, new_n1104, new_n1105,
    new_n1106, new_n1107, new_n1109, new_n1110, new_n1111, new_n1112,
    new_n1113, new_n1114, new_n1115, new_n1116, new_n1117, new_n1118,
    new_n1119, new_n1120, new_n1121, new_n1122, new_n1123, new_n1124,
    new_n1125, new_n1126, new_n1127, new_n1128, new_n1129, new_n1130,
    new_n1131, new_n1132, new_n1133, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1186, new_n1187, new_n1188, new_n1189, new_n1190, new_n1191,
    new_n1192, new_n1193, new_n1194, new_n1195, new_n1196, new_n1197,
    new_n1198, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1251, new_n1252,
    new_n1253, new_n1254, new_n1255, new_n1256, new_n1257, new_n1258,
    new_n1259, new_n1260, new_n1261, new_n1262, new_n1263, new_n1264,
    new_n1265, new_n1266, new_n1267, new_n1268, new_n1269, new_n1270,
    new_n1272, new_n1273, new_n1274, new_n1275, new_n1276, new_n1277,
    new_n1278, new_n1279, new_n1280, new_n1281, new_n1282, new_n1283,
    new_n1284, new_n1285, new_n1286, new_n1287, new_n1288, new_n1289,
    new_n1290, new_n1292, new_n1293, new_n1295, new_n1296, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1346,
    new_n1347, new_n1348, new_n1349, new_n1350, new_n1351, new_n1352,
    new_n1353, new_n1354, new_n1355, new_n1357, new_n1358, new_n1359,
    new_n1360, new_n1361, new_n1362, new_n1363, new_n1364, new_n1365,
    new_n1366, new_n1367, new_n1368, new_n1369, new_n1370, new_n1371,
    new_n1372, new_n1373, new_n1374;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  INV_X1    g0004(.A(G97), .ZN(new_n205));
  INV_X1    g0005(.A(G107), .ZN(new_n206));
  NAND2_X1  g0006(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  NAND2_X1  g0007(.A1(new_n207), .A2(G87), .ZN(G355));
  NAND2_X1  g0008(.A1(G1), .A2(G20), .ZN(new_n209));
  NOR2_X1   g0009(.A1(new_n209), .A2(G13), .ZN(new_n210));
  OAI211_X1 g0010(.A(new_n210), .B(G250), .C1(G257), .C2(G264), .ZN(new_n211));
  XNOR2_X1  g0011(.A(new_n211), .B(KEYINPUT0), .ZN(new_n212));
  AND2_X1   g0012(.A1(KEYINPUT64), .A2(G20), .ZN(new_n213));
  NOR2_X1   g0013(.A1(KEYINPUT64), .A2(G20), .ZN(new_n214));
  NOR2_X1   g0014(.A1(new_n213), .A2(new_n214), .ZN(new_n215));
  NAND2_X1  g0015(.A1(G1), .A2(G13), .ZN(new_n216));
  NOR2_X1   g0016(.A1(new_n215), .A2(new_n216), .ZN(new_n217));
  INV_X1    g0017(.A(new_n201), .ZN(new_n218));
  NAND2_X1  g0018(.A1(new_n218), .A2(G50), .ZN(new_n219));
  INV_X1    g0019(.A(new_n219), .ZN(new_n220));
  NAND2_X1  g0020(.A1(new_n217), .A2(new_n220), .ZN(new_n221));
  XNOR2_X1  g0021(.A(KEYINPUT65), .B(G68), .ZN(new_n222));
  INV_X1    g0022(.A(G238), .ZN(new_n223));
  NOR2_X1   g0023(.A1(new_n222), .A2(new_n223), .ZN(new_n224));
  AOI22_X1  g0024(.A1(G107), .A2(G264), .B1(G116), .B2(G270), .ZN(new_n225));
  AOI22_X1  g0025(.A1(G50), .A2(G226), .B1(G77), .B2(G244), .ZN(new_n226));
  AOI22_X1  g0026(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n227));
  NAND2_X1  g0027(.A1(G58), .A2(G232), .ZN(new_n228));
  NAND4_X1  g0028(.A1(new_n225), .A2(new_n226), .A3(new_n227), .A4(new_n228), .ZN(new_n229));
  OAI21_X1  g0029(.A(new_n209), .B1(new_n224), .B2(new_n229), .ZN(new_n230));
  OAI211_X1 g0030(.A(new_n212), .B(new_n221), .C1(KEYINPUT1), .C2(new_n230), .ZN(new_n231));
  AOI21_X1  g0031(.A(new_n231), .B1(KEYINPUT1), .B2(new_n230), .ZN(G361));
  XNOR2_X1  g0032(.A(G250), .B(G257), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n233), .B(KEYINPUT66), .ZN(new_n234));
  XOR2_X1   g0034(.A(G264), .B(G270), .Z(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XNOR2_X1  g0036(.A(G238), .B(G244), .ZN(new_n237));
  INV_X1    g0037(.A(G232), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XNOR2_X1  g0039(.A(KEYINPUT2), .B(G226), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n236), .B(new_n241), .ZN(G358));
  XNOR2_X1  g0042(.A(G50), .B(G68), .ZN(new_n243));
  XNOR2_X1  g0043(.A(G58), .B(G77), .ZN(new_n244));
  XOR2_X1   g0044(.A(new_n243), .B(new_n244), .Z(new_n245));
  NAND2_X1  g0045(.A1(new_n206), .A2(G97), .ZN(new_n246));
  NAND2_X1  g0046(.A1(new_n205), .A2(G107), .ZN(new_n247));
  NAND2_X1  g0047(.A1(new_n246), .A2(new_n247), .ZN(new_n248));
  XNOR2_X1  g0048(.A(G87), .B(G116), .ZN(new_n249));
  XNOR2_X1  g0049(.A(new_n248), .B(new_n249), .ZN(new_n250));
  XNOR2_X1  g0050(.A(new_n245), .B(new_n250), .ZN(G351));
  INV_X1    g0051(.A(KEYINPUT21), .ZN(new_n252));
  INV_X1    g0052(.A(G116), .ZN(new_n253));
  NAND2_X1  g0053(.A1(new_n253), .A2(KEYINPUT80), .ZN(new_n254));
  INV_X1    g0054(.A(KEYINPUT80), .ZN(new_n255));
  NAND2_X1  g0055(.A1(new_n255), .A2(G116), .ZN(new_n256));
  NAND2_X1  g0056(.A1(new_n254), .A2(new_n256), .ZN(new_n257));
  INV_X1    g0057(.A(G1), .ZN(new_n258));
  NAND3_X1  g0058(.A1(new_n258), .A2(G13), .A3(G20), .ZN(new_n259));
  OAI21_X1  g0059(.A(KEYINPUT82), .B1(new_n257), .B2(new_n259), .ZN(new_n260));
  XNOR2_X1  g0060(.A(KEYINPUT80), .B(G116), .ZN(new_n261));
  INV_X1    g0061(.A(new_n259), .ZN(new_n262));
  INV_X1    g0062(.A(KEYINPUT82), .ZN(new_n263));
  NAND3_X1  g0063(.A1(new_n261), .A2(new_n262), .A3(new_n263), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n260), .A2(new_n264), .ZN(new_n265));
  NAND3_X1  g0065(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n266));
  AND2_X1   g0066(.A1(new_n266), .A2(new_n216), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n258), .A2(G33), .ZN(new_n268));
  NAND3_X1  g0068(.A1(new_n267), .A2(new_n268), .A3(new_n259), .ZN(new_n269));
  OAI21_X1  g0069(.A(new_n265), .B1(new_n253), .B2(new_n269), .ZN(new_n270));
  AOI21_X1  g0070(.A(new_n267), .B1(G20), .B2(new_n261), .ZN(new_n271));
  INV_X1    g0071(.A(KEYINPUT83), .ZN(new_n272));
  NAND2_X1  g0072(.A1(G33), .A2(G283), .ZN(new_n273));
  OAI21_X1  g0073(.A(new_n273), .B1(new_n205), .B2(G33), .ZN(new_n274));
  INV_X1    g0074(.A(new_n274), .ZN(new_n275));
  AOI21_X1  g0075(.A(new_n272), .B1(new_n275), .B2(new_n215), .ZN(new_n276));
  OR2_X1    g0076(.A1(KEYINPUT64), .A2(G20), .ZN(new_n277));
  NAND2_X1  g0077(.A1(KEYINPUT64), .A2(G20), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n277), .A2(new_n278), .ZN(new_n279));
  NOR3_X1   g0079(.A1(new_n279), .A2(new_n274), .A3(KEYINPUT83), .ZN(new_n280));
  OAI21_X1  g0080(.A(new_n271), .B1(new_n276), .B2(new_n280), .ZN(new_n281));
  INV_X1    g0081(.A(KEYINPUT20), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n281), .A2(new_n282), .ZN(new_n283));
  NAND3_X1  g0083(.A1(new_n275), .A2(new_n272), .A3(new_n215), .ZN(new_n284));
  OAI21_X1  g0084(.A(KEYINPUT83), .B1(new_n279), .B2(new_n274), .ZN(new_n285));
  NAND2_X1  g0085(.A1(new_n284), .A2(new_n285), .ZN(new_n286));
  NAND3_X1  g0086(.A1(new_n286), .A2(KEYINPUT20), .A3(new_n271), .ZN(new_n287));
  AOI21_X1  g0087(.A(new_n270), .B1(new_n283), .B2(new_n287), .ZN(new_n288));
  AOI21_X1  g0088(.A(new_n216), .B1(G33), .B2(G41), .ZN(new_n289));
  INV_X1    g0089(.A(KEYINPUT3), .ZN(new_n290));
  INV_X1    g0090(.A(G33), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n290), .A2(new_n291), .ZN(new_n292));
  INV_X1    g0092(.A(G303), .ZN(new_n293));
  NAND2_X1  g0093(.A1(KEYINPUT3), .A2(G33), .ZN(new_n294));
  NAND3_X1  g0094(.A1(new_n292), .A2(new_n293), .A3(new_n294), .ZN(new_n295));
  MUX2_X1   g0095(.A(G257), .B(G264), .S(G1698), .Z(new_n296));
  AND2_X1   g0096(.A1(KEYINPUT3), .A2(G33), .ZN(new_n297));
  NOR2_X1   g0097(.A1(KEYINPUT3), .A2(G33), .ZN(new_n298));
  NOR2_X1   g0098(.A1(new_n297), .A2(new_n298), .ZN(new_n299));
  OAI211_X1 g0099(.A(new_n289), .B(new_n295), .C1(new_n296), .C2(new_n299), .ZN(new_n300));
  INV_X1    g0100(.A(G274), .ZN(new_n301));
  INV_X1    g0101(.A(new_n216), .ZN(new_n302));
  NAND2_X1  g0102(.A1(G33), .A2(G41), .ZN(new_n303));
  AOI21_X1  g0103(.A(new_n301), .B1(new_n302), .B2(new_n303), .ZN(new_n304));
  INV_X1    g0104(.A(G45), .ZN(new_n305));
  NOR2_X1   g0105(.A1(new_n305), .A2(G1), .ZN(new_n306));
  XNOR2_X1  g0106(.A(KEYINPUT5), .B(G41), .ZN(new_n307));
  NAND3_X1  g0107(.A1(new_n304), .A2(new_n306), .A3(new_n307), .ZN(new_n308));
  AND2_X1   g0108(.A1(KEYINPUT5), .A2(G41), .ZN(new_n309));
  NOR2_X1   g0109(.A1(KEYINPUT5), .A2(G41), .ZN(new_n310));
  OAI21_X1  g0110(.A(new_n306), .B1(new_n309), .B2(new_n310), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n302), .A2(new_n303), .ZN(new_n312));
  NAND3_X1  g0112(.A1(new_n311), .A2(G270), .A3(new_n312), .ZN(new_n313));
  NAND3_X1  g0113(.A1(new_n300), .A2(new_n308), .A3(new_n313), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n314), .A2(G169), .ZN(new_n315));
  OAI21_X1  g0115(.A(new_n252), .B1(new_n288), .B2(new_n315), .ZN(new_n316));
  INV_X1    g0116(.A(new_n270), .ZN(new_n317));
  INV_X1    g0117(.A(new_n287), .ZN(new_n318));
  AOI21_X1  g0118(.A(KEYINPUT20), .B1(new_n286), .B2(new_n271), .ZN(new_n319));
  OAI21_X1  g0119(.A(new_n317), .B1(new_n318), .B2(new_n319), .ZN(new_n320));
  INV_X1    g0120(.A(new_n315), .ZN(new_n321));
  NAND3_X1  g0121(.A1(new_n320), .A2(KEYINPUT21), .A3(new_n321), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n314), .A2(G200), .ZN(new_n323));
  INV_X1    g0123(.A(new_n314), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n324), .A2(G190), .ZN(new_n325));
  NAND3_X1  g0125(.A1(new_n288), .A2(new_n323), .A3(new_n325), .ZN(new_n326));
  NAND4_X1  g0126(.A1(new_n300), .A2(G179), .A3(new_n313), .A4(new_n308), .ZN(new_n327));
  INV_X1    g0127(.A(new_n327), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n320), .A2(new_n328), .ZN(new_n329));
  AND4_X1   g0129(.A1(new_n316), .A2(new_n322), .A3(new_n326), .A4(new_n329), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n266), .A2(new_n216), .ZN(new_n331));
  AOI21_X1  g0131(.A(new_n331), .B1(new_n258), .B2(G20), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n332), .A2(G50), .ZN(new_n333));
  OAI21_X1  g0133(.A(new_n333), .B1(G50), .B2(new_n259), .ZN(new_n334));
  INV_X1    g0134(.A(G20), .ZN(new_n335));
  NAND3_X1  g0135(.A1(new_n335), .A2(new_n291), .A3(KEYINPUT68), .ZN(new_n336));
  INV_X1    g0136(.A(KEYINPUT68), .ZN(new_n337));
  OAI21_X1  g0137(.A(new_n337), .B1(G20), .B2(G33), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n336), .A2(new_n338), .ZN(new_n339));
  AOI22_X1  g0139(.A1(new_n339), .A2(G150), .B1(G20), .B2(new_n203), .ZN(new_n340));
  XNOR2_X1  g0140(.A(KEYINPUT8), .B(G58), .ZN(new_n341));
  INV_X1    g0141(.A(KEYINPUT67), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n341), .A2(new_n342), .ZN(new_n343));
  INV_X1    g0143(.A(KEYINPUT8), .ZN(new_n344));
  NAND3_X1  g0144(.A1(new_n344), .A2(KEYINPUT67), .A3(G58), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n343), .A2(new_n345), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n215), .A2(G33), .ZN(new_n347));
  OAI21_X1  g0147(.A(new_n340), .B1(new_n346), .B2(new_n347), .ZN(new_n348));
  AOI21_X1  g0148(.A(new_n334), .B1(new_n331), .B2(new_n348), .ZN(new_n349));
  INV_X1    g0149(.A(G169), .ZN(new_n350));
  XNOR2_X1  g0150(.A(KEYINPUT3), .B(G33), .ZN(new_n351));
  INV_X1    g0151(.A(G1698), .ZN(new_n352));
  NAND3_X1  g0152(.A1(new_n351), .A2(G222), .A3(new_n352), .ZN(new_n353));
  NAND3_X1  g0153(.A1(new_n351), .A2(G223), .A3(G1698), .ZN(new_n354));
  INV_X1    g0154(.A(G77), .ZN(new_n355));
  OAI211_X1 g0155(.A(new_n353), .B(new_n354), .C1(new_n355), .C2(new_n351), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n356), .A2(new_n289), .ZN(new_n357));
  INV_X1    g0157(.A(G41), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n358), .A2(new_n305), .ZN(new_n359));
  AOI22_X1  g0159(.A1(new_n258), .A2(new_n359), .B1(new_n302), .B2(new_n303), .ZN(new_n360));
  OAI21_X1  g0160(.A(new_n258), .B1(G41), .B2(G45), .ZN(new_n361));
  INV_X1    g0161(.A(new_n361), .ZN(new_n362));
  AOI22_X1  g0162(.A1(new_n360), .A2(G226), .B1(new_n304), .B2(new_n362), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n357), .A2(new_n363), .ZN(new_n364));
  AOI21_X1  g0164(.A(new_n349), .B1(new_n350), .B2(new_n364), .ZN(new_n365));
  XOR2_X1   g0165(.A(KEYINPUT69), .B(G179), .Z(new_n366));
  INV_X1    g0166(.A(new_n366), .ZN(new_n367));
  OAI21_X1  g0167(.A(new_n365), .B1(new_n367), .B2(new_n364), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n349), .A2(KEYINPUT9), .ZN(new_n369));
  INV_X1    g0169(.A(G190), .ZN(new_n370));
  OAI21_X1  g0170(.A(new_n369), .B1(new_n370), .B2(new_n364), .ZN(new_n371));
  NOR2_X1   g0171(.A1(new_n371), .A2(KEYINPUT10), .ZN(new_n372));
  OR3_X1    g0172(.A1(new_n349), .A2(KEYINPUT72), .A3(KEYINPUT9), .ZN(new_n373));
  OAI21_X1  g0173(.A(KEYINPUT72), .B1(new_n349), .B2(KEYINPUT9), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n373), .A2(new_n374), .ZN(new_n375));
  INV_X1    g0175(.A(G200), .ZN(new_n376));
  AOI21_X1  g0176(.A(new_n376), .B1(new_n357), .B2(new_n363), .ZN(new_n377));
  XNOR2_X1  g0177(.A(new_n377), .B(KEYINPUT73), .ZN(new_n378));
  AND3_X1   g0178(.A1(new_n372), .A2(new_n375), .A3(new_n378), .ZN(new_n379));
  INV_X1    g0179(.A(KEYINPUT10), .ZN(new_n380));
  NOR2_X1   g0180(.A1(new_n371), .A2(new_n377), .ZN(new_n381));
  AOI21_X1  g0181(.A(new_n380), .B1(new_n381), .B2(new_n375), .ZN(new_n382));
  OAI21_X1  g0182(.A(new_n368), .B1(new_n379), .B2(new_n382), .ZN(new_n383));
  INV_X1    g0183(.A(KEYINPUT74), .ZN(new_n384));
  NAND2_X1  g0184(.A1(new_n238), .A2(G1698), .ZN(new_n385));
  OAI211_X1 g0185(.A(new_n351), .B(new_n385), .C1(G226), .C2(G1698), .ZN(new_n386));
  NAND2_X1  g0186(.A1(G33), .A2(G97), .ZN(new_n387));
  AOI21_X1  g0187(.A(new_n312), .B1(new_n386), .B2(new_n387), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n304), .A2(new_n362), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n312), .A2(new_n361), .ZN(new_n390));
  OAI21_X1  g0190(.A(new_n389), .B1(new_n390), .B2(new_n223), .ZN(new_n391));
  OAI21_X1  g0191(.A(KEYINPUT13), .B1(new_n388), .B2(new_n391), .ZN(new_n392));
  INV_X1    g0192(.A(new_n392), .ZN(new_n393));
  NOR3_X1   g0193(.A1(new_n388), .A2(new_n391), .A3(KEYINPUT13), .ZN(new_n394));
  NOR2_X1   g0194(.A1(new_n393), .A2(new_n394), .ZN(new_n395));
  OAI21_X1  g0195(.A(new_n384), .B1(new_n395), .B2(new_n376), .ZN(new_n396));
  OAI211_X1 g0196(.A(KEYINPUT74), .B(G200), .C1(new_n393), .C2(new_n394), .ZN(new_n397));
  NAND2_X1  g0197(.A1(new_n396), .A2(new_n397), .ZN(new_n398));
  AOI22_X1  g0198(.A1(new_n339), .A2(G50), .B1(new_n222), .B2(G20), .ZN(new_n399));
  OAI21_X1  g0199(.A(new_n399), .B1(new_n355), .B2(new_n347), .ZN(new_n400));
  AND3_X1   g0200(.A1(new_n400), .A2(KEYINPUT11), .A3(new_n331), .ZN(new_n401));
  AOI21_X1  g0201(.A(KEYINPUT11), .B1(new_n400), .B2(new_n331), .ZN(new_n402));
  NOR2_X1   g0202(.A1(new_n401), .A2(new_n402), .ZN(new_n403));
  INV_X1    g0203(.A(KEYINPUT12), .ZN(new_n404));
  AOI21_X1  g0204(.A(new_n404), .B1(new_n222), .B2(new_n262), .ZN(new_n405));
  INV_X1    g0205(.A(KEYINPUT75), .ZN(new_n406));
  AND2_X1   g0206(.A1(new_n405), .A2(new_n406), .ZN(new_n407));
  INV_X1    g0207(.A(G68), .ZN(new_n408));
  NAND3_X1  g0208(.A1(new_n262), .A2(new_n404), .A3(new_n408), .ZN(new_n409));
  OAI21_X1  g0209(.A(new_n409), .B1(new_n405), .B2(new_n406), .ZN(new_n410));
  INV_X1    g0210(.A(new_n332), .ZN(new_n411));
  OAI22_X1  g0211(.A1(new_n407), .A2(new_n410), .B1(new_n408), .B2(new_n411), .ZN(new_n412));
  INV_X1    g0212(.A(KEYINPUT76), .ZN(new_n413));
  NAND2_X1  g0213(.A1(new_n412), .A2(new_n413), .ZN(new_n414));
  OAI221_X1 g0214(.A(KEYINPUT76), .B1(new_n408), .B2(new_n411), .C1(new_n407), .C2(new_n410), .ZN(new_n415));
  AND3_X1   g0215(.A1(new_n403), .A2(new_n414), .A3(new_n415), .ZN(new_n416));
  INV_X1    g0216(.A(new_n388), .ZN(new_n417));
  INV_X1    g0217(.A(new_n391), .ZN(new_n418));
  INV_X1    g0218(.A(KEYINPUT13), .ZN(new_n419));
  NAND3_X1  g0219(.A1(new_n417), .A2(new_n418), .A3(new_n419), .ZN(new_n420));
  NAND3_X1  g0220(.A1(new_n420), .A2(G190), .A3(new_n392), .ZN(new_n421));
  NAND3_X1  g0221(.A1(new_n398), .A2(new_n416), .A3(new_n421), .ZN(new_n422));
  INV_X1    g0222(.A(new_n416), .ZN(new_n423));
  AOI21_X1  g0223(.A(new_n350), .B1(new_n420), .B2(new_n392), .ZN(new_n424));
  INV_X1    g0224(.A(KEYINPUT14), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n424), .A2(new_n425), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n395), .A2(G179), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n426), .A2(new_n427), .ZN(new_n428));
  NOR2_X1   g0228(.A1(new_n424), .A2(new_n425), .ZN(new_n429));
  OAI21_X1  g0229(.A(new_n423), .B1(new_n428), .B2(new_n429), .ZN(new_n430));
  XNOR2_X1  g0230(.A(KEYINPUT15), .B(G87), .ZN(new_n431));
  INV_X1    g0231(.A(new_n431), .ZN(new_n432));
  NAND3_X1  g0232(.A1(new_n432), .A2(G33), .A3(new_n215), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n344), .A2(G58), .ZN(new_n434));
  INV_X1    g0234(.A(G58), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n435), .A2(KEYINPUT8), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n434), .A2(new_n436), .ZN(new_n437));
  AOI22_X1  g0237(.A1(new_n339), .A2(new_n437), .B1(new_n279), .B2(G77), .ZN(new_n438));
  INV_X1    g0238(.A(KEYINPUT70), .ZN(new_n439));
  OAI21_X1  g0239(.A(new_n433), .B1(new_n438), .B2(new_n439), .ZN(new_n440));
  NAND2_X1  g0240(.A1(new_n339), .A2(new_n437), .ZN(new_n441));
  NAND2_X1  g0241(.A1(new_n279), .A2(G77), .ZN(new_n442));
  AND3_X1   g0242(.A1(new_n441), .A2(new_n439), .A3(new_n442), .ZN(new_n443));
  OAI21_X1  g0243(.A(new_n331), .B1(new_n440), .B2(new_n443), .ZN(new_n444));
  OAI211_X1 g0244(.A(G232), .B(new_n352), .C1(new_n297), .C2(new_n298), .ZN(new_n445));
  OAI211_X1 g0245(.A(G238), .B(G1698), .C1(new_n297), .C2(new_n298), .ZN(new_n446));
  NAND3_X1  g0246(.A1(new_n292), .A2(G107), .A3(new_n294), .ZN(new_n447));
  NAND3_X1  g0247(.A1(new_n445), .A2(new_n446), .A3(new_n447), .ZN(new_n448));
  NAND2_X1  g0248(.A1(new_n448), .A2(new_n289), .ZN(new_n449));
  AOI22_X1  g0249(.A1(new_n360), .A2(G244), .B1(new_n304), .B2(new_n362), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n449), .A2(new_n450), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n451), .A2(G200), .ZN(new_n452));
  NOR2_X1   g0252(.A1(new_n259), .A2(G77), .ZN(new_n453));
  AOI21_X1  g0253(.A(new_n453), .B1(new_n332), .B2(G77), .ZN(new_n454));
  NAND3_X1  g0254(.A1(new_n444), .A2(new_n452), .A3(new_n454), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n455), .A2(KEYINPUT71), .ZN(new_n456));
  INV_X1    g0256(.A(KEYINPUT71), .ZN(new_n457));
  NAND4_X1  g0257(.A1(new_n444), .A2(new_n452), .A3(new_n457), .A4(new_n454), .ZN(new_n458));
  NOR2_X1   g0258(.A1(new_n451), .A2(new_n370), .ZN(new_n459));
  INV_X1    g0259(.A(new_n459), .ZN(new_n460));
  NAND3_X1  g0260(.A1(new_n456), .A2(new_n458), .A3(new_n460), .ZN(new_n461));
  NAND2_X1  g0261(.A1(new_n444), .A2(new_n454), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n451), .A2(new_n350), .ZN(new_n463));
  NAND3_X1  g0263(.A1(new_n449), .A2(new_n366), .A3(new_n450), .ZN(new_n464));
  NAND3_X1  g0264(.A1(new_n462), .A2(new_n463), .A3(new_n464), .ZN(new_n465));
  NAND4_X1  g0265(.A1(new_n422), .A2(new_n430), .A3(new_n461), .A4(new_n465), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n346), .A2(new_n259), .ZN(new_n467));
  OAI21_X1  g0267(.A(new_n467), .B1(new_n332), .B2(new_n346), .ZN(new_n468));
  OAI21_X1  g0268(.A(new_n218), .B1(new_n222), .B2(new_n435), .ZN(new_n469));
  AOI22_X1  g0269(.A1(new_n469), .A2(G20), .B1(G159), .B2(new_n339), .ZN(new_n470));
  INV_X1    g0270(.A(KEYINPUT77), .ZN(new_n471));
  OAI21_X1  g0271(.A(new_n471), .B1(new_n297), .B2(new_n298), .ZN(new_n472));
  NAND3_X1  g0272(.A1(new_n292), .A2(KEYINPUT77), .A3(new_n294), .ZN(new_n473));
  INV_X1    g0273(.A(KEYINPUT7), .ZN(new_n474));
  NAND4_X1  g0274(.A1(new_n472), .A2(new_n473), .A3(new_n474), .A4(new_n215), .ZN(new_n475));
  NAND3_X1  g0275(.A1(new_n292), .A2(new_n335), .A3(new_n294), .ZN(new_n476));
  AOI21_X1  g0276(.A(new_n408), .B1(new_n476), .B2(KEYINPUT7), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n475), .A2(new_n477), .ZN(new_n478));
  NAND3_X1  g0278(.A1(new_n470), .A2(new_n478), .A3(KEYINPUT16), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n479), .A2(new_n331), .ZN(new_n480));
  NAND3_X1  g0280(.A1(new_n215), .A2(new_n299), .A3(KEYINPUT7), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n476), .A2(new_n474), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n481), .A2(new_n482), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n408), .A2(KEYINPUT65), .ZN(new_n484));
  INV_X1    g0284(.A(KEYINPUT65), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n485), .A2(G68), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n484), .A2(new_n486), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n483), .A2(new_n487), .ZN(new_n488));
  AOI21_X1  g0288(.A(KEYINPUT16), .B1(new_n488), .B2(new_n470), .ZN(new_n489));
  OAI21_X1  g0289(.A(new_n468), .B1(new_n480), .B2(new_n489), .ZN(new_n490));
  OAI211_X1 g0290(.A(G223), .B(new_n352), .C1(new_n297), .C2(new_n298), .ZN(new_n491));
  INV_X1    g0291(.A(KEYINPUT78), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n491), .A2(new_n492), .ZN(new_n493));
  NAND4_X1  g0293(.A1(new_n351), .A2(KEYINPUT78), .A3(G223), .A4(new_n352), .ZN(new_n494));
  NAND3_X1  g0294(.A1(new_n351), .A2(G226), .A3(G1698), .ZN(new_n495));
  NAND2_X1  g0295(.A1(G33), .A2(G87), .ZN(new_n496));
  XNOR2_X1  g0296(.A(new_n496), .B(KEYINPUT79), .ZN(new_n497));
  NAND4_X1  g0297(.A1(new_n493), .A2(new_n494), .A3(new_n495), .A4(new_n497), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n498), .A2(new_n289), .ZN(new_n499));
  OAI21_X1  g0299(.A(new_n389), .B1(new_n390), .B2(new_n238), .ZN(new_n500));
  INV_X1    g0300(.A(new_n500), .ZN(new_n501));
  NAND3_X1  g0301(.A1(new_n499), .A2(new_n367), .A3(new_n501), .ZN(new_n502));
  AOI21_X1  g0302(.A(new_n500), .B1(new_n498), .B2(new_n289), .ZN(new_n503));
  OAI21_X1  g0303(.A(new_n502), .B1(new_n350), .B2(new_n503), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n490), .A2(new_n504), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n505), .A2(KEYINPUT18), .ZN(new_n506));
  INV_X1    g0306(.A(KEYINPUT16), .ZN(new_n507));
  AOI21_X1  g0307(.A(new_n201), .B1(new_n487), .B2(G58), .ZN(new_n508));
  INV_X1    g0308(.A(G159), .ZN(new_n509));
  AND2_X1   g0309(.A1(new_n336), .A2(new_n338), .ZN(new_n510));
  OAI22_X1  g0310(.A1(new_n508), .A2(new_n335), .B1(new_n509), .B2(new_n510), .ZN(new_n511));
  AOI21_X1  g0311(.A(new_n222), .B1(new_n481), .B2(new_n482), .ZN(new_n512));
  OAI21_X1  g0312(.A(new_n507), .B1(new_n511), .B2(new_n512), .ZN(new_n513));
  NAND3_X1  g0313(.A1(new_n513), .A2(new_n331), .A3(new_n479), .ZN(new_n514));
  AND2_X1   g0314(.A1(new_n514), .A2(new_n468), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n503), .A2(new_n370), .ZN(new_n516));
  OAI21_X1  g0316(.A(new_n516), .B1(G200), .B2(new_n503), .ZN(new_n517));
  NAND3_X1  g0317(.A1(new_n515), .A2(KEYINPUT17), .A3(new_n517), .ZN(new_n518));
  AOI211_X1 g0318(.A(G190), .B(new_n500), .C1(new_n498), .C2(new_n289), .ZN(new_n519));
  AOI21_X1  g0319(.A(G200), .B1(new_n499), .B2(new_n501), .ZN(new_n520));
  OAI211_X1 g0320(.A(new_n514), .B(new_n468), .C1(new_n519), .C2(new_n520), .ZN(new_n521));
  INV_X1    g0321(.A(KEYINPUT17), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  INV_X1    g0323(.A(KEYINPUT18), .ZN(new_n524));
  NAND3_X1  g0324(.A1(new_n490), .A2(new_n504), .A3(new_n524), .ZN(new_n525));
  NAND4_X1  g0325(.A1(new_n506), .A2(new_n518), .A3(new_n523), .A4(new_n525), .ZN(new_n526));
  NOR3_X1   g0326(.A1(new_n383), .A2(new_n466), .A3(new_n526), .ZN(new_n527));
  OAI211_X1 g0327(.A(G257), .B(G1698), .C1(new_n297), .C2(new_n298), .ZN(new_n528));
  INV_X1    g0328(.A(KEYINPUT84), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  NAND4_X1  g0330(.A1(new_n351), .A2(KEYINPUT84), .A3(G257), .A4(G1698), .ZN(new_n531));
  NAND3_X1  g0331(.A1(new_n351), .A2(G250), .A3(new_n352), .ZN(new_n532));
  NAND2_X1  g0332(.A1(G33), .A2(G294), .ZN(new_n533));
  NAND4_X1  g0333(.A1(new_n530), .A2(new_n531), .A3(new_n532), .A4(new_n533), .ZN(new_n534));
  NAND2_X1  g0334(.A1(new_n534), .A2(new_n289), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n311), .A2(new_n312), .ZN(new_n536));
  INV_X1    g0336(.A(new_n536), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n537), .A2(G264), .ZN(new_n538));
  NAND3_X1  g0338(.A1(new_n535), .A2(new_n308), .A3(new_n538), .ZN(new_n539));
  NOR2_X1   g0339(.A1(new_n539), .A2(G179), .ZN(new_n540));
  OAI211_X1 g0340(.A(new_n277), .B(new_n278), .C1(new_n297), .C2(new_n298), .ZN(new_n541));
  INV_X1    g0341(.A(G87), .ZN(new_n542));
  OAI21_X1  g0342(.A(KEYINPUT22), .B1(new_n541), .B2(new_n542), .ZN(new_n543));
  INV_X1    g0343(.A(KEYINPUT22), .ZN(new_n544));
  NAND4_X1  g0344(.A1(new_n215), .A2(new_n351), .A3(new_n544), .A4(G87), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n543), .A2(new_n545), .ZN(new_n546));
  INV_X1    g0346(.A(KEYINPUT24), .ZN(new_n547));
  NOR3_X1   g0347(.A1(new_n261), .A2(G20), .A3(new_n291), .ZN(new_n548));
  OAI21_X1  g0348(.A(KEYINPUT23), .B1(new_n335), .B2(G107), .ZN(new_n549));
  OR2_X1    g0349(.A1(KEYINPUT23), .A2(G107), .ZN(new_n550));
  OAI21_X1  g0350(.A(new_n549), .B1(new_n215), .B2(new_n550), .ZN(new_n551));
  NOR2_X1   g0351(.A1(new_n548), .A2(new_n551), .ZN(new_n552));
  NAND3_X1  g0352(.A1(new_n546), .A2(new_n547), .A3(new_n552), .ZN(new_n553));
  INV_X1    g0353(.A(new_n553), .ZN(new_n554));
  AOI21_X1  g0354(.A(new_n547), .B1(new_n546), .B2(new_n552), .ZN(new_n555));
  OAI21_X1  g0355(.A(new_n331), .B1(new_n554), .B2(new_n555), .ZN(new_n556));
  INV_X1    g0356(.A(KEYINPUT25), .ZN(new_n557));
  OAI21_X1  g0357(.A(new_n557), .B1(new_n259), .B2(G107), .ZN(new_n558));
  INV_X1    g0358(.A(new_n558), .ZN(new_n559));
  NOR3_X1   g0359(.A1(new_n259), .A2(new_n557), .A3(G107), .ZN(new_n560));
  OAI22_X1  g0360(.A1(new_n269), .A2(new_n206), .B1(new_n559), .B2(new_n560), .ZN(new_n561));
  INV_X1    g0361(.A(new_n561), .ZN(new_n562));
  AOI21_X1  g0362(.A(new_n540), .B1(new_n556), .B2(new_n562), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n539), .A2(new_n350), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n539), .A2(new_n376), .ZN(new_n565));
  OAI21_X1  g0365(.A(new_n565), .B1(G190), .B2(new_n539), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n546), .A2(new_n552), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n567), .A2(KEYINPUT24), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n568), .A2(new_n553), .ZN(new_n569));
  AOI21_X1  g0369(.A(new_n561), .B1(new_n569), .B2(new_n331), .ZN(new_n570));
  AOI22_X1  g0370(.A1(new_n563), .A2(new_n564), .B1(new_n566), .B2(new_n570), .ZN(new_n571));
  INV_X1    g0371(.A(G257), .ZN(new_n572));
  OAI21_X1  g0372(.A(new_n308), .B1(new_n536), .B2(new_n572), .ZN(new_n573));
  OAI211_X1 g0373(.A(G244), .B(new_n352), .C1(new_n297), .C2(new_n298), .ZN(new_n574));
  INV_X1    g0374(.A(KEYINPUT4), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  NAND4_X1  g0376(.A1(new_n351), .A2(KEYINPUT4), .A3(G244), .A4(new_n352), .ZN(new_n577));
  NAND3_X1  g0377(.A1(new_n351), .A2(G250), .A3(G1698), .ZN(new_n578));
  NAND4_X1  g0378(.A1(new_n576), .A2(new_n577), .A3(new_n273), .A4(new_n578), .ZN(new_n579));
  AOI21_X1  g0379(.A(new_n573), .B1(new_n579), .B2(new_n289), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n580), .A2(new_n366), .ZN(new_n581));
  NAND2_X1  g0381(.A1(G97), .A2(G107), .ZN(new_n582));
  AOI21_X1  g0382(.A(KEYINPUT6), .B1(new_n207), .B2(new_n582), .ZN(new_n583));
  INV_X1    g0383(.A(KEYINPUT6), .ZN(new_n584));
  NOR2_X1   g0384(.A1(new_n246), .A2(new_n584), .ZN(new_n585));
  NOR2_X1   g0385(.A1(new_n583), .A2(new_n585), .ZN(new_n586));
  OAI22_X1  g0386(.A1(new_n586), .A2(new_n215), .B1(new_n355), .B2(new_n510), .ZN(new_n587));
  AOI21_X1  g0387(.A(new_n206), .B1(new_n481), .B2(new_n482), .ZN(new_n588));
  OAI21_X1  g0388(.A(new_n331), .B1(new_n587), .B2(new_n588), .ZN(new_n589));
  NOR2_X1   g0389(.A1(new_n259), .A2(G97), .ZN(new_n590));
  INV_X1    g0390(.A(new_n269), .ZN(new_n591));
  AOI21_X1  g0391(.A(new_n590), .B1(new_n591), .B2(G97), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n589), .A2(new_n592), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n581), .A2(new_n593), .ZN(new_n594));
  NOR2_X1   g0394(.A1(new_n580), .A2(G169), .ZN(new_n595));
  OAI211_X1 g0395(.A(new_n589), .B(new_n592), .C1(new_n580), .C2(new_n376), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n579), .A2(new_n289), .ZN(new_n597));
  INV_X1    g0397(.A(new_n573), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n597), .A2(new_n598), .ZN(new_n599));
  NOR2_X1   g0399(.A1(new_n599), .A2(new_n370), .ZN(new_n600));
  OAI22_X1  g0400(.A1(new_n594), .A2(new_n595), .B1(new_n596), .B2(new_n600), .ZN(new_n601));
  NOR2_X1   g0401(.A1(new_n432), .A2(new_n259), .ZN(new_n602));
  NAND4_X1  g0402(.A1(new_n277), .A2(G33), .A3(G97), .A4(new_n278), .ZN(new_n603));
  INV_X1    g0403(.A(KEYINPUT19), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  NAND3_X1  g0405(.A1(KEYINPUT19), .A2(G33), .A3(G97), .ZN(new_n606));
  NAND3_X1  g0406(.A1(new_n277), .A2(new_n278), .A3(new_n606), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n542), .A2(KEYINPUT81), .ZN(new_n608));
  INV_X1    g0408(.A(KEYINPUT81), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n609), .A2(G87), .ZN(new_n610));
  NOR2_X1   g0410(.A1(G97), .A2(G107), .ZN(new_n611));
  NAND3_X1  g0411(.A1(new_n608), .A2(new_n610), .A3(new_n611), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n607), .A2(new_n612), .ZN(new_n613));
  NAND3_X1  g0413(.A1(new_n215), .A2(new_n351), .A3(G68), .ZN(new_n614));
  NAND3_X1  g0414(.A1(new_n605), .A2(new_n613), .A3(new_n614), .ZN(new_n615));
  AOI21_X1  g0415(.A(new_n602), .B1(new_n615), .B2(new_n331), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n591), .A2(new_n432), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n257), .A2(G33), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n223), .A2(new_n352), .ZN(new_n619));
  INV_X1    g0419(.A(G244), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n620), .A2(G1698), .ZN(new_n621));
  OAI211_X1 g0421(.A(new_n619), .B(new_n621), .C1(new_n297), .C2(new_n298), .ZN(new_n622));
  AOI21_X1  g0422(.A(new_n312), .B1(new_n618), .B2(new_n622), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n304), .A2(new_n306), .ZN(new_n624));
  INV_X1    g0424(.A(G250), .ZN(new_n625));
  AOI21_X1  g0425(.A(new_n625), .B1(new_n258), .B2(G45), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n312), .A2(new_n626), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n624), .A2(new_n627), .ZN(new_n628));
  NOR2_X1   g0428(.A1(new_n623), .A2(new_n628), .ZN(new_n629));
  AOI22_X1  g0429(.A1(new_n616), .A2(new_n617), .B1(new_n629), .B2(new_n366), .ZN(new_n630));
  OAI21_X1  g0430(.A(new_n630), .B1(G169), .B2(new_n629), .ZN(new_n631));
  AND4_X1   g0431(.A1(G87), .A2(new_n267), .A3(new_n268), .A4(new_n259), .ZN(new_n632));
  AOI211_X1 g0432(.A(new_n602), .B(new_n632), .C1(new_n615), .C2(new_n331), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n629), .A2(G190), .ZN(new_n634));
  OAI211_X1 g0434(.A(new_n633), .B(new_n634), .C1(new_n376), .C2(new_n629), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n631), .A2(new_n635), .ZN(new_n636));
  NOR2_X1   g0436(.A1(new_n601), .A2(new_n636), .ZN(new_n637));
  AND4_X1   g0437(.A1(new_n330), .A2(new_n527), .A3(new_n571), .A4(new_n637), .ZN(G372));
  INV_X1    g0438(.A(new_n368), .ZN(new_n639));
  NOR2_X1   g0439(.A1(new_n379), .A2(new_n382), .ZN(new_n640));
  NAND4_X1  g0440(.A1(new_n403), .A2(new_n421), .A3(new_n414), .A4(new_n415), .ZN(new_n641));
  AOI21_X1  g0441(.A(new_n641), .B1(new_n396), .B2(new_n397), .ZN(new_n642));
  OAI21_X1  g0442(.A(new_n430), .B1(new_n642), .B2(new_n465), .ZN(new_n643));
  AND2_X1   g0443(.A1(new_n518), .A2(new_n523), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  AND2_X1   g0445(.A1(new_n506), .A2(new_n525), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  AOI21_X1  g0447(.A(new_n640), .B1(new_n647), .B2(KEYINPUT88), .ZN(new_n648));
  INV_X1    g0448(.A(KEYINPUT88), .ZN(new_n649));
  NAND3_X1  g0449(.A1(new_n645), .A2(new_n649), .A3(new_n646), .ZN(new_n650));
  AOI21_X1  g0450(.A(new_n639), .B1(new_n648), .B2(new_n650), .ZN(new_n651));
  INV_X1    g0451(.A(new_n651), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n283), .A2(new_n287), .ZN(new_n653));
  AOI21_X1  g0453(.A(new_n315), .B1(new_n653), .B2(new_n317), .ZN(new_n654));
  AOI22_X1  g0454(.A1(new_n654), .A2(KEYINPUT21), .B1(new_n320), .B2(new_n328), .ZN(new_n655));
  AOI22_X1  g0455(.A1(new_n534), .A2(new_n289), .B1(G264), .B2(new_n537), .ZN(new_n656));
  INV_X1    g0456(.A(G179), .ZN(new_n657));
  NAND3_X1  g0457(.A1(new_n656), .A2(new_n657), .A3(new_n308), .ZN(new_n658));
  AOI21_X1  g0458(.A(new_n267), .B1(new_n568), .B2(new_n553), .ZN(new_n659));
  OAI211_X1 g0459(.A(new_n564), .B(new_n658), .C1(new_n659), .C2(new_n561), .ZN(new_n660));
  NAND3_X1  g0460(.A1(new_n655), .A2(new_n660), .A3(new_n316), .ZN(new_n661));
  NOR2_X1   g0461(.A1(G238), .A2(G1698), .ZN(new_n662));
  AOI21_X1  g0462(.A(new_n662), .B1(new_n620), .B2(G1698), .ZN(new_n663));
  AOI22_X1  g0463(.A1(new_n663), .A2(new_n351), .B1(new_n257), .B2(G33), .ZN(new_n664));
  OAI21_X1  g0464(.A(KEYINPUT85), .B1(new_n664), .B2(new_n312), .ZN(new_n665));
  INV_X1    g0465(.A(KEYINPUT85), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n623), .A2(new_n666), .ZN(new_n667));
  AOI21_X1  g0467(.A(new_n628), .B1(new_n665), .B2(new_n667), .ZN(new_n668));
  OAI211_X1 g0468(.A(new_n633), .B(new_n634), .C1(new_n668), .C2(new_n376), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n629), .A2(new_n366), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n615), .A2(new_n331), .ZN(new_n671));
  INV_X1    g0471(.A(new_n602), .ZN(new_n672));
  NAND3_X1  g0472(.A1(new_n671), .A2(new_n672), .A3(new_n617), .ZN(new_n673));
  OAI211_X1 g0473(.A(new_n670), .B(new_n673), .C1(new_n668), .C2(G169), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n669), .A2(new_n674), .ZN(new_n675));
  AOI21_X1  g0475(.A(new_n675), .B1(new_n570), .B2(new_n566), .ZN(new_n676));
  INV_X1    g0476(.A(new_n601), .ZN(new_n677));
  NAND3_X1  g0477(.A1(new_n661), .A2(new_n676), .A3(new_n677), .ZN(new_n678));
  INV_X1    g0478(.A(new_n674), .ZN(new_n679));
  INV_X1    g0479(.A(KEYINPUT26), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n599), .A2(new_n350), .ZN(new_n681));
  NAND3_X1  g0481(.A1(new_n681), .A2(new_n593), .A3(new_n581), .ZN(new_n682));
  OAI21_X1  g0482(.A(new_n680), .B1(new_n675), .B2(new_n682), .ZN(new_n683));
  AND3_X1   g0483(.A1(new_n681), .A2(new_n593), .A3(new_n581), .ZN(new_n684));
  XNOR2_X1  g0484(.A(KEYINPUT86), .B(KEYINPUT26), .ZN(new_n685));
  INV_X1    g0485(.A(new_n685), .ZN(new_n686));
  NAND4_X1  g0486(.A1(new_n684), .A2(new_n631), .A3(new_n635), .A4(new_n686), .ZN(new_n687));
  AOI21_X1  g0487(.A(new_n679), .B1(new_n683), .B2(new_n687), .ZN(new_n688));
  OAI21_X1  g0488(.A(new_n678), .B1(new_n688), .B2(KEYINPUT87), .ZN(new_n689));
  INV_X1    g0489(.A(new_n689), .ZN(new_n690));
  INV_X1    g0490(.A(KEYINPUT87), .ZN(new_n691));
  AOI211_X1 g0491(.A(new_n691), .B(new_n679), .C1(new_n683), .C2(new_n687), .ZN(new_n692));
  INV_X1    g0492(.A(new_n692), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n690), .A2(new_n693), .ZN(new_n694));
  AOI21_X1  g0494(.A(new_n652), .B1(new_n527), .B2(new_n694), .ZN(new_n695));
  XOR2_X1   g0495(.A(new_n695), .B(KEYINPUT89), .Z(G369));
  NAND2_X1  g0496(.A1(new_n570), .A2(new_n566), .ZN(new_n697));
  INV_X1    g0497(.A(G213), .ZN(new_n698));
  NAND2_X1  g0498(.A1(new_n258), .A2(G13), .ZN(new_n699));
  NOR3_X1   g0499(.A1(new_n279), .A2(KEYINPUT27), .A3(new_n699), .ZN(new_n700));
  OR2_X1    g0500(.A1(new_n700), .A2(KEYINPUT90), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n700), .A2(KEYINPUT90), .ZN(new_n702));
  AOI21_X1  g0502(.A(new_n698), .B1(new_n701), .B2(new_n702), .ZN(new_n703));
  OAI21_X1  g0503(.A(KEYINPUT27), .B1(new_n279), .B2(new_n699), .ZN(new_n704));
  XNOR2_X1  g0504(.A(new_n704), .B(KEYINPUT91), .ZN(new_n705));
  AND3_X1   g0505(.A1(new_n703), .A2(G343), .A3(new_n705), .ZN(new_n706));
  INV_X1    g0506(.A(new_n706), .ZN(new_n707));
  OAI211_X1 g0507(.A(new_n697), .B(new_n660), .C1(new_n570), .C2(new_n707), .ZN(new_n708));
  NAND3_X1  g0508(.A1(new_n563), .A2(new_n564), .A3(new_n706), .ZN(new_n709));
  NAND2_X1  g0509(.A1(new_n708), .A2(new_n709), .ZN(new_n710));
  INV_X1    g0510(.A(KEYINPUT92), .ZN(new_n711));
  OAI21_X1  g0511(.A(new_n330), .B1(new_n288), .B2(new_n707), .ZN(new_n712));
  NAND3_X1  g0512(.A1(new_n316), .A2(new_n322), .A3(new_n329), .ZN(new_n713));
  NAND3_X1  g0513(.A1(new_n713), .A2(new_n320), .A3(new_n706), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n712), .A2(new_n714), .ZN(new_n715));
  AOI21_X1  g0515(.A(new_n711), .B1(new_n715), .B2(G330), .ZN(new_n716));
  INV_X1    g0516(.A(G330), .ZN(new_n717));
  AOI211_X1 g0517(.A(KEYINPUT92), .B(new_n717), .C1(new_n712), .C2(new_n714), .ZN(new_n718));
  OAI21_X1  g0518(.A(new_n710), .B1(new_n716), .B2(new_n718), .ZN(new_n719));
  NAND4_X1  g0519(.A1(new_n713), .A2(new_n697), .A3(new_n660), .A4(new_n707), .ZN(new_n720));
  NAND3_X1  g0520(.A1(new_n563), .A2(new_n564), .A3(new_n707), .ZN(new_n721));
  NAND2_X1  g0521(.A1(new_n720), .A2(new_n721), .ZN(new_n722));
  INV_X1    g0522(.A(new_n722), .ZN(new_n723));
  NAND2_X1  g0523(.A1(new_n719), .A2(new_n723), .ZN(G399));
  NOR2_X1   g0524(.A1(new_n612), .A2(G116), .ZN(new_n725));
  XOR2_X1   g0525(.A(new_n725), .B(KEYINPUT93), .Z(new_n726));
  INV_X1    g0526(.A(new_n210), .ZN(new_n727));
  NOR2_X1   g0527(.A1(new_n727), .A2(G41), .ZN(new_n728));
  NOR3_X1   g0528(.A1(new_n726), .A2(new_n258), .A3(new_n728), .ZN(new_n729));
  AOI21_X1  g0529(.A(new_n729), .B1(new_n220), .B2(new_n728), .ZN(new_n730));
  XOR2_X1   g0530(.A(new_n730), .B(KEYINPUT28), .Z(new_n731));
  OAI21_X1  g0531(.A(new_n685), .B1(new_n636), .B2(new_n682), .ZN(new_n732));
  NAND2_X1  g0532(.A1(new_n732), .A2(KEYINPUT96), .ZN(new_n733));
  INV_X1    g0533(.A(new_n675), .ZN(new_n734));
  NAND3_X1  g0534(.A1(new_n734), .A2(KEYINPUT26), .A3(new_n684), .ZN(new_n735));
  INV_X1    g0535(.A(KEYINPUT96), .ZN(new_n736));
  OAI211_X1 g0536(.A(new_n736), .B(new_n685), .C1(new_n636), .C2(new_n682), .ZN(new_n737));
  NAND3_X1  g0537(.A1(new_n733), .A2(new_n735), .A3(new_n737), .ZN(new_n738));
  NAND3_X1  g0538(.A1(new_n738), .A2(new_n674), .A3(new_n678), .ZN(new_n739));
  NAND3_X1  g0539(.A1(new_n739), .A2(KEYINPUT29), .A3(new_n707), .ZN(new_n740));
  AOI21_X1  g0540(.A(new_n706), .B1(new_n690), .B2(new_n693), .ZN(new_n741));
  XOR2_X1   g0541(.A(KEYINPUT95), .B(KEYINPUT29), .Z(new_n742));
  INV_X1    g0542(.A(new_n742), .ZN(new_n743));
  OAI21_X1  g0543(.A(new_n740), .B1(new_n741), .B2(new_n743), .ZN(new_n744));
  INV_X1    g0544(.A(KEYINPUT31), .ZN(new_n745));
  AOI22_X1  g0545(.A1(new_n304), .A2(new_n306), .B1(new_n312), .B2(new_n626), .ZN(new_n746));
  OAI21_X1  g0546(.A(new_n746), .B1(new_n664), .B2(new_n312), .ZN(new_n747));
  NOR2_X1   g0547(.A1(new_n327), .A2(new_n747), .ZN(new_n748));
  NAND3_X1  g0548(.A1(new_n748), .A2(new_n580), .A3(new_n656), .ZN(new_n749));
  INV_X1    g0549(.A(KEYINPUT30), .ZN(new_n750));
  NAND2_X1  g0550(.A1(new_n749), .A2(new_n750), .ZN(new_n751));
  INV_X1    g0551(.A(KEYINPUT94), .ZN(new_n752));
  NOR2_X1   g0552(.A1(new_n751), .A2(new_n752), .ZN(new_n753));
  NOR2_X1   g0553(.A1(new_n623), .A2(new_n666), .ZN(new_n754));
  NOR3_X1   g0554(.A1(new_n664), .A2(KEYINPUT85), .A3(new_n312), .ZN(new_n755));
  OAI21_X1  g0555(.A(new_n746), .B1(new_n754), .B2(new_n755), .ZN(new_n756));
  NOR2_X1   g0556(.A1(new_n324), .A2(new_n367), .ZN(new_n757));
  NAND4_X1  g0557(.A1(new_n756), .A2(new_n757), .A3(new_n539), .A4(new_n599), .ZN(new_n758));
  NAND4_X1  g0558(.A1(new_n748), .A2(new_n580), .A3(new_n656), .A4(KEYINPUT30), .ZN(new_n759));
  NAND2_X1  g0559(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  AOI21_X1  g0560(.A(KEYINPUT94), .B1(new_n749), .B2(new_n750), .ZN(new_n761));
  NOR3_X1   g0561(.A1(new_n753), .A2(new_n760), .A3(new_n761), .ZN(new_n762));
  OAI21_X1  g0562(.A(new_n745), .B1(new_n762), .B2(new_n707), .ZN(new_n763));
  NAND4_X1  g0563(.A1(new_n571), .A2(new_n637), .A3(new_n330), .A4(new_n707), .ZN(new_n764));
  AND2_X1   g0564(.A1(new_n749), .A2(new_n750), .ZN(new_n765));
  OAI211_X1 g0565(.A(KEYINPUT31), .B(new_n706), .C1(new_n760), .C2(new_n765), .ZN(new_n766));
  NAND3_X1  g0566(.A1(new_n763), .A2(new_n764), .A3(new_n766), .ZN(new_n767));
  NAND2_X1  g0567(.A1(new_n767), .A2(G330), .ZN(new_n768));
  NAND2_X1  g0568(.A1(new_n744), .A2(new_n768), .ZN(new_n769));
  INV_X1    g0569(.A(new_n769), .ZN(new_n770));
  OAI21_X1  g0570(.A(new_n731), .B1(new_n770), .B2(G1), .ZN(G364));
  NAND3_X1  g0571(.A1(new_n215), .A2(G13), .A3(G45), .ZN(new_n772));
  NAND2_X1  g0572(.A1(new_n772), .A2(G1), .ZN(new_n773));
  NOR2_X1   g0573(.A1(new_n773), .A2(new_n728), .ZN(new_n774));
  NOR2_X1   g0574(.A1(new_n727), .A2(new_n299), .ZN(new_n775));
  NAND2_X1  g0575(.A1(new_n775), .A2(G355), .ZN(new_n776));
  OAI21_X1  g0576(.A(new_n776), .B1(G116), .B2(new_n210), .ZN(new_n777));
  NAND2_X1  g0577(.A1(new_n472), .A2(new_n473), .ZN(new_n778));
  NOR2_X1   g0578(.A1(new_n778), .A2(new_n727), .ZN(new_n779));
  INV_X1    g0579(.A(new_n779), .ZN(new_n780));
  AOI21_X1  g0580(.A(new_n780), .B1(new_n305), .B2(new_n220), .ZN(new_n781));
  OR2_X1    g0581(.A1(new_n245), .A2(new_n305), .ZN(new_n782));
  AOI21_X1  g0582(.A(new_n777), .B1(new_n781), .B2(new_n782), .ZN(new_n783));
  NOR2_X1   g0583(.A1(G13), .A2(G33), .ZN(new_n784));
  INV_X1    g0584(.A(new_n784), .ZN(new_n785));
  NOR2_X1   g0585(.A1(new_n785), .A2(G20), .ZN(new_n786));
  AOI21_X1  g0586(.A(new_n216), .B1(G20), .B2(new_n350), .ZN(new_n787));
  NOR2_X1   g0587(.A1(new_n786), .A2(new_n787), .ZN(new_n788));
  INV_X1    g0588(.A(new_n788), .ZN(new_n789));
  OAI21_X1  g0589(.A(new_n774), .B1(new_n783), .B2(new_n789), .ZN(new_n790));
  NAND3_X1  g0590(.A1(new_n367), .A2(G200), .A3(new_n279), .ZN(new_n791));
  NOR2_X1   g0591(.A1(new_n791), .A2(G190), .ZN(new_n792));
  XNOR2_X1  g0592(.A(KEYINPUT33), .B(G317), .ZN(new_n793));
  NOR2_X1   g0593(.A1(new_n366), .A2(G200), .ZN(new_n794));
  NOR2_X1   g0594(.A1(new_n215), .A2(new_n370), .ZN(new_n795));
  NAND2_X1  g0595(.A1(new_n794), .A2(new_n795), .ZN(new_n796));
  INV_X1    g0596(.A(new_n796), .ZN(new_n797));
  AOI22_X1  g0597(.A1(new_n792), .A2(new_n793), .B1(new_n797), .B2(G322), .ZN(new_n798));
  XOR2_X1   g0598(.A(new_n798), .B(KEYINPUT98), .Z(new_n799));
  NOR2_X1   g0599(.A1(new_n215), .A2(G190), .ZN(new_n800));
  NOR2_X1   g0600(.A1(new_n376), .A2(G179), .ZN(new_n801));
  NAND2_X1  g0601(.A1(new_n800), .A2(new_n801), .ZN(new_n802));
  INV_X1    g0602(.A(G283), .ZN(new_n803));
  NOR2_X1   g0603(.A1(G179), .A2(G200), .ZN(new_n804));
  AOI21_X1  g0604(.A(new_n215), .B1(G190), .B2(new_n804), .ZN(new_n805));
  INV_X1    g0605(.A(G294), .ZN(new_n806));
  OAI22_X1  g0606(.A1(new_n802), .A2(new_n803), .B1(new_n805), .B2(new_n806), .ZN(new_n807));
  NAND2_X1  g0607(.A1(new_n800), .A2(new_n804), .ZN(new_n808));
  INV_X1    g0608(.A(new_n808), .ZN(new_n809));
  AOI21_X1  g0609(.A(new_n807), .B1(G329), .B2(new_n809), .ZN(new_n810));
  NAND3_X1  g0610(.A1(new_n801), .A2(G20), .A3(G190), .ZN(new_n811));
  NAND2_X1  g0611(.A1(new_n794), .A2(new_n800), .ZN(new_n812));
  INV_X1    g0612(.A(G311), .ZN(new_n813));
  OAI221_X1 g0613(.A(new_n299), .B1(new_n293), .B2(new_n811), .C1(new_n812), .C2(new_n813), .ZN(new_n814));
  NOR2_X1   g0614(.A1(new_n791), .A2(new_n370), .ZN(new_n815));
  AOI21_X1  g0615(.A(new_n814), .B1(G326), .B2(new_n815), .ZN(new_n816));
  NAND3_X1  g0616(.A1(new_n799), .A2(new_n810), .A3(new_n816), .ZN(new_n817));
  INV_X1    g0617(.A(new_n812), .ZN(new_n818));
  AOI22_X1  g0618(.A1(G58), .A2(new_n797), .B1(new_n818), .B2(G77), .ZN(new_n819));
  INV_X1    g0619(.A(new_n815), .ZN(new_n820));
  OAI21_X1  g0620(.A(new_n819), .B1(new_n202), .B2(new_n820), .ZN(new_n821));
  XOR2_X1   g0621(.A(new_n821), .B(KEYINPUT97), .Z(new_n822));
  NOR2_X1   g0622(.A1(new_n802), .A2(new_n206), .ZN(new_n823));
  NOR2_X1   g0623(.A1(new_n805), .A2(new_n205), .ZN(new_n824));
  AOI21_X1  g0624(.A(new_n811), .B1(new_n608), .B2(new_n610), .ZN(new_n825));
  OR4_X1    g0625(.A1(new_n299), .A2(new_n823), .A3(new_n824), .A4(new_n825), .ZN(new_n826));
  NOR3_X1   g0626(.A1(new_n808), .A2(KEYINPUT32), .A3(new_n509), .ZN(new_n827));
  OAI21_X1  g0627(.A(KEYINPUT32), .B1(new_n808), .B2(new_n509), .ZN(new_n828));
  INV_X1    g0628(.A(new_n792), .ZN(new_n829));
  OAI21_X1  g0629(.A(new_n828), .B1(new_n829), .B2(new_n408), .ZN(new_n830));
  OR3_X1    g0630(.A1(new_n826), .A2(new_n827), .A3(new_n830), .ZN(new_n831));
  OAI21_X1  g0631(.A(new_n817), .B1(new_n822), .B2(new_n831), .ZN(new_n832));
  AOI21_X1  g0632(.A(new_n790), .B1(new_n832), .B2(new_n787), .ZN(new_n833));
  INV_X1    g0633(.A(new_n786), .ZN(new_n834));
  OAI21_X1  g0634(.A(new_n833), .B1(new_n715), .B2(new_n834), .ZN(new_n835));
  XNOR2_X1  g0635(.A(new_n835), .B(KEYINPUT99), .ZN(new_n836));
  NOR2_X1   g0636(.A1(new_n716), .A2(new_n718), .ZN(new_n837));
  INV_X1    g0637(.A(new_n774), .ZN(new_n838));
  OAI211_X1 g0638(.A(new_n837), .B(new_n838), .C1(G330), .C2(new_n715), .ZN(new_n839));
  NAND2_X1  g0639(.A1(new_n836), .A2(new_n839), .ZN(G396));
  INV_X1    g0640(.A(new_n465), .ZN(new_n841));
  NAND2_X1  g0641(.A1(new_n706), .A2(new_n462), .ZN(new_n842));
  AOI21_X1  g0642(.A(new_n841), .B1(new_n461), .B2(new_n842), .ZN(new_n843));
  NOR2_X1   g0643(.A1(new_n465), .A2(new_n706), .ZN(new_n844));
  OAI21_X1  g0644(.A(KEYINPUT102), .B1(new_n843), .B2(new_n844), .ZN(new_n845));
  INV_X1    g0645(.A(KEYINPUT102), .ZN(new_n846));
  INV_X1    g0646(.A(new_n844), .ZN(new_n847));
  AOI21_X1  g0647(.A(new_n459), .B1(new_n455), .B2(KEYINPUT71), .ZN(new_n848));
  AOI22_X1  g0648(.A1(new_n848), .A2(new_n458), .B1(new_n462), .B2(new_n706), .ZN(new_n849));
  OAI211_X1 g0649(.A(new_n846), .B(new_n847), .C1(new_n849), .C2(new_n841), .ZN(new_n850));
  NAND2_X1  g0650(.A1(new_n845), .A2(new_n850), .ZN(new_n851));
  OAI211_X1 g0651(.A(new_n851), .B(new_n707), .C1(new_n689), .C2(new_n692), .ZN(new_n852));
  INV_X1    g0652(.A(KEYINPUT103), .ZN(new_n853));
  NAND2_X1  g0653(.A1(new_n851), .A2(new_n853), .ZN(new_n854));
  NAND3_X1  g0654(.A1(new_n845), .A2(KEYINPUT103), .A3(new_n850), .ZN(new_n855));
  NAND2_X1  g0655(.A1(new_n854), .A2(new_n855), .ZN(new_n856));
  OAI21_X1  g0656(.A(new_n852), .B1(new_n741), .B2(new_n856), .ZN(new_n857));
  AOI21_X1  g0657(.A(new_n774), .B1(new_n857), .B2(new_n768), .ZN(new_n858));
  OAI21_X1  g0658(.A(new_n858), .B1(new_n768), .B2(new_n857), .ZN(new_n859));
  NOR2_X1   g0659(.A1(new_n787), .A2(new_n784), .ZN(new_n860));
  INV_X1    g0660(.A(new_n860), .ZN(new_n861));
  OAI21_X1  g0661(.A(new_n774), .B1(G77), .B2(new_n861), .ZN(new_n862));
  OAI21_X1  g0662(.A(new_n299), .B1(new_n811), .B2(new_n206), .ZN(new_n863));
  XOR2_X1   g0663(.A(KEYINPUT100), .B(G283), .Z(new_n864));
  INV_X1    g0664(.A(new_n864), .ZN(new_n865));
  AOI211_X1 g0665(.A(new_n863), .B(new_n824), .C1(new_n792), .C2(new_n865), .ZN(new_n866));
  NOR2_X1   g0666(.A1(new_n802), .A2(new_n542), .ZN(new_n867));
  AOI21_X1  g0667(.A(new_n867), .B1(G294), .B2(new_n797), .ZN(new_n868));
  AOI22_X1  g0668(.A1(new_n818), .A2(new_n257), .B1(new_n809), .B2(G311), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n815), .A2(G303), .ZN(new_n870));
  NAND4_X1  g0670(.A1(new_n866), .A2(new_n868), .A3(new_n869), .A4(new_n870), .ZN(new_n871));
  AOI22_X1  g0671(.A1(G143), .A2(new_n797), .B1(new_n818), .B2(G159), .ZN(new_n872));
  INV_X1    g0672(.A(G137), .ZN(new_n873));
  INV_X1    g0673(.A(G150), .ZN(new_n874));
  OAI221_X1 g0674(.A(new_n872), .B1(new_n873), .B2(new_n820), .C1(new_n874), .C2(new_n829), .ZN(new_n875));
  XOR2_X1   g0675(.A(new_n875), .B(KEYINPUT101), .Z(new_n876));
  NAND2_X1  g0676(.A1(new_n876), .A2(KEYINPUT34), .ZN(new_n877));
  INV_X1    g0677(.A(new_n802), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n878), .A2(G68), .ZN(new_n879));
  INV_X1    g0679(.A(new_n778), .ZN(new_n880));
  INV_X1    g0680(.A(new_n811), .ZN(new_n881));
  AOI21_X1  g0681(.A(new_n880), .B1(G50), .B2(new_n881), .ZN(new_n882));
  INV_X1    g0682(.A(new_n805), .ZN(new_n883));
  AOI22_X1  g0683(.A1(new_n809), .A2(G132), .B1(new_n883), .B2(G58), .ZN(new_n884));
  NAND4_X1  g0684(.A1(new_n877), .A2(new_n879), .A3(new_n882), .A4(new_n884), .ZN(new_n885));
  NOR2_X1   g0685(.A1(new_n876), .A2(KEYINPUT34), .ZN(new_n886));
  OAI21_X1  g0686(.A(new_n871), .B1(new_n885), .B2(new_n886), .ZN(new_n887));
  AOI21_X1  g0687(.A(new_n862), .B1(new_n887), .B2(new_n787), .ZN(new_n888));
  OAI21_X1  g0688(.A(new_n888), .B1(new_n785), .B2(new_n851), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n859), .A2(new_n889), .ZN(G384));
  INV_X1    g0690(.A(new_n586), .ZN(new_n891));
  OR2_X1    g0691(.A1(new_n891), .A2(KEYINPUT35), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n891), .A2(KEYINPUT35), .ZN(new_n893));
  NAND4_X1  g0693(.A1(new_n892), .A2(G116), .A3(new_n217), .A4(new_n893), .ZN(new_n894));
  XOR2_X1   g0694(.A(new_n894), .B(KEYINPUT36), .Z(new_n895));
  OAI211_X1 g0695(.A(new_n220), .B(G77), .C1(new_n435), .C2(new_n222), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n202), .A2(G68), .ZN(new_n897));
  AOI211_X1 g0697(.A(new_n258), .B(G13), .C1(new_n896), .C2(new_n897), .ZN(new_n898));
  NOR2_X1   g0698(.A1(new_n895), .A2(new_n898), .ZN(new_n899));
  INV_X1    g0699(.A(KEYINPUT38), .ZN(new_n900));
  AOI21_X1  g0700(.A(KEYINPUT16), .B1(new_n470), .B2(new_n478), .ZN(new_n901));
  OAI21_X1  g0701(.A(new_n468), .B1(new_n480), .B2(new_n901), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n902), .A2(new_n504), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n703), .A2(new_n705), .ZN(new_n904));
  INV_X1    g0704(.A(new_n904), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n902), .A2(new_n905), .ZN(new_n906));
  NAND3_X1  g0706(.A1(new_n903), .A2(new_n906), .A3(new_n521), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n907), .A2(KEYINPUT37), .ZN(new_n908));
  INV_X1    g0708(.A(KEYINPUT105), .ZN(new_n909));
  INV_X1    g0709(.A(KEYINPUT104), .ZN(new_n910));
  NAND3_X1  g0710(.A1(new_n490), .A2(new_n905), .A3(new_n910), .ZN(new_n911));
  INV_X1    g0711(.A(new_n911), .ZN(new_n912));
  AOI21_X1  g0712(.A(new_n910), .B1(new_n490), .B2(new_n905), .ZN(new_n913));
  NOR2_X1   g0713(.A1(new_n912), .A2(new_n913), .ZN(new_n914));
  INV_X1    g0714(.A(KEYINPUT37), .ZN(new_n915));
  NAND3_X1  g0715(.A1(new_n505), .A2(new_n521), .A3(new_n915), .ZN(new_n916));
  OAI211_X1 g0716(.A(new_n908), .B(new_n909), .C1(new_n914), .C2(new_n916), .ZN(new_n917));
  NAND3_X1  g0717(.A1(new_n526), .A2(new_n905), .A3(new_n902), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n917), .A2(new_n918), .ZN(new_n919));
  INV_X1    g0719(.A(new_n913), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n920), .A2(new_n911), .ZN(new_n921));
  INV_X1    g0721(.A(new_n916), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n921), .A2(new_n922), .ZN(new_n923));
  AOI21_X1  g0723(.A(new_n909), .B1(new_n923), .B2(new_n908), .ZN(new_n924));
  OAI21_X1  g0724(.A(new_n900), .B1(new_n919), .B2(new_n924), .ZN(new_n925));
  AOI21_X1  g0725(.A(new_n916), .B1(new_n911), .B2(new_n920), .ZN(new_n926));
  AOI22_X1  g0726(.A1(new_n515), .A2(new_n517), .B1(new_n905), .B2(new_n902), .ZN(new_n927));
  AOI21_X1  g0727(.A(new_n915), .B1(new_n927), .B2(new_n903), .ZN(new_n928));
  OAI21_X1  g0728(.A(KEYINPUT105), .B1(new_n926), .B2(new_n928), .ZN(new_n929));
  NAND4_X1  g0729(.A1(new_n929), .A2(KEYINPUT38), .A3(new_n918), .A4(new_n917), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n925), .A2(new_n930), .ZN(new_n931));
  OAI211_X1 g0731(.A(new_n759), .B(new_n758), .C1(new_n765), .C2(KEYINPUT94), .ZN(new_n932));
  OAI211_X1 g0732(.A(KEYINPUT31), .B(new_n706), .C1(new_n932), .C2(new_n753), .ZN(new_n933));
  NAND3_X1  g0733(.A1(new_n763), .A2(new_n764), .A3(new_n933), .ZN(new_n934));
  AOI22_X1  g0734(.A1(new_n425), .A2(new_n424), .B1(new_n395), .B2(G179), .ZN(new_n935));
  OAI21_X1  g0735(.A(KEYINPUT14), .B1(new_n395), .B2(new_n350), .ZN(new_n936));
  AOI21_X1  g0736(.A(new_n416), .B1(new_n935), .B2(new_n936), .ZN(new_n937));
  OAI211_X1 g0737(.A(new_n423), .B(new_n706), .C1(new_n937), .C2(new_n642), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n423), .A2(new_n706), .ZN(new_n939));
  NAND3_X1  g0739(.A1(new_n422), .A2(new_n430), .A3(new_n939), .ZN(new_n940));
  NAND2_X1  g0740(.A1(new_n938), .A2(new_n940), .ZN(new_n941));
  AND3_X1   g0741(.A1(new_n934), .A2(new_n941), .A3(new_n851), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n931), .A2(new_n942), .ZN(new_n943));
  XOR2_X1   g0743(.A(KEYINPUT106), .B(KEYINPUT40), .Z(new_n944));
  INV_X1    g0744(.A(new_n944), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n943), .A2(new_n945), .ZN(new_n946));
  AOI21_X1  g0746(.A(new_n921), .B1(new_n646), .B2(new_n644), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n505), .A2(new_n521), .ZN(new_n948));
  OAI21_X1  g0748(.A(KEYINPUT37), .B1(new_n914), .B2(new_n948), .ZN(new_n949));
  OAI211_X1 g0749(.A(new_n900), .B(new_n923), .C1(new_n947), .C2(new_n949), .ZN(new_n950));
  NAND2_X1  g0750(.A1(new_n930), .A2(new_n950), .ZN(new_n951));
  NAND3_X1  g0751(.A1(new_n951), .A2(new_n942), .A3(KEYINPUT40), .ZN(new_n952));
  AND2_X1   g0752(.A1(new_n946), .A2(new_n952), .ZN(new_n953));
  AND2_X1   g0753(.A1(new_n527), .A2(new_n934), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n953), .A2(new_n954), .ZN(new_n955));
  INV_X1    g0755(.A(new_n955), .ZN(new_n956));
  NOR2_X1   g0756(.A1(new_n953), .A2(new_n954), .ZN(new_n957));
  NOR3_X1   g0757(.A1(new_n956), .A2(new_n717), .A3(new_n957), .ZN(new_n958));
  INV_X1    g0758(.A(KEYINPUT39), .ZN(new_n959));
  NAND2_X1  g0759(.A1(new_n951), .A2(new_n959), .ZN(new_n960));
  NAND3_X1  g0760(.A1(new_n925), .A2(KEYINPUT39), .A3(new_n930), .ZN(new_n961));
  NAND2_X1  g0761(.A1(new_n937), .A2(new_n707), .ZN(new_n962));
  INV_X1    g0762(.A(new_n962), .ZN(new_n963));
  NAND3_X1  g0763(.A1(new_n960), .A2(new_n961), .A3(new_n963), .ZN(new_n964));
  INV_X1    g0764(.A(new_n941), .ZN(new_n965));
  AOI21_X1  g0765(.A(new_n965), .B1(new_n852), .B2(new_n847), .ZN(new_n966));
  NAND2_X1  g0766(.A1(new_n966), .A2(new_n931), .ZN(new_n967));
  OR2_X1    g0767(.A1(new_n646), .A2(new_n905), .ZN(new_n968));
  AND3_X1   g0768(.A1(new_n964), .A2(new_n967), .A3(new_n968), .ZN(new_n969));
  OAI211_X1 g0769(.A(new_n527), .B(new_n740), .C1(new_n741), .C2(new_n743), .ZN(new_n970));
  NAND2_X1  g0770(.A1(new_n651), .A2(new_n970), .ZN(new_n971));
  XNOR2_X1  g0771(.A(new_n969), .B(new_n971), .ZN(new_n972));
  NAND2_X1  g0772(.A1(new_n958), .A2(new_n972), .ZN(new_n973));
  INV_X1    g0773(.A(G13), .ZN(new_n974));
  OAI21_X1  g0774(.A(G1), .B1(new_n279), .B2(new_n974), .ZN(new_n975));
  NAND3_X1  g0775(.A1(new_n973), .A2(KEYINPUT107), .A3(new_n975), .ZN(new_n976));
  OAI21_X1  g0776(.A(new_n976), .B1(new_n972), .B2(new_n958), .ZN(new_n977));
  AOI21_X1  g0777(.A(KEYINPUT107), .B1(new_n973), .B2(new_n975), .ZN(new_n978));
  OAI21_X1  g0778(.A(new_n899), .B1(new_n977), .B2(new_n978), .ZN(G367));
  AND2_X1   g0779(.A1(new_n236), .A2(new_n779), .ZN(new_n980));
  OAI21_X1  g0780(.A(new_n788), .B1(new_n210), .B2(new_n431), .ZN(new_n981));
  OAI21_X1  g0781(.A(new_n774), .B1(new_n980), .B2(new_n981), .ZN(new_n982));
  AOI22_X1  g0782(.A1(new_n797), .A2(G303), .B1(G107), .B2(new_n883), .ZN(new_n983));
  INV_X1    g0783(.A(KEYINPUT46), .ZN(new_n984));
  OAI21_X1  g0784(.A(new_n984), .B1(new_n811), .B2(new_n261), .ZN(new_n985));
  NAND3_X1  g0785(.A1(new_n881), .A2(KEYINPUT46), .A3(G116), .ZN(new_n986));
  AND4_X1   g0786(.A1(new_n880), .A2(new_n983), .A3(new_n985), .A4(new_n986), .ZN(new_n987));
  OAI221_X1 g0787(.A(new_n987), .B1(new_n806), .B2(new_n829), .C1(new_n813), .C2(new_n820), .ZN(new_n988));
  NAND2_X1  g0788(.A1(new_n878), .A2(G97), .ZN(new_n989));
  INV_X1    g0789(.A(G317), .ZN(new_n990));
  OAI221_X1 g0790(.A(new_n989), .B1(new_n990), .B2(new_n808), .C1(new_n812), .C2(new_n864), .ZN(new_n991));
  AOI22_X1  g0791(.A1(G50), .A2(new_n818), .B1(new_n797), .B2(G150), .ZN(new_n992));
  NAND2_X1  g0792(.A1(new_n883), .A2(G68), .ZN(new_n993));
  OAI211_X1 g0793(.A(new_n992), .B(new_n993), .C1(new_n873), .C2(new_n808), .ZN(new_n994));
  NAND2_X1  g0794(.A1(new_n792), .A2(G159), .ZN(new_n995));
  NAND2_X1  g0795(.A1(new_n815), .A2(G143), .ZN(new_n996));
  NOR2_X1   g0796(.A1(new_n802), .A2(new_n355), .ZN(new_n997));
  INV_X1    g0797(.A(new_n997), .ZN(new_n998));
  AOI21_X1  g0798(.A(new_n299), .B1(new_n881), .B2(G58), .ZN(new_n999));
  NAND4_X1  g0799(.A1(new_n995), .A2(new_n996), .A3(new_n998), .A4(new_n999), .ZN(new_n1000));
  OAI22_X1  g0800(.A1(new_n988), .A2(new_n991), .B1(new_n994), .B2(new_n1000), .ZN(new_n1001));
  XNOR2_X1  g0801(.A(new_n1001), .B(KEYINPUT47), .ZN(new_n1002));
  AOI21_X1  g0802(.A(new_n982), .B1(new_n1002), .B2(new_n787), .ZN(new_n1003));
  OR2_X1    g0803(.A1(new_n707), .A2(new_n633), .ZN(new_n1004));
  NOR2_X1   g0804(.A1(new_n1004), .A2(new_n674), .ZN(new_n1005));
  AOI21_X1  g0805(.A(new_n1005), .B1(new_n734), .B2(new_n1004), .ZN(new_n1006));
  NAND2_X1  g0806(.A1(new_n1006), .A2(new_n786), .ZN(new_n1007));
  NAND2_X1  g0807(.A1(new_n1003), .A2(new_n1007), .ZN(new_n1008));
  INV_X1    g0808(.A(new_n1008), .ZN(new_n1009));
  INV_X1    g0809(.A(new_n773), .ZN(new_n1010));
  NAND2_X1  g0810(.A1(KEYINPUT109), .A2(KEYINPUT44), .ZN(new_n1011));
  INV_X1    g0811(.A(new_n1011), .ZN(new_n1012));
  NAND2_X1  g0812(.A1(new_n706), .A2(new_n593), .ZN(new_n1013));
  OAI211_X1 g0813(.A(new_n1013), .B(new_n682), .C1(new_n600), .C2(new_n596), .ZN(new_n1014));
  NAND2_X1  g0814(.A1(new_n684), .A2(new_n706), .ZN(new_n1015));
  NAND2_X1  g0815(.A1(new_n1014), .A2(new_n1015), .ZN(new_n1016));
  INV_X1    g0816(.A(new_n1016), .ZN(new_n1017));
  NAND2_X1  g0817(.A1(new_n722), .A2(new_n1017), .ZN(new_n1018));
  NOR2_X1   g0818(.A1(KEYINPUT109), .A2(KEYINPUT44), .ZN(new_n1019));
  AOI21_X1  g0819(.A(new_n1012), .B1(new_n1018), .B2(new_n1019), .ZN(new_n1020));
  OAI21_X1  g0820(.A(new_n1020), .B1(new_n1018), .B2(new_n1019), .ZN(new_n1021));
  NOR2_X1   g0821(.A1(new_n722), .A2(new_n1017), .ZN(new_n1022));
  XNOR2_X1  g0822(.A(new_n1022), .B(KEYINPUT45), .ZN(new_n1023));
  NAND2_X1  g0823(.A1(new_n1021), .A2(new_n1023), .ZN(new_n1024));
  INV_X1    g0824(.A(KEYINPUT111), .ZN(new_n1025));
  NAND3_X1  g0825(.A1(new_n1024), .A2(new_n1025), .A3(new_n719), .ZN(new_n1026));
  NAND2_X1  g0826(.A1(new_n719), .A2(new_n1025), .ZN(new_n1027));
  OAI211_X1 g0827(.A(KEYINPUT111), .B(new_n710), .C1(new_n716), .C2(new_n718), .ZN(new_n1028));
  NAND4_X1  g0828(.A1(new_n1027), .A2(new_n1028), .A3(new_n1023), .A4(new_n1021), .ZN(new_n1029));
  NAND2_X1  g0829(.A1(new_n1026), .A2(new_n1029), .ZN(new_n1030));
  NOR2_X1   g0830(.A1(new_n720), .A2(KEYINPUT110), .ZN(new_n1031));
  INV_X1    g0831(.A(new_n720), .ZN(new_n1032));
  NAND2_X1  g0832(.A1(new_n713), .A2(new_n707), .ZN(new_n1033));
  NAND3_X1  g0833(.A1(new_n708), .A2(new_n709), .A3(new_n1033), .ZN(new_n1034));
  INV_X1    g0834(.A(KEYINPUT110), .ZN(new_n1035));
  AOI21_X1  g0835(.A(new_n1032), .B1(new_n1034), .B2(new_n1035), .ZN(new_n1036));
  OAI21_X1  g0836(.A(new_n837), .B1(new_n1031), .B2(new_n1036), .ZN(new_n1037));
  NOR2_X1   g0837(.A1(new_n1036), .A2(new_n1031), .ZN(new_n1038));
  OAI21_X1  g0838(.A(new_n1038), .B1(new_n718), .B2(new_n716), .ZN(new_n1039));
  NAND2_X1  g0839(.A1(new_n1037), .A2(new_n1039), .ZN(new_n1040));
  INV_X1    g0840(.A(new_n1040), .ZN(new_n1041));
  AOI21_X1  g0841(.A(new_n769), .B1(new_n1030), .B2(new_n1041), .ZN(new_n1042));
  XOR2_X1   g0842(.A(new_n728), .B(KEYINPUT41), .Z(new_n1043));
  OAI21_X1  g0843(.A(new_n1010), .B1(new_n1042), .B2(new_n1043), .ZN(new_n1044));
  NAND2_X1  g0844(.A1(new_n1032), .A2(new_n1016), .ZN(new_n1045));
  OR2_X1    g0845(.A1(new_n1045), .A2(KEYINPUT42), .ZN(new_n1046));
  OAI21_X1  g0846(.A(new_n682), .B1(new_n1014), .B2(new_n660), .ZN(new_n1047));
  AOI22_X1  g0847(.A1(new_n1045), .A2(KEYINPUT42), .B1(new_n707), .B2(new_n1047), .ZN(new_n1048));
  NAND2_X1  g0848(.A1(new_n1046), .A2(new_n1048), .ZN(new_n1049));
  INV_X1    g0849(.A(KEYINPUT43), .ZN(new_n1050));
  NAND2_X1  g0850(.A1(new_n1006), .A2(new_n1050), .ZN(new_n1051));
  OR2_X1    g0851(.A1(new_n1006), .A2(new_n1050), .ZN(new_n1052));
  NAND3_X1  g0852(.A1(new_n1049), .A2(new_n1051), .A3(new_n1052), .ZN(new_n1053));
  NAND4_X1  g0853(.A1(new_n1046), .A2(new_n1048), .A3(new_n1050), .A4(new_n1006), .ZN(new_n1054));
  NAND2_X1  g0854(.A1(new_n1053), .A2(new_n1054), .ZN(new_n1055));
  NOR2_X1   g0855(.A1(new_n719), .A2(new_n1017), .ZN(new_n1056));
  INV_X1    g0856(.A(new_n1056), .ZN(new_n1057));
  OAI21_X1  g0857(.A(KEYINPUT108), .B1(new_n1055), .B2(new_n1057), .ZN(new_n1058));
  NAND2_X1  g0858(.A1(new_n1055), .A2(new_n1057), .ZN(new_n1059));
  NAND2_X1  g0859(.A1(new_n1058), .A2(new_n1059), .ZN(new_n1060));
  NOR3_X1   g0860(.A1(new_n1055), .A2(new_n1057), .A3(KEYINPUT108), .ZN(new_n1061));
  NOR2_X1   g0861(.A1(new_n1060), .A2(new_n1061), .ZN(new_n1062));
  AOI21_X1  g0862(.A(new_n1009), .B1(new_n1044), .B2(new_n1062), .ZN(new_n1063));
  INV_X1    g0863(.A(KEYINPUT112), .ZN(new_n1064));
  AND2_X1   g0864(.A1(new_n1063), .A2(new_n1064), .ZN(new_n1065));
  NOR2_X1   g0865(.A1(new_n1063), .A2(new_n1064), .ZN(new_n1066));
  NOR2_X1   g0866(.A1(new_n1065), .A2(new_n1066), .ZN(G387));
  NOR2_X1   g0867(.A1(new_n769), .A2(new_n1040), .ZN(new_n1068));
  INV_X1    g0868(.A(new_n728), .ZN(new_n1069));
  OAI21_X1  g0869(.A(KEYINPUT114), .B1(new_n1068), .B2(new_n1069), .ZN(new_n1070));
  NAND2_X1  g0870(.A1(new_n769), .A2(new_n1040), .ZN(new_n1071));
  INV_X1    g0871(.A(KEYINPUT114), .ZN(new_n1072));
  OAI211_X1 g0872(.A(new_n1072), .B(new_n728), .C1(new_n769), .C2(new_n1040), .ZN(new_n1073));
  NAND3_X1  g0873(.A1(new_n1070), .A2(new_n1071), .A3(new_n1073), .ZN(new_n1074));
  NAND2_X1  g0874(.A1(new_n1041), .A2(new_n773), .ZN(new_n1075));
  NAND2_X1  g0875(.A1(new_n881), .A2(G77), .ZN(new_n1076));
  NAND3_X1  g0876(.A1(new_n989), .A2(new_n778), .A3(new_n1076), .ZN(new_n1077));
  AOI21_X1  g0877(.A(new_n1077), .B1(G159), .B2(new_n815), .ZN(new_n1078));
  AOI22_X1  g0878(.A1(new_n809), .A2(G150), .B1(new_n883), .B2(new_n432), .ZN(new_n1079));
  AOI22_X1  g0879(.A1(G50), .A2(new_n797), .B1(new_n818), .B2(G68), .ZN(new_n1080));
  INV_X1    g0880(.A(new_n346), .ZN(new_n1081));
  NAND2_X1  g0881(.A1(new_n792), .A2(new_n1081), .ZN(new_n1082));
  NAND4_X1  g0882(.A1(new_n1078), .A2(new_n1079), .A3(new_n1080), .A4(new_n1082), .ZN(new_n1083));
  AOI21_X1  g0883(.A(new_n778), .B1(new_n809), .B2(G326), .ZN(new_n1084));
  OAI22_X1  g0884(.A1(new_n805), .A2(new_n864), .B1(new_n806), .B2(new_n811), .ZN(new_n1085));
  AOI22_X1  g0885(.A1(G303), .A2(new_n818), .B1(new_n797), .B2(G317), .ZN(new_n1086));
  INV_X1    g0886(.A(G322), .ZN(new_n1087));
  OAI221_X1 g0887(.A(new_n1086), .B1(new_n813), .B2(new_n829), .C1(new_n1087), .C2(new_n820), .ZN(new_n1088));
  INV_X1    g0888(.A(KEYINPUT48), .ZN(new_n1089));
  AOI21_X1  g0889(.A(new_n1085), .B1(new_n1088), .B2(new_n1089), .ZN(new_n1090));
  OAI21_X1  g0890(.A(new_n1090), .B1(new_n1089), .B2(new_n1088), .ZN(new_n1091));
  INV_X1    g0891(.A(KEYINPUT49), .ZN(new_n1092));
  OAI221_X1 g0892(.A(new_n1084), .B1(new_n261), .B2(new_n802), .C1(new_n1091), .C2(new_n1092), .ZN(new_n1093));
  AND2_X1   g0893(.A1(new_n1091), .A2(new_n1092), .ZN(new_n1094));
  OAI21_X1  g0894(.A(new_n1083), .B1(new_n1093), .B2(new_n1094), .ZN(new_n1095));
  NAND2_X1  g0895(.A1(new_n1095), .A2(new_n787), .ZN(new_n1096));
  AOI21_X1  g0896(.A(new_n780), .B1(new_n241), .B2(G45), .ZN(new_n1097));
  AOI21_X1  g0897(.A(new_n1097), .B1(new_n726), .B2(new_n775), .ZN(new_n1098));
  NOR2_X1   g0898(.A1(new_n341), .A2(G50), .ZN(new_n1099));
  INV_X1    g0899(.A(KEYINPUT50), .ZN(new_n1100));
  OAI221_X1 g0900(.A(new_n305), .B1(new_n408), .B2(new_n355), .C1(new_n1099), .C2(new_n1100), .ZN(new_n1101));
  AOI211_X1 g0901(.A(new_n1101), .B(new_n726), .C1(new_n1100), .C2(new_n1099), .ZN(new_n1102));
  OAI22_X1  g0902(.A1(new_n1098), .A2(new_n1102), .B1(G107), .B2(new_n210), .ZN(new_n1103));
  AOI21_X1  g0903(.A(new_n838), .B1(new_n1103), .B2(new_n788), .ZN(new_n1104));
  XOR2_X1   g0904(.A(new_n1104), .B(KEYINPUT113), .Z(new_n1105));
  OAI211_X1 g0905(.A(new_n1096), .B(new_n1105), .C1(new_n710), .C2(new_n834), .ZN(new_n1106));
  AND2_X1   g0906(.A1(new_n1075), .A2(new_n1106), .ZN(new_n1107));
  NAND2_X1  g0907(.A1(new_n1074), .A2(new_n1107), .ZN(G393));
  NAND2_X1  g0908(.A1(new_n1030), .A2(new_n773), .ZN(new_n1109));
  OAI221_X1 g0909(.A(new_n788), .B1(new_n205), .B2(new_n210), .C1(new_n780), .C2(new_n250), .ZN(new_n1110));
  NAND2_X1  g0910(.A1(new_n1110), .A2(new_n774), .ZN(new_n1111));
  AOI22_X1  g0911(.A1(new_n815), .A2(G317), .B1(new_n797), .B2(G311), .ZN(new_n1112));
  XOR2_X1   g0912(.A(new_n1112), .B(KEYINPUT52), .Z(new_n1113));
  OAI22_X1  g0913(.A1(new_n808), .A2(new_n1087), .B1(new_n805), .B2(new_n261), .ZN(new_n1114));
  AOI21_X1  g0914(.A(new_n1114), .B1(G294), .B2(new_n818), .ZN(new_n1115));
  OAI21_X1  g0915(.A(new_n299), .B1(new_n864), .B2(new_n811), .ZN(new_n1116));
  AOI211_X1 g0916(.A(new_n1116), .B(new_n823), .C1(G303), .C2(new_n792), .ZN(new_n1117));
  NAND3_X1  g0917(.A1(new_n1113), .A2(new_n1115), .A3(new_n1117), .ZN(new_n1118));
  AOI22_X1  g0918(.A1(new_n815), .A2(G150), .B1(new_n797), .B2(G159), .ZN(new_n1119));
  XNOR2_X1  g0919(.A(new_n1119), .B(KEYINPUT51), .ZN(new_n1120));
  OAI21_X1  g0920(.A(new_n778), .B1(new_n222), .B2(new_n811), .ZN(new_n1121));
  AOI211_X1 g0921(.A(new_n1121), .B(new_n867), .C1(G50), .C2(new_n792), .ZN(new_n1122));
  AOI22_X1  g0922(.A1(new_n818), .A2(new_n437), .B1(new_n809), .B2(G143), .ZN(new_n1123));
  OAI211_X1 g0923(.A(new_n1122), .B(new_n1123), .C1(new_n355), .C2(new_n805), .ZN(new_n1124));
  OAI21_X1  g0924(.A(new_n1118), .B1(new_n1120), .B2(new_n1124), .ZN(new_n1125));
  AOI21_X1  g0925(.A(new_n1111), .B1(new_n1125), .B2(new_n787), .ZN(new_n1126));
  OAI21_X1  g0926(.A(new_n1126), .B1(new_n1016), .B2(new_n834), .ZN(new_n1127));
  AOI21_X1  g0927(.A(new_n1069), .B1(new_n1030), .B2(new_n1068), .ZN(new_n1128));
  INV_X1    g0928(.A(KEYINPUT115), .ZN(new_n1129));
  OAI211_X1 g0929(.A(new_n1026), .B(new_n1029), .C1(new_n769), .C2(new_n1040), .ZN(new_n1130));
  NAND3_X1  g0930(.A1(new_n1128), .A2(new_n1129), .A3(new_n1130), .ZN(new_n1131));
  INV_X1    g0931(.A(new_n1131), .ZN(new_n1132));
  AOI21_X1  g0932(.A(new_n1129), .B1(new_n1128), .B2(new_n1130), .ZN(new_n1133));
  OAI211_X1 g0933(.A(new_n1109), .B(new_n1127), .C1(new_n1132), .C2(new_n1133), .ZN(G390));
  NAND4_X1  g0934(.A1(new_n934), .A2(new_n941), .A3(new_n851), .A4(G330), .ZN(new_n1135));
  INV_X1    g0935(.A(new_n1135), .ZN(new_n1136));
  NAND2_X1  g0936(.A1(new_n852), .A2(new_n847), .ZN(new_n1137));
  NAND2_X1  g0937(.A1(new_n1137), .A2(new_n941), .ZN(new_n1138));
  AOI22_X1  g0938(.A1(new_n1138), .A2(new_n962), .B1(new_n960), .B2(new_n961), .ZN(new_n1139));
  NAND2_X1  g0939(.A1(new_n951), .A2(new_n962), .ZN(new_n1140));
  NAND3_X1  g0940(.A1(new_n739), .A2(new_n707), .A3(new_n851), .ZN(new_n1141));
  NAND2_X1  g0941(.A1(new_n1141), .A2(new_n847), .ZN(new_n1142));
  AOI21_X1  g0942(.A(new_n1140), .B1(new_n941), .B2(new_n1142), .ZN(new_n1143));
  OAI21_X1  g0943(.A(new_n1136), .B1(new_n1139), .B2(new_n1143), .ZN(new_n1144));
  AND3_X1   g0944(.A1(new_n925), .A2(KEYINPUT39), .A3(new_n930), .ZN(new_n1145));
  AOI21_X1  g0945(.A(KEYINPUT39), .B1(new_n930), .B2(new_n950), .ZN(new_n1146));
  OAI22_X1  g0946(.A1(new_n1145), .A2(new_n1146), .B1(new_n966), .B2(new_n963), .ZN(new_n1147));
  NAND2_X1  g0947(.A1(new_n1142), .A2(new_n941), .ZN(new_n1148));
  NAND3_X1  g0948(.A1(new_n1148), .A2(new_n962), .A3(new_n951), .ZN(new_n1149));
  NAND4_X1  g0949(.A1(new_n767), .A2(new_n941), .A3(new_n851), .A4(G330), .ZN(new_n1150));
  NAND3_X1  g0950(.A1(new_n1147), .A2(new_n1149), .A3(new_n1150), .ZN(new_n1151));
  NAND2_X1  g0951(.A1(new_n1144), .A2(new_n1151), .ZN(new_n1152));
  INV_X1    g0952(.A(KEYINPUT116), .ZN(new_n1153));
  INV_X1    g0953(.A(new_n851), .ZN(new_n1154));
  OAI21_X1  g0954(.A(new_n965), .B1(new_n768), .B2(new_n1154), .ZN(new_n1155));
  NAND2_X1  g0955(.A1(new_n1155), .A2(new_n1135), .ZN(new_n1156));
  NAND2_X1  g0956(.A1(new_n1156), .A2(new_n1137), .ZN(new_n1157));
  AND2_X1   g0957(.A1(new_n934), .A2(G330), .ZN(new_n1158));
  AOI21_X1  g0958(.A(new_n941), .B1(new_n856), .B2(new_n1158), .ZN(new_n1159));
  NAND3_X1  g0959(.A1(new_n1141), .A2(new_n1150), .A3(new_n847), .ZN(new_n1160));
  OAI21_X1  g0960(.A(new_n1157), .B1(new_n1159), .B2(new_n1160), .ZN(new_n1161));
  NAND2_X1  g0961(.A1(new_n1158), .A2(new_n527), .ZN(new_n1162));
  AND3_X1   g0962(.A1(new_n651), .A2(new_n970), .A3(new_n1162), .ZN(new_n1163));
  AOI21_X1  g0963(.A(new_n1153), .B1(new_n1161), .B2(new_n1163), .ZN(new_n1164));
  NAND2_X1  g0964(.A1(new_n1152), .A2(new_n1164), .ZN(new_n1165));
  INV_X1    g0965(.A(new_n1159), .ZN(new_n1166));
  INV_X1    g0966(.A(new_n1160), .ZN(new_n1167));
  AOI22_X1  g0967(.A1(new_n1166), .A2(new_n1167), .B1(new_n1156), .B2(new_n1137), .ZN(new_n1168));
  NAND3_X1  g0968(.A1(new_n651), .A2(new_n970), .A3(new_n1162), .ZN(new_n1169));
  OAI21_X1  g0969(.A(KEYINPUT116), .B1(new_n1168), .B2(new_n1169), .ZN(new_n1170));
  NAND3_X1  g0970(.A1(new_n1170), .A2(new_n1151), .A3(new_n1144), .ZN(new_n1171));
  NAND3_X1  g0971(.A1(new_n1165), .A2(new_n1171), .A3(new_n728), .ZN(new_n1172));
  AOI21_X1  g0972(.A(new_n785), .B1(new_n960), .B2(new_n961), .ZN(new_n1173));
  OAI21_X1  g0973(.A(new_n351), .B1(new_n802), .B2(new_n202), .ZN(new_n1174));
  AOI21_X1  g0974(.A(new_n1174), .B1(G125), .B2(new_n809), .ZN(new_n1175));
  XOR2_X1   g0975(.A(new_n1175), .B(KEYINPUT117), .Z(new_n1176));
  INV_X1    g0976(.A(G128), .ZN(new_n1177));
  OAI22_X1  g0977(.A1(new_n1177), .A2(new_n820), .B1(new_n829), .B2(new_n873), .ZN(new_n1178));
  OR3_X1    g0978(.A1(new_n811), .A2(KEYINPUT53), .A3(new_n874), .ZN(new_n1179));
  OAI21_X1  g0979(.A(KEYINPUT53), .B1(new_n811), .B2(new_n874), .ZN(new_n1180));
  INV_X1    g0980(.A(G132), .ZN(new_n1181));
  OAI211_X1 g0981(.A(new_n1179), .B(new_n1180), .C1(new_n796), .C2(new_n1181), .ZN(new_n1182));
  XNOR2_X1  g0982(.A(KEYINPUT54), .B(G143), .ZN(new_n1183));
  OAI22_X1  g0983(.A1(new_n812), .A2(new_n1183), .B1(new_n509), .B2(new_n805), .ZN(new_n1184));
  NOR3_X1   g0984(.A1(new_n1178), .A2(new_n1182), .A3(new_n1184), .ZN(new_n1185));
  OAI22_X1  g0985(.A1(new_n796), .A2(new_n253), .B1(new_n355), .B2(new_n805), .ZN(new_n1186));
  OAI22_X1  g0986(.A1(new_n812), .A2(new_n205), .B1(new_n808), .B2(new_n806), .ZN(new_n1187));
  NOR2_X1   g0987(.A1(new_n1186), .A2(new_n1187), .ZN(new_n1188));
  AOI21_X1  g0988(.A(new_n351), .B1(new_n881), .B2(G87), .ZN(new_n1189));
  OAI211_X1 g0989(.A(new_n879), .B(new_n1189), .C1(new_n829), .C2(new_n206), .ZN(new_n1190));
  AOI21_X1  g0990(.A(new_n1190), .B1(G283), .B2(new_n815), .ZN(new_n1191));
  AOI22_X1  g0991(.A1(new_n1176), .A2(new_n1185), .B1(new_n1188), .B2(new_n1191), .ZN(new_n1192));
  INV_X1    g0992(.A(new_n787), .ZN(new_n1193));
  OAI221_X1 g0993(.A(new_n774), .B1(new_n1081), .B2(new_n861), .C1(new_n1192), .C2(new_n1193), .ZN(new_n1194));
  NOR2_X1   g0994(.A1(new_n1173), .A2(new_n1194), .ZN(new_n1195));
  XNOR2_X1  g0995(.A(new_n1195), .B(KEYINPUT118), .ZN(new_n1196));
  NAND3_X1  g0996(.A1(new_n1144), .A2(new_n1151), .A3(new_n773), .ZN(new_n1197));
  AND2_X1   g0997(.A1(new_n1196), .A2(new_n1197), .ZN(new_n1198));
  NAND2_X1  g0998(.A1(new_n1172), .A2(new_n1198), .ZN(G378));
  NOR2_X1   g0999(.A1(new_n904), .A2(new_n349), .ZN(new_n1200));
  XNOR2_X1  g1000(.A(new_n1200), .B(KEYINPUT55), .ZN(new_n1201));
  OR2_X1    g1001(.A1(new_n383), .A2(new_n1201), .ZN(new_n1202));
  NAND2_X1  g1002(.A1(new_n383), .A2(new_n1201), .ZN(new_n1203));
  NAND2_X1  g1003(.A1(new_n1202), .A2(new_n1203), .ZN(new_n1204));
  XOR2_X1   g1004(.A(KEYINPUT122), .B(KEYINPUT56), .Z(new_n1205));
  INV_X1    g1005(.A(new_n1205), .ZN(new_n1206));
  NAND2_X1  g1006(.A1(new_n1204), .A2(new_n1206), .ZN(new_n1207));
  NAND3_X1  g1007(.A1(new_n1202), .A2(new_n1205), .A3(new_n1203), .ZN(new_n1208));
  NAND2_X1  g1008(.A1(new_n1207), .A2(new_n1208), .ZN(new_n1209));
  NAND4_X1  g1009(.A1(new_n946), .A2(new_n1209), .A3(G330), .A4(new_n952), .ZN(new_n1210));
  NAND3_X1  g1010(.A1(new_n934), .A2(new_n941), .A3(new_n851), .ZN(new_n1211));
  AOI21_X1  g1011(.A(new_n1211), .B1(new_n925), .B2(new_n930), .ZN(new_n1212));
  OAI211_X1 g1012(.A(new_n952), .B(G330), .C1(new_n1212), .C2(new_n944), .ZN(new_n1213));
  AND2_X1   g1013(.A1(new_n1207), .A2(new_n1208), .ZN(new_n1214));
  NAND2_X1  g1014(.A1(new_n1213), .A2(new_n1214), .ZN(new_n1215));
  NAND2_X1  g1015(.A1(new_n1210), .A2(new_n1215), .ZN(new_n1216));
  INV_X1    g1016(.A(new_n969), .ZN(new_n1217));
  NAND2_X1  g1017(.A1(new_n1216), .A2(new_n1217), .ZN(new_n1218));
  NAND3_X1  g1018(.A1(new_n969), .A2(new_n1210), .A3(new_n1215), .ZN(new_n1219));
  NAND2_X1  g1019(.A1(new_n1218), .A2(new_n1219), .ZN(new_n1220));
  NAND2_X1  g1020(.A1(new_n1214), .A2(new_n784), .ZN(new_n1221));
  OAI21_X1  g1021(.A(new_n774), .B1(G50), .B2(new_n861), .ZN(new_n1222));
  NAND2_X1  g1022(.A1(new_n878), .A2(G58), .ZN(new_n1223));
  AND2_X1   g1023(.A1(new_n1223), .A2(new_n993), .ZN(new_n1224));
  OAI221_X1 g1024(.A(new_n1224), .B1(new_n205), .B2(new_n829), .C1(new_n253), .C2(new_n820), .ZN(new_n1225));
  NAND3_X1  g1025(.A1(new_n880), .A2(new_n1076), .A3(new_n358), .ZN(new_n1226));
  NOR2_X1   g1026(.A1(new_n1226), .A2(KEYINPUT119), .ZN(new_n1227));
  AOI22_X1  g1027(.A1(G107), .A2(new_n797), .B1(new_n818), .B2(new_n432), .ZN(new_n1228));
  NAND2_X1  g1028(.A1(new_n1226), .A2(KEYINPUT119), .ZN(new_n1229));
  OAI211_X1 g1029(.A(new_n1228), .B(new_n1229), .C1(new_n803), .C2(new_n808), .ZN(new_n1230));
  NOR3_X1   g1030(.A1(new_n1225), .A2(new_n1227), .A3(new_n1230), .ZN(new_n1231));
  NOR2_X1   g1031(.A1(new_n1231), .A2(KEYINPUT58), .ZN(new_n1232));
  NAND2_X1  g1032(.A1(new_n880), .A2(new_n358), .ZN(new_n1233));
  NOR2_X1   g1033(.A1(G33), .A2(G41), .ZN(new_n1234));
  NOR2_X1   g1034(.A1(new_n1234), .A2(G50), .ZN(new_n1235));
  AOI21_X1  g1035(.A(new_n1232), .B1(new_n1233), .B2(new_n1235), .ZN(new_n1236));
  OR2_X1    g1036(.A1(new_n1236), .A2(KEYINPUT120), .ZN(new_n1237));
  NAND2_X1  g1037(.A1(new_n1236), .A2(KEYINPUT120), .ZN(new_n1238));
  NOR2_X1   g1038(.A1(new_n811), .A2(new_n1183), .ZN(new_n1239));
  XNOR2_X1  g1039(.A(new_n1239), .B(KEYINPUT121), .ZN(new_n1240));
  AOI21_X1  g1040(.A(new_n1240), .B1(G150), .B2(new_n883), .ZN(new_n1241));
  AOI22_X1  g1041(.A1(G128), .A2(new_n797), .B1(new_n818), .B2(G137), .ZN(new_n1242));
  AOI22_X1  g1042(.A1(G125), .A2(new_n815), .B1(new_n792), .B2(G132), .ZN(new_n1243));
  NAND3_X1  g1043(.A1(new_n1241), .A2(new_n1242), .A3(new_n1243), .ZN(new_n1244));
  OR2_X1    g1044(.A1(new_n1244), .A2(KEYINPUT59), .ZN(new_n1245));
  INV_X1    g1045(.A(G124), .ZN(new_n1246));
  OAI221_X1 g1046(.A(new_n1234), .B1(new_n808), .B2(new_n1246), .C1(new_n509), .C2(new_n802), .ZN(new_n1247));
  AOI21_X1  g1047(.A(new_n1247), .B1(new_n1244), .B2(KEYINPUT59), .ZN(new_n1248));
  AOI22_X1  g1048(.A1(new_n1231), .A2(KEYINPUT58), .B1(new_n1245), .B2(new_n1248), .ZN(new_n1249));
  NAND3_X1  g1049(.A1(new_n1237), .A2(new_n1238), .A3(new_n1249), .ZN(new_n1250));
  AOI21_X1  g1050(.A(new_n1222), .B1(new_n1250), .B2(new_n787), .ZN(new_n1251));
  AOI22_X1  g1051(.A1(new_n1220), .A2(new_n773), .B1(new_n1221), .B2(new_n1251), .ZN(new_n1252));
  AND3_X1   g1052(.A1(new_n969), .A2(new_n1210), .A3(new_n1215), .ZN(new_n1253));
  AOI21_X1  g1053(.A(new_n969), .B1(new_n1210), .B2(new_n1215), .ZN(new_n1254));
  OAI21_X1  g1054(.A(KEYINPUT57), .B1(new_n1253), .B2(new_n1254), .ZN(new_n1255));
  NAND3_X1  g1055(.A1(new_n1144), .A2(new_n1151), .A3(new_n1161), .ZN(new_n1256));
  AND2_X1   g1056(.A1(new_n1256), .A2(new_n1163), .ZN(new_n1257));
  OAI21_X1  g1057(.A(new_n728), .B1(new_n1255), .B2(new_n1257), .ZN(new_n1258));
  NAND2_X1  g1058(.A1(new_n1256), .A2(new_n1163), .ZN(new_n1259));
  AOI21_X1  g1059(.A(KEYINPUT57), .B1(new_n1220), .B2(new_n1259), .ZN(new_n1260));
  OAI21_X1  g1060(.A(new_n1252), .B1(new_n1258), .B2(new_n1260), .ZN(new_n1261));
  INV_X1    g1061(.A(KEYINPUT123), .ZN(new_n1262));
  NOR2_X1   g1062(.A1(new_n1261), .A2(new_n1262), .ZN(new_n1263));
  NAND2_X1  g1063(.A1(new_n1220), .A2(new_n1259), .ZN(new_n1264));
  INV_X1    g1064(.A(KEYINPUT57), .ZN(new_n1265));
  NAND2_X1  g1065(.A1(new_n1264), .A2(new_n1265), .ZN(new_n1266));
  AOI21_X1  g1066(.A(new_n1265), .B1(new_n1218), .B2(new_n1219), .ZN(new_n1267));
  AOI21_X1  g1067(.A(new_n1069), .B1(new_n1267), .B2(new_n1259), .ZN(new_n1268));
  NAND2_X1  g1068(.A1(new_n1266), .A2(new_n1268), .ZN(new_n1269));
  AOI21_X1  g1069(.A(KEYINPUT123), .B1(new_n1269), .B2(new_n1252), .ZN(new_n1270));
  NOR2_X1   g1070(.A1(new_n1263), .A2(new_n1270), .ZN(G375));
  NAND2_X1  g1071(.A1(new_n1161), .A2(new_n1163), .ZN(new_n1272));
  NAND2_X1  g1072(.A1(new_n1168), .A2(new_n1169), .ZN(new_n1273));
  XOR2_X1   g1073(.A(new_n1043), .B(KEYINPUT124), .Z(new_n1274));
  NAND3_X1  g1074(.A1(new_n1272), .A2(new_n1273), .A3(new_n1274), .ZN(new_n1275));
  NOR2_X1   g1075(.A1(new_n941), .A2(new_n785), .ZN(new_n1276));
  AOI211_X1 g1076(.A(new_n351), .B(new_n997), .C1(G97), .C2(new_n881), .ZN(new_n1277));
  OAI221_X1 g1077(.A(new_n1277), .B1(new_n806), .B2(new_n820), .C1(new_n261), .C2(new_n829), .ZN(new_n1278));
  AOI22_X1  g1078(.A1(new_n818), .A2(G107), .B1(new_n809), .B2(G303), .ZN(new_n1279));
  OAI221_X1 g1079(.A(new_n1279), .B1(new_n803), .B2(new_n796), .C1(new_n431), .C2(new_n805), .ZN(new_n1280));
  AOI22_X1  g1080(.A1(new_n818), .A2(G150), .B1(G50), .B2(new_n883), .ZN(new_n1281));
  OAI221_X1 g1081(.A(new_n1281), .B1(new_n1177), .B2(new_n808), .C1(new_n873), .C2(new_n796), .ZN(new_n1282));
  OAI21_X1  g1082(.A(new_n778), .B1(new_n509), .B2(new_n811), .ZN(new_n1283));
  AOI21_X1  g1083(.A(new_n1283), .B1(new_n878), .B2(G58), .ZN(new_n1284));
  OAI221_X1 g1084(.A(new_n1284), .B1(new_n829), .B2(new_n1183), .C1(new_n1181), .C2(new_n820), .ZN(new_n1285));
  OAI22_X1  g1085(.A1(new_n1278), .A2(new_n1280), .B1(new_n1282), .B2(new_n1285), .ZN(new_n1286));
  NAND2_X1  g1086(.A1(new_n1286), .A2(new_n787), .ZN(new_n1287));
  OAI211_X1 g1087(.A(new_n1287), .B(new_n774), .C1(G68), .C2(new_n861), .ZN(new_n1288));
  OAI22_X1  g1088(.A1(new_n1168), .A2(new_n1010), .B1(new_n1276), .B2(new_n1288), .ZN(new_n1289));
  INV_X1    g1089(.A(new_n1289), .ZN(new_n1290));
  NAND2_X1  g1090(.A1(new_n1275), .A2(new_n1290), .ZN(G381));
  NAND4_X1  g1091(.A1(new_n1074), .A2(new_n836), .A3(new_n839), .A4(new_n1107), .ZN(new_n1292));
  OR4_X1    g1092(.A1(G384), .A2(G390), .A3(G381), .A4(new_n1292), .ZN(new_n1293));
  OR4_X1    g1093(.A1(G387), .A2(G375), .A3(G378), .A4(new_n1293), .ZN(G407));
  AND2_X1   g1094(.A1(new_n1172), .A2(new_n1198), .ZN(new_n1295));
  OAI21_X1  g1095(.A(new_n1295), .B1(new_n1263), .B2(new_n1270), .ZN(new_n1296));
  OAI211_X1 g1096(.A(G407), .B(G213), .C1(G343), .C2(new_n1296), .ZN(G409));
  NAND2_X1  g1097(.A1(G393), .A2(G396), .ZN(new_n1298));
  NAND2_X1  g1098(.A1(new_n1298), .A2(new_n1292), .ZN(new_n1299));
  NAND2_X1  g1099(.A1(G390), .A2(new_n1063), .ZN(new_n1300));
  NAND2_X1  g1100(.A1(new_n1109), .A2(new_n1127), .ZN(new_n1301));
  INV_X1    g1101(.A(new_n1133), .ZN(new_n1302));
  AOI21_X1  g1102(.A(new_n1301), .B1(new_n1302), .B2(new_n1131), .ZN(new_n1303));
  NAND2_X1  g1103(.A1(new_n1044), .A2(new_n1062), .ZN(new_n1304));
  NAND2_X1  g1104(.A1(new_n1304), .A2(new_n1008), .ZN(new_n1305));
  NAND2_X1  g1105(.A1(new_n1303), .A2(new_n1305), .ZN(new_n1306));
  AOI21_X1  g1106(.A(new_n1299), .B1(new_n1300), .B2(new_n1306), .ZN(new_n1307));
  NOR3_X1   g1107(.A1(new_n1065), .A2(new_n1066), .A3(G390), .ZN(new_n1308));
  NAND2_X1  g1108(.A1(new_n1308), .A2(KEYINPUT126), .ZN(new_n1309));
  OAI21_X1  g1109(.A(new_n1299), .B1(new_n1303), .B2(new_n1305), .ZN(new_n1310));
  NAND2_X1  g1110(.A1(new_n1305), .A2(KEYINPUT112), .ZN(new_n1311));
  NAND2_X1  g1111(.A1(new_n1063), .A2(new_n1064), .ZN(new_n1312));
  NAND3_X1  g1112(.A1(new_n1311), .A2(new_n1312), .A3(new_n1303), .ZN(new_n1313));
  INV_X1    g1113(.A(KEYINPUT126), .ZN(new_n1314));
  AOI21_X1  g1114(.A(new_n1310), .B1(new_n1313), .B2(new_n1314), .ZN(new_n1315));
  AOI21_X1  g1115(.A(new_n1307), .B1(new_n1309), .B2(new_n1315), .ZN(new_n1316));
  OAI211_X1 g1116(.A(G378), .B(new_n1252), .C1(new_n1258), .C2(new_n1260), .ZN(new_n1317));
  NAND3_X1  g1117(.A1(new_n1220), .A2(new_n1259), .A3(new_n1274), .ZN(new_n1318));
  NAND2_X1  g1118(.A1(new_n1252), .A2(new_n1318), .ZN(new_n1319));
  NAND2_X1  g1119(.A1(new_n1319), .A2(new_n1295), .ZN(new_n1320));
  NAND2_X1  g1120(.A1(new_n1317), .A2(new_n1320), .ZN(new_n1321));
  NOR2_X1   g1121(.A1(new_n698), .A2(G343), .ZN(new_n1322));
  INV_X1    g1122(.A(new_n1322), .ZN(new_n1323));
  NAND3_X1  g1123(.A1(new_n1168), .A2(KEYINPUT60), .A3(new_n1169), .ZN(new_n1324));
  NAND2_X1  g1124(.A1(new_n1324), .A2(new_n728), .ZN(new_n1325));
  NAND2_X1  g1125(.A1(new_n1272), .A2(KEYINPUT60), .ZN(new_n1326));
  AOI21_X1  g1126(.A(new_n1325), .B1(new_n1273), .B2(new_n1326), .ZN(new_n1327));
  OAI211_X1 g1127(.A(new_n859), .B(new_n889), .C1(new_n1327), .C2(new_n1289), .ZN(new_n1328));
  AND2_X1   g1128(.A1(new_n1326), .A2(new_n1273), .ZN(new_n1329));
  OAI211_X1 g1129(.A(G384), .B(new_n1290), .C1(new_n1329), .C2(new_n1325), .ZN(new_n1330));
  NAND2_X1  g1130(.A1(new_n1328), .A2(new_n1330), .ZN(new_n1331));
  INV_X1    g1131(.A(new_n1331), .ZN(new_n1332));
  NAND3_X1  g1132(.A1(new_n1321), .A2(new_n1323), .A3(new_n1332), .ZN(new_n1333));
  INV_X1    g1133(.A(KEYINPUT125), .ZN(new_n1334));
  NAND2_X1  g1134(.A1(new_n1333), .A2(new_n1334), .ZN(new_n1335));
  NAND4_X1  g1135(.A1(new_n1321), .A2(KEYINPUT125), .A3(new_n1323), .A4(new_n1332), .ZN(new_n1336));
  AOI21_X1  g1136(.A(KEYINPUT62), .B1(new_n1335), .B2(new_n1336), .ZN(new_n1337));
  NAND2_X1  g1137(.A1(new_n1321), .A2(new_n1323), .ZN(new_n1338));
  NAND2_X1  g1138(.A1(new_n1322), .A2(G2897), .ZN(new_n1339));
  AND3_X1   g1139(.A1(new_n1328), .A2(new_n1330), .A3(new_n1339), .ZN(new_n1340));
  AOI21_X1  g1140(.A(new_n1339), .B1(new_n1328), .B2(new_n1330), .ZN(new_n1341));
  NOR2_X1   g1141(.A1(new_n1340), .A2(new_n1341), .ZN(new_n1342));
  AOI21_X1  g1142(.A(KEYINPUT61), .B1(new_n1338), .B2(new_n1342), .ZN(new_n1343));
  NAND2_X1  g1143(.A1(new_n1333), .A2(KEYINPUT62), .ZN(new_n1344));
  NAND2_X1  g1144(.A1(new_n1343), .A2(new_n1344), .ZN(new_n1345));
  OAI21_X1  g1145(.A(new_n1316), .B1(new_n1337), .B2(new_n1345), .ZN(new_n1346));
  INV_X1    g1146(.A(KEYINPUT63), .ZN(new_n1347));
  NAND3_X1  g1147(.A1(new_n1335), .A2(new_n1347), .A3(new_n1336), .ZN(new_n1348));
  INV_X1    g1148(.A(new_n1307), .ZN(new_n1349));
  INV_X1    g1149(.A(new_n1310), .ZN(new_n1350));
  OAI21_X1  g1150(.A(new_n1350), .B1(new_n1308), .B2(KEYINPUT126), .ZN(new_n1351));
  NOR2_X1   g1151(.A1(new_n1313), .A2(new_n1314), .ZN(new_n1352));
  OAI21_X1  g1152(.A(new_n1349), .B1(new_n1351), .B2(new_n1352), .ZN(new_n1353));
  OR2_X1    g1153(.A1(new_n1333), .A2(new_n1347), .ZN(new_n1354));
  NAND4_X1  g1154(.A1(new_n1348), .A2(new_n1353), .A3(new_n1343), .A4(new_n1354), .ZN(new_n1355));
  NAND2_X1  g1155(.A1(new_n1346), .A2(new_n1355), .ZN(G405));
  NAND2_X1  g1156(.A1(new_n1353), .A2(KEYINPUT127), .ZN(new_n1357));
  NAND2_X1  g1157(.A1(new_n1220), .A2(new_n773), .ZN(new_n1358));
  NAND2_X1  g1158(.A1(new_n1221), .A2(new_n1251), .ZN(new_n1359));
  NAND2_X1  g1159(.A1(new_n1358), .A2(new_n1359), .ZN(new_n1360));
  AOI21_X1  g1160(.A(new_n1360), .B1(new_n1266), .B2(new_n1268), .ZN(new_n1361));
  NOR2_X1   g1161(.A1(new_n1361), .A2(new_n1295), .ZN(new_n1362));
  INV_X1    g1162(.A(new_n1362), .ZN(new_n1363));
  NAND3_X1  g1163(.A1(new_n1296), .A2(new_n1331), .A3(new_n1363), .ZN(new_n1364));
  INV_X1    g1164(.A(KEYINPUT127), .ZN(new_n1365));
  NAND2_X1  g1165(.A1(new_n1316), .A2(new_n1365), .ZN(new_n1366));
  NAND2_X1  g1166(.A1(new_n1361), .A2(KEYINPUT123), .ZN(new_n1367));
  NAND2_X1  g1167(.A1(new_n1261), .A2(new_n1262), .ZN(new_n1368));
  AOI21_X1  g1168(.A(G378), .B1(new_n1367), .B2(new_n1368), .ZN(new_n1369));
  OAI21_X1  g1169(.A(new_n1332), .B1(new_n1369), .B2(new_n1362), .ZN(new_n1370));
  NAND4_X1  g1170(.A1(new_n1357), .A2(new_n1364), .A3(new_n1366), .A4(new_n1370), .ZN(new_n1371));
  NOR3_X1   g1171(.A1(new_n1369), .A2(new_n1332), .A3(new_n1362), .ZN(new_n1372));
  AOI21_X1  g1172(.A(new_n1331), .B1(new_n1296), .B2(new_n1363), .ZN(new_n1373));
  OAI211_X1 g1173(.A(KEYINPUT127), .B(new_n1353), .C1(new_n1372), .C2(new_n1373), .ZN(new_n1374));
  NAND2_X1  g1174(.A1(new_n1371), .A2(new_n1374), .ZN(G402));
endmodule


