//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 0 0 0 0 1 1 1 1 1 1 1 1 0 0 0 0 1 1 0 1 0 1 1 1 1 1 0 1 0 0 0 0 1 1 0 0 0 0 0 1 1 0 1 0 0 1 0 0 1 0 0 0 1 0 1 1 1 0 1 1 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:41:05 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n204, new_n205, new_n206, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1033, new_n1034,
    new_n1035, new_n1036, new_n1037, new_n1038, new_n1039, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1122, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1187,
    new_n1188, new_n1189, new_n1190, new_n1191, new_n1192, new_n1193,
    new_n1194, new_n1195, new_n1196, new_n1197, new_n1198, new_n1199,
    new_n1200, new_n1201, new_n1202, new_n1203, new_n1204, new_n1205,
    new_n1206, new_n1207, new_n1208, new_n1210, new_n1211, new_n1212,
    new_n1214, new_n1215, new_n1216, new_n1217, new_n1219, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1274, new_n1275,
    new_n1276;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(new_n201), .ZN(new_n202));
  NOR3_X1   g0002(.A1(new_n202), .A2(G50), .A3(G77), .ZN(G353));
  INV_X1    g0003(.A(G97), .ZN(new_n204));
  INV_X1    g0004(.A(G107), .ZN(new_n205));
  NAND2_X1  g0005(.A1(new_n204), .A2(new_n205), .ZN(new_n206));
  NAND2_X1  g0006(.A1(new_n206), .A2(G87), .ZN(G355));
  INV_X1    g0007(.A(G1), .ZN(new_n208));
  INV_X1    g0008(.A(G20), .ZN(new_n209));
  NOR2_X1   g0009(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  INV_X1    g0010(.A(new_n210), .ZN(new_n211));
  NOR2_X1   g0011(.A1(new_n211), .A2(G13), .ZN(new_n212));
  OAI211_X1 g0012(.A(new_n212), .B(G250), .C1(G257), .C2(G264), .ZN(new_n213));
  XNOR2_X1  g0013(.A(new_n213), .B(KEYINPUT64), .ZN(new_n214));
  XNOR2_X1  g0014(.A(new_n214), .B(KEYINPUT0), .ZN(new_n215));
  NAND2_X1  g0015(.A1(new_n202), .A2(G50), .ZN(new_n216));
  INV_X1    g0016(.A(new_n216), .ZN(new_n217));
  NAND2_X1  g0017(.A1(G1), .A2(G13), .ZN(new_n218));
  NOR2_X1   g0018(.A1(new_n218), .A2(new_n209), .ZN(new_n219));
  NAND2_X1  g0019(.A1(new_n217), .A2(new_n219), .ZN(new_n220));
  AOI22_X1  g0020(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n221));
  XNOR2_X1  g0021(.A(new_n221), .B(KEYINPUT65), .ZN(new_n222));
  AOI22_X1  g0022(.A1(G58), .A2(G232), .B1(G116), .B2(G270), .ZN(new_n223));
  AOI22_X1  g0023(.A1(G50), .A2(G226), .B1(G68), .B2(G238), .ZN(new_n224));
  AOI22_X1  g0024(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n225));
  NAND3_X1  g0025(.A1(new_n223), .A2(new_n224), .A3(new_n225), .ZN(new_n226));
  OAI21_X1  g0026(.A(new_n211), .B1(new_n222), .B2(new_n226), .ZN(new_n227));
  OAI211_X1 g0027(.A(new_n215), .B(new_n220), .C1(KEYINPUT1), .C2(new_n227), .ZN(new_n228));
  NAND2_X1  g0028(.A1(new_n227), .A2(KEYINPUT1), .ZN(new_n229));
  XNOR2_X1  g0029(.A(new_n229), .B(KEYINPUT66), .ZN(new_n230));
  NOR2_X1   g0030(.A1(new_n228), .A2(new_n230), .ZN(G361));
  XNOR2_X1  g0031(.A(G250), .B(G257), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n232), .B(KEYINPUT67), .ZN(new_n233));
  XOR2_X1   g0033(.A(G264), .B(G270), .Z(new_n234));
  XNOR2_X1  g0034(.A(new_n233), .B(new_n234), .ZN(new_n235));
  XNOR2_X1  g0035(.A(G238), .B(G244), .ZN(new_n236));
  INV_X1    g0036(.A(G232), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XNOR2_X1  g0038(.A(KEYINPUT2), .B(G226), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n235), .B(new_n240), .ZN(G358));
  XNOR2_X1  g0041(.A(G50), .B(G68), .ZN(new_n242));
  XNOR2_X1  g0042(.A(G58), .B(G77), .ZN(new_n243));
  XOR2_X1   g0043(.A(new_n242), .B(new_n243), .Z(new_n244));
  XOR2_X1   g0044(.A(G87), .B(G97), .Z(new_n245));
  XNOR2_X1  g0045(.A(G107), .B(G116), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n245), .B(new_n246), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n244), .B(new_n247), .ZN(G351));
  INV_X1    g0048(.A(G41), .ZN(new_n249));
  INV_X1    g0049(.A(G45), .ZN(new_n250));
  AOI21_X1  g0050(.A(G1), .B1(new_n249), .B2(new_n250), .ZN(new_n251));
  NAND2_X1  g0051(.A1(G33), .A2(G41), .ZN(new_n252));
  NAND2_X1  g0052(.A1(new_n252), .A2(KEYINPUT68), .ZN(new_n253));
  INV_X1    g0053(.A(KEYINPUT68), .ZN(new_n254));
  NAND3_X1  g0054(.A1(new_n254), .A2(G33), .A3(G41), .ZN(new_n255));
  INV_X1    g0055(.A(new_n218), .ZN(new_n256));
  NAND3_X1  g0056(.A1(new_n253), .A2(new_n255), .A3(new_n256), .ZN(new_n257));
  INV_X1    g0057(.A(KEYINPUT69), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n257), .A2(new_n258), .ZN(new_n259));
  AOI21_X1  g0059(.A(new_n218), .B1(KEYINPUT68), .B2(new_n252), .ZN(new_n260));
  NAND3_X1  g0060(.A1(new_n260), .A2(KEYINPUT69), .A3(new_n255), .ZN(new_n261));
  AOI21_X1  g0061(.A(new_n251), .B1(new_n259), .B2(new_n261), .ZN(new_n262));
  INV_X1    g0062(.A(KEYINPUT77), .ZN(new_n263));
  OAI21_X1  g0063(.A(G238), .B1(new_n262), .B2(new_n263), .ZN(new_n264));
  INV_X1    g0064(.A(new_n251), .ZN(new_n265));
  AOI21_X1  g0065(.A(KEYINPUT69), .B1(new_n260), .B2(new_n255), .ZN(new_n266));
  AND4_X1   g0066(.A1(KEYINPUT69), .A2(new_n253), .A3(new_n255), .A4(new_n256), .ZN(new_n267));
  OAI21_X1  g0067(.A(new_n265), .B1(new_n266), .B2(new_n267), .ZN(new_n268));
  NOR2_X1   g0068(.A1(new_n268), .A2(KEYINPUT77), .ZN(new_n269));
  NOR2_X1   g0069(.A1(new_n264), .A2(new_n269), .ZN(new_n270));
  NAND2_X1  g0070(.A1(G33), .A2(G97), .ZN(new_n271));
  INV_X1    g0071(.A(new_n271), .ZN(new_n272));
  NOR2_X1   g0072(.A1(G226), .A2(G1698), .ZN(new_n273));
  AOI21_X1  g0073(.A(new_n273), .B1(new_n237), .B2(G1698), .ZN(new_n274));
  OR2_X1    g0074(.A1(KEYINPUT3), .A2(G33), .ZN(new_n275));
  NAND2_X1  g0075(.A1(KEYINPUT3), .A2(G33), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n275), .A2(new_n276), .ZN(new_n277));
  AOI21_X1  g0077(.A(new_n272), .B1(new_n274), .B2(new_n277), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n256), .A2(new_n252), .ZN(new_n279));
  OAI21_X1  g0079(.A(KEYINPUT75), .B1(new_n278), .B2(new_n279), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n237), .A2(G1698), .ZN(new_n281));
  OAI21_X1  g0081(.A(new_n281), .B1(G226), .B2(G1698), .ZN(new_n282));
  AND2_X1   g0082(.A1(KEYINPUT3), .A2(G33), .ZN(new_n283));
  NOR2_X1   g0083(.A1(KEYINPUT3), .A2(G33), .ZN(new_n284));
  NOR2_X1   g0084(.A1(new_n283), .A2(new_n284), .ZN(new_n285));
  OAI21_X1  g0085(.A(new_n271), .B1(new_n282), .B2(new_n285), .ZN(new_n286));
  INV_X1    g0086(.A(KEYINPUT75), .ZN(new_n287));
  INV_X1    g0087(.A(new_n279), .ZN(new_n288));
  NAND3_X1  g0088(.A1(new_n286), .A2(new_n287), .A3(new_n288), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n280), .A2(new_n289), .ZN(new_n290));
  INV_X1    g0090(.A(KEYINPUT76), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n259), .A2(new_n261), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n251), .A2(G274), .ZN(new_n293));
  INV_X1    g0093(.A(new_n293), .ZN(new_n294));
  AOI21_X1  g0094(.A(new_n291), .B1(new_n292), .B2(new_n294), .ZN(new_n295));
  AOI211_X1 g0095(.A(KEYINPUT76), .B(new_n293), .C1(new_n259), .C2(new_n261), .ZN(new_n296));
  OAI21_X1  g0096(.A(new_n290), .B1(new_n295), .B2(new_n296), .ZN(new_n297));
  NOR3_X1   g0097(.A1(new_n270), .A2(new_n297), .A3(KEYINPUT13), .ZN(new_n298));
  INV_X1    g0098(.A(KEYINPUT13), .ZN(new_n299));
  OAI21_X1  g0099(.A(new_n294), .B1(new_n266), .B2(new_n267), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n300), .A2(KEYINPUT76), .ZN(new_n301));
  NAND3_X1  g0101(.A1(new_n292), .A2(new_n291), .A3(new_n294), .ZN(new_n302));
  AOI22_X1  g0102(.A1(new_n301), .A2(new_n302), .B1(new_n280), .B2(new_n289), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n268), .A2(KEYINPUT77), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n262), .A2(new_n263), .ZN(new_n305));
  NAND3_X1  g0105(.A1(new_n304), .A2(new_n305), .A3(G238), .ZN(new_n306));
  AOI21_X1  g0106(.A(new_n299), .B1(new_n303), .B2(new_n306), .ZN(new_n307));
  OAI21_X1  g0107(.A(G169), .B1(new_n298), .B2(new_n307), .ZN(new_n308));
  INV_X1    g0108(.A(KEYINPUT78), .ZN(new_n309));
  NAND3_X1  g0109(.A1(new_n308), .A2(new_n309), .A3(KEYINPUT14), .ZN(new_n310));
  INV_X1    g0110(.A(G169), .ZN(new_n311));
  OAI21_X1  g0111(.A(KEYINPUT13), .B1(new_n270), .B2(new_n297), .ZN(new_n312));
  NAND3_X1  g0112(.A1(new_n303), .A2(new_n299), .A3(new_n306), .ZN(new_n313));
  AOI21_X1  g0113(.A(new_n311), .B1(new_n312), .B2(new_n313), .ZN(new_n314));
  INV_X1    g0114(.A(KEYINPUT14), .ZN(new_n315));
  OAI21_X1  g0115(.A(KEYINPUT78), .B1(new_n314), .B2(new_n315), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n314), .A2(new_n315), .ZN(new_n317));
  NAND3_X1  g0117(.A1(new_n312), .A2(G179), .A3(new_n313), .ZN(new_n318));
  NAND4_X1  g0118(.A1(new_n310), .A2(new_n316), .A3(new_n317), .A4(new_n318), .ZN(new_n319));
  NAND3_X1  g0119(.A1(new_n208), .A2(G13), .A3(G20), .ZN(new_n320));
  INV_X1    g0120(.A(new_n320), .ZN(new_n321));
  INV_X1    g0121(.A(G68), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n321), .A2(new_n322), .ZN(new_n323));
  XNOR2_X1  g0123(.A(new_n323), .B(KEYINPUT12), .ZN(new_n324));
  NOR2_X1   g0124(.A1(G20), .A2(G33), .ZN(new_n325));
  AOI22_X1  g0125(.A1(new_n325), .A2(G50), .B1(G20), .B2(new_n322), .ZN(new_n326));
  INV_X1    g0126(.A(G33), .ZN(new_n327));
  NOR2_X1   g0127(.A1(new_n327), .A2(G20), .ZN(new_n328));
  INV_X1    g0128(.A(new_n328), .ZN(new_n329));
  INV_X1    g0129(.A(G77), .ZN(new_n330));
  OAI21_X1  g0130(.A(new_n326), .B1(new_n329), .B2(new_n330), .ZN(new_n331));
  NAND3_X1  g0131(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n332), .A2(new_n218), .ZN(new_n333));
  NAND3_X1  g0133(.A1(new_n331), .A2(KEYINPUT11), .A3(new_n333), .ZN(new_n334));
  NOR2_X1   g0134(.A1(new_n321), .A2(new_n333), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n208), .A2(G20), .ZN(new_n336));
  NAND3_X1  g0136(.A1(new_n335), .A2(G68), .A3(new_n336), .ZN(new_n337));
  NAND3_X1  g0137(.A1(new_n324), .A2(new_n334), .A3(new_n337), .ZN(new_n338));
  AOI21_X1  g0138(.A(KEYINPUT11), .B1(new_n331), .B2(new_n333), .ZN(new_n339));
  OR3_X1    g0139(.A1(new_n338), .A2(KEYINPUT79), .A3(new_n339), .ZN(new_n340));
  OAI21_X1  g0140(.A(KEYINPUT79), .B1(new_n338), .B2(new_n339), .ZN(new_n341));
  AND2_X1   g0141(.A1(new_n340), .A2(new_n341), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n319), .A2(new_n342), .ZN(new_n343));
  NAND3_X1  g0143(.A1(new_n312), .A2(G190), .A3(new_n313), .ZN(new_n344));
  NOR2_X1   g0144(.A1(new_n338), .A2(new_n339), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n344), .A2(new_n345), .ZN(new_n346));
  INV_X1    g0146(.A(G200), .ZN(new_n347));
  AOI21_X1  g0147(.A(new_n347), .B1(new_n312), .B2(new_n313), .ZN(new_n348));
  NOR2_X1   g0148(.A1(new_n346), .A2(new_n348), .ZN(new_n349));
  INV_X1    g0149(.A(new_n349), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n343), .A2(new_n350), .ZN(new_n351));
  INV_X1    g0151(.A(new_n333), .ZN(new_n352));
  XNOR2_X1  g0152(.A(KEYINPUT8), .B(G58), .ZN(new_n353));
  INV_X1    g0153(.A(new_n353), .ZN(new_n354));
  AOI22_X1  g0154(.A1(new_n354), .A2(new_n328), .B1(G150), .B2(new_n325), .ZN(new_n355));
  OAI21_X1  g0155(.A(G20), .B1(new_n202), .B2(G50), .ZN(new_n356));
  AOI21_X1  g0156(.A(new_n352), .B1(new_n355), .B2(new_n356), .ZN(new_n357));
  NAND3_X1  g0157(.A1(new_n335), .A2(G50), .A3(new_n336), .ZN(new_n358));
  OAI21_X1  g0158(.A(new_n358), .B1(G50), .B2(new_n320), .ZN(new_n359));
  NOR2_X1   g0159(.A1(new_n357), .A2(new_n359), .ZN(new_n360));
  XNOR2_X1  g0160(.A(new_n360), .B(KEYINPUT9), .ZN(new_n361));
  INV_X1    g0161(.A(G1698), .ZN(new_n362));
  AOI21_X1  g0162(.A(new_n362), .B1(new_n275), .B2(new_n276), .ZN(new_n363));
  AOI22_X1  g0163(.A1(new_n363), .A2(G223), .B1(new_n285), .B2(G77), .ZN(new_n364));
  AOI21_X1  g0164(.A(G1698), .B1(new_n275), .B2(new_n276), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n365), .A2(G222), .ZN(new_n366));
  AOI21_X1  g0166(.A(new_n279), .B1(new_n364), .B2(new_n366), .ZN(new_n367));
  AOI21_X1  g0167(.A(new_n367), .B1(new_n292), .B2(new_n294), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n262), .A2(G226), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n368), .A2(new_n369), .ZN(new_n370));
  INV_X1    g0170(.A(KEYINPUT70), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n370), .A2(new_n371), .ZN(new_n372));
  NAND3_X1  g0172(.A1(new_n368), .A2(KEYINPUT70), .A3(new_n369), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n372), .A2(new_n373), .ZN(new_n374));
  AOI21_X1  g0174(.A(new_n361), .B1(new_n374), .B2(G190), .ZN(new_n375));
  INV_X1    g0175(.A(KEYINPUT74), .ZN(new_n376));
  AOI21_X1  g0176(.A(KEYINPUT10), .B1(new_n375), .B2(new_n376), .ZN(new_n377));
  NAND3_X1  g0177(.A1(new_n372), .A2(G200), .A3(new_n373), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n375), .A2(new_n378), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n377), .A2(new_n379), .ZN(new_n380));
  OAI211_X1 g0180(.A(new_n375), .B(new_n378), .C1(new_n376), .C2(KEYINPUT10), .ZN(new_n381));
  AND2_X1   g0181(.A1(KEYINPUT71), .A2(G179), .ZN(new_n382));
  NOR2_X1   g0182(.A1(KEYINPUT71), .A2(G179), .ZN(new_n383));
  NOR2_X1   g0183(.A1(new_n382), .A2(new_n383), .ZN(new_n384));
  NAND2_X1  g0184(.A1(new_n374), .A2(new_n384), .ZN(new_n385));
  INV_X1    g0185(.A(new_n360), .ZN(new_n386));
  OAI211_X1 g0186(.A(new_n385), .B(new_n386), .C1(G169), .C2(new_n374), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n209), .A2(new_n327), .ZN(new_n388));
  OAI22_X1  g0188(.A1(new_n353), .A2(new_n388), .B1(new_n209), .B2(new_n330), .ZN(new_n389));
  XNOR2_X1  g0189(.A(KEYINPUT15), .B(G87), .ZN(new_n390));
  INV_X1    g0190(.A(new_n390), .ZN(new_n391));
  AOI22_X1  g0191(.A1(new_n389), .A2(KEYINPUT72), .B1(new_n328), .B2(new_n391), .ZN(new_n392));
  OAI21_X1  g0192(.A(new_n392), .B1(KEYINPUT72), .B2(new_n389), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n393), .A2(new_n333), .ZN(new_n394));
  OR3_X1    g0194(.A1(new_n320), .A2(KEYINPUT73), .A3(G77), .ZN(new_n395));
  OAI21_X1  g0195(.A(KEYINPUT73), .B1(new_n320), .B2(G77), .ZN(new_n396));
  AOI21_X1  g0196(.A(new_n330), .B1(new_n208), .B2(G20), .ZN(new_n397));
  AOI22_X1  g0197(.A1(new_n395), .A2(new_n396), .B1(new_n335), .B2(new_n397), .ZN(new_n398));
  AND2_X1   g0198(.A1(new_n394), .A2(new_n398), .ZN(new_n399));
  NOR2_X1   g0199(.A1(G232), .A2(G1698), .ZN(new_n400));
  NOR2_X1   g0200(.A1(new_n362), .A2(G238), .ZN(new_n401));
  OAI21_X1  g0201(.A(new_n277), .B1(new_n400), .B2(new_n401), .ZN(new_n402));
  OAI211_X1 g0202(.A(new_n402), .B(new_n288), .C1(G107), .C2(new_n277), .ZN(new_n403));
  INV_X1    g0203(.A(G244), .ZN(new_n404));
  OAI211_X1 g0204(.A(new_n300), .B(new_n403), .C1(new_n268), .C2(new_n404), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n405), .A2(G200), .ZN(new_n406));
  INV_X1    g0206(.A(G190), .ZN(new_n407));
  OAI211_X1 g0207(.A(new_n399), .B(new_n406), .C1(new_n407), .C2(new_n405), .ZN(new_n408));
  INV_X1    g0208(.A(new_n408), .ZN(new_n409));
  AOI22_X1  g0209(.A1(new_n394), .A2(new_n398), .B1(new_n405), .B2(new_n311), .ZN(new_n410));
  INV_X1    g0210(.A(new_n384), .ZN(new_n411));
  OR2_X1    g0211(.A1(new_n405), .A2(new_n411), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n410), .A2(new_n412), .ZN(new_n413));
  INV_X1    g0213(.A(new_n413), .ZN(new_n414));
  NOR2_X1   g0214(.A1(new_n409), .A2(new_n414), .ZN(new_n415));
  NAND4_X1  g0215(.A1(new_n380), .A2(new_n381), .A3(new_n387), .A4(new_n415), .ZN(new_n416));
  INV_X1    g0216(.A(KEYINPUT82), .ZN(new_n417));
  INV_X1    g0217(.A(new_n335), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n354), .A2(new_n336), .ZN(new_n419));
  OAI22_X1  g0219(.A1(new_n418), .A2(new_n419), .B1(new_n320), .B2(new_n354), .ZN(new_n420));
  INV_X1    g0220(.A(new_n420), .ZN(new_n421));
  INV_X1    g0221(.A(KEYINPUT80), .ZN(new_n422));
  INV_X1    g0222(.A(G159), .ZN(new_n423));
  OAI21_X1  g0223(.A(new_n422), .B1(new_n388), .B2(new_n423), .ZN(new_n424));
  NAND3_X1  g0224(.A1(new_n325), .A2(KEYINPUT80), .A3(G159), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n424), .A2(new_n425), .ZN(new_n426));
  INV_X1    g0226(.A(G58), .ZN(new_n427));
  NOR2_X1   g0227(.A1(new_n427), .A2(new_n322), .ZN(new_n428));
  OAI21_X1  g0228(.A(G20), .B1(new_n428), .B2(new_n201), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n426), .A2(new_n429), .ZN(new_n430));
  AOI21_X1  g0230(.A(KEYINPUT7), .B1(new_n285), .B2(new_n209), .ZN(new_n431));
  INV_X1    g0231(.A(KEYINPUT7), .ZN(new_n432));
  NOR4_X1   g0232(.A1(new_n283), .A2(new_n284), .A3(new_n432), .A4(G20), .ZN(new_n433));
  OAI21_X1  g0233(.A(G68), .B1(new_n431), .B2(new_n433), .ZN(new_n434));
  AOI21_X1  g0234(.A(new_n430), .B1(new_n434), .B2(KEYINPUT81), .ZN(new_n435));
  OAI21_X1  g0235(.A(new_n432), .B1(new_n277), .B2(G20), .ZN(new_n436));
  NAND3_X1  g0236(.A1(new_n285), .A2(KEYINPUT7), .A3(new_n209), .ZN(new_n437));
  AOI21_X1  g0237(.A(new_n322), .B1(new_n436), .B2(new_n437), .ZN(new_n438));
  INV_X1    g0238(.A(KEYINPUT81), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n438), .A2(new_n439), .ZN(new_n440));
  AOI21_X1  g0240(.A(KEYINPUT16), .B1(new_n435), .B2(new_n440), .ZN(new_n441));
  INV_X1    g0241(.A(new_n430), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n442), .A2(new_n434), .ZN(new_n443));
  INV_X1    g0243(.A(KEYINPUT16), .ZN(new_n444));
  OAI21_X1  g0244(.A(new_n333), .B1(new_n443), .B2(new_n444), .ZN(new_n445));
  OAI21_X1  g0245(.A(new_n421), .B1(new_n441), .B2(new_n445), .ZN(new_n446));
  OR2_X1    g0246(.A1(G223), .A2(G1698), .ZN(new_n447));
  OAI21_X1  g0247(.A(new_n447), .B1(G226), .B2(new_n362), .ZN(new_n448));
  INV_X1    g0248(.A(G87), .ZN(new_n449));
  OAI22_X1  g0249(.A1(new_n448), .A2(new_n285), .B1(new_n327), .B2(new_n449), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n450), .A2(new_n288), .ZN(new_n451));
  OAI211_X1 g0251(.A(new_n300), .B(new_n451), .C1(new_n268), .C2(new_n237), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n452), .A2(G200), .ZN(new_n453));
  OAI21_X1  g0253(.A(new_n453), .B1(new_n407), .B2(new_n452), .ZN(new_n454));
  OAI21_X1  g0254(.A(new_n417), .B1(new_n446), .B2(new_n454), .ZN(new_n455));
  OAI21_X1  g0255(.A(new_n442), .B1(new_n438), .B2(new_n439), .ZN(new_n456));
  NOR2_X1   g0256(.A1(new_n434), .A2(KEYINPUT81), .ZN(new_n457));
  OAI21_X1  g0257(.A(new_n444), .B1(new_n456), .B2(new_n457), .ZN(new_n458));
  NOR2_X1   g0258(.A1(new_n438), .A2(new_n430), .ZN(new_n459));
  AOI21_X1  g0259(.A(new_n352), .B1(new_n459), .B2(KEYINPUT16), .ZN(new_n460));
  AOI21_X1  g0260(.A(new_n420), .B1(new_n458), .B2(new_n460), .ZN(new_n461));
  AOI22_X1  g0261(.A1(new_n292), .A2(new_n294), .B1(new_n450), .B2(new_n288), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n262), .A2(G232), .ZN(new_n463));
  AND3_X1   g0263(.A1(new_n462), .A2(new_n463), .A3(G190), .ZN(new_n464));
  AOI21_X1  g0264(.A(new_n347), .B1(new_n462), .B2(new_n463), .ZN(new_n465));
  NOR2_X1   g0265(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  NAND3_X1  g0266(.A1(new_n461), .A2(KEYINPUT82), .A3(new_n466), .ZN(new_n467));
  NAND3_X1  g0267(.A1(new_n455), .A2(new_n467), .A3(KEYINPUT17), .ZN(new_n468));
  INV_X1    g0268(.A(KEYINPUT83), .ZN(new_n469));
  NOR2_X1   g0269(.A1(new_n446), .A2(new_n454), .ZN(new_n470));
  INV_X1    g0270(.A(KEYINPUT17), .ZN(new_n471));
  AOI21_X1  g0271(.A(new_n469), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  NAND2_X1  g0272(.A1(new_n468), .A2(new_n472), .ZN(new_n473));
  NAND4_X1  g0273(.A1(new_n455), .A2(new_n467), .A3(new_n469), .A4(KEYINPUT17), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n452), .A2(G169), .ZN(new_n475));
  OAI21_X1  g0275(.A(new_n475), .B1(new_n452), .B2(new_n384), .ZN(new_n476));
  INV_X1    g0276(.A(KEYINPUT18), .ZN(new_n477));
  NAND3_X1  g0277(.A1(new_n446), .A2(new_n476), .A3(new_n477), .ZN(new_n478));
  INV_X1    g0278(.A(new_n478), .ZN(new_n479));
  AOI21_X1  g0279(.A(new_n477), .B1(new_n446), .B2(new_n476), .ZN(new_n480));
  NOR2_X1   g0280(.A1(new_n479), .A2(new_n480), .ZN(new_n481));
  NAND3_X1  g0281(.A1(new_n473), .A2(new_n474), .A3(new_n481), .ZN(new_n482));
  NOR3_X1   g0282(.A1(new_n351), .A2(new_n416), .A3(new_n482), .ZN(new_n483));
  INV_X1    g0283(.A(KEYINPUT5), .ZN(new_n484));
  INV_X1    g0284(.A(KEYINPUT87), .ZN(new_n485));
  OAI21_X1  g0285(.A(new_n484), .B1(new_n485), .B2(G41), .ZN(new_n486));
  NAND3_X1  g0286(.A1(new_n249), .A2(KEYINPUT87), .A3(KEYINPUT5), .ZN(new_n487));
  NOR2_X1   g0287(.A1(new_n250), .A2(G1), .ZN(new_n488));
  AND3_X1   g0288(.A1(new_n486), .A2(new_n487), .A3(new_n488), .ZN(new_n489));
  AOI21_X1  g0289(.A(new_n489), .B1(new_n259), .B2(new_n261), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n490), .A2(G264), .ZN(new_n491));
  AND2_X1   g0291(.A1(new_n489), .A2(G274), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n492), .A2(new_n292), .ZN(new_n493));
  OAI211_X1 g0293(.A(G257), .B(G1698), .C1(new_n283), .C2(new_n284), .ZN(new_n494));
  OAI211_X1 g0294(.A(G250), .B(new_n362), .C1(new_n283), .C2(new_n284), .ZN(new_n495));
  INV_X1    g0295(.A(G294), .ZN(new_n496));
  OAI211_X1 g0296(.A(new_n494), .B(new_n495), .C1(new_n327), .C2(new_n496), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n497), .A2(new_n288), .ZN(new_n498));
  NAND4_X1  g0298(.A1(new_n491), .A2(new_n493), .A3(G179), .A4(new_n498), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n498), .A2(KEYINPUT97), .ZN(new_n500));
  INV_X1    g0300(.A(KEYINPUT97), .ZN(new_n501));
  NAND3_X1  g0301(.A1(new_n497), .A2(new_n501), .A3(new_n288), .ZN(new_n502));
  NAND4_X1  g0302(.A1(new_n500), .A2(new_n491), .A3(new_n493), .A4(new_n502), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n503), .A2(G169), .ZN(new_n504));
  NAND3_X1  g0304(.A1(new_n277), .A2(new_n209), .A3(G87), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n505), .A2(KEYINPUT22), .ZN(new_n506));
  INV_X1    g0306(.A(KEYINPUT22), .ZN(new_n507));
  NAND4_X1  g0307(.A1(new_n277), .A2(new_n507), .A3(new_n209), .A4(G87), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n506), .A2(new_n508), .ZN(new_n509));
  INV_X1    g0309(.A(KEYINPUT24), .ZN(new_n510));
  INV_X1    g0310(.A(G116), .ZN(new_n511));
  NOR3_X1   g0311(.A1(new_n327), .A2(new_n511), .A3(G20), .ZN(new_n512));
  INV_X1    g0312(.A(KEYINPUT23), .ZN(new_n513));
  OAI21_X1  g0313(.A(new_n513), .B1(new_n209), .B2(G107), .ZN(new_n514));
  NAND3_X1  g0314(.A1(new_n205), .A2(KEYINPUT23), .A3(G20), .ZN(new_n515));
  AOI21_X1  g0315(.A(new_n512), .B1(new_n514), .B2(new_n515), .ZN(new_n516));
  AND3_X1   g0316(.A1(new_n509), .A2(new_n510), .A3(new_n516), .ZN(new_n517));
  AOI21_X1  g0317(.A(new_n510), .B1(new_n509), .B2(new_n516), .ZN(new_n518));
  OAI21_X1  g0318(.A(new_n333), .B1(new_n517), .B2(new_n518), .ZN(new_n519));
  AOI21_X1  g0319(.A(KEYINPUT25), .B1(new_n321), .B2(new_n205), .ZN(new_n520));
  INV_X1    g0320(.A(new_n520), .ZN(new_n521));
  NAND3_X1  g0321(.A1(new_n321), .A2(KEYINPUT25), .A3(new_n205), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n208), .A2(G33), .ZN(new_n523));
  NAND4_X1  g0323(.A1(new_n320), .A2(new_n523), .A3(new_n218), .A4(new_n332), .ZN(new_n524));
  INV_X1    g0324(.A(new_n524), .ZN(new_n525));
  AOI22_X1  g0325(.A1(new_n521), .A2(new_n522), .B1(G107), .B2(new_n525), .ZN(new_n526));
  AOI22_X1  g0326(.A1(new_n499), .A2(new_n504), .B1(new_n519), .B2(new_n526), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n519), .A2(new_n526), .ZN(new_n528));
  INV_X1    g0328(.A(new_n528), .ZN(new_n529));
  INV_X1    g0329(.A(KEYINPUT98), .ZN(new_n530));
  OAI21_X1  g0330(.A(new_n530), .B1(new_n503), .B2(G190), .ZN(new_n531));
  AND2_X1   g0331(.A1(new_n491), .A2(new_n502), .ZN(new_n532));
  AOI22_X1  g0332(.A1(new_n498), .A2(KEYINPUT97), .B1(new_n492), .B2(new_n292), .ZN(new_n533));
  NAND4_X1  g0333(.A1(new_n532), .A2(KEYINPUT98), .A3(new_n407), .A4(new_n533), .ZN(new_n534));
  NAND3_X1  g0334(.A1(new_n491), .A2(new_n493), .A3(new_n498), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n535), .A2(new_n347), .ZN(new_n536));
  NAND3_X1  g0336(.A1(new_n531), .A2(new_n534), .A3(new_n536), .ZN(new_n537));
  AOI21_X1  g0337(.A(new_n527), .B1(new_n529), .B2(new_n537), .ZN(new_n538));
  OAI211_X1 g0338(.A(G264), .B(G1698), .C1(new_n283), .C2(new_n284), .ZN(new_n539));
  OAI211_X1 g0339(.A(G257), .B(new_n362), .C1(new_n283), .C2(new_n284), .ZN(new_n540));
  INV_X1    g0340(.A(G303), .ZN(new_n541));
  OAI211_X1 g0341(.A(new_n539), .B(new_n540), .C1(new_n541), .C2(new_n277), .ZN(new_n542));
  AOI22_X1  g0342(.A1(new_n492), .A2(new_n292), .B1(new_n542), .B2(new_n288), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n490), .A2(G270), .ZN(new_n544));
  AOI21_X1  g0344(.A(new_n311), .B1(new_n543), .B2(new_n544), .ZN(new_n545));
  AOI21_X1  g0345(.A(G20), .B1(new_n327), .B2(G97), .ZN(new_n546));
  AND3_X1   g0346(.A1(KEYINPUT86), .A2(G33), .A3(G283), .ZN(new_n547));
  AOI21_X1  g0347(.A(KEYINPUT86), .B1(G33), .B2(G283), .ZN(new_n548));
  OAI21_X1  g0348(.A(new_n546), .B1(new_n547), .B2(new_n548), .ZN(new_n549));
  AOI22_X1  g0349(.A1(new_n332), .A2(new_n218), .B1(G20), .B2(new_n511), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  INV_X1    g0351(.A(KEYINPUT20), .ZN(new_n552));
  OAI21_X1  g0352(.A(KEYINPUT95), .B1(new_n551), .B2(new_n552), .ZN(new_n553));
  INV_X1    g0353(.A(KEYINPUT95), .ZN(new_n554));
  NAND4_X1  g0354(.A1(new_n549), .A2(new_n554), .A3(KEYINPUT20), .A4(new_n550), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n551), .A2(new_n552), .ZN(new_n556));
  NAND3_X1  g0356(.A1(new_n553), .A2(new_n555), .A3(new_n556), .ZN(new_n557));
  NAND4_X1  g0357(.A1(new_n208), .A2(new_n511), .A3(G13), .A4(G20), .ZN(new_n558));
  XNOR2_X1  g0358(.A(new_n558), .B(KEYINPUT94), .ZN(new_n559));
  OR3_X1    g0359(.A1(new_n524), .A2(KEYINPUT93), .A3(new_n511), .ZN(new_n560));
  OAI21_X1  g0360(.A(KEYINPUT93), .B1(new_n524), .B2(new_n511), .ZN(new_n561));
  AOI21_X1  g0361(.A(new_n559), .B1(new_n560), .B2(new_n561), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n557), .A2(new_n562), .ZN(new_n563));
  AOI21_X1  g0363(.A(KEYINPUT96), .B1(new_n545), .B2(new_n563), .ZN(new_n564));
  INV_X1    g0364(.A(KEYINPUT21), .ZN(new_n565));
  INV_X1    g0365(.A(new_n563), .ZN(new_n566));
  NAND3_X1  g0366(.A1(new_n543), .A2(G179), .A3(new_n544), .ZN(new_n567));
  OAI22_X1  g0367(.A1(new_n564), .A2(new_n565), .B1(new_n566), .B2(new_n567), .ZN(new_n568));
  AOI21_X1  g0368(.A(new_n347), .B1(new_n543), .B2(new_n544), .ZN(new_n569));
  AND2_X1   g0369(.A1(new_n543), .A2(new_n544), .ZN(new_n570));
  AOI211_X1 g0370(.A(new_n563), .B(new_n569), .C1(G190), .C2(new_n570), .ZN(new_n571));
  AOI211_X1 g0371(.A(KEYINPUT96), .B(KEYINPUT21), .C1(new_n545), .C2(new_n563), .ZN(new_n572));
  NOR3_X1   g0372(.A1(new_n568), .A2(new_n571), .A3(new_n572), .ZN(new_n573));
  INV_X1    g0373(.A(KEYINPUT88), .ZN(new_n574));
  NAND4_X1  g0374(.A1(new_n277), .A2(KEYINPUT4), .A3(G244), .A4(new_n362), .ZN(new_n575));
  INV_X1    g0375(.A(KEYINPUT85), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n575), .A2(new_n576), .ZN(new_n577));
  NAND3_X1  g0377(.A1(new_n277), .A2(G244), .A3(new_n362), .ZN(new_n578));
  INV_X1    g0378(.A(KEYINPUT4), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  NAND4_X1  g0380(.A1(new_n365), .A2(KEYINPUT85), .A3(KEYINPUT4), .A4(G244), .ZN(new_n581));
  NOR2_X1   g0381(.A1(new_n547), .A2(new_n548), .ZN(new_n582));
  AOI21_X1  g0382(.A(new_n582), .B1(new_n363), .B2(G250), .ZN(new_n583));
  NAND4_X1  g0383(.A1(new_n577), .A2(new_n580), .A3(new_n581), .A4(new_n583), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n584), .A2(new_n288), .ZN(new_n585));
  AOI22_X1  g0385(.A1(new_n490), .A2(G257), .B1(new_n492), .B2(new_n292), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  OAI21_X1  g0387(.A(new_n574), .B1(new_n587), .B2(new_n407), .ZN(new_n588));
  XNOR2_X1  g0388(.A(KEYINPUT84), .B(KEYINPUT6), .ZN(new_n589));
  NAND2_X1  g0389(.A1(G97), .A2(G107), .ZN(new_n590));
  NAND3_X1  g0390(.A1(new_n589), .A2(new_n206), .A3(new_n590), .ZN(new_n591));
  NOR2_X1   g0391(.A1(new_n204), .A2(G107), .ZN(new_n592));
  OAI21_X1  g0392(.A(new_n591), .B1(new_n589), .B2(new_n592), .ZN(new_n593));
  OAI22_X1  g0393(.A1(new_n593), .A2(new_n209), .B1(new_n330), .B2(new_n388), .ZN(new_n594));
  AOI21_X1  g0394(.A(new_n205), .B1(new_n436), .B2(new_n437), .ZN(new_n595));
  OAI21_X1  g0395(.A(new_n333), .B1(new_n594), .B2(new_n595), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n321), .A2(new_n204), .ZN(new_n597));
  OAI21_X1  g0397(.A(new_n597), .B1(new_n524), .B2(new_n204), .ZN(new_n598));
  INV_X1    g0398(.A(new_n598), .ZN(new_n599));
  AND2_X1   g0399(.A1(new_n596), .A2(new_n599), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n587), .A2(G200), .ZN(new_n601));
  NAND4_X1  g0401(.A1(new_n585), .A2(new_n586), .A3(KEYINPUT88), .A4(G190), .ZN(new_n602));
  NAND4_X1  g0402(.A1(new_n588), .A2(new_n600), .A3(new_n601), .A4(new_n602), .ZN(new_n603));
  AOI22_X1  g0403(.A1(new_n587), .A2(new_n311), .B1(new_n596), .B2(new_n599), .ZN(new_n604));
  INV_X1    g0404(.A(KEYINPUT89), .ZN(new_n605));
  OAI21_X1  g0405(.A(new_n605), .B1(new_n587), .B2(new_n411), .ZN(new_n606));
  NAND4_X1  g0406(.A1(new_n585), .A2(new_n586), .A3(KEYINPUT89), .A4(new_n384), .ZN(new_n607));
  NAND3_X1  g0407(.A1(new_n604), .A2(new_n606), .A3(new_n607), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n603), .A2(new_n608), .ZN(new_n609));
  AOI22_X1  g0409(.A1(new_n365), .A2(G238), .B1(G33), .B2(G116), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n363), .A2(G244), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n612), .A2(new_n288), .ZN(new_n613));
  INV_X1    g0413(.A(KEYINPUT90), .ZN(new_n614));
  MUX2_X1   g0414(.A(G250), .B(G274), .S(new_n488), .Z(new_n615));
  AND3_X1   g0415(.A1(new_n292), .A2(new_n614), .A3(new_n615), .ZN(new_n616));
  AOI21_X1  g0416(.A(new_n614), .B1(new_n292), .B2(new_n615), .ZN(new_n617));
  OAI21_X1  g0417(.A(new_n613), .B1(new_n616), .B2(new_n617), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n618), .A2(new_n311), .ZN(new_n619));
  INV_X1    g0419(.A(new_n619), .ZN(new_n620));
  INV_X1    g0420(.A(KEYINPUT19), .ZN(new_n621));
  OAI21_X1  g0421(.A(new_n621), .B1(new_n329), .B2(new_n204), .ZN(new_n622));
  NAND3_X1  g0422(.A1(new_n277), .A2(new_n209), .A3(G68), .ZN(new_n623));
  OAI21_X1  g0423(.A(new_n209), .B1(new_n271), .B2(new_n621), .ZN(new_n624));
  OAI21_X1  g0424(.A(new_n624), .B1(G87), .B2(new_n206), .ZN(new_n625));
  NAND3_X1  g0425(.A1(new_n622), .A2(new_n623), .A3(new_n625), .ZN(new_n626));
  AOI22_X1  g0426(.A1(new_n626), .A2(new_n333), .B1(new_n321), .B2(new_n390), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n525), .A2(new_n391), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  INV_X1    g0429(.A(KEYINPUT91), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  OAI211_X1 g0431(.A(new_n613), .B(new_n384), .C1(new_n616), .C2(new_n617), .ZN(new_n632));
  NAND3_X1  g0432(.A1(new_n627), .A2(KEYINPUT91), .A3(new_n628), .ZN(new_n633));
  NAND3_X1  g0433(.A1(new_n631), .A2(new_n632), .A3(new_n633), .ZN(new_n634));
  NOR2_X1   g0434(.A1(new_n524), .A2(new_n449), .ZN(new_n635));
  XNOR2_X1  g0435(.A(new_n635), .B(KEYINPUT92), .ZN(new_n636));
  AND2_X1   g0436(.A1(new_n636), .A2(new_n627), .ZN(new_n637));
  OAI21_X1  g0437(.A(new_n637), .B1(new_n618), .B2(new_n407), .ZN(new_n638));
  INV_X1    g0438(.A(new_n617), .ZN(new_n639));
  NAND3_X1  g0439(.A1(new_n292), .A2(new_n615), .A3(new_n614), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  AOI21_X1  g0441(.A(new_n347), .B1(new_n641), .B2(new_n613), .ZN(new_n642));
  OAI22_X1  g0442(.A1(new_n620), .A2(new_n634), .B1(new_n638), .B2(new_n642), .ZN(new_n643));
  NOR2_X1   g0443(.A1(new_n609), .A2(new_n643), .ZN(new_n644));
  AND4_X1   g0444(.A1(new_n483), .A2(new_n538), .A3(new_n573), .A4(new_n644), .ZN(G372));
  NAND2_X1  g0445(.A1(new_n537), .A2(new_n529), .ZN(new_n646));
  NAND3_X1  g0446(.A1(new_n646), .A2(new_n608), .A3(new_n603), .ZN(new_n647));
  NOR3_X1   g0447(.A1(new_n568), .A2(new_n527), .A3(new_n572), .ZN(new_n648));
  INV_X1    g0448(.A(KEYINPUT99), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n619), .A2(new_n649), .ZN(new_n650));
  AND2_X1   g0450(.A1(new_n632), .A2(new_n629), .ZN(new_n651));
  NAND3_X1  g0451(.A1(new_n618), .A2(KEYINPUT99), .A3(new_n311), .ZN(new_n652));
  NAND3_X1  g0452(.A1(new_n650), .A2(new_n651), .A3(new_n652), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n618), .A2(G200), .ZN(new_n654));
  OAI211_X1 g0454(.A(new_n654), .B(new_n637), .C1(new_n407), .C2(new_n618), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n653), .A2(new_n655), .ZN(new_n656));
  NOR3_X1   g0456(.A1(new_n647), .A2(new_n648), .A3(new_n656), .ZN(new_n657));
  INV_X1    g0457(.A(new_n608), .ZN(new_n658));
  INV_X1    g0458(.A(KEYINPUT26), .ZN(new_n659));
  NAND4_X1  g0459(.A1(new_n658), .A2(new_n659), .A3(new_n655), .A4(new_n653), .ZN(new_n660));
  OAI21_X1  g0460(.A(KEYINPUT26), .B1(new_n643), .B2(new_n608), .ZN(new_n661));
  NAND3_X1  g0461(.A1(new_n660), .A2(new_n653), .A3(new_n661), .ZN(new_n662));
  OAI21_X1  g0462(.A(new_n483), .B1(new_n657), .B2(new_n662), .ZN(new_n663));
  INV_X1    g0463(.A(new_n387), .ZN(new_n664));
  INV_X1    g0464(.A(KEYINPUT100), .ZN(new_n665));
  OAI21_X1  g0465(.A(new_n665), .B1(new_n479), .B2(new_n480), .ZN(new_n666));
  INV_X1    g0466(.A(new_n480), .ZN(new_n667));
  NAND3_X1  g0467(.A1(new_n667), .A2(KEYINPUT100), .A3(new_n478), .ZN(new_n668));
  AND2_X1   g0468(.A1(new_n666), .A2(new_n668), .ZN(new_n669));
  AOI22_X1  g0469(.A1(new_n319), .A2(new_n342), .B1(new_n350), .B2(new_n414), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n473), .A2(new_n474), .ZN(new_n671));
  OAI21_X1  g0471(.A(new_n669), .B1(new_n670), .B2(new_n671), .ZN(new_n672));
  AND2_X1   g0472(.A1(new_n380), .A2(new_n381), .ZN(new_n673));
  AOI21_X1  g0473(.A(new_n664), .B1(new_n672), .B2(new_n673), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n663), .A2(new_n674), .ZN(G369));
  NAND3_X1  g0475(.A1(new_n208), .A2(new_n209), .A3(G13), .ZN(new_n676));
  OR2_X1    g0476(.A1(new_n676), .A2(KEYINPUT27), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n676), .A2(KEYINPUT27), .ZN(new_n678));
  NAND3_X1  g0478(.A1(new_n677), .A2(new_n678), .A3(G213), .ZN(new_n679));
  INV_X1    g0479(.A(new_n679), .ZN(new_n680));
  INV_X1    g0480(.A(KEYINPUT101), .ZN(new_n681));
  OR2_X1    g0481(.A1(new_n681), .A2(G343), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n681), .A2(G343), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n680), .A2(new_n684), .ZN(new_n685));
  INV_X1    g0485(.A(new_n685), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n563), .A2(new_n686), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n573), .A2(new_n687), .ZN(new_n688));
  NOR2_X1   g0488(.A1(new_n568), .A2(new_n572), .ZN(new_n689));
  OAI21_X1  g0489(.A(new_n688), .B1(new_n689), .B2(new_n687), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n690), .A2(G330), .ZN(new_n691));
  INV_X1    g0491(.A(new_n691), .ZN(new_n692));
  OAI21_X1  g0492(.A(new_n538), .B1(new_n529), .B2(new_n685), .ZN(new_n693));
  INV_X1    g0493(.A(new_n527), .ZN(new_n694));
  OAI21_X1  g0494(.A(new_n693), .B1(new_n694), .B2(new_n685), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n692), .A2(new_n695), .ZN(new_n696));
  NOR2_X1   g0496(.A1(new_n689), .A2(new_n686), .ZN(new_n697));
  AOI22_X1  g0497(.A1(new_n697), .A2(new_n538), .B1(new_n527), .B2(new_n685), .ZN(new_n698));
  NAND2_X1  g0498(.A1(new_n696), .A2(new_n698), .ZN(G399));
  NAND2_X1  g0499(.A1(new_n212), .A2(new_n249), .ZN(new_n700));
  NOR3_X1   g0500(.A1(new_n206), .A2(G87), .A3(G116), .ZN(new_n701));
  NAND3_X1  g0501(.A1(new_n700), .A2(G1), .A3(new_n701), .ZN(new_n702));
  OAI21_X1  g0502(.A(new_n702), .B1(new_n216), .B2(new_n700), .ZN(new_n703));
  XNOR2_X1  g0503(.A(new_n703), .B(KEYINPUT28), .ZN(new_n704));
  NAND4_X1  g0504(.A1(new_n644), .A2(new_n538), .A3(new_n573), .A4(new_n685), .ZN(new_n705));
  NAND2_X1  g0505(.A1(new_n491), .A2(new_n498), .ZN(new_n706));
  NOR2_X1   g0506(.A1(new_n567), .A2(new_n706), .ZN(new_n707));
  INV_X1    g0507(.A(new_n587), .ZN(new_n708));
  AOI22_X1  g0508(.A1(new_n639), .A2(new_n640), .B1(new_n288), .B2(new_n612), .ZN(new_n709));
  NAND3_X1  g0509(.A1(new_n707), .A2(new_n708), .A3(new_n709), .ZN(new_n710));
  INV_X1    g0510(.A(KEYINPUT30), .ZN(new_n711));
  NOR2_X1   g0511(.A1(new_n708), .A2(new_n709), .ZN(new_n712));
  AOI21_X1  g0512(.A(new_n411), .B1(new_n543), .B2(new_n544), .ZN(new_n713));
  AND2_X1   g0513(.A1(new_n713), .A2(new_n535), .ZN(new_n714));
  AOI22_X1  g0514(.A1(new_n710), .A2(new_n711), .B1(new_n712), .B2(new_n714), .ZN(new_n715));
  NAND4_X1  g0515(.A1(new_n707), .A2(new_n708), .A3(KEYINPUT30), .A4(new_n709), .ZN(new_n716));
  AOI21_X1  g0516(.A(new_n685), .B1(new_n715), .B2(new_n716), .ZN(new_n717));
  NAND2_X1  g0517(.A1(new_n717), .A2(KEYINPUT31), .ZN(new_n718));
  NAND2_X1  g0518(.A1(new_n710), .A2(new_n711), .ZN(new_n719));
  NAND2_X1  g0519(.A1(new_n712), .A2(new_n714), .ZN(new_n720));
  NAND3_X1  g0520(.A1(new_n719), .A2(new_n720), .A3(new_n716), .ZN(new_n721));
  NAND2_X1  g0521(.A1(new_n721), .A2(new_n686), .ZN(new_n722));
  INV_X1    g0522(.A(KEYINPUT31), .ZN(new_n723));
  NAND2_X1  g0523(.A1(new_n722), .A2(new_n723), .ZN(new_n724));
  NAND3_X1  g0524(.A1(new_n705), .A2(new_n718), .A3(new_n724), .ZN(new_n725));
  AND2_X1   g0525(.A1(new_n725), .A2(G330), .ZN(new_n726));
  OAI21_X1  g0526(.A(new_n685), .B1(new_n657), .B2(new_n662), .ZN(new_n727));
  INV_X1    g0527(.A(KEYINPUT29), .ZN(new_n728));
  NAND2_X1  g0528(.A1(new_n727), .A2(new_n728), .ZN(new_n729));
  AND2_X1   g0529(.A1(new_n653), .A2(new_n655), .ZN(new_n730));
  AND2_X1   g0530(.A1(new_n603), .A2(new_n608), .ZN(new_n731));
  NAND3_X1  g0531(.A1(new_n730), .A2(new_n731), .A3(new_n646), .ZN(new_n732));
  INV_X1    g0532(.A(new_n568), .ZN(new_n733));
  INV_X1    g0533(.A(new_n572), .ZN(new_n734));
  NAND3_X1  g0534(.A1(new_n733), .A2(new_n694), .A3(new_n734), .ZN(new_n735));
  INV_X1    g0535(.A(KEYINPUT102), .ZN(new_n736));
  NAND2_X1  g0536(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  NAND2_X1  g0537(.A1(new_n648), .A2(KEYINPUT102), .ZN(new_n738));
  AOI21_X1  g0538(.A(new_n732), .B1(new_n737), .B2(new_n738), .ZN(new_n739));
  OR3_X1    g0539(.A1(new_n643), .A2(KEYINPUT26), .A3(new_n608), .ZN(new_n740));
  OAI21_X1  g0540(.A(KEYINPUT26), .B1(new_n656), .B2(new_n608), .ZN(new_n741));
  NAND3_X1  g0541(.A1(new_n740), .A2(new_n741), .A3(new_n653), .ZN(new_n742));
  OAI211_X1 g0542(.A(KEYINPUT29), .B(new_n685), .C1(new_n739), .C2(new_n742), .ZN(new_n743));
  AOI21_X1  g0543(.A(new_n726), .B1(new_n729), .B2(new_n743), .ZN(new_n744));
  OAI21_X1  g0544(.A(new_n704), .B1(new_n744), .B2(G1), .ZN(G364));
  INV_X1    g0545(.A(new_n700), .ZN(new_n746));
  AND2_X1   g0546(.A1(new_n209), .A2(G13), .ZN(new_n747));
  AOI21_X1  g0547(.A(new_n208), .B1(new_n747), .B2(G45), .ZN(new_n748));
  INV_X1    g0548(.A(new_n748), .ZN(new_n749));
  NOR2_X1   g0549(.A1(new_n746), .A2(new_n749), .ZN(new_n750));
  NOR2_X1   g0550(.A1(new_n692), .A2(new_n750), .ZN(new_n751));
  OAI21_X1  g0551(.A(new_n751), .B1(G330), .B2(new_n690), .ZN(new_n752));
  NAND2_X1  g0552(.A1(new_n212), .A2(new_n277), .ZN(new_n753));
  INV_X1    g0553(.A(G355), .ZN(new_n754));
  OAI22_X1  g0554(.A1(new_n753), .A2(new_n754), .B1(G116), .B2(new_n212), .ZN(new_n755));
  OR2_X1    g0555(.A1(new_n244), .A2(new_n250), .ZN(new_n756));
  NAND2_X1  g0556(.A1(new_n212), .A2(new_n285), .ZN(new_n757));
  AOI21_X1  g0557(.A(new_n757), .B1(new_n250), .B2(new_n217), .ZN(new_n758));
  AOI21_X1  g0558(.A(new_n755), .B1(new_n756), .B2(new_n758), .ZN(new_n759));
  NOR2_X1   g0559(.A1(G13), .A2(G33), .ZN(new_n760));
  XNOR2_X1  g0560(.A(new_n760), .B(KEYINPUT103), .ZN(new_n761));
  NOR2_X1   g0561(.A1(new_n761), .A2(G20), .ZN(new_n762));
  AOI21_X1  g0562(.A(new_n218), .B1(G20), .B2(new_n311), .ZN(new_n763));
  NOR2_X1   g0563(.A1(new_n762), .A2(new_n763), .ZN(new_n764));
  INV_X1    g0564(.A(new_n764), .ZN(new_n765));
  OAI21_X1  g0565(.A(new_n750), .B1(new_n759), .B2(new_n765), .ZN(new_n766));
  NOR2_X1   g0566(.A1(new_n209), .A2(G190), .ZN(new_n767));
  NOR2_X1   g0567(.A1(G179), .A2(G200), .ZN(new_n768));
  NAND2_X1  g0568(.A1(new_n767), .A2(new_n768), .ZN(new_n769));
  NOR2_X1   g0569(.A1(new_n769), .A2(new_n423), .ZN(new_n770));
  XNOR2_X1  g0570(.A(new_n770), .B(KEYINPUT106), .ZN(new_n771));
  XNOR2_X1  g0571(.A(KEYINPUT105), .B(KEYINPUT32), .ZN(new_n772));
  XNOR2_X1  g0572(.A(new_n771), .B(new_n772), .ZN(new_n773));
  NOR2_X1   g0573(.A1(new_n209), .A2(new_n407), .ZN(new_n774));
  NAND3_X1  g0574(.A1(new_n411), .A2(new_n347), .A3(new_n774), .ZN(new_n775));
  XOR2_X1   g0575(.A(new_n775), .B(KEYINPUT104), .Z(new_n776));
  OAI21_X1  g0576(.A(new_n773), .B1(new_n427), .B2(new_n776), .ZN(new_n777));
  NOR2_X1   g0577(.A1(new_n347), .A2(G179), .ZN(new_n778));
  NAND2_X1  g0578(.A1(new_n774), .A2(new_n778), .ZN(new_n779));
  NOR2_X1   g0579(.A1(new_n779), .A2(new_n449), .ZN(new_n780));
  NOR2_X1   g0580(.A1(new_n780), .A2(new_n285), .ZN(new_n781));
  NOR2_X1   g0581(.A1(new_n781), .A2(KEYINPUT107), .ZN(new_n782));
  NOR2_X1   g0582(.A1(new_n209), .A2(new_n347), .ZN(new_n783));
  NAND3_X1  g0583(.A1(new_n411), .A2(G190), .A3(new_n783), .ZN(new_n784));
  INV_X1    g0584(.A(new_n784), .ZN(new_n785));
  AOI21_X1  g0585(.A(new_n782), .B1(G50), .B2(new_n785), .ZN(new_n786));
  NAND2_X1  g0586(.A1(new_n778), .A2(new_n767), .ZN(new_n787));
  NOR2_X1   g0587(.A1(new_n787), .A2(new_n205), .ZN(new_n788));
  NAND2_X1  g0588(.A1(new_n768), .A2(G190), .ZN(new_n789));
  NAND2_X1  g0589(.A1(new_n789), .A2(G20), .ZN(new_n790));
  INV_X1    g0590(.A(new_n790), .ZN(new_n791));
  NOR2_X1   g0591(.A1(new_n791), .A2(new_n204), .ZN(new_n792));
  NAND3_X1  g0592(.A1(new_n411), .A2(new_n347), .A3(new_n767), .ZN(new_n793));
  INV_X1    g0593(.A(new_n793), .ZN(new_n794));
  AOI211_X1 g0594(.A(new_n788), .B(new_n792), .C1(new_n794), .C2(G77), .ZN(new_n795));
  NAND3_X1  g0595(.A1(new_n411), .A2(new_n407), .A3(new_n783), .ZN(new_n796));
  INV_X1    g0596(.A(new_n796), .ZN(new_n797));
  AOI22_X1  g0597(.A1(new_n781), .A2(KEYINPUT107), .B1(new_n797), .B2(G68), .ZN(new_n798));
  NAND3_X1  g0598(.A1(new_n786), .A2(new_n795), .A3(new_n798), .ZN(new_n799));
  OR2_X1    g0599(.A1(new_n769), .A2(KEYINPUT108), .ZN(new_n800));
  NAND2_X1  g0600(.A1(new_n769), .A2(KEYINPUT108), .ZN(new_n801));
  NAND2_X1  g0601(.A1(new_n800), .A2(new_n801), .ZN(new_n802));
  INV_X1    g0602(.A(new_n802), .ZN(new_n803));
  INV_X1    g0603(.A(new_n787), .ZN(new_n804));
  AOI22_X1  g0604(.A1(new_n803), .A2(G329), .B1(G283), .B2(new_n804), .ZN(new_n805));
  XNOR2_X1  g0605(.A(new_n805), .B(KEYINPUT109), .ZN(new_n806));
  OAI221_X1 g0606(.A(new_n285), .B1(new_n779), .B2(new_n541), .C1(new_n791), .C2(new_n496), .ZN(new_n807));
  AOI21_X1  g0607(.A(new_n807), .B1(G311), .B2(new_n794), .ZN(new_n808));
  INV_X1    g0608(.A(new_n775), .ZN(new_n809));
  AOI22_X1  g0609(.A1(G322), .A2(new_n809), .B1(new_n785), .B2(G326), .ZN(new_n810));
  XOR2_X1   g0610(.A(KEYINPUT33), .B(G317), .Z(new_n811));
  OAI211_X1 g0611(.A(new_n808), .B(new_n810), .C1(new_n796), .C2(new_n811), .ZN(new_n812));
  OAI22_X1  g0612(.A1(new_n777), .A2(new_n799), .B1(new_n806), .B2(new_n812), .ZN(new_n813));
  AOI21_X1  g0613(.A(new_n766), .B1(new_n813), .B2(new_n763), .ZN(new_n814));
  INV_X1    g0614(.A(new_n762), .ZN(new_n815));
  OAI21_X1  g0615(.A(new_n814), .B1(new_n690), .B2(new_n815), .ZN(new_n816));
  AND2_X1   g0616(.A1(new_n752), .A2(new_n816), .ZN(new_n817));
  INV_X1    g0617(.A(new_n817), .ZN(G396));
  NOR2_X1   g0618(.A1(new_n399), .A2(new_n685), .ZN(new_n819));
  OAI21_X1  g0619(.A(new_n413), .B1(new_n409), .B2(new_n819), .ZN(new_n820));
  NAND2_X1  g0620(.A1(new_n414), .A2(new_n685), .ZN(new_n821));
  NAND2_X1  g0621(.A1(new_n820), .A2(new_n821), .ZN(new_n822));
  NAND2_X1  g0622(.A1(new_n727), .A2(new_n822), .ZN(new_n823));
  INV_X1    g0623(.A(new_n822), .ZN(new_n824));
  OAI211_X1 g0624(.A(new_n685), .B(new_n824), .C1(new_n657), .C2(new_n662), .ZN(new_n825));
  AOI21_X1  g0625(.A(new_n726), .B1(new_n823), .B2(new_n825), .ZN(new_n826));
  NOR2_X1   g0626(.A1(new_n826), .A2(new_n750), .ZN(new_n827));
  NAND3_X1  g0627(.A1(new_n726), .A2(new_n823), .A3(new_n825), .ZN(new_n828));
  NAND2_X1  g0628(.A1(new_n827), .A2(new_n828), .ZN(new_n829));
  NOR2_X1   g0629(.A1(new_n787), .A2(new_n322), .ZN(new_n830));
  INV_X1    g0630(.A(new_n779), .ZN(new_n831));
  AOI211_X1 g0631(.A(new_n285), .B(new_n830), .C1(G50), .C2(new_n831), .ZN(new_n832));
  OAI21_X1  g0632(.A(new_n832), .B1(new_n427), .B2(new_n791), .ZN(new_n833));
  AOI22_X1  g0633(.A1(G137), .A2(new_n785), .B1(new_n794), .B2(G159), .ZN(new_n834));
  INV_X1    g0634(.A(G150), .ZN(new_n835));
  INV_X1    g0635(.A(G143), .ZN(new_n836));
  OAI221_X1 g0636(.A(new_n834), .B1(new_n835), .B2(new_n796), .C1(new_n776), .C2(new_n836), .ZN(new_n837));
  XOR2_X1   g0637(.A(new_n837), .B(KEYINPUT34), .Z(new_n838));
  AOI211_X1 g0638(.A(new_n833), .B(new_n838), .C1(G132), .C2(new_n803), .ZN(new_n839));
  AOI22_X1  g0639(.A1(new_n803), .A2(G311), .B1(G294), .B2(new_n809), .ZN(new_n840));
  OAI21_X1  g0640(.A(new_n840), .B1(new_n541), .B2(new_n784), .ZN(new_n841));
  NOR2_X1   g0641(.A1(new_n787), .A2(new_n449), .ZN(new_n842));
  OAI21_X1  g0642(.A(new_n285), .B1(new_n779), .B2(new_n205), .ZN(new_n843));
  OR3_X1    g0643(.A1(new_n792), .A2(new_n842), .A3(new_n843), .ZN(new_n844));
  INV_X1    g0644(.A(G283), .ZN(new_n845));
  OAI22_X1  g0645(.A1(new_n511), .A2(new_n793), .B1(new_n796), .B2(new_n845), .ZN(new_n846));
  NOR3_X1   g0646(.A1(new_n841), .A2(new_n844), .A3(new_n846), .ZN(new_n847));
  OAI21_X1  g0647(.A(new_n763), .B1(new_n839), .B2(new_n847), .ZN(new_n848));
  INV_X1    g0648(.A(new_n750), .ZN(new_n849));
  NOR2_X1   g0649(.A1(new_n763), .A2(new_n760), .ZN(new_n850));
  AOI21_X1  g0650(.A(new_n849), .B1(new_n330), .B2(new_n850), .ZN(new_n851));
  OAI211_X1 g0651(.A(new_n848), .B(new_n851), .C1(new_n761), .C2(new_n824), .ZN(new_n852));
  AND2_X1   g0652(.A1(new_n829), .A2(new_n852), .ZN(new_n853));
  INV_X1    g0653(.A(new_n853), .ZN(G384));
  INV_X1    g0654(.A(KEYINPUT35), .ZN(new_n855));
  OAI211_X1 g0655(.A(G116), .B(new_n219), .C1(new_n593), .C2(new_n855), .ZN(new_n856));
  AOI21_X1  g0656(.A(new_n856), .B1(new_n855), .B2(new_n593), .ZN(new_n857));
  XNOR2_X1  g0657(.A(new_n857), .B(KEYINPUT36), .ZN(new_n858));
  OR3_X1    g0658(.A1(new_n216), .A2(new_n330), .A3(new_n428), .ZN(new_n859));
  INV_X1    g0659(.A(G50), .ZN(new_n860));
  NAND2_X1  g0660(.A1(new_n860), .A2(G68), .ZN(new_n861));
  AOI211_X1 g0661(.A(new_n208), .B(G13), .C1(new_n859), .C2(new_n861), .ZN(new_n862));
  NOR2_X1   g0662(.A1(new_n858), .A2(new_n862), .ZN(new_n863));
  NAND2_X1  g0663(.A1(new_n825), .A2(new_n821), .ZN(new_n864));
  NAND3_X1  g0664(.A1(new_n340), .A2(new_n341), .A3(new_n686), .ZN(new_n865));
  XNOR2_X1  g0665(.A(new_n865), .B(KEYINPUT110), .ZN(new_n866));
  AOI211_X1 g0666(.A(new_n349), .B(new_n866), .C1(new_n319), .C2(new_n342), .ZN(new_n867));
  INV_X1    g0667(.A(new_n866), .ZN(new_n868));
  AOI21_X1  g0668(.A(new_n868), .B1(new_n343), .B2(new_n350), .ZN(new_n869));
  OAI21_X1  g0669(.A(new_n864), .B1(new_n867), .B2(new_n869), .ZN(new_n870));
  INV_X1    g0670(.A(KEYINPUT38), .ZN(new_n871));
  NOR2_X1   g0671(.A1(new_n459), .A2(KEYINPUT16), .ZN(new_n872));
  OAI21_X1  g0672(.A(new_n421), .B1(new_n445), .B2(new_n872), .ZN(new_n873));
  OAI21_X1  g0673(.A(new_n873), .B1(new_n476), .B2(new_n680), .ZN(new_n874));
  NAND3_X1  g0674(.A1(new_n455), .A2(new_n467), .A3(new_n874), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n875), .A2(KEYINPUT37), .ZN(new_n876));
  AOI21_X1  g0676(.A(KEYINPUT37), .B1(new_n446), .B2(new_n476), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n446), .A2(new_n680), .ZN(new_n878));
  NAND4_X1  g0678(.A1(new_n455), .A2(new_n877), .A3(new_n467), .A4(new_n878), .ZN(new_n879));
  AND2_X1   g0679(.A1(new_n873), .A2(new_n680), .ZN(new_n880));
  AOI221_X4 g0680(.A(new_n871), .B1(new_n876), .B2(new_n879), .C1(new_n482), .C2(new_n880), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n482), .A2(new_n880), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n876), .A2(new_n879), .ZN(new_n883));
  AOI21_X1  g0683(.A(KEYINPUT38), .B1(new_n882), .B2(new_n883), .ZN(new_n884));
  NOR2_X1   g0684(.A1(new_n881), .A2(new_n884), .ZN(new_n885));
  NOR2_X1   g0685(.A1(new_n870), .A2(new_n885), .ZN(new_n886));
  NOR2_X1   g0686(.A1(new_n669), .A2(new_n680), .ZN(new_n887));
  NOR2_X1   g0687(.A1(new_n886), .A2(new_n887), .ZN(new_n888));
  NAND3_X1  g0688(.A1(new_n882), .A2(KEYINPUT38), .A3(new_n883), .ZN(new_n889));
  NAND4_X1  g0689(.A1(new_n473), .A2(new_n668), .A3(new_n666), .A4(new_n474), .ZN(new_n890));
  INV_X1    g0690(.A(new_n878), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n446), .A2(new_n476), .ZN(new_n892));
  XNOR2_X1  g0692(.A(new_n892), .B(KEYINPUT100), .ZN(new_n893));
  OAI21_X1  g0693(.A(new_n878), .B1(new_n446), .B2(new_n454), .ZN(new_n894));
  OAI21_X1  g0694(.A(KEYINPUT37), .B1(new_n893), .B2(new_n894), .ZN(new_n895));
  AOI22_X1  g0695(.A1(new_n890), .A2(new_n891), .B1(new_n895), .B2(new_n879), .ZN(new_n896));
  XOR2_X1   g0696(.A(KEYINPUT111), .B(KEYINPUT38), .Z(new_n897));
  INV_X1    g0697(.A(new_n897), .ZN(new_n898));
  OAI21_X1  g0698(.A(new_n889), .B1(new_n896), .B2(new_n898), .ZN(new_n899));
  INV_X1    g0699(.A(KEYINPUT39), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n899), .A2(new_n900), .ZN(new_n901));
  NAND3_X1  g0701(.A1(new_n319), .A2(new_n342), .A3(new_n685), .ZN(new_n902));
  INV_X1    g0702(.A(new_n902), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n882), .A2(new_n883), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n904), .A2(new_n871), .ZN(new_n905));
  NAND3_X1  g0705(.A1(new_n905), .A2(KEYINPUT39), .A3(new_n889), .ZN(new_n906));
  NAND3_X1  g0706(.A1(new_n901), .A2(new_n903), .A3(new_n906), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n888), .A2(new_n907), .ZN(new_n908));
  NAND3_X1  g0708(.A1(new_n483), .A2(new_n743), .A3(new_n729), .ZN(new_n909));
  AND2_X1   g0709(.A1(new_n909), .A2(new_n674), .ZN(new_n910));
  XOR2_X1   g0710(.A(new_n908), .B(new_n910), .Z(new_n911));
  INV_X1    g0711(.A(new_n911), .ZN(new_n912));
  XNOR2_X1  g0712(.A(KEYINPUT112), .B(KEYINPUT40), .ZN(new_n913));
  OAI21_X1  g0713(.A(KEYINPUT113), .B1(new_n717), .B2(KEYINPUT31), .ZN(new_n914));
  INV_X1    g0714(.A(KEYINPUT113), .ZN(new_n915));
  NAND3_X1  g0715(.A1(new_n722), .A2(new_n915), .A3(new_n723), .ZN(new_n916));
  NAND4_X1  g0716(.A1(new_n914), .A2(new_n705), .A3(new_n916), .A4(new_n718), .ZN(new_n917));
  OAI211_X1 g0717(.A(new_n824), .B(new_n917), .C1(new_n869), .C2(new_n867), .ZN(new_n918));
  OAI21_X1  g0718(.A(new_n913), .B1(new_n885), .B2(new_n918), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n351), .A2(new_n866), .ZN(new_n920));
  NAND3_X1  g0720(.A1(new_n343), .A2(new_n350), .A3(new_n868), .ZN(new_n921));
  AOI21_X1  g0721(.A(new_n822), .B1(new_n920), .B2(new_n921), .ZN(new_n922));
  NAND4_X1  g0722(.A1(new_n922), .A2(KEYINPUT40), .A3(new_n899), .A4(new_n917), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n919), .A2(new_n923), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n483), .A2(new_n917), .ZN(new_n925));
  OR2_X1    g0725(.A1(new_n924), .A2(new_n925), .ZN(new_n926));
  NAND2_X1  g0726(.A1(new_n926), .A2(G330), .ZN(new_n927));
  AOI21_X1  g0727(.A(new_n927), .B1(new_n924), .B2(new_n925), .ZN(new_n928));
  OAI22_X1  g0728(.A1(new_n912), .A2(new_n928), .B1(new_n208), .B2(new_n747), .ZN(new_n929));
  AND2_X1   g0729(.A1(new_n912), .A2(new_n928), .ZN(new_n930));
  OAI21_X1  g0730(.A(new_n863), .B1(new_n929), .B2(new_n930), .ZN(G367));
  AND3_X1   g0731(.A1(new_n235), .A2(new_n212), .A3(new_n285), .ZN(new_n932));
  OAI21_X1  g0732(.A(new_n764), .B1(new_n212), .B2(new_n390), .ZN(new_n933));
  INV_X1    g0733(.A(KEYINPUT115), .ZN(new_n934));
  OAI21_X1  g0734(.A(new_n934), .B1(new_n779), .B2(new_n511), .ZN(new_n935));
  AOI22_X1  g0735(.A1(new_n794), .A2(G283), .B1(KEYINPUT46), .B2(new_n935), .ZN(new_n936));
  OAI21_X1  g0736(.A(new_n936), .B1(KEYINPUT46), .B2(new_n935), .ZN(new_n937));
  INV_X1    g0737(.A(new_n769), .ZN(new_n938));
  AOI21_X1  g0738(.A(new_n277), .B1(new_n938), .B2(G317), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n804), .A2(G97), .ZN(new_n940));
  OAI211_X1 g0740(.A(new_n939), .B(new_n940), .C1(new_n205), .C2(new_n791), .ZN(new_n941));
  INV_X1    g0741(.A(G311), .ZN(new_n942));
  OAI22_X1  g0742(.A1(new_n496), .A2(new_n796), .B1(new_n784), .B2(new_n942), .ZN(new_n943));
  NOR3_X1   g0743(.A1(new_n937), .A2(new_n941), .A3(new_n943), .ZN(new_n944));
  OAI21_X1  g0744(.A(new_n944), .B1(new_n541), .B2(new_n776), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n790), .A2(G68), .ZN(new_n946));
  INV_X1    g0746(.A(G137), .ZN(new_n947));
  OAI221_X1 g0747(.A(new_n946), .B1(new_n427), .B2(new_n779), .C1(new_n947), .C2(new_n769), .ZN(new_n948));
  AOI21_X1  g0748(.A(new_n285), .B1(new_n804), .B2(G77), .ZN(new_n949));
  OAI22_X1  g0749(.A1(new_n949), .A2(KEYINPUT116), .B1(new_n784), .B2(new_n836), .ZN(new_n950));
  AOI211_X1 g0750(.A(new_n948), .B(new_n950), .C1(G159), .C2(new_n797), .ZN(new_n951));
  AOI22_X1  g0751(.A1(new_n809), .A2(G150), .B1(new_n949), .B2(KEYINPUT116), .ZN(new_n952));
  OAI211_X1 g0752(.A(new_n951), .B(new_n952), .C1(new_n860), .C2(new_n793), .ZN(new_n953));
  NAND2_X1  g0753(.A1(new_n945), .A2(new_n953), .ZN(new_n954));
  XOR2_X1   g0754(.A(new_n954), .B(KEYINPUT47), .Z(new_n955));
  INV_X1    g0755(.A(new_n763), .ZN(new_n956));
  OAI221_X1 g0756(.A(new_n750), .B1(new_n932), .B2(new_n933), .C1(new_n955), .C2(new_n956), .ZN(new_n957));
  XOR2_X1   g0757(.A(new_n957), .B(KEYINPUT117), .Z(new_n958));
  NOR2_X1   g0758(.A1(new_n637), .A2(new_n685), .ZN(new_n959));
  INV_X1    g0759(.A(new_n959), .ZN(new_n960));
  NAND2_X1  g0760(.A1(new_n730), .A2(new_n960), .ZN(new_n961));
  OAI21_X1  g0761(.A(new_n961), .B1(new_n653), .B2(new_n960), .ZN(new_n962));
  NOR2_X1   g0762(.A1(new_n962), .A2(new_n815), .ZN(new_n963));
  NOR2_X1   g0763(.A1(new_n958), .A2(new_n963), .ZN(new_n964));
  OAI21_X1  g0764(.A(new_n731), .B1(new_n600), .B2(new_n685), .ZN(new_n965));
  NAND2_X1  g0765(.A1(new_n658), .A2(new_n686), .ZN(new_n966));
  NAND2_X1  g0766(.A1(new_n965), .A2(new_n966), .ZN(new_n967));
  NOR2_X1   g0767(.A1(new_n698), .A2(new_n967), .ZN(new_n968));
  XOR2_X1   g0768(.A(KEYINPUT114), .B(KEYINPUT44), .Z(new_n969));
  XNOR2_X1  g0769(.A(new_n968), .B(new_n969), .ZN(new_n970));
  NAND2_X1  g0770(.A1(new_n698), .A2(new_n967), .ZN(new_n971));
  XNOR2_X1  g0771(.A(new_n971), .B(KEYINPUT45), .ZN(new_n972));
  NOR2_X1   g0772(.A1(new_n970), .A2(new_n972), .ZN(new_n973));
  XNOR2_X1  g0773(.A(new_n973), .B(new_n696), .ZN(new_n974));
  NAND2_X1  g0774(.A1(new_n697), .A2(new_n538), .ZN(new_n975));
  OAI21_X1  g0775(.A(new_n975), .B1(new_n695), .B2(new_n697), .ZN(new_n976));
  XNOR2_X1  g0776(.A(new_n692), .B(new_n976), .ZN(new_n977));
  NAND2_X1  g0777(.A1(new_n977), .A2(new_n744), .ZN(new_n978));
  OAI21_X1  g0778(.A(new_n744), .B1(new_n974), .B2(new_n978), .ZN(new_n979));
  XOR2_X1   g0779(.A(new_n700), .B(KEYINPUT41), .Z(new_n980));
  NAND2_X1  g0780(.A1(new_n979), .A2(new_n980), .ZN(new_n981));
  NAND2_X1  g0781(.A1(new_n981), .A2(new_n748), .ZN(new_n982));
  NAND3_X1  g0782(.A1(new_n967), .A2(new_n538), .A3(new_n697), .ZN(new_n983));
  OR2_X1    g0783(.A1(new_n983), .A2(KEYINPUT42), .ZN(new_n984));
  OAI21_X1  g0784(.A(new_n608), .B1(new_n965), .B2(new_n694), .ZN(new_n985));
  AOI22_X1  g0785(.A1(new_n983), .A2(KEYINPUT42), .B1(new_n685), .B2(new_n985), .ZN(new_n986));
  AOI22_X1  g0786(.A1(new_n984), .A2(new_n986), .B1(KEYINPUT43), .B2(new_n962), .ZN(new_n987));
  NOR2_X1   g0787(.A1(new_n962), .A2(KEYINPUT43), .ZN(new_n988));
  XOR2_X1   g0788(.A(new_n987), .B(new_n988), .Z(new_n989));
  INV_X1    g0789(.A(new_n967), .ZN(new_n990));
  NOR2_X1   g0790(.A1(new_n696), .A2(new_n990), .ZN(new_n991));
  XNOR2_X1  g0791(.A(new_n989), .B(new_n991), .ZN(new_n992));
  AOI21_X1  g0792(.A(new_n964), .B1(new_n982), .B2(new_n992), .ZN(new_n993));
  INV_X1    g0793(.A(new_n993), .ZN(G387));
  AOI21_X1  g0794(.A(KEYINPUT119), .B1(new_n978), .B2(new_n746), .ZN(new_n995));
  INV_X1    g0795(.A(new_n995), .ZN(new_n996));
  NAND3_X1  g0796(.A1(new_n978), .A2(KEYINPUT119), .A3(new_n746), .ZN(new_n997));
  OAI211_X1 g0797(.A(new_n996), .B(new_n997), .C1(new_n744), .C2(new_n977), .ZN(new_n998));
  OR2_X1    g0798(.A1(new_n695), .A2(new_n815), .ZN(new_n999));
  OAI22_X1  g0799(.A1(new_n753), .A2(new_n701), .B1(G107), .B2(new_n212), .ZN(new_n1000));
  NAND2_X1  g0800(.A1(new_n240), .A2(G45), .ZN(new_n1001));
  INV_X1    g0801(.A(new_n701), .ZN(new_n1002));
  AOI211_X1 g0802(.A(G45), .B(new_n1002), .C1(G68), .C2(G77), .ZN(new_n1003));
  NOR2_X1   g0803(.A1(new_n353), .A2(G50), .ZN(new_n1004));
  XNOR2_X1  g0804(.A(KEYINPUT118), .B(KEYINPUT50), .ZN(new_n1005));
  XNOR2_X1  g0805(.A(new_n1004), .B(new_n1005), .ZN(new_n1006));
  AOI21_X1  g0806(.A(new_n757), .B1(new_n1003), .B2(new_n1006), .ZN(new_n1007));
  AOI21_X1  g0807(.A(new_n1000), .B1(new_n1001), .B2(new_n1007), .ZN(new_n1008));
  OAI21_X1  g0808(.A(new_n750), .B1(new_n1008), .B2(new_n765), .ZN(new_n1009));
  AOI21_X1  g0809(.A(new_n277), .B1(new_n938), .B2(G326), .ZN(new_n1010));
  AOI22_X1  g0810(.A1(G303), .A2(new_n794), .B1(new_n797), .B2(G311), .ZN(new_n1011));
  INV_X1    g0811(.A(G322), .ZN(new_n1012));
  INV_X1    g0812(.A(G317), .ZN(new_n1013));
  OAI221_X1 g0813(.A(new_n1011), .B1(new_n1012), .B2(new_n784), .C1(new_n776), .C2(new_n1013), .ZN(new_n1014));
  INV_X1    g0814(.A(KEYINPUT48), .ZN(new_n1015));
  OR2_X1    g0815(.A1(new_n1014), .A2(new_n1015), .ZN(new_n1016));
  NAND2_X1  g0816(.A1(new_n1014), .A2(new_n1015), .ZN(new_n1017));
  AOI22_X1  g0817(.A1(new_n831), .A2(G294), .B1(new_n790), .B2(G283), .ZN(new_n1018));
  NAND3_X1  g0818(.A1(new_n1016), .A2(new_n1017), .A3(new_n1018), .ZN(new_n1019));
  INV_X1    g0819(.A(KEYINPUT49), .ZN(new_n1020));
  OAI221_X1 g0820(.A(new_n1010), .B1(new_n511), .B2(new_n787), .C1(new_n1019), .C2(new_n1020), .ZN(new_n1021));
  AND2_X1   g0821(.A1(new_n1019), .A2(new_n1020), .ZN(new_n1022));
  NOR2_X1   g0822(.A1(new_n791), .A2(new_n390), .ZN(new_n1023));
  INV_X1    g0823(.A(new_n1023), .ZN(new_n1024));
  AOI22_X1  g0824(.A1(new_n831), .A2(G77), .B1(new_n938), .B2(G150), .ZN(new_n1025));
  NAND4_X1  g0825(.A1(new_n1024), .A2(new_n277), .A3(new_n940), .A4(new_n1025), .ZN(new_n1026));
  AOI22_X1  g0826(.A1(G68), .A2(new_n794), .B1(new_n797), .B2(new_n354), .ZN(new_n1027));
  OAI221_X1 g0827(.A(new_n1027), .B1(new_n860), .B2(new_n775), .C1(new_n423), .C2(new_n784), .ZN(new_n1028));
  OAI22_X1  g0828(.A1(new_n1021), .A2(new_n1022), .B1(new_n1026), .B2(new_n1028), .ZN(new_n1029));
  AOI21_X1  g0829(.A(new_n1009), .B1(new_n1029), .B2(new_n763), .ZN(new_n1030));
  AOI22_X1  g0830(.A1(new_n977), .A2(new_n749), .B1(new_n999), .B2(new_n1030), .ZN(new_n1031));
  NAND2_X1  g0831(.A1(new_n998), .A2(new_n1031), .ZN(G393));
  NAND2_X1  g0832(.A1(new_n990), .A2(new_n762), .ZN(new_n1033));
  XNOR2_X1  g0833(.A(new_n1033), .B(KEYINPUT120), .ZN(new_n1034));
  OAI21_X1  g0834(.A(new_n764), .B1(new_n204), .B2(new_n212), .ZN(new_n1035));
  NOR2_X1   g0835(.A1(new_n247), .A2(new_n757), .ZN(new_n1036));
  OAI21_X1  g0836(.A(new_n750), .B1(new_n1035), .B2(new_n1036), .ZN(new_n1037));
  OAI22_X1  g0837(.A1(new_n942), .A2(new_n775), .B1(new_n784), .B2(new_n1013), .ZN(new_n1038));
  XNOR2_X1  g0838(.A(new_n1038), .B(KEYINPUT52), .ZN(new_n1039));
  NOR2_X1   g0839(.A1(new_n791), .A2(new_n511), .ZN(new_n1040));
  OAI22_X1  g0840(.A1(new_n779), .A2(new_n845), .B1(new_n769), .B2(new_n1012), .ZN(new_n1041));
  NOR4_X1   g0841(.A1(new_n1040), .A2(new_n1041), .A3(new_n277), .A4(new_n788), .ZN(new_n1042));
  AOI22_X1  g0842(.A1(G294), .A2(new_n794), .B1(new_n797), .B2(G303), .ZN(new_n1043));
  NAND3_X1  g0843(.A1(new_n1039), .A2(new_n1042), .A3(new_n1043), .ZN(new_n1044));
  OAI22_X1  g0844(.A1(new_n835), .A2(new_n784), .B1(new_n775), .B2(new_n423), .ZN(new_n1045));
  XNOR2_X1  g0845(.A(new_n1045), .B(KEYINPUT51), .ZN(new_n1046));
  NOR2_X1   g0846(.A1(new_n791), .A2(new_n330), .ZN(new_n1047));
  OAI22_X1  g0847(.A1(new_n779), .A2(new_n322), .B1(new_n769), .B2(new_n836), .ZN(new_n1048));
  NOR4_X1   g0848(.A1(new_n1047), .A2(new_n1048), .A3(new_n285), .A4(new_n842), .ZN(new_n1049));
  AOI22_X1  g0849(.A1(G50), .A2(new_n797), .B1(new_n794), .B2(new_n354), .ZN(new_n1050));
  NAND3_X1  g0850(.A1(new_n1046), .A2(new_n1049), .A3(new_n1050), .ZN(new_n1051));
  NAND2_X1  g0851(.A1(new_n1044), .A2(new_n1051), .ZN(new_n1052));
  AOI21_X1  g0852(.A(new_n1037), .B1(new_n1052), .B2(new_n763), .ZN(new_n1053));
  NAND2_X1  g0853(.A1(new_n1034), .A2(new_n1053), .ZN(new_n1054));
  OAI21_X1  g0854(.A(new_n1054), .B1(new_n974), .B2(new_n748), .ZN(new_n1055));
  NOR2_X1   g0855(.A1(new_n974), .A2(new_n978), .ZN(new_n1056));
  NOR2_X1   g0856(.A1(new_n1056), .A2(new_n700), .ZN(new_n1057));
  NAND2_X1  g0857(.A1(new_n974), .A2(new_n978), .ZN(new_n1058));
  AOI21_X1  g0858(.A(new_n1055), .B1(new_n1057), .B2(new_n1058), .ZN(new_n1059));
  INV_X1    g0859(.A(new_n1059), .ZN(G390));
  OAI21_X1  g0860(.A(new_n824), .B1(new_n869), .B2(new_n867), .ZN(new_n1061));
  NAND2_X1  g0861(.A1(new_n917), .A2(G330), .ZN(new_n1062));
  NOR2_X1   g0862(.A1(new_n1061), .A2(new_n1062), .ZN(new_n1063));
  AOI22_X1  g0863(.A1(new_n901), .A2(new_n906), .B1(new_n870), .B2(new_n902), .ZN(new_n1064));
  NAND2_X1  g0864(.A1(new_n899), .A2(new_n902), .ZN(new_n1065));
  OAI211_X1 g0865(.A(new_n685), .B(new_n820), .C1(new_n739), .C2(new_n742), .ZN(new_n1066));
  AOI22_X1  g0866(.A1(new_n1066), .A2(new_n821), .B1(new_n920), .B2(new_n921), .ZN(new_n1067));
  NOR2_X1   g0867(.A1(new_n1065), .A2(new_n1067), .ZN(new_n1068));
  OAI21_X1  g0868(.A(new_n1063), .B1(new_n1064), .B2(new_n1068), .ZN(new_n1069));
  AND2_X1   g0869(.A1(new_n825), .A2(new_n821), .ZN(new_n1070));
  NOR2_X1   g0870(.A1(new_n869), .A2(new_n867), .ZN(new_n1071));
  OAI21_X1  g0871(.A(new_n902), .B1(new_n1070), .B2(new_n1071), .ZN(new_n1072));
  NAND2_X1  g0872(.A1(new_n890), .A2(new_n891), .ZN(new_n1073));
  NAND2_X1  g0873(.A1(new_n895), .A2(new_n879), .ZN(new_n1074));
  NAND2_X1  g0874(.A1(new_n1073), .A2(new_n1074), .ZN(new_n1075));
  NAND2_X1  g0875(.A1(new_n1075), .A2(new_n897), .ZN(new_n1076));
  AOI21_X1  g0876(.A(KEYINPUT39), .B1(new_n1076), .B2(new_n889), .ZN(new_n1077));
  NOR3_X1   g0877(.A1(new_n881), .A2(new_n884), .A3(new_n900), .ZN(new_n1078));
  OAI21_X1  g0878(.A(new_n1072), .B1(new_n1077), .B2(new_n1078), .ZN(new_n1079));
  AND2_X1   g0879(.A1(new_n1066), .A2(new_n821), .ZN(new_n1080));
  OAI211_X1 g0880(.A(new_n902), .B(new_n899), .C1(new_n1080), .C2(new_n1071), .ZN(new_n1081));
  NAND2_X1  g0881(.A1(new_n922), .A2(new_n726), .ZN(new_n1082));
  NAND3_X1  g0882(.A1(new_n1079), .A2(new_n1081), .A3(new_n1082), .ZN(new_n1083));
  NAND2_X1  g0883(.A1(new_n1069), .A2(new_n1083), .ZN(new_n1084));
  NAND3_X1  g0884(.A1(new_n725), .A2(G330), .A3(new_n824), .ZN(new_n1085));
  NAND3_X1  g0885(.A1(new_n1085), .A2(new_n920), .A3(new_n921), .ZN(new_n1086));
  OAI21_X1  g0886(.A(new_n1086), .B1(new_n1061), .B2(new_n1062), .ZN(new_n1087));
  NAND2_X1  g0887(.A1(new_n1087), .A2(new_n864), .ZN(new_n1088));
  OAI21_X1  g0888(.A(new_n1071), .B1(new_n1062), .B2(new_n822), .ZN(new_n1089));
  NAND3_X1  g0889(.A1(new_n1082), .A2(new_n1080), .A3(new_n1089), .ZN(new_n1090));
  NAND2_X1  g0890(.A1(new_n1088), .A2(new_n1090), .ZN(new_n1091));
  NAND3_X1  g0891(.A1(new_n483), .A2(G330), .A3(new_n917), .ZN(new_n1092));
  NAND3_X1  g0892(.A1(new_n1092), .A2(new_n909), .A3(new_n674), .ZN(new_n1093));
  INV_X1    g0893(.A(new_n1093), .ZN(new_n1094));
  NAND2_X1  g0894(.A1(new_n1091), .A2(new_n1094), .ZN(new_n1095));
  NAND2_X1  g0895(.A1(new_n1084), .A2(new_n1095), .ZN(new_n1096));
  AOI21_X1  g0896(.A(new_n1093), .B1(new_n1088), .B2(new_n1090), .ZN(new_n1097));
  NAND3_X1  g0897(.A1(new_n1097), .A2(new_n1069), .A3(new_n1083), .ZN(new_n1098));
  NAND3_X1  g0898(.A1(new_n1096), .A2(new_n746), .A3(new_n1098), .ZN(new_n1099));
  NAND3_X1  g0899(.A1(new_n1069), .A2(new_n1083), .A3(new_n749), .ZN(new_n1100));
  INV_X1    g0900(.A(new_n761), .ZN(new_n1101));
  OAI21_X1  g0901(.A(new_n1101), .B1(new_n1077), .B2(new_n1078), .ZN(new_n1102));
  AOI21_X1  g0902(.A(new_n849), .B1(new_n353), .B2(new_n850), .ZN(new_n1103));
  OAI22_X1  g0903(.A1(new_n204), .A2(new_n793), .B1(new_n775), .B2(new_n511), .ZN(new_n1104));
  NOR4_X1   g0904(.A1(new_n1047), .A2(new_n780), .A3(new_n830), .A4(new_n277), .ZN(new_n1105));
  OAI221_X1 g0905(.A(new_n1105), .B1(new_n845), .B2(new_n784), .C1(new_n496), .C2(new_n802), .ZN(new_n1106));
  AOI211_X1 g0906(.A(new_n1104), .B(new_n1106), .C1(G107), .C2(new_n797), .ZN(new_n1107));
  OR2_X1    g0907(.A1(new_n1107), .A2(KEYINPUT121), .ZN(new_n1108));
  OAI21_X1  g0908(.A(new_n277), .B1(new_n787), .B2(new_n860), .ZN(new_n1109));
  NAND2_X1  g0909(.A1(new_n831), .A2(G150), .ZN(new_n1110));
  XNOR2_X1  g0910(.A(new_n1110), .B(KEYINPUT53), .ZN(new_n1111));
  AOI211_X1 g0911(.A(new_n1109), .B(new_n1111), .C1(G159), .C2(new_n790), .ZN(new_n1112));
  NAND2_X1  g0912(.A1(new_n797), .A2(G137), .ZN(new_n1113));
  XOR2_X1   g0913(.A(KEYINPUT54), .B(G143), .Z(new_n1114));
  AOI22_X1  g0914(.A1(G132), .A2(new_n809), .B1(new_n794), .B2(new_n1114), .ZN(new_n1115));
  AOI22_X1  g0915(.A1(new_n803), .A2(G125), .B1(G128), .B2(new_n785), .ZN(new_n1116));
  NAND4_X1  g0916(.A1(new_n1112), .A2(new_n1113), .A3(new_n1115), .A4(new_n1116), .ZN(new_n1117));
  NAND2_X1  g0917(.A1(new_n1108), .A2(new_n1117), .ZN(new_n1118));
  AOI21_X1  g0918(.A(new_n1118), .B1(KEYINPUT121), .B2(new_n1107), .ZN(new_n1119));
  OAI211_X1 g0919(.A(new_n1102), .B(new_n1103), .C1(new_n956), .C2(new_n1119), .ZN(new_n1120));
  NAND3_X1  g0920(.A1(new_n1099), .A2(new_n1100), .A3(new_n1120), .ZN(G378));
  AOI21_X1  g0921(.A(new_n849), .B1(new_n860), .B2(new_n850), .ZN(new_n1122));
  XNOR2_X1  g0922(.A(new_n1122), .B(KEYINPUT122), .ZN(new_n1123));
  INV_X1    g0923(.A(new_n1123), .ZN(new_n1124));
  OAI22_X1  g0924(.A1(new_n204), .A2(new_n796), .B1(new_n775), .B2(new_n205), .ZN(new_n1125));
  NAND2_X1  g0925(.A1(new_n831), .A2(G77), .ZN(new_n1126));
  NAND2_X1  g0926(.A1(new_n804), .A2(G58), .ZN(new_n1127));
  NOR2_X1   g0927(.A1(new_n277), .A2(G41), .ZN(new_n1128));
  AND4_X1   g0928(.A1(new_n946), .A2(new_n1126), .A3(new_n1127), .A4(new_n1128), .ZN(new_n1129));
  OAI221_X1 g0929(.A(new_n1129), .B1(new_n511), .B2(new_n784), .C1(new_n845), .C2(new_n802), .ZN(new_n1130));
  AOI211_X1 g0930(.A(new_n1125), .B(new_n1130), .C1(new_n391), .C2(new_n794), .ZN(new_n1131));
  OR2_X1    g0931(.A1(new_n1131), .A2(KEYINPUT58), .ZN(new_n1132));
  AOI22_X1  g0932(.A1(new_n831), .A2(new_n1114), .B1(new_n790), .B2(G150), .ZN(new_n1133));
  INV_X1    g0933(.A(G132), .ZN(new_n1134));
  OAI21_X1  g0934(.A(new_n1133), .B1(new_n1134), .B2(new_n796), .ZN(new_n1135));
  INV_X1    g0935(.A(G125), .ZN(new_n1136));
  INV_X1    g0936(.A(G128), .ZN(new_n1137));
  OAI22_X1  g0937(.A1(new_n1136), .A2(new_n784), .B1(new_n775), .B2(new_n1137), .ZN(new_n1138));
  AOI211_X1 g0938(.A(new_n1135), .B(new_n1138), .C1(G137), .C2(new_n794), .ZN(new_n1139));
  INV_X1    g0939(.A(new_n1139), .ZN(new_n1140));
  OR2_X1    g0940(.A1(new_n1140), .A2(KEYINPUT59), .ZN(new_n1141));
  NAND2_X1  g0941(.A1(new_n1140), .A2(KEYINPUT59), .ZN(new_n1142));
  OAI211_X1 g0942(.A(new_n327), .B(new_n249), .C1(new_n787), .C2(new_n423), .ZN(new_n1143));
  AOI21_X1  g0943(.A(new_n1143), .B1(G124), .B2(new_n938), .ZN(new_n1144));
  NAND3_X1  g0944(.A1(new_n1141), .A2(new_n1142), .A3(new_n1144), .ZN(new_n1145));
  NAND2_X1  g0945(.A1(new_n1131), .A2(KEYINPUT58), .ZN(new_n1146));
  INV_X1    g0946(.A(new_n1128), .ZN(new_n1147));
  OAI211_X1 g0947(.A(new_n1147), .B(new_n860), .C1(G33), .C2(G41), .ZN(new_n1148));
  NAND4_X1  g0948(.A1(new_n1132), .A2(new_n1145), .A3(new_n1146), .A4(new_n1148), .ZN(new_n1149));
  AOI21_X1  g0949(.A(new_n1124), .B1(new_n1149), .B2(new_n763), .ZN(new_n1150));
  NAND3_X1  g0950(.A1(new_n380), .A2(new_n381), .A3(new_n387), .ZN(new_n1151));
  NOR2_X1   g0951(.A1(new_n360), .A2(new_n679), .ZN(new_n1152));
  XNOR2_X1  g0952(.A(new_n1151), .B(new_n1152), .ZN(new_n1153));
  XNOR2_X1  g0953(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1154));
  XNOR2_X1  g0954(.A(new_n1153), .B(new_n1154), .ZN(new_n1155));
  INV_X1    g0955(.A(new_n1155), .ZN(new_n1156));
  OAI21_X1  g0956(.A(new_n1150), .B1(new_n1156), .B2(new_n761), .ZN(new_n1157));
  INV_X1    g0957(.A(new_n1157), .ZN(new_n1158));
  INV_X1    g0958(.A(new_n913), .ZN(new_n1159));
  INV_X1    g0959(.A(new_n918), .ZN(new_n1160));
  NAND2_X1  g0960(.A1(new_n905), .A2(new_n889), .ZN(new_n1161));
  AOI21_X1  g0961(.A(new_n1159), .B1(new_n1160), .B2(new_n1161), .ZN(new_n1162));
  AOI21_X1  g0962(.A(new_n898), .B1(new_n1073), .B2(new_n1074), .ZN(new_n1163));
  OAI21_X1  g0963(.A(KEYINPUT40), .B1(new_n1163), .B2(new_n881), .ZN(new_n1164));
  OAI21_X1  g0964(.A(G330), .B1(new_n1164), .B2(new_n918), .ZN(new_n1165));
  OAI21_X1  g0965(.A(KEYINPUT123), .B1(new_n1162), .B2(new_n1165), .ZN(new_n1166));
  INV_X1    g0966(.A(KEYINPUT123), .ZN(new_n1167));
  NAND4_X1  g0967(.A1(new_n919), .A2(new_n923), .A3(new_n1167), .A4(G330), .ZN(new_n1168));
  NAND3_X1  g0968(.A1(new_n1166), .A2(new_n1168), .A3(new_n1156), .ZN(new_n1169));
  INV_X1    g0969(.A(new_n908), .ZN(new_n1170));
  NOR2_X1   g0970(.A1(new_n1162), .A2(new_n1165), .ZN(new_n1171));
  NAND3_X1  g0971(.A1(new_n1171), .A2(new_n1167), .A3(new_n1155), .ZN(new_n1172));
  AND3_X1   g0972(.A1(new_n1169), .A2(new_n1170), .A3(new_n1172), .ZN(new_n1173));
  AOI21_X1  g0973(.A(new_n1170), .B1(new_n1169), .B2(new_n1172), .ZN(new_n1174));
  NOR2_X1   g0974(.A1(new_n1173), .A2(new_n1174), .ZN(new_n1175));
  AOI21_X1  g0975(.A(new_n1158), .B1(new_n1175), .B2(new_n749), .ZN(new_n1176));
  NAND2_X1  g0976(.A1(new_n1098), .A2(new_n1094), .ZN(new_n1177));
  AOI21_X1  g0977(.A(KEYINPUT57), .B1(new_n1175), .B2(new_n1177), .ZN(new_n1178));
  NAND2_X1  g0978(.A1(new_n1169), .A2(new_n1172), .ZN(new_n1179));
  NAND2_X1  g0979(.A1(new_n1179), .A2(new_n908), .ZN(new_n1180));
  INV_X1    g0980(.A(KEYINPUT57), .ZN(new_n1181));
  AOI21_X1  g0981(.A(new_n1181), .B1(new_n1098), .B2(new_n1094), .ZN(new_n1182));
  NAND3_X1  g0982(.A1(new_n1169), .A2(new_n1172), .A3(new_n1170), .ZN(new_n1183));
  NAND3_X1  g0983(.A1(new_n1180), .A2(new_n1182), .A3(new_n1183), .ZN(new_n1184));
  NAND2_X1  g0984(.A1(new_n1184), .A2(new_n746), .ZN(new_n1185));
  OAI21_X1  g0985(.A(new_n1176), .B1(new_n1178), .B2(new_n1185), .ZN(G375));
  NAND2_X1  g0986(.A1(new_n1071), .A2(new_n760), .ZN(new_n1187));
  AOI22_X1  g0987(.A1(G107), .A2(new_n794), .B1(new_n797), .B2(G116), .ZN(new_n1188));
  OAI21_X1  g0988(.A(new_n1188), .B1(new_n496), .B2(new_n784), .ZN(new_n1189));
  OAI22_X1  g0989(.A1(new_n802), .A2(new_n541), .B1(new_n845), .B2(new_n775), .ZN(new_n1190));
  OAI221_X1 g0990(.A(new_n285), .B1(new_n787), .B2(new_n330), .C1(new_n204), .C2(new_n779), .ZN(new_n1191));
  NOR4_X1   g0991(.A1(new_n1189), .A2(new_n1023), .A3(new_n1190), .A4(new_n1191), .ZN(new_n1192));
  OAI211_X1 g0992(.A(new_n1127), .B(new_n277), .C1(new_n860), .C2(new_n791), .ZN(new_n1193));
  AOI21_X1  g0993(.A(new_n1193), .B1(new_n797), .B2(new_n1114), .ZN(new_n1194));
  OAI21_X1  g0994(.A(new_n1194), .B1(new_n835), .B2(new_n793), .ZN(new_n1195));
  NOR2_X1   g0995(.A1(new_n776), .A2(new_n947), .ZN(new_n1196));
  NOR2_X1   g0996(.A1(new_n784), .A2(new_n1134), .ZN(new_n1197));
  XNOR2_X1  g0997(.A(new_n1197), .B(KEYINPUT124), .ZN(new_n1198));
  NOR3_X1   g0998(.A1(new_n1195), .A2(new_n1196), .A3(new_n1198), .ZN(new_n1199));
  OAI22_X1  g0999(.A1(new_n802), .A2(new_n1137), .B1(new_n423), .B2(new_n779), .ZN(new_n1200));
  XNOR2_X1  g1000(.A(new_n1200), .B(KEYINPUT125), .ZN(new_n1201));
  INV_X1    g1001(.A(new_n1201), .ZN(new_n1202));
  AOI21_X1  g1002(.A(new_n1192), .B1(new_n1199), .B2(new_n1202), .ZN(new_n1203));
  NOR2_X1   g1003(.A1(new_n1203), .A2(new_n956), .ZN(new_n1204));
  AOI211_X1 g1004(.A(new_n849), .B(new_n1204), .C1(new_n322), .C2(new_n850), .ZN(new_n1205));
  AOI22_X1  g1005(.A1(new_n1091), .A2(new_n749), .B1(new_n1187), .B2(new_n1205), .ZN(new_n1206));
  NAND2_X1  g1006(.A1(new_n1095), .A2(new_n980), .ZN(new_n1207));
  NOR2_X1   g1007(.A1(new_n1091), .A2(new_n1094), .ZN(new_n1208));
  OAI21_X1  g1008(.A(new_n1206), .B1(new_n1207), .B2(new_n1208), .ZN(G381));
  NAND3_X1  g1009(.A1(new_n998), .A2(new_n817), .A3(new_n1031), .ZN(new_n1210));
  NOR2_X1   g1010(.A1(new_n1210), .A2(G381), .ZN(new_n1211));
  NAND4_X1  g1011(.A1(new_n993), .A2(new_n853), .A3(new_n1059), .A4(new_n1211), .ZN(new_n1212));
  OR3_X1    g1012(.A1(G375), .A2(new_n1212), .A3(G378), .ZN(G407));
  INV_X1    g1013(.A(G378), .ZN(new_n1214));
  NAND3_X1  g1014(.A1(new_n682), .A2(new_n683), .A3(G213), .ZN(new_n1215));
  INV_X1    g1015(.A(new_n1215), .ZN(new_n1216));
  NAND2_X1  g1016(.A1(new_n1214), .A2(new_n1216), .ZN(new_n1217));
  OAI211_X1 g1017(.A(G407), .B(G213), .C1(G375), .C2(new_n1217), .ZN(G409));
  NAND2_X1  g1018(.A1(G393), .A2(G396), .ZN(new_n1219));
  NAND2_X1  g1019(.A1(new_n1219), .A2(new_n1210), .ZN(new_n1220));
  NOR2_X1   g1020(.A1(new_n1220), .A2(new_n1059), .ZN(new_n1221));
  INV_X1    g1021(.A(new_n1221), .ZN(new_n1222));
  NAND2_X1  g1022(.A1(new_n1220), .A2(new_n1059), .ZN(new_n1223));
  AND3_X1   g1023(.A1(new_n1222), .A2(new_n993), .A3(new_n1223), .ZN(new_n1224));
  AOI21_X1  g1024(.A(new_n993), .B1(new_n1222), .B2(new_n1223), .ZN(new_n1225));
  NOR2_X1   g1025(.A1(new_n1224), .A2(new_n1225), .ZN(new_n1226));
  INV_X1    g1026(.A(KEYINPUT61), .ZN(new_n1227));
  OAI211_X1 g1027(.A(G378), .B(new_n1176), .C1(new_n1178), .C2(new_n1185), .ZN(new_n1228));
  NAND4_X1  g1028(.A1(new_n1180), .A2(new_n980), .A3(new_n1177), .A4(new_n1183), .ZN(new_n1229));
  NAND3_X1  g1029(.A1(new_n1180), .A2(new_n749), .A3(new_n1183), .ZN(new_n1230));
  NAND3_X1  g1030(.A1(new_n1229), .A2(new_n1230), .A3(new_n1157), .ZN(new_n1231));
  NAND2_X1  g1031(.A1(new_n1231), .A2(new_n1214), .ZN(new_n1232));
  AOI21_X1  g1032(.A(new_n1216), .B1(new_n1228), .B2(new_n1232), .ZN(new_n1233));
  NAND2_X1  g1033(.A1(new_n1095), .A2(KEYINPUT60), .ZN(new_n1234));
  INV_X1    g1034(.A(new_n1208), .ZN(new_n1235));
  NAND2_X1  g1035(.A1(new_n1234), .A2(new_n1235), .ZN(new_n1236));
  NAND3_X1  g1036(.A1(new_n1208), .A2(KEYINPUT60), .A3(new_n1095), .ZN(new_n1237));
  NAND3_X1  g1037(.A1(new_n1236), .A2(new_n746), .A3(new_n1237), .ZN(new_n1238));
  NAND3_X1  g1038(.A1(new_n1238), .A2(G384), .A3(new_n1206), .ZN(new_n1239));
  INV_X1    g1039(.A(new_n1239), .ZN(new_n1240));
  AOI21_X1  g1040(.A(G384), .B1(new_n1238), .B2(new_n1206), .ZN(new_n1241));
  OAI211_X1 g1041(.A(G2897), .B(new_n1216), .C1(new_n1240), .C2(new_n1241), .ZN(new_n1242));
  NAND2_X1  g1042(.A1(new_n1238), .A2(new_n1206), .ZN(new_n1243));
  NAND2_X1  g1043(.A1(new_n1243), .A2(new_n853), .ZN(new_n1244));
  NAND2_X1  g1044(.A1(new_n1216), .A2(G2897), .ZN(new_n1245));
  NAND3_X1  g1045(.A1(new_n1244), .A2(new_n1239), .A3(new_n1245), .ZN(new_n1246));
  NAND2_X1  g1046(.A1(new_n1242), .A2(new_n1246), .ZN(new_n1247));
  OAI21_X1  g1047(.A(new_n1227), .B1(new_n1233), .B2(new_n1247), .ZN(new_n1248));
  INV_X1    g1048(.A(KEYINPUT126), .ZN(new_n1249));
  NAND2_X1  g1049(.A1(new_n1249), .A2(KEYINPUT62), .ZN(new_n1250));
  NAND2_X1  g1050(.A1(new_n1244), .A2(new_n1239), .ZN(new_n1251));
  INV_X1    g1051(.A(new_n1251), .ZN(new_n1252));
  AOI21_X1  g1052(.A(new_n1250), .B1(new_n1233), .B2(new_n1252), .ZN(new_n1253));
  NOR2_X1   g1053(.A1(new_n1248), .A2(new_n1253), .ZN(new_n1254));
  NAND2_X1  g1054(.A1(new_n1233), .A2(new_n1252), .ZN(new_n1255));
  XOR2_X1   g1055(.A(KEYINPUT126), .B(KEYINPUT62), .Z(new_n1256));
  OR2_X1    g1056(.A1(new_n1255), .A2(new_n1256), .ZN(new_n1257));
  AOI21_X1  g1057(.A(new_n1226), .B1(new_n1254), .B2(new_n1257), .ZN(new_n1258));
  NAND3_X1  g1058(.A1(new_n1233), .A2(KEYINPUT63), .A3(new_n1252), .ZN(new_n1259));
  OAI211_X1 g1059(.A(new_n1259), .B(new_n1227), .C1(new_n1233), .C2(new_n1247), .ZN(new_n1260));
  AOI211_X1 g1060(.A(new_n1216), .B(new_n1251), .C1(new_n1228), .C2(new_n1232), .ZN(new_n1261));
  OAI21_X1  g1061(.A(new_n1226), .B1(new_n1261), .B2(KEYINPUT63), .ZN(new_n1262));
  NOR2_X1   g1062(.A1(new_n1260), .A2(new_n1262), .ZN(new_n1263));
  OAI21_X1  g1063(.A(KEYINPUT127), .B1(new_n1258), .B2(new_n1263), .ZN(new_n1264));
  INV_X1    g1064(.A(KEYINPUT127), .ZN(new_n1265));
  INV_X1    g1065(.A(new_n1248), .ZN(new_n1266));
  INV_X1    g1066(.A(KEYINPUT63), .ZN(new_n1267));
  NAND2_X1  g1067(.A1(new_n1255), .A2(new_n1267), .ZN(new_n1268));
  NAND4_X1  g1068(.A1(new_n1266), .A2(new_n1268), .A3(new_n1226), .A4(new_n1259), .ZN(new_n1269));
  NOR2_X1   g1069(.A1(new_n1255), .A2(new_n1256), .ZN(new_n1270));
  NOR3_X1   g1070(.A1(new_n1270), .A2(new_n1248), .A3(new_n1253), .ZN(new_n1271));
  OAI211_X1 g1071(.A(new_n1265), .B(new_n1269), .C1(new_n1271), .C2(new_n1226), .ZN(new_n1272));
  NAND2_X1  g1072(.A1(new_n1264), .A2(new_n1272), .ZN(G405));
  NAND2_X1  g1073(.A1(G375), .A2(new_n1214), .ZN(new_n1274));
  NAND2_X1  g1074(.A1(new_n1274), .A2(new_n1228), .ZN(new_n1275));
  XNOR2_X1  g1075(.A(new_n1275), .B(new_n1251), .ZN(new_n1276));
  XNOR2_X1  g1076(.A(new_n1276), .B(new_n1226), .ZN(G402));
endmodule


