//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 0 0 0 1 1 0 0 0 0 1 0 1 1 1 1 0 0 0 1 0 1 1 0 0 0 1 0 1 1 1 0 1 1 1 0 0 1 1 0 1 1 0 0 1 0 1 0 1 0 1 1 0 0 1 0 0 0 0 1 0 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:22:15 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n620, new_n621, new_n622,
    new_n623, new_n624, new_n625, new_n626, new_n628, new_n629, new_n630,
    new_n631, new_n632, new_n633, new_n634, new_n635, new_n636, new_n637,
    new_n638, new_n640, new_n641, new_n642, new_n643, new_n644, new_n645,
    new_n646, new_n647, new_n648, new_n649, new_n650, new_n651, new_n652,
    new_n653, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n689, new_n691, new_n692,
    new_n694, new_n695, new_n696, new_n697, new_n698, new_n699, new_n700,
    new_n702, new_n703, new_n704, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n718, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n850, new_n851, new_n852, new_n853, new_n854, new_n855, new_n857,
    new_n858, new_n859, new_n860, new_n861, new_n862, new_n863, new_n864,
    new_n865, new_n866, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n919, new_n920, new_n921, new_n922, new_n923, new_n924,
    new_n925, new_n926, new_n927, new_n928, new_n929, new_n930;
  INV_X1    g000(.A(KEYINPUT87), .ZN(new_n187));
  INV_X1    g001(.A(G143), .ZN(new_n188));
  NOR2_X1   g002(.A1(new_n188), .A2(G146), .ZN(new_n189));
  INV_X1    g003(.A(G146), .ZN(new_n190));
  OAI21_X1  g004(.A(KEYINPUT64), .B1(new_n190), .B2(G143), .ZN(new_n191));
  INV_X1    g005(.A(KEYINPUT64), .ZN(new_n192));
  NAND3_X1  g006(.A1(new_n192), .A2(new_n188), .A3(G146), .ZN(new_n193));
  AOI21_X1  g007(.A(new_n189), .B1(new_n191), .B2(new_n193), .ZN(new_n194));
  AND2_X1   g008(.A1(KEYINPUT0), .A2(G128), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n190), .A2(G143), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n188), .A2(G146), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n196), .A2(new_n197), .ZN(new_n198));
  NOR2_X1   g012(.A1(KEYINPUT0), .A2(G128), .ZN(new_n199));
  NOR2_X1   g013(.A1(new_n195), .A2(new_n199), .ZN(new_n200));
  AOI22_X1  g014(.A1(new_n194), .A2(new_n195), .B1(new_n198), .B2(new_n200), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n201), .A2(G125), .ZN(new_n202));
  OAI21_X1  g016(.A(KEYINPUT1), .B1(new_n188), .B2(G146), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n203), .A2(KEYINPUT66), .ZN(new_n204));
  INV_X1    g018(.A(KEYINPUT66), .ZN(new_n205));
  OAI211_X1 g019(.A(new_n205), .B(KEYINPUT1), .C1(new_n188), .C2(G146), .ZN(new_n206));
  NAND3_X1  g020(.A1(new_n204), .A2(G128), .A3(new_n206), .ZN(new_n207));
  INV_X1    g021(.A(G128), .ZN(new_n208));
  AOI21_X1  g022(.A(new_n208), .B1(new_n196), .B2(KEYINPUT1), .ZN(new_n209));
  AOI22_X1  g023(.A1(new_n207), .A2(new_n198), .B1(new_n194), .B2(new_n209), .ZN(new_n210));
  OAI21_X1  g024(.A(new_n202), .B1(new_n210), .B2(G125), .ZN(new_n211));
  XNOR2_X1  g025(.A(KEYINPUT81), .B(G224), .ZN(new_n212));
  NOR2_X1   g026(.A1(new_n212), .A2(G953), .ZN(new_n213));
  INV_X1    g027(.A(new_n213), .ZN(new_n214));
  AND2_X1   g028(.A1(new_n214), .A2(KEYINPUT7), .ZN(new_n215));
  NOR2_X1   g029(.A1(new_n211), .A2(new_n215), .ZN(new_n216));
  XNOR2_X1  g030(.A(KEYINPUT2), .B(G113), .ZN(new_n217));
  INV_X1    g031(.A(G116), .ZN(new_n218));
  OR2_X1    g032(.A1(KEYINPUT67), .A2(G119), .ZN(new_n219));
  NAND2_X1  g033(.A1(KEYINPUT67), .A2(G119), .ZN(new_n220));
  AOI21_X1  g034(.A(new_n218), .B1(new_n219), .B2(new_n220), .ZN(new_n221));
  INV_X1    g035(.A(G119), .ZN(new_n222));
  NOR2_X1   g036(.A1(new_n222), .A2(G116), .ZN(new_n223));
  OAI21_X1  g037(.A(new_n217), .B1(new_n221), .B2(new_n223), .ZN(new_n224));
  INV_X1    g038(.A(new_n217), .ZN(new_n225));
  AND2_X1   g039(.A1(KEYINPUT67), .A2(G119), .ZN(new_n226));
  NOR2_X1   g040(.A1(KEYINPUT67), .A2(G119), .ZN(new_n227));
  OAI21_X1  g041(.A(G116), .B1(new_n226), .B2(new_n227), .ZN(new_n228));
  INV_X1    g042(.A(new_n223), .ZN(new_n229));
  NAND3_X1  g043(.A1(new_n225), .A2(new_n228), .A3(new_n229), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n224), .A2(new_n230), .ZN(new_n231));
  INV_X1    g045(.A(G104), .ZN(new_n232));
  OAI21_X1  g046(.A(KEYINPUT3), .B1(new_n232), .B2(G107), .ZN(new_n233));
  INV_X1    g047(.A(KEYINPUT77), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n233), .A2(new_n234), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n232), .A2(G107), .ZN(new_n236));
  OR3_X1    g050(.A1(new_n232), .A2(KEYINPUT3), .A3(G107), .ZN(new_n237));
  OAI211_X1 g051(.A(KEYINPUT77), .B(KEYINPUT3), .C1(new_n232), .C2(G107), .ZN(new_n238));
  NAND4_X1  g052(.A1(new_n235), .A2(new_n236), .A3(new_n237), .A4(new_n238), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n239), .A2(G101), .ZN(new_n240));
  NOR3_X1   g054(.A1(new_n232), .A2(KEYINPUT3), .A3(G107), .ZN(new_n241));
  AOI21_X1  g055(.A(new_n241), .B1(new_n234), .B2(new_n233), .ZN(new_n242));
  INV_X1    g056(.A(G101), .ZN(new_n243));
  NAND4_X1  g057(.A1(new_n242), .A2(new_n243), .A3(new_n236), .A4(new_n238), .ZN(new_n244));
  NAND3_X1  g058(.A1(new_n240), .A2(new_n244), .A3(KEYINPUT4), .ZN(new_n245));
  INV_X1    g059(.A(KEYINPUT4), .ZN(new_n246));
  NAND3_X1  g060(.A1(new_n239), .A2(new_n246), .A3(G101), .ZN(new_n247));
  AND2_X1   g061(.A1(new_n245), .A2(new_n247), .ZN(new_n248));
  AOI21_X1  g062(.A(KEYINPUT78), .B1(new_n232), .B2(G107), .ZN(new_n249));
  NOR2_X1   g063(.A1(new_n232), .A2(G107), .ZN(new_n250));
  NOR2_X1   g064(.A1(new_n249), .A2(new_n250), .ZN(new_n251));
  NAND3_X1  g065(.A1(new_n232), .A2(KEYINPUT78), .A3(G107), .ZN(new_n252));
  AOI21_X1  g066(.A(new_n243), .B1(new_n251), .B2(new_n252), .ZN(new_n253));
  AND4_X1   g067(.A1(new_n236), .A2(new_n235), .A3(new_n238), .A4(new_n237), .ZN(new_n254));
  AOI21_X1  g068(.A(new_n253), .B1(new_n254), .B2(new_n243), .ZN(new_n255));
  INV_X1    g069(.A(KEYINPUT80), .ZN(new_n256));
  NAND3_X1  g070(.A1(new_n228), .A2(KEYINPUT5), .A3(new_n229), .ZN(new_n257));
  XNOR2_X1  g071(.A(KEYINPUT67), .B(G119), .ZN(new_n258));
  INV_X1    g072(.A(KEYINPUT5), .ZN(new_n259));
  NAND3_X1  g073(.A1(new_n258), .A2(new_n259), .A3(G116), .ZN(new_n260));
  NAND3_X1  g074(.A1(new_n257), .A2(G113), .A3(new_n260), .ZN(new_n261));
  NAND4_X1  g075(.A1(new_n255), .A2(new_n256), .A3(new_n230), .A4(new_n261), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n261), .A2(new_n230), .ZN(new_n263));
  INV_X1    g077(.A(KEYINPUT78), .ZN(new_n264));
  INV_X1    g078(.A(G107), .ZN(new_n265));
  OAI21_X1  g079(.A(new_n264), .B1(new_n265), .B2(G104), .ZN(new_n266));
  OAI211_X1 g080(.A(new_n266), .B(new_n252), .C1(new_n232), .C2(G107), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n267), .A2(G101), .ZN(new_n268));
  OAI21_X1  g082(.A(new_n268), .B1(new_n239), .B2(G101), .ZN(new_n269));
  OAI21_X1  g083(.A(KEYINPUT80), .B1(new_n263), .B2(new_n269), .ZN(new_n270));
  AOI22_X1  g084(.A1(new_n231), .A2(new_n248), .B1(new_n262), .B2(new_n270), .ZN(new_n271));
  XOR2_X1   g085(.A(G110), .B(G122), .Z(new_n272));
  INV_X1    g086(.A(new_n272), .ZN(new_n273));
  AOI21_X1  g087(.A(new_n216), .B1(new_n271), .B2(new_n273), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n211), .A2(new_n215), .ZN(new_n275));
  XNOR2_X1  g089(.A(new_n275), .B(KEYINPUT86), .ZN(new_n276));
  AND2_X1   g090(.A1(new_n261), .A2(new_n230), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n277), .A2(new_n255), .ZN(new_n278));
  INV_X1    g092(.A(KEYINPUT84), .ZN(new_n279));
  AND3_X1   g093(.A1(new_n263), .A2(new_n279), .A3(new_n269), .ZN(new_n280));
  AOI21_X1  g094(.A(new_n279), .B1(new_n263), .B2(new_n269), .ZN(new_n281));
  OAI21_X1  g095(.A(new_n278), .B1(new_n280), .B2(new_n281), .ZN(new_n282));
  XOR2_X1   g096(.A(KEYINPUT83), .B(KEYINPUT8), .Z(new_n283));
  XNOR2_X1  g097(.A(new_n272), .B(new_n283), .ZN(new_n284));
  INV_X1    g098(.A(new_n284), .ZN(new_n285));
  AND3_X1   g099(.A1(new_n282), .A2(KEYINPUT85), .A3(new_n285), .ZN(new_n286));
  AOI21_X1  g100(.A(KEYINPUT85), .B1(new_n282), .B2(new_n285), .ZN(new_n287));
  OAI211_X1 g101(.A(new_n274), .B(new_n276), .C1(new_n286), .C2(new_n287), .ZN(new_n288));
  INV_X1    g102(.A(G902), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n288), .A2(new_n289), .ZN(new_n290));
  NAND3_X1  g104(.A1(new_n245), .A2(new_n231), .A3(new_n247), .ZN(new_n291));
  AOI21_X1  g105(.A(new_n256), .B1(new_n277), .B2(new_n255), .ZN(new_n292));
  NOR3_X1   g106(.A1(new_n263), .A2(new_n269), .A3(KEYINPUT80), .ZN(new_n293));
  OAI21_X1  g107(.A(new_n291), .B1(new_n292), .B2(new_n293), .ZN(new_n294));
  NAND2_X1  g108(.A1(new_n294), .A2(new_n272), .ZN(new_n295));
  OAI211_X1 g109(.A(new_n273), .B(new_n291), .C1(new_n292), .C2(new_n293), .ZN(new_n296));
  NAND3_X1  g110(.A1(new_n295), .A2(KEYINPUT6), .A3(new_n296), .ZN(new_n297));
  INV_X1    g111(.A(KEYINPUT6), .ZN(new_n298));
  NAND3_X1  g112(.A1(new_n294), .A2(new_n298), .A3(new_n272), .ZN(new_n299));
  XNOR2_X1  g113(.A(new_n211), .B(new_n214), .ZN(new_n300));
  NAND3_X1  g114(.A1(new_n297), .A2(new_n299), .A3(new_n300), .ZN(new_n301));
  INV_X1    g115(.A(KEYINPUT82), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n301), .A2(new_n302), .ZN(new_n303));
  NAND4_X1  g117(.A1(new_n297), .A2(KEYINPUT82), .A3(new_n299), .A4(new_n300), .ZN(new_n304));
  AOI21_X1  g118(.A(new_n290), .B1(new_n303), .B2(new_n304), .ZN(new_n305));
  OAI21_X1  g119(.A(G210), .B1(G237), .B2(G902), .ZN(new_n306));
  AOI21_X1  g120(.A(new_n187), .B1(new_n305), .B2(new_n306), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n303), .A2(new_n304), .ZN(new_n308));
  INV_X1    g122(.A(new_n290), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n308), .A2(new_n309), .ZN(new_n310));
  INV_X1    g124(.A(new_n306), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n310), .A2(new_n311), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n307), .A2(new_n312), .ZN(new_n313));
  NAND3_X1  g127(.A1(new_n310), .A2(new_n187), .A3(new_n311), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n313), .A2(new_n314), .ZN(new_n315));
  OAI21_X1  g129(.A(G214), .B1(G237), .B2(G902), .ZN(new_n316));
  INV_X1    g130(.A(new_n316), .ZN(new_n317));
  OAI21_X1  g131(.A(KEYINPUT88), .B1(new_n315), .B2(new_n317), .ZN(new_n318));
  INV_X1    g132(.A(KEYINPUT88), .ZN(new_n319));
  NAND4_X1  g133(.A1(new_n313), .A2(new_n319), .A3(new_n316), .A4(new_n314), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n318), .A2(new_n320), .ZN(new_n321));
  INV_X1    g135(.A(G125), .ZN(new_n322));
  NOR3_X1   g136(.A1(new_n322), .A2(KEYINPUT16), .A3(G140), .ZN(new_n323));
  XNOR2_X1  g137(.A(G125), .B(G140), .ZN(new_n324));
  AOI21_X1  g138(.A(new_n323), .B1(new_n324), .B2(KEYINPUT16), .ZN(new_n325));
  XNOR2_X1  g139(.A(new_n325), .B(new_n190), .ZN(new_n326));
  INV_X1    g140(.A(new_n326), .ZN(new_n327));
  NOR2_X1   g141(.A1(new_n222), .A2(G128), .ZN(new_n328));
  AOI21_X1  g142(.A(new_n328), .B1(new_n258), .B2(G128), .ZN(new_n329));
  XOR2_X1   g143(.A(KEYINPUT24), .B(G110), .Z(new_n330));
  NAND2_X1  g144(.A1(new_n329), .A2(new_n330), .ZN(new_n331));
  INV_X1    g145(.A(KEYINPUT75), .ZN(new_n332));
  OAI21_X1  g146(.A(new_n332), .B1(new_n258), .B2(G128), .ZN(new_n333));
  OAI21_X1  g147(.A(G128), .B1(new_n226), .B2(new_n227), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n334), .A2(KEYINPUT23), .ZN(new_n335));
  NAND4_X1  g149(.A1(new_n219), .A2(KEYINPUT75), .A3(new_n208), .A4(new_n220), .ZN(new_n336));
  NAND3_X1  g150(.A1(new_n333), .A2(new_n335), .A3(new_n336), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n328), .A2(KEYINPUT23), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n337), .A2(new_n338), .ZN(new_n339));
  AOI21_X1  g153(.A(KEYINPUT76), .B1(new_n339), .B2(G110), .ZN(new_n340));
  INV_X1    g154(.A(KEYINPUT76), .ZN(new_n341));
  INV_X1    g155(.A(G110), .ZN(new_n342));
  AOI211_X1 g156(.A(new_n341), .B(new_n342), .C1(new_n337), .C2(new_n338), .ZN(new_n343));
  OAI211_X1 g157(.A(new_n327), .B(new_n331), .C1(new_n340), .C2(new_n343), .ZN(new_n344));
  OAI22_X1  g158(.A1(new_n339), .A2(G110), .B1(new_n329), .B2(new_n330), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n325), .A2(G146), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n324), .A2(new_n190), .ZN(new_n347));
  NAND3_X1  g161(.A1(new_n345), .A2(new_n346), .A3(new_n347), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n344), .A2(new_n348), .ZN(new_n349));
  XNOR2_X1  g163(.A(KEYINPUT22), .B(G137), .ZN(new_n350));
  INV_X1    g164(.A(G953), .ZN(new_n351));
  NAND3_X1  g165(.A1(new_n351), .A2(G221), .A3(G234), .ZN(new_n352));
  XNOR2_X1  g166(.A(new_n350), .B(new_n352), .ZN(new_n353));
  INV_X1    g167(.A(new_n353), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n349), .A2(new_n354), .ZN(new_n355));
  NAND3_X1  g169(.A1(new_n344), .A2(new_n348), .A3(new_n353), .ZN(new_n356));
  NAND3_X1  g170(.A1(new_n355), .A2(new_n289), .A3(new_n356), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n357), .A2(KEYINPUT25), .ZN(new_n358));
  INV_X1    g172(.A(G217), .ZN(new_n359));
  AOI21_X1  g173(.A(new_n359), .B1(G234), .B2(new_n289), .ZN(new_n360));
  INV_X1    g174(.A(KEYINPUT25), .ZN(new_n361));
  NAND4_X1  g175(.A1(new_n355), .A2(new_n361), .A3(new_n289), .A4(new_n356), .ZN(new_n362));
  NAND3_X1  g176(.A1(new_n358), .A2(new_n360), .A3(new_n362), .ZN(new_n363));
  OR2_X1    g177(.A1(new_n357), .A2(new_n360), .ZN(new_n364));
  NAND2_X1  g178(.A1(new_n363), .A2(new_n364), .ZN(new_n365));
  INV_X1    g179(.A(KEYINPUT31), .ZN(new_n366));
  INV_X1    g180(.A(new_n231), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n206), .A2(G128), .ZN(new_n368));
  AOI21_X1  g182(.A(new_n205), .B1(new_n196), .B2(KEYINPUT1), .ZN(new_n369));
  OAI21_X1  g183(.A(new_n198), .B1(new_n368), .B2(new_n369), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n194), .A2(new_n209), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n370), .A2(new_n371), .ZN(new_n372));
  INV_X1    g186(.A(G137), .ZN(new_n373));
  NAND3_X1  g187(.A1(new_n373), .A2(KEYINPUT65), .A3(G134), .ZN(new_n374));
  INV_X1    g188(.A(KEYINPUT65), .ZN(new_n375));
  OAI21_X1  g189(.A(new_n375), .B1(new_n373), .B2(G134), .ZN(new_n376));
  INV_X1    g190(.A(G134), .ZN(new_n377));
  NOR2_X1   g191(.A1(new_n377), .A2(G137), .ZN(new_n378));
  OAI211_X1 g192(.A(G131), .B(new_n374), .C1(new_n376), .C2(new_n378), .ZN(new_n379));
  INV_X1    g193(.A(KEYINPUT11), .ZN(new_n380));
  OAI21_X1  g194(.A(new_n380), .B1(new_n377), .B2(G137), .ZN(new_n381));
  NAND3_X1  g195(.A1(new_n373), .A2(KEYINPUT11), .A3(G134), .ZN(new_n382));
  INV_X1    g196(.A(G131), .ZN(new_n383));
  NAND2_X1  g197(.A1(new_n377), .A2(G137), .ZN(new_n384));
  NAND4_X1  g198(.A1(new_n381), .A2(new_n382), .A3(new_n383), .A4(new_n384), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n379), .A2(new_n385), .ZN(new_n386));
  INV_X1    g200(.A(new_n386), .ZN(new_n387));
  NAND3_X1  g201(.A1(new_n381), .A2(new_n384), .A3(new_n382), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n388), .A2(G131), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n389), .A2(new_n385), .ZN(new_n390));
  AOI22_X1  g204(.A1(new_n372), .A2(new_n387), .B1(new_n390), .B2(new_n201), .ZN(new_n391));
  INV_X1    g205(.A(KEYINPUT30), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n391), .A2(new_n392), .ZN(new_n393));
  AND2_X1   g207(.A1(new_n390), .A2(new_n201), .ZN(new_n394));
  AOI21_X1  g208(.A(new_n386), .B1(new_n371), .B2(new_n370), .ZN(new_n395));
  OAI21_X1  g209(.A(KEYINPUT30), .B1(new_n394), .B2(new_n395), .ZN(new_n396));
  AOI21_X1  g210(.A(new_n367), .B1(new_n393), .B2(new_n396), .ZN(new_n397));
  AND3_X1   g211(.A1(new_n224), .A2(new_n230), .A3(KEYINPUT68), .ZN(new_n398));
  AOI21_X1  g212(.A(KEYINPUT68), .B1(new_n224), .B2(new_n230), .ZN(new_n399));
  NOR2_X1   g213(.A1(new_n398), .A2(new_n399), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n400), .A2(new_n391), .ZN(new_n401));
  INV_X1    g215(.A(new_n401), .ZN(new_n402));
  NOR2_X1   g216(.A1(new_n397), .A2(new_n402), .ZN(new_n403));
  INV_X1    g217(.A(G237), .ZN(new_n404));
  NAND3_X1  g218(.A1(new_n404), .A2(new_n351), .A3(G210), .ZN(new_n405));
  XNOR2_X1  g219(.A(new_n405), .B(G101), .ZN(new_n406));
  XNOR2_X1  g220(.A(KEYINPUT26), .B(KEYINPUT27), .ZN(new_n407));
  XNOR2_X1  g221(.A(new_n406), .B(new_n407), .ZN(new_n408));
  AOI21_X1  g222(.A(new_n366), .B1(new_n403), .B2(new_n408), .ZN(new_n409));
  INV_X1    g223(.A(new_n408), .ZN(new_n410));
  NOR4_X1   g224(.A1(new_n397), .A2(new_n402), .A3(KEYINPUT31), .A4(new_n410), .ZN(new_n411));
  NOR2_X1   g225(.A1(new_n409), .A2(new_n411), .ZN(new_n412));
  AOI21_X1  g226(.A(KEYINPUT28), .B1(new_n400), .B2(new_n391), .ZN(new_n413));
  INV_X1    g227(.A(KEYINPUT70), .ZN(new_n414));
  NOR2_X1   g228(.A1(new_n413), .A2(new_n414), .ZN(new_n415));
  INV_X1    g229(.A(KEYINPUT69), .ZN(new_n416));
  OAI21_X1  g230(.A(new_n416), .B1(new_n391), .B2(new_n367), .ZN(new_n417));
  OAI211_X1 g231(.A(KEYINPUT69), .B(new_n231), .C1(new_n394), .C2(new_n395), .ZN(new_n418));
  NAND3_X1  g232(.A1(new_n417), .A2(new_n401), .A3(new_n418), .ZN(new_n419));
  AOI21_X1  g233(.A(new_n415), .B1(KEYINPUT28), .B2(new_n419), .ZN(new_n420));
  NAND3_X1  g234(.A1(new_n419), .A2(KEYINPUT70), .A3(KEYINPUT28), .ZN(new_n421));
  INV_X1    g235(.A(new_n421), .ZN(new_n422));
  OAI21_X1  g236(.A(new_n410), .B1(new_n420), .B2(new_n422), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n412), .A2(new_n423), .ZN(new_n424));
  NOR2_X1   g238(.A1(G472), .A2(G902), .ZN(new_n425));
  AND3_X1   g239(.A1(new_n424), .A2(KEYINPUT32), .A3(new_n425), .ZN(new_n426));
  INV_X1    g240(.A(KEYINPUT28), .ZN(new_n427));
  OAI21_X1  g241(.A(new_n231), .B1(new_n394), .B2(new_n395), .ZN(new_n428));
  AOI22_X1  g242(.A1(new_n428), .A2(new_n416), .B1(new_n391), .B2(new_n400), .ZN(new_n429));
  AOI21_X1  g243(.A(new_n427), .B1(new_n429), .B2(new_n418), .ZN(new_n430));
  OAI211_X1 g244(.A(new_n408), .B(new_n421), .C1(new_n430), .C2(new_n415), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n431), .A2(KEYINPUT72), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n419), .A2(KEYINPUT28), .ZN(new_n433));
  OAI21_X1  g247(.A(new_n433), .B1(new_n414), .B2(new_n413), .ZN(new_n434));
  INV_X1    g248(.A(KEYINPUT72), .ZN(new_n435));
  NAND4_X1  g249(.A1(new_n434), .A2(new_n435), .A3(new_n408), .A4(new_n421), .ZN(new_n436));
  INV_X1    g250(.A(new_n403), .ZN(new_n437));
  AOI21_X1  g251(.A(KEYINPUT29), .B1(new_n437), .B2(new_n410), .ZN(new_n438));
  NAND3_X1  g252(.A1(new_n432), .A2(new_n436), .A3(new_n438), .ZN(new_n439));
  INV_X1    g253(.A(KEYINPUT74), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n408), .A2(KEYINPUT29), .ZN(new_n441));
  INV_X1    g255(.A(KEYINPUT73), .ZN(new_n442));
  OAI221_X1 g256(.A(new_n442), .B1(new_n398), .B2(new_n399), .C1(new_n394), .C2(new_n395), .ZN(new_n443));
  OAI21_X1  g257(.A(KEYINPUT73), .B1(new_n400), .B2(new_n391), .ZN(new_n444));
  NAND3_X1  g258(.A1(new_n443), .A2(new_n444), .A3(new_n401), .ZN(new_n445));
  AOI211_X1 g259(.A(new_n413), .B(new_n441), .C1(new_n445), .C2(KEYINPUT28), .ZN(new_n446));
  OAI21_X1  g260(.A(new_n440), .B1(new_n446), .B2(G902), .ZN(new_n447));
  AOI21_X1  g261(.A(new_n413), .B1(new_n445), .B2(KEYINPUT28), .ZN(new_n448));
  INV_X1    g262(.A(new_n441), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n448), .A2(new_n449), .ZN(new_n450));
  NAND3_X1  g264(.A1(new_n450), .A2(KEYINPUT74), .A3(new_n289), .ZN(new_n451));
  NAND3_X1  g265(.A1(new_n439), .A2(new_n447), .A3(new_n451), .ZN(new_n452));
  AOI21_X1  g266(.A(new_n426), .B1(new_n452), .B2(G472), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n424), .A2(new_n425), .ZN(new_n454));
  NOR2_X1   g268(.A1(KEYINPUT71), .A2(KEYINPUT32), .ZN(new_n455));
  AND2_X1   g269(.A1(KEYINPUT71), .A2(KEYINPUT32), .ZN(new_n456));
  OAI21_X1  g270(.A(new_n454), .B1(new_n455), .B2(new_n456), .ZN(new_n457));
  AOI21_X1  g271(.A(new_n365), .B1(new_n453), .B2(new_n457), .ZN(new_n458));
  INV_X1    g272(.A(G475), .ZN(new_n459));
  NAND3_X1  g273(.A1(new_n404), .A2(new_n351), .A3(G214), .ZN(new_n460));
  NAND2_X1  g274(.A1(new_n460), .A2(new_n188), .ZN(new_n461));
  NAND4_X1  g275(.A1(new_n404), .A2(new_n351), .A3(G143), .A4(G214), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n463), .A2(G131), .ZN(new_n464));
  INV_X1    g278(.A(KEYINPUT90), .ZN(new_n465));
  NAND2_X1  g279(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  NAND3_X1  g280(.A1(new_n463), .A2(KEYINPUT90), .A3(G131), .ZN(new_n467));
  NAND3_X1  g281(.A1(new_n466), .A2(KEYINPUT17), .A3(new_n467), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n468), .A2(new_n326), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n469), .A2(KEYINPUT91), .ZN(new_n470));
  NAND2_X1  g284(.A1(new_n466), .A2(new_n467), .ZN(new_n471));
  INV_X1    g285(.A(KEYINPUT17), .ZN(new_n472));
  INV_X1    g286(.A(new_n463), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n473), .A2(new_n383), .ZN(new_n474));
  NAND3_X1  g288(.A1(new_n471), .A2(new_n472), .A3(new_n474), .ZN(new_n475));
  INV_X1    g289(.A(KEYINPUT91), .ZN(new_n476));
  NAND3_X1  g290(.A1(new_n468), .A2(new_n476), .A3(new_n326), .ZN(new_n477));
  NAND3_X1  g291(.A1(new_n470), .A2(new_n475), .A3(new_n477), .ZN(new_n478));
  NAND2_X1  g292(.A1(KEYINPUT18), .A2(G131), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n473), .A2(new_n479), .ZN(new_n480));
  INV_X1    g294(.A(KEYINPUT89), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n480), .A2(new_n481), .ZN(new_n482));
  NAND3_X1  g296(.A1(new_n473), .A2(KEYINPUT89), .A3(new_n479), .ZN(new_n483));
  OR2_X1    g297(.A1(new_n324), .A2(new_n190), .ZN(new_n484));
  AOI22_X1  g298(.A1(new_n482), .A2(new_n483), .B1(new_n347), .B2(new_n484), .ZN(new_n485));
  NAND3_X1  g299(.A1(new_n463), .A2(KEYINPUT18), .A3(G131), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n485), .A2(new_n486), .ZN(new_n487));
  NAND2_X1  g301(.A1(new_n478), .A2(new_n487), .ZN(new_n488));
  XNOR2_X1  g302(.A(G113), .B(G122), .ZN(new_n489));
  XNOR2_X1  g303(.A(new_n489), .B(new_n232), .ZN(new_n490));
  INV_X1    g304(.A(new_n490), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n488), .A2(new_n491), .ZN(new_n492));
  NAND3_X1  g306(.A1(new_n478), .A2(new_n490), .A3(new_n487), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  AOI21_X1  g308(.A(new_n459), .B1(new_n494), .B2(new_n289), .ZN(new_n495));
  INV_X1    g309(.A(new_n487), .ZN(new_n496));
  XOR2_X1   g310(.A(new_n324), .B(KEYINPUT19), .Z(new_n497));
  OAI21_X1  g311(.A(new_n346), .B1(new_n497), .B2(G146), .ZN(new_n498));
  AOI21_X1  g312(.A(new_n498), .B1(new_n471), .B2(new_n474), .ZN(new_n499));
  OAI21_X1  g313(.A(new_n491), .B1(new_n496), .B2(new_n499), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n493), .A2(new_n500), .ZN(new_n501));
  NAND3_X1  g315(.A1(new_n501), .A2(new_n459), .A3(new_n289), .ZN(new_n502));
  INV_X1    g316(.A(KEYINPUT92), .ZN(new_n503));
  AOI21_X1  g317(.A(new_n503), .B1(new_n493), .B2(new_n500), .ZN(new_n504));
  OAI21_X1  g318(.A(new_n502), .B1(KEYINPUT20), .B2(new_n504), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n501), .A2(KEYINPUT92), .ZN(new_n506));
  INV_X1    g320(.A(KEYINPUT20), .ZN(new_n507));
  AOI21_X1  g321(.A(G475), .B1(new_n493), .B2(new_n500), .ZN(new_n508));
  NAND4_X1  g322(.A1(new_n506), .A2(new_n507), .A3(new_n289), .A4(new_n508), .ZN(new_n509));
  AOI21_X1  g323(.A(new_n495), .B1(new_n505), .B2(new_n509), .ZN(new_n510));
  INV_X1    g324(.A(new_n510), .ZN(new_n511));
  XNOR2_X1  g325(.A(G128), .B(G143), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n512), .A2(KEYINPUT13), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n188), .A2(G128), .ZN(new_n514));
  OAI211_X1 g328(.A(new_n513), .B(G134), .C1(KEYINPUT13), .C2(new_n514), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n512), .A2(new_n377), .ZN(new_n516));
  INV_X1    g330(.A(G122), .ZN(new_n517));
  AND2_X1   g331(.A1(new_n517), .A2(KEYINPUT93), .ZN(new_n518));
  NOR2_X1   g332(.A1(new_n517), .A2(KEYINPUT93), .ZN(new_n519));
  OAI21_X1  g333(.A(G116), .B1(new_n518), .B2(new_n519), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n218), .A2(G122), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n522), .A2(KEYINPUT94), .ZN(new_n523));
  INV_X1    g337(.A(KEYINPUT94), .ZN(new_n524));
  NAND3_X1  g338(.A1(new_n520), .A2(new_n524), .A3(new_n521), .ZN(new_n525));
  NAND3_X1  g339(.A1(new_n523), .A2(new_n265), .A3(new_n525), .ZN(new_n526));
  INV_X1    g340(.A(new_n526), .ZN(new_n527));
  AOI21_X1  g341(.A(new_n265), .B1(new_n523), .B2(new_n525), .ZN(new_n528));
  OAI211_X1 g342(.A(new_n515), .B(new_n516), .C1(new_n527), .C2(new_n528), .ZN(new_n529));
  XNOR2_X1  g343(.A(new_n512), .B(new_n377), .ZN(new_n530));
  XNOR2_X1  g344(.A(new_n530), .B(KEYINPUT95), .ZN(new_n531));
  INV_X1    g345(.A(new_n520), .ZN(new_n532));
  XNOR2_X1  g346(.A(new_n521), .B(KEYINPUT14), .ZN(new_n533));
  OAI21_X1  g347(.A(G107), .B1(new_n532), .B2(new_n533), .ZN(new_n534));
  NAND3_X1  g348(.A1(new_n531), .A2(new_n526), .A3(new_n534), .ZN(new_n535));
  XOR2_X1   g349(.A(KEYINPUT9), .B(G234), .Z(new_n536));
  INV_X1    g350(.A(new_n536), .ZN(new_n537));
  NOR3_X1   g351(.A1(new_n537), .A2(new_n359), .A3(G953), .ZN(new_n538));
  NAND3_X1  g352(.A1(new_n529), .A2(new_n535), .A3(new_n538), .ZN(new_n539));
  INV_X1    g353(.A(new_n539), .ZN(new_n540));
  AOI21_X1  g354(.A(new_n538), .B1(new_n529), .B2(new_n535), .ZN(new_n541));
  OAI21_X1  g355(.A(new_n289), .B1(new_n540), .B2(new_n541), .ZN(new_n542));
  XNOR2_X1  g356(.A(new_n542), .B(KEYINPUT96), .ZN(new_n543));
  INV_X1    g357(.A(KEYINPUT15), .ZN(new_n544));
  NAND2_X1  g358(.A1(new_n544), .A2(G478), .ZN(new_n545));
  NAND2_X1  g359(.A1(new_n543), .A2(new_n545), .ZN(new_n546));
  OAI211_X1 g360(.A(new_n544), .B(G478), .C1(new_n542), .C2(KEYINPUT96), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n546), .A2(new_n547), .ZN(new_n548));
  NAND2_X1  g362(.A1(G234), .A2(G237), .ZN(new_n549));
  NAND3_X1  g363(.A1(new_n549), .A2(G952), .A3(new_n351), .ZN(new_n550));
  INV_X1    g364(.A(new_n550), .ZN(new_n551));
  XOR2_X1   g365(.A(KEYINPUT21), .B(G898), .Z(new_n552));
  INV_X1    g366(.A(new_n552), .ZN(new_n553));
  NAND3_X1  g367(.A1(new_n549), .A2(G902), .A3(G953), .ZN(new_n554));
  INV_X1    g368(.A(new_n554), .ZN(new_n555));
  AOI21_X1  g369(.A(new_n551), .B1(new_n553), .B2(new_n555), .ZN(new_n556));
  NOR3_X1   g370(.A1(new_n511), .A2(new_n548), .A3(new_n556), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n269), .A2(new_n210), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n203), .A2(G128), .ZN(new_n559));
  XNOR2_X1  g373(.A(new_n194), .B(new_n559), .ZN(new_n560));
  OAI21_X1  g374(.A(new_n558), .B1(new_n269), .B2(new_n560), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n561), .A2(new_n390), .ZN(new_n562));
  INV_X1    g376(.A(KEYINPUT12), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  NAND3_X1  g378(.A1(new_n561), .A2(KEYINPUT12), .A3(new_n390), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  XOR2_X1   g380(.A(G110), .B(G140), .Z(new_n567));
  AND2_X1   g381(.A1(new_n351), .A2(G227), .ZN(new_n568));
  XNOR2_X1  g382(.A(new_n567), .B(new_n568), .ZN(new_n569));
  NAND3_X1  g383(.A1(new_n245), .A2(new_n201), .A3(new_n247), .ZN(new_n570));
  INV_X1    g384(.A(new_n390), .ZN(new_n571));
  INV_X1    g385(.A(KEYINPUT10), .ZN(new_n572));
  OAI21_X1  g386(.A(new_n572), .B1(new_n560), .B2(new_n269), .ZN(new_n573));
  NAND4_X1  g387(.A1(new_n372), .A2(KEYINPUT10), .A3(new_n244), .A4(new_n268), .ZN(new_n574));
  NAND4_X1  g388(.A1(new_n570), .A2(new_n571), .A3(new_n573), .A4(new_n574), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n575), .A2(KEYINPUT79), .ZN(new_n576));
  INV_X1    g390(.A(new_n576), .ZN(new_n577));
  NOR2_X1   g391(.A1(new_n575), .A2(KEYINPUT79), .ZN(new_n578));
  OAI211_X1 g392(.A(new_n566), .B(new_n569), .C1(new_n577), .C2(new_n578), .ZN(new_n579));
  OR2_X1    g393(.A1(new_n575), .A2(KEYINPUT79), .ZN(new_n580));
  NAND3_X1  g394(.A1(new_n570), .A2(new_n573), .A3(new_n574), .ZN(new_n581));
  AOI22_X1  g395(.A1(new_n580), .A2(new_n576), .B1(new_n390), .B2(new_n581), .ZN(new_n582));
  OAI21_X1  g396(.A(new_n579), .B1(new_n582), .B2(new_n569), .ZN(new_n583));
  INV_X1    g397(.A(G469), .ZN(new_n584));
  NAND3_X1  g398(.A1(new_n583), .A2(new_n584), .A3(new_n289), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n581), .A2(new_n390), .ZN(new_n586));
  OAI211_X1 g400(.A(new_n586), .B(new_n569), .C1(new_n577), .C2(new_n578), .ZN(new_n587));
  AOI22_X1  g401(.A1(new_n580), .A2(new_n576), .B1(new_n565), .B2(new_n564), .ZN(new_n588));
  OAI211_X1 g402(.A(new_n587), .B(G469), .C1(new_n588), .C2(new_n569), .ZN(new_n589));
  NAND2_X1  g403(.A1(G469), .A2(G902), .ZN(new_n590));
  NAND3_X1  g404(.A1(new_n585), .A2(new_n589), .A3(new_n590), .ZN(new_n591));
  OAI21_X1  g405(.A(G221), .B1(new_n537), .B2(G902), .ZN(new_n592));
  AND2_X1   g406(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  AND2_X1   g407(.A1(new_n557), .A2(new_n593), .ZN(new_n594));
  NAND3_X1  g408(.A1(new_n321), .A2(new_n458), .A3(new_n594), .ZN(new_n595));
  XNOR2_X1  g409(.A(new_n595), .B(G101), .ZN(G3));
  INV_X1    g410(.A(KEYINPUT97), .ZN(new_n597));
  AOI21_X1  g411(.A(new_n597), .B1(new_n305), .B2(new_n306), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n598), .A2(new_n312), .ZN(new_n599));
  AOI21_X1  g413(.A(new_n306), .B1(new_n308), .B2(new_n309), .ZN(new_n600));
  AOI21_X1  g414(.A(new_n317), .B1(new_n600), .B2(new_n597), .ZN(new_n601));
  AND3_X1   g415(.A1(new_n599), .A2(new_n593), .A3(new_n601), .ZN(new_n602));
  OAI21_X1  g416(.A(KEYINPUT33), .B1(new_n540), .B2(new_n541), .ZN(new_n603));
  INV_X1    g417(.A(new_n541), .ZN(new_n604));
  INV_X1    g418(.A(KEYINPUT33), .ZN(new_n605));
  NAND3_X1  g419(.A1(new_n604), .A2(new_n605), .A3(new_n539), .ZN(new_n606));
  AOI21_X1  g420(.A(G902), .B1(new_n603), .B2(new_n606), .ZN(new_n607));
  XOR2_X1   g421(.A(KEYINPUT98), .B(G478), .Z(new_n608));
  AOI22_X1  g422(.A1(new_n607), .A2(G478), .B1(new_n542), .B2(new_n608), .ZN(new_n609));
  INV_X1    g423(.A(new_n609), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n511), .A2(new_n610), .ZN(new_n611));
  NOR2_X1   g425(.A1(new_n611), .A2(new_n556), .ZN(new_n612));
  AND2_X1   g426(.A1(new_n412), .A2(new_n423), .ZN(new_n613));
  OAI21_X1  g427(.A(G472), .B1(new_n613), .B2(G902), .ZN(new_n614));
  NAND2_X1  g428(.A1(new_n614), .A2(new_n454), .ZN(new_n615));
  NOR2_X1   g429(.A1(new_n615), .A2(new_n365), .ZN(new_n616));
  NAND3_X1  g430(.A1(new_n602), .A2(new_n612), .A3(new_n616), .ZN(new_n617));
  XOR2_X1   g431(.A(KEYINPUT34), .B(G104), .Z(new_n618));
  XNOR2_X1  g432(.A(new_n617), .B(new_n618), .ZN(G6));
  XNOR2_X1  g433(.A(new_n502), .B(new_n507), .ZN(new_n620));
  OR2_X1    g434(.A1(new_n620), .A2(new_n495), .ZN(new_n621));
  INV_X1    g435(.A(new_n547), .ZN(new_n622));
  AOI21_X1  g436(.A(new_n622), .B1(new_n543), .B2(new_n545), .ZN(new_n623));
  NOR3_X1   g437(.A1(new_n621), .A2(new_n623), .A3(new_n556), .ZN(new_n624));
  NAND3_X1  g438(.A1(new_n602), .A2(new_n616), .A3(new_n624), .ZN(new_n625));
  XOR2_X1   g439(.A(KEYINPUT35), .B(G107), .Z(new_n626));
  XNOR2_X1  g440(.A(new_n625), .B(new_n626), .ZN(G9));
  NOR2_X1   g441(.A1(new_n354), .A2(KEYINPUT36), .ZN(new_n628));
  XNOR2_X1  g442(.A(new_n349), .B(new_n628), .ZN(new_n629));
  OAI211_X1 g443(.A(new_n629), .B(new_n289), .C1(new_n359), .C2(G234), .ZN(new_n630));
  AOI21_X1  g444(.A(KEYINPUT99), .B1(new_n363), .B2(new_n630), .ZN(new_n631));
  INV_X1    g445(.A(new_n631), .ZN(new_n632));
  NAND3_X1  g446(.A1(new_n363), .A2(KEYINPUT99), .A3(new_n630), .ZN(new_n633));
  NAND2_X1  g447(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  NOR2_X1   g448(.A1(new_n634), .A2(new_n615), .ZN(new_n635));
  NAND3_X1  g449(.A1(new_n321), .A2(new_n594), .A3(new_n635), .ZN(new_n636));
  XNOR2_X1  g450(.A(KEYINPUT37), .B(G110), .ZN(new_n637));
  XNOR2_X1  g451(.A(new_n637), .B(KEYINPUT100), .ZN(new_n638));
  XNOR2_X1  g452(.A(new_n636), .B(new_n638), .ZN(G12));
  NAND3_X1  g453(.A1(new_n599), .A2(new_n593), .A3(new_n601), .ZN(new_n640));
  AND3_X1   g454(.A1(new_n432), .A2(new_n438), .A3(new_n436), .ZN(new_n641));
  NAND2_X1  g455(.A1(new_n447), .A2(new_n451), .ZN(new_n642));
  OAI21_X1  g456(.A(G472), .B1(new_n641), .B2(new_n642), .ZN(new_n643));
  NAND3_X1  g457(.A1(new_n424), .A2(KEYINPUT32), .A3(new_n425), .ZN(new_n644));
  NAND3_X1  g458(.A1(new_n643), .A2(new_n457), .A3(new_n644), .ZN(new_n645));
  INV_X1    g459(.A(new_n633), .ZN(new_n646));
  NOR2_X1   g460(.A1(new_n646), .A2(new_n631), .ZN(new_n647));
  NAND2_X1  g461(.A1(new_n645), .A2(new_n647), .ZN(new_n648));
  NOR2_X1   g462(.A1(new_n640), .A2(new_n648), .ZN(new_n649));
  INV_X1    g463(.A(G900), .ZN(new_n650));
  AOI21_X1  g464(.A(new_n551), .B1(new_n555), .B2(new_n650), .ZN(new_n651));
  NOR3_X1   g465(.A1(new_n621), .A2(new_n623), .A3(new_n651), .ZN(new_n652));
  NAND2_X1  g466(.A1(new_n649), .A2(new_n652), .ZN(new_n653));
  XNOR2_X1  g467(.A(new_n653), .B(G128), .ZN(G30));
  XOR2_X1   g468(.A(new_n651), .B(KEYINPUT39), .Z(new_n655));
  NAND2_X1  g469(.A1(new_n593), .A2(new_n655), .ZN(new_n656));
  XOR2_X1   g470(.A(new_n656), .B(KEYINPUT101), .Z(new_n657));
  XOR2_X1   g471(.A(new_n657), .B(KEYINPUT40), .Z(new_n658));
  XNOR2_X1  g472(.A(new_n315), .B(KEYINPUT38), .ZN(new_n659));
  NAND2_X1  g473(.A1(new_n403), .A2(new_n408), .ZN(new_n660));
  NAND2_X1  g474(.A1(new_n445), .A2(new_n410), .ZN(new_n661));
  AND2_X1   g475(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  OAI21_X1  g476(.A(G472), .B1(new_n662), .B2(G902), .ZN(new_n663));
  NAND3_X1  g477(.A1(new_n457), .A2(new_n644), .A3(new_n663), .ZN(new_n664));
  INV_X1    g478(.A(new_n664), .ZN(new_n665));
  NOR4_X1   g479(.A1(new_n659), .A2(new_n510), .A3(new_n623), .A4(new_n665), .ZN(new_n666));
  NAND4_X1  g480(.A1(new_n658), .A2(new_n316), .A3(new_n634), .A4(new_n666), .ZN(new_n667));
  XNOR2_X1  g481(.A(KEYINPUT102), .B(G143), .ZN(new_n668));
  XNOR2_X1  g482(.A(new_n667), .B(new_n668), .ZN(G45));
  AOI21_X1  g483(.A(new_n634), .B1(new_n453), .B2(new_n457), .ZN(new_n670));
  NOR3_X1   g484(.A1(new_n510), .A2(new_n609), .A3(new_n651), .ZN(new_n671));
  NAND3_X1  g485(.A1(new_n602), .A2(new_n670), .A3(new_n671), .ZN(new_n672));
  NAND2_X1  g486(.A1(new_n672), .A2(KEYINPUT103), .ZN(new_n673));
  INV_X1    g487(.A(KEYINPUT103), .ZN(new_n674));
  NAND3_X1  g488(.A1(new_n649), .A2(new_n674), .A3(new_n671), .ZN(new_n675));
  NAND2_X1  g489(.A1(new_n673), .A2(new_n675), .ZN(new_n676));
  XNOR2_X1  g490(.A(new_n676), .B(G146), .ZN(G48));
  INV_X1    g491(.A(new_n585), .ZN(new_n678));
  AOI21_X1  g492(.A(new_n584), .B1(new_n583), .B2(new_n289), .ZN(new_n679));
  INV_X1    g493(.A(new_n592), .ZN(new_n680));
  NOR3_X1   g494(.A1(new_n678), .A2(new_n679), .A3(new_n680), .ZN(new_n681));
  NAND3_X1  g495(.A1(new_n599), .A2(new_n601), .A3(new_n681), .ZN(new_n682));
  INV_X1    g496(.A(new_n365), .ZN(new_n683));
  NAND2_X1  g497(.A1(new_n645), .A2(new_n683), .ZN(new_n684));
  NOR2_X1   g498(.A1(new_n682), .A2(new_n684), .ZN(new_n685));
  NAND2_X1  g499(.A1(new_n685), .A2(new_n612), .ZN(new_n686));
  XNOR2_X1  g500(.A(KEYINPUT41), .B(G113), .ZN(new_n687));
  XNOR2_X1  g501(.A(new_n686), .B(new_n687), .ZN(G15));
  NAND2_X1  g502(.A1(new_n685), .A2(new_n624), .ZN(new_n689));
  XNOR2_X1  g503(.A(new_n689), .B(G116), .ZN(G18));
  INV_X1    g504(.A(new_n682), .ZN(new_n691));
  NAND3_X1  g505(.A1(new_n691), .A2(new_n557), .A3(new_n670), .ZN(new_n692));
  XNOR2_X1  g506(.A(new_n692), .B(G119), .ZN(G21));
  NOR2_X1   g507(.A1(new_n623), .A2(new_n510), .ZN(new_n694));
  AND4_X1   g508(.A1(new_n601), .A2(new_n599), .A3(new_n694), .A4(new_n681), .ZN(new_n695));
  OAI21_X1  g509(.A(new_n412), .B1(new_n408), .B2(new_n448), .ZN(new_n696));
  NAND2_X1  g510(.A1(new_n696), .A2(new_n425), .ZN(new_n697));
  NAND2_X1  g511(.A1(new_n614), .A2(new_n697), .ZN(new_n698));
  NOR3_X1   g512(.A1(new_n698), .A2(new_n365), .A3(new_n556), .ZN(new_n699));
  NAND2_X1  g513(.A1(new_n695), .A2(new_n699), .ZN(new_n700));
  XNOR2_X1  g514(.A(new_n700), .B(G122), .ZN(G24));
  AND4_X1   g515(.A1(new_n601), .A2(new_n599), .A3(new_n671), .A4(new_n681), .ZN(new_n702));
  NOR2_X1   g516(.A1(new_n634), .A2(new_n698), .ZN(new_n703));
  NAND2_X1  g517(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  XNOR2_X1  g518(.A(new_n704), .B(G125), .ZN(G27));
  AOI21_X1  g519(.A(new_n317), .B1(new_n313), .B2(new_n314), .ZN(new_n706));
  NAND4_X1  g520(.A1(new_n706), .A2(new_n458), .A3(new_n593), .A4(new_n671), .ZN(new_n707));
  XNOR2_X1  g521(.A(KEYINPUT104), .B(KEYINPUT42), .ZN(new_n708));
  NAND2_X1  g522(.A1(new_n707), .A2(new_n708), .ZN(new_n709));
  NAND2_X1  g523(.A1(new_n591), .A2(new_n592), .ZN(new_n710));
  AOI211_X1 g524(.A(new_n317), .B(new_n710), .C1(new_n313), .C2(new_n314), .ZN(new_n711));
  INV_X1    g525(.A(KEYINPUT32), .ZN(new_n712));
  NAND2_X1  g526(.A1(new_n454), .A2(new_n712), .ZN(new_n713));
  AOI21_X1  g527(.A(new_n365), .B1(new_n453), .B2(new_n713), .ZN(new_n714));
  NAND4_X1  g528(.A1(new_n711), .A2(KEYINPUT42), .A3(new_n671), .A4(new_n714), .ZN(new_n715));
  NAND2_X1  g529(.A1(new_n709), .A2(new_n715), .ZN(new_n716));
  XNOR2_X1  g530(.A(new_n716), .B(G131), .ZN(G33));
  NAND3_X1  g531(.A1(new_n711), .A2(new_n458), .A3(new_n652), .ZN(new_n718));
  XNOR2_X1  g532(.A(new_n718), .B(G134), .ZN(G36));
  NAND2_X1  g533(.A1(new_n610), .A2(new_n510), .ZN(new_n720));
  XOR2_X1   g534(.A(new_n720), .B(KEYINPUT43), .Z(new_n721));
  NAND3_X1  g535(.A1(new_n721), .A2(new_n615), .A3(new_n647), .ZN(new_n722));
  INV_X1    g536(.A(KEYINPUT44), .ZN(new_n723));
  NAND2_X1  g537(.A1(new_n722), .A2(new_n723), .ZN(new_n724));
  XOR2_X1   g538(.A(new_n724), .B(KEYINPUT107), .Z(new_n725));
  OAI211_X1 g539(.A(new_n725), .B(new_n706), .C1(new_n723), .C2(new_n722), .ZN(new_n726));
  OAI21_X1  g540(.A(new_n587), .B1(new_n588), .B2(new_n569), .ZN(new_n727));
  XNOR2_X1  g541(.A(new_n727), .B(KEYINPUT45), .ZN(new_n728));
  OAI21_X1  g542(.A(G469), .B1(new_n728), .B2(G902), .ZN(new_n729));
  NAND2_X1  g543(.A1(new_n729), .A2(KEYINPUT46), .ZN(new_n730));
  INV_X1    g544(.A(KEYINPUT105), .ZN(new_n731));
  AOI21_X1  g545(.A(new_n678), .B1(new_n730), .B2(new_n731), .ZN(new_n732));
  OR2_X1    g546(.A1(new_n729), .A2(KEYINPUT46), .ZN(new_n733));
  OAI211_X1 g547(.A(new_n732), .B(new_n733), .C1(new_n731), .C2(new_n730), .ZN(new_n734));
  NAND3_X1  g548(.A1(new_n734), .A2(new_n592), .A3(new_n655), .ZN(new_n735));
  XNOR2_X1  g549(.A(new_n735), .B(KEYINPUT106), .ZN(new_n736));
  NOR2_X1   g550(.A1(new_n726), .A2(new_n736), .ZN(new_n737));
  XNOR2_X1  g551(.A(new_n737), .B(new_n373), .ZN(G39));
  NAND2_X1  g552(.A1(new_n734), .A2(new_n592), .ZN(new_n739));
  INV_X1    g553(.A(KEYINPUT47), .ZN(new_n740));
  XNOR2_X1  g554(.A(new_n739), .B(new_n740), .ZN(new_n741));
  INV_X1    g555(.A(new_n706), .ZN(new_n742));
  NOR3_X1   g556(.A1(new_n742), .A2(new_n645), .A3(new_n683), .ZN(new_n743));
  NAND3_X1  g557(.A1(new_n741), .A2(new_n671), .A3(new_n743), .ZN(new_n744));
  XNOR2_X1  g558(.A(new_n744), .B(G140), .ZN(G42));
  INV_X1    g559(.A(KEYINPUT110), .ZN(new_n746));
  INV_X1    g560(.A(KEYINPUT53), .ZN(new_n747));
  NAND2_X1  g561(.A1(new_n548), .A2(new_n510), .ZN(new_n748));
  NAND2_X1  g562(.A1(new_n611), .A2(new_n748), .ZN(new_n749));
  INV_X1    g563(.A(new_n556), .ZN(new_n750));
  AND4_X1   g564(.A1(new_n593), .A2(new_n749), .A3(new_n750), .A4(new_n616), .ZN(new_n751));
  AOI22_X1  g565(.A1(new_n321), .A2(new_n751), .B1(new_n624), .B2(new_n685), .ZN(new_n752));
  NAND2_X1  g566(.A1(new_n752), .A2(new_n636), .ZN(new_n753));
  AOI22_X1  g567(.A1(new_n685), .A2(new_n612), .B1(new_n695), .B2(new_n699), .ZN(new_n754));
  NAND3_X1  g568(.A1(new_n595), .A2(new_n692), .A3(new_n754), .ZN(new_n755));
  NOR2_X1   g569(.A1(new_n753), .A2(new_n755), .ZN(new_n756));
  AOI22_X1  g570(.A1(new_n649), .A2(new_n652), .B1(new_n702), .B2(new_n703), .ZN(new_n757));
  NAND2_X1  g571(.A1(new_n363), .A2(new_n630), .ZN(new_n758));
  NOR3_X1   g572(.A1(new_n665), .A2(new_n758), .A3(new_n651), .ZN(new_n759));
  AND2_X1   g573(.A1(new_n599), .A2(new_n601), .ZN(new_n760));
  NAND4_X1  g574(.A1(new_n759), .A2(new_n593), .A3(new_n760), .A4(new_n694), .ZN(new_n761));
  AOI21_X1  g575(.A(new_n674), .B1(new_n649), .B2(new_n671), .ZN(new_n762));
  INV_X1    g576(.A(new_n671), .ZN(new_n763));
  NOR4_X1   g577(.A1(new_n640), .A2(new_n648), .A3(KEYINPUT103), .A4(new_n763), .ZN(new_n764));
  OAI211_X1 g578(.A(new_n757), .B(new_n761), .C1(new_n762), .C2(new_n764), .ZN(new_n765));
  INV_X1    g579(.A(KEYINPUT109), .ZN(new_n766));
  INV_X1    g580(.A(KEYINPUT52), .ZN(new_n767));
  NAND3_X1  g581(.A1(new_n765), .A2(new_n766), .A3(new_n767), .ZN(new_n768));
  INV_X1    g582(.A(KEYINPUT108), .ZN(new_n769));
  NOR2_X1   g583(.A1(new_n621), .A2(new_n651), .ZN(new_n770));
  NAND3_X1  g584(.A1(new_n706), .A2(new_n593), .A3(new_n770), .ZN(new_n771));
  NAND2_X1  g585(.A1(new_n670), .A2(new_n623), .ZN(new_n772));
  OAI21_X1  g586(.A(new_n769), .B1(new_n771), .B2(new_n772), .ZN(new_n773));
  NOR2_X1   g587(.A1(new_n648), .A2(new_n548), .ZN(new_n774));
  NAND4_X1  g588(.A1(new_n774), .A2(new_n711), .A3(KEYINPUT108), .A4(new_n770), .ZN(new_n775));
  NAND2_X1  g589(.A1(new_n773), .A2(new_n775), .ZN(new_n776));
  AND3_X1   g590(.A1(new_n776), .A2(new_n716), .A3(new_n718), .ZN(new_n777));
  AND2_X1   g591(.A1(new_n711), .A2(new_n671), .ZN(new_n778));
  NAND2_X1  g592(.A1(new_n778), .A2(new_n703), .ZN(new_n779));
  NAND4_X1  g593(.A1(new_n756), .A2(new_n768), .A3(new_n777), .A4(new_n779), .ZN(new_n780));
  NAND2_X1  g594(.A1(new_n765), .A2(new_n767), .ZN(new_n781));
  NAND4_X1  g595(.A1(new_n676), .A2(KEYINPUT52), .A3(new_n757), .A4(new_n761), .ZN(new_n782));
  AND3_X1   g596(.A1(new_n781), .A2(KEYINPUT109), .A3(new_n782), .ZN(new_n783));
  OAI21_X1  g597(.A(new_n747), .B1(new_n780), .B2(new_n783), .ZN(new_n784));
  AND2_X1   g598(.A1(new_n754), .A2(new_n692), .ZN(new_n785));
  NAND4_X1  g599(.A1(new_n785), .A2(new_n752), .A3(new_n595), .A4(new_n636), .ZN(new_n786));
  INV_X1    g600(.A(new_n779), .ZN(new_n787));
  NOR2_X1   g601(.A1(new_n786), .A2(new_n787), .ZN(new_n788));
  NAND2_X1  g602(.A1(new_n781), .A2(new_n782), .ZN(new_n789));
  NAND4_X1  g603(.A1(new_n788), .A2(new_n789), .A3(KEYINPUT53), .A4(new_n777), .ZN(new_n790));
  NAND2_X1  g604(.A1(new_n784), .A2(new_n790), .ZN(new_n791));
  AOI21_X1  g605(.A(new_n746), .B1(new_n791), .B2(KEYINPUT54), .ZN(new_n792));
  INV_X1    g606(.A(KEYINPUT54), .ZN(new_n793));
  AOI211_X1 g607(.A(KEYINPUT110), .B(new_n793), .C1(new_n784), .C2(new_n790), .ZN(new_n794));
  XNOR2_X1  g608(.A(KEYINPUT111), .B(KEYINPUT54), .ZN(new_n795));
  OAI21_X1  g609(.A(KEYINPUT53), .B1(new_n780), .B2(new_n783), .ZN(new_n796));
  NAND4_X1  g610(.A1(new_n788), .A2(new_n789), .A3(new_n747), .A4(new_n777), .ZN(new_n797));
  AOI21_X1  g611(.A(new_n795), .B1(new_n796), .B2(new_n797), .ZN(new_n798));
  NOR3_X1   g612(.A1(new_n792), .A2(new_n794), .A3(new_n798), .ZN(new_n799));
  AND2_X1   g613(.A1(new_n706), .A2(new_n681), .ZN(new_n800));
  NAND4_X1  g614(.A1(new_n800), .A2(new_n683), .A3(new_n551), .A4(new_n665), .ZN(new_n801));
  XNOR2_X1  g615(.A(new_n801), .B(KEYINPUT113), .ZN(new_n802));
  NOR2_X1   g616(.A1(new_n802), .A2(new_n611), .ZN(new_n803));
  AND2_X1   g617(.A1(new_n721), .A2(new_n551), .ZN(new_n804));
  AND2_X1   g618(.A1(new_n804), .A2(new_n800), .ZN(new_n805));
  NAND2_X1  g619(.A1(new_n805), .A2(new_n714), .ZN(new_n806));
  XNOR2_X1  g620(.A(new_n806), .B(KEYINPUT48), .ZN(new_n807));
  NAND3_X1  g621(.A1(new_n807), .A2(G952), .A3(new_n351), .ZN(new_n808));
  NAND4_X1  g622(.A1(new_n804), .A2(new_n683), .A3(new_n614), .A4(new_n697), .ZN(new_n809));
  INV_X1    g623(.A(new_n809), .ZN(new_n810));
  NAND4_X1  g624(.A1(new_n810), .A2(new_n317), .A3(new_n659), .A4(new_n681), .ZN(new_n811));
  OR2_X1    g625(.A1(KEYINPUT112), .A2(KEYINPUT50), .ZN(new_n812));
  NOR2_X1   g626(.A1(new_n811), .A2(new_n812), .ZN(new_n813));
  XOR2_X1   g627(.A(KEYINPUT112), .B(KEYINPUT50), .Z(new_n814));
  AOI21_X1  g628(.A(new_n813), .B1(new_n814), .B2(new_n811), .ZN(new_n815));
  NOR3_X1   g629(.A1(new_n678), .A2(new_n679), .A3(new_n592), .ZN(new_n816));
  OAI211_X1 g630(.A(new_n706), .B(new_n810), .C1(new_n741), .C2(new_n816), .ZN(new_n817));
  NAND2_X1  g631(.A1(new_n805), .A2(new_n703), .ZN(new_n818));
  OR3_X1    g632(.A1(new_n802), .A2(new_n511), .A3(new_n610), .ZN(new_n819));
  NAND4_X1  g633(.A1(new_n815), .A2(new_n817), .A3(new_n818), .A4(new_n819), .ZN(new_n820));
  INV_X1    g634(.A(KEYINPUT51), .ZN(new_n821));
  AOI211_X1 g635(.A(new_n803), .B(new_n808), .C1(new_n820), .C2(new_n821), .ZN(new_n822));
  OAI211_X1 g636(.A(new_n799), .B(new_n822), .C1(new_n821), .C2(new_n820), .ZN(new_n823));
  NAND2_X1  g637(.A1(new_n810), .A2(new_n691), .ZN(new_n824));
  XNOR2_X1  g638(.A(new_n824), .B(KEYINPUT114), .ZN(new_n825));
  OAI22_X1  g639(.A1(new_n823), .A2(new_n825), .B1(G952), .B2(G953), .ZN(new_n826));
  NOR2_X1   g640(.A1(new_n678), .A2(new_n679), .ZN(new_n827));
  XOR2_X1   g641(.A(new_n827), .B(KEYINPUT49), .Z(new_n828));
  NOR4_X1   g642(.A1(new_n828), .A2(new_n365), .A3(new_n317), .A4(new_n680), .ZN(new_n829));
  NAND4_X1  g643(.A1(new_n829), .A2(new_n510), .A3(new_n610), .A4(new_n659), .ZN(new_n830));
  OAI21_X1  g644(.A(new_n826), .B1(new_n664), .B2(new_n830), .ZN(G75));
  NOR2_X1   g645(.A1(new_n351), .A2(G952), .ZN(new_n832));
  AND2_X1   g646(.A1(new_n297), .A2(new_n299), .ZN(new_n833));
  XNOR2_X1  g647(.A(new_n833), .B(new_n300), .ZN(new_n834));
  XNOR2_X1  g648(.A(new_n834), .B(KEYINPUT55), .ZN(new_n835));
  NAND4_X1  g649(.A1(new_n796), .A2(G210), .A3(G902), .A4(new_n797), .ZN(new_n836));
  INV_X1    g650(.A(KEYINPUT56), .ZN(new_n837));
  NAND2_X1  g651(.A1(new_n836), .A2(new_n837), .ZN(new_n838));
  AOI21_X1  g652(.A(new_n835), .B1(new_n838), .B2(KEYINPUT115), .ZN(new_n839));
  XNOR2_X1  g653(.A(new_n838), .B(KEYINPUT115), .ZN(new_n840));
  AOI211_X1 g654(.A(new_n832), .B(new_n839), .C1(new_n840), .C2(new_n835), .ZN(G51));
  XNOR2_X1  g655(.A(new_n583), .B(KEYINPUT116), .ZN(new_n842));
  AND3_X1   g656(.A1(new_n796), .A2(new_n795), .A3(new_n797), .ZN(new_n843));
  NOR2_X1   g657(.A1(new_n843), .A2(new_n798), .ZN(new_n844));
  XNOR2_X1  g658(.A(new_n590), .B(KEYINPUT57), .ZN(new_n845));
  OAI21_X1  g659(.A(new_n842), .B1(new_n844), .B2(new_n845), .ZN(new_n846));
  AND3_X1   g660(.A1(new_n796), .A2(G902), .A3(new_n797), .ZN(new_n847));
  NAND3_X1  g661(.A1(new_n847), .A2(G469), .A3(new_n728), .ZN(new_n848));
  AOI21_X1  g662(.A(new_n832), .B1(new_n846), .B2(new_n848), .ZN(G54));
  AND2_X1   g663(.A1(new_n847), .A2(KEYINPUT58), .ZN(new_n850));
  AOI21_X1  g664(.A(new_n501), .B1(new_n850), .B2(G475), .ZN(new_n851));
  NAND3_X1  g665(.A1(new_n850), .A2(G475), .A3(new_n501), .ZN(new_n852));
  INV_X1    g666(.A(KEYINPUT117), .ZN(new_n853));
  OR2_X1    g667(.A1(new_n852), .A2(new_n853), .ZN(new_n854));
  NAND2_X1  g668(.A1(new_n852), .A2(new_n853), .ZN(new_n855));
  AOI211_X1 g669(.A(new_n832), .B(new_n851), .C1(new_n854), .C2(new_n855), .ZN(G60));
  AND2_X1   g670(.A1(new_n603), .A2(new_n606), .ZN(new_n857));
  NAND2_X1  g671(.A1(G478), .A2(G902), .ZN(new_n858));
  XOR2_X1   g672(.A(new_n858), .B(KEYINPUT59), .Z(new_n859));
  OAI21_X1  g673(.A(new_n857), .B1(new_n799), .B2(new_n859), .ZN(new_n860));
  INV_X1    g674(.A(new_n832), .ZN(new_n861));
  OR3_X1    g675(.A1(new_n844), .A2(new_n857), .A3(new_n859), .ZN(new_n862));
  NAND3_X1  g676(.A1(new_n860), .A2(new_n861), .A3(new_n862), .ZN(new_n863));
  NAND2_X1  g677(.A1(new_n863), .A2(KEYINPUT118), .ZN(new_n864));
  INV_X1    g678(.A(KEYINPUT118), .ZN(new_n865));
  NAND4_X1  g679(.A1(new_n860), .A2(new_n865), .A3(new_n861), .A4(new_n862), .ZN(new_n866));
  NAND2_X1  g680(.A1(new_n864), .A2(new_n866), .ZN(G63));
  NAND2_X1  g681(.A1(G217), .A2(G902), .ZN(new_n868));
  XOR2_X1   g682(.A(new_n868), .B(KEYINPUT60), .Z(new_n869));
  NAND3_X1  g683(.A1(new_n796), .A2(new_n797), .A3(new_n869), .ZN(new_n870));
  INV_X1    g684(.A(KEYINPUT119), .ZN(new_n871));
  NAND2_X1  g685(.A1(new_n870), .A2(new_n871), .ZN(new_n872));
  NAND4_X1  g686(.A1(new_n796), .A2(KEYINPUT119), .A3(new_n797), .A4(new_n869), .ZN(new_n873));
  NAND2_X1  g687(.A1(new_n872), .A2(new_n873), .ZN(new_n874));
  AOI21_X1  g688(.A(new_n832), .B1(new_n874), .B2(new_n629), .ZN(new_n875));
  NAND2_X1  g689(.A1(new_n355), .A2(new_n356), .ZN(new_n876));
  NAND3_X1  g690(.A1(new_n872), .A2(new_n876), .A3(new_n873), .ZN(new_n877));
  NAND2_X1  g691(.A1(new_n877), .A2(KEYINPUT120), .ZN(new_n878));
  INV_X1    g692(.A(KEYINPUT120), .ZN(new_n879));
  NAND4_X1  g693(.A1(new_n872), .A2(new_n879), .A3(new_n876), .A4(new_n873), .ZN(new_n880));
  NAND4_X1  g694(.A1(new_n875), .A2(new_n878), .A3(KEYINPUT61), .A4(new_n880), .ZN(new_n881));
  INV_X1    g695(.A(KEYINPUT121), .ZN(new_n882));
  NAND2_X1  g696(.A1(new_n881), .A2(new_n882), .ZN(new_n883));
  AND2_X1   g697(.A1(new_n880), .A2(KEYINPUT61), .ZN(new_n884));
  NAND4_X1  g698(.A1(new_n884), .A2(KEYINPUT121), .A3(new_n875), .A4(new_n878), .ZN(new_n885));
  NAND2_X1  g699(.A1(new_n883), .A2(new_n885), .ZN(new_n886));
  AND2_X1   g700(.A1(new_n875), .A2(new_n877), .ZN(new_n887));
  OR2_X1    g701(.A1(new_n887), .A2(KEYINPUT61), .ZN(new_n888));
  NAND2_X1  g702(.A1(new_n886), .A2(new_n888), .ZN(G66));
  NOR2_X1   g703(.A1(new_n756), .A2(G953), .ZN(new_n890));
  XNOR2_X1  g704(.A(new_n890), .B(KEYINPUT122), .ZN(new_n891));
  OAI21_X1  g705(.A(G953), .B1(new_n553), .B2(new_n212), .ZN(new_n892));
  NAND2_X1  g706(.A1(new_n891), .A2(new_n892), .ZN(new_n893));
  XNOR2_X1  g707(.A(new_n893), .B(KEYINPUT123), .ZN(new_n894));
  INV_X1    g708(.A(G898), .ZN(new_n895));
  AOI21_X1  g709(.A(new_n833), .B1(new_n895), .B2(G953), .ZN(new_n896));
  XNOR2_X1  g710(.A(new_n894), .B(new_n896), .ZN(G69));
  NAND2_X1  g711(.A1(new_n393), .A2(new_n396), .ZN(new_n898));
  XOR2_X1   g712(.A(new_n898), .B(new_n497), .Z(new_n899));
  NAND2_X1  g713(.A1(G900), .A2(G953), .ZN(new_n900));
  NAND2_X1  g714(.A1(new_n676), .A2(new_n757), .ZN(new_n901));
  INV_X1    g715(.A(KEYINPUT124), .ZN(new_n902));
  XNOR2_X1  g716(.A(new_n901), .B(new_n902), .ZN(new_n903));
  AND3_X1   g717(.A1(new_n744), .A2(new_n716), .A3(new_n718), .ZN(new_n904));
  NAND3_X1  g718(.A1(new_n760), .A2(new_n714), .A3(new_n694), .ZN(new_n905));
  AND2_X1   g719(.A1(new_n726), .A2(new_n905), .ZN(new_n906));
  OAI211_X1 g720(.A(new_n903), .B(new_n904), .C1(new_n906), .C2(new_n736), .ZN(new_n907));
  OAI211_X1 g721(.A(new_n899), .B(new_n900), .C1(new_n907), .C2(G953), .ZN(new_n908));
  NAND2_X1  g722(.A1(new_n667), .A2(new_n903), .ZN(new_n909));
  XNOR2_X1  g723(.A(new_n909), .B(KEYINPUT62), .ZN(new_n910));
  INV_X1    g724(.A(new_n744), .ZN(new_n911));
  NOR2_X1   g725(.A1(new_n910), .A2(new_n911), .ZN(new_n912));
  AOI211_X1 g726(.A(new_n742), .B(new_n657), .C1(new_n611), .C2(new_n748), .ZN(new_n913));
  AOI21_X1  g727(.A(new_n737), .B1(new_n458), .B2(new_n913), .ZN(new_n914));
  AOI21_X1  g728(.A(G953), .B1(new_n912), .B2(new_n914), .ZN(new_n915));
  OAI21_X1  g729(.A(new_n908), .B1(new_n915), .B2(new_n899), .ZN(new_n916));
  AOI21_X1  g730(.A(new_n351), .B1(G227), .B2(G900), .ZN(new_n917));
  XNOR2_X1  g731(.A(new_n916), .B(new_n917), .ZN(G72));
  XOR2_X1   g732(.A(KEYINPUT125), .B(KEYINPUT63), .Z(new_n919));
  AND2_X1   g733(.A1(G472), .A2(G902), .ZN(new_n920));
  XNOR2_X1  g734(.A(new_n919), .B(new_n920), .ZN(new_n921));
  XNOR2_X1  g735(.A(new_n921), .B(KEYINPUT126), .ZN(new_n922));
  OAI21_X1  g736(.A(new_n922), .B1(new_n907), .B2(new_n786), .ZN(new_n923));
  XOR2_X1   g737(.A(new_n403), .B(KEYINPUT127), .Z(new_n924));
  NAND3_X1  g738(.A1(new_n923), .A2(new_n410), .A3(new_n924), .ZN(new_n925));
  XNOR2_X1  g739(.A(new_n403), .B(new_n408), .ZN(new_n926));
  NAND3_X1  g740(.A1(new_n791), .A2(new_n921), .A3(new_n926), .ZN(new_n927));
  NAND3_X1  g741(.A1(new_n925), .A2(new_n861), .A3(new_n927), .ZN(new_n928));
  NAND3_X1  g742(.A1(new_n912), .A2(new_n756), .A3(new_n914), .ZN(new_n929));
  AOI21_X1  g743(.A(new_n924), .B1(new_n929), .B2(new_n922), .ZN(new_n930));
  AOI21_X1  g744(.A(new_n928), .B1(new_n408), .B2(new_n930), .ZN(G57));
endmodule


