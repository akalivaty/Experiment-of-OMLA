//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 1 1 1 0 1 0 0 1 1 0 1 0 1 0 1 1 0 1 0 0 0 0 1 0 1 1 0 1 0 1 1 1 1 1 1 0 0 0 1 1 1 1 1 0 1 1 0 0 1 1 0 0 0 1 1 1 1 1 1 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:19:40 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n693, new_n694, new_n695, new_n696, new_n697, new_n699, new_n700,
    new_n701, new_n703, new_n704, new_n705, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n737, new_n738,
    new_n739, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n770,
    new_n771, new_n772, new_n773, new_n775, new_n776, new_n777, new_n778,
    new_n779, new_n781, new_n782, new_n784, new_n785, new_n786, new_n787,
    new_n788, new_n789, new_n790, new_n791, new_n792, new_n793, new_n794,
    new_n795, new_n796, new_n797, new_n798, new_n799, new_n800, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n813, new_n814, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n880, new_n881, new_n883, new_n884,
    new_n885, new_n886, new_n887, new_n889, new_n890, new_n891, new_n892,
    new_n893, new_n894, new_n895, new_n896, new_n897, new_n898, new_n899,
    new_n900, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n938, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n948, new_n949, new_n951,
    new_n952, new_n953, new_n955, new_n956, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n977, new_n978, new_n979, new_n981, new_n982, new_n983,
    new_n985, new_n986, new_n987, new_n988, new_n989, new_n990, new_n991,
    new_n992, new_n994, new_n995, new_n996, new_n997, new_n998, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014;
  XNOR2_X1  g000(.A(G8gat), .B(G36gat), .ZN(new_n202));
  XNOR2_X1  g001(.A(G64gat), .B(G92gat), .ZN(new_n203));
  XOR2_X1   g002(.A(new_n202), .B(new_n203), .Z(new_n204));
  INV_X1    g003(.A(new_n204), .ZN(new_n205));
  NAND2_X1  g004(.A1(G226gat), .A2(G233gat), .ZN(new_n206));
  INV_X1    g005(.A(new_n206), .ZN(new_n207));
  NOR2_X1   g006(.A1(G169gat), .A2(G176gat), .ZN(new_n208));
  INV_X1    g007(.A(KEYINPUT23), .ZN(new_n209));
  NAND2_X1  g008(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  OAI21_X1  g009(.A(KEYINPUT23), .B1(G169gat), .B2(G176gat), .ZN(new_n211));
  NAND2_X1  g010(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  AND2_X1   g011(.A1(G183gat), .A2(G190gat), .ZN(new_n213));
  INV_X1    g012(.A(KEYINPUT24), .ZN(new_n214));
  AOI22_X1  g013(.A1(new_n213), .A2(new_n214), .B1(G169gat), .B2(G176gat), .ZN(new_n215));
  INV_X1    g014(.A(G183gat), .ZN(new_n216));
  INV_X1    g015(.A(G190gat), .ZN(new_n217));
  NAND2_X1  g016(.A1(new_n216), .A2(new_n217), .ZN(new_n218));
  NAND2_X1  g017(.A1(G183gat), .A2(G190gat), .ZN(new_n219));
  NAND3_X1  g018(.A1(new_n218), .A2(KEYINPUT24), .A3(new_n219), .ZN(new_n220));
  NAND3_X1  g019(.A1(new_n212), .A2(new_n215), .A3(new_n220), .ZN(new_n221));
  INV_X1    g020(.A(KEYINPUT25), .ZN(new_n222));
  NAND2_X1  g021(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  NAND4_X1  g022(.A1(new_n212), .A2(new_n215), .A3(new_n220), .A4(KEYINPUT25), .ZN(new_n224));
  AND2_X1   g023(.A1(new_n223), .A2(new_n224), .ZN(new_n225));
  NAND2_X1  g024(.A1(new_n208), .A2(KEYINPUT26), .ZN(new_n226));
  INV_X1    g025(.A(KEYINPUT26), .ZN(new_n227));
  INV_X1    g026(.A(G169gat), .ZN(new_n228));
  INV_X1    g027(.A(G176gat), .ZN(new_n229));
  OAI21_X1  g028(.A(new_n227), .B1(new_n228), .B2(new_n229), .ZN(new_n230));
  OAI211_X1 g029(.A(new_n219), .B(new_n226), .C1(new_n230), .C2(new_n208), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n216), .A2(KEYINPUT27), .ZN(new_n232));
  INV_X1    g031(.A(KEYINPUT27), .ZN(new_n233));
  NAND2_X1  g032(.A1(new_n233), .A2(G183gat), .ZN(new_n234));
  NAND3_X1  g033(.A1(new_n232), .A2(new_n234), .A3(new_n217), .ZN(new_n235));
  INV_X1    g034(.A(KEYINPUT65), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n235), .A2(new_n236), .ZN(new_n237));
  XNOR2_X1  g036(.A(KEYINPUT27), .B(G183gat), .ZN(new_n238));
  NAND3_X1  g037(.A1(new_n238), .A2(KEYINPUT65), .A3(new_n217), .ZN(new_n239));
  XOR2_X1   g038(.A(KEYINPUT66), .B(KEYINPUT28), .Z(new_n240));
  NAND3_X1  g039(.A1(new_n237), .A2(new_n239), .A3(new_n240), .ZN(new_n241));
  NAND2_X1  g040(.A1(new_n232), .A2(new_n234), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n242), .A2(KEYINPUT67), .ZN(new_n243));
  INV_X1    g042(.A(KEYINPUT67), .ZN(new_n244));
  NAND2_X1  g043(.A1(new_n238), .A2(new_n244), .ZN(new_n245));
  NAND4_X1  g044(.A1(new_n243), .A2(new_n245), .A3(KEYINPUT28), .A4(new_n217), .ZN(new_n246));
  AOI21_X1  g045(.A(new_n231), .B1(new_n241), .B2(new_n246), .ZN(new_n247));
  OAI21_X1  g046(.A(new_n207), .B1(new_n225), .B2(new_n247), .ZN(new_n248));
  XOR2_X1   g047(.A(G211gat), .B(G218gat), .Z(new_n249));
  NAND2_X1  g048(.A1(new_n249), .A2(KEYINPUT73), .ZN(new_n250));
  INV_X1    g049(.A(G204gat), .ZN(new_n251));
  AND2_X1   g050(.A1(KEYINPUT72), .A2(G197gat), .ZN(new_n252));
  NOR2_X1   g051(.A1(KEYINPUT72), .A2(G197gat), .ZN(new_n253));
  OAI21_X1  g052(.A(new_n251), .B1(new_n252), .B2(new_n253), .ZN(new_n254));
  INV_X1    g053(.A(KEYINPUT72), .ZN(new_n255));
  INV_X1    g054(.A(G197gat), .ZN(new_n256));
  NAND2_X1  g055(.A1(new_n255), .A2(new_n256), .ZN(new_n257));
  NAND2_X1  g056(.A1(KEYINPUT72), .A2(G197gat), .ZN(new_n258));
  NAND3_X1  g057(.A1(new_n257), .A2(G204gat), .A3(new_n258), .ZN(new_n259));
  NAND2_X1  g058(.A1(new_n254), .A2(new_n259), .ZN(new_n260));
  NAND2_X1  g059(.A1(G211gat), .A2(G218gat), .ZN(new_n261));
  INV_X1    g060(.A(KEYINPUT22), .ZN(new_n262));
  NAND2_X1  g061(.A1(new_n261), .A2(new_n262), .ZN(new_n263));
  AND3_X1   g062(.A1(new_n250), .A2(new_n260), .A3(new_n263), .ZN(new_n264));
  AOI21_X1  g063(.A(new_n250), .B1(new_n263), .B2(new_n260), .ZN(new_n265));
  NOR2_X1   g064(.A1(new_n264), .A2(new_n265), .ZN(new_n266));
  INV_X1    g065(.A(new_n266), .ZN(new_n267));
  INV_X1    g066(.A(new_n231), .ZN(new_n268));
  AND3_X1   g067(.A1(new_n237), .A2(new_n239), .A3(new_n240), .ZN(new_n269));
  AND2_X1   g068(.A1(new_n217), .A2(KEYINPUT28), .ZN(new_n270));
  AND3_X1   g069(.A1(new_n243), .A2(new_n245), .A3(new_n270), .ZN(new_n271));
  OAI21_X1  g070(.A(new_n268), .B1(new_n269), .B2(new_n271), .ZN(new_n272));
  NAND2_X1  g071(.A1(new_n223), .A2(new_n224), .ZN(new_n273));
  AOI21_X1  g072(.A(KEYINPUT29), .B1(new_n272), .B2(new_n273), .ZN(new_n274));
  OAI211_X1 g073(.A(new_n248), .B(new_n267), .C1(new_n274), .C2(new_n207), .ZN(new_n275));
  INV_X1    g074(.A(new_n275), .ZN(new_n276));
  INV_X1    g075(.A(KEYINPUT29), .ZN(new_n277));
  OAI21_X1  g076(.A(new_n277), .B1(new_n225), .B2(new_n247), .ZN(new_n278));
  NAND2_X1  g077(.A1(new_n278), .A2(new_n206), .ZN(new_n279));
  AOI21_X1  g078(.A(new_n267), .B1(new_n279), .B2(new_n248), .ZN(new_n280));
  OAI21_X1  g079(.A(new_n205), .B1(new_n276), .B2(new_n280), .ZN(new_n281));
  OAI21_X1  g080(.A(new_n248), .B1(new_n274), .B2(new_n207), .ZN(new_n282));
  NAND2_X1  g081(.A1(new_n282), .A2(new_n266), .ZN(new_n283));
  NAND3_X1  g082(.A1(new_n283), .A2(new_n204), .A3(new_n275), .ZN(new_n284));
  NAND3_X1  g083(.A1(new_n281), .A2(KEYINPUT30), .A3(new_n284), .ZN(new_n285));
  INV_X1    g084(.A(KEYINPUT30), .ZN(new_n286));
  NAND4_X1  g085(.A1(new_n283), .A2(new_n286), .A3(new_n204), .A4(new_n275), .ZN(new_n287));
  NAND2_X1  g086(.A1(new_n285), .A2(new_n287), .ZN(new_n288));
  XOR2_X1   g087(.A(KEYINPUT69), .B(G113gat), .Z(new_n289));
  NAND2_X1  g088(.A1(new_n289), .A2(G120gat), .ZN(new_n290));
  INV_X1    g089(.A(G113gat), .ZN(new_n291));
  INV_X1    g090(.A(G120gat), .ZN(new_n292));
  AOI22_X1  g091(.A1(new_n291), .A2(new_n292), .B1(KEYINPUT70), .B2(KEYINPUT1), .ZN(new_n293));
  OR2_X1    g092(.A1(KEYINPUT70), .A2(KEYINPUT1), .ZN(new_n294));
  AND2_X1   g093(.A1(new_n293), .A2(new_n294), .ZN(new_n295));
  XNOR2_X1  g094(.A(G127gat), .B(G134gat), .ZN(new_n296));
  NAND3_X1  g095(.A1(new_n290), .A2(new_n295), .A3(new_n296), .ZN(new_n297));
  INV_X1    g096(.A(G155gat), .ZN(new_n298));
  INV_X1    g097(.A(G162gat), .ZN(new_n299));
  INV_X1    g098(.A(KEYINPUT2), .ZN(new_n300));
  OAI211_X1 g099(.A(new_n298), .B(new_n299), .C1(new_n300), .C2(KEYINPUT75), .ZN(new_n301));
  NAND2_X1  g100(.A1(G155gat), .A2(G162gat), .ZN(new_n302));
  NAND2_X1  g101(.A1(new_n301), .A2(new_n302), .ZN(new_n303));
  XOR2_X1   g102(.A(G141gat), .B(G148gat), .Z(new_n304));
  NAND2_X1  g103(.A1(new_n302), .A2(KEYINPUT2), .ZN(new_n305));
  NAND2_X1  g104(.A1(new_n305), .A2(KEYINPUT75), .ZN(new_n306));
  NAND3_X1  g105(.A1(new_n303), .A2(new_n304), .A3(new_n306), .ZN(new_n307));
  INV_X1    g106(.A(G141gat), .ZN(new_n308));
  INV_X1    g107(.A(G148gat), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n308), .A2(new_n309), .ZN(new_n310));
  NAND2_X1  g109(.A1(G141gat), .A2(G148gat), .ZN(new_n311));
  NAND3_X1  g110(.A1(new_n305), .A2(new_n310), .A3(new_n311), .ZN(new_n312));
  NAND3_X1  g111(.A1(new_n298), .A2(new_n299), .A3(KEYINPUT74), .ZN(new_n313));
  INV_X1    g112(.A(KEYINPUT74), .ZN(new_n314));
  OAI21_X1  g113(.A(new_n314), .B1(G155gat), .B2(G162gat), .ZN(new_n315));
  NAND4_X1  g114(.A1(new_n312), .A2(new_n302), .A3(new_n313), .A4(new_n315), .ZN(new_n316));
  OR2_X1    g115(.A1(KEYINPUT68), .A2(G134gat), .ZN(new_n317));
  NAND2_X1  g116(.A1(KEYINPUT68), .A2(G134gat), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n317), .A2(new_n318), .ZN(new_n319));
  NAND2_X1  g118(.A1(new_n319), .A2(G127gat), .ZN(new_n320));
  NAND2_X1  g119(.A1(new_n291), .A2(new_n292), .ZN(new_n321));
  INV_X1    g120(.A(KEYINPUT1), .ZN(new_n322));
  NAND2_X1  g121(.A1(G113gat), .A2(G120gat), .ZN(new_n323));
  NAND3_X1  g122(.A1(new_n321), .A2(new_n322), .A3(new_n323), .ZN(new_n324));
  OR2_X1    g123(.A1(G127gat), .A2(G134gat), .ZN(new_n325));
  NAND3_X1  g124(.A1(new_n320), .A2(new_n324), .A3(new_n325), .ZN(new_n326));
  NAND4_X1  g125(.A1(new_n297), .A2(new_n307), .A3(new_n316), .A4(new_n326), .ZN(new_n327));
  XNOR2_X1  g126(.A(new_n327), .B(KEYINPUT4), .ZN(new_n328));
  NAND2_X1  g127(.A1(G225gat), .A2(G233gat), .ZN(new_n329));
  NAND2_X1  g128(.A1(new_n316), .A2(new_n307), .ZN(new_n330));
  NAND2_X1  g129(.A1(new_n330), .A2(KEYINPUT3), .ZN(new_n331));
  INV_X1    g130(.A(KEYINPUT3), .ZN(new_n332));
  NAND3_X1  g131(.A1(new_n316), .A2(new_n307), .A3(new_n332), .ZN(new_n333));
  NAND3_X1  g132(.A1(new_n296), .A2(new_n294), .A3(new_n293), .ZN(new_n334));
  XNOR2_X1  g133(.A(KEYINPUT69), .B(G113gat), .ZN(new_n335));
  NOR2_X1   g134(.A1(new_n335), .A2(new_n292), .ZN(new_n336));
  OAI21_X1  g135(.A(new_n322), .B1(G113gat), .B2(G120gat), .ZN(new_n337));
  INV_X1    g136(.A(new_n323), .ZN(new_n338));
  OAI21_X1  g137(.A(new_n325), .B1(new_n337), .B2(new_n338), .ZN(new_n339));
  INV_X1    g138(.A(G127gat), .ZN(new_n340));
  AOI21_X1  g139(.A(new_n340), .B1(new_n317), .B2(new_n318), .ZN(new_n341));
  OAI22_X1  g140(.A1(new_n334), .A2(new_n336), .B1(new_n339), .B2(new_n341), .ZN(new_n342));
  NAND3_X1  g141(.A1(new_n331), .A2(new_n333), .A3(new_n342), .ZN(new_n343));
  NAND4_X1  g142(.A1(new_n328), .A2(KEYINPUT5), .A3(new_n329), .A4(new_n343), .ZN(new_n344));
  INV_X1    g143(.A(new_n329), .ZN(new_n345));
  NOR2_X1   g144(.A1(new_n330), .A2(new_n342), .ZN(new_n346));
  AOI22_X1  g145(.A1(new_n297), .A2(new_n326), .B1(new_n307), .B2(new_n316), .ZN(new_n347));
  OAI21_X1  g146(.A(new_n345), .B1(new_n346), .B2(new_n347), .ZN(new_n348));
  NAND2_X1  g147(.A1(new_n348), .A2(KEYINPUT5), .ZN(new_n349));
  NAND2_X1  g148(.A1(new_n346), .A2(KEYINPUT4), .ZN(new_n350));
  INV_X1    g149(.A(KEYINPUT4), .ZN(new_n351));
  NAND2_X1  g150(.A1(new_n327), .A2(new_n351), .ZN(new_n352));
  NAND4_X1  g151(.A1(new_n350), .A2(new_n343), .A3(new_n352), .A4(new_n329), .ZN(new_n353));
  NAND2_X1  g152(.A1(new_n349), .A2(new_n353), .ZN(new_n354));
  NAND2_X1  g153(.A1(new_n344), .A2(new_n354), .ZN(new_n355));
  XNOR2_X1  g154(.A(G1gat), .B(G29gat), .ZN(new_n356));
  XNOR2_X1  g155(.A(new_n356), .B(KEYINPUT0), .ZN(new_n357));
  XNOR2_X1  g156(.A(G57gat), .B(G85gat), .ZN(new_n358));
  XOR2_X1   g157(.A(new_n357), .B(new_n358), .Z(new_n359));
  AOI21_X1  g158(.A(KEYINPUT6), .B1(new_n355), .B2(new_n359), .ZN(new_n360));
  INV_X1    g159(.A(new_n359), .ZN(new_n361));
  NAND3_X1  g160(.A1(new_n344), .A2(new_n354), .A3(new_n361), .ZN(new_n362));
  NAND2_X1  g161(.A1(new_n360), .A2(new_n362), .ZN(new_n363));
  INV_X1    g162(.A(KEYINPUT6), .ZN(new_n364));
  NOR2_X1   g163(.A1(new_n362), .A2(new_n364), .ZN(new_n365));
  INV_X1    g164(.A(new_n365), .ZN(new_n366));
  NAND2_X1  g165(.A1(new_n363), .A2(new_n366), .ZN(new_n367));
  INV_X1    g166(.A(KEYINPUT35), .ZN(new_n368));
  INV_X1    g167(.A(new_n342), .ZN(new_n369));
  OAI21_X1  g168(.A(new_n369), .B1(new_n225), .B2(new_n247), .ZN(new_n370));
  NAND3_X1  g169(.A1(new_n272), .A2(new_n273), .A3(new_n342), .ZN(new_n371));
  NAND2_X1  g170(.A1(G227gat), .A2(G233gat), .ZN(new_n372));
  XNOR2_X1  g171(.A(new_n372), .B(KEYINPUT64), .ZN(new_n373));
  NAND3_X1  g172(.A1(new_n370), .A2(new_n371), .A3(new_n373), .ZN(new_n374));
  INV_X1    g173(.A(KEYINPUT32), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n375), .A2(KEYINPUT33), .ZN(new_n376));
  NAND2_X1  g175(.A1(new_n374), .A2(new_n376), .ZN(new_n377));
  XNOR2_X1  g176(.A(G15gat), .B(G43gat), .ZN(new_n378));
  XNOR2_X1  g177(.A(G71gat), .B(G99gat), .ZN(new_n379));
  XOR2_X1   g178(.A(new_n378), .B(new_n379), .Z(new_n380));
  NAND2_X1  g179(.A1(new_n377), .A2(new_n380), .ZN(new_n381));
  AOI21_X1  g180(.A(new_n375), .B1(new_n380), .B2(KEYINPUT33), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n374), .A2(new_n382), .ZN(new_n383));
  NAND2_X1  g182(.A1(new_n383), .A2(KEYINPUT71), .ZN(new_n384));
  INV_X1    g183(.A(KEYINPUT71), .ZN(new_n385));
  NAND3_X1  g184(.A1(new_n374), .A2(new_n385), .A3(new_n382), .ZN(new_n386));
  NAND3_X1  g185(.A1(new_n381), .A2(new_n384), .A3(new_n386), .ZN(new_n387));
  INV_X1    g186(.A(KEYINPUT34), .ZN(new_n388));
  NAND2_X1  g187(.A1(new_n370), .A2(new_n371), .ZN(new_n389));
  INV_X1    g188(.A(new_n373), .ZN(new_n390));
  AOI21_X1  g189(.A(new_n388), .B1(new_n389), .B2(new_n390), .ZN(new_n391));
  AOI211_X1 g190(.A(KEYINPUT34), .B(new_n373), .C1(new_n370), .C2(new_n371), .ZN(new_n392));
  OR2_X1    g191(.A1(new_n391), .A2(new_n392), .ZN(new_n393));
  NOR2_X1   g192(.A1(new_n387), .A2(new_n393), .ZN(new_n394));
  NOR2_X1   g193(.A1(new_n391), .A2(new_n392), .ZN(new_n395));
  INV_X1    g194(.A(new_n380), .ZN(new_n396));
  AOI21_X1  g195(.A(new_n396), .B1(new_n374), .B2(new_n376), .ZN(new_n397));
  AOI21_X1  g196(.A(new_n385), .B1(new_n374), .B2(new_n382), .ZN(new_n398));
  NOR2_X1   g197(.A1(new_n397), .A2(new_n398), .ZN(new_n399));
  AOI21_X1  g198(.A(new_n395), .B1(new_n399), .B2(new_n386), .ZN(new_n400));
  NOR2_X1   g199(.A1(new_n394), .A2(new_n400), .ZN(new_n401));
  NAND2_X1  g200(.A1(new_n333), .A2(new_n277), .ZN(new_n402));
  NAND2_X1  g201(.A1(new_n266), .A2(new_n402), .ZN(new_n403));
  INV_X1    g202(.A(G228gat), .ZN(new_n404));
  INV_X1    g203(.A(G233gat), .ZN(new_n405));
  NOR2_X1   g204(.A1(new_n404), .A2(new_n405), .ZN(new_n406));
  NAND2_X1  g205(.A1(new_n403), .A2(new_n406), .ZN(new_n407));
  INV_X1    g206(.A(new_n330), .ZN(new_n408));
  OAI21_X1  g207(.A(new_n277), .B1(new_n264), .B2(new_n265), .ZN(new_n409));
  AOI21_X1  g208(.A(new_n408), .B1(new_n409), .B2(new_n332), .ZN(new_n410));
  NOR2_X1   g209(.A1(new_n407), .A2(new_n410), .ZN(new_n411));
  AOI22_X1  g210(.A1(new_n254), .A2(new_n259), .B1(new_n262), .B2(new_n261), .ZN(new_n412));
  OAI21_X1  g211(.A(new_n277), .B1(new_n412), .B2(new_n249), .ZN(new_n413));
  AND3_X1   g212(.A1(new_n260), .A2(new_n249), .A3(new_n263), .ZN(new_n414));
  OAI21_X1  g213(.A(new_n332), .B1(new_n413), .B2(new_n414), .ZN(new_n415));
  NAND2_X1  g214(.A1(new_n415), .A2(new_n330), .ZN(new_n416));
  NAND2_X1  g215(.A1(new_n416), .A2(new_n403), .ZN(new_n417));
  INV_X1    g216(.A(KEYINPUT76), .ZN(new_n418));
  INV_X1    g217(.A(new_n406), .ZN(new_n419));
  NAND3_X1  g218(.A1(new_n417), .A2(new_n418), .A3(new_n419), .ZN(new_n420));
  AOI22_X1  g219(.A1(new_n415), .A2(new_n330), .B1(new_n266), .B2(new_n402), .ZN(new_n421));
  OAI21_X1  g220(.A(KEYINPUT76), .B1(new_n421), .B2(new_n406), .ZN(new_n422));
  AOI21_X1  g221(.A(new_n411), .B1(new_n420), .B2(new_n422), .ZN(new_n423));
  INV_X1    g222(.A(G22gat), .ZN(new_n424));
  NOR2_X1   g223(.A1(new_n423), .A2(new_n424), .ZN(new_n425));
  AOI211_X1 g224(.A(G22gat), .B(new_n411), .C1(new_n420), .C2(new_n422), .ZN(new_n426));
  XNOR2_X1  g225(.A(G78gat), .B(G106gat), .ZN(new_n427));
  XNOR2_X1  g226(.A(KEYINPUT31), .B(G50gat), .ZN(new_n428));
  XNOR2_X1  g227(.A(new_n427), .B(new_n428), .ZN(new_n429));
  INV_X1    g228(.A(new_n429), .ZN(new_n430));
  NOR3_X1   g229(.A1(new_n425), .A2(new_n426), .A3(new_n430), .ZN(new_n431));
  AOI21_X1  g230(.A(new_n418), .B1(new_n417), .B2(new_n419), .ZN(new_n432));
  NOR3_X1   g231(.A1(new_n421), .A2(KEYINPUT76), .A3(new_n406), .ZN(new_n433));
  OAI22_X1  g232(.A1(new_n432), .A2(new_n433), .B1(new_n410), .B2(new_n407), .ZN(new_n434));
  NAND2_X1  g233(.A1(new_n434), .A2(G22gat), .ZN(new_n435));
  NAND2_X1  g234(.A1(new_n423), .A2(new_n424), .ZN(new_n436));
  AOI21_X1  g235(.A(new_n429), .B1(new_n435), .B2(new_n436), .ZN(new_n437));
  OAI21_X1  g236(.A(new_n401), .B1(new_n431), .B2(new_n437), .ZN(new_n438));
  NAND2_X1  g237(.A1(new_n438), .A2(KEYINPUT82), .ZN(new_n439));
  OAI21_X1  g238(.A(new_n430), .B1(new_n425), .B2(new_n426), .ZN(new_n440));
  NAND3_X1  g239(.A1(new_n435), .A2(new_n436), .A3(new_n429), .ZN(new_n441));
  NAND2_X1  g240(.A1(new_n440), .A2(new_n441), .ZN(new_n442));
  INV_X1    g241(.A(KEYINPUT82), .ZN(new_n443));
  NAND3_X1  g242(.A1(new_n442), .A2(new_n443), .A3(new_n401), .ZN(new_n444));
  AOI21_X1  g243(.A(new_n368), .B1(new_n439), .B2(new_n444), .ZN(new_n445));
  NAND2_X1  g244(.A1(new_n387), .A2(new_n393), .ZN(new_n446));
  NAND3_X1  g245(.A1(new_n399), .A2(new_n395), .A3(new_n386), .ZN(new_n447));
  NAND2_X1  g246(.A1(new_n446), .A2(new_n447), .ZN(new_n448));
  INV_X1    g247(.A(KEYINPUT36), .ZN(new_n449));
  NAND2_X1  g248(.A1(new_n448), .A2(new_n449), .ZN(new_n450));
  NAND3_X1  g249(.A1(new_n446), .A2(KEYINPUT36), .A3(new_n447), .ZN(new_n451));
  AOI21_X1  g250(.A(new_n442), .B1(new_n450), .B2(new_n451), .ZN(new_n452));
  OAI211_X1 g251(.A(new_n288), .B(new_n367), .C1(new_n445), .C2(new_n452), .ZN(new_n453));
  INV_X1    g252(.A(new_n288), .ZN(new_n454));
  INV_X1    g253(.A(KEYINPUT79), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n355), .A2(new_n455), .ZN(new_n456));
  NAND3_X1  g255(.A1(new_n344), .A2(new_n354), .A3(KEYINPUT79), .ZN(new_n457));
  NAND3_X1  g256(.A1(new_n456), .A2(new_n361), .A3(new_n457), .ZN(new_n458));
  AOI21_X1  g257(.A(new_n365), .B1(new_n458), .B2(new_n360), .ZN(new_n459));
  OAI21_X1  g258(.A(KEYINPUT81), .B1(new_n454), .B2(new_n459), .ZN(new_n460));
  INV_X1    g259(.A(new_n457), .ZN(new_n461));
  AOI21_X1  g260(.A(KEYINPUT79), .B1(new_n344), .B2(new_n354), .ZN(new_n462));
  NOR3_X1   g261(.A1(new_n461), .A2(new_n462), .A3(new_n359), .ZN(new_n463));
  INV_X1    g262(.A(new_n360), .ZN(new_n464));
  OAI21_X1  g263(.A(new_n366), .B1(new_n463), .B2(new_n464), .ZN(new_n465));
  INV_X1    g264(.A(KEYINPUT81), .ZN(new_n466));
  NAND3_X1  g265(.A1(new_n465), .A2(new_n466), .A3(new_n288), .ZN(new_n467));
  AOI21_X1  g266(.A(new_n448), .B1(new_n441), .B2(new_n440), .ZN(new_n468));
  NAND3_X1  g267(.A1(new_n460), .A2(new_n467), .A3(new_n468), .ZN(new_n469));
  INV_X1    g268(.A(KEYINPUT40), .ZN(new_n470));
  NAND3_X1  g269(.A1(new_n350), .A2(new_n343), .A3(new_n352), .ZN(new_n471));
  NAND2_X1  g270(.A1(new_n471), .A2(new_n345), .ZN(new_n472));
  NAND2_X1  g271(.A1(new_n472), .A2(KEYINPUT39), .ZN(new_n473));
  NAND2_X1  g272(.A1(new_n330), .A2(new_n342), .ZN(new_n474));
  NAND3_X1  g273(.A1(new_n327), .A2(new_n474), .A3(new_n329), .ZN(new_n475));
  XNOR2_X1  g274(.A(new_n475), .B(KEYINPUT77), .ZN(new_n476));
  NOR2_X1   g275(.A1(new_n473), .A2(new_n476), .ZN(new_n477));
  OAI21_X1  g276(.A(new_n359), .B1(new_n472), .B2(KEYINPUT39), .ZN(new_n478));
  OAI21_X1  g277(.A(new_n470), .B1(new_n477), .B2(new_n478), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n479), .A2(KEYINPUT78), .ZN(new_n480));
  INV_X1    g279(.A(KEYINPUT78), .ZN(new_n481));
  OAI211_X1 g280(.A(new_n481), .B(new_n470), .C1(new_n477), .C2(new_n478), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n480), .A2(new_n482), .ZN(new_n483));
  NOR3_X1   g282(.A1(new_n477), .A2(new_n470), .A3(new_n478), .ZN(new_n484));
  NOR2_X1   g283(.A1(new_n463), .A2(new_n484), .ZN(new_n485));
  NAND3_X1  g284(.A1(new_n483), .A2(new_n454), .A3(new_n485), .ZN(new_n486));
  OAI21_X1  g285(.A(KEYINPUT37), .B1(new_n276), .B2(new_n280), .ZN(new_n487));
  INV_X1    g286(.A(KEYINPUT38), .ZN(new_n488));
  INV_X1    g287(.A(KEYINPUT37), .ZN(new_n489));
  NAND3_X1  g288(.A1(new_n283), .A2(new_n489), .A3(new_n275), .ZN(new_n490));
  NAND4_X1  g289(.A1(new_n487), .A2(new_n488), .A3(new_n490), .A4(new_n205), .ZN(new_n491));
  INV_X1    g290(.A(KEYINPUT80), .ZN(new_n492));
  XNOR2_X1  g291(.A(new_n491), .B(new_n492), .ZN(new_n493));
  NAND3_X1  g292(.A1(new_n487), .A2(new_n205), .A3(new_n490), .ZN(new_n494));
  NAND2_X1  g293(.A1(new_n494), .A2(KEYINPUT38), .ZN(new_n495));
  NAND3_X1  g294(.A1(new_n459), .A2(new_n284), .A3(new_n495), .ZN(new_n496));
  OAI21_X1  g295(.A(new_n486), .B1(new_n493), .B2(new_n496), .ZN(new_n497));
  AOI22_X1  g296(.A1(new_n450), .A2(new_n451), .B1(new_n441), .B2(new_n440), .ZN(new_n498));
  AOI22_X1  g297(.A1(new_n368), .A2(new_n469), .B1(new_n497), .B2(new_n498), .ZN(new_n499));
  NAND2_X1  g298(.A1(new_n453), .A2(new_n499), .ZN(new_n500));
  AND2_X1   g299(.A1(G57gat), .A2(G64gat), .ZN(new_n501));
  NOR2_X1   g300(.A1(G57gat), .A2(G64gat), .ZN(new_n502));
  NOR2_X1   g301(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  INV_X1    g302(.A(KEYINPUT91), .ZN(new_n504));
  NAND2_X1  g303(.A1(G71gat), .A2(G78gat), .ZN(new_n505));
  OR2_X1    g304(.A1(G71gat), .A2(G78gat), .ZN(new_n506));
  AOI22_X1  g305(.A1(new_n503), .A2(new_n504), .B1(new_n505), .B2(new_n506), .ZN(new_n507));
  INV_X1    g306(.A(KEYINPUT90), .ZN(new_n508));
  INV_X1    g307(.A(KEYINPUT9), .ZN(new_n509));
  AND3_X1   g308(.A1(new_n505), .A2(new_n508), .A3(new_n509), .ZN(new_n510));
  AOI21_X1  g309(.A(new_n508), .B1(new_n505), .B2(new_n509), .ZN(new_n511));
  OAI21_X1  g310(.A(new_n503), .B1(new_n510), .B2(new_n511), .ZN(new_n512));
  NAND2_X1  g311(.A1(new_n507), .A2(new_n512), .ZN(new_n513));
  OR2_X1    g312(.A1(G57gat), .A2(G64gat), .ZN(new_n514));
  NAND2_X1  g313(.A1(G57gat), .A2(G64gat), .ZN(new_n515));
  NAND3_X1  g314(.A1(new_n514), .A2(new_n504), .A3(new_n515), .ZN(new_n516));
  NAND2_X1  g315(.A1(new_n506), .A2(new_n505), .ZN(new_n517));
  NAND2_X1  g316(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  NAND2_X1  g317(.A1(new_n505), .A2(new_n509), .ZN(new_n519));
  NAND2_X1  g318(.A1(new_n519), .A2(KEYINPUT90), .ZN(new_n520));
  NAND3_X1  g319(.A1(new_n505), .A2(new_n508), .A3(new_n509), .ZN(new_n521));
  NAND2_X1  g320(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  NAND3_X1  g321(.A1(new_n518), .A2(new_n522), .A3(new_n503), .ZN(new_n523));
  AND3_X1   g322(.A1(new_n513), .A2(new_n523), .A3(KEYINPUT93), .ZN(new_n524));
  INV_X1    g323(.A(new_n524), .ZN(new_n525));
  AOI21_X1  g324(.A(KEYINPUT93), .B1(new_n513), .B2(new_n523), .ZN(new_n526));
  INV_X1    g325(.A(new_n526), .ZN(new_n527));
  NAND3_X1  g326(.A1(new_n525), .A2(KEYINPUT21), .A3(new_n527), .ZN(new_n528));
  INV_X1    g327(.A(G1gat), .ZN(new_n529));
  NAND2_X1  g328(.A1(new_n529), .A2(KEYINPUT16), .ZN(new_n530));
  NAND2_X1  g329(.A1(new_n424), .A2(G15gat), .ZN(new_n531));
  INV_X1    g330(.A(G15gat), .ZN(new_n532));
  NAND2_X1  g331(.A1(new_n532), .A2(G22gat), .ZN(new_n533));
  INV_X1    g332(.A(KEYINPUT86), .ZN(new_n534));
  NAND3_X1  g333(.A1(new_n531), .A2(new_n533), .A3(new_n534), .ZN(new_n535));
  INV_X1    g334(.A(new_n535), .ZN(new_n536));
  AOI21_X1  g335(.A(new_n534), .B1(new_n531), .B2(new_n533), .ZN(new_n537));
  OAI21_X1  g336(.A(new_n530), .B1(new_n536), .B2(new_n537), .ZN(new_n538));
  NAND2_X1  g337(.A1(new_n531), .A2(new_n533), .ZN(new_n539));
  NAND2_X1  g338(.A1(new_n539), .A2(KEYINPUT86), .ZN(new_n540));
  NAND3_X1  g339(.A1(new_n540), .A2(new_n529), .A3(new_n535), .ZN(new_n541));
  INV_X1    g340(.A(G8gat), .ZN(new_n542));
  AND3_X1   g341(.A1(new_n538), .A2(new_n541), .A3(new_n542), .ZN(new_n543));
  AOI21_X1  g342(.A(new_n542), .B1(new_n538), .B2(new_n541), .ZN(new_n544));
  NOR2_X1   g343(.A1(new_n543), .A2(new_n544), .ZN(new_n545));
  NAND2_X1  g344(.A1(new_n528), .A2(new_n545), .ZN(new_n546));
  NAND2_X1  g345(.A1(new_n513), .A2(new_n523), .ZN(new_n547));
  NOR2_X1   g346(.A1(new_n547), .A2(KEYINPUT21), .ZN(new_n548));
  XOR2_X1   g347(.A(G127gat), .B(G155gat), .Z(new_n549));
  XNOR2_X1  g348(.A(new_n548), .B(new_n549), .ZN(new_n550));
  XNOR2_X1  g349(.A(new_n546), .B(new_n550), .ZN(new_n551));
  NAND2_X1  g350(.A1(G231gat), .A2(G233gat), .ZN(new_n552));
  XNOR2_X1  g351(.A(new_n552), .B(KEYINPUT92), .ZN(new_n553));
  XOR2_X1   g352(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n554));
  XNOR2_X1  g353(.A(new_n553), .B(new_n554), .ZN(new_n555));
  XNOR2_X1  g354(.A(G183gat), .B(G211gat), .ZN(new_n556));
  XNOR2_X1  g355(.A(new_n555), .B(new_n556), .ZN(new_n557));
  OR2_X1    g356(.A1(new_n551), .A2(new_n557), .ZN(new_n558));
  NAND2_X1  g357(.A1(new_n551), .A2(new_n557), .ZN(new_n559));
  NAND2_X1  g358(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  AND2_X1   g359(.A1(G232gat), .A2(G233gat), .ZN(new_n561));
  NOR2_X1   g360(.A1(new_n561), .A2(KEYINPUT41), .ZN(new_n562));
  XNOR2_X1  g361(.A(new_n562), .B(KEYINPUT94), .ZN(new_n563));
  XNOR2_X1  g362(.A(G134gat), .B(G162gat), .ZN(new_n564));
  XNOR2_X1  g363(.A(new_n563), .B(new_n564), .ZN(new_n565));
  INV_X1    g364(.A(new_n565), .ZN(new_n566));
  INV_X1    g365(.A(G50gat), .ZN(new_n567));
  NAND2_X1  g366(.A1(new_n567), .A2(G43gat), .ZN(new_n568));
  INV_X1    g367(.A(G43gat), .ZN(new_n569));
  NAND2_X1  g368(.A1(new_n569), .A2(G50gat), .ZN(new_n570));
  INV_X1    g369(.A(KEYINPUT84), .ZN(new_n571));
  AND3_X1   g370(.A1(new_n568), .A2(new_n570), .A3(new_n571), .ZN(new_n572));
  NAND3_X1  g371(.A1(new_n567), .A2(KEYINPUT84), .A3(G43gat), .ZN(new_n573));
  INV_X1    g372(.A(KEYINPUT15), .ZN(new_n574));
  NAND2_X1  g373(.A1(new_n573), .A2(new_n574), .ZN(new_n575));
  OAI21_X1  g374(.A(KEYINPUT85), .B1(new_n572), .B2(new_n575), .ZN(new_n576));
  NAND3_X1  g375(.A1(new_n568), .A2(new_n570), .A3(KEYINPUT15), .ZN(new_n577));
  XNOR2_X1  g376(.A(KEYINPUT14), .B(G29gat), .ZN(new_n578));
  INV_X1    g377(.A(G36gat), .ZN(new_n579));
  NAND2_X1  g378(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  INV_X1    g379(.A(G29gat), .ZN(new_n581));
  NAND3_X1  g380(.A1(new_n581), .A2(KEYINPUT14), .A3(G36gat), .ZN(new_n582));
  AOI22_X1  g381(.A1(new_n576), .A2(new_n577), .B1(new_n580), .B2(new_n582), .ZN(new_n583));
  INV_X1    g382(.A(new_n577), .ZN(new_n584));
  NAND2_X1  g383(.A1(new_n580), .A2(new_n582), .ZN(new_n585));
  NAND3_X1  g384(.A1(new_n568), .A2(new_n570), .A3(new_n571), .ZN(new_n586));
  INV_X1    g385(.A(KEYINPUT85), .ZN(new_n587));
  NAND4_X1  g386(.A1(new_n586), .A2(new_n587), .A3(new_n574), .A4(new_n573), .ZN(new_n588));
  AOI21_X1  g387(.A(new_n584), .B1(new_n585), .B2(new_n588), .ZN(new_n589));
  NOR2_X1   g388(.A1(new_n583), .A2(new_n589), .ZN(new_n590));
  NAND2_X1  g389(.A1(G99gat), .A2(G106gat), .ZN(new_n591));
  NAND2_X1  g390(.A1(new_n591), .A2(KEYINPUT8), .ZN(new_n592));
  NAND2_X1  g391(.A1(G85gat), .A2(G92gat), .ZN(new_n593));
  INV_X1    g392(.A(KEYINPUT7), .ZN(new_n594));
  NAND2_X1  g393(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  INV_X1    g394(.A(G85gat), .ZN(new_n596));
  INV_X1    g395(.A(G92gat), .ZN(new_n597));
  NAND2_X1  g396(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  NAND3_X1  g397(.A1(KEYINPUT7), .A2(G85gat), .A3(G92gat), .ZN(new_n599));
  NAND4_X1  g398(.A1(new_n592), .A2(new_n595), .A3(new_n598), .A4(new_n599), .ZN(new_n600));
  XNOR2_X1  g399(.A(G99gat), .B(G106gat), .ZN(new_n601));
  INV_X1    g400(.A(new_n601), .ZN(new_n602));
  NOR2_X1   g401(.A1(new_n600), .A2(new_n602), .ZN(new_n603));
  AND3_X1   g402(.A1(KEYINPUT7), .A2(G85gat), .A3(G92gat), .ZN(new_n604));
  AOI21_X1  g403(.A(KEYINPUT7), .B1(G85gat), .B2(G92gat), .ZN(new_n605));
  NOR2_X1   g404(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  AOI22_X1  g405(.A1(KEYINPUT8), .A2(new_n591), .B1(new_n596), .B2(new_n597), .ZN(new_n607));
  AOI21_X1  g406(.A(new_n601), .B1(new_n606), .B2(new_n607), .ZN(new_n608));
  NOR2_X1   g407(.A1(new_n603), .A2(new_n608), .ZN(new_n609));
  AOI22_X1  g408(.A1(new_n590), .A2(new_n609), .B1(KEYINPUT41), .B2(new_n561), .ZN(new_n610));
  OAI21_X1  g409(.A(KEYINPUT17), .B1(new_n583), .B2(new_n589), .ZN(new_n611));
  NAND2_X1  g410(.A1(new_n585), .A2(new_n588), .ZN(new_n612));
  NAND2_X1  g411(.A1(new_n612), .A2(new_n577), .ZN(new_n613));
  INV_X1    g412(.A(new_n575), .ZN(new_n614));
  AOI21_X1  g413(.A(new_n587), .B1(new_n614), .B2(new_n586), .ZN(new_n615));
  OAI21_X1  g414(.A(new_n585), .B1(new_n615), .B2(new_n584), .ZN(new_n616));
  INV_X1    g415(.A(KEYINPUT17), .ZN(new_n617));
  NAND3_X1  g416(.A1(new_n613), .A2(new_n616), .A3(new_n617), .ZN(new_n618));
  INV_X1    g417(.A(new_n609), .ZN(new_n619));
  NAND3_X1  g418(.A1(new_n611), .A2(new_n618), .A3(new_n619), .ZN(new_n620));
  XNOR2_X1  g419(.A(G190gat), .B(G218gat), .ZN(new_n621));
  XNOR2_X1  g420(.A(new_n621), .B(KEYINPUT95), .ZN(new_n622));
  INV_X1    g421(.A(new_n622), .ZN(new_n623));
  NAND3_X1  g422(.A1(new_n610), .A2(new_n620), .A3(new_n623), .ZN(new_n624));
  INV_X1    g423(.A(new_n624), .ZN(new_n625));
  AOI21_X1  g424(.A(new_n623), .B1(new_n610), .B2(new_n620), .ZN(new_n626));
  OAI21_X1  g425(.A(new_n566), .B1(new_n625), .B2(new_n626), .ZN(new_n627));
  INV_X1    g426(.A(new_n627), .ZN(new_n628));
  NOR3_X1   g427(.A1(new_n625), .A2(new_n566), .A3(new_n626), .ZN(new_n629));
  NOR2_X1   g428(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  NOR2_X1   g429(.A1(new_n560), .A2(new_n630), .ZN(new_n631));
  NAND2_X1  g430(.A1(G230gat), .A2(G233gat), .ZN(new_n632));
  INV_X1    g431(.A(KEYINPUT96), .ZN(new_n633));
  OAI21_X1  g432(.A(new_n633), .B1(new_n603), .B2(new_n608), .ZN(new_n634));
  NAND2_X1  g433(.A1(new_n600), .A2(new_n602), .ZN(new_n635));
  NAND3_X1  g434(.A1(new_n606), .A2(new_n601), .A3(new_n607), .ZN(new_n636));
  NAND3_X1  g435(.A1(new_n635), .A2(KEYINPUT96), .A3(new_n636), .ZN(new_n637));
  NAND3_X1  g436(.A1(new_n547), .A2(new_n634), .A3(new_n637), .ZN(new_n638));
  NAND4_X1  g437(.A1(new_n609), .A2(KEYINPUT96), .A3(new_n523), .A4(new_n513), .ZN(new_n639));
  AOI21_X1  g438(.A(KEYINPUT10), .B1(new_n638), .B2(new_n639), .ZN(new_n640));
  NAND3_X1  g439(.A1(new_n635), .A2(KEYINPUT10), .A3(new_n636), .ZN(new_n641));
  NOR3_X1   g440(.A1(new_n524), .A2(new_n526), .A3(new_n641), .ZN(new_n642));
  OAI21_X1  g441(.A(new_n632), .B1(new_n640), .B2(new_n642), .ZN(new_n643));
  INV_X1    g442(.A(new_n643), .ZN(new_n644));
  NAND2_X1  g443(.A1(new_n638), .A2(new_n639), .ZN(new_n645));
  NOR2_X1   g444(.A1(new_n645), .A2(new_n632), .ZN(new_n646));
  XNOR2_X1  g445(.A(G120gat), .B(G148gat), .ZN(new_n647));
  XNOR2_X1  g446(.A(G176gat), .B(G204gat), .ZN(new_n648));
  XOR2_X1   g447(.A(new_n647), .B(new_n648), .Z(new_n649));
  INV_X1    g448(.A(new_n649), .ZN(new_n650));
  NOR3_X1   g449(.A1(new_n644), .A2(new_n646), .A3(new_n650), .ZN(new_n651));
  INV_X1    g450(.A(new_n651), .ZN(new_n652));
  OAI21_X1  g451(.A(new_n650), .B1(new_n644), .B2(new_n646), .ZN(new_n653));
  NAND2_X1  g452(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  INV_X1    g453(.A(new_n654), .ZN(new_n655));
  NAND2_X1  g454(.A1(new_n631), .A2(new_n655), .ZN(new_n656));
  XNOR2_X1  g455(.A(G113gat), .B(G141gat), .ZN(new_n657));
  XNOR2_X1  g456(.A(G169gat), .B(G197gat), .ZN(new_n658));
  XNOR2_X1  g457(.A(new_n657), .B(new_n658), .ZN(new_n659));
  XOR2_X1   g458(.A(KEYINPUT83), .B(KEYINPUT11), .Z(new_n660));
  XNOR2_X1  g459(.A(new_n659), .B(new_n660), .ZN(new_n661));
  XNOR2_X1  g460(.A(new_n661), .B(KEYINPUT12), .ZN(new_n662));
  INV_X1    g461(.A(new_n662), .ZN(new_n663));
  NAND3_X1  g462(.A1(new_n545), .A2(new_n611), .A3(new_n618), .ZN(new_n664));
  OAI21_X1  g463(.A(new_n590), .B1(new_n544), .B2(new_n543), .ZN(new_n665));
  NAND2_X1  g464(.A1(G229gat), .A2(G233gat), .ZN(new_n666));
  NAND4_X1  g465(.A1(new_n664), .A2(KEYINPUT18), .A3(new_n665), .A4(new_n666), .ZN(new_n667));
  INV_X1    g466(.A(KEYINPUT88), .ZN(new_n668));
  XNOR2_X1  g467(.A(new_n667), .B(new_n668), .ZN(new_n669));
  NAND2_X1  g468(.A1(new_n613), .A2(new_n616), .ZN(new_n670));
  AOI21_X1  g469(.A(KEYINPUT89), .B1(new_n545), .B2(new_n670), .ZN(new_n671));
  NAND2_X1  g470(.A1(new_n671), .A2(new_n665), .ZN(new_n672));
  OAI211_X1 g471(.A(new_n590), .B(KEYINPUT89), .C1(new_n544), .C2(new_n543), .ZN(new_n673));
  XOR2_X1   g472(.A(new_n666), .B(KEYINPUT13), .Z(new_n674));
  NAND3_X1  g473(.A1(new_n672), .A2(new_n673), .A3(new_n674), .ZN(new_n675));
  NAND3_X1  g474(.A1(new_n664), .A2(new_n666), .A3(new_n665), .ZN(new_n676));
  XNOR2_X1  g475(.A(KEYINPUT87), .B(KEYINPUT18), .ZN(new_n677));
  NAND2_X1  g476(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  NAND2_X1  g477(.A1(new_n675), .A2(new_n678), .ZN(new_n679));
  OAI21_X1  g478(.A(new_n663), .B1(new_n669), .B2(new_n679), .ZN(new_n680));
  XNOR2_X1  g479(.A(new_n667), .B(KEYINPUT88), .ZN(new_n681));
  NAND4_X1  g480(.A1(new_n681), .A2(new_n675), .A3(new_n678), .A4(new_n662), .ZN(new_n682));
  NAND2_X1  g481(.A1(new_n680), .A2(new_n682), .ZN(new_n683));
  INV_X1    g482(.A(new_n683), .ZN(new_n684));
  NOR2_X1   g483(.A1(new_n656), .A2(new_n684), .ZN(new_n685));
  AND2_X1   g484(.A1(new_n500), .A2(new_n685), .ZN(new_n686));
  OR2_X1    g485(.A1(new_n367), .A2(KEYINPUT97), .ZN(new_n687));
  NAND2_X1  g486(.A1(new_n367), .A2(KEYINPUT97), .ZN(new_n688));
  NAND2_X1  g487(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  INV_X1    g488(.A(new_n689), .ZN(new_n690));
  NAND2_X1  g489(.A1(new_n686), .A2(new_n690), .ZN(new_n691));
  XNOR2_X1  g490(.A(new_n691), .B(G1gat), .ZN(G1324gat));
  INV_X1    g491(.A(new_n686), .ZN(new_n693));
  XNOR2_X1  g492(.A(KEYINPUT16), .B(G8gat), .ZN(new_n694));
  NOR3_X1   g493(.A1(new_n693), .A2(new_n288), .A3(new_n694), .ZN(new_n695));
  AOI21_X1  g494(.A(new_n542), .B1(new_n686), .B2(new_n454), .ZN(new_n696));
  OAI21_X1  g495(.A(KEYINPUT42), .B1(new_n695), .B2(new_n696), .ZN(new_n697));
  OAI21_X1  g496(.A(new_n697), .B1(KEYINPUT42), .B2(new_n695), .ZN(G1325gat));
  NAND2_X1  g497(.A1(new_n450), .A2(new_n451), .ZN(new_n699));
  OAI21_X1  g498(.A(G15gat), .B1(new_n693), .B2(new_n699), .ZN(new_n700));
  NAND3_X1  g499(.A1(new_n686), .A2(new_n532), .A3(new_n401), .ZN(new_n701));
  NAND2_X1  g500(.A1(new_n700), .A2(new_n701), .ZN(G1326gat));
  INV_X1    g501(.A(new_n442), .ZN(new_n703));
  NAND2_X1  g502(.A1(new_n686), .A2(new_n703), .ZN(new_n704));
  XNOR2_X1  g503(.A(KEYINPUT43), .B(G22gat), .ZN(new_n705));
  XNOR2_X1  g504(.A(new_n704), .B(new_n705), .ZN(G1327gat));
  NAND2_X1  g505(.A1(new_n367), .A2(new_n288), .ZN(new_n707));
  AND3_X1   g506(.A1(new_n442), .A2(new_n443), .A3(new_n401), .ZN(new_n708));
  AOI21_X1  g507(.A(new_n443), .B1(new_n442), .B2(new_n401), .ZN(new_n709));
  OAI21_X1  g508(.A(KEYINPUT35), .B1(new_n708), .B2(new_n709), .ZN(new_n710));
  INV_X1    g509(.A(new_n452), .ZN(new_n711));
  AOI21_X1  g510(.A(new_n707), .B1(new_n710), .B2(new_n711), .ZN(new_n712));
  NAND2_X1  g511(.A1(new_n469), .A2(new_n368), .ZN(new_n713));
  NAND2_X1  g512(.A1(new_n497), .A2(new_n498), .ZN(new_n714));
  NAND2_X1  g513(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  OAI21_X1  g514(.A(new_n630), .B1(new_n712), .B2(new_n715), .ZN(new_n716));
  INV_X1    g515(.A(new_n560), .ZN(new_n717));
  NOR3_X1   g516(.A1(new_n684), .A2(new_n717), .A3(new_n654), .ZN(new_n718));
  INV_X1    g517(.A(new_n718), .ZN(new_n719));
  NOR2_X1   g518(.A1(new_n716), .A2(new_n719), .ZN(new_n720));
  NAND3_X1  g519(.A1(new_n720), .A2(new_n581), .A3(new_n690), .ZN(new_n721));
  XNOR2_X1  g520(.A(new_n721), .B(KEYINPUT45), .ZN(new_n722));
  INV_X1    g521(.A(KEYINPUT98), .ZN(new_n723));
  OAI21_X1  g522(.A(new_n723), .B1(new_n712), .B2(new_n715), .ZN(new_n724));
  NAND2_X1  g523(.A1(new_n439), .A2(new_n444), .ZN(new_n725));
  AOI21_X1  g524(.A(new_n452), .B1(new_n725), .B2(KEYINPUT35), .ZN(new_n726));
  OAI211_X1 g525(.A(new_n499), .B(KEYINPUT98), .C1(new_n726), .C2(new_n707), .ZN(new_n727));
  XNOR2_X1  g526(.A(new_n630), .B(KEYINPUT99), .ZN(new_n728));
  INV_X1    g527(.A(new_n728), .ZN(new_n729));
  NOR2_X1   g528(.A1(new_n729), .A2(KEYINPUT44), .ZN(new_n730));
  NAND3_X1  g529(.A1(new_n724), .A2(new_n727), .A3(new_n730), .ZN(new_n731));
  NAND2_X1  g530(.A1(new_n716), .A2(KEYINPUT44), .ZN(new_n732));
  AOI21_X1  g531(.A(new_n719), .B1(new_n731), .B2(new_n732), .ZN(new_n733));
  INV_X1    g532(.A(new_n733), .ZN(new_n734));
  OAI21_X1  g533(.A(G29gat), .B1(new_n734), .B2(new_n689), .ZN(new_n735));
  NAND2_X1  g534(.A1(new_n722), .A2(new_n735), .ZN(G1328gat));
  NAND3_X1  g535(.A1(new_n720), .A2(new_n579), .A3(new_n454), .ZN(new_n737));
  XOR2_X1   g536(.A(new_n737), .B(KEYINPUT46), .Z(new_n738));
  OAI21_X1  g537(.A(G36gat), .B1(new_n734), .B2(new_n288), .ZN(new_n739));
  NAND2_X1  g538(.A1(new_n738), .A2(new_n739), .ZN(G1329gat));
  INV_X1    g539(.A(new_n699), .ZN(new_n741));
  NAND3_X1  g540(.A1(new_n733), .A2(G43gat), .A3(new_n741), .ZN(new_n742));
  INV_X1    g541(.A(new_n720), .ZN(new_n743));
  OAI21_X1  g542(.A(new_n569), .B1(new_n743), .B2(new_n448), .ZN(new_n744));
  INV_X1    g543(.A(KEYINPUT47), .ZN(new_n745));
  OAI211_X1 g544(.A(new_n742), .B(new_n744), .C1(KEYINPUT100), .C2(new_n745), .ZN(new_n746));
  NAND2_X1  g545(.A1(new_n745), .A2(KEYINPUT100), .ZN(new_n747));
  XNOR2_X1  g546(.A(new_n746), .B(new_n747), .ZN(G1330gat));
  INV_X1    g547(.A(KEYINPUT48), .ZN(new_n749));
  NAND3_X1  g548(.A1(new_n720), .A2(new_n567), .A3(new_n703), .ZN(new_n750));
  AOI21_X1  g549(.A(new_n567), .B1(new_n733), .B2(new_n703), .ZN(new_n751));
  INV_X1    g550(.A(KEYINPUT101), .ZN(new_n752));
  OAI21_X1  g551(.A(new_n750), .B1(new_n751), .B2(new_n752), .ZN(new_n753));
  AOI211_X1 g552(.A(new_n442), .B(new_n719), .C1(new_n731), .C2(new_n732), .ZN(new_n754));
  NOR3_X1   g553(.A1(new_n754), .A2(KEYINPUT101), .A3(new_n567), .ZN(new_n755));
  OAI21_X1  g554(.A(new_n749), .B1(new_n753), .B2(new_n755), .ZN(new_n756));
  INV_X1    g555(.A(KEYINPUT102), .ZN(new_n757));
  AND2_X1   g556(.A1(new_n754), .A2(new_n757), .ZN(new_n758));
  OAI21_X1  g557(.A(G50gat), .B1(new_n754), .B2(new_n757), .ZN(new_n759));
  OAI211_X1 g558(.A(KEYINPUT48), .B(new_n750), .C1(new_n758), .C2(new_n759), .ZN(new_n760));
  NAND2_X1  g559(.A1(new_n756), .A2(new_n760), .ZN(G1331gat));
  AND2_X1   g560(.A1(new_n724), .A2(new_n727), .ZN(new_n762));
  NOR4_X1   g561(.A1(new_n683), .A2(new_n560), .A3(new_n655), .A4(new_n630), .ZN(new_n763));
  AND2_X1   g562(.A1(new_n762), .A2(new_n763), .ZN(new_n764));
  NOR2_X1   g563(.A1(new_n690), .A2(KEYINPUT103), .ZN(new_n765));
  AND3_X1   g564(.A1(new_n687), .A2(KEYINPUT103), .A3(new_n688), .ZN(new_n766));
  NOR2_X1   g565(.A1(new_n765), .A2(new_n766), .ZN(new_n767));
  NAND2_X1  g566(.A1(new_n764), .A2(new_n767), .ZN(new_n768));
  XNOR2_X1  g567(.A(new_n768), .B(G57gat), .ZN(G1332gat));
  AOI21_X1  g568(.A(new_n288), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n770));
  XNOR2_X1  g569(.A(new_n770), .B(KEYINPUT104), .ZN(new_n771));
  NAND2_X1  g570(.A1(new_n764), .A2(new_n771), .ZN(new_n772));
  NOR2_X1   g571(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n773));
  XOR2_X1   g572(.A(new_n772), .B(new_n773), .Z(G1333gat));
  NOR2_X1   g573(.A1(new_n448), .A2(G71gat), .ZN(new_n775));
  NAND2_X1  g574(.A1(new_n764), .A2(new_n775), .ZN(new_n776));
  NAND2_X1  g575(.A1(new_n762), .A2(new_n763), .ZN(new_n777));
  OAI21_X1  g576(.A(G71gat), .B1(new_n777), .B2(new_n699), .ZN(new_n778));
  AND2_X1   g577(.A1(new_n776), .A2(new_n778), .ZN(new_n779));
  XNOR2_X1  g578(.A(new_n779), .B(KEYINPUT50), .ZN(G1334gat));
  NOR2_X1   g579(.A1(new_n777), .A2(new_n442), .ZN(new_n781));
  XOR2_X1   g580(.A(KEYINPUT105), .B(G78gat), .Z(new_n782));
  XNOR2_X1  g581(.A(new_n781), .B(new_n782), .ZN(G1335gat));
  NOR2_X1   g582(.A1(new_n717), .A2(new_n683), .ZN(new_n784));
  NAND2_X1  g583(.A1(new_n784), .A2(new_n654), .ZN(new_n785));
  AOI21_X1  g584(.A(new_n785), .B1(new_n731), .B2(new_n732), .ZN(new_n786));
  INV_X1    g585(.A(new_n786), .ZN(new_n787));
  OAI21_X1  g586(.A(G85gat), .B1(new_n787), .B2(new_n689), .ZN(new_n788));
  INV_X1    g587(.A(new_n630), .ZN(new_n789));
  AOI21_X1  g588(.A(new_n789), .B1(new_n453), .B2(new_n499), .ZN(new_n790));
  NAND4_X1  g589(.A1(new_n790), .A2(KEYINPUT106), .A3(KEYINPUT51), .A4(new_n784), .ZN(new_n791));
  INV_X1    g590(.A(KEYINPUT106), .ZN(new_n792));
  OAI211_X1 g591(.A(new_n630), .B(new_n784), .C1(new_n712), .C2(new_n715), .ZN(new_n793));
  INV_X1    g592(.A(KEYINPUT51), .ZN(new_n794));
  OAI21_X1  g593(.A(new_n792), .B1(new_n793), .B2(new_n794), .ZN(new_n795));
  NAND2_X1  g594(.A1(new_n793), .A2(new_n794), .ZN(new_n796));
  NAND3_X1  g595(.A1(new_n791), .A2(new_n795), .A3(new_n796), .ZN(new_n797));
  INV_X1    g596(.A(new_n797), .ZN(new_n798));
  NAND3_X1  g597(.A1(new_n690), .A2(new_n596), .A3(new_n654), .ZN(new_n799));
  XNOR2_X1  g598(.A(new_n799), .B(KEYINPUT107), .ZN(new_n800));
  OAI21_X1  g599(.A(new_n788), .B1(new_n798), .B2(new_n800), .ZN(G1336gat));
  AOI21_X1  g600(.A(new_n597), .B1(new_n786), .B2(new_n454), .ZN(new_n802));
  NOR2_X1   g601(.A1(new_n802), .A2(KEYINPUT52), .ZN(new_n803));
  NOR3_X1   g602(.A1(new_n655), .A2(G92gat), .A3(new_n288), .ZN(new_n804));
  INV_X1    g603(.A(new_n804), .ZN(new_n805));
  OAI21_X1  g604(.A(new_n803), .B1(new_n798), .B2(new_n805), .ZN(new_n806));
  NAND2_X1  g605(.A1(new_n793), .A2(KEYINPUT108), .ZN(new_n807));
  NAND2_X1  g606(.A1(new_n807), .A2(new_n794), .ZN(new_n808));
  NAND3_X1  g607(.A1(new_n793), .A2(KEYINPUT108), .A3(KEYINPUT51), .ZN(new_n809));
  AND3_X1   g608(.A1(new_n808), .A2(new_n809), .A3(new_n804), .ZN(new_n810));
  OAI21_X1  g609(.A(KEYINPUT52), .B1(new_n802), .B2(new_n810), .ZN(new_n811));
  NAND2_X1  g610(.A1(new_n806), .A2(new_n811), .ZN(G1337gat));
  OAI21_X1  g611(.A(G99gat), .B1(new_n787), .B2(new_n699), .ZN(new_n813));
  OR3_X1    g612(.A1(new_n655), .A2(new_n448), .A3(G99gat), .ZN(new_n814));
  OAI21_X1  g613(.A(new_n813), .B1(new_n798), .B2(new_n814), .ZN(G1338gat));
  INV_X1    g614(.A(G106gat), .ZN(new_n816));
  AOI21_X1  g615(.A(new_n816), .B1(new_n786), .B2(new_n703), .ZN(new_n817));
  NOR2_X1   g616(.A1(new_n817), .A2(KEYINPUT53), .ZN(new_n818));
  INV_X1    g617(.A(KEYINPUT110), .ZN(new_n819));
  NOR3_X1   g618(.A1(new_n442), .A2(G106gat), .A3(new_n655), .ZN(new_n820));
  AOI21_X1  g619(.A(new_n819), .B1(new_n797), .B2(new_n820), .ZN(new_n821));
  AND3_X1   g620(.A1(new_n797), .A2(new_n819), .A3(new_n820), .ZN(new_n822));
  OAI21_X1  g621(.A(new_n818), .B1(new_n821), .B2(new_n822), .ZN(new_n823));
  AND3_X1   g622(.A1(new_n808), .A2(new_n809), .A3(new_n820), .ZN(new_n824));
  OAI211_X1 g623(.A(KEYINPUT109), .B(KEYINPUT53), .C1(new_n817), .C2(new_n824), .ZN(new_n825));
  INV_X1    g624(.A(new_n825), .ZN(new_n826));
  NAND3_X1  g625(.A1(new_n808), .A2(new_n809), .A3(new_n820), .ZN(new_n827));
  AOI211_X1 g626(.A(new_n442), .B(new_n785), .C1(new_n731), .C2(new_n732), .ZN(new_n828));
  OAI21_X1  g627(.A(new_n827), .B1(new_n828), .B2(new_n816), .ZN(new_n829));
  AOI21_X1  g628(.A(KEYINPUT109), .B1(new_n829), .B2(KEYINPUT53), .ZN(new_n830));
  OAI21_X1  g629(.A(new_n823), .B1(new_n826), .B2(new_n830), .ZN(G1339gat));
  NAND3_X1  g630(.A1(new_n631), .A2(new_n684), .A3(new_n655), .ZN(new_n832));
  INV_X1    g631(.A(new_n832), .ZN(new_n833));
  INV_X1    g632(.A(KEYINPUT10), .ZN(new_n834));
  NAND2_X1  g633(.A1(new_n645), .A2(new_n834), .ZN(new_n835));
  INV_X1    g634(.A(new_n632), .ZN(new_n836));
  NAND4_X1  g635(.A1(new_n525), .A2(new_n527), .A3(KEYINPUT10), .A4(new_n609), .ZN(new_n837));
  NAND3_X1  g636(.A1(new_n835), .A2(new_n836), .A3(new_n837), .ZN(new_n838));
  NAND3_X1  g637(.A1(new_n838), .A2(KEYINPUT54), .A3(new_n643), .ZN(new_n839));
  NAND2_X1  g638(.A1(new_n839), .A2(KEYINPUT111), .ZN(new_n840));
  INV_X1    g639(.A(KEYINPUT111), .ZN(new_n841));
  NAND4_X1  g640(.A1(new_n838), .A2(new_n643), .A3(new_n841), .A4(KEYINPUT54), .ZN(new_n842));
  NAND2_X1  g641(.A1(new_n840), .A2(new_n842), .ZN(new_n843));
  INV_X1    g642(.A(KEYINPUT54), .ZN(new_n844));
  AOI21_X1  g643(.A(new_n649), .B1(new_n644), .B2(new_n844), .ZN(new_n845));
  AOI21_X1  g644(.A(KEYINPUT55), .B1(new_n843), .B2(new_n845), .ZN(new_n846));
  OAI211_X1 g645(.A(KEYINPUT55), .B(new_n650), .C1(new_n643), .C2(KEYINPUT54), .ZN(new_n847));
  INV_X1    g646(.A(new_n847), .ZN(new_n848));
  NAND2_X1  g647(.A1(new_n835), .A2(new_n837), .ZN(new_n849));
  AOI21_X1  g648(.A(new_n844), .B1(new_n849), .B2(new_n632), .ZN(new_n850));
  AOI21_X1  g649(.A(new_n841), .B1(new_n850), .B2(new_n838), .ZN(new_n851));
  INV_X1    g650(.A(new_n842), .ZN(new_n852));
  OAI21_X1  g651(.A(new_n848), .B1(new_n851), .B2(new_n852), .ZN(new_n853));
  INV_X1    g652(.A(KEYINPUT112), .ZN(new_n854));
  NAND3_X1  g653(.A1(new_n853), .A2(new_n854), .A3(new_n652), .ZN(new_n855));
  AOI21_X1  g654(.A(new_n847), .B1(new_n840), .B2(new_n842), .ZN(new_n856));
  OAI21_X1  g655(.A(KEYINPUT112), .B1(new_n856), .B2(new_n651), .ZN(new_n857));
  AOI21_X1  g656(.A(new_n846), .B1(new_n855), .B2(new_n857), .ZN(new_n858));
  AOI21_X1  g657(.A(new_n674), .B1(new_n672), .B2(new_n673), .ZN(new_n859));
  INV_X1    g658(.A(KEYINPUT113), .ZN(new_n860));
  AND2_X1   g659(.A1(new_n664), .A2(new_n665), .ZN(new_n861));
  OAI22_X1  g660(.A1(new_n859), .A2(new_n860), .B1(new_n666), .B2(new_n861), .ZN(new_n862));
  AND2_X1   g661(.A1(new_n859), .A2(new_n860), .ZN(new_n863));
  OAI21_X1  g662(.A(new_n661), .B1(new_n862), .B2(new_n863), .ZN(new_n864));
  AND2_X1   g663(.A1(new_n864), .A2(new_n682), .ZN(new_n865));
  NAND3_X1  g664(.A1(new_n858), .A2(new_n728), .A3(new_n865), .ZN(new_n866));
  NAND3_X1  g665(.A1(new_n864), .A2(new_n682), .A3(new_n654), .ZN(new_n867));
  INV_X1    g666(.A(new_n867), .ZN(new_n868));
  AOI21_X1  g667(.A(new_n868), .B1(new_n858), .B2(new_n683), .ZN(new_n869));
  OAI21_X1  g668(.A(new_n866), .B1(new_n869), .B2(new_n728), .ZN(new_n870));
  AOI21_X1  g669(.A(new_n833), .B1(new_n870), .B2(new_n560), .ZN(new_n871));
  NOR2_X1   g670(.A1(new_n871), .A2(new_n703), .ZN(new_n872));
  NAND4_X1  g671(.A1(new_n872), .A2(new_n401), .A3(new_n288), .A4(new_n690), .ZN(new_n873));
  OAI21_X1  g672(.A(G113gat), .B1(new_n873), .B2(new_n684), .ZN(new_n874));
  NOR3_X1   g673(.A1(new_n871), .A2(new_n766), .A3(new_n765), .ZN(new_n875));
  AND2_X1   g674(.A1(new_n875), .A2(new_n725), .ZN(new_n876));
  NAND2_X1  g675(.A1(new_n876), .A2(new_n288), .ZN(new_n877));
  NAND2_X1  g676(.A1(new_n683), .A2(new_n335), .ZN(new_n878));
  OAI21_X1  g677(.A(new_n874), .B1(new_n877), .B2(new_n878), .ZN(G1340gat));
  NOR3_X1   g678(.A1(new_n873), .A2(new_n292), .A3(new_n655), .ZN(new_n880));
  NAND3_X1  g679(.A1(new_n876), .A2(new_n288), .A3(new_n654), .ZN(new_n881));
  AOI21_X1  g680(.A(new_n880), .B1(new_n881), .B2(new_n292), .ZN(G1341gat));
  NOR3_X1   g681(.A1(new_n873), .A2(new_n340), .A3(new_n560), .ZN(new_n883));
  NOR2_X1   g682(.A1(new_n877), .A2(new_n560), .ZN(new_n884));
  AOI21_X1  g683(.A(G127gat), .B1(new_n884), .B2(KEYINPUT114), .ZN(new_n885));
  INV_X1    g684(.A(KEYINPUT114), .ZN(new_n886));
  OAI21_X1  g685(.A(new_n886), .B1(new_n877), .B2(new_n560), .ZN(new_n887));
  AOI21_X1  g686(.A(new_n883), .B1(new_n885), .B2(new_n887), .ZN(G1342gat));
  INV_X1    g687(.A(KEYINPUT56), .ZN(new_n889));
  INV_X1    g688(.A(KEYINPUT116), .ZN(new_n890));
  NAND2_X1  g689(.A1(new_n288), .A2(new_n630), .ZN(new_n891));
  XNOR2_X1  g690(.A(new_n891), .B(KEYINPUT115), .ZN(new_n892));
  NOR2_X1   g691(.A1(new_n892), .A2(new_n319), .ZN(new_n893));
  NAND3_X1  g692(.A1(new_n876), .A2(new_n890), .A3(new_n893), .ZN(new_n894));
  INV_X1    g693(.A(new_n894), .ZN(new_n895));
  AOI21_X1  g694(.A(new_n890), .B1(new_n876), .B2(new_n893), .ZN(new_n896));
  OAI21_X1  g695(.A(new_n889), .B1(new_n895), .B2(new_n896), .ZN(new_n897));
  INV_X1    g696(.A(new_n896), .ZN(new_n898));
  NAND3_X1  g697(.A1(new_n898), .A2(KEYINPUT56), .A3(new_n894), .ZN(new_n899));
  OAI21_X1  g698(.A(G134gat), .B1(new_n873), .B2(new_n789), .ZN(new_n900));
  NAND3_X1  g699(.A1(new_n897), .A2(new_n899), .A3(new_n900), .ZN(G1343gat));
  NAND2_X1  g700(.A1(new_n690), .A2(new_n288), .ZN(new_n902));
  NOR2_X1   g701(.A1(new_n902), .A2(new_n741), .ZN(new_n903));
  INV_X1    g702(.A(new_n903), .ZN(new_n904));
  INV_X1    g703(.A(KEYINPUT57), .ZN(new_n905));
  NOR2_X1   g704(.A1(new_n442), .A2(new_n905), .ZN(new_n906));
  INV_X1    g705(.A(new_n906), .ZN(new_n907));
  NAND2_X1  g706(.A1(new_n843), .A2(new_n845), .ZN(new_n908));
  INV_X1    g707(.A(KEYINPUT55), .ZN(new_n909));
  NAND2_X1  g708(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  NOR2_X1   g709(.A1(new_n856), .A2(new_n651), .ZN(new_n911));
  NAND3_X1  g710(.A1(new_n910), .A2(new_n683), .A3(new_n911), .ZN(new_n912));
  AOI21_X1  g711(.A(new_n630), .B1(new_n912), .B2(new_n867), .ZN(new_n913));
  INV_X1    g712(.A(KEYINPUT118), .ZN(new_n914));
  OAI21_X1  g713(.A(new_n866), .B1(new_n913), .B2(new_n914), .ZN(new_n915));
  AOI211_X1 g714(.A(KEYINPUT118), .B(new_n630), .C1(new_n912), .C2(new_n867), .ZN(new_n916));
  OAI21_X1  g715(.A(new_n560), .B1(new_n915), .B2(new_n916), .ZN(new_n917));
  AOI21_X1  g716(.A(new_n907), .B1(new_n917), .B2(new_n832), .ZN(new_n918));
  OAI21_X1  g717(.A(new_n905), .B1(new_n871), .B2(new_n442), .ZN(new_n919));
  AOI21_X1  g718(.A(new_n918), .B1(new_n919), .B2(KEYINPUT117), .ZN(new_n920));
  INV_X1    g719(.A(KEYINPUT117), .ZN(new_n921));
  OAI211_X1 g720(.A(new_n921), .B(new_n905), .C1(new_n871), .C2(new_n442), .ZN(new_n922));
  AOI21_X1  g721(.A(new_n904), .B1(new_n920), .B2(new_n922), .ZN(new_n923));
  AOI21_X1  g722(.A(new_n308), .B1(new_n923), .B2(new_n683), .ZN(new_n924));
  NOR2_X1   g723(.A1(new_n684), .A2(G141gat), .ZN(new_n925));
  NAND4_X1  g724(.A1(new_n875), .A2(new_n452), .A3(new_n288), .A4(new_n925), .ZN(new_n926));
  NAND2_X1  g725(.A1(new_n926), .A2(KEYINPUT119), .ZN(new_n927));
  OAI21_X1  g726(.A(KEYINPUT58), .B1(new_n924), .B2(new_n927), .ZN(new_n928));
  NAND2_X1  g727(.A1(new_n919), .A2(KEYINPUT117), .ZN(new_n929));
  INV_X1    g728(.A(new_n918), .ZN(new_n930));
  NAND3_X1  g729(.A1(new_n929), .A2(new_n922), .A3(new_n930), .ZN(new_n931));
  NAND3_X1  g730(.A1(new_n931), .A2(new_n683), .A3(new_n903), .ZN(new_n932));
  NAND2_X1  g731(.A1(new_n932), .A2(G141gat), .ZN(new_n933));
  INV_X1    g732(.A(KEYINPUT58), .ZN(new_n934));
  INV_X1    g733(.A(new_n927), .ZN(new_n935));
  NAND3_X1  g734(.A1(new_n933), .A2(new_n934), .A3(new_n935), .ZN(new_n936));
  NAND2_X1  g735(.A1(new_n928), .A2(new_n936), .ZN(G1344gat));
  NAND2_X1  g736(.A1(new_n875), .A2(new_n452), .ZN(new_n938));
  NOR2_X1   g737(.A1(new_n938), .A2(new_n454), .ZN(new_n939));
  NAND3_X1  g738(.A1(new_n939), .A2(new_n309), .A3(new_n654), .ZN(new_n940));
  AOI211_X1 g739(.A(KEYINPUT59), .B(new_n309), .C1(new_n923), .C2(new_n654), .ZN(new_n941));
  INV_X1    g740(.A(KEYINPUT59), .ZN(new_n942));
  AND3_X1   g741(.A1(new_n858), .A2(new_n630), .A3(new_n865), .ZN(new_n943));
  OAI21_X1  g742(.A(new_n560), .B1(new_n943), .B2(new_n913), .ZN(new_n944));
  XNOR2_X1  g743(.A(new_n832), .B(KEYINPUT120), .ZN(new_n945));
  AOI21_X1  g744(.A(new_n442), .B1(new_n944), .B2(new_n945), .ZN(new_n946));
  OAI22_X1  g745(.A1(new_n946), .A2(KEYINPUT57), .B1(new_n871), .B2(new_n907), .ZN(new_n947));
  NAND3_X1  g746(.A1(new_n947), .A2(new_n654), .A3(new_n903), .ZN(new_n948));
  AOI21_X1  g747(.A(new_n942), .B1(new_n948), .B2(G148gat), .ZN(new_n949));
  OAI21_X1  g748(.A(new_n940), .B1(new_n941), .B2(new_n949), .ZN(G1345gat));
  AOI21_X1  g749(.A(G155gat), .B1(new_n939), .B2(new_n717), .ZN(new_n951));
  NOR2_X1   g750(.A1(new_n560), .A2(new_n298), .ZN(new_n952));
  XNOR2_X1  g751(.A(new_n952), .B(KEYINPUT121), .ZN(new_n953));
  AOI21_X1  g752(.A(new_n951), .B1(new_n923), .B2(new_n953), .ZN(G1346gat));
  AOI21_X1  g753(.A(new_n299), .B1(new_n923), .B2(new_n728), .ZN(new_n955));
  NOR3_X1   g754(.A1(new_n938), .A2(G162gat), .A3(new_n892), .ZN(new_n956));
  OR2_X1    g755(.A1(new_n955), .A2(new_n956), .ZN(G1347gat));
  OAI21_X1  g756(.A(KEYINPUT122), .B1(new_n871), .B2(new_n690), .ZN(new_n958));
  AND2_X1   g757(.A1(new_n958), .A2(new_n454), .ZN(new_n959));
  INV_X1    g758(.A(KEYINPUT123), .ZN(new_n960));
  INV_X1    g759(.A(KEYINPUT122), .ZN(new_n961));
  AND2_X1   g760(.A1(new_n870), .A2(new_n560), .ZN(new_n962));
  OAI211_X1 g761(.A(new_n961), .B(new_n689), .C1(new_n962), .C2(new_n833), .ZN(new_n963));
  NAND4_X1  g762(.A1(new_n959), .A2(new_n960), .A3(new_n725), .A4(new_n963), .ZN(new_n964));
  NAND4_X1  g763(.A1(new_n963), .A2(new_n958), .A3(new_n725), .A4(new_n454), .ZN(new_n965));
  NAND2_X1  g764(.A1(new_n965), .A2(KEYINPUT123), .ZN(new_n966));
  NOR2_X1   g765(.A1(new_n684), .A2(G169gat), .ZN(new_n967));
  NAND3_X1  g766(.A1(new_n964), .A2(new_n966), .A3(new_n967), .ZN(new_n968));
  INV_X1    g767(.A(KEYINPUT124), .ZN(new_n969));
  OAI211_X1 g768(.A(new_n401), .B(new_n454), .C1(new_n765), .C2(new_n766), .ZN(new_n970));
  XNOR2_X1  g769(.A(new_n970), .B(KEYINPUT125), .ZN(new_n971));
  NAND3_X1  g770(.A1(new_n971), .A2(new_n683), .A3(new_n872), .ZN(new_n972));
  AOI21_X1  g771(.A(new_n969), .B1(new_n972), .B2(G169gat), .ZN(new_n973));
  NAND2_X1  g772(.A1(new_n968), .A2(new_n973), .ZN(new_n974));
  NAND4_X1  g773(.A1(new_n964), .A2(new_n966), .A3(new_n969), .A4(new_n967), .ZN(new_n975));
  AND2_X1   g774(.A1(new_n974), .A2(new_n975), .ZN(G1348gat));
  NAND4_X1  g775(.A1(new_n964), .A2(new_n966), .A3(new_n229), .A4(new_n654), .ZN(new_n977));
  NAND2_X1  g776(.A1(new_n971), .A2(new_n872), .ZN(new_n978));
  OAI21_X1  g777(.A(G176gat), .B1(new_n978), .B2(new_n655), .ZN(new_n979));
  NAND2_X1  g778(.A1(new_n977), .A2(new_n979), .ZN(G1349gat));
  OAI21_X1  g779(.A(G183gat), .B1(new_n978), .B2(new_n560), .ZN(new_n981));
  NAND3_X1  g780(.A1(new_n717), .A2(new_n243), .A3(new_n245), .ZN(new_n982));
  OAI21_X1  g781(.A(new_n981), .B1(new_n965), .B2(new_n982), .ZN(new_n983));
  XNOR2_X1  g782(.A(new_n983), .B(KEYINPUT60), .ZN(G1350gat));
  NAND2_X1  g783(.A1(KEYINPUT126), .A2(KEYINPUT61), .ZN(new_n985));
  NAND3_X1  g784(.A1(new_n971), .A2(new_n630), .A3(new_n872), .ZN(new_n986));
  NOR2_X1   g785(.A1(KEYINPUT126), .A2(KEYINPUT61), .ZN(new_n987));
  INV_X1    g786(.A(new_n987), .ZN(new_n988));
  AND3_X1   g787(.A1(new_n986), .A2(G190gat), .A3(new_n988), .ZN(new_n989));
  AOI21_X1  g788(.A(new_n988), .B1(new_n986), .B2(G190gat), .ZN(new_n990));
  OAI21_X1  g789(.A(new_n985), .B1(new_n989), .B2(new_n990), .ZN(new_n991));
  NAND4_X1  g790(.A1(new_n964), .A2(new_n966), .A3(new_n217), .A4(new_n728), .ZN(new_n992));
  NAND2_X1  g791(.A1(new_n991), .A2(new_n992), .ZN(G1351gat));
  NOR3_X1   g792(.A1(new_n767), .A2(new_n741), .A3(new_n288), .ZN(new_n994));
  NAND2_X1  g793(.A1(new_n947), .A2(new_n994), .ZN(new_n995));
  NOR3_X1   g794(.A1(new_n995), .A2(new_n256), .A3(new_n684), .ZN(new_n996));
  NAND3_X1  g795(.A1(new_n959), .A2(new_n452), .A3(new_n963), .ZN(new_n997));
  OR2_X1    g796(.A1(new_n997), .A2(new_n684), .ZN(new_n998));
  AOI21_X1  g797(.A(new_n996), .B1(new_n998), .B2(new_n256), .ZN(G1352gat));
  NAND2_X1  g798(.A1(new_n654), .A2(new_n251), .ZN(new_n1000));
  OR3_X1    g799(.A1(new_n997), .A2(KEYINPUT62), .A3(new_n1000), .ZN(new_n1001));
  OAI21_X1  g800(.A(G204gat), .B1(new_n995), .B2(new_n655), .ZN(new_n1002));
  OAI21_X1  g801(.A(KEYINPUT62), .B1(new_n997), .B2(new_n1000), .ZN(new_n1003));
  NAND3_X1  g802(.A1(new_n1001), .A2(new_n1002), .A3(new_n1003), .ZN(G1353gat));
  NAND3_X1  g803(.A1(new_n947), .A2(new_n717), .A3(new_n994), .ZN(new_n1005));
  AND3_X1   g804(.A1(new_n1005), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n1006));
  AOI21_X1  g805(.A(KEYINPUT63), .B1(new_n1005), .B2(G211gat), .ZN(new_n1007));
  OR2_X1    g806(.A1(new_n560), .A2(G211gat), .ZN(new_n1008));
  OAI22_X1  g807(.A1(new_n1006), .A2(new_n1007), .B1(new_n997), .B2(new_n1008), .ZN(G1354gat));
  NAND2_X1  g808(.A1(new_n630), .A2(G218gat), .ZN(new_n1010));
  XNOR2_X1  g809(.A(new_n1010), .B(KEYINPUT127), .ZN(new_n1011));
  NOR2_X1   g810(.A1(new_n995), .A2(new_n1011), .ZN(new_n1012));
  OR2_X1    g811(.A1(new_n997), .A2(new_n729), .ZN(new_n1013));
  INV_X1    g812(.A(G218gat), .ZN(new_n1014));
  AOI21_X1  g813(.A(new_n1012), .B1(new_n1013), .B2(new_n1014), .ZN(G1355gat));
endmodule


