

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359,
         n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370,
         n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381,
         n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392,
         n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403,
         n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414,
         n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425,
         n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436,
         n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447,
         n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458,
         n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469,
         n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480,
         n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491,
         n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502,
         n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n513,
         n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
         n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
         n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590,
         n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601,
         n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612,
         n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623,
         n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634,
         n635, n636, n637, n638, n639, n640, n641, n642, n643, n644, n645,
         n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, n656,
         n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n667,
         n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678,
         n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689,
         n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700,
         n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711,
         n712, n713, n714, n715, n716, n717, n718, n719, n720, n721, n722,
         n723, n724, n725, n726, n727, n728, n729, n730, n731, n732, n733,
         n734;

  XNOR2_X1 U370 ( .A(n717), .B(n451), .ZN(n478) );
  NAND2_X1 U371 ( .A1(n381), .A2(n377), .ZN(n645) );
  INV_X2 U372 ( .A(G953), .ZN(n719) );
  OR2_X1 U373 ( .A1(n614), .A2(n613), .ZN(n349) );
  OR2_X1 U374 ( .A1(n635), .A2(n620), .ZN(n350) );
  INV_X1 U375 ( .A(n563), .ZN(n647) );
  XNOR2_X2 U376 ( .A(n506), .B(KEYINPUT0), .ZN(n544) );
  NOR2_X2 U377 ( .A1(n595), .A2(n505), .ZN(n506) );
  XNOR2_X2 U378 ( .A(n373), .B(n356), .ZN(n672) );
  XNOR2_X1 U379 ( .A(G902), .B(KEYINPUT15), .ZN(n610) );
  INV_X1 U380 ( .A(G469), .ZN(n472) );
  AND2_X1 U381 ( .A1(n445), .A2(n444), .ZN(n617) );
  NAND2_X1 U382 ( .A1(n402), .A2(n349), .ZN(n448) );
  NAND2_X1 U383 ( .A1(n384), .A2(n357), .ZN(n402) );
  NOR2_X1 U384 ( .A1(n675), .A2(n610), .ZN(n555) );
  XNOR2_X1 U385 ( .A(n580), .B(KEYINPUT40), .ZN(n731) );
  XNOR2_X1 U386 ( .A(n542), .B(n541), .ZN(n635) );
  XNOR2_X1 U387 ( .A(KEYINPUT108), .B(n549), .ZN(n734) );
  XNOR2_X1 U388 ( .A(n546), .B(KEYINPUT104), .ZN(n620) );
  AND2_X1 U389 ( .A1(n544), .A2(n399), .ZN(n542) );
  AND2_X1 U390 ( .A1(n544), .A2(n404), .ZN(n546) );
  INV_X1 U391 ( .A(n652), .ZN(n399) );
  AND2_X1 U392 ( .A1(n545), .A2(n405), .ZN(n404) );
  INV_X1 U393 ( .A(n584), .ZN(n405) );
  XNOR2_X1 U394 ( .A(n465), .B(n352), .ZN(n434) );
  XNOR2_X1 U395 ( .A(n491), .B(G134), .ZN(n519) );
  INV_X1 U396 ( .A(n647), .ZN(n351) );
  XNOR2_X1 U397 ( .A(n481), .B(n480), .ZN(n563) );
  XNOR2_X1 U398 ( .A(n554), .B(n553), .ZN(n675) );
  XNOR2_X1 U399 ( .A(n519), .B(n470), .ZN(n717) );
  XNOR2_X1 U400 ( .A(G131), .B(KEYINPUT69), .ZN(n400) );
  XNOR2_X1 U401 ( .A(n568), .B(KEYINPUT1), .ZN(n607) );
  OR2_X1 U402 ( .A1(n701), .A2(n378), .ZN(n377) );
  NAND2_X1 U403 ( .A1(n380), .A2(n379), .ZN(n378) );
  INV_X1 U404 ( .A(G902), .ZN(n379) );
  INV_X1 U405 ( .A(n434), .ZN(n380) );
  AND2_X1 U406 ( .A1(n383), .A2(n382), .ZN(n381) );
  NAND2_X1 U407 ( .A1(n434), .A2(G902), .ZN(n382) );
  XNOR2_X1 U408 ( .A(n647), .B(n410), .ZN(n573) );
  INV_X1 U409 ( .A(KEYINPUT6), .ZN(n410) );
  XNOR2_X1 U410 ( .A(n485), .B(n484), .ZN(n442) );
  XNOR2_X1 U411 ( .A(n514), .B(n424), .ZN(n694) );
  XNOR2_X1 U412 ( .A(n427), .B(n425), .ZN(n424) );
  XNOR2_X1 U413 ( .A(n515), .B(n426), .ZN(n425) );
  NOR2_X1 U414 ( .A1(n629), .A2(n423), .ZN(n422) );
  INV_X1 U415 ( .A(KEYINPUT74), .ZN(n423) );
  XNOR2_X1 U416 ( .A(n361), .B(KEYINPUT77), .ZN(n508) );
  NAND2_X1 U417 ( .A1(n719), .A2(n362), .ZN(n361) );
  INV_X1 U418 ( .A(G237), .ZN(n362) );
  XNOR2_X1 U419 ( .A(G146), .B(G125), .ZN(n494) );
  INV_X1 U420 ( .A(KEYINPUT107), .ZN(n416) );
  XOR2_X1 U421 ( .A(KEYINPUT5), .B(KEYINPUT102), .Z(n475) );
  XNOR2_X1 U422 ( .A(n440), .B(n439), .ZN(n486) );
  XNOR2_X1 U423 ( .A(G119), .B(G116), .ZN(n439) );
  XNOR2_X1 U424 ( .A(n441), .B(G113), .ZN(n440) );
  XNOR2_X1 U425 ( .A(KEYINPUT92), .B(KEYINPUT3), .ZN(n441) );
  XNOR2_X1 U426 ( .A(n494), .B(n371), .ZN(n513) );
  XNOR2_X1 U427 ( .A(KEYINPUT10), .B(KEYINPUT68), .ZN(n371) );
  XOR2_X1 U428 ( .A(G137), .B(G140), .Z(n468) );
  XNOR2_X1 U429 ( .A(n413), .B(n412), .ZN(n485) );
  XNOR2_X1 U430 ( .A(G107), .B(G104), .ZN(n412) );
  XNOR2_X1 U431 ( .A(n414), .B(G110), .ZN(n413) );
  INV_X1 U432 ( .A(KEYINPUT76), .ZN(n414) );
  XNOR2_X1 U433 ( .A(n471), .B(G146), .ZN(n451) );
  XOR2_X1 U434 ( .A(G101), .B(KEYINPUT67), .Z(n487) );
  XNOR2_X1 U435 ( .A(KEYINPUT4), .B(KEYINPUT17), .ZN(n488) );
  OR2_X1 U436 ( .A1(n605), .A2(n395), .ZN(n614) );
  INV_X1 U437 ( .A(n640), .ZN(n396) );
  NOR2_X1 U438 ( .A1(n644), .A2(n561), .ZN(n571) );
  XNOR2_X1 U439 ( .A(G119), .B(KEYINPUT97), .ZN(n454) );
  XNOR2_X1 U440 ( .A(G128), .B(G110), .ZN(n457) );
  XNOR2_X1 U441 ( .A(n513), .B(n468), .ZN(n716) );
  XNOR2_X1 U442 ( .A(n436), .B(n435), .ZN(n522) );
  INV_X1 U443 ( .A(KEYINPUT8), .ZN(n435) );
  NAND2_X1 U444 ( .A1(n719), .A2(G234), .ZN(n436) );
  NAND2_X1 U445 ( .A1(n370), .A2(n369), .ZN(n368) );
  NOR2_X1 U446 ( .A1(n401), .A2(n657), .ZN(n369) );
  XNOR2_X1 U447 ( .A(n586), .B(KEYINPUT41), .ZN(n671) );
  NOR2_X1 U448 ( .A1(n592), .A2(n658), .ZN(n570) );
  XNOR2_X1 U449 ( .A(n372), .B(KEYINPUT34), .ZN(n527) );
  INV_X1 U450 ( .A(KEYINPUT81), .ZN(n409) );
  XNOR2_X1 U451 ( .A(n495), .B(KEYINPUT93), .ZN(n443) );
  NOR2_X1 U452 ( .A1(n584), .A2(n583), .ZN(n597) );
  NOR2_X1 U453 ( .A1(n647), .A2(n581), .ZN(n582) );
  XNOR2_X1 U454 ( .A(n516), .B(n429), .ZN(n537) );
  XNOR2_X1 U455 ( .A(KEYINPUT13), .B(G475), .ZN(n429) );
  XNOR2_X1 U456 ( .A(n531), .B(n355), .ZN(n388) );
  AND2_X1 U457 ( .A1(n544), .A2(n353), .ZN(n531) );
  NOR2_X1 U458 ( .A1(n448), .A2(n420), .ZN(n419) );
  INV_X1 U459 ( .A(G475), .ZN(n420) );
  XNOR2_X1 U460 ( .A(n682), .B(n681), .ZN(n683) );
  INV_X1 U461 ( .A(n637), .ZN(n408) );
  XNOR2_X1 U462 ( .A(n421), .B(KEYINPUT47), .ZN(n601) );
  XNOR2_X1 U463 ( .A(n556), .B(n397), .ZN(n557) );
  INV_X1 U464 ( .A(KEYINPUT111), .ZN(n397) );
  NOR2_X1 U465 ( .A1(n375), .A2(n374), .ZN(n543) );
  INV_X1 U466 ( .A(n381), .ZN(n374) );
  NAND2_X1 U467 ( .A1(n377), .A2(n376), .ZN(n375) );
  XNOR2_X1 U468 ( .A(G104), .B(G140), .ZN(n507) );
  INV_X1 U469 ( .A(KEYINPUT106), .ZN(n426) );
  XNOR2_X1 U470 ( .A(n512), .B(n511), .ZN(n427) );
  XNOR2_X1 U471 ( .A(G143), .B(G131), .ZN(n509) );
  XNOR2_X1 U472 ( .A(n552), .B(KEYINPUT87), .ZN(n553) );
  OR2_X1 U473 ( .A1(G237), .A2(G902), .ZN(n496) );
  XNOR2_X1 U474 ( .A(n411), .B(n486), .ZN(n479) );
  XNOR2_X1 U475 ( .A(n477), .B(n476), .ZN(n411) );
  XNOR2_X1 U476 ( .A(G116), .B(G107), .ZN(n517) );
  XNOR2_X1 U477 ( .A(n469), .B(n468), .ZN(n450) );
  XNOR2_X1 U478 ( .A(n709), .B(n390), .ZN(n680) );
  XNOR2_X1 U479 ( .A(n493), .B(n391), .ZN(n390) );
  XNOR2_X1 U480 ( .A(n392), .B(n487), .ZN(n391) );
  XNOR2_X1 U481 ( .A(n564), .B(n565), .ZN(n406) );
  INV_X1 U482 ( .A(G472), .ZN(n447) );
  XNOR2_X1 U483 ( .A(n461), .B(n460), .ZN(n462) );
  INV_X1 U484 ( .A(n448), .ZN(n699) );
  XNOR2_X1 U485 ( .A(n363), .B(KEYINPUT84), .ZN(n676) );
  NAND2_X1 U486 ( .A1(n349), .A2(n364), .ZN(n363) );
  NAND2_X1 U487 ( .A1(n365), .A2(n612), .ZN(n364) );
  NAND2_X1 U488 ( .A1(n385), .A2(n704), .ZN(n365) );
  AND2_X1 U489 ( .A1(n367), .A2(n366), .ZN(n609) );
  INV_X1 U490 ( .A(n608), .ZN(n366) );
  XNOR2_X1 U491 ( .A(n368), .B(KEYINPUT43), .ZN(n367) );
  XNOR2_X1 U492 ( .A(n587), .B(KEYINPUT42), .ZN(n733) );
  NOR2_X1 U493 ( .A1(n527), .A2(n526), .ZN(n529) );
  NOR2_X1 U494 ( .A1(n642), .A2(n533), .ZN(n534) );
  NAND2_X1 U495 ( .A1(n597), .A2(n596), .ZN(n629) );
  INV_X1 U496 ( .A(n537), .ZN(n538) );
  OR2_X1 U497 ( .A1(n437), .A2(n394), .ZN(n393) );
  INV_X1 U498 ( .A(n645), .ZN(n394) );
  AND2_X1 U499 ( .A1(n537), .A2(n428), .ZN(n632) );
  INV_X1 U500 ( .A(n539), .ZN(n428) );
  NAND2_X1 U501 ( .A1(n548), .A2(n642), .ZN(n438) );
  INV_X1 U502 ( .A(KEYINPUT60), .ZN(n359) );
  XNOR2_X1 U503 ( .A(n389), .B(n683), .ZN(n684) );
  INV_X1 U504 ( .A(n644), .ZN(n376) );
  INV_X1 U505 ( .A(n401), .ZN(n642) );
  XOR2_X1 U506 ( .A(KEYINPUT101), .B(KEYINPUT25), .Z(n352) );
  AND2_X1 U507 ( .A1(n659), .A2(n376), .ZN(n353) );
  XNOR2_X1 U508 ( .A(n614), .B(KEYINPUT86), .ZN(n718) );
  AND2_X1 U509 ( .A1(n349), .A2(G210), .ZN(n354) );
  NAND2_X1 U510 ( .A1(n630), .A2(n625), .ZN(n661) );
  XOR2_X1 U511 ( .A(n530), .B(KEYINPUT22), .Z(n355) );
  XNOR2_X1 U512 ( .A(n482), .B(KEYINPUT110), .ZN(n356) );
  OR2_X1 U513 ( .A1(n612), .A2(n611), .ZN(n357) );
  XNOR2_X1 U514 ( .A(n442), .B(n486), .ZN(n709) );
  XNOR2_X1 U515 ( .A(n478), .B(n449), .ZN(n687) );
  XNOR2_X1 U516 ( .A(KEYINPUT62), .B(n615), .ZN(n358) );
  NOR2_X1 U517 ( .A1(G952), .A2(n719), .ZN(n703) );
  INV_X1 U518 ( .A(n703), .ZN(n444) );
  XNOR2_X1 U519 ( .A(n573), .B(n409), .ZN(n532) );
  XNOR2_X1 U520 ( .A(n360), .B(n359), .ZN(G60) );
  NAND2_X1 U521 ( .A1(n418), .A2(n444), .ZN(n360) );
  INV_X1 U522 ( .A(n606), .ZN(n370) );
  NAND2_X1 U523 ( .A1(n672), .A2(n544), .ZN(n372) );
  NAND2_X1 U524 ( .A1(n540), .A2(n547), .ZN(n373) );
  NAND2_X1 U525 ( .A1(n701), .A2(n434), .ZN(n383) );
  XNOR2_X1 U526 ( .A(n462), .B(n463), .ZN(n701) );
  NAND2_X1 U527 ( .A1(n386), .A2(n385), .ZN(n384) );
  INV_X1 U528 ( .A(n718), .ZN(n385) );
  XNOR2_X1 U529 ( .A(n555), .B(n387), .ZN(n386) );
  INV_X1 U530 ( .A(KEYINPUT83), .ZN(n387) );
  NOR2_X1 U531 ( .A1(n388), .A2(n535), .ZN(n536) );
  OR2_X1 U532 ( .A1(n388), .A2(n438), .ZN(n549) );
  OR2_X1 U533 ( .A1(n388), .A2(n393), .ZN(n624) );
  NAND2_X1 U534 ( .A1(n402), .A2(n354), .ZN(n389) );
  NAND2_X1 U535 ( .A1(n680), .A2(n610), .ZN(n415) );
  XNOR2_X1 U536 ( .A(n492), .B(n494), .ZN(n392) );
  NOR2_X1 U537 ( .A1(n684), .A2(n703), .ZN(n686) );
  NAND2_X1 U538 ( .A1(n661), .A2(n422), .ZN(n421) );
  NAND2_X1 U539 ( .A1(n729), .A2(n396), .ZN(n395) );
  NAND2_X1 U540 ( .A1(n502), .A2(G953), .ZN(n556) );
  NAND2_X1 U541 ( .A1(n551), .A2(n398), .ZN(n554) );
  XNOR2_X1 U542 ( .A(n550), .B(KEYINPUT109), .ZN(n398) );
  INV_X1 U543 ( .A(n400), .ZN(n453) );
  BUF_X1 U544 ( .A(n607), .Z(n401) );
  XNOR2_X1 U545 ( .A(n536), .B(KEYINPUT32), .ZN(n730) );
  NAND2_X1 U546 ( .A1(n403), .A2(n734), .ZN(n550) );
  XNOR2_X1 U547 ( .A(n417), .B(n416), .ZN(n403) );
  NAND2_X1 U548 ( .A1(n406), .A2(n571), .ZN(n566) );
  NOR2_X1 U549 ( .A1(n407), .A2(n590), .ZN(n604) );
  NAND2_X1 U550 ( .A1(n603), .A2(n408), .ZN(n407) );
  NAND2_X1 U551 ( .A1(n350), .A2(n661), .ZN(n417) );
  NOR2_X1 U552 ( .A1(n730), .A2(n433), .ZN(n432) );
  NAND2_X1 U553 ( .A1(n608), .A2(n562), .ZN(n576) );
  XNOR2_X2 U554 ( .A(n415), .B(n443), .ZN(n608) );
  XNOR2_X1 U555 ( .A(n419), .B(n695), .ZN(n418) );
  XNOR2_X1 U556 ( .A(n431), .B(n430), .ZN(n551) );
  INV_X1 U557 ( .A(KEYINPUT44), .ZN(n430) );
  NAND2_X1 U558 ( .A1(n432), .A2(n726), .ZN(n431) );
  XNOR2_X1 U559 ( .A(n529), .B(n528), .ZN(n726) );
  INV_X1 U560 ( .A(n624), .ZN(n433) );
  OR2_X1 U561 ( .A1(n351), .A2(n401), .ZN(n437) );
  NAND2_X1 U562 ( .A1(n543), .A2(n607), .ZN(n474) );
  XNOR2_X2 U563 ( .A(n473), .B(n472), .ZN(n568) );
  XNOR2_X1 U564 ( .A(n446), .B(n358), .ZN(n445) );
  NOR2_X2 U565 ( .A1(n448), .A2(n447), .ZN(n446) );
  XNOR2_X1 U566 ( .A(n485), .B(n450), .ZN(n449) );
  NOR2_X2 U567 ( .A1(G902), .A2(n687), .ZN(n473) );
  XOR2_X1 U568 ( .A(KEYINPUT48), .B(KEYINPUT90), .Z(n452) );
  XNOR2_X1 U569 ( .A(n483), .B(KEYINPUT16), .ZN(n484) );
  XNOR2_X1 U570 ( .A(n475), .B(G137), .ZN(n476) );
  INV_X1 U571 ( .A(n487), .ZN(n471) );
  INV_X1 U572 ( .A(KEYINPUT19), .ZN(n498) );
  INV_X1 U573 ( .A(n568), .ZN(n584) );
  XNOR2_X1 U574 ( .A(n694), .B(n693), .ZN(n695) );
  INV_X1 U575 ( .A(KEYINPUT39), .ZN(n569) );
  XNOR2_X1 U576 ( .A(KEYINPUT63), .B(KEYINPUT117), .ZN(n616) );
  XOR2_X1 U577 ( .A(KEYINPUT99), .B(KEYINPUT100), .Z(n455) );
  XNOR2_X1 U578 ( .A(n455), .B(n454), .ZN(n456) );
  XNOR2_X1 U579 ( .A(n716), .B(n456), .ZN(n463) );
  XOR2_X1 U580 ( .A(KEYINPUT98), .B(KEYINPUT23), .Z(n458) );
  XNOR2_X1 U581 ( .A(n458), .B(n457), .ZN(n459) );
  XOR2_X1 U582 ( .A(n459), .B(KEYINPUT24), .Z(n461) );
  NAND2_X1 U583 ( .A1(n522), .A2(G221), .ZN(n460) );
  NAND2_X1 U584 ( .A1(G234), .A2(n610), .ZN(n464) );
  XNOR2_X1 U585 ( .A(KEYINPUT20), .B(n464), .ZN(n466) );
  NAND2_X1 U586 ( .A1(n466), .A2(G217), .ZN(n465) );
  NAND2_X1 U587 ( .A1(n466), .A2(G221), .ZN(n467) );
  XNOR2_X1 U588 ( .A(n467), .B(KEYINPUT21), .ZN(n644) );
  NAND2_X1 U589 ( .A1(G227), .A2(n719), .ZN(n469) );
  XNOR2_X2 U590 ( .A(G143), .B(G128), .ZN(n491) );
  XNOR2_X1 U591 ( .A(KEYINPUT4), .B(n453), .ZN(n470) );
  XNOR2_X1 U592 ( .A(n474), .B(KEYINPUT75), .ZN(n540) );
  NAND2_X1 U593 ( .A1(n508), .A2(G210), .ZN(n477) );
  XNOR2_X1 U594 ( .A(n478), .B(n479), .ZN(n615) );
  NOR2_X1 U595 ( .A1(n615), .A2(G902), .ZN(n481) );
  XNOR2_X1 U596 ( .A(G472), .B(KEYINPUT103), .ZN(n480) );
  INV_X1 U597 ( .A(n573), .ZN(n547) );
  XOR2_X1 U598 ( .A(KEYINPUT33), .B(KEYINPUT71), .Z(n482) );
  XNOR2_X1 U599 ( .A(KEYINPUT73), .B(G122), .ZN(n483) );
  XOR2_X1 U600 ( .A(KEYINPUT78), .B(KEYINPUT18), .Z(n489) );
  XNOR2_X1 U601 ( .A(n489), .B(n488), .ZN(n490) );
  XNOR2_X1 U602 ( .A(n491), .B(n490), .ZN(n493) );
  NAND2_X1 U603 ( .A1(G224), .A2(n719), .ZN(n492) );
  NAND2_X1 U604 ( .A1(n496), .A2(G210), .ZN(n495) );
  NAND2_X1 U605 ( .A1(G214), .A2(n496), .ZN(n497) );
  XOR2_X1 U606 ( .A(KEYINPUT94), .B(n497), .Z(n657) );
  INV_X1 U607 ( .A(n657), .ZN(n562) );
  XNOR2_X1 U608 ( .A(n576), .B(n498), .ZN(n595) );
  NAND2_X1 U609 ( .A1(G234), .A2(G237), .ZN(n499) );
  XNOR2_X1 U610 ( .A(n499), .B(KEYINPUT14), .ZN(n500) );
  NAND2_X1 U611 ( .A1(G952), .A2(n500), .ZN(n670) );
  NOR2_X1 U612 ( .A1(G953), .A2(n670), .ZN(n559) );
  NAND2_X1 U613 ( .A1(G902), .A2(n500), .ZN(n501) );
  XNOR2_X1 U614 ( .A(KEYINPUT95), .B(n501), .ZN(n502) );
  NOR2_X1 U615 ( .A1(G898), .A2(n556), .ZN(n503) );
  NOR2_X1 U616 ( .A1(n559), .A2(n503), .ZN(n504) );
  XNOR2_X1 U617 ( .A(n504), .B(KEYINPUT96), .ZN(n505) );
  XNOR2_X1 U618 ( .A(n507), .B(KEYINPUT11), .ZN(n515) );
  NAND2_X1 U619 ( .A1(G214), .A2(n508), .ZN(n512) );
  XOR2_X1 U620 ( .A(G122), .B(G113), .Z(n510) );
  XNOR2_X1 U621 ( .A(n510), .B(n509), .ZN(n511) );
  XOR2_X1 U622 ( .A(n513), .B(KEYINPUT12), .Z(n514) );
  NOR2_X1 U623 ( .A1(G902), .A2(n694), .ZN(n516) );
  XNOR2_X1 U624 ( .A(n517), .B(KEYINPUT7), .ZN(n518) );
  XOR2_X1 U625 ( .A(n518), .B(KEYINPUT9), .Z(n521) );
  XNOR2_X1 U626 ( .A(n519), .B(G122), .ZN(n520) );
  XNOR2_X1 U627 ( .A(n521), .B(n520), .ZN(n524) );
  NAND2_X1 U628 ( .A1(n522), .A2(G217), .ZN(n523) );
  XOR2_X1 U629 ( .A(n524), .B(n523), .Z(n697) );
  NOR2_X1 U630 ( .A1(G902), .A2(n697), .ZN(n525) );
  XOR2_X1 U631 ( .A(G478), .B(n525), .Z(n539) );
  NAND2_X1 U632 ( .A1(n537), .A2(n539), .ZN(n591) );
  XOR2_X1 U633 ( .A(n591), .B(KEYINPUT79), .Z(n526) );
  XNOR2_X1 U634 ( .A(KEYINPUT88), .B(KEYINPUT35), .ZN(n528) );
  NOR2_X1 U635 ( .A1(n537), .A2(n539), .ZN(n659) );
  XOR2_X1 U636 ( .A(KEYINPUT72), .B(KEYINPUT65), .Z(n530) );
  NAND2_X1 U637 ( .A1(n532), .A2(n645), .ZN(n533) );
  XOR2_X1 U638 ( .A(KEYINPUT80), .B(n534), .Z(n535) );
  INV_X1 U639 ( .A(n632), .ZN(n630) );
  NAND2_X1 U640 ( .A1(n539), .A2(n538), .ZN(n625) );
  INV_X1 U641 ( .A(n661), .ZN(n599) );
  NAND2_X1 U642 ( .A1(n351), .A2(n540), .ZN(n652) );
  XNOR2_X1 U643 ( .A(KEYINPUT105), .B(KEYINPUT31), .ZN(n541) );
  INV_X1 U644 ( .A(n543), .ZN(n641) );
  NOR2_X1 U645 ( .A1(n351), .A2(n641), .ZN(n545) );
  NOR2_X1 U646 ( .A1(n547), .A2(n645), .ZN(n548) );
  XNOR2_X1 U647 ( .A(KEYINPUT45), .B(KEYINPUT64), .ZN(n552) );
  NOR2_X1 U648 ( .A1(G900), .A2(n557), .ZN(n558) );
  NOR2_X1 U649 ( .A1(n559), .A2(n558), .ZN(n560) );
  XNOR2_X1 U650 ( .A(n560), .B(KEYINPUT82), .ZN(n561) );
  XOR2_X1 U651 ( .A(KEYINPUT114), .B(KEYINPUT30), .Z(n565) );
  NAND2_X1 U652 ( .A1(n563), .A2(n562), .ZN(n564) );
  NOR2_X1 U653 ( .A1(n645), .A2(n566), .ZN(n567) );
  NAND2_X1 U654 ( .A1(n568), .A2(n567), .ZN(n592) );
  XNOR2_X1 U655 ( .A(n608), .B(KEYINPUT38), .ZN(n658) );
  XNOR2_X1 U656 ( .A(n570), .B(n569), .ZN(n579) );
  INV_X1 U657 ( .A(n625), .ZN(n634) );
  AND2_X1 U658 ( .A1(n579), .A2(n634), .ZN(n640) );
  XNOR2_X1 U659 ( .A(KEYINPUT70), .B(n571), .ZN(n572) );
  NAND2_X1 U660 ( .A1(n572), .A2(n645), .ZN(n581) );
  NOR2_X1 U661 ( .A1(n573), .A2(n581), .ZN(n574) );
  XNOR2_X1 U662 ( .A(KEYINPUT112), .B(n574), .ZN(n575) );
  NAND2_X1 U663 ( .A1(n575), .A2(n632), .ZN(n606) );
  NOR2_X1 U664 ( .A1(n606), .A2(n576), .ZN(n577) );
  XOR2_X1 U665 ( .A(KEYINPUT36), .B(n577), .Z(n578) );
  NOR2_X1 U666 ( .A1(n642), .A2(n578), .ZN(n637) );
  NAND2_X1 U667 ( .A1(n579), .A2(n632), .ZN(n580) );
  XOR2_X1 U668 ( .A(KEYINPUT28), .B(n582), .Z(n583) );
  NOR2_X1 U669 ( .A1(n658), .A2(n657), .ZN(n585) );
  XNOR2_X1 U670 ( .A(n585), .B(KEYINPUT116), .ZN(n662) );
  NAND2_X1 U671 ( .A1(n662), .A2(n659), .ZN(n586) );
  NAND2_X1 U672 ( .A1(n597), .A2(n671), .ZN(n587) );
  NAND2_X1 U673 ( .A1(n731), .A2(n733), .ZN(n589) );
  XOR2_X1 U674 ( .A(KEYINPUT46), .B(KEYINPUT91), .Z(n588) );
  XNOR2_X1 U675 ( .A(n589), .B(n588), .ZN(n590) );
  NOR2_X1 U676 ( .A1(n592), .A2(n591), .ZN(n593) );
  NAND2_X1 U677 ( .A1(n593), .A2(n608), .ZN(n594) );
  XOR2_X1 U678 ( .A(KEYINPUT115), .B(n594), .Z(n728) );
  INV_X1 U679 ( .A(n595), .ZN(n596) );
  NOR2_X1 U680 ( .A1(KEYINPUT74), .A2(n629), .ZN(n598) );
  NAND2_X1 U681 ( .A1(n599), .A2(n598), .ZN(n600) );
  NAND2_X1 U682 ( .A1(n728), .A2(n600), .ZN(n602) );
  NOR2_X1 U683 ( .A1(n602), .A2(n601), .ZN(n603) );
  XNOR2_X1 U684 ( .A(n604), .B(n452), .ZN(n605) );
  XNOR2_X1 U685 ( .A(KEYINPUT113), .B(n609), .ZN(n729) );
  INV_X1 U686 ( .A(KEYINPUT2), .ZN(n612) );
  XOR2_X1 U687 ( .A(KEYINPUT85), .B(n610), .Z(n611) );
  INV_X1 U688 ( .A(n675), .ZN(n704) );
  NAND2_X1 U689 ( .A1(KEYINPUT2), .A2(n704), .ZN(n613) );
  XNOR2_X1 U690 ( .A(n617), .B(n616), .ZN(G57) );
  NAND2_X1 U691 ( .A1(n620), .A2(n632), .ZN(n618) );
  XNOR2_X1 U692 ( .A(n618), .B(KEYINPUT118), .ZN(n619) );
  XNOR2_X1 U693 ( .A(G104), .B(n619), .ZN(G6) );
  XOR2_X1 U694 ( .A(KEYINPUT27), .B(KEYINPUT26), .Z(n622) );
  NAND2_X1 U695 ( .A1(n634), .A2(n620), .ZN(n621) );
  XNOR2_X1 U696 ( .A(n622), .B(n621), .ZN(n623) );
  XNOR2_X1 U697 ( .A(G107), .B(n623), .ZN(G9) );
  XNOR2_X1 U698 ( .A(n624), .B(G110), .ZN(G12) );
  NOR2_X1 U699 ( .A1(n629), .A2(n625), .ZN(n627) );
  XNOR2_X1 U700 ( .A(KEYINPUT29), .B(KEYINPUT119), .ZN(n626) );
  XNOR2_X1 U701 ( .A(n627), .B(n626), .ZN(n628) );
  XOR2_X1 U702 ( .A(G128), .B(n628), .Z(G30) );
  NOR2_X1 U703 ( .A1(n630), .A2(n629), .ZN(n631) );
  XOR2_X1 U704 ( .A(G146), .B(n631), .Z(G48) );
  NAND2_X1 U705 ( .A1(n635), .A2(n632), .ZN(n633) );
  XNOR2_X1 U706 ( .A(n633), .B(G113), .ZN(G15) );
  NAND2_X1 U707 ( .A1(n635), .A2(n634), .ZN(n636) );
  XNOR2_X1 U708 ( .A(n636), .B(G116), .ZN(G18) );
  XNOR2_X1 U709 ( .A(n637), .B(KEYINPUT120), .ZN(n638) );
  XNOR2_X1 U710 ( .A(n638), .B(KEYINPUT37), .ZN(n639) );
  XNOR2_X1 U711 ( .A(G125), .B(n639), .ZN(G27) );
  XOR2_X1 U712 ( .A(G134), .B(n640), .Z(G36) );
  NAND2_X1 U713 ( .A1(n642), .A2(n641), .ZN(n643) );
  XNOR2_X1 U714 ( .A(n643), .B(KEYINPUT50), .ZN(n651) );
  NAND2_X1 U715 ( .A1(n645), .A2(n644), .ZN(n646) );
  XOR2_X1 U716 ( .A(KEYINPUT49), .B(n646), .Z(n648) );
  NAND2_X1 U717 ( .A1(n648), .A2(n647), .ZN(n649) );
  XNOR2_X1 U718 ( .A(KEYINPUT121), .B(n649), .ZN(n650) );
  NAND2_X1 U719 ( .A1(n651), .A2(n650), .ZN(n653) );
  NAND2_X1 U720 ( .A1(n653), .A2(n652), .ZN(n655) );
  XOR2_X1 U721 ( .A(KEYINPUT122), .B(KEYINPUT51), .Z(n654) );
  XNOR2_X1 U722 ( .A(n655), .B(n654), .ZN(n656) );
  NAND2_X1 U723 ( .A1(n671), .A2(n656), .ZN(n667) );
  NAND2_X1 U724 ( .A1(n658), .A2(n657), .ZN(n660) );
  NAND2_X1 U725 ( .A1(n660), .A2(n659), .ZN(n664) );
  NAND2_X1 U726 ( .A1(n662), .A2(n661), .ZN(n663) );
  NAND2_X1 U727 ( .A1(n664), .A2(n663), .ZN(n665) );
  NAND2_X1 U728 ( .A1(n665), .A2(n672), .ZN(n666) );
  NAND2_X1 U729 ( .A1(n667), .A2(n666), .ZN(n668) );
  XOR2_X1 U730 ( .A(KEYINPUT52), .B(n668), .Z(n669) );
  NOR2_X1 U731 ( .A1(n670), .A2(n669), .ZN(n674) );
  AND2_X1 U732 ( .A1(n672), .A2(n671), .ZN(n673) );
  NOR2_X1 U733 ( .A1(n674), .A2(n673), .ZN(n677) );
  NAND2_X1 U734 ( .A1(n677), .A2(n676), .ZN(n678) );
  NOR2_X1 U735 ( .A1(n678), .A2(G953), .ZN(n679) );
  XNOR2_X1 U736 ( .A(n679), .B(KEYINPUT53), .ZN(G75) );
  INV_X1 U737 ( .A(n680), .ZN(n682) );
  XOR2_X1 U738 ( .A(KEYINPUT54), .B(KEYINPUT55), .Z(n681) );
  XOR2_X1 U739 ( .A(KEYINPUT89), .B(KEYINPUT56), .Z(n685) );
  XNOR2_X1 U740 ( .A(n686), .B(n685), .ZN(G51) );
  XNOR2_X1 U741 ( .A(KEYINPUT58), .B(KEYINPUT123), .ZN(n689) );
  XNOR2_X1 U742 ( .A(n687), .B(KEYINPUT57), .ZN(n688) );
  XNOR2_X1 U743 ( .A(n689), .B(n688), .ZN(n691) );
  NAND2_X1 U744 ( .A1(n699), .A2(G469), .ZN(n690) );
  XNOR2_X1 U745 ( .A(n691), .B(n690), .ZN(n692) );
  NOR2_X1 U746 ( .A1(n703), .A2(n692), .ZN(G54) );
  XOR2_X1 U747 ( .A(KEYINPUT59), .B(KEYINPUT66), .Z(n693) );
  NAND2_X1 U748 ( .A1(G478), .A2(n699), .ZN(n696) );
  XNOR2_X1 U749 ( .A(n697), .B(n696), .ZN(n698) );
  NOR2_X1 U750 ( .A1(n703), .A2(n698), .ZN(G63) );
  NAND2_X1 U751 ( .A1(G217), .A2(n699), .ZN(n700) );
  XNOR2_X1 U752 ( .A(n701), .B(n700), .ZN(n702) );
  NOR2_X1 U753 ( .A1(n703), .A2(n702), .ZN(G66) );
  NAND2_X1 U754 ( .A1(n719), .A2(n704), .ZN(n708) );
  NAND2_X1 U755 ( .A1(G953), .A2(G224), .ZN(n705) );
  XNOR2_X1 U756 ( .A(KEYINPUT61), .B(n705), .ZN(n706) );
  NAND2_X1 U757 ( .A1(n706), .A2(G898), .ZN(n707) );
  NAND2_X1 U758 ( .A1(n708), .A2(n707), .ZN(n714) );
  XOR2_X1 U759 ( .A(G101), .B(n709), .Z(n710) );
  XNOR2_X1 U760 ( .A(KEYINPUT125), .B(n710), .ZN(n712) );
  NOR2_X1 U761 ( .A1(G898), .A2(n719), .ZN(n711) );
  NOR2_X1 U762 ( .A1(n712), .A2(n711), .ZN(n713) );
  XNOR2_X1 U763 ( .A(n714), .B(n713), .ZN(n715) );
  XNOR2_X1 U764 ( .A(KEYINPUT124), .B(n715), .ZN(G69) );
  XNOR2_X1 U765 ( .A(n717), .B(n716), .ZN(n721) );
  XNOR2_X1 U766 ( .A(n721), .B(n718), .ZN(n720) );
  NAND2_X1 U767 ( .A1(n720), .A2(n719), .ZN(n725) );
  XNOR2_X1 U768 ( .A(G227), .B(n721), .ZN(n722) );
  NAND2_X1 U769 ( .A1(n722), .A2(G900), .ZN(n723) );
  NAND2_X1 U770 ( .A1(n723), .A2(G953), .ZN(n724) );
  NAND2_X1 U771 ( .A1(n725), .A2(n724), .ZN(G72) );
  XNOR2_X1 U772 ( .A(n726), .B(G122), .ZN(n727) );
  XNOR2_X1 U773 ( .A(n727), .B(KEYINPUT126), .ZN(G24) );
  XNOR2_X1 U774 ( .A(G143), .B(n728), .ZN(G45) );
  XNOR2_X1 U775 ( .A(G140), .B(n729), .ZN(G42) );
  XOR2_X1 U776 ( .A(n730), .B(G119), .Z(G21) );
  XOR2_X1 U777 ( .A(G131), .B(n731), .Z(n732) );
  XNOR2_X1 U778 ( .A(KEYINPUT127), .B(n732), .ZN(G33) );
  XNOR2_X1 U779 ( .A(G137), .B(n733), .ZN(G39) );
  XNOR2_X1 U780 ( .A(G101), .B(n734), .ZN(G3) );
endmodule

