//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 1 0 1 1 0 1 1 0 0 1 0 1 0 0 1 0 1 1 0 0 0 0 1 0 1 1 0 1 1 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 0 1 1 1 0 0 0 0 0 0 0 0 1 1 1 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:17:27 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n608,
    new_n609, new_n610, new_n611, new_n612, new_n613, new_n614, new_n615,
    new_n616, new_n617, new_n619, new_n620, new_n621, new_n622, new_n623,
    new_n624, new_n625, new_n626, new_n628, new_n629, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n681, new_n682, new_n683, new_n684, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n692, new_n693,
    new_n694, new_n695, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n705, new_n706, new_n708, new_n709, new_n710,
    new_n711, new_n712, new_n713, new_n714, new_n715, new_n716, new_n717,
    new_n718, new_n719, new_n720, new_n721, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n743, new_n744, new_n745, new_n746, new_n747, new_n748, new_n749,
    new_n750, new_n751, new_n752, new_n753, new_n754, new_n755, new_n756,
    new_n757, new_n758, new_n759, new_n760, new_n761, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n790, new_n791, new_n793,
    new_n794, new_n796, new_n797, new_n798, new_n799, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n866, new_n867,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n881, new_n882, new_n884, new_n885,
    new_n886, new_n887, new_n888, new_n889, new_n890, new_n891, new_n893,
    new_n894, new_n895, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n903, new_n904, new_n905, new_n906, new_n908, new_n909, new_n910,
    new_n911, new_n913, new_n914, new_n915;
  INV_X1    g000(.A(KEYINPUT69), .ZN(new_n202));
  NAND2_X1  g001(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n203));
  INV_X1    g002(.A(new_n203), .ZN(new_n204));
  NOR2_X1   g003(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n205));
  NOR2_X1   g004(.A1(new_n204), .A2(new_n205), .ZN(new_n206));
  XNOR2_X1  g005(.A(KEYINPUT68), .B(G190gat), .ZN(new_n207));
  OAI21_X1  g006(.A(new_n202), .B1(new_n206), .B2(new_n207), .ZN(new_n208));
  INV_X1    g007(.A(G190gat), .ZN(new_n209));
  NAND2_X1  g008(.A1(new_n209), .A2(KEYINPUT68), .ZN(new_n210));
  INV_X1    g009(.A(KEYINPUT68), .ZN(new_n211));
  NAND2_X1  g010(.A1(new_n211), .A2(G190gat), .ZN(new_n212));
  NAND2_X1  g011(.A1(new_n210), .A2(new_n212), .ZN(new_n213));
  XNOR2_X1  g012(.A(KEYINPUT27), .B(G183gat), .ZN(new_n214));
  NAND3_X1  g013(.A1(new_n213), .A2(new_n214), .A3(KEYINPUT69), .ZN(new_n215));
  AOI21_X1  g014(.A(KEYINPUT28), .B1(new_n208), .B2(new_n215), .ZN(new_n216));
  INV_X1    g015(.A(KEYINPUT28), .ZN(new_n217));
  INV_X1    g016(.A(KEYINPUT70), .ZN(new_n218));
  OAI21_X1  g017(.A(new_n218), .B1(new_n204), .B2(new_n205), .ZN(new_n219));
  INV_X1    g018(.A(KEYINPUT27), .ZN(new_n220));
  INV_X1    g019(.A(G183gat), .ZN(new_n221));
  NAND2_X1  g020(.A1(new_n220), .A2(new_n221), .ZN(new_n222));
  NAND3_X1  g021(.A1(new_n222), .A2(KEYINPUT70), .A3(new_n203), .ZN(new_n223));
  NAND2_X1  g022(.A1(new_n219), .A2(new_n223), .ZN(new_n224));
  AOI21_X1  g023(.A(new_n217), .B1(new_n224), .B2(new_n213), .ZN(new_n225));
  OAI21_X1  g024(.A(KEYINPUT71), .B1(new_n216), .B2(new_n225), .ZN(new_n226));
  AND3_X1   g025(.A1(new_n213), .A2(new_n214), .A3(KEYINPUT69), .ZN(new_n227));
  AOI21_X1  g026(.A(KEYINPUT69), .B1(new_n213), .B2(new_n214), .ZN(new_n228));
  OAI21_X1  g027(.A(new_n217), .B1(new_n227), .B2(new_n228), .ZN(new_n229));
  NOR3_X1   g028(.A1(new_n204), .A2(new_n205), .A3(new_n218), .ZN(new_n230));
  AOI21_X1  g029(.A(KEYINPUT70), .B1(new_n222), .B2(new_n203), .ZN(new_n231));
  OAI21_X1  g030(.A(new_n213), .B1(new_n230), .B2(new_n231), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n232), .A2(KEYINPUT28), .ZN(new_n233));
  INV_X1    g032(.A(KEYINPUT71), .ZN(new_n234));
  NAND3_X1  g033(.A1(new_n229), .A2(new_n233), .A3(new_n234), .ZN(new_n235));
  NOR2_X1   g034(.A1(new_n221), .A2(new_n209), .ZN(new_n236));
  AND3_X1   g035(.A1(KEYINPUT65), .A2(G169gat), .A3(G176gat), .ZN(new_n237));
  AOI21_X1  g036(.A(KEYINPUT65), .B1(G169gat), .B2(G176gat), .ZN(new_n238));
  NOR2_X1   g037(.A1(new_n237), .A2(new_n238), .ZN(new_n239));
  NOR2_X1   g038(.A1(G169gat), .A2(G176gat), .ZN(new_n240));
  NAND2_X1  g039(.A1(new_n240), .A2(KEYINPUT72), .ZN(new_n241));
  AOI21_X1  g040(.A(new_n239), .B1(KEYINPUT26), .B2(new_n241), .ZN(new_n242));
  OR2_X1    g041(.A1(new_n241), .A2(KEYINPUT26), .ZN(new_n243));
  AOI21_X1  g042(.A(new_n236), .B1(new_n242), .B2(new_n243), .ZN(new_n244));
  NAND3_X1  g043(.A1(new_n226), .A2(new_n235), .A3(new_n244), .ZN(new_n245));
  INV_X1    g044(.A(KEYINPUT25), .ZN(new_n246));
  OR2_X1    g045(.A1(new_n240), .A2(KEYINPUT23), .ZN(new_n247));
  AOI21_X1  g046(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n248));
  XNOR2_X1  g047(.A(new_n248), .B(KEYINPUT64), .ZN(new_n249));
  NAND3_X1  g048(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n250));
  OAI21_X1  g049(.A(new_n250), .B1(G183gat), .B2(G190gat), .ZN(new_n251));
  OAI211_X1 g050(.A(new_n246), .B(new_n247), .C1(new_n249), .C2(new_n251), .ZN(new_n252));
  OR2_X1    g051(.A1(new_n246), .A2(KEYINPUT66), .ZN(new_n253));
  NAND2_X1  g052(.A1(new_n252), .A2(new_n253), .ZN(new_n254));
  NAND2_X1  g053(.A1(new_n240), .A2(KEYINPUT23), .ZN(new_n255));
  OAI21_X1  g054(.A(new_n255), .B1(new_n237), .B2(new_n238), .ZN(new_n256));
  INV_X1    g055(.A(new_n256), .ZN(new_n257));
  NAND2_X1  g056(.A1(new_n256), .A2(KEYINPUT66), .ZN(new_n258));
  OAI22_X1  g057(.A1(new_n207), .A2(G183gat), .B1(KEYINPUT24), .B2(new_n236), .ZN(new_n259));
  XNOR2_X1  g058(.A(new_n250), .B(KEYINPUT67), .ZN(new_n260));
  OAI211_X1 g059(.A(new_n258), .B(new_n247), .C1(new_n259), .C2(new_n260), .ZN(new_n261));
  AOI22_X1  g060(.A1(new_n254), .A2(new_n257), .B1(new_n261), .B2(KEYINPUT25), .ZN(new_n262));
  NAND2_X1  g061(.A1(new_n245), .A2(new_n262), .ZN(new_n263));
  XNOR2_X1  g062(.A(G113gat), .B(G120gat), .ZN(new_n264));
  NAND2_X1  g063(.A1(new_n264), .A2(KEYINPUT75), .ZN(new_n265));
  INV_X1    g064(.A(G134gat), .ZN(new_n266));
  NAND2_X1  g065(.A1(new_n266), .A2(G127gat), .ZN(new_n267));
  INV_X1    g066(.A(G127gat), .ZN(new_n268));
  AOI21_X1  g067(.A(KEYINPUT1), .B1(new_n268), .B2(G134gat), .ZN(new_n269));
  INV_X1    g068(.A(G113gat), .ZN(new_n270));
  OR3_X1    g069(.A1(new_n270), .A2(KEYINPUT75), .A3(G120gat), .ZN(new_n271));
  NAND4_X1  g070(.A1(new_n265), .A2(new_n267), .A3(new_n269), .A4(new_n271), .ZN(new_n272));
  OR2_X1    g071(.A1(KEYINPUT74), .A2(G127gat), .ZN(new_n273));
  NAND2_X1  g072(.A1(KEYINPUT74), .A2(G127gat), .ZN(new_n274));
  AOI21_X1  g073(.A(new_n266), .B1(new_n273), .B2(new_n274), .ZN(new_n275));
  OAI21_X1  g074(.A(KEYINPUT73), .B1(new_n268), .B2(G134gat), .ZN(new_n276));
  INV_X1    g075(.A(KEYINPUT73), .ZN(new_n277));
  NAND3_X1  g076(.A1(new_n277), .A2(new_n266), .A3(G127gat), .ZN(new_n278));
  NAND2_X1  g077(.A1(new_n276), .A2(new_n278), .ZN(new_n279));
  OAI22_X1  g078(.A1(new_n275), .A2(new_n279), .B1(KEYINPUT1), .B2(new_n264), .ZN(new_n280));
  NAND2_X1  g079(.A1(new_n272), .A2(new_n280), .ZN(new_n281));
  NAND2_X1  g080(.A1(new_n263), .A2(new_n281), .ZN(new_n282));
  INV_X1    g081(.A(new_n281), .ZN(new_n283));
  NAND3_X1  g082(.A1(new_n245), .A2(new_n283), .A3(new_n262), .ZN(new_n284));
  NAND2_X1  g083(.A1(new_n282), .A2(new_n284), .ZN(new_n285));
  AND2_X1   g084(.A1(G227gat), .A2(G233gat), .ZN(new_n286));
  AOI21_X1  g085(.A(KEYINPUT76), .B1(new_n285), .B2(new_n286), .ZN(new_n287));
  AND3_X1   g086(.A1(new_n245), .A2(new_n283), .A3(new_n262), .ZN(new_n288));
  AOI21_X1  g087(.A(new_n283), .B1(new_n245), .B2(new_n262), .ZN(new_n289));
  OAI211_X1 g088(.A(KEYINPUT76), .B(new_n286), .C1(new_n288), .C2(new_n289), .ZN(new_n290));
  INV_X1    g089(.A(new_n290), .ZN(new_n291));
  OAI21_X1  g090(.A(KEYINPUT32), .B1(new_n287), .B2(new_n291), .ZN(new_n292));
  NAND2_X1  g091(.A1(new_n292), .A2(KEYINPUT34), .ZN(new_n293));
  INV_X1    g092(.A(KEYINPUT33), .ZN(new_n294));
  OAI21_X1  g093(.A(new_n294), .B1(new_n287), .B2(new_n291), .ZN(new_n295));
  XNOR2_X1  g094(.A(G15gat), .B(G43gat), .ZN(new_n296));
  INV_X1    g095(.A(G71gat), .ZN(new_n297));
  XNOR2_X1  g096(.A(new_n296), .B(new_n297), .ZN(new_n298));
  XOR2_X1   g097(.A(KEYINPUT77), .B(G99gat), .Z(new_n299));
  XOR2_X1   g098(.A(new_n298), .B(new_n299), .Z(new_n300));
  NAND2_X1  g099(.A1(new_n295), .A2(new_n300), .ZN(new_n301));
  OAI21_X1  g100(.A(new_n286), .B1(new_n288), .B2(new_n289), .ZN(new_n302));
  INV_X1    g101(.A(KEYINPUT76), .ZN(new_n303));
  NAND2_X1  g102(.A1(new_n302), .A2(new_n303), .ZN(new_n304));
  NAND2_X1  g103(.A1(new_n304), .A2(new_n290), .ZN(new_n305));
  INV_X1    g104(.A(KEYINPUT34), .ZN(new_n306));
  NAND3_X1  g105(.A1(new_n305), .A2(KEYINPUT32), .A3(new_n306), .ZN(new_n307));
  NAND3_X1  g106(.A1(new_n293), .A2(new_n301), .A3(new_n307), .ZN(new_n308));
  INV_X1    g107(.A(new_n300), .ZN(new_n309));
  AOI21_X1  g108(.A(new_n309), .B1(new_n305), .B2(new_n294), .ZN(new_n310));
  AOI21_X1  g109(.A(new_n306), .B1(new_n305), .B2(KEYINPUT32), .ZN(new_n311));
  INV_X1    g110(.A(KEYINPUT32), .ZN(new_n312));
  AOI211_X1 g111(.A(new_n312), .B(KEYINPUT34), .C1(new_n304), .C2(new_n290), .ZN(new_n313));
  OAI21_X1  g112(.A(new_n310), .B1(new_n311), .B2(new_n313), .ZN(new_n314));
  NOR2_X1   g113(.A1(new_n285), .A2(new_n286), .ZN(new_n315));
  AND3_X1   g114(.A1(new_n308), .A2(new_n314), .A3(new_n315), .ZN(new_n316));
  AOI21_X1  g115(.A(new_n315), .B1(new_n308), .B2(new_n314), .ZN(new_n317));
  NAND2_X1  g116(.A1(G228gat), .A2(G233gat), .ZN(new_n318));
  INV_X1    g117(.A(KEYINPUT3), .ZN(new_n319));
  XNOR2_X1  g118(.A(KEYINPUT78), .B(G197gat), .ZN(new_n320));
  OR2_X1    g119(.A1(new_n320), .A2(G204gat), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n320), .A2(G204gat), .ZN(new_n322));
  AND2_X1   g121(.A1(G211gat), .A2(G218gat), .ZN(new_n323));
  OAI211_X1 g122(.A(new_n321), .B(new_n322), .C1(KEYINPUT22), .C2(new_n323), .ZN(new_n324));
  NOR2_X1   g123(.A1(G211gat), .A2(G218gat), .ZN(new_n325));
  NOR2_X1   g124(.A1(new_n323), .A2(new_n325), .ZN(new_n326));
  INV_X1    g125(.A(new_n326), .ZN(new_n327));
  XNOR2_X1  g126(.A(new_n324), .B(new_n327), .ZN(new_n328));
  OAI21_X1  g127(.A(new_n319), .B1(new_n328), .B2(KEYINPUT29), .ZN(new_n329));
  NAND2_X1  g128(.A1(G155gat), .A2(G162gat), .ZN(new_n330));
  INV_X1    g129(.A(G155gat), .ZN(new_n331));
  INV_X1    g130(.A(G162gat), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n331), .A2(new_n332), .ZN(new_n333));
  OAI21_X1  g132(.A(new_n330), .B1(new_n333), .B2(KEYINPUT2), .ZN(new_n334));
  XOR2_X1   g133(.A(G141gat), .B(G148gat), .Z(new_n335));
  NAND2_X1  g134(.A1(new_n334), .A2(new_n335), .ZN(new_n336));
  NAND2_X1  g135(.A1(new_n336), .A2(KEYINPUT81), .ZN(new_n337));
  INV_X1    g136(.A(KEYINPUT81), .ZN(new_n338));
  NAND3_X1  g137(.A1(new_n334), .A2(new_n335), .A3(new_n338), .ZN(new_n339));
  XNOR2_X1  g138(.A(G141gat), .B(G148gat), .ZN(new_n340));
  OAI211_X1 g139(.A(new_n330), .B(new_n333), .C1(new_n340), .C2(KEYINPUT2), .ZN(new_n341));
  NAND3_X1  g140(.A1(new_n337), .A2(new_n339), .A3(new_n341), .ZN(new_n342));
  NAND2_X1  g141(.A1(new_n329), .A2(new_n342), .ZN(new_n343));
  AOI21_X1  g142(.A(new_n318), .B1(new_n343), .B2(KEYINPUT84), .ZN(new_n344));
  AND3_X1   g143(.A1(new_n334), .A2(new_n335), .A3(new_n338), .ZN(new_n345));
  AOI21_X1  g144(.A(new_n338), .B1(new_n334), .B2(new_n335), .ZN(new_n346));
  NOR2_X1   g145(.A1(new_n345), .A2(new_n346), .ZN(new_n347));
  INV_X1    g146(.A(KEYINPUT82), .ZN(new_n348));
  NAND4_X1  g147(.A1(new_n347), .A2(new_n348), .A3(new_n319), .A4(new_n341), .ZN(new_n349));
  NAND4_X1  g148(.A1(new_n337), .A2(new_n319), .A3(new_n339), .A4(new_n341), .ZN(new_n350));
  NAND2_X1  g149(.A1(new_n350), .A2(KEYINPUT82), .ZN(new_n351));
  AOI21_X1  g150(.A(KEYINPUT29), .B1(new_n349), .B2(new_n351), .ZN(new_n352));
  INV_X1    g151(.A(new_n328), .ZN(new_n353));
  OAI21_X1  g152(.A(new_n343), .B1(new_n352), .B2(new_n353), .ZN(new_n354));
  XNOR2_X1  g153(.A(new_n344), .B(new_n354), .ZN(new_n355));
  XNOR2_X1  g154(.A(G78gat), .B(G106gat), .ZN(new_n356));
  XNOR2_X1  g155(.A(KEYINPUT31), .B(G50gat), .ZN(new_n357));
  XNOR2_X1  g156(.A(new_n356), .B(new_n357), .ZN(new_n358));
  NOR2_X1   g157(.A1(new_n358), .A2(G22gat), .ZN(new_n359));
  INV_X1    g158(.A(G22gat), .ZN(new_n360));
  NOR2_X1   g159(.A1(new_n360), .A2(KEYINPUT85), .ZN(new_n361));
  AOI21_X1  g160(.A(new_n359), .B1(new_n358), .B2(new_n361), .ZN(new_n362));
  XNOR2_X1  g161(.A(new_n355), .B(new_n362), .ZN(new_n363));
  NOR3_X1   g162(.A1(new_n316), .A2(new_n317), .A3(new_n363), .ZN(new_n364));
  AOI21_X1  g163(.A(KEYINPUT29), .B1(new_n245), .B2(new_n262), .ZN(new_n365));
  NAND2_X1  g164(.A1(G226gat), .A2(G233gat), .ZN(new_n366));
  INV_X1    g165(.A(new_n366), .ZN(new_n367));
  OAI21_X1  g166(.A(KEYINPUT79), .B1(new_n365), .B2(new_n367), .ZN(new_n368));
  AOI21_X1  g167(.A(new_n366), .B1(new_n245), .B2(new_n262), .ZN(new_n369));
  INV_X1    g168(.A(KEYINPUT29), .ZN(new_n370));
  NAND2_X1  g169(.A1(new_n263), .A2(new_n370), .ZN(new_n371));
  AOI21_X1  g170(.A(new_n369), .B1(new_n371), .B2(new_n366), .ZN(new_n372));
  OAI211_X1 g171(.A(new_n328), .B(new_n368), .C1(new_n372), .C2(KEYINPUT79), .ZN(new_n373));
  NOR2_X1   g172(.A1(new_n365), .A2(new_n367), .ZN(new_n374));
  OAI21_X1  g173(.A(new_n353), .B1(new_n374), .B2(new_n369), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n373), .A2(new_n375), .ZN(new_n376));
  XNOR2_X1  g175(.A(KEYINPUT80), .B(G64gat), .ZN(new_n377));
  XNOR2_X1  g176(.A(new_n377), .B(G92gat), .ZN(new_n378));
  XNOR2_X1  g177(.A(G8gat), .B(G36gat), .ZN(new_n379));
  XOR2_X1   g178(.A(new_n378), .B(new_n379), .Z(new_n380));
  NAND2_X1  g179(.A1(new_n376), .A2(new_n380), .ZN(new_n381));
  INV_X1    g180(.A(KEYINPUT30), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n381), .A2(new_n382), .ZN(new_n383));
  XNOR2_X1  g182(.A(G1gat), .B(G29gat), .ZN(new_n384));
  INV_X1    g183(.A(G85gat), .ZN(new_n385));
  XNOR2_X1  g184(.A(new_n384), .B(new_n385), .ZN(new_n386));
  XNOR2_X1  g185(.A(KEYINPUT0), .B(G57gat), .ZN(new_n387));
  XOR2_X1   g186(.A(new_n386), .B(new_n387), .Z(new_n388));
  INV_X1    g187(.A(KEYINPUT5), .ZN(new_n389));
  OAI21_X1  g188(.A(KEYINPUT4), .B1(new_n342), .B2(new_n281), .ZN(new_n390));
  NOR3_X1   g189(.A1(new_n342), .A2(new_n281), .A3(KEYINPUT4), .ZN(new_n391));
  INV_X1    g190(.A(KEYINPUT83), .ZN(new_n392));
  OAI21_X1  g191(.A(new_n390), .B1(new_n391), .B2(new_n392), .ZN(new_n393));
  NAND3_X1  g192(.A1(new_n283), .A2(new_n347), .A3(new_n341), .ZN(new_n394));
  NAND3_X1  g193(.A1(new_n394), .A2(KEYINPUT83), .A3(KEYINPUT4), .ZN(new_n395));
  NAND2_X1  g194(.A1(new_n393), .A2(new_n395), .ZN(new_n396));
  NAND2_X1  g195(.A1(G225gat), .A2(G233gat), .ZN(new_n397));
  AOI21_X1  g196(.A(new_n283), .B1(new_n349), .B2(new_n351), .ZN(new_n398));
  NAND2_X1  g197(.A1(new_n342), .A2(KEYINPUT3), .ZN(new_n399));
  NAND2_X1  g198(.A1(new_n398), .A2(new_n399), .ZN(new_n400));
  AND4_X1   g199(.A1(new_n389), .A2(new_n396), .A3(new_n397), .A4(new_n400), .ZN(new_n401));
  NAND2_X1  g200(.A1(new_n342), .A2(new_n281), .ZN(new_n402));
  AOI21_X1  g201(.A(new_n397), .B1(new_n394), .B2(new_n402), .ZN(new_n403));
  OR3_X1    g202(.A1(new_n342), .A2(new_n281), .A3(KEYINPUT4), .ZN(new_n404));
  INV_X1    g203(.A(new_n397), .ZN(new_n405));
  OAI21_X1  g204(.A(new_n404), .B1(new_n390), .B2(new_n405), .ZN(new_n406));
  AOI211_X1 g205(.A(new_n389), .B(new_n403), .C1(new_n400), .C2(new_n406), .ZN(new_n407));
  OAI21_X1  g206(.A(new_n388), .B1(new_n401), .B2(new_n407), .ZN(new_n408));
  AOI22_X1  g207(.A1(new_n393), .A2(new_n395), .B1(new_n398), .B2(new_n399), .ZN(new_n409));
  NAND3_X1  g208(.A1(new_n409), .A2(new_n389), .A3(new_n397), .ZN(new_n410));
  INV_X1    g209(.A(new_n388), .ZN(new_n411));
  NAND2_X1  g210(.A1(new_n400), .A2(new_n406), .ZN(new_n412));
  NAND2_X1  g211(.A1(new_n412), .A2(KEYINPUT5), .ZN(new_n413));
  OAI211_X1 g212(.A(new_n410), .B(new_n411), .C1(new_n413), .C2(new_n403), .ZN(new_n414));
  INV_X1    g213(.A(KEYINPUT6), .ZN(new_n415));
  NAND3_X1  g214(.A1(new_n408), .A2(new_n414), .A3(new_n415), .ZN(new_n416));
  OAI211_X1 g215(.A(KEYINPUT6), .B(new_n388), .C1(new_n401), .C2(new_n407), .ZN(new_n417));
  NAND2_X1  g216(.A1(new_n416), .A2(new_n417), .ZN(new_n418));
  INV_X1    g217(.A(new_n380), .ZN(new_n419));
  NAND3_X1  g218(.A1(new_n373), .A2(new_n375), .A3(new_n419), .ZN(new_n420));
  NAND3_X1  g219(.A1(new_n376), .A2(KEYINPUT30), .A3(new_n380), .ZN(new_n421));
  NAND4_X1  g220(.A1(new_n383), .A2(new_n418), .A3(new_n420), .A4(new_n421), .ZN(new_n422));
  INV_X1    g221(.A(new_n422), .ZN(new_n423));
  INV_X1    g222(.A(KEYINPUT88), .ZN(new_n424));
  OAI211_X1 g223(.A(new_n364), .B(new_n423), .C1(new_n424), .C2(KEYINPUT35), .ZN(new_n425));
  NAND2_X1  g224(.A1(new_n308), .A2(new_n314), .ZN(new_n426));
  INV_X1    g225(.A(new_n315), .ZN(new_n427));
  NAND2_X1  g226(.A1(new_n426), .A2(new_n427), .ZN(new_n428));
  INV_X1    g227(.A(new_n363), .ZN(new_n429));
  NAND3_X1  g228(.A1(new_n308), .A2(new_n314), .A3(new_n315), .ZN(new_n430));
  NAND4_X1  g229(.A1(new_n428), .A2(new_n423), .A3(new_n429), .A4(new_n430), .ZN(new_n431));
  INV_X1    g230(.A(KEYINPUT35), .ZN(new_n432));
  NAND3_X1  g231(.A1(new_n428), .A2(new_n429), .A3(new_n430), .ZN(new_n433));
  OAI211_X1 g232(.A(new_n431), .B(new_n432), .C1(new_n433), .C2(KEYINPUT88), .ZN(new_n434));
  INV_X1    g233(.A(KEYINPUT36), .ZN(new_n435));
  OAI21_X1  g234(.A(new_n435), .B1(new_n316), .B2(new_n317), .ZN(new_n436));
  NAND3_X1  g235(.A1(new_n428), .A2(KEYINPUT36), .A3(new_n430), .ZN(new_n437));
  NAND2_X1  g236(.A1(new_n436), .A2(new_n437), .ZN(new_n438));
  INV_X1    g237(.A(KEYINPUT37), .ZN(new_n439));
  NAND3_X1  g238(.A1(new_n373), .A2(new_n439), .A3(new_n375), .ZN(new_n440));
  OAI211_X1 g239(.A(new_n353), .B(new_n368), .C1(new_n372), .C2(KEYINPUT79), .ZN(new_n441));
  OAI21_X1  g240(.A(new_n441), .B1(new_n353), .B2(new_n372), .ZN(new_n442));
  OAI21_X1  g241(.A(new_n440), .B1(new_n442), .B2(new_n439), .ZN(new_n443));
  NOR2_X1   g242(.A1(new_n380), .A2(KEYINPUT38), .ZN(new_n444));
  AOI21_X1  g243(.A(new_n418), .B1(new_n443), .B2(new_n444), .ZN(new_n445));
  INV_X1    g244(.A(KEYINPUT38), .ZN(new_n446));
  NAND2_X1  g245(.A1(new_n376), .A2(KEYINPUT37), .ZN(new_n447));
  AOI21_X1  g246(.A(new_n380), .B1(new_n447), .B2(new_n440), .ZN(new_n448));
  OAI211_X1 g247(.A(new_n445), .B(new_n381), .C1(new_n446), .C2(new_n448), .ZN(new_n449));
  AOI21_X1  g248(.A(new_n397), .B1(new_n396), .B2(new_n400), .ZN(new_n450));
  INV_X1    g249(.A(KEYINPUT39), .ZN(new_n451));
  AOI21_X1  g250(.A(new_n388), .B1(new_n450), .B2(new_n451), .ZN(new_n452));
  INV_X1    g251(.A(KEYINPUT86), .ZN(new_n453));
  NAND3_X1  g252(.A1(new_n394), .A2(new_n397), .A3(new_n402), .ZN(new_n454));
  OAI211_X1 g253(.A(KEYINPUT39), .B(new_n454), .C1(new_n409), .C2(new_n397), .ZN(new_n455));
  AND3_X1   g254(.A1(new_n452), .A2(new_n453), .A3(new_n455), .ZN(new_n456));
  AOI21_X1  g255(.A(new_n453), .B1(new_n452), .B2(new_n455), .ZN(new_n457));
  NOR3_X1   g256(.A1(new_n456), .A2(new_n457), .A3(KEYINPUT40), .ZN(new_n458));
  NAND3_X1  g257(.A1(new_n452), .A2(KEYINPUT40), .A3(new_n455), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n459), .A2(KEYINPUT87), .ZN(new_n460));
  INV_X1    g259(.A(KEYINPUT87), .ZN(new_n461));
  NAND4_X1  g260(.A1(new_n452), .A2(new_n461), .A3(KEYINPUT40), .A4(new_n455), .ZN(new_n462));
  NAND2_X1  g261(.A1(new_n460), .A2(new_n462), .ZN(new_n463));
  NOR2_X1   g262(.A1(new_n458), .A2(new_n463), .ZN(new_n464));
  NAND3_X1  g263(.A1(new_n383), .A2(new_n420), .A3(new_n421), .ZN(new_n465));
  NAND3_X1  g264(.A1(new_n464), .A2(new_n465), .A3(new_n408), .ZN(new_n466));
  NAND3_X1  g265(.A1(new_n449), .A2(new_n429), .A3(new_n466), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n438), .A2(new_n467), .ZN(new_n468));
  NOR2_X1   g267(.A1(new_n423), .A2(new_n429), .ZN(new_n469));
  OAI211_X1 g268(.A(new_n425), .B(new_n434), .C1(new_n468), .C2(new_n469), .ZN(new_n470));
  INV_X1    g269(.A(KEYINPUT89), .ZN(new_n471));
  NAND2_X1  g270(.A1(new_n471), .A2(KEYINPUT14), .ZN(new_n472));
  INV_X1    g271(.A(KEYINPUT14), .ZN(new_n473));
  NAND2_X1  g272(.A1(new_n473), .A2(KEYINPUT89), .ZN(new_n474));
  OAI211_X1 g273(.A(new_n472), .B(new_n474), .C1(G29gat), .C2(G36gat), .ZN(new_n475));
  INV_X1    g274(.A(G29gat), .ZN(new_n476));
  INV_X1    g275(.A(G36gat), .ZN(new_n477));
  NAND4_X1  g276(.A1(new_n471), .A2(new_n476), .A3(new_n477), .A4(KEYINPUT14), .ZN(new_n478));
  OAI211_X1 g277(.A(new_n475), .B(new_n478), .C1(new_n476), .C2(new_n477), .ZN(new_n479));
  INV_X1    g278(.A(G43gat), .ZN(new_n480));
  NAND2_X1  g279(.A1(new_n480), .A2(G50gat), .ZN(new_n481));
  INV_X1    g280(.A(G50gat), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n482), .A2(G43gat), .ZN(new_n483));
  NAND3_X1  g282(.A1(new_n481), .A2(new_n483), .A3(KEYINPUT15), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n479), .A2(new_n484), .ZN(new_n485));
  INV_X1    g284(.A(KEYINPUT91), .ZN(new_n486));
  OAI21_X1  g285(.A(new_n486), .B1(new_n480), .B2(G50gat), .ZN(new_n487));
  NAND3_X1  g286(.A1(new_n482), .A2(KEYINPUT91), .A3(G43gat), .ZN(new_n488));
  NAND3_X1  g287(.A1(new_n487), .A2(new_n481), .A3(new_n488), .ZN(new_n489));
  XOR2_X1   g288(.A(KEYINPUT90), .B(KEYINPUT15), .Z(new_n490));
  NAND2_X1  g289(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  AND2_X1   g290(.A1(new_n491), .A2(new_n484), .ZN(new_n492));
  OAI21_X1  g291(.A(new_n485), .B1(new_n492), .B2(new_n479), .ZN(new_n493));
  NAND2_X1  g292(.A1(new_n493), .A2(KEYINPUT17), .ZN(new_n494));
  XNOR2_X1  g293(.A(G15gat), .B(G22gat), .ZN(new_n495));
  INV_X1    g294(.A(G1gat), .ZN(new_n496));
  NAND2_X1  g295(.A1(new_n496), .A2(KEYINPUT16), .ZN(new_n497));
  NAND2_X1  g296(.A1(new_n495), .A2(new_n497), .ZN(new_n498));
  OAI21_X1  g297(.A(new_n498), .B1(G1gat), .B2(new_n495), .ZN(new_n499));
  INV_X1    g298(.A(G8gat), .ZN(new_n500));
  XNOR2_X1  g299(.A(new_n499), .B(new_n500), .ZN(new_n501));
  INV_X1    g300(.A(KEYINPUT17), .ZN(new_n502));
  OAI211_X1 g301(.A(new_n502), .B(new_n485), .C1(new_n492), .C2(new_n479), .ZN(new_n503));
  NAND3_X1  g302(.A1(new_n494), .A2(new_n501), .A3(new_n503), .ZN(new_n504));
  OR2_X1    g303(.A1(new_n501), .A2(new_n493), .ZN(new_n505));
  NAND2_X1  g304(.A1(G229gat), .A2(G233gat), .ZN(new_n506));
  NAND3_X1  g305(.A1(new_n504), .A2(new_n505), .A3(new_n506), .ZN(new_n507));
  INV_X1    g306(.A(KEYINPUT18), .ZN(new_n508));
  NAND2_X1  g307(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n501), .A2(new_n493), .ZN(new_n510));
  NAND2_X1  g309(.A1(new_n505), .A2(new_n510), .ZN(new_n511));
  XNOR2_X1  g310(.A(new_n506), .B(KEYINPUT13), .ZN(new_n512));
  INV_X1    g311(.A(new_n512), .ZN(new_n513));
  NAND2_X1  g312(.A1(new_n511), .A2(new_n513), .ZN(new_n514));
  NAND4_X1  g313(.A1(new_n504), .A2(KEYINPUT18), .A3(new_n505), .A4(new_n506), .ZN(new_n515));
  NAND3_X1  g314(.A1(new_n509), .A2(new_n514), .A3(new_n515), .ZN(new_n516));
  XOR2_X1   g315(.A(G113gat), .B(G141gat), .Z(new_n517));
  XNOR2_X1  g316(.A(new_n517), .B(G197gat), .ZN(new_n518));
  XNOR2_X1  g317(.A(KEYINPUT11), .B(G169gat), .ZN(new_n519));
  XNOR2_X1  g318(.A(new_n518), .B(new_n519), .ZN(new_n520));
  XOR2_X1   g319(.A(new_n520), .B(KEYINPUT12), .Z(new_n521));
  NAND2_X1  g320(.A1(new_n516), .A2(new_n521), .ZN(new_n522));
  INV_X1    g321(.A(new_n521), .ZN(new_n523));
  NAND4_X1  g322(.A1(new_n523), .A2(new_n509), .A3(new_n514), .A4(new_n515), .ZN(new_n524));
  NAND2_X1  g323(.A1(new_n522), .A2(new_n524), .ZN(new_n525));
  AND2_X1   g324(.A1(new_n470), .A2(new_n525), .ZN(new_n526));
  INV_X1    g325(.A(KEYINPUT21), .ZN(new_n527));
  INV_X1    g326(.A(KEYINPUT92), .ZN(new_n528));
  XNOR2_X1  g327(.A(G57gat), .B(G64gat), .ZN(new_n529));
  AOI21_X1  g328(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n530));
  OAI21_X1  g329(.A(new_n528), .B1(new_n529), .B2(new_n530), .ZN(new_n531));
  XNOR2_X1  g330(.A(G71gat), .B(G78gat), .ZN(new_n532));
  XNOR2_X1  g331(.A(new_n531), .B(new_n532), .ZN(new_n533));
  OAI21_X1  g332(.A(new_n501), .B1(new_n527), .B2(new_n533), .ZN(new_n534));
  XNOR2_X1  g333(.A(new_n534), .B(new_n221), .ZN(new_n535));
  XNOR2_X1  g334(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n536));
  XNOR2_X1  g335(.A(new_n535), .B(new_n536), .ZN(new_n537));
  NAND2_X1  g336(.A1(G231gat), .A2(G233gat), .ZN(new_n538));
  INV_X1    g337(.A(G211gat), .ZN(new_n539));
  XNOR2_X1  g338(.A(new_n538), .B(new_n539), .ZN(new_n540));
  OR2_X1    g339(.A1(new_n537), .A2(new_n540), .ZN(new_n541));
  XOR2_X1   g340(.A(KEYINPUT93), .B(KEYINPUT21), .Z(new_n542));
  NAND2_X1  g341(.A1(new_n533), .A2(new_n542), .ZN(new_n543));
  XNOR2_X1  g342(.A(G127gat), .B(G155gat), .ZN(new_n544));
  XNOR2_X1  g343(.A(new_n543), .B(new_n544), .ZN(new_n545));
  NAND2_X1  g344(.A1(new_n537), .A2(new_n540), .ZN(new_n546));
  AND3_X1   g345(.A1(new_n541), .A2(new_n545), .A3(new_n546), .ZN(new_n547));
  AOI21_X1  g346(.A(new_n545), .B1(new_n541), .B2(new_n546), .ZN(new_n548));
  NOR2_X1   g347(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  INV_X1    g348(.A(KEYINPUT95), .ZN(new_n550));
  INV_X1    g349(.A(KEYINPUT7), .ZN(new_n551));
  NAND2_X1  g350(.A1(new_n550), .A2(new_n551), .ZN(new_n552));
  NAND2_X1  g351(.A1(KEYINPUT95), .A2(KEYINPUT7), .ZN(new_n553));
  NAND4_X1  g352(.A1(new_n552), .A2(G85gat), .A3(G92gat), .A4(new_n553), .ZN(new_n554));
  NOR2_X1   g353(.A1(KEYINPUT95), .A2(KEYINPUT7), .ZN(new_n555));
  NAND2_X1  g354(.A1(G85gat), .A2(G92gat), .ZN(new_n556));
  NAND2_X1  g355(.A1(G99gat), .A2(G106gat), .ZN(new_n557));
  AOI22_X1  g356(.A1(new_n555), .A2(new_n556), .B1(new_n557), .B2(KEYINPUT8), .ZN(new_n558));
  OAI211_X1 g357(.A(new_n554), .B(new_n558), .C1(G85gat), .C2(G92gat), .ZN(new_n559));
  XOR2_X1   g358(.A(G99gat), .B(G106gat), .Z(new_n560));
  XNOR2_X1  g359(.A(new_n559), .B(new_n560), .ZN(new_n561));
  AND3_X1   g360(.A1(new_n494), .A2(new_n503), .A3(new_n561), .ZN(new_n562));
  NAND2_X1  g361(.A1(G232gat), .A2(G233gat), .ZN(new_n563));
  INV_X1    g362(.A(new_n563), .ZN(new_n564));
  NAND2_X1  g363(.A1(new_n564), .A2(KEYINPUT41), .ZN(new_n565));
  OAI21_X1  g364(.A(new_n565), .B1(new_n561), .B2(new_n493), .ZN(new_n566));
  NOR2_X1   g365(.A1(new_n562), .A2(new_n566), .ZN(new_n567));
  XOR2_X1   g366(.A(G190gat), .B(G218gat), .Z(new_n568));
  NOR2_X1   g367(.A1(new_n567), .A2(new_n568), .ZN(new_n569));
  INV_X1    g368(.A(new_n569), .ZN(new_n570));
  NAND2_X1  g369(.A1(new_n567), .A2(new_n568), .ZN(new_n571));
  NOR2_X1   g370(.A1(new_n564), .A2(KEYINPUT41), .ZN(new_n572));
  XNOR2_X1  g371(.A(new_n572), .B(KEYINPUT94), .ZN(new_n573));
  XNOR2_X1  g372(.A(new_n573), .B(new_n266), .ZN(new_n574));
  XNOR2_X1  g373(.A(new_n574), .B(new_n332), .ZN(new_n575));
  NAND4_X1  g374(.A1(new_n570), .A2(KEYINPUT96), .A3(new_n571), .A4(new_n575), .ZN(new_n576));
  INV_X1    g375(.A(new_n571), .ZN(new_n577));
  AOI21_X1  g376(.A(KEYINPUT96), .B1(new_n567), .B2(new_n568), .ZN(new_n578));
  INV_X1    g377(.A(new_n575), .ZN(new_n579));
  OAI22_X1  g378(.A1(new_n577), .A2(new_n569), .B1(new_n578), .B2(new_n579), .ZN(new_n580));
  NAND2_X1  g379(.A1(new_n576), .A2(new_n580), .ZN(new_n581));
  NAND2_X1  g380(.A1(G230gat), .A2(G233gat), .ZN(new_n582));
  INV_X1    g381(.A(new_n582), .ZN(new_n583));
  NAND2_X1  g382(.A1(new_n561), .A2(new_n533), .ZN(new_n584));
  INV_X1    g383(.A(new_n560), .ZN(new_n585));
  XNOR2_X1  g384(.A(new_n559), .B(new_n585), .ZN(new_n586));
  XOR2_X1   g385(.A(new_n531), .B(new_n532), .Z(new_n587));
  NAND2_X1  g386(.A1(new_n586), .A2(new_n587), .ZN(new_n588));
  INV_X1    g387(.A(KEYINPUT10), .ZN(new_n589));
  NAND3_X1  g388(.A1(new_n584), .A2(new_n588), .A3(new_n589), .ZN(new_n590));
  NAND3_X1  g389(.A1(new_n586), .A2(new_n587), .A3(KEYINPUT10), .ZN(new_n591));
  AOI21_X1  g390(.A(new_n583), .B1(new_n590), .B2(new_n591), .ZN(new_n592));
  AOI21_X1  g391(.A(new_n582), .B1(new_n584), .B2(new_n588), .ZN(new_n593));
  OR2_X1    g392(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  XNOR2_X1  g393(.A(G120gat), .B(G148gat), .ZN(new_n595));
  XNOR2_X1  g394(.A(new_n595), .B(KEYINPUT97), .ZN(new_n596));
  XNOR2_X1  g395(.A(G176gat), .B(G204gat), .ZN(new_n597));
  XOR2_X1   g396(.A(new_n596), .B(new_n597), .Z(new_n598));
  INV_X1    g397(.A(new_n598), .ZN(new_n599));
  XNOR2_X1  g398(.A(new_n594), .B(new_n599), .ZN(new_n600));
  INV_X1    g399(.A(new_n600), .ZN(new_n601));
  NOR3_X1   g400(.A1(new_n549), .A2(new_n581), .A3(new_n601), .ZN(new_n602));
  AND2_X1   g401(.A1(new_n526), .A2(new_n602), .ZN(new_n603));
  INV_X1    g402(.A(new_n418), .ZN(new_n604));
  NAND2_X1  g403(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  XNOR2_X1  g404(.A(KEYINPUT98), .B(G1gat), .ZN(new_n606));
  XNOR2_X1  g405(.A(new_n605), .B(new_n606), .ZN(G1324gat));
  NAND2_X1  g406(.A1(new_n603), .A2(new_n465), .ZN(new_n608));
  NOR2_X1   g407(.A1(KEYINPUT100), .A2(KEYINPUT42), .ZN(new_n609));
  XNOR2_X1  g408(.A(KEYINPUT99), .B(KEYINPUT16), .ZN(new_n610));
  XNOR2_X1  g409(.A(new_n610), .B(new_n500), .ZN(new_n611));
  OR3_X1    g410(.A1(new_n608), .A2(new_n609), .A3(new_n611), .ZN(new_n612));
  AND2_X1   g411(.A1(KEYINPUT100), .A2(KEYINPUT42), .ZN(new_n613));
  OAI22_X1  g412(.A1(new_n608), .A2(new_n611), .B1(new_n609), .B2(new_n613), .ZN(new_n614));
  AOI211_X1 g413(.A(KEYINPUT101), .B(new_n500), .C1(new_n603), .C2(new_n465), .ZN(new_n615));
  INV_X1    g414(.A(KEYINPUT101), .ZN(new_n616));
  AOI21_X1  g415(.A(new_n616), .B1(new_n608), .B2(G8gat), .ZN(new_n617));
  OAI211_X1 g416(.A(new_n612), .B(new_n614), .C1(new_n615), .C2(new_n617), .ZN(G1325gat));
  NOR2_X1   g417(.A1(new_n316), .A2(new_n317), .ZN(new_n619));
  NAND2_X1  g418(.A1(new_n603), .A2(new_n619), .ZN(new_n620));
  INV_X1    g419(.A(G15gat), .ZN(new_n621));
  NAND2_X1  g420(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  NAND2_X1  g421(.A1(new_n622), .A2(KEYINPUT102), .ZN(new_n623));
  INV_X1    g422(.A(KEYINPUT102), .ZN(new_n624));
  NAND3_X1  g423(.A1(new_n620), .A2(new_n624), .A3(new_n621), .ZN(new_n625));
  NOR2_X1   g424(.A1(new_n438), .A2(new_n621), .ZN(new_n626));
  AOI22_X1  g425(.A1(new_n623), .A2(new_n625), .B1(new_n603), .B2(new_n626), .ZN(G1326gat));
  NAND2_X1  g426(.A1(new_n603), .A2(new_n363), .ZN(new_n628));
  XNOR2_X1  g427(.A(KEYINPUT43), .B(G22gat), .ZN(new_n629));
  XNOR2_X1  g428(.A(new_n628), .B(new_n629), .ZN(G1327gat));
  INV_X1    g429(.A(new_n549), .ZN(new_n631));
  INV_X1    g430(.A(new_n581), .ZN(new_n632));
  NOR3_X1   g431(.A1(new_n631), .A2(new_n632), .A3(new_n601), .ZN(new_n633));
  NAND2_X1  g432(.A1(new_n526), .A2(new_n633), .ZN(new_n634));
  NOR3_X1   g433(.A1(new_n634), .A2(G29gat), .A3(new_n418), .ZN(new_n635));
  XNOR2_X1  g434(.A(KEYINPUT103), .B(KEYINPUT45), .ZN(new_n636));
  XNOR2_X1  g435(.A(new_n635), .B(new_n636), .ZN(new_n637));
  AND3_X1   g436(.A1(new_n422), .A2(KEYINPUT105), .A3(new_n363), .ZN(new_n638));
  AOI21_X1  g437(.A(KEYINPUT105), .B1(new_n422), .B2(new_n363), .ZN(new_n639));
  NOR2_X1   g438(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  NAND3_X1  g439(.A1(new_n438), .A2(new_n640), .A3(new_n467), .ZN(new_n641));
  NAND3_X1  g440(.A1(new_n641), .A2(new_n425), .A3(new_n434), .ZN(new_n642));
  NAND2_X1  g441(.A1(new_n642), .A2(new_n581), .ZN(new_n643));
  INV_X1    g442(.A(KEYINPUT44), .ZN(new_n644));
  NAND2_X1  g443(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  NOR2_X1   g444(.A1(new_n631), .A2(new_n601), .ZN(new_n646));
  NAND3_X1  g445(.A1(new_n470), .A2(KEYINPUT44), .A3(new_n581), .ZN(new_n647));
  AND3_X1   g446(.A1(new_n522), .A2(KEYINPUT104), .A3(new_n524), .ZN(new_n648));
  AOI21_X1  g447(.A(KEYINPUT104), .B1(new_n522), .B2(new_n524), .ZN(new_n649));
  NOR2_X1   g448(.A1(new_n648), .A2(new_n649), .ZN(new_n650));
  NAND4_X1  g449(.A1(new_n645), .A2(new_n646), .A3(new_n647), .A4(new_n650), .ZN(new_n651));
  OAI21_X1  g450(.A(G29gat), .B1(new_n651), .B2(new_n418), .ZN(new_n652));
  NAND2_X1  g451(.A1(new_n637), .A2(new_n652), .ZN(G1328gat));
  INV_X1    g452(.A(new_n465), .ZN(new_n654));
  NOR2_X1   g453(.A1(new_n654), .A2(G36gat), .ZN(new_n655));
  NAND3_X1  g454(.A1(new_n526), .A2(new_n633), .A3(new_n655), .ZN(new_n656));
  NOR2_X1   g455(.A1(new_n656), .A2(KEYINPUT46), .ZN(new_n657));
  INV_X1    g456(.A(KEYINPUT106), .ZN(new_n658));
  XNOR2_X1  g457(.A(new_n657), .B(new_n658), .ZN(new_n659));
  OR2_X1    g458(.A1(new_n651), .A2(new_n654), .ZN(new_n660));
  AOI21_X1  g459(.A(KEYINPUT46), .B1(new_n660), .B2(G36gat), .ZN(new_n661));
  INV_X1    g460(.A(new_n656), .ZN(new_n662));
  OAI21_X1  g461(.A(new_n659), .B1(new_n661), .B2(new_n662), .ZN(G1329gat));
  INV_X1    g462(.A(KEYINPUT47), .ZN(new_n664));
  INV_X1    g463(.A(new_n619), .ZN(new_n665));
  OAI21_X1  g464(.A(new_n480), .B1(new_n634), .B2(new_n665), .ZN(new_n666));
  OR2_X1    g465(.A1(new_n651), .A2(new_n480), .ZN(new_n667));
  OAI211_X1 g466(.A(new_n664), .B(new_n666), .C1(new_n667), .C2(new_n438), .ZN(new_n668));
  NOR3_X1   g467(.A1(new_n651), .A2(new_n480), .A3(new_n438), .ZN(new_n669));
  INV_X1    g468(.A(new_n666), .ZN(new_n670));
  OAI21_X1  g469(.A(KEYINPUT47), .B1(new_n669), .B2(new_n670), .ZN(new_n671));
  NAND2_X1  g470(.A1(new_n668), .A2(new_n671), .ZN(G1330gat));
  OAI21_X1  g471(.A(G50gat), .B1(new_n651), .B2(new_n429), .ZN(new_n673));
  NAND4_X1  g472(.A1(new_n526), .A2(new_n482), .A3(new_n363), .A4(new_n633), .ZN(new_n674));
  NAND2_X1  g473(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  XOR2_X1   g474(.A(KEYINPUT107), .B(KEYINPUT48), .Z(new_n676));
  NAND2_X1  g475(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  INV_X1    g476(.A(new_n676), .ZN(new_n678));
  NAND3_X1  g477(.A1(new_n673), .A2(new_n678), .A3(new_n674), .ZN(new_n679));
  NAND2_X1  g478(.A1(new_n677), .A2(new_n679), .ZN(G1331gat));
  AND2_X1   g479(.A1(new_n642), .A2(new_n601), .ZN(new_n681));
  NOR3_X1   g480(.A1(new_n549), .A2(new_n581), .A3(new_n650), .ZN(new_n682));
  AND2_X1   g481(.A1(new_n681), .A2(new_n682), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n683), .A2(new_n604), .ZN(new_n684));
  XNOR2_X1  g483(.A(new_n684), .B(G57gat), .ZN(G1332gat));
  AND3_X1   g484(.A1(new_n681), .A2(new_n465), .A3(new_n682), .ZN(new_n686));
  INV_X1    g485(.A(KEYINPUT108), .ZN(new_n687));
  NAND2_X1  g486(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n688));
  NAND3_X1  g487(.A1(new_n686), .A2(new_n687), .A3(new_n688), .ZN(new_n689));
  INV_X1    g488(.A(new_n689), .ZN(new_n690));
  AOI21_X1  g489(.A(new_n687), .B1(new_n686), .B2(new_n688), .ZN(new_n691));
  OAI22_X1  g490(.A1(new_n690), .A2(new_n691), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n692));
  INV_X1    g491(.A(new_n691), .ZN(new_n693));
  NOR2_X1   g492(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n694));
  NAND3_X1  g493(.A1(new_n693), .A2(new_n689), .A3(new_n694), .ZN(new_n695));
  NAND2_X1  g494(.A1(new_n692), .A2(new_n695), .ZN(G1333gat));
  NAND2_X1  g495(.A1(new_n683), .A2(new_n619), .ZN(new_n697));
  NAND2_X1  g496(.A1(new_n697), .A2(new_n297), .ZN(new_n698));
  NAND4_X1  g497(.A1(new_n683), .A2(G71gat), .A3(new_n437), .A4(new_n436), .ZN(new_n699));
  NAND2_X1  g498(.A1(new_n698), .A2(new_n699), .ZN(new_n700));
  NAND2_X1  g499(.A1(new_n700), .A2(KEYINPUT50), .ZN(new_n701));
  INV_X1    g500(.A(KEYINPUT50), .ZN(new_n702));
  NAND3_X1  g501(.A1(new_n698), .A2(new_n702), .A3(new_n699), .ZN(new_n703));
  NAND2_X1  g502(.A1(new_n701), .A2(new_n703), .ZN(G1334gat));
  NAND2_X1  g503(.A1(new_n683), .A2(new_n363), .ZN(new_n705));
  XNOR2_X1  g504(.A(KEYINPUT109), .B(G78gat), .ZN(new_n706));
  XNOR2_X1  g505(.A(new_n705), .B(new_n706), .ZN(G1335gat));
  NOR2_X1   g506(.A1(new_n631), .A2(new_n650), .ZN(new_n708));
  NAND4_X1  g507(.A1(new_n645), .A2(new_n601), .A3(new_n647), .A4(new_n708), .ZN(new_n709));
  NOR3_X1   g508(.A1(new_n709), .A2(new_n385), .A3(new_n418), .ZN(new_n710));
  INV_X1    g509(.A(new_n710), .ZN(new_n711));
  INV_X1    g510(.A(KEYINPUT110), .ZN(new_n712));
  NAND3_X1  g511(.A1(new_n642), .A2(new_n581), .A3(new_n708), .ZN(new_n713));
  NAND2_X1  g512(.A1(new_n713), .A2(KEYINPUT51), .ZN(new_n714));
  INV_X1    g513(.A(KEYINPUT51), .ZN(new_n715));
  NAND4_X1  g514(.A1(new_n642), .A2(new_n715), .A3(new_n581), .A4(new_n708), .ZN(new_n716));
  NAND4_X1  g515(.A1(new_n714), .A2(new_n604), .A3(new_n601), .A4(new_n716), .ZN(new_n717));
  NAND2_X1  g516(.A1(new_n717), .A2(new_n385), .ZN(new_n718));
  NAND3_X1  g517(.A1(new_n711), .A2(new_n712), .A3(new_n718), .ZN(new_n719));
  INV_X1    g518(.A(new_n718), .ZN(new_n720));
  OAI21_X1  g519(.A(KEYINPUT110), .B1(new_n720), .B2(new_n710), .ZN(new_n721));
  NAND2_X1  g520(.A1(new_n719), .A2(new_n721), .ZN(G1336gat));
  OAI21_X1  g521(.A(G92gat), .B1(new_n709), .B2(new_n654), .ZN(new_n723));
  NAND4_X1  g522(.A1(new_n714), .A2(new_n465), .A3(new_n601), .A4(new_n716), .ZN(new_n724));
  OAI21_X1  g523(.A(new_n723), .B1(G92gat), .B2(new_n724), .ZN(new_n725));
  NAND2_X1  g524(.A1(new_n725), .A2(KEYINPUT52), .ZN(new_n726));
  INV_X1    g525(.A(KEYINPUT52), .ZN(new_n727));
  OAI211_X1 g526(.A(new_n723), .B(new_n727), .C1(G92gat), .C2(new_n724), .ZN(new_n728));
  NAND2_X1  g527(.A1(new_n726), .A2(new_n728), .ZN(G1337gat));
  XNOR2_X1  g528(.A(KEYINPUT111), .B(G99gat), .ZN(new_n730));
  OAI21_X1  g529(.A(new_n730), .B1(new_n709), .B2(new_n438), .ZN(new_n731));
  AND2_X1   g530(.A1(new_n714), .A2(new_n716), .ZN(new_n732));
  INV_X1    g531(.A(new_n730), .ZN(new_n733));
  NAND3_X1  g532(.A1(new_n732), .A2(new_n601), .A3(new_n733), .ZN(new_n734));
  OAI21_X1  g533(.A(new_n731), .B1(new_n734), .B2(new_n665), .ZN(G1338gat));
  INV_X1    g534(.A(G106gat), .ZN(new_n736));
  NAND4_X1  g535(.A1(new_n732), .A2(new_n736), .A3(new_n363), .A4(new_n601), .ZN(new_n737));
  XNOR2_X1  g536(.A(KEYINPUT112), .B(KEYINPUT53), .ZN(new_n738));
  OAI21_X1  g537(.A(G106gat), .B1(new_n709), .B2(new_n429), .ZN(new_n739));
  AND3_X1   g538(.A1(new_n737), .A2(new_n738), .A3(new_n739), .ZN(new_n740));
  AOI21_X1  g539(.A(new_n738), .B1(new_n737), .B2(new_n739), .ZN(new_n741));
  NOR2_X1   g540(.A1(new_n740), .A2(new_n741), .ZN(G1339gat));
  NOR2_X1   g541(.A1(new_n594), .A2(new_n598), .ZN(new_n743));
  NAND3_X1  g542(.A1(new_n590), .A2(new_n591), .A3(new_n583), .ZN(new_n744));
  INV_X1    g543(.A(KEYINPUT113), .ZN(new_n745));
  NAND2_X1  g544(.A1(new_n744), .A2(new_n745), .ZN(new_n746));
  NAND2_X1  g545(.A1(new_n590), .A2(new_n591), .ZN(new_n747));
  NAND2_X1  g546(.A1(new_n747), .A2(new_n582), .ZN(new_n748));
  NAND4_X1  g547(.A1(new_n590), .A2(new_n591), .A3(KEYINPUT113), .A4(new_n583), .ZN(new_n749));
  NAND4_X1  g548(.A1(new_n746), .A2(new_n748), .A3(KEYINPUT54), .A4(new_n749), .ZN(new_n750));
  INV_X1    g549(.A(KEYINPUT54), .ZN(new_n751));
  AOI21_X1  g550(.A(new_n599), .B1(new_n592), .B2(new_n751), .ZN(new_n752));
  NAND2_X1  g551(.A1(new_n750), .A2(new_n752), .ZN(new_n753));
  INV_X1    g552(.A(KEYINPUT55), .ZN(new_n754));
  AOI21_X1  g553(.A(new_n743), .B1(new_n753), .B2(new_n754), .ZN(new_n755));
  NAND3_X1  g554(.A1(new_n750), .A2(KEYINPUT55), .A3(new_n752), .ZN(new_n756));
  NAND2_X1  g555(.A1(new_n756), .A2(KEYINPUT114), .ZN(new_n757));
  INV_X1    g556(.A(KEYINPUT114), .ZN(new_n758));
  NAND4_X1  g557(.A1(new_n750), .A2(new_n758), .A3(KEYINPUT55), .A4(new_n752), .ZN(new_n759));
  OAI21_X1  g558(.A(KEYINPUT115), .B1(new_n511), .B2(new_n513), .ZN(new_n760));
  INV_X1    g559(.A(KEYINPUT115), .ZN(new_n761));
  NAND4_X1  g560(.A1(new_n505), .A2(new_n761), .A3(new_n510), .A4(new_n512), .ZN(new_n762));
  NAND2_X1  g561(.A1(new_n760), .A2(new_n762), .ZN(new_n763));
  AOI21_X1  g562(.A(new_n506), .B1(new_n504), .B2(new_n505), .ZN(new_n764));
  OAI21_X1  g563(.A(new_n520), .B1(new_n763), .B2(new_n764), .ZN(new_n765));
  NAND3_X1  g564(.A1(new_n765), .A2(KEYINPUT116), .A3(new_n524), .ZN(new_n766));
  AND4_X1   g565(.A1(new_n755), .A2(new_n757), .A3(new_n759), .A4(new_n766), .ZN(new_n767));
  NAND2_X1  g566(.A1(new_n765), .A2(new_n524), .ZN(new_n768));
  INV_X1    g567(.A(KEYINPUT116), .ZN(new_n769));
  NAND2_X1  g568(.A1(new_n768), .A2(new_n769), .ZN(new_n770));
  NAND2_X1  g569(.A1(new_n770), .A2(new_n581), .ZN(new_n771));
  INV_X1    g570(.A(new_n771), .ZN(new_n772));
  AOI21_X1  g571(.A(KEYINPUT117), .B1(new_n767), .B2(new_n772), .ZN(new_n773));
  NAND4_X1  g572(.A1(new_n755), .A2(new_n757), .A3(new_n759), .A4(new_n766), .ZN(new_n774));
  INV_X1    g573(.A(KEYINPUT117), .ZN(new_n775));
  NOR3_X1   g574(.A1(new_n774), .A2(new_n771), .A3(new_n775), .ZN(new_n776));
  NOR2_X1   g575(.A1(new_n600), .A2(new_n768), .ZN(new_n777));
  AND3_X1   g576(.A1(new_n755), .A2(new_n757), .A3(new_n759), .ZN(new_n778));
  AOI21_X1  g577(.A(new_n777), .B1(new_n778), .B2(new_n650), .ZN(new_n779));
  OAI22_X1  g578(.A1(new_n773), .A2(new_n776), .B1(new_n779), .B2(new_n581), .ZN(new_n780));
  NAND2_X1  g579(.A1(new_n780), .A2(new_n549), .ZN(new_n781));
  NAND2_X1  g580(.A1(new_n682), .A2(new_n600), .ZN(new_n782));
  AOI21_X1  g581(.A(new_n433), .B1(new_n781), .B2(new_n782), .ZN(new_n783));
  NOR2_X1   g582(.A1(new_n465), .A2(new_n418), .ZN(new_n784));
  NAND2_X1  g583(.A1(new_n783), .A2(new_n784), .ZN(new_n785));
  INV_X1    g584(.A(new_n525), .ZN(new_n786));
  OAI21_X1  g585(.A(G113gat), .B1(new_n785), .B2(new_n786), .ZN(new_n787));
  NAND2_X1  g586(.A1(new_n650), .A2(new_n270), .ZN(new_n788));
  OAI21_X1  g587(.A(new_n787), .B1(new_n785), .B2(new_n788), .ZN(G1340gat));
  INV_X1    g588(.A(new_n785), .ZN(new_n790));
  NAND2_X1  g589(.A1(new_n790), .A2(new_n601), .ZN(new_n791));
  XNOR2_X1  g590(.A(new_n791), .B(G120gat), .ZN(G1341gat));
  NOR2_X1   g591(.A1(new_n785), .A2(new_n549), .ZN(new_n793));
  NAND2_X1  g592(.A1(new_n273), .A2(new_n274), .ZN(new_n794));
  XNOR2_X1  g593(.A(new_n793), .B(new_n794), .ZN(G1342gat));
  NAND2_X1  g594(.A1(new_n790), .A2(new_n581), .ZN(new_n796));
  NOR2_X1   g595(.A1(new_n796), .A2(G134gat), .ZN(new_n797));
  XNOR2_X1  g596(.A(new_n797), .B(KEYINPUT56), .ZN(new_n798));
  NAND2_X1  g597(.A1(new_n796), .A2(G134gat), .ZN(new_n799));
  NAND2_X1  g598(.A1(new_n798), .A2(new_n799), .ZN(G1343gat));
  AOI21_X1  g599(.A(new_n429), .B1(new_n781), .B2(new_n782), .ZN(new_n801));
  OAI21_X1  g600(.A(KEYINPUT119), .B1(new_n801), .B2(KEYINPUT57), .ZN(new_n802));
  AND2_X1   g601(.A1(new_n778), .A2(new_n650), .ZN(new_n803));
  OAI21_X1  g602(.A(new_n632), .B1(new_n803), .B2(new_n777), .ZN(new_n804));
  NAND3_X1  g603(.A1(new_n767), .A2(new_n772), .A3(KEYINPUT117), .ZN(new_n805));
  OAI21_X1  g604(.A(new_n775), .B1(new_n774), .B2(new_n771), .ZN(new_n806));
  NAND2_X1  g605(.A1(new_n805), .A2(new_n806), .ZN(new_n807));
  AOI21_X1  g606(.A(new_n631), .B1(new_n804), .B2(new_n807), .ZN(new_n808));
  INV_X1    g607(.A(new_n782), .ZN(new_n809));
  OAI21_X1  g608(.A(new_n363), .B1(new_n808), .B2(new_n809), .ZN(new_n810));
  INV_X1    g609(.A(KEYINPUT119), .ZN(new_n811));
  INV_X1    g610(.A(KEYINPUT57), .ZN(new_n812));
  NAND3_X1  g611(.A1(new_n810), .A2(new_n811), .A3(new_n812), .ZN(new_n813));
  INV_X1    g612(.A(KEYINPUT121), .ZN(new_n814));
  NAND4_X1  g613(.A1(new_n755), .A2(new_n757), .A3(new_n525), .A4(new_n759), .ZN(new_n815));
  OR2_X1    g614(.A1(new_n600), .A2(new_n768), .ZN(new_n816));
  AND3_X1   g615(.A1(new_n815), .A2(new_n816), .A3(KEYINPUT120), .ZN(new_n817));
  AOI21_X1  g616(.A(KEYINPUT120), .B1(new_n815), .B2(new_n816), .ZN(new_n818));
  OAI21_X1  g617(.A(new_n632), .B1(new_n817), .B2(new_n818), .ZN(new_n819));
  NAND2_X1  g618(.A1(new_n819), .A2(new_n807), .ZN(new_n820));
  AOI21_X1  g619(.A(new_n814), .B1(new_n820), .B2(new_n549), .ZN(new_n821));
  AOI211_X1 g620(.A(KEYINPUT121), .B(new_n631), .C1(new_n819), .C2(new_n807), .ZN(new_n822));
  NOR3_X1   g621(.A1(new_n821), .A2(new_n822), .A3(new_n809), .ZN(new_n823));
  NAND2_X1  g622(.A1(new_n363), .A2(KEYINPUT57), .ZN(new_n824));
  OAI211_X1 g623(.A(new_n802), .B(new_n813), .C1(new_n823), .C2(new_n824), .ZN(new_n825));
  AND2_X1   g624(.A1(new_n438), .A2(new_n784), .ZN(new_n826));
  XNOR2_X1  g625(.A(new_n826), .B(KEYINPUT118), .ZN(new_n827));
  INV_X1    g626(.A(new_n827), .ZN(new_n828));
  NAND3_X1  g627(.A1(new_n825), .A2(new_n525), .A3(new_n828), .ZN(new_n829));
  INV_X1    g628(.A(KEYINPUT123), .ZN(new_n830));
  NAND2_X1  g629(.A1(new_n829), .A2(new_n830), .ZN(new_n831));
  NAND4_X1  g630(.A1(new_n825), .A2(KEYINPUT123), .A3(new_n525), .A4(new_n828), .ZN(new_n832));
  NAND3_X1  g631(.A1(new_n831), .A2(G141gat), .A3(new_n832), .ZN(new_n833));
  INV_X1    g632(.A(G141gat), .ZN(new_n834));
  NAND4_X1  g633(.A1(new_n801), .A2(new_n834), .A3(new_n525), .A4(new_n826), .ZN(new_n835));
  INV_X1    g634(.A(new_n835), .ZN(new_n836));
  XNOR2_X1  g635(.A(KEYINPUT122), .B(KEYINPUT58), .ZN(new_n837));
  NOR2_X1   g636(.A1(new_n836), .A2(new_n837), .ZN(new_n838));
  NAND2_X1  g637(.A1(new_n833), .A2(new_n838), .ZN(new_n839));
  AND2_X1   g638(.A1(new_n802), .A2(new_n813), .ZN(new_n840));
  INV_X1    g639(.A(new_n821), .ZN(new_n841));
  INV_X1    g640(.A(new_n822), .ZN(new_n842));
  NAND3_X1  g641(.A1(new_n841), .A2(new_n842), .A3(new_n782), .ZN(new_n843));
  NAND3_X1  g642(.A1(new_n843), .A2(KEYINPUT57), .A3(new_n363), .ZN(new_n844));
  AOI21_X1  g643(.A(new_n827), .B1(new_n840), .B2(new_n844), .ZN(new_n845));
  AOI21_X1  g644(.A(new_n834), .B1(new_n845), .B2(new_n650), .ZN(new_n846));
  OAI21_X1  g645(.A(KEYINPUT58), .B1(new_n846), .B2(new_n836), .ZN(new_n847));
  NAND2_X1  g646(.A1(new_n839), .A2(new_n847), .ZN(G1344gat));
  INV_X1    g647(.A(KEYINPUT59), .ZN(new_n849));
  NAND2_X1  g648(.A1(new_n825), .A2(new_n828), .ZN(new_n850));
  OAI211_X1 g649(.A(new_n849), .B(G148gat), .C1(new_n850), .C2(new_n600), .ZN(new_n851));
  INV_X1    g650(.A(G148gat), .ZN(new_n852));
  NAND2_X1  g651(.A1(new_n767), .A2(new_n772), .ZN(new_n853));
  AOI21_X1  g652(.A(new_n631), .B1(new_n819), .B2(new_n853), .ZN(new_n854));
  AND2_X1   g653(.A1(new_n602), .A2(new_n786), .ZN(new_n855));
  OAI211_X1 g654(.A(new_n812), .B(new_n363), .C1(new_n854), .C2(new_n855), .ZN(new_n856));
  INV_X1    g655(.A(new_n856), .ZN(new_n857));
  AOI21_X1  g656(.A(new_n857), .B1(KEYINPUT57), .B2(new_n810), .ZN(new_n858));
  AND2_X1   g657(.A1(new_n858), .A2(new_n601), .ZN(new_n859));
  AOI21_X1  g658(.A(new_n852), .B1(new_n859), .B2(new_n828), .ZN(new_n860));
  XOR2_X1   g659(.A(KEYINPUT124), .B(KEYINPUT59), .Z(new_n861));
  OAI21_X1  g660(.A(new_n851), .B1(new_n860), .B2(new_n861), .ZN(new_n862));
  NAND2_X1  g661(.A1(new_n801), .A2(new_n826), .ZN(new_n863));
  NAND2_X1  g662(.A1(new_n601), .A2(new_n852), .ZN(new_n864));
  OAI21_X1  g663(.A(new_n862), .B1(new_n863), .B2(new_n864), .ZN(G1345gat));
  NAND3_X1  g664(.A1(new_n845), .A2(G155gat), .A3(new_n631), .ZN(new_n866));
  OAI21_X1  g665(.A(new_n331), .B1(new_n863), .B2(new_n549), .ZN(new_n867));
  AND2_X1   g666(.A1(new_n866), .A2(new_n867), .ZN(G1346gat));
  INV_X1    g667(.A(KEYINPUT125), .ZN(new_n869));
  NAND3_X1  g668(.A1(new_n845), .A2(new_n869), .A3(new_n581), .ZN(new_n870));
  OAI21_X1  g669(.A(KEYINPUT125), .B1(new_n850), .B2(new_n632), .ZN(new_n871));
  NAND3_X1  g670(.A1(new_n870), .A2(new_n871), .A3(G162gat), .ZN(new_n872));
  NAND3_X1  g671(.A1(new_n801), .A2(new_n332), .A3(new_n826), .ZN(new_n873));
  OAI21_X1  g672(.A(new_n872), .B1(new_n632), .B2(new_n873), .ZN(G1347gat));
  NOR2_X1   g673(.A1(new_n654), .A2(new_n604), .ZN(new_n875));
  NAND2_X1  g674(.A1(new_n783), .A2(new_n875), .ZN(new_n876));
  OAI21_X1  g675(.A(G169gat), .B1(new_n876), .B2(new_n786), .ZN(new_n877));
  INV_X1    g676(.A(new_n650), .ZN(new_n878));
  OR2_X1    g677(.A1(new_n878), .A2(G169gat), .ZN(new_n879));
  OAI21_X1  g678(.A(new_n877), .B1(new_n876), .B2(new_n879), .ZN(G1348gat));
  INV_X1    g679(.A(new_n876), .ZN(new_n881));
  NAND2_X1  g680(.A1(new_n881), .A2(new_n601), .ZN(new_n882));
  XNOR2_X1  g681(.A(new_n882), .B(G176gat), .ZN(G1349gat));
  AOI21_X1  g682(.A(new_n221), .B1(new_n881), .B2(new_n631), .ZN(new_n884));
  NOR2_X1   g683(.A1(new_n876), .A2(new_n549), .ZN(new_n885));
  AOI21_X1  g684(.A(new_n884), .B1(new_n224), .B2(new_n885), .ZN(new_n886));
  INV_X1    g685(.A(KEYINPUT127), .ZN(new_n887));
  OAI21_X1  g686(.A(new_n886), .B1(new_n887), .B2(KEYINPUT60), .ZN(new_n888));
  INV_X1    g687(.A(KEYINPUT126), .ZN(new_n889));
  NAND2_X1  g688(.A1(new_n889), .A2(KEYINPUT60), .ZN(new_n890));
  NOR2_X1   g689(.A1(new_n890), .A2(KEYINPUT127), .ZN(new_n891));
  AOI22_X1  g690(.A1(new_n888), .A2(new_n890), .B1(new_n886), .B2(new_n891), .ZN(G1350gat));
  NAND2_X1  g691(.A1(new_n881), .A2(new_n581), .ZN(new_n893));
  OAI21_X1  g692(.A(KEYINPUT61), .B1(new_n893), .B2(new_n207), .ZN(new_n894));
  NAND2_X1  g693(.A1(new_n893), .A2(G190gat), .ZN(new_n895));
  MUX2_X1   g694(.A(KEYINPUT61), .B(new_n894), .S(new_n895), .Z(G1351gat));
  AND2_X1   g695(.A1(new_n438), .A2(new_n875), .ZN(new_n897));
  NAND3_X1  g696(.A1(new_n858), .A2(new_n525), .A3(new_n897), .ZN(new_n898));
  NAND2_X1  g697(.A1(new_n898), .A2(G197gat), .ZN(new_n899));
  NAND2_X1  g698(.A1(new_n801), .A2(new_n897), .ZN(new_n900));
  OR2_X1    g699(.A1(new_n900), .A2(G197gat), .ZN(new_n901));
  OAI21_X1  g700(.A(new_n899), .B1(new_n878), .B2(new_n901), .ZN(G1352gat));
  NAND2_X1  g701(.A1(new_n859), .A2(new_n897), .ZN(new_n903));
  NAND2_X1  g702(.A1(new_n903), .A2(G204gat), .ZN(new_n904));
  NOR3_X1   g703(.A1(new_n900), .A2(G204gat), .A3(new_n600), .ZN(new_n905));
  XNOR2_X1  g704(.A(new_n905), .B(KEYINPUT62), .ZN(new_n906));
  NAND2_X1  g705(.A1(new_n904), .A2(new_n906), .ZN(G1353gat));
  NAND3_X1  g706(.A1(new_n858), .A2(new_n631), .A3(new_n897), .ZN(new_n908));
  AND3_X1   g707(.A1(new_n908), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n909));
  AOI21_X1  g708(.A(KEYINPUT63), .B1(new_n908), .B2(G211gat), .ZN(new_n910));
  NAND2_X1  g709(.A1(new_n631), .A2(new_n539), .ZN(new_n911));
  OAI22_X1  g710(.A1(new_n909), .A2(new_n910), .B1(new_n900), .B2(new_n911), .ZN(G1354gat));
  NAND3_X1  g711(.A1(new_n858), .A2(new_n581), .A3(new_n897), .ZN(new_n913));
  NAND2_X1  g712(.A1(new_n913), .A2(G218gat), .ZN(new_n914));
  OR2_X1    g713(.A1(new_n900), .A2(G218gat), .ZN(new_n915));
  OAI21_X1  g714(.A(new_n914), .B1(new_n632), .B2(new_n915), .ZN(G1355gat));
endmodule


