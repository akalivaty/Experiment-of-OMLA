//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 1 0 1 1 0 1 1 1 1 0 1 0 0 1 1 1 0 1 0 0 1 1 1 0 1 0 0 0 1 0 1 0 1 0 0 1 0 0 1 0 1 0 1 1 0 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:27:38 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n713, new_n714, new_n715, new_n716, new_n717,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n731, new_n732, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n744, new_n745, new_n746, new_n747, new_n748, new_n749,
    new_n750, new_n751, new_n752, new_n753, new_n755, new_n756, new_n757,
    new_n758, new_n759, new_n760, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n786, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n805, new_n806, new_n807, new_n808, new_n809, new_n810,
    new_n811, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n929, new_n930, new_n931,
    new_n932, new_n933, new_n934, new_n935, new_n936, new_n937, new_n938,
    new_n939, new_n940, new_n941, new_n942, new_n943, new_n944, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n955, new_n956, new_n957, new_n959, new_n960, new_n961, new_n962,
    new_n963, new_n964, new_n965, new_n966, new_n967, new_n969, new_n970,
    new_n971, new_n972, new_n973, new_n974, new_n975, new_n976, new_n978,
    new_n979, new_n980, new_n981, new_n982, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1017, new_n1018, new_n1019,
    new_n1020, new_n1021, new_n1022, new_n1023, new_n1024, new_n1025,
    new_n1026;
  INV_X1    g000(.A(G472), .ZN(new_n187));
  INV_X1    g001(.A(G237), .ZN(new_n188));
  INV_X1    g002(.A(G953), .ZN(new_n189));
  NAND3_X1  g003(.A1(new_n188), .A2(new_n189), .A3(G210), .ZN(new_n190));
  XNOR2_X1  g004(.A(new_n190), .B(KEYINPUT27), .ZN(new_n191));
  XNOR2_X1  g005(.A(KEYINPUT26), .B(G101), .ZN(new_n192));
  XNOR2_X1  g006(.A(new_n191), .B(new_n192), .ZN(new_n193));
  INV_X1    g007(.A(new_n193), .ZN(new_n194));
  INV_X1    g008(.A(G113), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n195), .A2(KEYINPUT2), .ZN(new_n196));
  INV_X1    g010(.A(KEYINPUT2), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n197), .A2(G113), .ZN(new_n198));
  INV_X1    g012(.A(G116), .ZN(new_n199));
  NOR2_X1   g013(.A1(new_n199), .A2(G119), .ZN(new_n200));
  INV_X1    g014(.A(G119), .ZN(new_n201));
  NOR2_X1   g015(.A1(new_n201), .A2(G116), .ZN(new_n202));
  OAI211_X1 g016(.A(new_n196), .B(new_n198), .C1(new_n200), .C2(new_n202), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n196), .A2(new_n198), .ZN(new_n204));
  XNOR2_X1  g018(.A(G116), .B(G119), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n204), .A2(new_n205), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n203), .A2(new_n206), .ZN(new_n207));
  INV_X1    g021(.A(new_n207), .ZN(new_n208));
  INV_X1    g022(.A(G137), .ZN(new_n209));
  NAND3_X1  g023(.A1(new_n209), .A2(KEYINPUT11), .A3(G134), .ZN(new_n210));
  INV_X1    g024(.A(KEYINPUT11), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n211), .A2(G137), .ZN(new_n212));
  AND2_X1   g026(.A1(new_n210), .A2(new_n212), .ZN(new_n213));
  INV_X1    g027(.A(G134), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n214), .A2(KEYINPUT65), .ZN(new_n215));
  INV_X1    g029(.A(KEYINPUT65), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n216), .A2(G134), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n209), .A2(KEYINPUT11), .ZN(new_n218));
  NAND3_X1  g032(.A1(new_n215), .A2(new_n217), .A3(new_n218), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n213), .A2(new_n219), .ZN(new_n220));
  NAND2_X1  g034(.A1(KEYINPUT66), .A2(G131), .ZN(new_n221));
  INV_X1    g035(.A(new_n221), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n220), .A2(new_n222), .ZN(new_n223));
  NAND3_X1  g037(.A1(new_n213), .A2(new_n221), .A3(new_n219), .ZN(new_n224));
  INV_X1    g038(.A(KEYINPUT64), .ZN(new_n225));
  INV_X1    g039(.A(KEYINPUT0), .ZN(new_n226));
  INV_X1    g040(.A(G128), .ZN(new_n227));
  NAND3_X1  g041(.A1(new_n225), .A2(new_n226), .A3(new_n227), .ZN(new_n228));
  OAI21_X1  g042(.A(KEYINPUT64), .B1(KEYINPUT0), .B2(G128), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n228), .A2(new_n229), .ZN(new_n230));
  NOR2_X1   g044(.A1(new_n226), .A2(new_n227), .ZN(new_n231));
  INV_X1    g045(.A(new_n231), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n230), .A2(new_n232), .ZN(new_n233));
  INV_X1    g047(.A(G146), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n234), .A2(G143), .ZN(new_n235));
  INV_X1    g049(.A(G143), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n236), .A2(G146), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n235), .A2(new_n237), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n233), .A2(new_n238), .ZN(new_n239));
  XNOR2_X1  g053(.A(G143), .B(G146), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n232), .A2(new_n240), .ZN(new_n241));
  AOI22_X1  g055(.A1(new_n223), .A2(new_n224), .B1(new_n239), .B2(new_n241), .ZN(new_n242));
  INV_X1    g056(.A(KEYINPUT1), .ZN(new_n243));
  NAND4_X1  g057(.A1(new_n235), .A2(new_n237), .A3(new_n243), .A4(G128), .ZN(new_n244));
  NOR2_X1   g058(.A1(new_n234), .A2(G143), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n245), .A2(KEYINPUT1), .ZN(new_n246));
  OAI211_X1 g060(.A(new_n244), .B(new_n246), .C1(G128), .C2(new_n240), .ZN(new_n247));
  AOI21_X1  g061(.A(G137), .B1(new_n215), .B2(new_n217), .ZN(new_n248));
  NOR2_X1   g062(.A1(new_n209), .A2(G134), .ZN(new_n249));
  OAI21_X1  g063(.A(G131), .B1(new_n248), .B2(new_n249), .ZN(new_n250));
  INV_X1    g064(.A(G131), .ZN(new_n251));
  NAND3_X1  g065(.A1(new_n213), .A2(new_n251), .A3(new_n219), .ZN(new_n252));
  AND3_X1   g066(.A1(new_n247), .A2(new_n250), .A3(new_n252), .ZN(new_n253));
  OAI21_X1  g067(.A(KEYINPUT30), .B1(new_n242), .B2(new_n253), .ZN(new_n254));
  AOI21_X1  g068(.A(new_n231), .B1(new_n228), .B2(new_n229), .ZN(new_n255));
  OAI21_X1  g069(.A(new_n241), .B1(new_n255), .B2(new_n240), .ZN(new_n256));
  AND3_X1   g070(.A1(new_n213), .A2(new_n221), .A3(new_n219), .ZN(new_n257));
  AOI21_X1  g071(.A(new_n221), .B1(new_n213), .B2(new_n219), .ZN(new_n258));
  OAI21_X1  g072(.A(new_n256), .B1(new_n257), .B2(new_n258), .ZN(new_n259));
  INV_X1    g073(.A(KEYINPUT30), .ZN(new_n260));
  NAND3_X1  g074(.A1(new_n247), .A2(new_n250), .A3(new_n252), .ZN(new_n261));
  NAND3_X1  g075(.A1(new_n259), .A2(new_n260), .A3(new_n261), .ZN(new_n262));
  AOI21_X1  g076(.A(new_n208), .B1(new_n254), .B2(new_n262), .ZN(new_n263));
  NAND3_X1  g077(.A1(new_n259), .A2(new_n208), .A3(new_n261), .ZN(new_n264));
  INV_X1    g078(.A(new_n264), .ZN(new_n265));
  OAI21_X1  g079(.A(new_n194), .B1(new_n263), .B2(new_n265), .ZN(new_n266));
  AOI21_X1  g080(.A(new_n208), .B1(new_n259), .B2(new_n261), .ZN(new_n267));
  OAI21_X1  g081(.A(KEYINPUT28), .B1(new_n265), .B2(new_n267), .ZN(new_n268));
  INV_X1    g082(.A(KEYINPUT28), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n264), .A2(new_n269), .ZN(new_n270));
  NAND3_X1  g084(.A1(new_n268), .A2(new_n270), .A3(new_n193), .ZN(new_n271));
  INV_X1    g085(.A(KEYINPUT29), .ZN(new_n272));
  AND3_X1   g086(.A1(new_n266), .A2(new_n271), .A3(new_n272), .ZN(new_n273));
  OAI21_X1  g087(.A(new_n207), .B1(new_n242), .B2(new_n253), .ZN(new_n274));
  AOI21_X1  g088(.A(new_n269), .B1(new_n274), .B2(new_n264), .ZN(new_n275));
  INV_X1    g089(.A(new_n270), .ZN(new_n276));
  OAI21_X1  g090(.A(KEYINPUT68), .B1(new_n275), .B2(new_n276), .ZN(new_n277));
  INV_X1    g091(.A(KEYINPUT68), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n270), .A2(new_n278), .ZN(new_n279));
  NOR2_X1   g093(.A1(new_n194), .A2(new_n272), .ZN(new_n280));
  NAND3_X1  g094(.A1(new_n277), .A2(new_n279), .A3(new_n280), .ZN(new_n281));
  INV_X1    g095(.A(G902), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n281), .A2(new_n282), .ZN(new_n283));
  AOI21_X1  g097(.A(new_n273), .B1(new_n283), .B2(KEYINPUT69), .ZN(new_n284));
  INV_X1    g098(.A(KEYINPUT69), .ZN(new_n285));
  NAND3_X1  g099(.A1(new_n281), .A2(new_n285), .A3(new_n282), .ZN(new_n286));
  AOI21_X1  g100(.A(new_n187), .B1(new_n284), .B2(new_n286), .ZN(new_n287));
  AND3_X1   g101(.A1(new_n259), .A2(new_n260), .A3(new_n261), .ZN(new_n288));
  AOI21_X1  g102(.A(new_n260), .B1(new_n259), .B2(new_n261), .ZN(new_n289));
  OAI21_X1  g103(.A(new_n207), .B1(new_n288), .B2(new_n289), .ZN(new_n290));
  NAND3_X1  g104(.A1(new_n290), .A2(new_n264), .A3(new_n193), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n291), .A2(KEYINPUT31), .ZN(new_n292));
  OAI21_X1  g106(.A(new_n194), .B1(new_n275), .B2(new_n276), .ZN(new_n293));
  INV_X1    g107(.A(KEYINPUT31), .ZN(new_n294));
  NAND4_X1  g108(.A1(new_n290), .A2(new_n294), .A3(new_n264), .A4(new_n193), .ZN(new_n295));
  NAND3_X1  g109(.A1(new_n292), .A2(new_n293), .A3(new_n295), .ZN(new_n296));
  NOR2_X1   g110(.A1(G472), .A2(G902), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n296), .A2(new_n297), .ZN(new_n298));
  INV_X1    g112(.A(KEYINPUT32), .ZN(new_n299));
  NAND3_X1  g113(.A1(new_n298), .A2(KEYINPUT67), .A3(new_n299), .ZN(new_n300));
  NAND2_X1  g114(.A1(new_n298), .A2(new_n299), .ZN(new_n301));
  INV_X1    g115(.A(KEYINPUT67), .ZN(new_n302));
  NAND3_X1  g116(.A1(new_n296), .A2(KEYINPUT32), .A3(new_n297), .ZN(new_n303));
  NAND3_X1  g117(.A1(new_n301), .A2(new_n302), .A3(new_n303), .ZN(new_n304));
  AOI21_X1  g118(.A(new_n287), .B1(new_n300), .B2(new_n304), .ZN(new_n305));
  INV_X1    g119(.A(KEYINPUT16), .ZN(new_n306));
  INV_X1    g120(.A(G140), .ZN(new_n307));
  NAND3_X1  g121(.A1(new_n306), .A2(new_n307), .A3(G125), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n308), .A2(KEYINPUT73), .ZN(new_n309));
  INV_X1    g123(.A(G125), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n310), .A2(G140), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n307), .A2(G125), .ZN(new_n312));
  NAND3_X1  g126(.A1(new_n311), .A2(new_n312), .A3(KEYINPUT72), .ZN(new_n313));
  INV_X1    g127(.A(KEYINPUT72), .ZN(new_n314));
  NAND3_X1  g128(.A1(new_n314), .A2(new_n310), .A3(G140), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n313), .A2(new_n315), .ZN(new_n316));
  AOI21_X1  g130(.A(new_n309), .B1(new_n316), .B2(KEYINPUT16), .ZN(new_n317));
  AOI211_X1 g131(.A(KEYINPUT73), .B(new_n306), .C1(new_n313), .C2(new_n315), .ZN(new_n318));
  OAI21_X1  g132(.A(G146), .B1(new_n317), .B2(new_n318), .ZN(new_n319));
  INV_X1    g133(.A(KEYINPUT74), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n319), .A2(new_n320), .ZN(new_n321));
  OAI211_X1 g135(.A(KEYINPUT74), .B(G146), .C1(new_n317), .C2(new_n318), .ZN(new_n322));
  XNOR2_X1  g136(.A(G125), .B(G140), .ZN(new_n323));
  AOI21_X1  g137(.A(KEYINPUT75), .B1(new_n323), .B2(new_n234), .ZN(new_n324));
  AND4_X1   g138(.A1(KEYINPUT75), .A2(new_n311), .A3(new_n312), .A4(new_n234), .ZN(new_n325));
  NOR2_X1   g139(.A1(new_n324), .A2(new_n325), .ZN(new_n326));
  XNOR2_X1  g140(.A(G119), .B(G128), .ZN(new_n327));
  XNOR2_X1  g141(.A(new_n327), .B(KEYINPUT70), .ZN(new_n328));
  XNOR2_X1  g142(.A(KEYINPUT24), .B(G110), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n328), .A2(new_n329), .ZN(new_n330));
  INV_X1    g144(.A(KEYINPUT23), .ZN(new_n331));
  OAI21_X1  g145(.A(new_n331), .B1(new_n201), .B2(G128), .ZN(new_n332));
  NAND3_X1  g146(.A1(new_n227), .A2(KEYINPUT23), .A3(G119), .ZN(new_n333));
  OAI211_X1 g147(.A(new_n332), .B(new_n333), .C1(G119), .C2(new_n227), .ZN(new_n334));
  OR2_X1    g148(.A1(new_n334), .A2(G110), .ZN(new_n335));
  AOI21_X1  g149(.A(new_n326), .B1(new_n330), .B2(new_n335), .ZN(new_n336));
  NAND3_X1  g150(.A1(new_n321), .A2(new_n322), .A3(new_n336), .ZN(new_n337));
  INV_X1    g151(.A(KEYINPUT73), .ZN(new_n338));
  NAND3_X1  g152(.A1(new_n316), .A2(new_n338), .A3(KEYINPUT16), .ZN(new_n339));
  NOR3_X1   g153(.A1(new_n307), .A2(KEYINPUT72), .A3(G125), .ZN(new_n340));
  AOI21_X1  g154(.A(new_n340), .B1(new_n323), .B2(KEYINPUT72), .ZN(new_n341));
  NOR2_X1   g155(.A1(new_n341), .A2(new_n306), .ZN(new_n342));
  OAI211_X1 g156(.A(new_n234), .B(new_n339), .C1(new_n342), .C2(new_n309), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n343), .A2(new_n319), .ZN(new_n344));
  INV_X1    g158(.A(new_n328), .ZN(new_n345));
  INV_X1    g159(.A(new_n329), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n334), .A2(G110), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n347), .A2(KEYINPUT71), .ZN(new_n348));
  INV_X1    g162(.A(KEYINPUT71), .ZN(new_n349));
  NAND3_X1  g163(.A1(new_n334), .A2(new_n349), .A3(G110), .ZN(new_n350));
  AOI22_X1  g164(.A1(new_n345), .A2(new_n346), .B1(new_n348), .B2(new_n350), .ZN(new_n351));
  NAND2_X1  g165(.A1(new_n344), .A2(new_n351), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n337), .A2(new_n352), .ZN(new_n353));
  XNOR2_X1  g167(.A(KEYINPUT22), .B(G137), .ZN(new_n354));
  NAND3_X1  g168(.A1(new_n189), .A2(G221), .A3(G234), .ZN(new_n355));
  XNOR2_X1  g169(.A(new_n354), .B(new_n355), .ZN(new_n356));
  INV_X1    g170(.A(new_n356), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n353), .A2(new_n357), .ZN(new_n358));
  NAND3_X1  g172(.A1(new_n337), .A2(new_n352), .A3(new_n356), .ZN(new_n359));
  NAND3_X1  g173(.A1(new_n358), .A2(new_n282), .A3(new_n359), .ZN(new_n360));
  INV_X1    g174(.A(KEYINPUT25), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n360), .A2(new_n361), .ZN(new_n362));
  NAND4_X1  g176(.A1(new_n358), .A2(KEYINPUT25), .A3(new_n282), .A4(new_n359), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n362), .A2(new_n363), .ZN(new_n364));
  INV_X1    g178(.A(G217), .ZN(new_n365));
  AOI21_X1  g179(.A(new_n365), .B1(G234), .B2(new_n282), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n364), .A2(new_n366), .ZN(new_n367));
  NOR2_X1   g181(.A1(new_n366), .A2(G902), .ZN(new_n368));
  XOR2_X1   g182(.A(new_n368), .B(KEYINPUT76), .Z(new_n369));
  NAND2_X1  g183(.A1(new_n358), .A2(new_n359), .ZN(new_n370));
  OAI21_X1  g184(.A(new_n367), .B1(new_n369), .B2(new_n370), .ZN(new_n371));
  OAI21_X1  g185(.A(KEYINPUT77), .B1(new_n305), .B2(new_n371), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n283), .A2(KEYINPUT69), .ZN(new_n373));
  INV_X1    g187(.A(new_n273), .ZN(new_n374));
  NAND3_X1  g188(.A1(new_n373), .A2(new_n286), .A3(new_n374), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n375), .A2(G472), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n303), .A2(new_n302), .ZN(new_n377));
  AOI21_X1  g191(.A(KEYINPUT32), .B1(new_n296), .B2(new_n297), .ZN(new_n378));
  NOR2_X1   g192(.A1(new_n377), .A2(new_n378), .ZN(new_n379));
  INV_X1    g193(.A(new_n300), .ZN(new_n380));
  OAI21_X1  g194(.A(new_n376), .B1(new_n379), .B2(new_n380), .ZN(new_n381));
  INV_X1    g195(.A(KEYINPUT77), .ZN(new_n382));
  INV_X1    g196(.A(new_n366), .ZN(new_n383));
  AOI21_X1  g197(.A(new_n383), .B1(new_n362), .B2(new_n363), .ZN(new_n384));
  INV_X1    g198(.A(new_n369), .ZN(new_n385));
  INV_X1    g199(.A(new_n370), .ZN(new_n386));
  AOI21_X1  g200(.A(new_n384), .B1(new_n385), .B2(new_n386), .ZN(new_n387));
  NAND3_X1  g201(.A1(new_n381), .A2(new_n382), .A3(new_n387), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n372), .A2(new_n388), .ZN(new_n389));
  OAI21_X1  g203(.A(G214), .B1(G237), .B2(G902), .ZN(new_n390));
  INV_X1    g204(.A(new_n390), .ZN(new_n391));
  OAI21_X1  g205(.A(G210), .B1(G237), .B2(G902), .ZN(new_n392));
  INV_X1    g206(.A(new_n392), .ZN(new_n393));
  XNOR2_X1  g207(.A(G110), .B(G122), .ZN(new_n394));
  XOR2_X1   g208(.A(new_n394), .B(KEYINPUT81), .Z(new_n395));
  INV_X1    g209(.A(G104), .ZN(new_n396));
  OAI21_X1  g210(.A(KEYINPUT3), .B1(new_n396), .B2(G107), .ZN(new_n397));
  INV_X1    g211(.A(KEYINPUT3), .ZN(new_n398));
  INV_X1    g212(.A(G107), .ZN(new_n399));
  NAND3_X1  g213(.A1(new_n398), .A2(new_n399), .A3(G104), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n396), .A2(G107), .ZN(new_n401));
  NAND3_X1  g215(.A1(new_n397), .A2(new_n400), .A3(new_n401), .ZN(new_n402));
  INV_X1    g216(.A(KEYINPUT4), .ZN(new_n403));
  NAND3_X1  g217(.A1(new_n402), .A2(new_n403), .A3(G101), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n207), .A2(new_n404), .ZN(new_n405));
  AOI21_X1  g219(.A(G101), .B1(new_n396), .B2(G107), .ZN(new_n406));
  NAND3_X1  g220(.A1(new_n397), .A2(new_n406), .A3(new_n400), .ZN(new_n407));
  INV_X1    g221(.A(KEYINPUT78), .ZN(new_n408));
  NAND2_X1  g222(.A1(new_n407), .A2(new_n408), .ZN(new_n409));
  NAND4_X1  g223(.A1(new_n397), .A2(new_n406), .A3(new_n400), .A4(KEYINPUT78), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n409), .A2(new_n410), .ZN(new_n411));
  AOI21_X1  g225(.A(new_n403), .B1(new_n402), .B2(G101), .ZN(new_n412));
  AOI21_X1  g226(.A(new_n405), .B1(new_n411), .B2(new_n412), .ZN(new_n413));
  INV_X1    g227(.A(G101), .ZN(new_n414));
  NAND2_X1  g228(.A1(new_n399), .A2(G104), .ZN(new_n415));
  AOI21_X1  g229(.A(new_n414), .B1(new_n415), .B2(new_n401), .ZN(new_n416));
  AOI21_X1  g230(.A(new_n416), .B1(new_n409), .B2(new_n410), .ZN(new_n417));
  NAND2_X1  g231(.A1(new_n205), .A2(KEYINPUT5), .ZN(new_n418));
  INV_X1    g232(.A(KEYINPUT5), .ZN(new_n419));
  AOI21_X1  g233(.A(new_n195), .B1(new_n200), .B2(new_n419), .ZN(new_n420));
  AOI22_X1  g234(.A1(new_n418), .A2(new_n420), .B1(new_n205), .B2(new_n204), .ZN(new_n421));
  AND2_X1   g235(.A1(new_n417), .A2(new_n421), .ZN(new_n422));
  OAI21_X1  g236(.A(new_n395), .B1(new_n413), .B2(new_n422), .ZN(new_n423));
  NOR2_X1   g237(.A1(new_n423), .A2(KEYINPUT6), .ZN(new_n424));
  OAI211_X1 g238(.A(G125), .B(new_n241), .C1(new_n255), .C2(new_n240), .ZN(new_n425));
  AND2_X1   g239(.A1(new_n425), .A2(KEYINPUT84), .ZN(new_n426));
  INV_X1    g240(.A(KEYINPUT84), .ZN(new_n427));
  OAI21_X1  g241(.A(new_n425), .B1(G125), .B2(new_n247), .ZN(new_n428));
  AOI21_X1  g242(.A(new_n426), .B1(new_n427), .B2(new_n428), .ZN(new_n429));
  INV_X1    g243(.A(G224), .ZN(new_n430));
  NOR2_X1   g244(.A1(new_n430), .A2(G953), .ZN(new_n431));
  XNOR2_X1  g245(.A(new_n429), .B(new_n431), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n411), .A2(new_n412), .ZN(new_n433));
  AND2_X1   g247(.A1(new_n207), .A2(new_n404), .ZN(new_n434));
  AOI22_X1  g248(.A1(new_n433), .A2(new_n434), .B1(new_n417), .B2(new_n421), .ZN(new_n435));
  INV_X1    g249(.A(new_n395), .ZN(new_n436));
  OAI21_X1  g250(.A(KEYINPUT82), .B1(new_n435), .B2(new_n436), .ZN(new_n437));
  INV_X1    g251(.A(KEYINPUT6), .ZN(new_n438));
  AOI21_X1  g252(.A(new_n438), .B1(new_n435), .B2(new_n394), .ZN(new_n439));
  INV_X1    g253(.A(KEYINPUT82), .ZN(new_n440));
  OAI211_X1 g254(.A(new_n440), .B(new_n395), .C1(new_n413), .C2(new_n422), .ZN(new_n441));
  NAND3_X1  g255(.A1(new_n437), .A2(new_n439), .A3(new_n441), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n442), .A2(KEYINPUT83), .ZN(new_n443));
  INV_X1    g257(.A(KEYINPUT83), .ZN(new_n444));
  NAND4_X1  g258(.A1(new_n437), .A2(new_n439), .A3(new_n444), .A4(new_n441), .ZN(new_n445));
  AOI211_X1 g259(.A(new_n424), .B(new_n432), .C1(new_n443), .C2(new_n445), .ZN(new_n446));
  INV_X1    g260(.A(KEYINPUT86), .ZN(new_n447));
  INV_X1    g261(.A(KEYINPUT85), .ZN(new_n448));
  AOI21_X1  g262(.A(new_n447), .B1(new_n417), .B2(new_n448), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n449), .A2(new_n421), .ZN(new_n450));
  XNOR2_X1  g264(.A(new_n394), .B(KEYINPUT8), .ZN(new_n451));
  INV_X1    g265(.A(new_n421), .ZN(new_n452));
  INV_X1    g266(.A(new_n416), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n411), .A2(new_n453), .ZN(new_n454));
  OAI21_X1  g268(.A(new_n452), .B1(new_n454), .B2(KEYINPUT86), .ZN(new_n455));
  OAI211_X1 g269(.A(new_n450), .B(new_n451), .C1(new_n455), .C2(new_n449), .ZN(new_n456));
  OAI21_X1  g270(.A(KEYINPUT7), .B1(new_n430), .B2(G953), .ZN(new_n457));
  AOI22_X1  g271(.A1(new_n435), .A2(new_n394), .B1(new_n428), .B2(new_n457), .ZN(new_n458));
  AND2_X1   g272(.A1(new_n456), .A2(new_n458), .ZN(new_n459));
  INV_X1    g273(.A(new_n457), .ZN(new_n460));
  NAND2_X1  g274(.A1(new_n429), .A2(new_n460), .ZN(new_n461));
  AND2_X1   g275(.A1(new_n461), .A2(KEYINPUT87), .ZN(new_n462));
  NOR2_X1   g276(.A1(new_n461), .A2(KEYINPUT87), .ZN(new_n463));
  OAI21_X1  g277(.A(new_n459), .B1(new_n462), .B2(new_n463), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n464), .A2(new_n282), .ZN(new_n465));
  OAI21_X1  g279(.A(new_n393), .B1(new_n446), .B2(new_n465), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n443), .A2(new_n445), .ZN(new_n467));
  INV_X1    g281(.A(new_n432), .ZN(new_n468));
  INV_X1    g282(.A(new_n424), .ZN(new_n469));
  NAND3_X1  g283(.A1(new_n467), .A2(new_n468), .A3(new_n469), .ZN(new_n470));
  XNOR2_X1  g284(.A(new_n461), .B(KEYINPUT87), .ZN(new_n471));
  AOI21_X1  g285(.A(G902), .B1(new_n471), .B2(new_n459), .ZN(new_n472));
  NAND3_X1  g286(.A1(new_n470), .A2(new_n472), .A3(new_n392), .ZN(new_n473));
  AOI21_X1  g287(.A(new_n391), .B1(new_n466), .B2(new_n473), .ZN(new_n474));
  XNOR2_X1  g288(.A(KEYINPUT9), .B(G234), .ZN(new_n475));
  OAI21_X1  g289(.A(G221), .B1(new_n475), .B2(G902), .ZN(new_n476));
  INV_X1    g290(.A(new_n476), .ZN(new_n477));
  AOI21_X1  g291(.A(G128), .B1(new_n235), .B2(new_n237), .ZN(new_n478));
  NOR2_X1   g292(.A1(new_n237), .A2(new_n243), .ZN(new_n479));
  OAI21_X1  g293(.A(KEYINPUT79), .B1(new_n478), .B2(new_n479), .ZN(new_n480));
  INV_X1    g294(.A(KEYINPUT79), .ZN(new_n481));
  OAI211_X1 g295(.A(new_n246), .B(new_n481), .C1(new_n240), .C2(G128), .ZN(new_n482));
  NAND3_X1  g296(.A1(new_n480), .A2(new_n244), .A3(new_n482), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n483), .A2(new_n417), .ZN(new_n484));
  INV_X1    g298(.A(KEYINPUT10), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n484), .A2(new_n485), .ZN(new_n486));
  AOI22_X1  g300(.A1(new_n238), .A2(new_n227), .B1(KEYINPUT1), .B2(new_n245), .ZN(new_n487));
  AOI21_X1  g301(.A(new_n485), .B1(new_n487), .B2(new_n244), .ZN(new_n488));
  NAND2_X1  g302(.A1(new_n417), .A2(new_n488), .ZN(new_n489));
  INV_X1    g303(.A(KEYINPUT80), .ZN(new_n490));
  NAND2_X1  g304(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  AND2_X1   g305(.A1(new_n256), .A2(new_n404), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n492), .A2(new_n433), .ZN(new_n493));
  NAND3_X1  g307(.A1(new_n417), .A2(new_n488), .A3(KEYINPUT80), .ZN(new_n494));
  NAND4_X1  g308(.A1(new_n486), .A2(new_n491), .A3(new_n493), .A4(new_n494), .ZN(new_n495));
  NOR2_X1   g309(.A1(new_n257), .A2(new_n258), .ZN(new_n496));
  INV_X1    g310(.A(new_n496), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n495), .A2(new_n497), .ZN(new_n498));
  AND3_X1   g312(.A1(new_n417), .A2(new_n488), .A3(KEYINPUT80), .ZN(new_n499));
  AOI21_X1  g313(.A(KEYINPUT80), .B1(new_n417), .B2(new_n488), .ZN(new_n500));
  NOR2_X1   g314(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  AOI22_X1  g315(.A1(new_n484), .A2(new_n485), .B1(new_n492), .B2(new_n433), .ZN(new_n502));
  NAND3_X1  g316(.A1(new_n501), .A2(new_n502), .A3(new_n496), .ZN(new_n503));
  XNOR2_X1  g317(.A(G110), .B(G140), .ZN(new_n504));
  INV_X1    g318(.A(G227), .ZN(new_n505));
  NOR2_X1   g319(.A1(new_n505), .A2(G953), .ZN(new_n506));
  XNOR2_X1  g320(.A(new_n504), .B(new_n506), .ZN(new_n507));
  INV_X1    g321(.A(new_n507), .ZN(new_n508));
  AND2_X1   g322(.A1(new_n503), .A2(new_n508), .ZN(new_n509));
  INV_X1    g323(.A(new_n247), .ZN(new_n510));
  NAND2_X1  g324(.A1(new_n454), .A2(new_n510), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n511), .A2(new_n484), .ZN(new_n512));
  AOI21_X1  g326(.A(KEYINPUT12), .B1(new_n512), .B2(new_n497), .ZN(new_n513));
  INV_X1    g327(.A(KEYINPUT12), .ZN(new_n514));
  AOI211_X1 g328(.A(new_n514), .B(new_n496), .C1(new_n511), .C2(new_n484), .ZN(new_n515));
  OAI21_X1  g329(.A(new_n503), .B1(new_n513), .B2(new_n515), .ZN(new_n516));
  AOI22_X1  g330(.A1(new_n498), .A2(new_n509), .B1(new_n516), .B2(new_n507), .ZN(new_n517));
  OAI21_X1  g331(.A(G469), .B1(new_n517), .B2(G902), .ZN(new_n518));
  INV_X1    g332(.A(G469), .ZN(new_n519));
  OAI211_X1 g333(.A(new_n503), .B(new_n508), .C1(new_n513), .C2(new_n515), .ZN(new_n520));
  INV_X1    g334(.A(new_n520), .ZN(new_n521));
  AOI21_X1  g335(.A(new_n508), .B1(new_n498), .B2(new_n503), .ZN(new_n522));
  OAI211_X1 g336(.A(new_n519), .B(new_n282), .C1(new_n521), .C2(new_n522), .ZN(new_n523));
  AOI21_X1  g337(.A(new_n477), .B1(new_n518), .B2(new_n523), .ZN(new_n524));
  OAI22_X1  g338(.A1(new_n324), .A2(new_n325), .B1(new_n316), .B2(new_n234), .ZN(new_n525));
  XNOR2_X1  g339(.A(KEYINPUT88), .B(G143), .ZN(new_n526));
  AND3_X1   g340(.A1(new_n188), .A2(new_n189), .A3(G214), .ZN(new_n527));
  NOR2_X1   g341(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  NAND3_X1  g342(.A1(new_n188), .A2(new_n189), .A3(G214), .ZN(new_n529));
  AOI21_X1  g343(.A(new_n529), .B1(KEYINPUT88), .B2(new_n236), .ZN(new_n530));
  OAI211_X1 g344(.A(KEYINPUT18), .B(G131), .C1(new_n528), .C2(new_n530), .ZN(new_n531));
  INV_X1    g345(.A(KEYINPUT88), .ZN(new_n532));
  OAI21_X1  g346(.A(new_n527), .B1(new_n532), .B2(G143), .ZN(new_n533));
  NAND2_X1  g347(.A1(KEYINPUT18), .A2(G131), .ZN(new_n534));
  OAI211_X1 g348(.A(new_n533), .B(new_n534), .C1(new_n527), .C2(new_n526), .ZN(new_n535));
  NAND3_X1  g349(.A1(new_n525), .A2(new_n531), .A3(new_n535), .ZN(new_n536));
  INV_X1    g350(.A(KEYINPUT89), .ZN(new_n537));
  NAND2_X1  g351(.A1(new_n536), .A2(new_n537), .ZN(new_n538));
  NAND4_X1  g352(.A1(new_n525), .A2(new_n531), .A3(KEYINPUT89), .A4(new_n535), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n538), .A2(new_n539), .ZN(new_n540));
  XNOR2_X1  g354(.A(G113), .B(G122), .ZN(new_n541));
  XNOR2_X1  g355(.A(new_n541), .B(new_n396), .ZN(new_n542));
  OAI21_X1  g356(.A(G131), .B1(new_n528), .B2(new_n530), .ZN(new_n543));
  INV_X1    g357(.A(KEYINPUT17), .ZN(new_n544));
  OR2_X1    g358(.A1(new_n543), .A2(new_n544), .ZN(new_n545));
  OAI211_X1 g359(.A(new_n533), .B(new_n251), .C1(new_n527), .C2(new_n526), .ZN(new_n546));
  NAND3_X1  g360(.A1(new_n546), .A2(new_n543), .A3(new_n544), .ZN(new_n547));
  NAND4_X1  g361(.A1(new_n545), .A2(new_n343), .A3(new_n319), .A4(new_n547), .ZN(new_n548));
  NAND3_X1  g362(.A1(new_n540), .A2(new_n542), .A3(new_n548), .ZN(new_n549));
  INV_X1    g363(.A(new_n549), .ZN(new_n550));
  OR2_X1    g364(.A1(new_n323), .A2(KEYINPUT19), .ZN(new_n551));
  INV_X1    g365(.A(KEYINPUT19), .ZN(new_n552));
  OAI21_X1  g366(.A(new_n551), .B1(new_n341), .B2(new_n552), .ZN(new_n553));
  AOI22_X1  g367(.A1(new_n234), .A2(new_n553), .B1(new_n546), .B2(new_n543), .ZN(new_n554));
  NAND3_X1  g368(.A1(new_n321), .A2(new_n322), .A3(new_n554), .ZN(new_n555));
  AOI21_X1  g369(.A(new_n542), .B1(new_n555), .B2(new_n540), .ZN(new_n556));
  NOR2_X1   g370(.A1(new_n550), .A2(new_n556), .ZN(new_n557));
  NOR2_X1   g371(.A1(G475), .A2(G902), .ZN(new_n558));
  INV_X1    g372(.A(new_n558), .ZN(new_n559));
  OAI21_X1  g373(.A(KEYINPUT20), .B1(new_n557), .B2(new_n559), .ZN(new_n560));
  INV_X1    g374(.A(KEYINPUT20), .ZN(new_n561));
  OAI211_X1 g375(.A(new_n561), .B(new_n558), .C1(new_n550), .C2(new_n556), .ZN(new_n562));
  AOI21_X1  g376(.A(new_n542), .B1(new_n540), .B2(new_n548), .ZN(new_n563));
  OAI21_X1  g377(.A(new_n282), .B1(new_n550), .B2(new_n563), .ZN(new_n564));
  AOI22_X1  g378(.A1(new_n560), .A2(new_n562), .B1(G475), .B2(new_n564), .ZN(new_n565));
  INV_X1    g379(.A(G122), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n566), .A2(G116), .ZN(new_n567));
  AOI21_X1  g381(.A(new_n399), .B1(new_n567), .B2(KEYINPUT14), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n199), .A2(G122), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n567), .A2(new_n569), .ZN(new_n570));
  OR2_X1    g384(.A1(new_n568), .A2(new_n570), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n568), .A2(new_n570), .ZN(new_n572));
  OAI21_X1  g386(.A(KEYINPUT90), .B1(new_n236), .B2(G128), .ZN(new_n573));
  INV_X1    g387(.A(KEYINPUT90), .ZN(new_n574));
  NAND3_X1  g388(.A1(new_n574), .A2(new_n227), .A3(G143), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n573), .A2(new_n575), .ZN(new_n576));
  XNOR2_X1  g390(.A(KEYINPUT65), .B(G134), .ZN(new_n577));
  NAND2_X1  g391(.A1(new_n236), .A2(G128), .ZN(new_n578));
  AND3_X1   g392(.A1(new_n576), .A2(new_n577), .A3(new_n578), .ZN(new_n579));
  AOI21_X1  g393(.A(new_n577), .B1(new_n576), .B2(new_n578), .ZN(new_n580));
  OAI211_X1 g394(.A(new_n571), .B(new_n572), .C1(new_n579), .C2(new_n580), .ZN(new_n581));
  AND2_X1   g395(.A1(new_n573), .A2(new_n575), .ZN(new_n582));
  INV_X1    g396(.A(KEYINPUT13), .ZN(new_n583));
  NAND2_X1  g397(.A1(new_n578), .A2(new_n583), .ZN(new_n584));
  NAND3_X1  g398(.A1(new_n236), .A2(KEYINPUT13), .A3(G128), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n584), .A2(new_n585), .ZN(new_n586));
  OAI21_X1  g400(.A(G134), .B1(new_n582), .B2(new_n586), .ZN(new_n587));
  XNOR2_X1  g401(.A(G116), .B(G122), .ZN(new_n588));
  XNOR2_X1  g402(.A(new_n588), .B(new_n399), .ZN(new_n589));
  NAND3_X1  g403(.A1(new_n576), .A2(new_n577), .A3(new_n578), .ZN(new_n590));
  NAND3_X1  g404(.A1(new_n587), .A2(new_n589), .A3(new_n590), .ZN(new_n591));
  NOR3_X1   g405(.A1(new_n475), .A2(new_n365), .A3(G953), .ZN(new_n592));
  NAND3_X1  g406(.A1(new_n581), .A2(new_n591), .A3(new_n592), .ZN(new_n593));
  INV_X1    g407(.A(KEYINPUT91), .ZN(new_n594));
  NAND2_X1  g408(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  NAND4_X1  g409(.A1(new_n581), .A2(new_n591), .A3(KEYINPUT91), .A4(new_n592), .ZN(new_n596));
  NAND2_X1  g410(.A1(new_n595), .A2(new_n596), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n581), .A2(new_n591), .ZN(new_n598));
  INV_X1    g412(.A(new_n592), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  NAND2_X1  g414(.A1(new_n600), .A2(KEYINPUT92), .ZN(new_n601));
  INV_X1    g415(.A(KEYINPUT92), .ZN(new_n602));
  NAND3_X1  g416(.A1(new_n598), .A2(new_n602), .A3(new_n599), .ZN(new_n603));
  NAND3_X1  g417(.A1(new_n597), .A2(new_n601), .A3(new_n603), .ZN(new_n604));
  INV_X1    g418(.A(G478), .ZN(new_n605));
  NOR2_X1   g419(.A1(KEYINPUT93), .A2(KEYINPUT15), .ZN(new_n606));
  INV_X1    g420(.A(new_n606), .ZN(new_n607));
  NAND2_X1  g421(.A1(KEYINPUT93), .A2(KEYINPUT15), .ZN(new_n608));
  AOI21_X1  g422(.A(new_n605), .B1(new_n607), .B2(new_n608), .ZN(new_n609));
  INV_X1    g423(.A(new_n609), .ZN(new_n610));
  NAND3_X1  g424(.A1(new_n604), .A2(new_n282), .A3(new_n610), .ZN(new_n611));
  INV_X1    g425(.A(new_n611), .ZN(new_n612));
  AOI21_X1  g426(.A(new_n610), .B1(new_n604), .B2(new_n282), .ZN(new_n613));
  NOR2_X1   g427(.A1(new_n612), .A2(new_n613), .ZN(new_n614));
  INV_X1    g428(.A(new_n614), .ZN(new_n615));
  INV_X1    g429(.A(G952), .ZN(new_n616));
  NOR2_X1   g430(.A1(new_n616), .A2(G953), .ZN(new_n617));
  NAND2_X1  g431(.A1(G234), .A2(G237), .ZN(new_n618));
  NAND2_X1  g432(.A1(new_n617), .A2(new_n618), .ZN(new_n619));
  XNOR2_X1  g433(.A(KEYINPUT21), .B(G898), .ZN(new_n620));
  INV_X1    g434(.A(new_n620), .ZN(new_n621));
  NAND3_X1  g435(.A1(new_n618), .A2(G902), .A3(G953), .ZN(new_n622));
  OAI21_X1  g436(.A(new_n619), .B1(new_n621), .B2(new_n622), .ZN(new_n623));
  XNOR2_X1  g437(.A(new_n623), .B(KEYINPUT94), .ZN(new_n624));
  INV_X1    g438(.A(new_n624), .ZN(new_n625));
  NOR2_X1   g439(.A1(new_n615), .A2(new_n625), .ZN(new_n626));
  AND4_X1   g440(.A1(new_n474), .A2(new_n524), .A3(new_n565), .A4(new_n626), .ZN(new_n627));
  NAND2_X1  g441(.A1(new_n389), .A2(new_n627), .ZN(new_n628));
  XNOR2_X1  g442(.A(new_n628), .B(G101), .ZN(G3));
  NAND3_X1  g443(.A1(new_n600), .A2(KEYINPUT33), .A3(new_n593), .ZN(new_n630));
  NOR2_X1   g444(.A1(new_n605), .A2(G902), .ZN(new_n631));
  INV_X1    g445(.A(KEYINPUT96), .ZN(new_n632));
  INV_X1    g446(.A(KEYINPUT33), .ZN(new_n633));
  AND3_X1   g447(.A1(new_n604), .A2(new_n632), .A3(new_n633), .ZN(new_n634));
  AOI21_X1  g448(.A(new_n632), .B1(new_n604), .B2(new_n633), .ZN(new_n635));
  OAI211_X1 g449(.A(new_n630), .B(new_n631), .C1(new_n634), .C2(new_n635), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n604), .A2(new_n282), .ZN(new_n637));
  XNOR2_X1  g451(.A(KEYINPUT97), .B(G478), .ZN(new_n638));
  NAND2_X1  g452(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  NAND2_X1  g453(.A1(new_n636), .A2(new_n639), .ZN(new_n640));
  NAND2_X1  g454(.A1(new_n564), .A2(G475), .ZN(new_n641));
  AND2_X1   g455(.A1(new_n555), .A2(new_n540), .ZN(new_n642));
  OAI21_X1  g456(.A(new_n549), .B1(new_n642), .B2(new_n542), .ZN(new_n643));
  AOI21_X1  g457(.A(new_n561), .B1(new_n643), .B2(new_n558), .ZN(new_n644));
  INV_X1    g458(.A(new_n562), .ZN(new_n645));
  OAI21_X1  g459(.A(new_n641), .B1(new_n644), .B2(new_n645), .ZN(new_n646));
  AND3_X1   g460(.A1(new_n640), .A2(new_n646), .A3(new_n624), .ZN(new_n647));
  INV_X1    g461(.A(KEYINPUT95), .ZN(new_n648));
  NAND3_X1  g462(.A1(new_n466), .A2(new_n648), .A3(new_n473), .ZN(new_n649));
  AOI21_X1  g463(.A(new_n392), .B1(new_n470), .B2(new_n472), .ZN(new_n650));
  AOI21_X1  g464(.A(new_n391), .B1(new_n650), .B2(KEYINPUT95), .ZN(new_n651));
  NAND3_X1  g465(.A1(new_n647), .A2(new_n649), .A3(new_n651), .ZN(new_n652));
  INV_X1    g466(.A(KEYINPUT98), .ZN(new_n653));
  NAND2_X1  g467(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  NAND4_X1  g468(.A1(new_n647), .A2(new_n651), .A3(KEYINPUT98), .A4(new_n649), .ZN(new_n655));
  NAND2_X1  g469(.A1(new_n654), .A2(new_n655), .ZN(new_n656));
  INV_X1    g470(.A(new_n524), .ZN(new_n657));
  AOI21_X1  g471(.A(new_n187), .B1(new_n296), .B2(new_n282), .ZN(new_n658));
  INV_X1    g472(.A(new_n658), .ZN(new_n659));
  NAND2_X1  g473(.A1(new_n659), .A2(new_n298), .ZN(new_n660));
  NOR3_X1   g474(.A1(new_n657), .A2(new_n371), .A3(new_n660), .ZN(new_n661));
  NAND2_X1  g475(.A1(new_n656), .A2(new_n661), .ZN(new_n662));
  XOR2_X1   g476(.A(KEYINPUT34), .B(G104), .Z(new_n663));
  XNOR2_X1  g477(.A(new_n662), .B(new_n663), .ZN(G6));
  AND2_X1   g478(.A1(new_n651), .A2(new_n649), .ZN(new_n665));
  NOR3_X1   g479(.A1(new_n646), .A2(new_n614), .A3(new_n625), .ZN(new_n666));
  NAND3_X1  g480(.A1(new_n661), .A2(new_n665), .A3(new_n666), .ZN(new_n667));
  XNOR2_X1  g481(.A(new_n667), .B(KEYINPUT99), .ZN(new_n668));
  XNOR2_X1  g482(.A(KEYINPUT35), .B(G107), .ZN(new_n669));
  XNOR2_X1  g483(.A(new_n668), .B(new_n669), .ZN(G9));
  INV_X1    g484(.A(KEYINPUT100), .ZN(new_n671));
  NOR2_X1   g485(.A1(new_n357), .A2(KEYINPUT36), .ZN(new_n672));
  XNOR2_X1  g486(.A(new_n353), .B(new_n672), .ZN(new_n673));
  NAND2_X1  g487(.A1(new_n673), .A2(new_n385), .ZN(new_n674));
  NAND3_X1  g488(.A1(new_n367), .A2(new_n671), .A3(new_n674), .ZN(new_n675));
  INV_X1    g489(.A(new_n674), .ZN(new_n676));
  OAI21_X1  g490(.A(KEYINPUT100), .B1(new_n384), .B2(new_n676), .ZN(new_n677));
  NAND2_X1  g491(.A1(new_n675), .A2(new_n677), .ZN(new_n678));
  NOR2_X1   g492(.A1(new_n678), .A2(new_n660), .ZN(new_n679));
  NAND2_X1  g493(.A1(new_n627), .A2(new_n679), .ZN(new_n680));
  XOR2_X1   g494(.A(KEYINPUT37), .B(G110), .Z(new_n681));
  XNOR2_X1  g495(.A(new_n681), .B(KEYINPUT101), .ZN(new_n682));
  XNOR2_X1  g496(.A(new_n680), .B(new_n682), .ZN(G12));
  INV_X1    g497(.A(new_n678), .ZN(new_n684));
  INV_X1    g498(.A(new_n619), .ZN(new_n685));
  INV_X1    g499(.A(new_n622), .ZN(new_n686));
  XNOR2_X1  g500(.A(KEYINPUT102), .B(G900), .ZN(new_n687));
  AOI21_X1  g501(.A(new_n685), .B1(new_n686), .B2(new_n687), .ZN(new_n688));
  NOR3_X1   g502(.A1(new_n646), .A2(new_n614), .A3(new_n688), .ZN(new_n689));
  NAND3_X1  g503(.A1(new_n684), .A2(new_n381), .A3(new_n689), .ZN(new_n690));
  AND3_X1   g504(.A1(new_n651), .A2(new_n649), .A3(new_n524), .ZN(new_n691));
  INV_X1    g505(.A(new_n691), .ZN(new_n692));
  NOR2_X1   g506(.A1(new_n690), .A2(new_n692), .ZN(new_n693));
  XNOR2_X1  g507(.A(new_n693), .B(new_n227), .ZN(G30));
  XOR2_X1   g508(.A(new_n688), .B(KEYINPUT39), .Z(new_n695));
  NAND2_X1  g509(.A1(new_n524), .A2(new_n695), .ZN(new_n696));
  XNOR2_X1  g510(.A(new_n696), .B(KEYINPUT40), .ZN(new_n697));
  NOR4_X1   g511(.A1(new_n697), .A2(new_n391), .A3(new_n565), .A4(new_n614), .ZN(new_n698));
  NAND2_X1  g512(.A1(new_n367), .A2(new_n674), .ZN(new_n699));
  NAND2_X1  g513(.A1(new_n304), .A2(new_n300), .ZN(new_n700));
  NAND2_X1  g514(.A1(new_n290), .A2(new_n264), .ZN(new_n701));
  NAND2_X1  g515(.A1(new_n701), .A2(new_n193), .ZN(new_n702));
  NAND3_X1  g516(.A1(new_n274), .A2(new_n264), .A3(new_n194), .ZN(new_n703));
  NAND2_X1  g517(.A1(new_n703), .A2(new_n282), .ZN(new_n704));
  INV_X1    g518(.A(new_n704), .ZN(new_n705));
  AOI21_X1  g519(.A(new_n187), .B1(new_n702), .B2(new_n705), .ZN(new_n706));
  INV_X1    g520(.A(new_n706), .ZN(new_n707));
  AOI21_X1  g521(.A(new_n699), .B1(new_n700), .B2(new_n707), .ZN(new_n708));
  NAND2_X1  g522(.A1(new_n466), .A2(new_n473), .ZN(new_n709));
  XNOR2_X1  g523(.A(new_n709), .B(KEYINPUT38), .ZN(new_n710));
  AND3_X1   g524(.A1(new_n698), .A2(new_n708), .A3(new_n710), .ZN(new_n711));
  XNOR2_X1  g525(.A(new_n711), .B(new_n236), .ZN(G45));
  INV_X1    g526(.A(new_n688), .ZN(new_n713));
  NAND3_X1  g527(.A1(new_n640), .A2(new_n646), .A3(new_n713), .ZN(new_n714));
  INV_X1    g528(.A(new_n714), .ZN(new_n715));
  NAND3_X1  g529(.A1(new_n684), .A2(new_n381), .A3(new_n715), .ZN(new_n716));
  NOR2_X1   g530(.A1(new_n716), .A2(new_n692), .ZN(new_n717));
  XNOR2_X1  g531(.A(new_n717), .B(new_n234), .ZN(G48));
  NOR2_X1   g532(.A1(new_n495), .A2(new_n497), .ZN(new_n719));
  AOI21_X1  g533(.A(new_n496), .B1(new_n501), .B2(new_n502), .ZN(new_n720));
  OAI21_X1  g534(.A(new_n507), .B1(new_n719), .B2(new_n720), .ZN(new_n721));
  NAND2_X1  g535(.A1(new_n721), .A2(new_n520), .ZN(new_n722));
  AOI21_X1  g536(.A(new_n519), .B1(new_n722), .B2(new_n282), .ZN(new_n723));
  AOI211_X1 g537(.A(G469), .B(G902), .C1(new_n721), .C2(new_n520), .ZN(new_n724));
  NOR3_X1   g538(.A1(new_n723), .A2(new_n724), .A3(new_n477), .ZN(new_n725));
  INV_X1    g539(.A(new_n725), .ZN(new_n726));
  NOR3_X1   g540(.A1(new_n305), .A2(new_n371), .A3(new_n726), .ZN(new_n727));
  NAND2_X1  g541(.A1(new_n656), .A2(new_n727), .ZN(new_n728));
  XNOR2_X1  g542(.A(KEYINPUT41), .B(G113), .ZN(new_n729));
  XNOR2_X1  g543(.A(new_n728), .B(new_n729), .ZN(G15));
  AOI21_X1  g544(.A(new_n371), .B1(new_n700), .B2(new_n376), .ZN(new_n731));
  NAND4_X1  g545(.A1(new_n731), .A2(new_n665), .A3(new_n666), .A4(new_n725), .ZN(new_n732));
  XNOR2_X1  g546(.A(new_n732), .B(G116), .ZN(G18));
  NAND3_X1  g547(.A1(new_n651), .A2(new_n649), .A3(new_n725), .ZN(new_n734));
  NAND2_X1  g548(.A1(new_n734), .A2(KEYINPUT103), .ZN(new_n735));
  INV_X1    g549(.A(KEYINPUT103), .ZN(new_n736));
  NAND4_X1  g550(.A1(new_n651), .A2(new_n649), .A3(new_n725), .A4(new_n736), .ZN(new_n737));
  NAND2_X1  g551(.A1(new_n735), .A2(new_n737), .ZN(new_n738));
  NAND2_X1  g552(.A1(new_n626), .A2(new_n565), .ZN(new_n739));
  INV_X1    g553(.A(new_n739), .ZN(new_n740));
  AOI21_X1  g554(.A(new_n678), .B1(new_n376), .B2(new_n700), .ZN(new_n741));
  NAND3_X1  g555(.A1(new_n738), .A2(new_n740), .A3(new_n741), .ZN(new_n742));
  XNOR2_X1  g556(.A(new_n742), .B(G119), .ZN(G21));
  NOR2_X1   g557(.A1(new_n565), .A2(new_n614), .ZN(new_n744));
  AND3_X1   g558(.A1(new_n651), .A2(new_n649), .A3(new_n744), .ZN(new_n745));
  INV_X1    g559(.A(new_n297), .ZN(new_n746));
  AND2_X1   g560(.A1(new_n292), .A2(new_n295), .ZN(new_n747));
  NAND2_X1  g561(.A1(new_n277), .A2(new_n279), .ZN(new_n748));
  NAND2_X1  g562(.A1(new_n748), .A2(new_n194), .ZN(new_n749));
  AOI21_X1  g563(.A(new_n746), .B1(new_n747), .B2(new_n749), .ZN(new_n750));
  NOR2_X1   g564(.A1(new_n750), .A2(new_n658), .ZN(new_n751));
  AND4_X1   g565(.A1(new_n387), .A2(new_n725), .A3(new_n624), .A4(new_n751), .ZN(new_n752));
  NAND2_X1  g566(.A1(new_n745), .A2(new_n752), .ZN(new_n753));
  XNOR2_X1  g567(.A(new_n753), .B(G122), .ZN(G24));
  AND2_X1   g568(.A1(new_n751), .A2(new_n699), .ZN(new_n755));
  NAND2_X1  g569(.A1(new_n714), .A2(KEYINPUT104), .ZN(new_n756));
  INV_X1    g570(.A(KEYINPUT104), .ZN(new_n757));
  NAND4_X1  g571(.A1(new_n640), .A2(new_n757), .A3(new_n646), .A4(new_n713), .ZN(new_n758));
  NAND3_X1  g572(.A1(new_n755), .A2(new_n756), .A3(new_n758), .ZN(new_n759));
  AOI21_X1  g573(.A(new_n759), .B1(new_n735), .B2(new_n737), .ZN(new_n760));
  XNOR2_X1  g574(.A(new_n760), .B(new_n310), .ZN(G27));
  NAND2_X1  g575(.A1(new_n516), .A2(new_n507), .ZN(new_n762));
  NAND3_X1  g576(.A1(new_n498), .A2(new_n503), .A3(new_n508), .ZN(new_n763));
  NAND3_X1  g577(.A1(new_n762), .A2(G469), .A3(new_n763), .ZN(new_n764));
  NAND2_X1  g578(.A1(G469), .A2(G902), .ZN(new_n765));
  NAND2_X1  g579(.A1(new_n764), .A2(new_n765), .ZN(new_n766));
  OAI21_X1  g580(.A(KEYINPUT105), .B1(new_n766), .B2(new_n724), .ZN(new_n767));
  INV_X1    g581(.A(KEYINPUT105), .ZN(new_n768));
  NAND4_X1  g582(.A1(new_n523), .A2(new_n768), .A3(new_n765), .A4(new_n764), .ZN(new_n769));
  NAND3_X1  g583(.A1(new_n767), .A2(new_n476), .A3(new_n769), .ZN(new_n770));
  INV_X1    g584(.A(new_n770), .ZN(new_n771));
  NAND3_X1  g585(.A1(new_n466), .A2(new_n390), .A3(new_n473), .ZN(new_n772));
  INV_X1    g586(.A(new_n772), .ZN(new_n773));
  NAND4_X1  g587(.A1(new_n771), .A2(new_n756), .A3(new_n758), .A4(new_n773), .ZN(new_n774));
  OR2_X1    g588(.A1(new_n378), .A2(KEYINPUT106), .ZN(new_n775));
  NAND2_X1  g589(.A1(new_n378), .A2(KEYINPUT106), .ZN(new_n776));
  NAND3_X1  g590(.A1(new_n775), .A2(new_n303), .A3(new_n776), .ZN(new_n777));
  OAI21_X1  g591(.A(new_n387), .B1(new_n777), .B2(new_n287), .ZN(new_n778));
  OAI21_X1  g592(.A(KEYINPUT42), .B1(new_n774), .B2(new_n778), .ZN(new_n779));
  AND2_X1   g593(.A1(new_n756), .A2(new_n758), .ZN(new_n780));
  INV_X1    g594(.A(KEYINPUT42), .ZN(new_n781));
  NOR2_X1   g595(.A1(new_n770), .A2(new_n772), .ZN(new_n782));
  NAND4_X1  g596(.A1(new_n780), .A2(new_n781), .A3(new_n731), .A4(new_n782), .ZN(new_n783));
  NAND2_X1  g597(.A1(new_n779), .A2(new_n783), .ZN(new_n784));
  XNOR2_X1  g598(.A(new_n784), .B(new_n251), .ZN(G33));
  NAND3_X1  g599(.A1(new_n731), .A2(new_n689), .A3(new_n782), .ZN(new_n786));
  XNOR2_X1  g600(.A(new_n786), .B(G134), .ZN(G36));
  NAND2_X1  g601(.A1(new_n762), .A2(new_n763), .ZN(new_n788));
  INV_X1    g602(.A(KEYINPUT45), .ZN(new_n789));
  AOI21_X1  g603(.A(new_n519), .B1(new_n788), .B2(new_n789), .ZN(new_n790));
  OAI21_X1  g604(.A(new_n790), .B1(new_n789), .B2(new_n788), .ZN(new_n791));
  AND2_X1   g605(.A1(new_n791), .A2(new_n765), .ZN(new_n792));
  OR2_X1    g606(.A1(new_n792), .A2(KEYINPUT46), .ZN(new_n793));
  NAND2_X1  g607(.A1(new_n792), .A2(KEYINPUT46), .ZN(new_n794));
  NAND3_X1  g608(.A1(new_n793), .A2(new_n523), .A3(new_n794), .ZN(new_n795));
  NAND3_X1  g609(.A1(new_n795), .A2(new_n476), .A3(new_n695), .ZN(new_n796));
  XNOR2_X1  g610(.A(new_n796), .B(KEYINPUT107), .ZN(new_n797));
  AOI21_X1  g611(.A(new_n646), .B1(new_n639), .B2(new_n636), .ZN(new_n798));
  XNOR2_X1  g612(.A(new_n798), .B(KEYINPUT43), .ZN(new_n799));
  NAND3_X1  g613(.A1(new_n799), .A2(new_n660), .A3(new_n699), .ZN(new_n800));
  INV_X1    g614(.A(KEYINPUT44), .ZN(new_n801));
  AOI21_X1  g615(.A(new_n772), .B1(new_n800), .B2(new_n801), .ZN(new_n802));
  OAI211_X1 g616(.A(new_n797), .B(new_n802), .C1(new_n801), .C2(new_n800), .ZN(new_n803));
  XNOR2_X1  g617(.A(new_n803), .B(G137), .ZN(G39));
  NAND2_X1  g618(.A1(new_n795), .A2(new_n476), .ZN(new_n805));
  INV_X1    g619(.A(KEYINPUT47), .ZN(new_n806));
  NAND2_X1  g620(.A1(new_n805), .A2(new_n806), .ZN(new_n807));
  NAND3_X1  g621(.A1(new_n795), .A2(KEYINPUT47), .A3(new_n476), .ZN(new_n808));
  NAND2_X1  g622(.A1(new_n807), .A2(new_n808), .ZN(new_n809));
  NOR3_X1   g623(.A1(new_n772), .A2(new_n714), .A3(new_n387), .ZN(new_n810));
  NAND3_X1  g624(.A1(new_n809), .A2(new_n305), .A3(new_n810), .ZN(new_n811));
  XNOR2_X1  g625(.A(new_n811), .B(G140), .ZN(G42));
  XOR2_X1   g626(.A(KEYINPUT112), .B(KEYINPUT53), .Z(new_n813));
  NAND4_X1  g627(.A1(new_n767), .A2(new_n476), .A3(new_n713), .A4(new_n769), .ZN(new_n814));
  INV_X1    g628(.A(new_n814), .ZN(new_n815));
  AND4_X1   g629(.A1(KEYINPUT111), .A2(new_n708), .A3(new_n745), .A4(new_n815), .ZN(new_n816));
  AOI21_X1  g630(.A(new_n706), .B1(new_n304), .B2(new_n300), .ZN(new_n817));
  NOR3_X1   g631(.A1(new_n817), .A2(new_n814), .A3(new_n699), .ZN(new_n818));
  AOI21_X1  g632(.A(KEYINPUT111), .B1(new_n818), .B2(new_n745), .ZN(new_n819));
  NOR2_X1   g633(.A1(new_n816), .A2(new_n819), .ZN(new_n820));
  AND3_X1   g634(.A1(new_n755), .A2(new_n756), .A3(new_n758), .ZN(new_n821));
  NAND2_X1  g635(.A1(new_n738), .A2(new_n821), .ZN(new_n822));
  OAI211_X1 g636(.A(new_n741), .B(new_n691), .C1(new_n689), .C2(new_n715), .ZN(new_n823));
  NAND2_X1  g637(.A1(new_n822), .A2(new_n823), .ZN(new_n824));
  OAI21_X1  g638(.A(KEYINPUT52), .B1(new_n820), .B2(new_n824), .ZN(new_n825));
  NAND3_X1  g639(.A1(new_n708), .A2(new_n745), .A3(new_n815), .ZN(new_n826));
  INV_X1    g640(.A(KEYINPUT111), .ZN(new_n827));
  NAND2_X1  g641(.A1(new_n826), .A2(new_n827), .ZN(new_n828));
  NAND3_X1  g642(.A1(new_n818), .A2(KEYINPUT111), .A3(new_n745), .ZN(new_n829));
  NAND2_X1  g643(.A1(new_n828), .A2(new_n829), .ZN(new_n830));
  INV_X1    g644(.A(KEYINPUT52), .ZN(new_n831));
  NAND4_X1  g645(.A1(new_n830), .A2(new_n831), .A3(new_n822), .A4(new_n823), .ZN(new_n832));
  NAND2_X1  g646(.A1(new_n825), .A2(new_n832), .ZN(new_n833));
  AND3_X1   g647(.A1(new_n628), .A2(new_n728), .A3(new_n742), .ZN(new_n834));
  INV_X1    g648(.A(new_n613), .ZN(new_n835));
  NAND3_X1  g649(.A1(new_n835), .A2(new_n611), .A3(new_n713), .ZN(new_n836));
  OAI21_X1  g650(.A(KEYINPUT109), .B1(new_n646), .B2(new_n836), .ZN(new_n837));
  NOR3_X1   g651(.A1(new_n612), .A2(new_n613), .A3(new_n688), .ZN(new_n838));
  INV_X1    g652(.A(KEYINPUT109), .ZN(new_n839));
  NAND3_X1  g653(.A1(new_n565), .A2(new_n838), .A3(new_n839), .ZN(new_n840));
  NAND3_X1  g654(.A1(new_n837), .A2(new_n840), .A3(new_n524), .ZN(new_n841));
  NOR2_X1   g655(.A1(new_n841), .A2(new_n772), .ZN(new_n842));
  NAND2_X1  g656(.A1(new_n741), .A2(new_n842), .ZN(new_n843));
  INV_X1    g657(.A(new_n782), .ZN(new_n844));
  OAI211_X1 g658(.A(new_n843), .B(new_n786), .C1(new_n759), .C2(new_n844), .ZN(new_n845));
  NOR2_X1   g659(.A1(new_n784), .A2(new_n845), .ZN(new_n846));
  AOI22_X1  g660(.A1(new_n627), .A2(new_n679), .B1(new_n745), .B2(new_n752), .ZN(new_n847));
  INV_X1    g661(.A(KEYINPUT108), .ZN(new_n848));
  OR2_X1    g662(.A1(new_n474), .A2(new_n848), .ZN(new_n849));
  NOR2_X1   g663(.A1(new_n646), .A2(new_n614), .ZN(new_n850));
  NAND2_X1  g664(.A1(new_n850), .A2(new_n624), .ZN(new_n851));
  AOI21_X1  g665(.A(new_n851), .B1(new_n474), .B2(new_n848), .ZN(new_n852));
  NAND3_X1  g666(.A1(new_n640), .A2(new_n646), .A3(new_n624), .ZN(new_n853));
  OAI21_X1  g667(.A(new_n853), .B1(new_n666), .B2(KEYINPUT108), .ZN(new_n854));
  OAI211_X1 g668(.A(new_n849), .B(new_n661), .C1(new_n852), .C2(new_n854), .ZN(new_n855));
  AND3_X1   g669(.A1(new_n847), .A2(new_n855), .A3(new_n732), .ZN(new_n856));
  NAND3_X1  g670(.A1(new_n834), .A2(new_n846), .A3(new_n856), .ZN(new_n857));
  OAI21_X1  g671(.A(new_n813), .B1(new_n833), .B2(new_n857), .ZN(new_n858));
  INV_X1    g672(.A(KEYINPUT54), .ZN(new_n859));
  NAND3_X1  g673(.A1(new_n628), .A2(new_n728), .A3(new_n742), .ZN(new_n860));
  AOI22_X1  g674(.A1(new_n821), .A2(new_n782), .B1(new_n741), .B2(new_n842), .ZN(new_n861));
  NAND4_X1  g675(.A1(new_n861), .A2(new_n779), .A3(new_n783), .A4(new_n786), .ZN(new_n862));
  NAND3_X1  g676(.A1(new_n847), .A2(new_n855), .A3(new_n732), .ZN(new_n863));
  NOR3_X1   g677(.A1(new_n860), .A2(new_n862), .A3(new_n863), .ZN(new_n864));
  NAND4_X1  g678(.A1(new_n864), .A2(KEYINPUT53), .A3(new_n832), .A4(new_n825), .ZN(new_n865));
  NAND3_X1  g679(.A1(new_n858), .A2(new_n859), .A3(new_n865), .ZN(new_n866));
  NAND2_X1  g680(.A1(new_n866), .A2(KEYINPUT113), .ZN(new_n867));
  INV_X1    g681(.A(KEYINPUT113), .ZN(new_n868));
  NAND4_X1  g682(.A1(new_n858), .A2(new_n865), .A3(new_n868), .A4(new_n859), .ZN(new_n869));
  INV_X1    g683(.A(KEYINPUT110), .ZN(new_n870));
  NAND2_X1  g684(.A1(new_n857), .A2(new_n870), .ZN(new_n871));
  AND2_X1   g685(.A1(new_n825), .A2(new_n832), .ZN(new_n872));
  NOR2_X1   g686(.A1(new_n860), .A2(new_n863), .ZN(new_n873));
  NAND3_X1  g687(.A1(new_n873), .A2(KEYINPUT110), .A3(new_n846), .ZN(new_n874));
  NAND3_X1  g688(.A1(new_n871), .A2(new_n872), .A3(new_n874), .ZN(new_n875));
  INV_X1    g689(.A(KEYINPUT53), .ZN(new_n876));
  NOR2_X1   g690(.A1(new_n833), .A2(new_n857), .ZN(new_n877));
  INV_X1    g691(.A(new_n813), .ZN(new_n878));
  AOI22_X1  g692(.A1(new_n875), .A2(new_n876), .B1(new_n877), .B2(new_n878), .ZN(new_n879));
  OAI211_X1 g693(.A(new_n867), .B(new_n869), .C1(new_n879), .C2(new_n859), .ZN(new_n880));
  NOR2_X1   g694(.A1(new_n723), .A2(new_n724), .ZN(new_n881));
  INV_X1    g695(.A(new_n881), .ZN(new_n882));
  OAI211_X1 g696(.A(new_n807), .B(new_n808), .C1(new_n476), .C2(new_n882), .ZN(new_n883));
  AND3_X1   g697(.A1(new_n387), .A2(new_n685), .A3(new_n751), .ZN(new_n884));
  NAND2_X1  g698(.A1(new_n799), .A2(new_n884), .ZN(new_n885));
  NOR2_X1   g699(.A1(new_n885), .A2(new_n772), .ZN(new_n886));
  NAND2_X1  g700(.A1(new_n773), .A2(new_n725), .ZN(new_n887));
  OR2_X1    g701(.A1(new_n887), .A2(KEYINPUT114), .ZN(new_n888));
  AOI21_X1  g702(.A(new_n619), .B1(new_n887), .B2(KEYINPUT114), .ZN(new_n889));
  AND4_X1   g703(.A1(new_n387), .A2(new_n888), .A3(new_n817), .A4(new_n889), .ZN(new_n890));
  NOR2_X1   g704(.A1(new_n640), .A2(new_n646), .ZN(new_n891));
  AOI22_X1  g705(.A1(new_n883), .A2(new_n886), .B1(new_n890), .B2(new_n891), .ZN(new_n892));
  INV_X1    g706(.A(new_n885), .ZN(new_n893));
  NOR3_X1   g707(.A1(new_n710), .A2(new_n390), .A3(new_n726), .ZN(new_n894));
  NAND2_X1  g708(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  OR2_X1    g709(.A1(new_n895), .A2(KEYINPUT50), .ZN(new_n896));
  NAND4_X1  g710(.A1(new_n888), .A2(new_n799), .A3(new_n755), .A4(new_n889), .ZN(new_n897));
  NAND2_X1  g711(.A1(new_n895), .A2(KEYINPUT50), .ZN(new_n898));
  NAND3_X1  g712(.A1(new_n896), .A2(new_n897), .A3(new_n898), .ZN(new_n899));
  INV_X1    g713(.A(new_n899), .ZN(new_n900));
  AND3_X1   g714(.A1(new_n892), .A2(new_n900), .A3(KEYINPUT51), .ZN(new_n901));
  AOI21_X1  g715(.A(KEYINPUT51), .B1(new_n892), .B2(new_n900), .ZN(new_n902));
  INV_X1    g716(.A(new_n778), .ZN(new_n903));
  AND4_X1   g717(.A1(new_n903), .A2(new_n888), .A3(new_n799), .A4(new_n889), .ZN(new_n904));
  INV_X1    g718(.A(KEYINPUT48), .ZN(new_n905));
  XNOR2_X1  g719(.A(new_n904), .B(new_n905), .ZN(new_n906));
  NAND3_X1  g720(.A1(new_n890), .A2(new_n646), .A3(new_n640), .ZN(new_n907));
  NAND2_X1  g721(.A1(new_n893), .A2(new_n738), .ZN(new_n908));
  NAND4_X1  g722(.A1(new_n906), .A2(new_n617), .A3(new_n907), .A4(new_n908), .ZN(new_n909));
  OR3_X1    g723(.A1(new_n901), .A2(new_n902), .A3(new_n909), .ZN(new_n910));
  OAI21_X1  g724(.A(KEYINPUT115), .B1(new_n880), .B2(new_n910), .ZN(new_n911));
  AND2_X1   g725(.A1(new_n867), .A2(new_n869), .ZN(new_n912));
  INV_X1    g726(.A(KEYINPUT115), .ZN(new_n913));
  NAND2_X1  g727(.A1(new_n875), .A2(new_n876), .ZN(new_n914));
  NAND2_X1  g728(.A1(new_n877), .A2(new_n878), .ZN(new_n915));
  NAND2_X1  g729(.A1(new_n914), .A2(new_n915), .ZN(new_n916));
  NAND2_X1  g730(.A1(new_n916), .A2(KEYINPUT54), .ZN(new_n917));
  NOR3_X1   g731(.A1(new_n901), .A2(new_n902), .A3(new_n909), .ZN(new_n918));
  NAND4_X1  g732(.A1(new_n912), .A2(new_n913), .A3(new_n917), .A4(new_n918), .ZN(new_n919));
  NAND2_X1  g733(.A1(new_n616), .A2(new_n189), .ZN(new_n920));
  NAND3_X1  g734(.A1(new_n911), .A2(new_n919), .A3(new_n920), .ZN(new_n921));
  OR2_X1    g735(.A1(new_n882), .A2(KEYINPUT49), .ZN(new_n922));
  NAND2_X1  g736(.A1(new_n882), .A2(KEYINPUT49), .ZN(new_n923));
  AND3_X1   g737(.A1(new_n922), .A2(new_n798), .A3(new_n923), .ZN(new_n924));
  INV_X1    g738(.A(new_n710), .ZN(new_n925));
  NOR3_X1   g739(.A1(new_n371), .A2(new_n391), .A3(new_n477), .ZN(new_n926));
  NAND4_X1  g740(.A1(new_n924), .A2(new_n925), .A3(new_n817), .A4(new_n926), .ZN(new_n927));
  NAND2_X1  g741(.A1(new_n921), .A2(new_n927), .ZN(G75));
  AOI21_X1  g742(.A(new_n282), .B1(new_n858), .B2(new_n865), .ZN(new_n929));
  INV_X1    g743(.A(KEYINPUT117), .ZN(new_n930));
  NAND3_X1  g744(.A1(new_n929), .A2(new_n930), .A3(G210), .ZN(new_n931));
  INV_X1    g745(.A(KEYINPUT56), .ZN(new_n932));
  NAND2_X1  g746(.A1(new_n467), .A2(new_n469), .ZN(new_n933));
  NAND2_X1  g747(.A1(new_n933), .A2(new_n432), .ZN(new_n934));
  NAND2_X1  g748(.A1(new_n934), .A2(new_n470), .ZN(new_n935));
  XNOR2_X1  g749(.A(KEYINPUT116), .B(KEYINPUT55), .ZN(new_n936));
  XNOR2_X1  g750(.A(new_n935), .B(new_n936), .ZN(new_n937));
  NAND3_X1  g751(.A1(new_n931), .A2(new_n932), .A3(new_n937), .ZN(new_n938));
  AOI21_X1  g752(.A(new_n930), .B1(new_n929), .B2(G210), .ZN(new_n939));
  NOR2_X1   g753(.A1(new_n938), .A2(new_n939), .ZN(new_n940));
  NOR2_X1   g754(.A1(new_n189), .A2(G952), .ZN(new_n941));
  INV_X1    g755(.A(new_n941), .ZN(new_n942));
  AOI21_X1  g756(.A(KEYINPUT56), .B1(new_n929), .B2(G210), .ZN(new_n943));
  OAI21_X1  g757(.A(new_n942), .B1(new_n943), .B2(new_n937), .ZN(new_n944));
  NOR2_X1   g758(.A1(new_n940), .A2(new_n944), .ZN(G51));
  XOR2_X1   g759(.A(new_n765), .B(KEYINPUT57), .Z(new_n946));
  AND3_X1   g760(.A1(new_n858), .A2(new_n859), .A3(new_n865), .ZN(new_n947));
  AOI21_X1  g761(.A(new_n859), .B1(new_n858), .B2(new_n865), .ZN(new_n948));
  OAI21_X1  g762(.A(new_n946), .B1(new_n947), .B2(new_n948), .ZN(new_n949));
  NAND2_X1  g763(.A1(new_n949), .A2(new_n722), .ZN(new_n950));
  OR2_X1    g764(.A1(new_n950), .A2(KEYINPUT118), .ZN(new_n951));
  XOR2_X1   g765(.A(new_n791), .B(KEYINPUT119), .Z(new_n952));
  AOI22_X1  g766(.A1(new_n950), .A2(KEYINPUT118), .B1(new_n929), .B2(new_n952), .ZN(new_n953));
  AOI21_X1  g767(.A(new_n941), .B1(new_n951), .B2(new_n953), .ZN(G54));
  NAND3_X1  g768(.A1(new_n929), .A2(KEYINPUT58), .A3(G475), .ZN(new_n955));
  AND2_X1   g769(.A1(new_n955), .A2(new_n557), .ZN(new_n956));
  NOR2_X1   g770(.A1(new_n955), .A2(new_n557), .ZN(new_n957));
  NOR3_X1   g771(.A1(new_n956), .A2(new_n957), .A3(new_n941), .ZN(G60));
  OR2_X1    g772(.A1(new_n634), .A2(new_n635), .ZN(new_n959));
  AND2_X1   g773(.A1(new_n959), .A2(new_n630), .ZN(new_n960));
  NAND2_X1  g774(.A1(G478), .A2(G902), .ZN(new_n961));
  XNOR2_X1  g775(.A(new_n961), .B(KEYINPUT59), .ZN(new_n962));
  AOI21_X1  g776(.A(new_n960), .B1(new_n880), .B2(new_n962), .ZN(new_n963));
  OAI211_X1 g777(.A(new_n960), .B(new_n962), .C1(new_n947), .C2(new_n948), .ZN(new_n964));
  INV_X1    g778(.A(KEYINPUT120), .ZN(new_n965));
  AND3_X1   g779(.A1(new_n964), .A2(new_n965), .A3(new_n942), .ZN(new_n966));
  AOI21_X1  g780(.A(new_n965), .B1(new_n964), .B2(new_n942), .ZN(new_n967));
  NOR3_X1   g781(.A1(new_n963), .A2(new_n966), .A3(new_n967), .ZN(G63));
  NAND2_X1  g782(.A1(new_n858), .A2(new_n865), .ZN(new_n969));
  NAND2_X1  g783(.A1(G217), .A2(G902), .ZN(new_n970));
  XNOR2_X1  g784(.A(new_n970), .B(KEYINPUT121), .ZN(new_n971));
  XNOR2_X1  g785(.A(new_n971), .B(KEYINPUT60), .ZN(new_n972));
  NAND3_X1  g786(.A1(new_n969), .A2(new_n673), .A3(new_n972), .ZN(new_n973));
  AND2_X1   g787(.A1(new_n969), .A2(new_n972), .ZN(new_n974));
  OAI211_X1 g788(.A(new_n973), .B(new_n942), .C1(new_n386), .C2(new_n974), .ZN(new_n975));
  XNOR2_X1  g789(.A(KEYINPUT122), .B(KEYINPUT61), .ZN(new_n976));
  XNOR2_X1  g790(.A(new_n975), .B(new_n976), .ZN(G66));
  OAI21_X1  g791(.A(G953), .B1(new_n620), .B2(new_n430), .ZN(new_n978));
  XNOR2_X1  g792(.A(new_n978), .B(KEYINPUT123), .ZN(new_n979));
  OAI21_X1  g793(.A(new_n979), .B1(new_n873), .B2(G953), .ZN(new_n980));
  XOR2_X1   g794(.A(new_n980), .B(KEYINPUT124), .Z(new_n981));
  OAI21_X1  g795(.A(new_n933), .B1(G898), .B2(new_n189), .ZN(new_n982));
  XNOR2_X1  g796(.A(new_n981), .B(new_n982), .ZN(G69));
  NOR2_X1   g797(.A1(new_n288), .A2(new_n289), .ZN(new_n984));
  XNOR2_X1  g798(.A(new_n984), .B(new_n553), .ZN(new_n985));
  OR3_X1    g799(.A1(new_n711), .A2(KEYINPUT62), .A3(new_n824), .ZN(new_n986));
  AOI21_X1  g800(.A(new_n850), .B1(new_n646), .B2(new_n640), .ZN(new_n987));
  NOR3_X1   g801(.A1(new_n987), .A2(new_n696), .A3(new_n772), .ZN(new_n988));
  NAND2_X1  g802(.A1(new_n389), .A2(new_n988), .ZN(new_n989));
  NAND4_X1  g803(.A1(new_n803), .A2(new_n986), .A3(new_n811), .A4(new_n989), .ZN(new_n990));
  OR2_X1    g804(.A1(new_n711), .A2(new_n824), .ZN(new_n991));
  NAND2_X1  g805(.A1(new_n991), .A2(KEYINPUT62), .ZN(new_n992));
  INV_X1    g806(.A(KEYINPUT125), .ZN(new_n993));
  NAND2_X1  g807(.A1(new_n992), .A2(new_n993), .ZN(new_n994));
  NAND3_X1  g808(.A1(new_n991), .A2(KEYINPUT125), .A3(KEYINPUT62), .ZN(new_n995));
  AOI21_X1  g809(.A(new_n990), .B1(new_n994), .B2(new_n995), .ZN(new_n996));
  OAI21_X1  g810(.A(new_n985), .B1(new_n996), .B2(G953), .ZN(new_n997));
  AOI21_X1  g811(.A(new_n985), .B1(G900), .B2(G953), .ZN(new_n998));
  NAND3_X1  g812(.A1(new_n797), .A2(new_n745), .A3(new_n903), .ZN(new_n999));
  INV_X1    g813(.A(new_n786), .ZN(new_n1000));
  NOR3_X1   g814(.A1(new_n824), .A2(new_n784), .A3(new_n1000), .ZN(new_n1001));
  NAND4_X1  g815(.A1(new_n803), .A2(new_n811), .A3(new_n999), .A4(new_n1001), .ZN(new_n1002));
  OAI21_X1  g816(.A(new_n998), .B1(new_n1002), .B2(G953), .ZN(new_n1003));
  NAND2_X1  g817(.A1(new_n997), .A2(new_n1003), .ZN(new_n1004));
  INV_X1    g818(.A(G900), .ZN(new_n1005));
  OAI221_X1 g819(.A(G953), .B1(new_n505), .B2(new_n1005), .C1(new_n985), .C2(KEYINPUT126), .ZN(new_n1006));
  INV_X1    g820(.A(new_n1006), .ZN(new_n1007));
  NAND2_X1  g821(.A1(new_n1004), .A2(new_n1007), .ZN(new_n1008));
  NAND3_X1  g822(.A1(new_n997), .A2(new_n1003), .A3(new_n1006), .ZN(new_n1009));
  NAND2_X1  g823(.A1(new_n1008), .A2(new_n1009), .ZN(G72));
  NAND2_X1  g824(.A1(G472), .A2(G902), .ZN(new_n1011));
  XOR2_X1   g825(.A(new_n1011), .B(KEYINPUT63), .Z(new_n1012));
  NAND4_X1  g826(.A1(new_n856), .A2(new_n628), .A3(new_n728), .A4(new_n742), .ZN(new_n1013));
  OAI21_X1  g827(.A(new_n1012), .B1(new_n1002), .B2(new_n1013), .ZN(new_n1014));
  NAND4_X1  g828(.A1(new_n1014), .A2(new_n264), .A3(new_n194), .A4(new_n290), .ZN(new_n1015));
  NAND2_X1  g829(.A1(new_n266), .A2(new_n291), .ZN(new_n1016));
  NAND3_X1  g830(.A1(new_n916), .A2(new_n1012), .A3(new_n1016), .ZN(new_n1017));
  NAND3_X1  g831(.A1(new_n1015), .A2(new_n942), .A3(new_n1017), .ZN(new_n1018));
  NAND2_X1  g832(.A1(new_n996), .A2(new_n873), .ZN(new_n1019));
  NAND2_X1  g833(.A1(new_n1019), .A2(new_n1012), .ZN(new_n1020));
  INV_X1    g834(.A(KEYINPUT127), .ZN(new_n1021));
  INV_X1    g835(.A(new_n702), .ZN(new_n1022));
  NAND3_X1  g836(.A1(new_n1020), .A2(new_n1021), .A3(new_n1022), .ZN(new_n1023));
  INV_X1    g837(.A(new_n1012), .ZN(new_n1024));
  AOI21_X1  g838(.A(new_n1024), .B1(new_n996), .B2(new_n873), .ZN(new_n1025));
  OAI21_X1  g839(.A(KEYINPUT127), .B1(new_n1025), .B2(new_n702), .ZN(new_n1026));
  AOI21_X1  g840(.A(new_n1018), .B1(new_n1023), .B2(new_n1026), .ZN(G57));
endmodule


