//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 1 1 1 1 0 1 0 1 1 1 0 0 1 1 1 0 0 1 1 0 1 0 1 1 0 1 1 1 0 1 0 0 1 1 1 0 0 1 1 1 0 1 1 0 0 1 1 0 0 1 1 1 0 0 0 1 0 1 1 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:16:17 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n685, new_n686, new_n687,
    new_n688, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n722, new_n723, new_n724,
    new_n725, new_n726, new_n727, new_n728, new_n729, new_n730, new_n731,
    new_n732, new_n733, new_n734, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n759, new_n760, new_n762, new_n763,
    new_n764, new_n765, new_n767, new_n768, new_n769, new_n770, new_n771,
    new_n772, new_n773, new_n774, new_n776, new_n778, new_n779, new_n780,
    new_n781, new_n782, new_n783, new_n784, new_n785, new_n786, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n797, new_n798, new_n799, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n870, new_n871, new_n873, new_n874, new_n876, new_n877, new_n878,
    new_n879, new_n880, new_n881, new_n882, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n916,
    new_n917, new_n919, new_n920, new_n921, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n932, new_n933,
    new_n935, new_n936, new_n937, new_n938, new_n939, new_n940, new_n942,
    new_n943, new_n944, new_n945, new_n947, new_n948, new_n949, new_n950,
    new_n951, new_n952, new_n953, new_n955, new_n956, new_n957, new_n958,
    new_n960, new_n961, new_n962, new_n963, new_n964, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974;
  NOR2_X1   g000(.A1(G169gat), .A2(G176gat), .ZN(new_n202));
  OAI21_X1  g001(.A(KEYINPUT25), .B1(new_n202), .B2(KEYINPUT23), .ZN(new_n203));
  INV_X1    g002(.A(G183gat), .ZN(new_n204));
  INV_X1    g003(.A(G190gat), .ZN(new_n205));
  NAND2_X1  g004(.A1(new_n204), .A2(new_n205), .ZN(new_n206));
  NAND3_X1  g005(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n207));
  NAND2_X1  g006(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  AOI21_X1  g007(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n209));
  AOI21_X1  g008(.A(new_n208), .B1(KEYINPUT67), .B2(new_n209), .ZN(new_n210));
  OR2_X1    g009(.A1(new_n209), .A2(KEYINPUT67), .ZN(new_n211));
  AOI21_X1  g010(.A(new_n203), .B1(new_n210), .B2(new_n211), .ZN(new_n212));
  INV_X1    g011(.A(G169gat), .ZN(new_n213));
  INV_X1    g012(.A(G176gat), .ZN(new_n214));
  NOR2_X1   g013(.A1(new_n213), .A2(new_n214), .ZN(new_n215));
  INV_X1    g014(.A(new_n215), .ZN(new_n216));
  NAND2_X1  g015(.A1(new_n202), .A2(KEYINPUT65), .ZN(new_n217));
  INV_X1    g016(.A(KEYINPUT65), .ZN(new_n218));
  OAI21_X1  g017(.A(new_n218), .B1(G169gat), .B2(G176gat), .ZN(new_n219));
  NAND2_X1  g018(.A1(new_n217), .A2(new_n219), .ZN(new_n220));
  INV_X1    g019(.A(KEYINPUT23), .ZN(new_n221));
  OAI21_X1  g020(.A(new_n216), .B1(new_n220), .B2(new_n221), .ZN(new_n222));
  NAND2_X1  g021(.A1(new_n222), .A2(KEYINPUT66), .ZN(new_n223));
  INV_X1    g022(.A(KEYINPUT66), .ZN(new_n224));
  OAI211_X1 g023(.A(new_n224), .B(new_n216), .C1(new_n220), .C2(new_n221), .ZN(new_n225));
  NAND3_X1  g024(.A1(new_n212), .A2(new_n223), .A3(new_n225), .ZN(new_n226));
  INV_X1    g025(.A(KEYINPUT25), .ZN(new_n227));
  OR2_X1    g026(.A1(new_n206), .A2(KEYINPUT64), .ZN(new_n228));
  AOI21_X1  g027(.A(new_n209), .B1(new_n206), .B2(KEYINPUT64), .ZN(new_n229));
  AND3_X1   g028(.A1(new_n228), .A2(new_n229), .A3(new_n207), .ZN(new_n230));
  AOI21_X1  g029(.A(new_n215), .B1(KEYINPUT23), .B2(new_n202), .ZN(new_n231));
  OAI21_X1  g030(.A(new_n231), .B1(KEYINPUT23), .B2(new_n202), .ZN(new_n232));
  OAI21_X1  g031(.A(new_n227), .B1(new_n230), .B2(new_n232), .ZN(new_n233));
  NAND2_X1  g032(.A1(new_n226), .A2(new_n233), .ZN(new_n234));
  INV_X1    g033(.A(new_n202), .ZN(new_n235));
  AOI21_X1  g034(.A(new_n215), .B1(KEYINPUT26), .B2(new_n235), .ZN(new_n236));
  INV_X1    g035(.A(KEYINPUT26), .ZN(new_n237));
  NAND3_X1  g036(.A1(new_n217), .A2(new_n237), .A3(new_n219), .ZN(new_n238));
  AOI22_X1  g037(.A1(new_n236), .A2(new_n238), .B1(G183gat), .B2(G190gat), .ZN(new_n239));
  INV_X1    g038(.A(KEYINPUT68), .ZN(new_n240));
  OR2_X1    g039(.A1(new_n239), .A2(new_n240), .ZN(new_n241));
  NAND2_X1  g040(.A1(new_n204), .A2(KEYINPUT27), .ZN(new_n242));
  INV_X1    g041(.A(KEYINPUT27), .ZN(new_n243));
  NAND2_X1  g042(.A1(new_n243), .A2(G183gat), .ZN(new_n244));
  NAND3_X1  g043(.A1(new_n242), .A2(new_n244), .A3(new_n205), .ZN(new_n245));
  NAND2_X1  g044(.A1(new_n245), .A2(KEYINPUT28), .ZN(new_n246));
  XNOR2_X1  g045(.A(KEYINPUT27), .B(G183gat), .ZN(new_n247));
  INV_X1    g046(.A(KEYINPUT28), .ZN(new_n248));
  NAND3_X1  g047(.A1(new_n247), .A2(new_n248), .A3(new_n205), .ZN(new_n249));
  NAND2_X1  g048(.A1(new_n246), .A2(new_n249), .ZN(new_n250));
  AOI21_X1  g049(.A(new_n250), .B1(new_n239), .B2(new_n240), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n241), .A2(new_n251), .ZN(new_n252));
  NAND2_X1  g051(.A1(new_n234), .A2(new_n252), .ZN(new_n253));
  XNOR2_X1  g052(.A(G127gat), .B(G134gat), .ZN(new_n254));
  INV_X1    g053(.A(G113gat), .ZN(new_n255));
  INV_X1    g054(.A(G120gat), .ZN(new_n256));
  NAND2_X1  g055(.A1(new_n255), .A2(new_n256), .ZN(new_n257));
  NAND2_X1  g056(.A1(G113gat), .A2(G120gat), .ZN(new_n258));
  NAND2_X1  g057(.A1(new_n257), .A2(new_n258), .ZN(new_n259));
  AOI21_X1  g058(.A(KEYINPUT1), .B1(new_n259), .B2(KEYINPUT69), .ZN(new_n260));
  INV_X1    g059(.A(KEYINPUT69), .ZN(new_n261));
  NAND3_X1  g060(.A1(new_n257), .A2(new_n261), .A3(new_n258), .ZN(new_n262));
  AOI21_X1  g061(.A(new_n254), .B1(new_n260), .B2(new_n262), .ZN(new_n263));
  INV_X1    g062(.A(G134gat), .ZN(new_n264));
  NAND2_X1  g063(.A1(new_n264), .A2(G127gat), .ZN(new_n265));
  INV_X1    g064(.A(G127gat), .ZN(new_n266));
  NAND2_X1  g065(.A1(new_n266), .A2(G134gat), .ZN(new_n267));
  INV_X1    g066(.A(KEYINPUT1), .ZN(new_n268));
  NAND3_X1  g067(.A1(new_n265), .A2(new_n267), .A3(new_n268), .ZN(new_n269));
  OAI21_X1  g068(.A(KEYINPUT70), .B1(new_n269), .B2(new_n259), .ZN(new_n270));
  AND2_X1   g069(.A1(G113gat), .A2(G120gat), .ZN(new_n271));
  NOR2_X1   g070(.A1(G113gat), .A2(G120gat), .ZN(new_n272));
  NOR2_X1   g071(.A1(new_n271), .A2(new_n272), .ZN(new_n273));
  INV_X1    g072(.A(KEYINPUT70), .ZN(new_n274));
  NAND4_X1  g073(.A1(new_n273), .A2(new_n254), .A3(new_n274), .A4(new_n268), .ZN(new_n275));
  NAND2_X1  g074(.A1(new_n270), .A2(new_n275), .ZN(new_n276));
  OAI21_X1  g075(.A(KEYINPUT71), .B1(new_n263), .B2(new_n276), .ZN(new_n277));
  OAI21_X1  g076(.A(KEYINPUT69), .B1(new_n271), .B2(new_n272), .ZN(new_n278));
  NAND3_X1  g077(.A1(new_n278), .A2(new_n262), .A3(new_n268), .ZN(new_n279));
  INV_X1    g078(.A(new_n254), .ZN(new_n280));
  NAND2_X1  g079(.A1(new_n279), .A2(new_n280), .ZN(new_n281));
  INV_X1    g080(.A(KEYINPUT71), .ZN(new_n282));
  NAND4_X1  g081(.A1(new_n281), .A2(new_n282), .A3(new_n270), .A4(new_n275), .ZN(new_n283));
  NAND2_X1  g082(.A1(new_n277), .A2(new_n283), .ZN(new_n284));
  NAND2_X1  g083(.A1(new_n253), .A2(new_n284), .ZN(new_n285));
  INV_X1    g084(.A(G227gat), .ZN(new_n286));
  INV_X1    g085(.A(G233gat), .ZN(new_n287));
  NOR2_X1   g086(.A1(new_n286), .A2(new_n287), .ZN(new_n288));
  INV_X1    g087(.A(new_n288), .ZN(new_n289));
  NAND4_X1  g088(.A1(new_n234), .A2(new_n252), .A3(new_n277), .A4(new_n283), .ZN(new_n290));
  NAND3_X1  g089(.A1(new_n285), .A2(new_n289), .A3(new_n290), .ZN(new_n291));
  XOR2_X1   g090(.A(new_n291), .B(KEYINPUT34), .Z(new_n292));
  XOR2_X1   g091(.A(G15gat), .B(G43gat), .Z(new_n293));
  XNOR2_X1  g092(.A(G71gat), .B(G99gat), .ZN(new_n294));
  XNOR2_X1  g093(.A(new_n293), .B(new_n294), .ZN(new_n295));
  AOI21_X1  g094(.A(new_n289), .B1(new_n285), .B2(new_n290), .ZN(new_n296));
  XNOR2_X1  g095(.A(KEYINPUT72), .B(KEYINPUT33), .ZN(new_n297));
  INV_X1    g096(.A(new_n297), .ZN(new_n298));
  OAI21_X1  g097(.A(new_n295), .B1(new_n296), .B2(new_n298), .ZN(new_n299));
  INV_X1    g098(.A(KEYINPUT32), .ZN(new_n300));
  NOR2_X1   g099(.A1(new_n296), .A2(new_n300), .ZN(new_n301));
  OR2_X1    g100(.A1(new_n299), .A2(new_n301), .ZN(new_n302));
  INV_X1    g101(.A(KEYINPUT73), .ZN(new_n303));
  NAND2_X1  g102(.A1(new_n285), .A2(new_n290), .ZN(new_n304));
  AOI221_X4 g103(.A(new_n300), .B1(new_n298), .B2(new_n295), .C1(new_n304), .C2(new_n288), .ZN(new_n305));
  INV_X1    g104(.A(new_n305), .ZN(new_n306));
  NAND3_X1  g105(.A1(new_n302), .A2(new_n303), .A3(new_n306), .ZN(new_n307));
  NOR2_X1   g106(.A1(new_n299), .A2(new_n301), .ZN(new_n308));
  OAI21_X1  g107(.A(KEYINPUT73), .B1(new_n308), .B2(new_n305), .ZN(new_n309));
  AOI21_X1  g108(.A(new_n292), .B1(new_n307), .B2(new_n309), .ZN(new_n310));
  NAND3_X1  g109(.A1(new_n302), .A2(new_n292), .A3(new_n306), .ZN(new_n311));
  INV_X1    g110(.A(new_n311), .ZN(new_n312));
  NOR2_X1   g111(.A1(new_n310), .A2(new_n312), .ZN(new_n313));
  XOR2_X1   g112(.A(G78gat), .B(G106gat), .Z(new_n314));
  XNOR2_X1  g113(.A(new_n314), .B(G50gat), .ZN(new_n315));
  XNOR2_X1  g114(.A(new_n315), .B(G22gat), .ZN(new_n316));
  INV_X1    g115(.A(new_n316), .ZN(new_n317));
  NAND2_X1  g116(.A1(G228gat), .A2(G233gat), .ZN(new_n318));
  INV_X1    g117(.A(new_n318), .ZN(new_n319));
  XOR2_X1   g118(.A(G141gat), .B(G148gat), .Z(new_n320));
  XNOR2_X1  g119(.A(G155gat), .B(G162gat), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n320), .A2(new_n321), .ZN(new_n322));
  XOR2_X1   g121(.A(KEYINPUT81), .B(G155gat), .Z(new_n323));
  NAND2_X1  g122(.A1(new_n323), .A2(G162gat), .ZN(new_n324));
  AOI21_X1  g123(.A(new_n322), .B1(KEYINPUT2), .B2(new_n324), .ZN(new_n325));
  INV_X1    g124(.A(KEYINPUT80), .ZN(new_n326));
  NAND2_X1  g125(.A1(new_n321), .A2(new_n326), .ZN(new_n327));
  INV_X1    g126(.A(G155gat), .ZN(new_n328));
  INV_X1    g127(.A(G162gat), .ZN(new_n329));
  NAND2_X1  g128(.A1(new_n328), .A2(new_n329), .ZN(new_n330));
  NAND2_X1  g129(.A1(G155gat), .A2(G162gat), .ZN(new_n331));
  NAND3_X1  g130(.A1(new_n330), .A2(KEYINPUT80), .A3(new_n331), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n331), .A2(KEYINPUT2), .ZN(new_n333));
  AOI22_X1  g132(.A1(new_n327), .A2(new_n332), .B1(new_n320), .B2(new_n333), .ZN(new_n334));
  OAI21_X1  g133(.A(KEYINPUT82), .B1(new_n325), .B2(new_n334), .ZN(new_n335));
  NAND2_X1  g134(.A1(new_n327), .A2(new_n332), .ZN(new_n336));
  NAND2_X1  g135(.A1(new_n320), .A2(new_n333), .ZN(new_n337));
  NAND2_X1  g136(.A1(new_n336), .A2(new_n337), .ZN(new_n338));
  INV_X1    g137(.A(KEYINPUT82), .ZN(new_n339));
  XNOR2_X1  g138(.A(KEYINPUT81), .B(G155gat), .ZN(new_n340));
  OAI21_X1  g139(.A(KEYINPUT2), .B1(new_n340), .B2(new_n329), .ZN(new_n341));
  NAND3_X1  g140(.A1(new_n341), .A2(new_n320), .A3(new_n321), .ZN(new_n342));
  NAND3_X1  g141(.A1(new_n338), .A2(new_n339), .A3(new_n342), .ZN(new_n343));
  NAND2_X1  g142(.A1(new_n335), .A2(new_n343), .ZN(new_n344));
  XNOR2_X1  g143(.A(G211gat), .B(G218gat), .ZN(new_n345));
  INV_X1    g144(.A(new_n345), .ZN(new_n346));
  XNOR2_X1  g145(.A(G197gat), .B(G204gat), .ZN(new_n347));
  INV_X1    g146(.A(new_n347), .ZN(new_n348));
  OR2_X1    g147(.A1(KEYINPUT75), .A2(G218gat), .ZN(new_n349));
  NAND2_X1  g148(.A1(KEYINPUT75), .A2(G218gat), .ZN(new_n350));
  NAND2_X1  g149(.A1(new_n349), .A2(new_n350), .ZN(new_n351));
  NAND2_X1  g150(.A1(new_n351), .A2(G211gat), .ZN(new_n352));
  XNOR2_X1  g151(.A(KEYINPUT74), .B(KEYINPUT22), .ZN(new_n353));
  INV_X1    g152(.A(new_n353), .ZN(new_n354));
  AOI21_X1  g153(.A(new_n348), .B1(new_n352), .B2(new_n354), .ZN(new_n355));
  INV_X1    g154(.A(KEYINPUT76), .ZN(new_n356));
  OAI21_X1  g155(.A(new_n346), .B1(new_n355), .B2(new_n356), .ZN(new_n357));
  INV_X1    g156(.A(G211gat), .ZN(new_n358));
  AOI21_X1  g157(.A(new_n358), .B1(new_n349), .B2(new_n350), .ZN(new_n359));
  OAI21_X1  g158(.A(new_n347), .B1(new_n359), .B2(new_n353), .ZN(new_n360));
  NOR2_X1   g159(.A1(new_n360), .A2(KEYINPUT76), .ZN(new_n361));
  OAI21_X1  g160(.A(KEYINPUT77), .B1(new_n357), .B2(new_n361), .ZN(new_n362));
  AOI21_X1  g161(.A(new_n345), .B1(new_n360), .B2(KEYINPUT76), .ZN(new_n363));
  INV_X1    g162(.A(KEYINPUT77), .ZN(new_n364));
  OAI211_X1 g163(.A(new_n363), .B(new_n364), .C1(KEYINPUT76), .C2(new_n360), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n355), .A2(new_n345), .ZN(new_n366));
  NAND3_X1  g165(.A1(new_n362), .A2(new_n365), .A3(new_n366), .ZN(new_n367));
  INV_X1    g166(.A(KEYINPUT29), .ZN(new_n368));
  NAND2_X1  g167(.A1(new_n367), .A2(new_n368), .ZN(new_n369));
  INV_X1    g168(.A(KEYINPUT3), .ZN(new_n370));
  AOI21_X1  g169(.A(new_n344), .B1(new_n369), .B2(new_n370), .ZN(new_n371));
  NAND3_X1  g170(.A1(new_n338), .A2(new_n370), .A3(new_n342), .ZN(new_n372));
  XOR2_X1   g171(.A(KEYINPUT78), .B(KEYINPUT29), .Z(new_n373));
  AND2_X1   g172(.A1(new_n372), .A2(new_n373), .ZN(new_n374));
  NOR2_X1   g173(.A1(new_n367), .A2(new_n374), .ZN(new_n375));
  OAI21_X1  g174(.A(new_n319), .B1(new_n371), .B2(new_n375), .ZN(new_n376));
  NAND2_X1  g175(.A1(new_n338), .A2(new_n342), .ZN(new_n377));
  INV_X1    g176(.A(new_n373), .ZN(new_n378));
  NAND2_X1  g177(.A1(new_n360), .A2(new_n346), .ZN(new_n379));
  AOI21_X1  g178(.A(new_n378), .B1(new_n366), .B2(new_n379), .ZN(new_n380));
  AND2_X1   g179(.A1(new_n380), .A2(KEYINPUT88), .ZN(new_n381));
  OAI21_X1  g180(.A(new_n370), .B1(new_n380), .B2(KEYINPUT88), .ZN(new_n382));
  OAI21_X1  g181(.A(new_n377), .B1(new_n381), .B2(new_n382), .ZN(new_n383));
  OAI211_X1 g182(.A(new_n383), .B(new_n318), .C1(new_n367), .C2(new_n374), .ZN(new_n384));
  XNOR2_X1  g183(.A(KEYINPUT87), .B(KEYINPUT31), .ZN(new_n385));
  INV_X1    g184(.A(new_n385), .ZN(new_n386));
  AND3_X1   g185(.A1(new_n376), .A2(new_n384), .A3(new_n386), .ZN(new_n387));
  AOI21_X1  g186(.A(new_n386), .B1(new_n376), .B2(new_n384), .ZN(new_n388));
  OAI21_X1  g187(.A(new_n317), .B1(new_n387), .B2(new_n388), .ZN(new_n389));
  NAND2_X1  g188(.A1(new_n376), .A2(new_n384), .ZN(new_n390));
  NAND2_X1  g189(.A1(new_n390), .A2(new_n385), .ZN(new_n391));
  NAND3_X1  g190(.A1(new_n376), .A2(new_n384), .A3(new_n386), .ZN(new_n392));
  NAND3_X1  g191(.A1(new_n391), .A2(new_n316), .A3(new_n392), .ZN(new_n393));
  AND2_X1   g192(.A1(new_n389), .A2(new_n393), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n313), .A2(new_n394), .ZN(new_n395));
  INV_X1    g194(.A(new_n367), .ZN(new_n396));
  NAND2_X1  g195(.A1(G226gat), .A2(G233gat), .ZN(new_n397));
  INV_X1    g196(.A(new_n397), .ZN(new_n398));
  AOI21_X1  g197(.A(new_n398), .B1(new_n253), .B2(new_n373), .ZN(new_n399));
  AOI22_X1  g198(.A1(new_n233), .A2(new_n226), .B1(new_n241), .B2(new_n251), .ZN(new_n400));
  NOR2_X1   g199(.A1(new_n400), .A2(new_n397), .ZN(new_n401));
  OAI21_X1  g200(.A(new_n396), .B1(new_n399), .B2(new_n401), .ZN(new_n402));
  NAND2_X1  g201(.A1(new_n253), .A2(new_n398), .ZN(new_n403));
  NOR2_X1   g202(.A1(new_n400), .A2(KEYINPUT29), .ZN(new_n404));
  OAI211_X1 g203(.A(new_n403), .B(new_n367), .C1(new_n404), .C2(new_n398), .ZN(new_n405));
  XNOR2_X1  g204(.A(G8gat), .B(G36gat), .ZN(new_n406));
  XNOR2_X1  g205(.A(G64gat), .B(G92gat), .ZN(new_n407));
  XOR2_X1   g206(.A(new_n406), .B(new_n407), .Z(new_n408));
  NAND3_X1  g207(.A1(new_n402), .A2(new_n405), .A3(new_n408), .ZN(new_n409));
  INV_X1    g208(.A(KEYINPUT30), .ZN(new_n410));
  NAND2_X1  g209(.A1(new_n409), .A2(new_n410), .ZN(new_n411));
  NAND4_X1  g210(.A1(new_n402), .A2(new_n405), .A3(KEYINPUT30), .A4(new_n408), .ZN(new_n412));
  INV_X1    g211(.A(KEYINPUT79), .ZN(new_n413));
  NAND2_X1  g212(.A1(new_n402), .A2(new_n405), .ZN(new_n414));
  INV_X1    g213(.A(new_n408), .ZN(new_n415));
  AOI21_X1  g214(.A(new_n413), .B1(new_n414), .B2(new_n415), .ZN(new_n416));
  AOI211_X1 g215(.A(KEYINPUT79), .B(new_n408), .C1(new_n402), .C2(new_n405), .ZN(new_n417));
  OAI211_X1 g216(.A(new_n411), .B(new_n412), .C1(new_n416), .C2(new_n417), .ZN(new_n418));
  INV_X1    g217(.A(new_n418), .ZN(new_n419));
  NAND2_X1  g218(.A1(G225gat), .A2(G233gat), .ZN(new_n420));
  INV_X1    g219(.A(new_n420), .ZN(new_n421));
  NAND3_X1  g220(.A1(new_n335), .A2(KEYINPUT3), .A3(new_n343), .ZN(new_n422));
  NAND3_X1  g221(.A1(new_n281), .A2(new_n270), .A3(new_n275), .ZN(new_n423));
  AND2_X1   g222(.A1(new_n372), .A2(new_n423), .ZN(new_n424));
  AOI21_X1  g223(.A(new_n421), .B1(new_n422), .B2(new_n424), .ZN(new_n425));
  XOR2_X1   g224(.A(KEYINPUT84), .B(KEYINPUT5), .Z(new_n426));
  INV_X1    g225(.A(new_n322), .ZN(new_n427));
  AOI21_X1  g226(.A(new_n334), .B1(new_n341), .B2(new_n427), .ZN(new_n428));
  INV_X1    g227(.A(KEYINPUT4), .ZN(new_n429));
  NAND4_X1  g228(.A1(new_n277), .A2(new_n428), .A3(new_n429), .A4(new_n283), .ZN(new_n430));
  OAI21_X1  g229(.A(KEYINPUT4), .B1(new_n423), .B2(new_n377), .ZN(new_n431));
  AND3_X1   g230(.A1(new_n430), .A2(KEYINPUT85), .A3(new_n431), .ZN(new_n432));
  AOI21_X1  g231(.A(KEYINPUT85), .B1(new_n430), .B2(new_n431), .ZN(new_n433));
  OAI211_X1 g232(.A(new_n425), .B(new_n426), .C1(new_n432), .C2(new_n433), .ZN(new_n434));
  NAND2_X1  g233(.A1(new_n422), .A2(new_n424), .ZN(new_n435));
  NAND2_X1  g234(.A1(new_n435), .A2(new_n420), .ZN(new_n436));
  NOR3_X1   g235(.A1(new_n423), .A2(new_n377), .A3(KEYINPUT4), .ZN(new_n437));
  NAND3_X1  g236(.A1(new_n277), .A2(new_n428), .A3(new_n283), .ZN(new_n438));
  NAND2_X1  g237(.A1(new_n438), .A2(KEYINPUT4), .ZN(new_n439));
  INV_X1    g238(.A(KEYINPUT83), .ZN(new_n440));
  AOI21_X1  g239(.A(new_n437), .B1(new_n439), .B2(new_n440), .ZN(new_n441));
  NAND3_X1  g240(.A1(new_n438), .A2(KEYINPUT83), .A3(KEYINPUT4), .ZN(new_n442));
  AOI21_X1  g241(.A(new_n436), .B1(new_n441), .B2(new_n442), .ZN(new_n443));
  NAND3_X1  g242(.A1(new_n335), .A2(new_n343), .A3(new_n423), .ZN(new_n444));
  OAI21_X1  g243(.A(new_n444), .B1(new_n377), .B2(new_n423), .ZN(new_n445));
  AOI21_X1  g244(.A(new_n426), .B1(new_n445), .B2(new_n421), .ZN(new_n446));
  INV_X1    g245(.A(new_n446), .ZN(new_n447));
  OAI21_X1  g246(.A(new_n434), .B1(new_n443), .B2(new_n447), .ZN(new_n448));
  XNOR2_X1  g247(.A(G1gat), .B(G29gat), .ZN(new_n449));
  XNOR2_X1  g248(.A(new_n449), .B(KEYINPUT0), .ZN(new_n450));
  XNOR2_X1  g249(.A(G57gat), .B(G85gat), .ZN(new_n451));
  XOR2_X1   g250(.A(new_n450), .B(new_n451), .Z(new_n452));
  INV_X1    g251(.A(new_n452), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n448), .A2(new_n453), .ZN(new_n454));
  AND3_X1   g253(.A1(new_n438), .A2(KEYINPUT83), .A3(KEYINPUT4), .ZN(new_n455));
  AOI21_X1  g254(.A(KEYINPUT83), .B1(new_n438), .B2(KEYINPUT4), .ZN(new_n456));
  NOR3_X1   g255(.A1(new_n455), .A2(new_n456), .A3(new_n437), .ZN(new_n457));
  OAI21_X1  g256(.A(new_n446), .B1(new_n457), .B2(new_n436), .ZN(new_n458));
  NAND3_X1  g257(.A1(new_n458), .A2(new_n452), .A3(new_n434), .ZN(new_n459));
  XOR2_X1   g258(.A(KEYINPUT86), .B(KEYINPUT6), .Z(new_n460));
  NAND3_X1  g259(.A1(new_n454), .A2(new_n459), .A3(new_n460), .ZN(new_n461));
  INV_X1    g260(.A(new_n460), .ZN(new_n462));
  NAND3_X1  g261(.A1(new_n448), .A2(new_n453), .A3(new_n462), .ZN(new_n463));
  NAND2_X1  g262(.A1(new_n461), .A2(new_n463), .ZN(new_n464));
  NAND2_X1  g263(.A1(new_n419), .A2(new_n464), .ZN(new_n465));
  OAI21_X1  g264(.A(KEYINPUT35), .B1(new_n395), .B2(new_n465), .ZN(new_n466));
  NAND2_X1  g265(.A1(new_n389), .A2(new_n393), .ZN(new_n467));
  INV_X1    g266(.A(new_n292), .ZN(new_n468));
  OAI21_X1  g267(.A(new_n468), .B1(new_n308), .B2(new_n305), .ZN(new_n469));
  NAND2_X1  g268(.A1(new_n469), .A2(new_n311), .ZN(new_n470));
  NOR2_X1   g269(.A1(new_n467), .A2(new_n470), .ZN(new_n471));
  AOI21_X1  g270(.A(new_n452), .B1(new_n458), .B2(new_n434), .ZN(new_n472));
  INV_X1    g271(.A(KEYINPUT89), .ZN(new_n473));
  NAND3_X1  g272(.A1(new_n472), .A2(new_n473), .A3(new_n462), .ZN(new_n474));
  NAND2_X1  g273(.A1(new_n463), .A2(KEYINPUT89), .ZN(new_n475));
  NAND2_X1  g274(.A1(new_n474), .A2(new_n475), .ZN(new_n476));
  NAND2_X1  g275(.A1(new_n476), .A2(new_n461), .ZN(new_n477));
  NOR2_X1   g276(.A1(new_n418), .A2(KEYINPUT35), .ZN(new_n478));
  NAND3_X1  g277(.A1(new_n471), .A2(new_n477), .A3(new_n478), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n466), .A2(new_n479), .ZN(new_n480));
  AND2_X1   g279(.A1(new_n307), .A2(new_n309), .ZN(new_n481));
  OAI211_X1 g280(.A(KEYINPUT36), .B(new_n311), .C1(new_n481), .C2(new_n292), .ZN(new_n482));
  AOI21_X1  g281(.A(KEYINPUT36), .B1(new_n469), .B2(new_n311), .ZN(new_n483));
  INV_X1    g282(.A(new_n483), .ZN(new_n484));
  AOI22_X1  g283(.A1(new_n482), .A2(new_n484), .B1(new_n465), .B2(new_n467), .ZN(new_n485));
  OAI21_X1  g284(.A(new_n435), .B1(new_n432), .B2(new_n433), .ZN(new_n486));
  NAND2_X1  g285(.A1(new_n486), .A2(new_n421), .ZN(new_n487));
  OR2_X1    g286(.A1(new_n445), .A2(new_n421), .ZN(new_n488));
  NAND3_X1  g287(.A1(new_n487), .A2(KEYINPUT39), .A3(new_n488), .ZN(new_n489));
  INV_X1    g288(.A(KEYINPUT39), .ZN(new_n490));
  NAND3_X1  g289(.A1(new_n486), .A2(new_n490), .A3(new_n421), .ZN(new_n491));
  NAND3_X1  g290(.A1(new_n489), .A2(new_n452), .A3(new_n491), .ZN(new_n492));
  INV_X1    g291(.A(KEYINPUT40), .ZN(new_n493));
  NAND2_X1  g292(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  NAND4_X1  g293(.A1(new_n489), .A2(KEYINPUT40), .A3(new_n452), .A4(new_n491), .ZN(new_n495));
  NAND4_X1  g294(.A1(new_n418), .A2(new_n494), .A3(new_n454), .A4(new_n495), .ZN(new_n496));
  NAND2_X1  g295(.A1(new_n394), .A2(new_n496), .ZN(new_n497));
  AOI21_X1  g296(.A(new_n398), .B1(new_n253), .B2(new_n368), .ZN(new_n498));
  NOR3_X1   g297(.A1(new_n498), .A2(new_n401), .A3(new_n396), .ZN(new_n499));
  OAI21_X1  g298(.A(new_n397), .B1(new_n400), .B2(new_n378), .ZN(new_n500));
  AOI21_X1  g299(.A(new_n367), .B1(new_n500), .B2(new_n403), .ZN(new_n501));
  OAI21_X1  g300(.A(new_n415), .B1(new_n499), .B2(new_n501), .ZN(new_n502));
  NAND2_X1  g301(.A1(new_n415), .A2(KEYINPUT37), .ZN(new_n503));
  NAND2_X1  g302(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  NAND2_X1  g303(.A1(new_n414), .A2(KEYINPUT37), .ZN(new_n505));
  NAND2_X1  g304(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  NAND2_X1  g305(.A1(new_n506), .A2(KEYINPUT38), .ZN(new_n507));
  INV_X1    g306(.A(new_n507), .ZN(new_n508));
  INV_X1    g307(.A(new_n409), .ZN(new_n509));
  INV_X1    g308(.A(KEYINPUT37), .ZN(new_n510));
  NAND2_X1  g309(.A1(new_n500), .A2(new_n403), .ZN(new_n511));
  AOI21_X1  g310(.A(new_n510), .B1(new_n511), .B2(new_n367), .ZN(new_n512));
  OAI211_X1 g311(.A(new_n403), .B(new_n396), .C1(new_n404), .C2(new_n398), .ZN(new_n513));
  AOI21_X1  g312(.A(KEYINPUT38), .B1(new_n512), .B2(new_n513), .ZN(new_n514));
  AOI21_X1  g313(.A(new_n509), .B1(new_n504), .B2(new_n514), .ZN(new_n515));
  AOI21_X1  g314(.A(new_n473), .B1(new_n472), .B2(new_n462), .ZN(new_n516));
  AND4_X1   g315(.A1(new_n473), .A2(new_n448), .A3(new_n453), .A4(new_n462), .ZN(new_n517));
  OAI211_X1 g316(.A(new_n461), .B(new_n515), .C1(new_n516), .C2(new_n517), .ZN(new_n518));
  INV_X1    g317(.A(KEYINPUT90), .ZN(new_n519));
  AOI21_X1  g318(.A(new_n508), .B1(new_n518), .B2(new_n519), .ZN(new_n520));
  NAND4_X1  g319(.A1(new_n476), .A2(KEYINPUT90), .A3(new_n461), .A4(new_n515), .ZN(new_n521));
  AOI21_X1  g320(.A(new_n497), .B1(new_n520), .B2(new_n521), .ZN(new_n522));
  OAI21_X1  g321(.A(new_n485), .B1(new_n522), .B2(KEYINPUT91), .ZN(new_n523));
  NAND2_X1  g322(.A1(new_n518), .A2(new_n519), .ZN(new_n524));
  NAND3_X1  g323(.A1(new_n524), .A2(new_n521), .A3(new_n507), .ZN(new_n525));
  INV_X1    g324(.A(new_n497), .ZN(new_n526));
  AND3_X1   g325(.A1(new_n525), .A2(KEYINPUT91), .A3(new_n526), .ZN(new_n527));
  OAI21_X1  g326(.A(new_n480), .B1(new_n523), .B2(new_n527), .ZN(new_n528));
  NOR2_X1   g327(.A1(G29gat), .A2(G36gat), .ZN(new_n529));
  XOR2_X1   g328(.A(new_n529), .B(KEYINPUT14), .Z(new_n530));
  NAND2_X1  g329(.A1(G29gat), .A2(G36gat), .ZN(new_n531));
  XNOR2_X1  g330(.A(new_n531), .B(KEYINPUT92), .ZN(new_n532));
  NAND2_X1  g331(.A1(new_n530), .A2(new_n532), .ZN(new_n533));
  NAND2_X1  g332(.A1(G43gat), .A2(G50gat), .ZN(new_n534));
  INV_X1    g333(.A(new_n534), .ZN(new_n535));
  NOR2_X1   g334(.A1(G43gat), .A2(G50gat), .ZN(new_n536));
  OAI21_X1  g335(.A(KEYINPUT15), .B1(new_n535), .B2(new_n536), .ZN(new_n537));
  OR2_X1    g336(.A1(new_n533), .A2(new_n537), .ZN(new_n538));
  AND2_X1   g337(.A1(KEYINPUT93), .A2(KEYINPUT15), .ZN(new_n539));
  OAI21_X1  g338(.A(new_n534), .B1(KEYINPUT93), .B2(KEYINPUT15), .ZN(new_n540));
  INV_X1    g339(.A(G43gat), .ZN(new_n541));
  XNOR2_X1  g340(.A(KEYINPUT94), .B(G50gat), .ZN(new_n542));
  AOI211_X1 g341(.A(new_n539), .B(new_n540), .C1(new_n541), .C2(new_n542), .ZN(new_n543));
  OAI21_X1  g342(.A(new_n537), .B1(new_n533), .B2(new_n543), .ZN(new_n544));
  NAND2_X1  g343(.A1(new_n538), .A2(new_n544), .ZN(new_n545));
  OR2_X1    g344(.A1(new_n545), .A2(KEYINPUT17), .ZN(new_n546));
  XNOR2_X1  g345(.A(G15gat), .B(G22gat), .ZN(new_n547));
  INV_X1    g346(.A(G1gat), .ZN(new_n548));
  NAND3_X1  g347(.A1(new_n547), .A2(KEYINPUT16), .A3(new_n548), .ZN(new_n549));
  OAI221_X1 g348(.A(new_n549), .B1(KEYINPUT95), .B2(G8gat), .C1(new_n548), .C2(new_n547), .ZN(new_n550));
  NAND2_X1  g349(.A1(KEYINPUT95), .A2(G8gat), .ZN(new_n551));
  XOR2_X1   g350(.A(new_n550), .B(new_n551), .Z(new_n552));
  NAND2_X1  g351(.A1(new_n545), .A2(KEYINPUT17), .ZN(new_n553));
  NAND3_X1  g352(.A1(new_n546), .A2(new_n552), .A3(new_n553), .ZN(new_n554));
  NAND2_X1  g353(.A1(G229gat), .A2(G233gat), .ZN(new_n555));
  AND2_X1   g354(.A1(new_n538), .A2(new_n544), .ZN(new_n556));
  XNOR2_X1  g355(.A(new_n550), .B(new_n551), .ZN(new_n557));
  NAND2_X1  g356(.A1(new_n556), .A2(new_n557), .ZN(new_n558));
  NAND3_X1  g357(.A1(new_n554), .A2(new_n555), .A3(new_n558), .ZN(new_n559));
  NOR2_X1   g358(.A1(KEYINPUT96), .A2(KEYINPUT18), .ZN(new_n560));
  OR2_X1    g359(.A1(new_n559), .A2(new_n560), .ZN(new_n561));
  NAND2_X1  g360(.A1(new_n559), .A2(new_n560), .ZN(new_n562));
  NAND2_X1  g361(.A1(new_n552), .A2(new_n545), .ZN(new_n563));
  NAND3_X1  g362(.A1(new_n563), .A2(KEYINPUT98), .A3(new_n558), .ZN(new_n564));
  XNOR2_X1  g363(.A(KEYINPUT97), .B(KEYINPUT13), .ZN(new_n565));
  XNOR2_X1  g364(.A(new_n565), .B(new_n555), .ZN(new_n566));
  OR3_X1    g365(.A1(new_n556), .A2(new_n557), .A3(KEYINPUT98), .ZN(new_n567));
  NAND3_X1  g366(.A1(new_n564), .A2(new_n566), .A3(new_n567), .ZN(new_n568));
  AND3_X1   g367(.A1(new_n561), .A2(new_n562), .A3(new_n568), .ZN(new_n569));
  XNOR2_X1  g368(.A(G113gat), .B(G141gat), .ZN(new_n570));
  XNOR2_X1  g369(.A(new_n570), .B(G197gat), .ZN(new_n571));
  XOR2_X1   g370(.A(KEYINPUT11), .B(G169gat), .Z(new_n572));
  XNOR2_X1  g371(.A(new_n571), .B(new_n572), .ZN(new_n573));
  XNOR2_X1  g372(.A(new_n573), .B(KEYINPUT12), .ZN(new_n574));
  OR2_X1    g373(.A1(new_n569), .A2(new_n574), .ZN(new_n575));
  NAND4_X1  g374(.A1(new_n561), .A2(new_n574), .A3(new_n562), .A4(new_n568), .ZN(new_n576));
  NAND2_X1  g375(.A1(new_n575), .A2(new_n576), .ZN(new_n577));
  INV_X1    g376(.A(KEYINPUT106), .ZN(new_n578));
  AOI21_X1  g377(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n579));
  INV_X1    g378(.A(KEYINPUT99), .ZN(new_n580));
  XNOR2_X1  g379(.A(new_n579), .B(new_n580), .ZN(new_n581));
  XNOR2_X1  g380(.A(G71gat), .B(G78gat), .ZN(new_n582));
  XOR2_X1   g381(.A(G57gat), .B(G64gat), .Z(new_n583));
  NAND3_X1  g382(.A1(new_n581), .A2(new_n582), .A3(new_n583), .ZN(new_n584));
  OR2_X1    g383(.A1(new_n584), .A2(KEYINPUT100), .ZN(new_n585));
  AND2_X1   g384(.A1(new_n583), .A2(KEYINPUT9), .ZN(new_n586));
  OAI211_X1 g385(.A(new_n584), .B(KEYINPUT100), .C1(new_n582), .C2(new_n586), .ZN(new_n587));
  NAND2_X1  g386(.A1(new_n585), .A2(new_n587), .ZN(new_n588));
  NOR2_X1   g387(.A1(new_n588), .A2(KEYINPUT101), .ZN(new_n589));
  INV_X1    g388(.A(KEYINPUT101), .ZN(new_n590));
  AOI21_X1  g389(.A(new_n590), .B1(new_n585), .B2(new_n587), .ZN(new_n591));
  NOR2_X1   g390(.A1(new_n589), .A2(new_n591), .ZN(new_n592));
  AOI21_X1  g391(.A(new_n557), .B1(new_n592), .B2(KEYINPUT21), .ZN(new_n593));
  OAI211_X1 g392(.A(G231gat), .B(G233gat), .C1(new_n592), .C2(KEYINPUT21), .ZN(new_n594));
  INV_X1    g393(.A(KEYINPUT21), .ZN(new_n595));
  NAND2_X1  g394(.A1(G231gat), .A2(G233gat), .ZN(new_n596));
  OAI211_X1 g395(.A(new_n595), .B(new_n596), .C1(new_n589), .C2(new_n591), .ZN(new_n597));
  NAND3_X1  g396(.A1(new_n594), .A2(new_n266), .A3(new_n597), .ZN(new_n598));
  INV_X1    g397(.A(new_n598), .ZN(new_n599));
  AOI21_X1  g398(.A(new_n266), .B1(new_n594), .B2(new_n597), .ZN(new_n600));
  OAI21_X1  g399(.A(new_n593), .B1(new_n599), .B2(new_n600), .ZN(new_n601));
  INV_X1    g400(.A(new_n600), .ZN(new_n602));
  INV_X1    g401(.A(new_n593), .ZN(new_n603));
  NAND3_X1  g402(.A1(new_n602), .A2(new_n603), .A3(new_n598), .ZN(new_n604));
  NAND2_X1  g403(.A1(new_n601), .A2(new_n604), .ZN(new_n605));
  XNOR2_X1  g404(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n606));
  XNOR2_X1  g405(.A(new_n606), .B(new_n328), .ZN(new_n607));
  XNOR2_X1  g406(.A(G183gat), .B(G211gat), .ZN(new_n608));
  XOR2_X1   g407(.A(new_n607), .B(new_n608), .Z(new_n609));
  INV_X1    g408(.A(new_n609), .ZN(new_n610));
  NAND2_X1  g409(.A1(new_n605), .A2(new_n610), .ZN(new_n611));
  NAND3_X1  g410(.A1(new_n601), .A2(new_n604), .A3(new_n609), .ZN(new_n612));
  NAND2_X1  g411(.A1(new_n611), .A2(new_n612), .ZN(new_n613));
  NAND2_X1  g412(.A1(G85gat), .A2(G92gat), .ZN(new_n614));
  XNOR2_X1  g413(.A(new_n614), .B(KEYINPUT7), .ZN(new_n615));
  NAND2_X1  g414(.A1(G99gat), .A2(G106gat), .ZN(new_n616));
  INV_X1    g415(.A(G85gat), .ZN(new_n617));
  INV_X1    g416(.A(G92gat), .ZN(new_n618));
  AOI22_X1  g417(.A1(KEYINPUT8), .A2(new_n616), .B1(new_n617), .B2(new_n618), .ZN(new_n619));
  NAND2_X1  g418(.A1(new_n615), .A2(new_n619), .ZN(new_n620));
  INV_X1    g419(.A(KEYINPUT102), .ZN(new_n621));
  XNOR2_X1  g420(.A(new_n620), .B(new_n621), .ZN(new_n622));
  XOR2_X1   g421(.A(G99gat), .B(G106gat), .Z(new_n623));
  NAND2_X1  g422(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  XNOR2_X1  g423(.A(new_n620), .B(KEYINPUT102), .ZN(new_n625));
  INV_X1    g424(.A(new_n623), .ZN(new_n626));
  NAND2_X1  g425(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  NAND2_X1  g426(.A1(new_n624), .A2(new_n627), .ZN(new_n628));
  NAND3_X1  g427(.A1(new_n546), .A2(new_n553), .A3(new_n628), .ZN(new_n629));
  INV_X1    g428(.A(new_n628), .ZN(new_n630));
  NAND2_X1  g429(.A1(new_n630), .A2(new_n556), .ZN(new_n631));
  NAND3_X1  g430(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n632));
  NAND3_X1  g431(.A1(new_n629), .A2(new_n631), .A3(new_n632), .ZN(new_n633));
  XOR2_X1   g432(.A(G190gat), .B(G218gat), .Z(new_n634));
  INV_X1    g433(.A(new_n634), .ZN(new_n635));
  XNOR2_X1  g434(.A(new_n633), .B(new_n635), .ZN(new_n636));
  XNOR2_X1  g435(.A(G134gat), .B(G162gat), .ZN(new_n637));
  AOI21_X1  g436(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n638));
  XNOR2_X1  g437(.A(new_n637), .B(new_n638), .ZN(new_n639));
  XNOR2_X1  g438(.A(new_n636), .B(new_n639), .ZN(new_n640));
  NAND2_X1  g439(.A1(new_n613), .A2(new_n640), .ZN(new_n641));
  OAI21_X1  g440(.A(new_n628), .B1(new_n589), .B2(new_n591), .ZN(new_n642));
  INV_X1    g441(.A(KEYINPUT10), .ZN(new_n643));
  NAND3_X1  g442(.A1(new_n588), .A2(new_n624), .A3(new_n627), .ZN(new_n644));
  INV_X1    g443(.A(KEYINPUT103), .ZN(new_n645));
  NAND2_X1  g444(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  NAND4_X1  g445(.A1(new_n588), .A2(new_n624), .A3(new_n627), .A4(KEYINPUT103), .ZN(new_n647));
  NAND4_X1  g446(.A1(new_n642), .A2(new_n643), .A3(new_n646), .A4(new_n647), .ZN(new_n648));
  NAND3_X1  g447(.A1(new_n592), .A2(KEYINPUT10), .A3(new_n630), .ZN(new_n649));
  AND3_X1   g448(.A1(new_n648), .A2(KEYINPUT104), .A3(new_n649), .ZN(new_n650));
  AOI21_X1  g449(.A(KEYINPUT104), .B1(new_n648), .B2(new_n649), .ZN(new_n651));
  NAND2_X1  g450(.A1(G230gat), .A2(G233gat), .ZN(new_n652));
  INV_X1    g451(.A(new_n652), .ZN(new_n653));
  NOR3_X1   g452(.A1(new_n650), .A2(new_n651), .A3(new_n653), .ZN(new_n654));
  NAND3_X1  g453(.A1(new_n642), .A2(new_n647), .A3(new_n646), .ZN(new_n655));
  NAND2_X1  g454(.A1(new_n655), .A2(new_n653), .ZN(new_n656));
  XNOR2_X1  g455(.A(G120gat), .B(G148gat), .ZN(new_n657));
  XNOR2_X1  g456(.A(G176gat), .B(G204gat), .ZN(new_n658));
  XOR2_X1   g457(.A(new_n657), .B(new_n658), .Z(new_n659));
  NAND2_X1  g458(.A1(new_n656), .A2(new_n659), .ZN(new_n660));
  AOI21_X1  g459(.A(new_n653), .B1(new_n648), .B2(new_n649), .ZN(new_n661));
  AOI21_X1  g460(.A(new_n661), .B1(new_n655), .B2(new_n653), .ZN(new_n662));
  XOR2_X1   g461(.A(new_n659), .B(KEYINPUT105), .Z(new_n663));
  INV_X1    g462(.A(new_n663), .ZN(new_n664));
  OAI22_X1  g463(.A1(new_n654), .A2(new_n660), .B1(new_n662), .B2(new_n664), .ZN(new_n665));
  OAI21_X1  g464(.A(new_n578), .B1(new_n641), .B2(new_n665), .ZN(new_n666));
  INV_X1    g465(.A(new_n665), .ZN(new_n667));
  NAND4_X1  g466(.A1(new_n613), .A2(KEYINPUT106), .A3(new_n640), .A4(new_n667), .ZN(new_n668));
  NAND4_X1  g467(.A1(new_n528), .A2(new_n577), .A3(new_n666), .A4(new_n668), .ZN(new_n669));
  NOR2_X1   g468(.A1(new_n669), .A2(new_n464), .ZN(new_n670));
  XNOR2_X1  g469(.A(new_n670), .B(new_n548), .ZN(G1324gat));
  NOR2_X1   g470(.A1(new_n669), .A2(new_n419), .ZN(new_n672));
  XOR2_X1   g471(.A(KEYINPUT16), .B(G8gat), .Z(new_n673));
  NAND2_X1  g472(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  INV_X1    g473(.A(G8gat), .ZN(new_n675));
  OAI21_X1  g474(.A(new_n674), .B1(new_n675), .B2(new_n672), .ZN(new_n676));
  MUX2_X1   g475(.A(new_n674), .B(new_n676), .S(KEYINPUT42), .Z(G1325gat));
  INV_X1    g476(.A(KEYINPUT36), .ZN(new_n678));
  NOR3_X1   g477(.A1(new_n310), .A2(new_n678), .A3(new_n312), .ZN(new_n679));
  NOR2_X1   g478(.A1(new_n679), .A2(new_n483), .ZN(new_n680));
  INV_X1    g479(.A(new_n680), .ZN(new_n681));
  OAI21_X1  g480(.A(G15gat), .B1(new_n669), .B2(new_n681), .ZN(new_n682));
  OR2_X1    g481(.A1(new_n470), .A2(G15gat), .ZN(new_n683));
  OAI21_X1  g482(.A(new_n682), .B1(new_n669), .B2(new_n683), .ZN(G1326gat));
  OR3_X1    g483(.A1(new_n669), .A2(KEYINPUT107), .A3(new_n394), .ZN(new_n685));
  OAI21_X1  g484(.A(KEYINPUT107), .B1(new_n669), .B2(new_n394), .ZN(new_n686));
  NAND2_X1  g485(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  XNOR2_X1  g486(.A(KEYINPUT43), .B(G22gat), .ZN(new_n688));
  XNOR2_X1  g487(.A(new_n687), .B(new_n688), .ZN(G1327gat));
  INV_X1    g488(.A(KEYINPUT44), .ZN(new_n690));
  NAND2_X1  g489(.A1(new_n465), .A2(new_n467), .ZN(new_n691));
  OAI21_X1  g490(.A(new_n691), .B1(new_n679), .B2(new_n483), .ZN(new_n692));
  NAND2_X1  g491(.A1(new_n525), .A2(new_n526), .ZN(new_n693));
  INV_X1    g492(.A(KEYINPUT91), .ZN(new_n694));
  AOI21_X1  g493(.A(new_n692), .B1(new_n693), .B2(new_n694), .ZN(new_n695));
  NAND2_X1  g494(.A1(new_n522), .A2(KEYINPUT91), .ZN(new_n696));
  AOI22_X1  g495(.A1(new_n695), .A2(new_n696), .B1(new_n466), .B2(new_n479), .ZN(new_n697));
  OAI21_X1  g496(.A(new_n690), .B1(new_n697), .B2(new_n640), .ZN(new_n698));
  INV_X1    g497(.A(new_n464), .ZN(new_n699));
  INV_X1    g498(.A(new_n640), .ZN(new_n700));
  NAND3_X1  g499(.A1(new_n528), .A2(KEYINPUT44), .A3(new_n700), .ZN(new_n701));
  XNOR2_X1  g500(.A(new_n613), .B(KEYINPUT110), .ZN(new_n702));
  INV_X1    g501(.A(new_n702), .ZN(new_n703));
  AND2_X1   g502(.A1(new_n575), .A2(new_n576), .ZN(new_n704));
  XOR2_X1   g503(.A(new_n665), .B(KEYINPUT111), .Z(new_n705));
  INV_X1    g504(.A(new_n705), .ZN(new_n706));
  NOR3_X1   g505(.A1(new_n703), .A2(new_n704), .A3(new_n706), .ZN(new_n707));
  NAND4_X1  g506(.A1(new_n698), .A2(new_n699), .A3(new_n701), .A4(new_n707), .ZN(new_n708));
  NAND2_X1  g507(.A1(new_n708), .A2(G29gat), .ZN(new_n709));
  NOR2_X1   g508(.A1(new_n613), .A2(new_n640), .ZN(new_n710));
  NAND2_X1  g509(.A1(new_n710), .A2(new_n667), .ZN(new_n711));
  XOR2_X1   g510(.A(new_n711), .B(KEYINPUT108), .Z(new_n712));
  NOR2_X1   g511(.A1(new_n464), .A2(G29gat), .ZN(new_n713));
  NAND4_X1  g512(.A1(new_n712), .A2(new_n528), .A3(new_n577), .A4(new_n713), .ZN(new_n714));
  XOR2_X1   g513(.A(KEYINPUT109), .B(KEYINPUT45), .Z(new_n715));
  XNOR2_X1  g514(.A(new_n714), .B(new_n715), .ZN(new_n716));
  NAND2_X1  g515(.A1(new_n709), .A2(new_n716), .ZN(new_n717));
  NAND2_X1  g516(.A1(new_n717), .A2(KEYINPUT112), .ZN(new_n718));
  INV_X1    g517(.A(KEYINPUT112), .ZN(new_n719));
  NAND3_X1  g518(.A1(new_n709), .A2(new_n716), .A3(new_n719), .ZN(new_n720));
  NAND2_X1  g519(.A1(new_n718), .A2(new_n720), .ZN(G1328gat));
  NAND2_X1  g520(.A1(new_n693), .A2(new_n694), .ZN(new_n722));
  NAND3_X1  g521(.A1(new_n722), .A2(new_n696), .A3(new_n485), .ZN(new_n723));
  AOI21_X1  g522(.A(new_n704), .B1(new_n723), .B2(new_n480), .ZN(new_n724));
  NOR2_X1   g523(.A1(new_n419), .A2(G36gat), .ZN(new_n725));
  NAND3_X1  g524(.A1(new_n724), .A2(new_n712), .A3(new_n725), .ZN(new_n726));
  AND2_X1   g525(.A1(new_n726), .A2(KEYINPUT113), .ZN(new_n727));
  NOR2_X1   g526(.A1(new_n726), .A2(KEYINPUT113), .ZN(new_n728));
  INV_X1    g527(.A(KEYINPUT46), .ZN(new_n729));
  OR3_X1    g528(.A1(new_n727), .A2(new_n728), .A3(new_n729), .ZN(new_n730));
  AND2_X1   g529(.A1(new_n698), .A2(new_n701), .ZN(new_n731));
  NAND3_X1  g530(.A1(new_n731), .A2(new_n418), .A3(new_n707), .ZN(new_n732));
  NAND2_X1  g531(.A1(new_n732), .A2(G36gat), .ZN(new_n733));
  OAI21_X1  g532(.A(new_n729), .B1(new_n727), .B2(new_n728), .ZN(new_n734));
  NAND3_X1  g533(.A1(new_n730), .A2(new_n733), .A3(new_n734), .ZN(G1329gat));
  NOR2_X1   g534(.A1(new_n681), .A2(new_n541), .ZN(new_n736));
  NAND4_X1  g535(.A1(new_n698), .A2(new_n701), .A3(new_n707), .A4(new_n736), .ZN(new_n737));
  INV_X1    g536(.A(new_n470), .ZN(new_n738));
  AND3_X1   g537(.A1(new_n724), .A2(new_n738), .A3(new_n712), .ZN(new_n739));
  OAI21_X1  g538(.A(new_n737), .B1(G43gat), .B2(new_n739), .ZN(new_n740));
  XNOR2_X1  g539(.A(new_n740), .B(KEYINPUT47), .ZN(G1330gat));
  NAND4_X1  g540(.A1(new_n698), .A2(new_n467), .A3(new_n701), .A4(new_n707), .ZN(new_n742));
  INV_X1    g541(.A(KEYINPUT114), .ZN(new_n743));
  INV_X1    g542(.A(new_n542), .ZN(new_n744));
  NAND3_X1  g543(.A1(new_n742), .A2(new_n743), .A3(new_n744), .ZN(new_n745));
  NOR2_X1   g544(.A1(new_n394), .A2(new_n744), .ZN(new_n746));
  NAND4_X1  g545(.A1(new_n712), .A2(new_n528), .A3(new_n577), .A4(new_n746), .ZN(new_n747));
  XNOR2_X1  g546(.A(new_n747), .B(KEYINPUT115), .ZN(new_n748));
  NAND2_X1  g547(.A1(new_n745), .A2(new_n748), .ZN(new_n749));
  INV_X1    g548(.A(KEYINPUT48), .ZN(new_n750));
  NAND2_X1  g549(.A1(new_n749), .A2(new_n750), .ZN(new_n751));
  AOI22_X1  g550(.A1(new_n742), .A2(new_n744), .B1(new_n743), .B2(new_n750), .ZN(new_n752));
  INV_X1    g551(.A(KEYINPUT116), .ZN(new_n753));
  AND2_X1   g552(.A1(new_n747), .A2(new_n753), .ZN(new_n754));
  NOR2_X1   g553(.A1(new_n747), .A2(new_n753), .ZN(new_n755));
  OAI21_X1  g554(.A(KEYINPUT48), .B1(new_n754), .B2(new_n755), .ZN(new_n756));
  NAND2_X1  g555(.A1(new_n752), .A2(new_n756), .ZN(new_n757));
  NAND2_X1  g556(.A1(new_n751), .A2(new_n757), .ZN(G1331gat));
  NOR4_X1   g557(.A1(new_n697), .A2(new_n577), .A3(new_n641), .A4(new_n705), .ZN(new_n759));
  NAND2_X1  g558(.A1(new_n759), .A2(new_n699), .ZN(new_n760));
  XNOR2_X1  g559(.A(new_n760), .B(G57gat), .ZN(G1332gat));
  XNOR2_X1  g560(.A(new_n418), .B(KEYINPUT117), .ZN(new_n762));
  NAND2_X1  g561(.A1(new_n759), .A2(new_n762), .ZN(new_n763));
  OAI21_X1  g562(.A(new_n763), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n764));
  XOR2_X1   g563(.A(KEYINPUT49), .B(G64gat), .Z(new_n765));
  OAI21_X1  g564(.A(new_n764), .B1(new_n763), .B2(new_n765), .ZN(G1333gat));
  NAND2_X1  g565(.A1(new_n759), .A2(new_n680), .ZN(new_n767));
  NAND2_X1  g566(.A1(new_n767), .A2(G71gat), .ZN(new_n768));
  INV_X1    g567(.A(G71gat), .ZN(new_n769));
  NAND3_X1  g568(.A1(new_n759), .A2(new_n769), .A3(new_n738), .ZN(new_n770));
  NAND2_X1  g569(.A1(new_n768), .A2(new_n770), .ZN(new_n771));
  INV_X1    g570(.A(KEYINPUT50), .ZN(new_n772));
  NAND2_X1  g571(.A1(new_n771), .A2(new_n772), .ZN(new_n773));
  NAND3_X1  g572(.A1(new_n768), .A2(KEYINPUT50), .A3(new_n770), .ZN(new_n774));
  NAND2_X1  g573(.A1(new_n773), .A2(new_n774), .ZN(G1334gat));
  NAND2_X1  g574(.A1(new_n759), .A2(new_n467), .ZN(new_n776));
  XNOR2_X1  g575(.A(new_n776), .B(G78gat), .ZN(G1335gat));
  NOR3_X1   g576(.A1(new_n613), .A2(new_n577), .A3(new_n667), .ZN(new_n778));
  NAND2_X1  g577(.A1(new_n731), .A2(new_n778), .ZN(new_n779));
  OAI21_X1  g578(.A(G85gat), .B1(new_n779), .B2(new_n464), .ZN(new_n780));
  NAND3_X1  g579(.A1(new_n528), .A2(new_n704), .A3(new_n710), .ZN(new_n781));
  INV_X1    g580(.A(KEYINPUT51), .ZN(new_n782));
  NAND2_X1  g581(.A1(new_n781), .A2(new_n782), .ZN(new_n783));
  NAND4_X1  g582(.A1(new_n528), .A2(KEYINPUT51), .A3(new_n704), .A4(new_n710), .ZN(new_n784));
  NAND2_X1  g583(.A1(new_n783), .A2(new_n784), .ZN(new_n785));
  NAND4_X1  g584(.A1(new_n785), .A2(new_n617), .A3(new_n699), .A4(new_n665), .ZN(new_n786));
  NAND2_X1  g585(.A1(new_n780), .A2(new_n786), .ZN(G1336gat));
  NAND4_X1  g586(.A1(new_n698), .A2(new_n701), .A3(new_n762), .A4(new_n778), .ZN(new_n788));
  NAND2_X1  g587(.A1(new_n788), .A2(G92gat), .ZN(new_n789));
  AND3_X1   g588(.A1(new_n706), .A2(new_n618), .A3(new_n762), .ZN(new_n790));
  NAND2_X1  g589(.A1(new_n785), .A2(new_n790), .ZN(new_n791));
  INV_X1    g590(.A(KEYINPUT52), .ZN(new_n792));
  NAND3_X1  g591(.A1(new_n789), .A2(new_n791), .A3(new_n792), .ZN(new_n793));
  NAND4_X1  g592(.A1(new_n698), .A2(new_n418), .A3(new_n701), .A4(new_n778), .ZN(new_n794));
  AOI22_X1  g593(.A1(G92gat), .A2(new_n794), .B1(new_n785), .B2(new_n790), .ZN(new_n795));
  OAI21_X1  g594(.A(new_n793), .B1(new_n795), .B2(new_n792), .ZN(G1337gat));
  OAI21_X1  g595(.A(G99gat), .B1(new_n779), .B2(new_n681), .ZN(new_n797));
  NOR2_X1   g596(.A1(new_n470), .A2(G99gat), .ZN(new_n798));
  NAND3_X1  g597(.A1(new_n785), .A2(new_n665), .A3(new_n798), .ZN(new_n799));
  NAND2_X1  g598(.A1(new_n797), .A2(new_n799), .ZN(G1338gat));
  NAND4_X1  g599(.A1(new_n698), .A2(new_n467), .A3(new_n701), .A4(new_n778), .ZN(new_n801));
  NAND2_X1  g600(.A1(new_n801), .A2(G106gat), .ZN(new_n802));
  NAND2_X1  g601(.A1(KEYINPUT118), .A2(KEYINPUT53), .ZN(new_n803));
  NOR3_X1   g602(.A1(new_n705), .A2(G106gat), .A3(new_n394), .ZN(new_n804));
  AOI21_X1  g603(.A(new_n577), .B1(new_n723), .B2(new_n480), .ZN(new_n805));
  AOI21_X1  g604(.A(KEYINPUT51), .B1(new_n805), .B2(new_n710), .ZN(new_n806));
  INV_X1    g605(.A(new_n784), .ZN(new_n807));
  OAI21_X1  g606(.A(new_n804), .B1(new_n806), .B2(new_n807), .ZN(new_n808));
  NOR2_X1   g607(.A1(KEYINPUT118), .A2(KEYINPUT53), .ZN(new_n809));
  XNOR2_X1  g608(.A(new_n809), .B(KEYINPUT119), .ZN(new_n810));
  AND4_X1   g609(.A1(new_n802), .A2(new_n803), .A3(new_n808), .A4(new_n810), .ZN(new_n811));
  INV_X1    g610(.A(new_n803), .ZN(new_n812));
  AOI21_X1  g611(.A(new_n812), .B1(new_n785), .B2(new_n804), .ZN(new_n813));
  AOI21_X1  g612(.A(new_n810), .B1(new_n813), .B2(new_n802), .ZN(new_n814));
  NOR2_X1   g613(.A1(new_n811), .A2(new_n814), .ZN(G1339gat));
  AOI21_X1  g614(.A(new_n566), .B1(new_n564), .B2(new_n567), .ZN(new_n816));
  INV_X1    g615(.A(KEYINPUT122), .ZN(new_n817));
  AND2_X1   g616(.A1(new_n816), .A2(new_n817), .ZN(new_n818));
  NAND2_X1  g617(.A1(new_n554), .A2(new_n558), .ZN(new_n819));
  INV_X1    g618(.A(new_n555), .ZN(new_n820));
  NAND2_X1  g619(.A1(new_n819), .A2(new_n820), .ZN(new_n821));
  OAI21_X1  g620(.A(new_n821), .B1(new_n816), .B2(new_n817), .ZN(new_n822));
  OAI21_X1  g621(.A(new_n573), .B1(new_n818), .B2(new_n822), .ZN(new_n823));
  AND2_X1   g622(.A1(new_n823), .A2(new_n576), .ZN(new_n824));
  AND3_X1   g623(.A1(new_n824), .A2(KEYINPUT123), .A3(new_n665), .ZN(new_n825));
  AOI21_X1  g624(.A(KEYINPUT123), .B1(new_n824), .B2(new_n665), .ZN(new_n826));
  NOR2_X1   g625(.A1(new_n825), .A2(new_n826), .ZN(new_n827));
  NOR2_X1   g626(.A1(new_n654), .A2(new_n660), .ZN(new_n828));
  INV_X1    g627(.A(KEYINPUT54), .ZN(new_n829));
  AOI21_X1  g628(.A(new_n659), .B1(new_n661), .B2(new_n829), .ZN(new_n830));
  NAND3_X1  g629(.A1(new_n648), .A2(new_n649), .A3(new_n653), .ZN(new_n831));
  NAND2_X1  g630(.A1(new_n831), .A2(KEYINPUT54), .ZN(new_n832));
  OAI21_X1  g631(.A(new_n830), .B1(new_n654), .B2(new_n832), .ZN(new_n833));
  INV_X1    g632(.A(KEYINPUT55), .ZN(new_n834));
  AOI21_X1  g633(.A(new_n828), .B1(new_n833), .B2(new_n834), .ZN(new_n835));
  INV_X1    g634(.A(KEYINPUT121), .ZN(new_n836));
  NAND2_X1  g635(.A1(new_n648), .A2(new_n649), .ZN(new_n837));
  NAND3_X1  g636(.A1(new_n837), .A2(new_n829), .A3(new_n652), .ZN(new_n838));
  INV_X1    g637(.A(new_n659), .ZN(new_n839));
  NAND2_X1  g638(.A1(new_n838), .A2(new_n839), .ZN(new_n840));
  INV_X1    g639(.A(KEYINPUT104), .ZN(new_n841));
  AOI21_X1  g640(.A(new_n653), .B1(new_n837), .B2(new_n841), .ZN(new_n842));
  NAND3_X1  g641(.A1(new_n648), .A2(KEYINPUT104), .A3(new_n649), .ZN(new_n843));
  NAND2_X1  g642(.A1(new_n842), .A2(new_n843), .ZN(new_n844));
  INV_X1    g643(.A(new_n832), .ZN(new_n845));
  AOI21_X1  g644(.A(new_n840), .B1(new_n844), .B2(new_n845), .ZN(new_n846));
  AOI21_X1  g645(.A(new_n836), .B1(new_n846), .B2(KEYINPUT55), .ZN(new_n847));
  AOI21_X1  g646(.A(new_n832), .B1(new_n842), .B2(new_n843), .ZN(new_n848));
  NOR4_X1   g647(.A1(new_n848), .A2(new_n840), .A3(KEYINPUT121), .A4(new_n834), .ZN(new_n849));
  OAI211_X1 g648(.A(new_n577), .B(new_n835), .C1(new_n847), .C2(new_n849), .ZN(new_n850));
  AOI21_X1  g649(.A(new_n700), .B1(new_n827), .B2(new_n850), .ZN(new_n851));
  NAND2_X1  g650(.A1(new_n823), .A2(new_n576), .ZN(new_n852));
  NOR2_X1   g651(.A1(new_n640), .A2(new_n852), .ZN(new_n853));
  OAI211_X1 g652(.A(new_n853), .B(new_n835), .C1(new_n847), .C2(new_n849), .ZN(new_n854));
  INV_X1    g653(.A(new_n854), .ZN(new_n855));
  OAI21_X1  g654(.A(new_n702), .B1(new_n851), .B2(new_n855), .ZN(new_n856));
  NAND4_X1  g655(.A1(new_n704), .A2(new_n613), .A3(new_n640), .A4(new_n667), .ZN(new_n857));
  INV_X1    g656(.A(KEYINPUT120), .ZN(new_n858));
  XNOR2_X1  g657(.A(new_n857), .B(new_n858), .ZN(new_n859));
  NAND2_X1  g658(.A1(new_n856), .A2(new_n859), .ZN(new_n860));
  NOR2_X1   g659(.A1(new_n762), .A2(new_n464), .ZN(new_n861));
  INV_X1    g660(.A(new_n861), .ZN(new_n862));
  NOR2_X1   g661(.A1(new_n862), .A2(new_n395), .ZN(new_n863));
  NAND2_X1  g662(.A1(new_n860), .A2(new_n863), .ZN(new_n864));
  INV_X1    g663(.A(new_n864), .ZN(new_n865));
  AOI21_X1  g664(.A(G113gat), .B1(new_n865), .B2(new_n577), .ZN(new_n866));
  AND3_X1   g665(.A1(new_n860), .A2(new_n471), .A3(new_n861), .ZN(new_n867));
  NOR2_X1   g666(.A1(new_n704), .A2(new_n255), .ZN(new_n868));
  AOI21_X1  g667(.A(new_n866), .B1(new_n867), .B2(new_n868), .ZN(G1340gat));
  AOI21_X1  g668(.A(G120gat), .B1(new_n865), .B2(new_n665), .ZN(new_n870));
  NOR2_X1   g669(.A1(new_n705), .A2(new_n256), .ZN(new_n871));
  AOI21_X1  g670(.A(new_n870), .B1(new_n867), .B2(new_n871), .ZN(G1341gat));
  NAND3_X1  g671(.A1(new_n865), .A2(new_n266), .A3(new_n613), .ZN(new_n873));
  AND2_X1   g672(.A1(new_n867), .A2(new_n703), .ZN(new_n874));
  OAI21_X1  g673(.A(new_n873), .B1(new_n874), .B2(new_n266), .ZN(G1342gat));
  AND4_X1   g674(.A1(new_n699), .A2(new_n860), .A3(new_n419), .A4(new_n700), .ZN(new_n876));
  NOR2_X1   g675(.A1(new_n395), .A2(G134gat), .ZN(new_n877));
  NAND2_X1  g676(.A1(new_n876), .A2(new_n877), .ZN(new_n878));
  INV_X1    g677(.A(KEYINPUT56), .ZN(new_n879));
  XNOR2_X1  g678(.A(new_n878), .B(new_n879), .ZN(new_n880));
  NAND2_X1  g679(.A1(new_n867), .A2(new_n700), .ZN(new_n881));
  NAND2_X1  g680(.A1(new_n881), .A2(G134gat), .ZN(new_n882));
  NAND2_X1  g681(.A1(new_n880), .A2(new_n882), .ZN(G1343gat));
  AOI21_X1  g682(.A(new_n394), .B1(new_n856), .B2(new_n859), .ZN(new_n884));
  NOR2_X1   g683(.A1(new_n862), .A2(new_n680), .ZN(new_n885));
  AND2_X1   g684(.A1(new_n884), .A2(new_n885), .ZN(new_n886));
  INV_X1    g685(.A(G141gat), .ZN(new_n887));
  NAND3_X1  g686(.A1(new_n886), .A2(new_n887), .A3(new_n577), .ZN(new_n888));
  INV_X1    g687(.A(new_n613), .ZN(new_n889));
  NAND2_X1  g688(.A1(new_n824), .A2(new_n665), .ZN(new_n890));
  AOI21_X1  g689(.A(new_n700), .B1(new_n850), .B2(new_n890), .ZN(new_n891));
  OAI21_X1  g690(.A(new_n889), .B1(new_n891), .B2(new_n855), .ZN(new_n892));
  AOI21_X1  g691(.A(new_n394), .B1(new_n892), .B2(new_n859), .ZN(new_n893));
  INV_X1    g692(.A(KEYINPUT57), .ZN(new_n894));
  OAI21_X1  g693(.A(new_n885), .B1(new_n893), .B2(new_n894), .ZN(new_n895));
  AOI211_X1 g694(.A(KEYINPUT57), .B(new_n394), .C1(new_n856), .C2(new_n859), .ZN(new_n896));
  NOR3_X1   g695(.A1(new_n895), .A2(new_n896), .A3(new_n704), .ZN(new_n897));
  OAI21_X1  g696(.A(new_n888), .B1(new_n897), .B2(new_n887), .ZN(new_n898));
  NAND2_X1  g697(.A1(new_n898), .A2(KEYINPUT58), .ZN(new_n899));
  INV_X1    g698(.A(KEYINPUT58), .ZN(new_n900));
  OAI211_X1 g699(.A(new_n900), .B(new_n888), .C1(new_n897), .C2(new_n887), .ZN(new_n901));
  NAND2_X1  g700(.A1(new_n899), .A2(new_n901), .ZN(G1344gat));
  INV_X1    g701(.A(G148gat), .ZN(new_n903));
  NAND3_X1  g702(.A1(new_n886), .A2(new_n903), .A3(new_n665), .ZN(new_n904));
  NOR3_X1   g703(.A1(new_n895), .A2(new_n896), .A3(new_n667), .ZN(new_n905));
  NOR3_X1   g704(.A1(new_n905), .A2(KEYINPUT59), .A3(new_n903), .ZN(new_n906));
  INV_X1    g705(.A(KEYINPUT59), .ZN(new_n907));
  NAND2_X1  g706(.A1(new_n860), .A2(new_n467), .ZN(new_n908));
  NAND2_X1  g707(.A1(new_n908), .A2(KEYINPUT57), .ZN(new_n909));
  NAND3_X1  g708(.A1(new_n666), .A2(new_n704), .A3(new_n668), .ZN(new_n910));
  NAND2_X1  g709(.A1(new_n892), .A2(new_n910), .ZN(new_n911));
  NAND3_X1  g710(.A1(new_n911), .A2(new_n894), .A3(new_n467), .ZN(new_n912));
  NAND4_X1  g711(.A1(new_n909), .A2(new_n665), .A3(new_n885), .A4(new_n912), .ZN(new_n913));
  AOI21_X1  g712(.A(new_n907), .B1(new_n913), .B2(G148gat), .ZN(new_n914));
  OAI21_X1  g713(.A(new_n904), .B1(new_n906), .B2(new_n914), .ZN(G1345gat));
  NAND3_X1  g714(.A1(new_n886), .A2(new_n340), .A3(new_n613), .ZN(new_n916));
  NOR3_X1   g715(.A1(new_n895), .A2(new_n896), .A3(new_n702), .ZN(new_n917));
  OAI21_X1  g716(.A(new_n916), .B1(new_n917), .B2(new_n340), .ZN(G1346gat));
  NOR2_X1   g717(.A1(new_n680), .A2(new_n394), .ZN(new_n919));
  NAND3_X1  g718(.A1(new_n876), .A2(new_n329), .A3(new_n919), .ZN(new_n920));
  NOR3_X1   g719(.A1(new_n895), .A2(new_n896), .A3(new_n640), .ZN(new_n921));
  OAI21_X1  g720(.A(new_n920), .B1(new_n921), .B2(new_n329), .ZN(G1347gat));
  NAND4_X1  g721(.A1(new_n860), .A2(new_n464), .A3(new_n418), .A4(new_n471), .ZN(new_n923));
  NOR3_X1   g722(.A1(new_n923), .A2(new_n213), .A3(new_n704), .ZN(new_n924));
  AOI21_X1  g723(.A(new_n699), .B1(new_n856), .B2(new_n859), .ZN(new_n925));
  NAND3_X1  g724(.A1(new_n762), .A2(new_n394), .A3(new_n313), .ZN(new_n926));
  XOR2_X1   g725(.A(new_n926), .B(KEYINPUT124), .Z(new_n927));
  NAND2_X1  g726(.A1(new_n925), .A2(new_n927), .ZN(new_n928));
  INV_X1    g727(.A(new_n928), .ZN(new_n929));
  NAND2_X1  g728(.A1(new_n929), .A2(new_n577), .ZN(new_n930));
  AOI21_X1  g729(.A(new_n924), .B1(new_n930), .B2(new_n213), .ZN(G1348gat));
  OAI21_X1  g730(.A(G176gat), .B1(new_n923), .B2(new_n705), .ZN(new_n932));
  NAND2_X1  g731(.A1(new_n665), .A2(new_n214), .ZN(new_n933));
  OAI21_X1  g732(.A(new_n932), .B1(new_n928), .B2(new_n933), .ZN(G1349gat));
  NAND3_X1  g733(.A1(new_n929), .A2(new_n247), .A3(new_n613), .ZN(new_n935));
  OAI21_X1  g734(.A(G183gat), .B1(new_n923), .B2(new_n702), .ZN(new_n936));
  NAND3_X1  g735(.A1(new_n935), .A2(KEYINPUT125), .A3(new_n936), .ZN(new_n937));
  NAND2_X1  g736(.A1(new_n937), .A2(KEYINPUT60), .ZN(new_n938));
  INV_X1    g737(.A(KEYINPUT60), .ZN(new_n939));
  NAND4_X1  g738(.A1(new_n935), .A2(KEYINPUT125), .A3(new_n939), .A4(new_n936), .ZN(new_n940));
  NAND2_X1  g739(.A1(new_n938), .A2(new_n940), .ZN(G1350gat));
  NAND3_X1  g740(.A1(new_n929), .A2(new_n205), .A3(new_n700), .ZN(new_n942));
  OAI21_X1  g741(.A(G190gat), .B1(new_n923), .B2(new_n640), .ZN(new_n943));
  AND2_X1   g742(.A1(new_n943), .A2(KEYINPUT61), .ZN(new_n944));
  NOR2_X1   g743(.A1(new_n943), .A2(KEYINPUT61), .ZN(new_n945));
  OAI21_X1  g744(.A(new_n942), .B1(new_n944), .B2(new_n945), .ZN(G1351gat));
  AND2_X1   g745(.A1(new_n919), .A2(new_n762), .ZN(new_n947));
  NAND2_X1  g746(.A1(new_n925), .A2(new_n947), .ZN(new_n948));
  INV_X1    g747(.A(new_n948), .ZN(new_n949));
  AOI21_X1  g748(.A(G197gat), .B1(new_n949), .B2(new_n577), .ZN(new_n950));
  NOR3_X1   g749(.A1(new_n680), .A2(new_n699), .A3(new_n419), .ZN(new_n951));
  AND3_X1   g750(.A1(new_n909), .A2(new_n912), .A3(new_n951), .ZN(new_n952));
  AND2_X1   g751(.A1(new_n577), .A2(G197gat), .ZN(new_n953));
  AOI21_X1  g752(.A(new_n950), .B1(new_n952), .B2(new_n953), .ZN(G1352gat));
  NOR3_X1   g753(.A1(new_n948), .A2(G204gat), .A3(new_n667), .ZN(new_n955));
  XNOR2_X1  g754(.A(new_n955), .B(KEYINPUT62), .ZN(new_n956));
  NAND3_X1  g755(.A1(new_n909), .A2(new_n912), .A3(new_n951), .ZN(new_n957));
  OAI21_X1  g756(.A(G204gat), .B1(new_n957), .B2(new_n705), .ZN(new_n958));
  NAND2_X1  g757(.A1(new_n956), .A2(new_n958), .ZN(G1353gat));
  NAND3_X1  g758(.A1(new_n949), .A2(new_n358), .A3(new_n613), .ZN(new_n960));
  NAND4_X1  g759(.A1(new_n909), .A2(new_n613), .A3(new_n912), .A4(new_n951), .ZN(new_n961));
  NAND3_X1  g760(.A1(new_n961), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n962));
  INV_X1    g761(.A(new_n962), .ZN(new_n963));
  AOI21_X1  g762(.A(KEYINPUT63), .B1(new_n961), .B2(G211gat), .ZN(new_n964));
  OAI21_X1  g763(.A(new_n960), .B1(new_n963), .B2(new_n964), .ZN(G1354gat));
  NAND2_X1  g764(.A1(new_n700), .A2(new_n351), .ZN(new_n966));
  INV_X1    g765(.A(KEYINPUT127), .ZN(new_n967));
  AOI21_X1  g766(.A(new_n966), .B1(new_n952), .B2(new_n967), .ZN(new_n968));
  NAND2_X1  g767(.A1(new_n957), .A2(KEYINPUT127), .ZN(new_n969));
  INV_X1    g768(.A(G218gat), .ZN(new_n970));
  OAI21_X1  g769(.A(new_n970), .B1(new_n948), .B2(new_n640), .ZN(new_n971));
  INV_X1    g770(.A(KEYINPUT126), .ZN(new_n972));
  OR2_X1    g771(.A1(new_n971), .A2(new_n972), .ZN(new_n973));
  NAND2_X1  g772(.A1(new_n971), .A2(new_n972), .ZN(new_n974));
  AOI22_X1  g773(.A1(new_n968), .A2(new_n969), .B1(new_n973), .B2(new_n974), .ZN(G1355gat));
endmodule


