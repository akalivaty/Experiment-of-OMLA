//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 1 1 1 0 0 0 1 1 1 1 1 1 1 0 0 0 1 1 0 1 1 1 1 0 0 0 1 0 1 0 0 1 0 1 0 1 0 0 1 1 1 1 1 0 1 0 1 1 1 0 0 1 1 0 0 1 0 0 0 1 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:25:23 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n681, new_n682, new_n683, new_n684, new_n685,
    new_n686, new_n687, new_n689, new_n690, new_n691, new_n692, new_n693,
    new_n694, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n731,
    new_n732, new_n733, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n743, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n752, new_n753, new_n754, new_n755, new_n756,
    new_n757, new_n758, new_n759, new_n760, new_n761, new_n762, new_n763,
    new_n764, new_n765, new_n767, new_n768, new_n769, new_n770, new_n771,
    new_n772, new_n773, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n799, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n823, new_n824,
    new_n825, new_n826, new_n827, new_n828, new_n829, new_n830, new_n831,
    new_n832, new_n833, new_n834, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n945,
    new_n946, new_n947, new_n948, new_n949, new_n950, new_n951, new_n952,
    new_n953, new_n955, new_n956, new_n957, new_n958, new_n959, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n967, new_n968, new_n969,
    new_n970, new_n971, new_n972, new_n974, new_n975, new_n976, new_n977,
    new_n978, new_n979, new_n980, new_n981, new_n982, new_n983, new_n985,
    new_n986, new_n987, new_n988, new_n989, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1015, new_n1016, new_n1017, new_n1018, new_n1019,
    new_n1020, new_n1021, new_n1022, new_n1023, new_n1024;
  INV_X1    g000(.A(KEYINPUT97), .ZN(new_n187));
  OAI21_X1  g001(.A(G210), .B1(G237), .B2(G902), .ZN(new_n188));
  INV_X1    g002(.A(new_n188), .ZN(new_n189));
  INV_X1    g003(.A(G146), .ZN(new_n190));
  NAND2_X1  g004(.A1(new_n190), .A2(G143), .ZN(new_n191));
  INV_X1    g005(.A(G143), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n192), .A2(G146), .ZN(new_n193));
  NAND4_X1  g007(.A1(new_n191), .A2(new_n193), .A3(KEYINPUT0), .A4(G128), .ZN(new_n194));
  XNOR2_X1  g008(.A(G143), .B(G146), .ZN(new_n195));
  XNOR2_X1  g009(.A(KEYINPUT0), .B(G128), .ZN(new_n196));
  OAI211_X1 g010(.A(new_n194), .B(G125), .C1(new_n195), .C2(new_n196), .ZN(new_n197));
  INV_X1    g011(.A(new_n197), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n191), .A2(new_n193), .ZN(new_n199));
  INV_X1    g013(.A(KEYINPUT1), .ZN(new_n200));
  AOI21_X1  g014(.A(new_n200), .B1(G143), .B2(new_n190), .ZN(new_n201));
  INV_X1    g015(.A(G128), .ZN(new_n202));
  OAI21_X1  g016(.A(new_n199), .B1(new_n201), .B2(new_n202), .ZN(new_n203));
  NAND3_X1  g017(.A1(new_n195), .A2(new_n200), .A3(G128), .ZN(new_n204));
  AOI21_X1  g018(.A(G125), .B1(new_n203), .B2(new_n204), .ZN(new_n205));
  NOR2_X1   g019(.A1(new_n198), .A2(new_n205), .ZN(new_n206));
  INV_X1    g020(.A(G953), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n207), .A2(G224), .ZN(new_n208));
  XNOR2_X1  g022(.A(new_n206), .B(new_n208), .ZN(new_n209));
  XNOR2_X1  g023(.A(G110), .B(G122), .ZN(new_n210));
  INV_X1    g024(.A(new_n210), .ZN(new_n211));
  INV_X1    g025(.A(KEYINPUT6), .ZN(new_n212));
  NOR2_X1   g026(.A1(new_n212), .A2(KEYINPUT91), .ZN(new_n213));
  INV_X1    g027(.A(KEYINPUT90), .ZN(new_n214));
  OR2_X1    g028(.A1(KEYINPUT66), .A2(G119), .ZN(new_n215));
  NAND2_X1  g029(.A1(KEYINPUT66), .A2(G119), .ZN(new_n216));
  NAND3_X1  g030(.A1(new_n215), .A2(G116), .A3(new_n216), .ZN(new_n217));
  OR2_X1    g031(.A1(KEYINPUT67), .A2(G116), .ZN(new_n218));
  NAND2_X1  g032(.A1(KEYINPUT67), .A2(G116), .ZN(new_n219));
  NAND3_X1  g033(.A1(new_n218), .A2(G119), .A3(new_n219), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n217), .A2(new_n220), .ZN(new_n221));
  XNOR2_X1  g035(.A(KEYINPUT2), .B(G113), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  INV_X1    g037(.A(new_n222), .ZN(new_n224));
  NAND3_X1  g038(.A1(new_n224), .A2(new_n217), .A3(new_n220), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n223), .A2(new_n225), .ZN(new_n226));
  INV_X1    g040(.A(G104), .ZN(new_n227));
  OAI21_X1  g041(.A(KEYINPUT3), .B1(new_n227), .B2(G107), .ZN(new_n228));
  INV_X1    g042(.A(KEYINPUT83), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n228), .A2(new_n229), .ZN(new_n230));
  OAI211_X1 g044(.A(KEYINPUT83), .B(KEYINPUT3), .C1(new_n227), .C2(G107), .ZN(new_n231));
  INV_X1    g045(.A(KEYINPUT3), .ZN(new_n232));
  INV_X1    g046(.A(G107), .ZN(new_n233));
  NAND3_X1  g047(.A1(new_n232), .A2(new_n233), .A3(G104), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n227), .A2(G107), .ZN(new_n235));
  NAND4_X1  g049(.A1(new_n230), .A2(new_n231), .A3(new_n234), .A4(new_n235), .ZN(new_n236));
  INV_X1    g050(.A(KEYINPUT4), .ZN(new_n237));
  NAND3_X1  g051(.A1(new_n236), .A2(new_n237), .A3(G101), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n226), .A2(new_n238), .ZN(new_n239));
  INV_X1    g053(.A(new_n239), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n236), .A2(G101), .ZN(new_n241));
  AND2_X1   g055(.A1(new_n234), .A2(new_n235), .ZN(new_n242));
  XNOR2_X1  g056(.A(KEYINPUT84), .B(G101), .ZN(new_n243));
  NAND4_X1  g057(.A1(new_n242), .A2(new_n243), .A3(new_n231), .A4(new_n230), .ZN(new_n244));
  NAND3_X1  g058(.A1(new_n241), .A2(KEYINPUT4), .A3(new_n244), .ZN(new_n245));
  AOI21_X1  g059(.A(new_n214), .B1(new_n240), .B2(new_n245), .ZN(new_n246));
  NAND4_X1  g060(.A1(new_n245), .A2(new_n214), .A3(new_n238), .A4(new_n226), .ZN(new_n247));
  INV_X1    g061(.A(KEYINPUT5), .ZN(new_n248));
  NAND4_X1  g062(.A1(new_n215), .A2(new_n248), .A3(G116), .A4(new_n216), .ZN(new_n249));
  OAI211_X1 g063(.A(G113), .B(new_n249), .C1(new_n221), .C2(new_n248), .ZN(new_n250));
  XNOR2_X1  g064(.A(G104), .B(G107), .ZN(new_n251));
  INV_X1    g065(.A(G101), .ZN(new_n252));
  OAI21_X1  g066(.A(KEYINPUT86), .B1(new_n251), .B2(new_n252), .ZN(new_n253));
  INV_X1    g067(.A(KEYINPUT86), .ZN(new_n254));
  NOR2_X1   g068(.A1(new_n227), .A2(G107), .ZN(new_n255));
  NOR2_X1   g069(.A1(new_n233), .A2(G104), .ZN(new_n256));
  OAI211_X1 g070(.A(new_n254), .B(G101), .C1(new_n255), .C2(new_n256), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n253), .A2(new_n257), .ZN(new_n258));
  NAND4_X1  g072(.A1(new_n250), .A2(new_n244), .A3(new_n258), .A4(new_n225), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n247), .A2(new_n259), .ZN(new_n260));
  OAI211_X1 g074(.A(new_n211), .B(new_n213), .C1(new_n246), .C2(new_n260), .ZN(new_n261));
  INV_X1    g075(.A(new_n261), .ZN(new_n262));
  AND3_X1   g076(.A1(new_n241), .A2(KEYINPUT4), .A3(new_n244), .ZN(new_n263));
  OAI21_X1  g077(.A(KEYINPUT90), .B1(new_n263), .B2(new_n239), .ZN(new_n264));
  NAND3_X1  g078(.A1(new_n264), .A2(new_n259), .A3(new_n247), .ZN(new_n265));
  AOI21_X1  g079(.A(new_n213), .B1(new_n265), .B2(new_n211), .ZN(new_n266));
  NOR2_X1   g080(.A1(new_n262), .A2(new_n266), .ZN(new_n267));
  INV_X1    g081(.A(new_n260), .ZN(new_n268));
  INV_X1    g082(.A(KEYINPUT92), .ZN(new_n269));
  NAND4_X1  g083(.A1(new_n268), .A2(new_n269), .A3(new_n210), .A4(new_n264), .ZN(new_n270));
  NAND4_X1  g084(.A1(new_n264), .A2(new_n210), .A3(new_n259), .A4(new_n247), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n271), .A2(KEYINPUT92), .ZN(new_n272));
  NAND3_X1  g086(.A1(new_n270), .A2(new_n272), .A3(KEYINPUT6), .ZN(new_n273));
  AOI21_X1  g087(.A(new_n209), .B1(new_n267), .B2(new_n273), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n270), .A2(new_n272), .ZN(new_n275));
  INV_X1    g089(.A(new_n206), .ZN(new_n276));
  NAND4_X1  g090(.A1(new_n276), .A2(KEYINPUT96), .A3(KEYINPUT7), .A4(new_n208), .ZN(new_n277));
  OAI211_X1 g091(.A(KEYINPUT7), .B(new_n208), .C1(new_n198), .C2(new_n205), .ZN(new_n278));
  INV_X1    g092(.A(KEYINPUT96), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n278), .A2(new_n279), .ZN(new_n280));
  INV_X1    g094(.A(KEYINPUT95), .ZN(new_n281));
  INV_X1    g095(.A(KEYINPUT7), .ZN(new_n282));
  AOI22_X1  g096(.A1(new_n281), .A2(new_n282), .B1(new_n207), .B2(G224), .ZN(new_n283));
  OAI21_X1  g097(.A(new_n283), .B1(new_n281), .B2(new_n282), .ZN(new_n284));
  AOI22_X1  g098(.A1(new_n277), .A2(new_n280), .B1(new_n206), .B2(new_n284), .ZN(new_n285));
  XOR2_X1   g099(.A(KEYINPUT93), .B(KEYINPUT8), .Z(new_n286));
  XNOR2_X1  g100(.A(new_n286), .B(new_n210), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n250), .A2(new_n225), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n258), .A2(new_n244), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n288), .A2(new_n289), .ZN(new_n290));
  INV_X1    g104(.A(KEYINPUT94), .ZN(new_n291));
  OAI21_X1  g105(.A(new_n290), .B1(new_n291), .B2(new_n259), .ZN(new_n292));
  AND2_X1   g106(.A1(new_n259), .A2(new_n291), .ZN(new_n293));
  OAI21_X1  g107(.A(new_n287), .B1(new_n292), .B2(new_n293), .ZN(new_n294));
  AND2_X1   g108(.A1(new_n285), .A2(new_n294), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n275), .A2(new_n295), .ZN(new_n296));
  INV_X1    g110(.A(G902), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n296), .A2(new_n297), .ZN(new_n298));
  OAI21_X1  g112(.A(new_n189), .B1(new_n274), .B2(new_n298), .ZN(new_n299));
  INV_X1    g113(.A(new_n209), .ZN(new_n300));
  AND3_X1   g114(.A1(new_n270), .A2(new_n272), .A3(KEYINPUT6), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n265), .A2(new_n211), .ZN(new_n302));
  INV_X1    g116(.A(new_n213), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n302), .A2(new_n303), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n304), .A2(new_n261), .ZN(new_n305));
  OAI21_X1  g119(.A(new_n300), .B1(new_n301), .B2(new_n305), .ZN(new_n306));
  AOI21_X1  g120(.A(G902), .B1(new_n275), .B2(new_n295), .ZN(new_n307));
  NAND3_X1  g121(.A1(new_n306), .A2(new_n307), .A3(new_n188), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n299), .A2(new_n308), .ZN(new_n309));
  OAI21_X1  g123(.A(G214), .B1(G237), .B2(G902), .ZN(new_n310));
  AOI21_X1  g124(.A(new_n187), .B1(new_n309), .B2(new_n310), .ZN(new_n311));
  INV_X1    g125(.A(new_n310), .ZN(new_n312));
  AOI211_X1 g126(.A(KEYINPUT97), .B(new_n312), .C1(new_n299), .C2(new_n308), .ZN(new_n313));
  INV_X1    g127(.A(G469), .ZN(new_n314));
  XNOR2_X1  g128(.A(G110), .B(G140), .ZN(new_n315));
  XNOR2_X1  g129(.A(new_n315), .B(KEYINPUT81), .ZN(new_n316));
  XNOR2_X1  g130(.A(KEYINPUT70), .B(G953), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n317), .A2(G227), .ZN(new_n318));
  XNOR2_X1  g132(.A(new_n316), .B(new_n318), .ZN(new_n319));
  INV_X1    g133(.A(KEYINPUT10), .ZN(new_n320));
  NOR3_X1   g134(.A1(new_n199), .A2(KEYINPUT1), .A3(new_n202), .ZN(new_n321));
  OAI21_X1  g135(.A(KEYINPUT1), .B1(new_n192), .B2(G146), .ZN(new_n322));
  INV_X1    g136(.A(KEYINPUT87), .ZN(new_n323));
  NAND2_X1  g137(.A1(new_n322), .A2(new_n323), .ZN(new_n324));
  NAND3_X1  g138(.A1(new_n191), .A2(KEYINPUT87), .A3(KEYINPUT1), .ZN(new_n325));
  NAND3_X1  g139(.A1(new_n324), .A2(G128), .A3(new_n325), .ZN(new_n326));
  AOI21_X1  g140(.A(new_n321), .B1(new_n326), .B2(new_n199), .ZN(new_n327));
  OAI21_X1  g141(.A(new_n320), .B1(new_n289), .B2(new_n327), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n203), .A2(new_n204), .ZN(new_n329));
  NAND4_X1  g143(.A1(new_n244), .A2(new_n258), .A3(new_n329), .A4(KEYINPUT10), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n328), .A2(new_n330), .ZN(new_n331));
  OAI21_X1  g145(.A(new_n194), .B1(new_n195), .B2(new_n196), .ZN(new_n332));
  INV_X1    g146(.A(new_n332), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n238), .A2(new_n333), .ZN(new_n334));
  OAI21_X1  g148(.A(KEYINPUT85), .B1(new_n263), .B2(new_n334), .ZN(new_n335));
  INV_X1    g149(.A(KEYINPUT85), .ZN(new_n336));
  NAND4_X1  g150(.A1(new_n245), .A2(new_n336), .A3(new_n333), .A4(new_n238), .ZN(new_n337));
  AOI21_X1  g151(.A(new_n331), .B1(new_n335), .B2(new_n337), .ZN(new_n338));
  INV_X1    g152(.A(G137), .ZN(new_n339));
  NAND3_X1  g153(.A1(new_n339), .A2(KEYINPUT11), .A3(G134), .ZN(new_n340));
  XNOR2_X1  g154(.A(KEYINPUT64), .B(G134), .ZN(new_n341));
  OAI21_X1  g155(.A(new_n340), .B1(new_n341), .B2(new_n339), .ZN(new_n342));
  INV_X1    g156(.A(new_n342), .ZN(new_n343));
  AND2_X1   g157(.A1(KEYINPUT64), .A2(G134), .ZN(new_n344));
  NOR2_X1   g158(.A1(KEYINPUT64), .A2(G134), .ZN(new_n345));
  OAI21_X1  g159(.A(new_n339), .B1(new_n344), .B2(new_n345), .ZN(new_n346));
  INV_X1    g160(.A(KEYINPUT11), .ZN(new_n347));
  AND3_X1   g161(.A1(new_n346), .A2(KEYINPUT65), .A3(new_n347), .ZN(new_n348));
  AOI21_X1  g162(.A(KEYINPUT65), .B1(new_n346), .B2(new_n347), .ZN(new_n349));
  OAI21_X1  g163(.A(new_n343), .B1(new_n348), .B2(new_n349), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n350), .A2(G131), .ZN(new_n351));
  INV_X1    g165(.A(KEYINPUT65), .ZN(new_n352));
  OR2_X1    g166(.A1(KEYINPUT64), .A2(G134), .ZN(new_n353));
  NAND2_X1  g167(.A1(KEYINPUT64), .A2(G134), .ZN(new_n354));
  AOI21_X1  g168(.A(G137), .B1(new_n353), .B2(new_n354), .ZN(new_n355));
  OAI21_X1  g169(.A(new_n352), .B1(new_n355), .B2(KEYINPUT11), .ZN(new_n356));
  NAND3_X1  g170(.A1(new_n346), .A2(KEYINPUT65), .A3(new_n347), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n356), .A2(new_n357), .ZN(new_n358));
  INV_X1    g172(.A(G131), .ZN(new_n359));
  NAND3_X1  g173(.A1(new_n358), .A2(new_n359), .A3(new_n343), .ZN(new_n360));
  NAND2_X1  g174(.A1(new_n351), .A2(new_n360), .ZN(new_n361));
  INV_X1    g175(.A(new_n361), .ZN(new_n362));
  AOI21_X1  g176(.A(new_n319), .B1(new_n338), .B2(new_n362), .ZN(new_n363));
  NAND3_X1  g177(.A1(new_n289), .A2(new_n204), .A3(new_n203), .ZN(new_n364));
  AOI21_X1  g178(.A(new_n202), .B1(new_n201), .B2(KEYINPUT87), .ZN(new_n365));
  AOI21_X1  g179(.A(new_n195), .B1(new_n365), .B2(new_n324), .ZN(new_n366));
  OAI211_X1 g180(.A(new_n244), .B(new_n258), .C1(new_n366), .C2(new_n321), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n364), .A2(new_n367), .ZN(new_n368));
  XNOR2_X1  g182(.A(KEYINPUT88), .B(KEYINPUT12), .ZN(new_n369));
  NAND3_X1  g183(.A1(new_n368), .A2(new_n361), .A3(new_n369), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n370), .A2(KEYINPUT89), .ZN(new_n371));
  INV_X1    g185(.A(KEYINPUT89), .ZN(new_n372));
  NAND4_X1  g186(.A1(new_n368), .A2(new_n361), .A3(new_n372), .A4(new_n369), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n368), .A2(new_n361), .ZN(new_n374));
  INV_X1    g188(.A(KEYINPUT12), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n374), .A2(new_n375), .ZN(new_n376));
  NAND3_X1  g190(.A1(new_n371), .A2(new_n373), .A3(new_n376), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n363), .A2(new_n377), .ZN(new_n378));
  INV_X1    g192(.A(new_n378), .ZN(new_n379));
  INV_X1    g193(.A(new_n319), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n335), .A2(new_n337), .ZN(new_n381));
  INV_X1    g195(.A(new_n331), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n381), .A2(new_n382), .ZN(new_n383));
  NAND2_X1  g197(.A1(new_n383), .A2(new_n361), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n338), .A2(new_n362), .ZN(new_n385));
  AOI21_X1  g199(.A(new_n380), .B1(new_n384), .B2(new_n385), .ZN(new_n386));
  OAI211_X1 g200(.A(new_n314), .B(new_n297), .C1(new_n379), .C2(new_n386), .ZN(new_n387));
  NOR2_X1   g201(.A1(new_n314), .A2(new_n297), .ZN(new_n388));
  INV_X1    g202(.A(new_n388), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n363), .A2(new_n384), .ZN(new_n390));
  AOI22_X1  g204(.A1(new_n370), .A2(KEYINPUT89), .B1(new_n374), .B2(new_n375), .ZN(new_n391));
  AOI22_X1  g205(.A1(new_n391), .A2(new_n373), .B1(new_n362), .B2(new_n338), .ZN(new_n392));
  XOR2_X1   g206(.A(new_n319), .B(KEYINPUT82), .Z(new_n393));
  OAI211_X1 g207(.A(new_n390), .B(G469), .C1(new_n392), .C2(new_n393), .ZN(new_n394));
  NAND3_X1  g208(.A1(new_n387), .A2(new_n389), .A3(new_n394), .ZN(new_n395));
  XOR2_X1   g209(.A(KEYINPUT9), .B(G234), .Z(new_n396));
  XNOR2_X1  g210(.A(new_n396), .B(KEYINPUT80), .ZN(new_n397));
  OAI21_X1  g211(.A(G221), .B1(new_n397), .B2(G902), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n395), .A2(new_n398), .ZN(new_n399));
  NOR3_X1   g213(.A1(new_n311), .A2(new_n313), .A3(new_n399), .ZN(new_n400));
  NOR2_X1   g214(.A1(new_n339), .A2(G134), .ZN(new_n401));
  OAI21_X1  g215(.A(G131), .B1(new_n355), .B2(new_n401), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n329), .A2(new_n402), .ZN(new_n403));
  AOI21_X1  g217(.A(new_n342), .B1(new_n356), .B2(new_n357), .ZN(new_n404));
  AOI21_X1  g218(.A(new_n403), .B1(new_n404), .B2(new_n359), .ZN(new_n405));
  AOI21_X1  g219(.A(new_n405), .B1(new_n361), .B2(new_n333), .ZN(new_n406));
  OAI21_X1  g220(.A(new_n226), .B1(new_n406), .B2(KEYINPUT30), .ZN(new_n407));
  INV_X1    g221(.A(new_n407), .ZN(new_n408));
  INV_X1    g222(.A(KEYINPUT68), .ZN(new_n409));
  NAND3_X1  g223(.A1(new_n406), .A2(new_n409), .A3(KEYINPUT30), .ZN(new_n410));
  INV_X1    g224(.A(new_n410), .ZN(new_n411));
  AOI21_X1  g225(.A(new_n409), .B1(new_n406), .B2(KEYINPUT30), .ZN(new_n412));
  OAI21_X1  g226(.A(new_n408), .B1(new_n411), .B2(new_n412), .ZN(new_n413));
  INV_X1    g227(.A(KEYINPUT29), .ZN(new_n414));
  AOI21_X1  g228(.A(new_n359), .B1(new_n358), .B2(new_n343), .ZN(new_n415));
  AOI211_X1 g229(.A(G131), .B(new_n342), .C1(new_n356), .C2(new_n357), .ZN(new_n416));
  OAI21_X1  g230(.A(new_n333), .B1(new_n415), .B2(new_n416), .ZN(new_n417));
  INV_X1    g231(.A(new_n226), .ZN(new_n418));
  INV_X1    g232(.A(new_n405), .ZN(new_n419));
  NAND3_X1  g233(.A1(new_n417), .A2(new_n418), .A3(new_n419), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n420), .A2(KEYINPUT69), .ZN(new_n421));
  INV_X1    g235(.A(KEYINPUT69), .ZN(new_n422));
  NAND4_X1  g236(.A1(new_n417), .A2(new_n419), .A3(new_n422), .A4(new_n418), .ZN(new_n423));
  AND2_X1   g237(.A1(new_n421), .A2(new_n423), .ZN(new_n424));
  XOR2_X1   g238(.A(KEYINPUT71), .B(KEYINPUT27), .Z(new_n425));
  XNOR2_X1  g239(.A(new_n425), .B(KEYINPUT72), .ZN(new_n426));
  INV_X1    g240(.A(G237), .ZN(new_n427));
  NAND3_X1  g241(.A1(new_n317), .A2(G210), .A3(new_n427), .ZN(new_n428));
  XNOR2_X1  g242(.A(new_n426), .B(new_n428), .ZN(new_n429));
  XNOR2_X1  g243(.A(KEYINPUT26), .B(G101), .ZN(new_n430));
  XNOR2_X1  g244(.A(new_n429), .B(new_n430), .ZN(new_n431));
  INV_X1    g245(.A(new_n431), .ZN(new_n432));
  NAND4_X1  g246(.A1(new_n413), .A2(new_n414), .A3(new_n424), .A4(new_n432), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n417), .A2(new_n419), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n434), .A2(new_n226), .ZN(new_n435));
  NAND3_X1  g249(.A1(new_n421), .A2(new_n435), .A3(new_n423), .ZN(new_n436));
  INV_X1    g250(.A(KEYINPUT74), .ZN(new_n437));
  NAND3_X1  g251(.A1(new_n436), .A2(new_n437), .A3(KEYINPUT28), .ZN(new_n438));
  INV_X1    g252(.A(new_n438), .ZN(new_n439));
  INV_X1    g253(.A(KEYINPUT28), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n420), .A2(new_n440), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n441), .A2(KEYINPUT74), .ZN(new_n442));
  AOI21_X1  g256(.A(new_n442), .B1(new_n436), .B2(KEYINPUT28), .ZN(new_n443));
  NOR3_X1   g257(.A1(new_n439), .A2(new_n414), .A3(new_n443), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n436), .A2(KEYINPUT28), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n445), .A2(new_n441), .ZN(new_n446));
  OAI21_X1  g260(.A(new_n431), .B1(new_n446), .B2(KEYINPUT29), .ZN(new_n447));
  OAI211_X1 g261(.A(new_n297), .B(new_n433), .C1(new_n444), .C2(new_n447), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n448), .A2(G472), .ZN(new_n449));
  INV_X1    g263(.A(KEYINPUT30), .ZN(new_n450));
  OAI21_X1  g264(.A(KEYINPUT68), .B1(new_n434), .B2(new_n450), .ZN(new_n451));
  AOI21_X1  g265(.A(new_n407), .B1(new_n410), .B2(new_n451), .ZN(new_n452));
  NAND3_X1  g266(.A1(new_n421), .A2(new_n431), .A3(new_n423), .ZN(new_n453));
  OAI21_X1  g267(.A(KEYINPUT31), .B1(new_n452), .B2(new_n453), .ZN(new_n454));
  INV_X1    g268(.A(KEYINPUT73), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n454), .A2(new_n455), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n446), .A2(new_n432), .ZN(new_n457));
  OR3_X1    g271(.A1(new_n452), .A2(KEYINPUT31), .A3(new_n453), .ZN(new_n458));
  OAI211_X1 g272(.A(KEYINPUT73), .B(KEYINPUT31), .C1(new_n452), .C2(new_n453), .ZN(new_n459));
  NAND4_X1  g273(.A1(new_n456), .A2(new_n457), .A3(new_n458), .A4(new_n459), .ZN(new_n460));
  INV_X1    g274(.A(KEYINPUT32), .ZN(new_n461));
  NOR2_X1   g275(.A1(G472), .A2(G902), .ZN(new_n462));
  AND3_X1   g276(.A1(new_n460), .A2(new_n461), .A3(new_n462), .ZN(new_n463));
  AOI21_X1  g277(.A(new_n461), .B1(new_n460), .B2(new_n462), .ZN(new_n464));
  OAI21_X1  g278(.A(new_n449), .B1(new_n463), .B2(new_n464), .ZN(new_n465));
  NAND3_X1  g279(.A1(new_n317), .A2(G221), .A3(G234), .ZN(new_n466));
  XNOR2_X1  g280(.A(KEYINPUT22), .B(G137), .ZN(new_n467));
  XOR2_X1   g281(.A(new_n466), .B(new_n467), .Z(new_n468));
  INV_X1    g282(.A(new_n468), .ZN(new_n469));
  XNOR2_X1  g283(.A(KEYINPUT24), .B(G110), .ZN(new_n470));
  XOR2_X1   g284(.A(new_n470), .B(KEYINPUT75), .Z(new_n471));
  NOR2_X1   g285(.A1(G119), .A2(G128), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n215), .A2(new_n216), .ZN(new_n473));
  AOI21_X1  g287(.A(new_n472), .B1(new_n473), .B2(G128), .ZN(new_n474));
  INV_X1    g288(.A(new_n474), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n471), .A2(new_n475), .ZN(new_n476));
  INV_X1    g290(.A(G140), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n477), .A2(G125), .ZN(new_n478));
  INV_X1    g292(.A(G125), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n479), .A2(G140), .ZN(new_n480));
  NAND3_X1  g294(.A1(new_n478), .A2(new_n480), .A3(KEYINPUT16), .ZN(new_n481));
  OR3_X1    g295(.A1(new_n479), .A2(KEYINPUT16), .A3(G140), .ZN(new_n482));
  NAND2_X1  g296(.A1(new_n481), .A2(new_n482), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n483), .A2(new_n190), .ZN(new_n484));
  NAND3_X1  g298(.A1(new_n481), .A2(new_n482), .A3(G146), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n484), .A2(new_n485), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n476), .A2(new_n486), .ZN(new_n487));
  INV_X1    g301(.A(G110), .ZN(new_n488));
  NAND2_X1  g302(.A1(new_n474), .A2(KEYINPUT23), .ZN(new_n489));
  AOI21_X1  g303(.A(G128), .B1(new_n215), .B2(new_n216), .ZN(new_n490));
  OR2_X1    g304(.A1(new_n490), .A2(KEYINPUT23), .ZN(new_n491));
  AOI21_X1  g305(.A(new_n488), .B1(new_n489), .B2(new_n491), .ZN(new_n492));
  OR3_X1    g306(.A1(new_n487), .A2(KEYINPUT76), .A3(new_n492), .ZN(new_n493));
  OAI21_X1  g307(.A(KEYINPUT76), .B1(new_n487), .B2(new_n492), .ZN(new_n494));
  NAND2_X1  g308(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  XNOR2_X1  g309(.A(G125), .B(G140), .ZN(new_n496));
  INV_X1    g310(.A(KEYINPUT77), .ZN(new_n497));
  OAI21_X1  g311(.A(new_n190), .B1(new_n496), .B2(new_n497), .ZN(new_n498));
  AND3_X1   g312(.A1(new_n478), .A2(new_n480), .A3(new_n497), .ZN(new_n499));
  OR2_X1    g313(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n500), .A2(new_n485), .ZN(new_n501));
  OR2_X1    g315(.A1(new_n471), .A2(new_n475), .ZN(new_n502));
  NAND3_X1  g316(.A1(new_n489), .A2(new_n488), .A3(new_n491), .ZN(new_n503));
  AOI21_X1  g317(.A(new_n501), .B1(new_n502), .B2(new_n503), .ZN(new_n504));
  INV_X1    g318(.A(new_n504), .ZN(new_n505));
  AOI21_X1  g319(.A(new_n469), .B1(new_n495), .B2(new_n505), .ZN(new_n506));
  AOI211_X1 g320(.A(new_n504), .B(new_n468), .C1(new_n493), .C2(new_n494), .ZN(new_n507));
  NOR2_X1   g321(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  INV_X1    g322(.A(new_n508), .ZN(new_n509));
  INV_X1    g323(.A(G217), .ZN(new_n510));
  AOI21_X1  g324(.A(new_n510), .B1(G234), .B2(new_n297), .ZN(new_n511));
  NOR2_X1   g325(.A1(new_n511), .A2(G902), .ZN(new_n512));
  INV_X1    g326(.A(new_n512), .ZN(new_n513));
  OR3_X1    g327(.A1(new_n509), .A2(KEYINPUT79), .A3(new_n513), .ZN(new_n514));
  OAI21_X1  g328(.A(KEYINPUT79), .B1(new_n509), .B2(new_n513), .ZN(new_n515));
  INV_X1    g329(.A(new_n511), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n495), .A2(new_n505), .ZN(new_n517));
  NAND2_X1  g331(.A1(new_n517), .A2(new_n468), .ZN(new_n518));
  NAND3_X1  g332(.A1(new_n495), .A2(new_n505), .A3(new_n469), .ZN(new_n519));
  INV_X1    g333(.A(KEYINPUT78), .ZN(new_n520));
  INV_X1    g334(.A(KEYINPUT25), .ZN(new_n521));
  AOI21_X1  g335(.A(G902), .B1(new_n520), .B2(new_n521), .ZN(new_n522));
  NAND3_X1  g336(.A1(new_n518), .A2(new_n519), .A3(new_n522), .ZN(new_n523));
  NOR2_X1   g337(.A1(new_n520), .A2(new_n521), .ZN(new_n524));
  AOI21_X1  g338(.A(new_n516), .B1(new_n523), .B2(new_n524), .ZN(new_n525));
  INV_X1    g339(.A(new_n525), .ZN(new_n526));
  INV_X1    g340(.A(new_n522), .ZN(new_n527));
  NOR3_X1   g341(.A1(new_n506), .A2(new_n507), .A3(new_n527), .ZN(new_n528));
  INV_X1    g342(.A(new_n524), .ZN(new_n529));
  NAND2_X1  g343(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  INV_X1    g344(.A(new_n530), .ZN(new_n531));
  OAI211_X1 g345(.A(new_n514), .B(new_n515), .C1(new_n526), .C2(new_n531), .ZN(new_n532));
  INV_X1    g346(.A(new_n532), .ZN(new_n533));
  INV_X1    g347(.A(G116), .ZN(new_n534));
  INV_X1    g348(.A(G122), .ZN(new_n535));
  OR2_X1    g349(.A1(new_n535), .A2(KEYINPUT106), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n535), .A2(KEYINPUT106), .ZN(new_n537));
  AOI21_X1  g351(.A(new_n534), .B1(new_n536), .B2(new_n537), .ZN(new_n538));
  NAND3_X1  g352(.A1(new_n218), .A2(G122), .A3(new_n219), .ZN(new_n539));
  AOI21_X1  g353(.A(new_n538), .B1(new_n539), .B2(KEYINPUT14), .ZN(new_n540));
  OAI21_X1  g354(.A(new_n540), .B1(KEYINPUT14), .B2(new_n539), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n541), .A2(G107), .ZN(new_n542));
  INV_X1    g356(.A(new_n539), .ZN(new_n543));
  NOR3_X1   g357(.A1(new_n538), .A2(new_n543), .A3(G107), .ZN(new_n544));
  INV_X1    g358(.A(new_n544), .ZN(new_n545));
  NAND2_X1  g359(.A1(new_n192), .A2(G128), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n202), .A2(G143), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n546), .A2(new_n547), .ZN(new_n548));
  XNOR2_X1  g362(.A(new_n548), .B(new_n341), .ZN(new_n549));
  NAND3_X1  g363(.A1(new_n542), .A2(new_n545), .A3(new_n549), .ZN(new_n550));
  NAND3_X1  g364(.A1(new_n192), .A2(KEYINPUT13), .A3(G128), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n551), .A2(new_n547), .ZN(new_n552));
  AOI21_X1  g366(.A(KEYINPUT13), .B1(new_n192), .B2(G128), .ZN(new_n553));
  OAI21_X1  g367(.A(G134), .B1(new_n552), .B2(new_n553), .ZN(new_n554));
  XNOR2_X1  g368(.A(new_n554), .B(KEYINPUT107), .ZN(new_n555));
  NOR2_X1   g369(.A1(new_n538), .A2(new_n543), .ZN(new_n556));
  NOR2_X1   g370(.A1(new_n556), .A2(new_n233), .ZN(new_n557));
  OAI221_X1 g371(.A(new_n555), .B1(new_n341), .B2(new_n548), .C1(new_n557), .C2(new_n544), .ZN(new_n558));
  NOR3_X1   g372(.A1(new_n397), .A2(new_n510), .A3(G953), .ZN(new_n559));
  NAND3_X1  g373(.A1(new_n550), .A2(new_n558), .A3(new_n559), .ZN(new_n560));
  INV_X1    g374(.A(new_n560), .ZN(new_n561));
  AOI21_X1  g375(.A(new_n559), .B1(new_n550), .B2(new_n558), .ZN(new_n562));
  OAI21_X1  g376(.A(new_n297), .B1(new_n561), .B2(new_n562), .ZN(new_n563));
  INV_X1    g377(.A(G478), .ZN(new_n564));
  NOR2_X1   g378(.A1(new_n564), .A2(KEYINPUT15), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n563), .A2(new_n565), .ZN(new_n566));
  OAI221_X1 g380(.A(new_n297), .B1(KEYINPUT15), .B2(new_n564), .C1(new_n561), .C2(new_n562), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  INV_X1    g382(.A(G952), .ZN(new_n569));
  NOR2_X1   g383(.A1(new_n569), .A2(G953), .ZN(new_n570));
  NAND2_X1  g384(.A1(G234), .A2(G237), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n570), .A2(new_n571), .ZN(new_n572));
  XNOR2_X1  g386(.A(new_n572), .B(KEYINPUT108), .ZN(new_n573));
  INV_X1    g387(.A(new_n573), .ZN(new_n574));
  INV_X1    g388(.A(new_n317), .ZN(new_n575));
  NAND3_X1  g389(.A1(new_n575), .A2(G902), .A3(new_n571), .ZN(new_n576));
  INV_X1    g390(.A(new_n576), .ZN(new_n577));
  XNOR2_X1  g391(.A(KEYINPUT21), .B(G898), .ZN(new_n578));
  AOI21_X1  g392(.A(new_n574), .B1(new_n577), .B2(new_n578), .ZN(new_n579));
  NOR2_X1   g393(.A1(new_n568), .A2(new_n579), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n207), .A2(KEYINPUT70), .ZN(new_n581));
  INV_X1    g395(.A(KEYINPUT70), .ZN(new_n582));
  NAND2_X1  g396(.A1(new_n582), .A2(G953), .ZN(new_n583));
  NAND4_X1  g397(.A1(new_n581), .A2(new_n583), .A3(G214), .A4(new_n427), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n584), .A2(new_n192), .ZN(new_n585));
  NAND4_X1  g399(.A1(new_n317), .A2(G143), .A3(G214), .A4(new_n427), .ZN(new_n586));
  NAND2_X1  g400(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  INV_X1    g401(.A(KEYINPUT18), .ZN(new_n588));
  NOR2_X1   g402(.A1(new_n588), .A2(KEYINPUT98), .ZN(new_n589));
  NAND3_X1  g403(.A1(new_n587), .A2(G131), .A3(new_n589), .ZN(new_n590));
  OAI22_X1  g404(.A1(new_n498), .A2(new_n499), .B1(new_n190), .B2(new_n496), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n589), .A2(G131), .ZN(new_n592));
  NAND3_X1  g406(.A1(new_n585), .A2(new_n586), .A3(new_n592), .ZN(new_n593));
  NAND3_X1  g407(.A1(new_n590), .A2(new_n591), .A3(new_n593), .ZN(new_n594));
  XNOR2_X1  g408(.A(G113), .B(G122), .ZN(new_n595));
  XNOR2_X1  g409(.A(KEYINPUT100), .B(G104), .ZN(new_n596));
  XNOR2_X1  g410(.A(new_n595), .B(new_n596), .ZN(new_n597));
  AND3_X1   g411(.A1(new_n585), .A2(new_n586), .A3(new_n359), .ZN(new_n598));
  AOI21_X1  g412(.A(new_n359), .B1(new_n585), .B2(new_n586), .ZN(new_n599));
  NOR3_X1   g413(.A1(new_n598), .A2(new_n599), .A3(KEYINPUT17), .ZN(new_n600));
  NAND3_X1  g414(.A1(new_n587), .A2(KEYINPUT17), .A3(G131), .ZN(new_n601));
  INV_X1    g415(.A(new_n485), .ZN(new_n602));
  AOI21_X1  g416(.A(G146), .B1(new_n481), .B2(new_n482), .ZN(new_n603));
  NOR2_X1   g417(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  NAND2_X1  g418(.A1(new_n601), .A2(new_n604), .ZN(new_n605));
  OAI211_X1 g419(.A(new_n594), .B(new_n597), .C1(new_n600), .C2(new_n605), .ZN(new_n606));
  NAND2_X1  g420(.A1(new_n606), .A2(KEYINPUT101), .ZN(new_n607));
  AOI21_X1  g421(.A(new_n486), .B1(KEYINPUT17), .B2(new_n599), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n587), .A2(G131), .ZN(new_n609));
  INV_X1    g423(.A(KEYINPUT17), .ZN(new_n610));
  NAND3_X1  g424(.A1(new_n585), .A2(new_n586), .A3(new_n359), .ZN(new_n611));
  NAND3_X1  g425(.A1(new_n609), .A2(new_n610), .A3(new_n611), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n608), .A2(new_n612), .ZN(new_n613));
  INV_X1    g427(.A(KEYINPUT101), .ZN(new_n614));
  NAND4_X1  g428(.A1(new_n613), .A2(new_n614), .A3(new_n594), .A4(new_n597), .ZN(new_n615));
  AND2_X1   g429(.A1(new_n607), .A2(new_n615), .ZN(new_n616));
  INV_X1    g430(.A(KEYINPUT104), .ZN(new_n617));
  AND2_X1   g431(.A1(new_n591), .A2(new_n593), .ZN(new_n618));
  AOI22_X1  g432(.A1(new_n608), .A2(new_n612), .B1(new_n618), .B2(new_n590), .ZN(new_n619));
  OAI21_X1  g433(.A(new_n617), .B1(new_n619), .B2(new_n597), .ZN(new_n620));
  OAI21_X1  g434(.A(new_n594), .B1(new_n600), .B2(new_n605), .ZN(new_n621));
  INV_X1    g435(.A(new_n597), .ZN(new_n622));
  NAND3_X1  g436(.A1(new_n621), .A2(KEYINPUT104), .A3(new_n622), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n620), .A2(new_n623), .ZN(new_n624));
  OAI21_X1  g438(.A(new_n297), .B1(new_n616), .B2(new_n624), .ZN(new_n625));
  INV_X1    g439(.A(KEYINPUT105), .ZN(new_n626));
  NAND2_X1  g440(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  OAI211_X1 g441(.A(KEYINPUT105), .B(new_n297), .C1(new_n616), .C2(new_n624), .ZN(new_n628));
  NAND3_X1  g442(.A1(new_n627), .A2(G475), .A3(new_n628), .ZN(new_n629));
  INV_X1    g443(.A(KEYINPUT103), .ZN(new_n630));
  INV_X1    g444(.A(G475), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n631), .A2(new_n297), .ZN(new_n632));
  INV_X1    g446(.A(KEYINPUT102), .ZN(new_n633));
  NAND2_X1  g447(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  INV_X1    g448(.A(KEYINPUT20), .ZN(new_n635));
  NAND3_X1  g449(.A1(new_n631), .A2(new_n297), .A3(KEYINPUT102), .ZN(new_n636));
  NAND3_X1  g450(.A1(new_n634), .A2(new_n635), .A3(new_n636), .ZN(new_n637));
  INV_X1    g451(.A(new_n637), .ZN(new_n638));
  OAI21_X1  g452(.A(KEYINPUT99), .B1(new_n496), .B2(new_n497), .ZN(new_n639));
  INV_X1    g453(.A(KEYINPUT19), .ZN(new_n640));
  INV_X1    g454(.A(KEYINPUT99), .ZN(new_n641));
  OAI21_X1  g455(.A(KEYINPUT77), .B1(new_n641), .B2(new_n640), .ZN(new_n642));
  AOI22_X1  g456(.A1(new_n639), .A2(new_n640), .B1(new_n496), .B2(new_n642), .ZN(new_n643));
  OAI221_X1 g457(.A(new_n485), .B1(new_n643), .B2(G146), .C1(new_n598), .C2(new_n599), .ZN(new_n644));
  AOI21_X1  g458(.A(new_n597), .B1(new_n644), .B2(new_n594), .ZN(new_n645));
  OAI211_X1 g459(.A(new_n630), .B(new_n638), .C1(new_n616), .C2(new_n645), .ZN(new_n646));
  AOI21_X1  g460(.A(new_n645), .B1(new_n607), .B2(new_n615), .ZN(new_n647));
  OAI21_X1  g461(.A(KEYINPUT103), .B1(new_n647), .B2(new_n637), .ZN(new_n648));
  OAI21_X1  g462(.A(KEYINPUT20), .B1(new_n647), .B2(new_n632), .ZN(new_n649));
  NAND3_X1  g463(.A1(new_n646), .A2(new_n648), .A3(new_n649), .ZN(new_n650));
  NAND3_X1  g464(.A1(new_n580), .A2(new_n629), .A3(new_n650), .ZN(new_n651));
  INV_X1    g465(.A(new_n651), .ZN(new_n652));
  AND4_X1   g466(.A1(new_n400), .A2(new_n465), .A3(new_n533), .A4(new_n652), .ZN(new_n653));
  XNOR2_X1  g467(.A(new_n653), .B(new_n243), .ZN(G3));
  NAND2_X1  g468(.A1(new_n460), .A2(new_n297), .ZN(new_n655));
  AOI22_X1  g469(.A1(new_n655), .A2(G472), .B1(new_n462), .B2(new_n460), .ZN(new_n656));
  NOR2_X1   g470(.A1(new_n532), .A2(new_n399), .ZN(new_n657));
  NAND2_X1  g471(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  INV_X1    g472(.A(new_n658), .ZN(new_n659));
  NAND2_X1  g473(.A1(new_n309), .A2(new_n310), .ZN(new_n660));
  NAND2_X1  g474(.A1(new_n628), .A2(G475), .ZN(new_n661));
  AOI21_X1  g475(.A(new_n614), .B1(new_n619), .B2(new_n597), .ZN(new_n662));
  NOR2_X1   g476(.A1(new_n606), .A2(KEYINPUT101), .ZN(new_n663));
  OAI211_X1 g477(.A(new_n620), .B(new_n623), .C1(new_n662), .C2(new_n663), .ZN(new_n664));
  AOI21_X1  g478(.A(KEYINPUT105), .B1(new_n664), .B2(new_n297), .ZN(new_n665));
  OAI21_X1  g479(.A(new_n650), .B1(new_n661), .B2(new_n665), .ZN(new_n666));
  INV_X1    g480(.A(new_n562), .ZN(new_n667));
  INV_X1    g481(.A(KEYINPUT33), .ZN(new_n668));
  NAND3_X1  g482(.A1(new_n667), .A2(new_n668), .A3(new_n560), .ZN(new_n669));
  OAI21_X1  g483(.A(KEYINPUT33), .B1(new_n561), .B2(new_n562), .ZN(new_n670));
  NAND3_X1  g484(.A1(new_n669), .A2(new_n670), .A3(G478), .ZN(new_n671));
  OAI211_X1 g485(.A(new_n564), .B(new_n297), .C1(new_n561), .C2(new_n562), .ZN(new_n672));
  NAND2_X1  g486(.A1(G478), .A2(G902), .ZN(new_n673));
  NAND3_X1  g487(.A1(new_n671), .A2(new_n672), .A3(new_n673), .ZN(new_n674));
  INV_X1    g488(.A(new_n674), .ZN(new_n675));
  NAND2_X1  g489(.A1(new_n666), .A2(new_n675), .ZN(new_n676));
  NOR3_X1   g490(.A1(new_n660), .A2(new_n579), .A3(new_n676), .ZN(new_n677));
  NAND2_X1  g491(.A1(new_n659), .A2(new_n677), .ZN(new_n678));
  XOR2_X1   g492(.A(KEYINPUT34), .B(G104), .Z(new_n679));
  XNOR2_X1  g493(.A(new_n678), .B(new_n679), .ZN(G6));
  NOR2_X1   g494(.A1(new_n647), .A2(new_n632), .ZN(new_n681));
  NAND2_X1  g495(.A1(new_n681), .A2(new_n635), .ZN(new_n682));
  NAND2_X1  g496(.A1(new_n682), .A2(new_n649), .ZN(new_n683));
  NAND3_X1  g497(.A1(new_n629), .A2(new_n683), .A3(new_n568), .ZN(new_n684));
  NOR3_X1   g498(.A1(new_n660), .A2(new_n579), .A3(new_n684), .ZN(new_n685));
  NAND2_X1  g499(.A1(new_n659), .A2(new_n685), .ZN(new_n686));
  XOR2_X1   g500(.A(KEYINPUT35), .B(G107), .Z(new_n687));
  XNOR2_X1  g501(.A(new_n686), .B(new_n687), .ZN(G9));
  NOR2_X1   g502(.A1(new_n468), .A2(KEYINPUT36), .ZN(new_n689));
  XNOR2_X1  g503(.A(new_n517), .B(new_n689), .ZN(new_n690));
  AOI22_X1  g504(.A1(new_n525), .A2(new_n530), .B1(new_n512), .B2(new_n690), .ZN(new_n691));
  NOR2_X1   g505(.A1(new_n691), .A2(new_n651), .ZN(new_n692));
  NAND3_X1  g506(.A1(new_n400), .A2(new_n656), .A3(new_n692), .ZN(new_n693));
  XOR2_X1   g507(.A(KEYINPUT37), .B(G110), .Z(new_n694));
  XNOR2_X1  g508(.A(new_n693), .B(new_n694), .ZN(G12));
  NOR3_X1   g509(.A1(new_n660), .A2(new_n399), .A3(new_n691), .ZN(new_n696));
  AND2_X1   g510(.A1(new_n465), .A2(new_n696), .ZN(new_n697));
  INV_X1    g511(.A(new_n629), .ZN(new_n698));
  XOR2_X1   g512(.A(new_n573), .B(KEYINPUT109), .Z(new_n699));
  INV_X1    g513(.A(new_n699), .ZN(new_n700));
  INV_X1    g514(.A(G900), .ZN(new_n701));
  AOI21_X1  g515(.A(new_n700), .B1(new_n701), .B2(new_n577), .ZN(new_n702));
  INV_X1    g516(.A(new_n702), .ZN(new_n703));
  NAND2_X1  g517(.A1(new_n683), .A2(new_n703), .ZN(new_n704));
  INV_X1    g518(.A(new_n568), .ZN(new_n705));
  NOR3_X1   g519(.A1(new_n698), .A2(new_n704), .A3(new_n705), .ZN(new_n706));
  NAND2_X1  g520(.A1(new_n697), .A2(new_n706), .ZN(new_n707));
  XNOR2_X1  g521(.A(new_n707), .B(G128), .ZN(G30));
  INV_X1    g522(.A(new_n399), .ZN(new_n709));
  XNOR2_X1  g523(.A(KEYINPUT111), .B(KEYINPUT39), .ZN(new_n710));
  XOR2_X1   g524(.A(new_n702), .B(new_n710), .Z(new_n711));
  INV_X1    g525(.A(new_n711), .ZN(new_n712));
  NAND2_X1  g526(.A1(new_n709), .A2(new_n712), .ZN(new_n713));
  NAND2_X1  g527(.A1(new_n713), .A2(KEYINPUT40), .ZN(new_n714));
  INV_X1    g528(.A(KEYINPUT38), .ZN(new_n715));
  NAND2_X1  g529(.A1(new_n309), .A2(new_n715), .ZN(new_n716));
  NAND3_X1  g530(.A1(new_n299), .A2(new_n308), .A3(KEYINPUT38), .ZN(new_n717));
  AND2_X1   g531(.A1(new_n716), .A2(new_n717), .ZN(new_n718));
  NAND2_X1  g532(.A1(new_n714), .A2(new_n718), .ZN(new_n719));
  NOR2_X1   g533(.A1(new_n713), .A2(KEYINPUT40), .ZN(new_n720));
  AOI21_X1  g534(.A(new_n705), .B1(new_n629), .B2(new_n650), .ZN(new_n721));
  NAND2_X1  g535(.A1(new_n721), .A2(new_n310), .ZN(new_n722));
  NOR3_X1   g536(.A1(new_n719), .A2(new_n720), .A3(new_n722), .ZN(new_n723));
  AOI21_X1  g537(.A(new_n432), .B1(new_n413), .B2(new_n424), .ZN(new_n724));
  OAI21_X1  g538(.A(new_n297), .B1(new_n436), .B2(new_n431), .ZN(new_n725));
  OAI21_X1  g539(.A(G472), .B1(new_n724), .B2(new_n725), .ZN(new_n726));
  XNOR2_X1  g540(.A(new_n726), .B(KEYINPUT110), .ZN(new_n727));
  OAI21_X1  g541(.A(new_n727), .B1(new_n463), .B2(new_n464), .ZN(new_n728));
  NAND3_X1  g542(.A1(new_n723), .A2(new_n691), .A3(new_n728), .ZN(new_n729));
  XNOR2_X1  g543(.A(new_n729), .B(G143), .ZN(G45));
  NOR2_X1   g544(.A1(new_n676), .A2(new_n702), .ZN(new_n731));
  NAND2_X1  g545(.A1(new_n697), .A2(new_n731), .ZN(new_n732));
  XNOR2_X1  g546(.A(KEYINPUT112), .B(G146), .ZN(new_n733));
  XNOR2_X1  g547(.A(new_n732), .B(new_n733), .ZN(G48));
  NAND2_X1  g548(.A1(new_n384), .A2(new_n385), .ZN(new_n735));
  AOI22_X1  g549(.A1(new_n735), .A2(new_n319), .B1(new_n377), .B2(new_n363), .ZN(new_n736));
  OAI21_X1  g550(.A(G469), .B1(new_n736), .B2(G902), .ZN(new_n737));
  NAND3_X1  g551(.A1(new_n737), .A2(new_n398), .A3(new_n387), .ZN(new_n738));
  INV_X1    g552(.A(new_n738), .ZN(new_n739));
  NAND4_X1  g553(.A1(new_n465), .A2(new_n533), .A3(new_n677), .A4(new_n739), .ZN(new_n740));
  XNOR2_X1  g554(.A(KEYINPUT41), .B(G113), .ZN(new_n741));
  XNOR2_X1  g555(.A(new_n740), .B(new_n741), .ZN(G15));
  NAND4_X1  g556(.A1(new_n465), .A2(new_n685), .A3(new_n533), .A4(new_n739), .ZN(new_n743));
  XNOR2_X1  g557(.A(new_n743), .B(G116), .ZN(G18));
  NOR4_X1   g558(.A1(new_n660), .A2(new_n651), .A3(new_n691), .A4(new_n738), .ZN(new_n745));
  NAND2_X1  g559(.A1(new_n745), .A2(new_n465), .ZN(new_n746));
  NAND2_X1  g560(.A1(new_n746), .A2(KEYINPUT113), .ZN(new_n747));
  INV_X1    g561(.A(KEYINPUT113), .ZN(new_n748));
  NAND3_X1  g562(.A1(new_n745), .A2(new_n465), .A3(new_n748), .ZN(new_n749));
  NAND2_X1  g563(.A1(new_n747), .A2(new_n749), .ZN(new_n750));
  XNOR2_X1  g564(.A(new_n750), .B(G119), .ZN(G21));
  INV_X1    g565(.A(new_n462), .ZN(new_n752));
  OAI21_X1  g566(.A(KEYINPUT114), .B1(new_n439), .B2(new_n443), .ZN(new_n753));
  INV_X1    g567(.A(new_n443), .ZN(new_n754));
  INV_X1    g568(.A(KEYINPUT114), .ZN(new_n755));
  NAND3_X1  g569(.A1(new_n754), .A2(new_n755), .A3(new_n438), .ZN(new_n756));
  NAND3_X1  g570(.A1(new_n753), .A2(new_n756), .A3(new_n432), .ZN(new_n757));
  AND2_X1   g571(.A1(new_n458), .A2(new_n454), .ZN(new_n758));
  AOI21_X1  g572(.A(new_n752), .B1(new_n757), .B2(new_n758), .ZN(new_n759));
  INV_X1    g573(.A(G472), .ZN(new_n760));
  AOI21_X1  g574(.A(new_n760), .B1(new_n460), .B2(new_n297), .ZN(new_n761));
  NOR3_X1   g575(.A1(new_n759), .A2(new_n761), .A3(new_n532), .ZN(new_n762));
  NAND3_X1  g576(.A1(new_n721), .A2(new_n309), .A3(new_n310), .ZN(new_n763));
  NOR3_X1   g577(.A1(new_n763), .A2(new_n579), .A3(new_n738), .ZN(new_n764));
  NAND2_X1  g578(.A1(new_n762), .A2(new_n764), .ZN(new_n765));
  XNOR2_X1  g579(.A(new_n765), .B(G122), .ZN(G24));
  NOR3_X1   g580(.A1(new_n759), .A2(new_n761), .A3(new_n691), .ZN(new_n767));
  NOR2_X1   g581(.A1(new_n660), .A2(new_n738), .ZN(new_n768));
  AOI21_X1  g582(.A(new_n674), .B1(new_n629), .B2(new_n650), .ZN(new_n769));
  AOI21_X1  g583(.A(KEYINPUT115), .B1(new_n769), .B2(new_n703), .ZN(new_n770));
  AND4_X1   g584(.A1(KEYINPUT115), .A2(new_n666), .A3(new_n675), .A4(new_n703), .ZN(new_n771));
  NOR2_X1   g585(.A1(new_n770), .A2(new_n771), .ZN(new_n772));
  NAND3_X1  g586(.A1(new_n767), .A2(new_n768), .A3(new_n772), .ZN(new_n773));
  XNOR2_X1  g587(.A(new_n773), .B(G125), .ZN(G27));
  NAND2_X1  g588(.A1(new_n394), .A2(new_n389), .ZN(new_n775));
  AND3_X1   g589(.A1(new_n381), .A2(new_n362), .A3(new_n382), .ZN(new_n776));
  AOI21_X1  g590(.A(new_n362), .B1(new_n381), .B2(new_n382), .ZN(new_n777));
  OAI21_X1  g591(.A(new_n319), .B1(new_n776), .B2(new_n777), .ZN(new_n778));
  AOI211_X1 g592(.A(G469), .B(G902), .C1(new_n778), .C2(new_n378), .ZN(new_n779));
  OAI21_X1  g593(.A(KEYINPUT116), .B1(new_n775), .B2(new_n779), .ZN(new_n780));
  INV_X1    g594(.A(KEYINPUT116), .ZN(new_n781));
  NAND4_X1  g595(.A1(new_n387), .A2(new_n781), .A3(new_n389), .A4(new_n394), .ZN(new_n782));
  NAND3_X1  g596(.A1(new_n780), .A2(new_n398), .A3(new_n782), .ZN(new_n783));
  NAND3_X1  g597(.A1(new_n299), .A2(new_n308), .A3(new_n310), .ZN(new_n784));
  NOR2_X1   g598(.A1(new_n783), .A2(new_n784), .ZN(new_n785));
  NAND4_X1  g599(.A1(new_n465), .A2(new_n772), .A3(new_n533), .A4(new_n785), .ZN(new_n786));
  INV_X1    g600(.A(KEYINPUT42), .ZN(new_n787));
  NAND2_X1  g601(.A1(new_n786), .A2(new_n787), .ZN(new_n788));
  INV_X1    g602(.A(KEYINPUT115), .ZN(new_n789));
  OAI21_X1  g603(.A(new_n789), .B1(new_n676), .B2(new_n702), .ZN(new_n790));
  NAND3_X1  g604(.A1(new_n769), .A2(KEYINPUT115), .A3(new_n703), .ZN(new_n791));
  NAND2_X1  g605(.A1(new_n790), .A2(new_n791), .ZN(new_n792));
  AND3_X1   g606(.A1(new_n299), .A2(new_n308), .A3(new_n310), .ZN(new_n793));
  NAND4_X1  g607(.A1(new_n793), .A2(new_n398), .A3(new_n782), .A4(new_n780), .ZN(new_n794));
  NOR2_X1   g608(.A1(new_n792), .A2(new_n794), .ZN(new_n795));
  NAND4_X1  g609(.A1(new_n795), .A2(KEYINPUT42), .A3(new_n465), .A4(new_n533), .ZN(new_n796));
  NAND2_X1  g610(.A1(new_n788), .A2(new_n796), .ZN(new_n797));
  XNOR2_X1  g611(.A(new_n797), .B(G131), .ZN(G33));
  NAND4_X1  g612(.A1(new_n465), .A2(new_n533), .A3(new_n706), .A4(new_n785), .ZN(new_n799));
  XNOR2_X1  g613(.A(new_n799), .B(G134), .ZN(G36));
  OAI21_X1  g614(.A(new_n390), .B1(new_n392), .B2(new_n393), .ZN(new_n801));
  INV_X1    g615(.A(KEYINPUT45), .ZN(new_n802));
  NAND2_X1  g616(.A1(new_n801), .A2(new_n802), .ZN(new_n803));
  OAI211_X1 g617(.A(KEYINPUT45), .B(new_n390), .C1(new_n392), .C2(new_n393), .ZN(new_n804));
  NAND3_X1  g618(.A1(new_n803), .A2(G469), .A3(new_n804), .ZN(new_n805));
  AOI21_X1  g619(.A(KEYINPUT46), .B1(new_n805), .B2(new_n389), .ZN(new_n806));
  OR2_X1    g620(.A1(new_n806), .A2(new_n779), .ZN(new_n807));
  AND3_X1   g621(.A1(new_n805), .A2(KEYINPUT46), .A3(new_n389), .ZN(new_n808));
  OAI211_X1 g622(.A(new_n398), .B(new_n712), .C1(new_n807), .C2(new_n808), .ZN(new_n809));
  OR2_X1    g623(.A1(new_n656), .A2(new_n691), .ZN(new_n810));
  INV_X1    g624(.A(new_n666), .ZN(new_n811));
  NAND2_X1  g625(.A1(new_n811), .A2(new_n675), .ZN(new_n812));
  NAND2_X1  g626(.A1(new_n812), .A2(KEYINPUT43), .ZN(new_n813));
  OR3_X1    g627(.A1(new_n666), .A2(KEYINPUT43), .A3(new_n674), .ZN(new_n814));
  NAND2_X1  g628(.A1(new_n813), .A2(new_n814), .ZN(new_n815));
  OR2_X1    g629(.A1(new_n810), .A2(new_n815), .ZN(new_n816));
  INV_X1    g630(.A(KEYINPUT44), .ZN(new_n817));
  AOI21_X1  g631(.A(new_n809), .B1(new_n816), .B2(new_n817), .ZN(new_n818));
  OR3_X1    g632(.A1(new_n810), .A2(new_n817), .A3(new_n815), .ZN(new_n819));
  NAND3_X1  g633(.A1(new_n818), .A2(new_n793), .A3(new_n819), .ZN(new_n820));
  XNOR2_X1  g634(.A(KEYINPUT117), .B(G137), .ZN(new_n821));
  XNOR2_X1  g635(.A(new_n820), .B(new_n821), .ZN(G39));
  INV_X1    g636(.A(KEYINPUT47), .ZN(new_n823));
  NOR3_X1   g637(.A1(new_n808), .A2(new_n806), .A3(new_n779), .ZN(new_n824));
  INV_X1    g638(.A(new_n398), .ZN(new_n825));
  OAI21_X1  g639(.A(new_n823), .B1(new_n824), .B2(new_n825), .ZN(new_n826));
  OAI211_X1 g640(.A(KEYINPUT47), .B(new_n398), .C1(new_n807), .C2(new_n808), .ZN(new_n827));
  NAND2_X1  g641(.A1(new_n826), .A2(new_n827), .ZN(new_n828));
  NAND2_X1  g642(.A1(new_n460), .A2(new_n462), .ZN(new_n829));
  NAND2_X1  g643(.A1(new_n829), .A2(KEYINPUT32), .ZN(new_n830));
  NAND3_X1  g644(.A1(new_n460), .A2(new_n461), .A3(new_n462), .ZN(new_n831));
  AOI22_X1  g645(.A1(new_n830), .A2(new_n831), .B1(G472), .B2(new_n448), .ZN(new_n832));
  AND3_X1   g646(.A1(new_n731), .A2(new_n532), .A3(new_n793), .ZN(new_n833));
  NAND3_X1  g647(.A1(new_n828), .A2(new_n832), .A3(new_n833), .ZN(new_n834));
  XNOR2_X1  g648(.A(new_n834), .B(G140), .ZN(G42));
  NOR3_X1   g649(.A1(new_n532), .A2(new_n825), .A3(new_n312), .ZN(new_n836));
  NAND2_X1  g650(.A1(new_n737), .A2(new_n387), .ZN(new_n837));
  OR2_X1    g651(.A1(new_n837), .A2(KEYINPUT49), .ZN(new_n838));
  NAND2_X1  g652(.A1(new_n837), .A2(KEYINPUT49), .ZN(new_n839));
  NAND3_X1  g653(.A1(new_n836), .A2(new_n838), .A3(new_n839), .ZN(new_n840));
  OR4_X1    g654(.A1(new_n728), .A2(new_n840), .A3(new_n718), .A4(new_n812), .ZN(new_n841));
  AND3_X1   g655(.A1(new_n813), .A2(new_n700), .A3(new_n814), .ZN(new_n842));
  AOI211_X1 g656(.A(new_n310), .B(new_n738), .C1(new_n716), .C2(new_n717), .ZN(new_n843));
  NAND3_X1  g657(.A1(new_n842), .A2(new_n762), .A3(new_n843), .ZN(new_n844));
  INV_X1    g658(.A(KEYINPUT119), .ZN(new_n845));
  INV_X1    g659(.A(KEYINPUT50), .ZN(new_n846));
  NAND3_X1  g660(.A1(new_n844), .A2(new_n845), .A3(new_n846), .ZN(new_n847));
  NAND2_X1  g661(.A1(new_n845), .A2(new_n846), .ZN(new_n848));
  NAND4_X1  g662(.A1(new_n842), .A2(new_n762), .A3(new_n848), .A4(new_n843), .ZN(new_n849));
  NAND2_X1  g663(.A1(new_n847), .A2(new_n849), .ZN(new_n850));
  AND3_X1   g664(.A1(new_n842), .A2(new_n762), .A3(new_n793), .ZN(new_n851));
  NOR2_X1   g665(.A1(new_n837), .A2(new_n398), .ZN(new_n852));
  OAI21_X1  g666(.A(new_n851), .B1(new_n828), .B2(new_n852), .ZN(new_n853));
  NAND2_X1  g667(.A1(new_n793), .A2(new_n739), .ZN(new_n854));
  NOR3_X1   g668(.A1(new_n815), .A2(new_n699), .A3(new_n854), .ZN(new_n855));
  NAND2_X1  g669(.A1(new_n855), .A2(new_n767), .ZN(new_n856));
  INV_X1    g670(.A(new_n728), .ZN(new_n857));
  NOR3_X1   g671(.A1(new_n854), .A2(new_n532), .A3(new_n573), .ZN(new_n858));
  NAND4_X1  g672(.A1(new_n857), .A2(new_n811), .A3(new_n858), .A4(new_n674), .ZN(new_n859));
  AND2_X1   g673(.A1(new_n856), .A2(new_n859), .ZN(new_n860));
  NAND3_X1  g674(.A1(new_n850), .A2(new_n853), .A3(new_n860), .ZN(new_n861));
  INV_X1    g675(.A(KEYINPUT51), .ZN(new_n862));
  OR2_X1    g676(.A1(new_n861), .A2(new_n862), .ZN(new_n863));
  NAND3_X1  g677(.A1(new_n857), .A2(new_n769), .A3(new_n858), .ZN(new_n864));
  NAND3_X1  g678(.A1(new_n842), .A2(new_n768), .A3(new_n762), .ZN(new_n865));
  NAND3_X1  g679(.A1(new_n864), .A2(new_n865), .A3(new_n570), .ZN(new_n866));
  OR2_X1    g680(.A1(new_n866), .A2(KEYINPUT120), .ZN(new_n867));
  NAND2_X1  g681(.A1(new_n866), .A2(KEYINPUT120), .ZN(new_n868));
  AOI22_X1  g682(.A1(new_n861), .A2(new_n862), .B1(new_n867), .B2(new_n868), .ZN(new_n869));
  NOR2_X1   g683(.A1(new_n832), .A2(new_n532), .ZN(new_n870));
  NAND2_X1  g684(.A1(new_n870), .A2(new_n855), .ZN(new_n871));
  NAND2_X1  g685(.A1(new_n871), .A2(KEYINPUT121), .ZN(new_n872));
  INV_X1    g686(.A(KEYINPUT121), .ZN(new_n873));
  NAND3_X1  g687(.A1(new_n870), .A2(new_n855), .A3(new_n873), .ZN(new_n874));
  AOI21_X1  g688(.A(KEYINPUT122), .B1(new_n872), .B2(new_n874), .ZN(new_n875));
  NAND3_X1  g689(.A1(new_n872), .A2(KEYINPUT122), .A3(new_n874), .ZN(new_n876));
  AOI21_X1  g690(.A(new_n875), .B1(KEYINPUT48), .B2(new_n876), .ZN(new_n877));
  AND3_X1   g691(.A1(new_n875), .A2(KEYINPUT48), .A3(new_n876), .ZN(new_n878));
  OAI211_X1 g692(.A(new_n863), .B(new_n869), .C1(new_n877), .C2(new_n878), .ZN(new_n879));
  INV_X1    g693(.A(KEYINPUT54), .ZN(new_n880));
  NAND2_X1  g694(.A1(new_n660), .A2(KEYINPUT97), .ZN(new_n881));
  NAND3_X1  g695(.A1(new_n309), .A2(new_n187), .A3(new_n310), .ZN(new_n882));
  NAND3_X1  g696(.A1(new_n629), .A2(new_n650), .A3(new_n568), .ZN(new_n883));
  AOI21_X1  g697(.A(new_n579), .B1(new_n676), .B2(new_n883), .ZN(new_n884));
  NAND3_X1  g698(.A1(new_n881), .A2(new_n882), .A3(new_n884), .ZN(new_n885));
  NAND3_X1  g699(.A1(new_n881), .A2(new_n709), .A3(new_n882), .ZN(new_n886));
  NAND2_X1  g700(.A1(new_n655), .A2(G472), .ZN(new_n887));
  NAND3_X1  g701(.A1(new_n887), .A2(new_n829), .A3(new_n692), .ZN(new_n888));
  OAI22_X1  g702(.A1(new_n658), .A2(new_n885), .B1(new_n886), .B2(new_n888), .ZN(new_n889));
  NOR2_X1   g703(.A1(new_n653), .A2(new_n889), .ZN(new_n890));
  NOR2_X1   g704(.A1(new_n399), .A2(new_n691), .ZN(new_n891));
  NOR3_X1   g705(.A1(new_n698), .A2(new_n704), .A3(new_n568), .ZN(new_n892));
  NAND4_X1  g706(.A1(new_n465), .A2(new_n891), .A3(new_n793), .A4(new_n892), .ZN(new_n893));
  NAND2_X1  g707(.A1(new_n893), .A2(new_n799), .ZN(new_n894));
  INV_X1    g708(.A(new_n894), .ZN(new_n895));
  INV_X1    g709(.A(KEYINPUT118), .ZN(new_n896));
  NAND3_X1  g710(.A1(new_n795), .A2(new_n896), .A3(new_n767), .ZN(new_n897));
  INV_X1    g711(.A(new_n783), .ZN(new_n898));
  NAND4_X1  g712(.A1(new_n898), .A2(new_n790), .A3(new_n791), .A4(new_n793), .ZN(new_n899));
  INV_X1    g713(.A(new_n691), .ZN(new_n900));
  AND2_X1   g714(.A1(new_n757), .A2(new_n758), .ZN(new_n901));
  OAI211_X1 g715(.A(new_n887), .B(new_n900), .C1(new_n901), .C2(new_n752), .ZN(new_n902));
  OAI21_X1  g716(.A(KEYINPUT118), .B1(new_n899), .B2(new_n902), .ZN(new_n903));
  NAND2_X1  g717(.A1(new_n897), .A2(new_n903), .ZN(new_n904));
  NAND4_X1  g718(.A1(new_n890), .A2(new_n797), .A3(new_n895), .A4(new_n904), .ZN(new_n905));
  OAI211_X1 g719(.A(new_n465), .B(new_n696), .C1(new_n706), .C2(new_n731), .ZN(new_n906));
  NOR3_X1   g720(.A1(new_n763), .A2(new_n783), .A3(new_n702), .ZN(new_n907));
  NAND3_X1  g721(.A1(new_n907), .A2(new_n691), .A3(new_n728), .ZN(new_n908));
  INV_X1    g722(.A(KEYINPUT52), .ZN(new_n909));
  NAND4_X1  g723(.A1(new_n906), .A2(new_n908), .A3(new_n773), .A4(new_n909), .ZN(new_n910));
  AND2_X1   g724(.A1(new_n740), .A2(new_n765), .ZN(new_n911));
  NAND4_X1  g725(.A1(new_n910), .A2(new_n750), .A3(new_n911), .A4(new_n743), .ZN(new_n912));
  NOR2_X1   g726(.A1(new_n905), .A2(new_n912), .ZN(new_n913));
  NAND3_X1  g727(.A1(new_n906), .A2(new_n908), .A3(new_n773), .ZN(new_n914));
  AND2_X1   g728(.A1(new_n914), .A2(KEYINPUT52), .ZN(new_n915));
  INV_X1    g729(.A(new_n915), .ZN(new_n916));
  AOI21_X1  g730(.A(KEYINPUT53), .B1(new_n913), .B2(new_n916), .ZN(new_n917));
  INV_X1    g731(.A(KEYINPUT53), .ZN(new_n918));
  NOR4_X1   g732(.A1(new_n905), .A2(new_n912), .A3(new_n915), .A4(new_n918), .ZN(new_n919));
  OAI21_X1  g733(.A(new_n880), .B1(new_n917), .B2(new_n919), .ZN(new_n920));
  AND2_X1   g734(.A1(new_n897), .A2(new_n903), .ZN(new_n921));
  NOR2_X1   g735(.A1(new_n311), .A2(new_n313), .ZN(new_n922));
  NAND4_X1  g736(.A1(new_n922), .A2(new_n656), .A3(new_n657), .A4(new_n884), .ZN(new_n923));
  NAND3_X1  g737(.A1(new_n465), .A2(new_n533), .A3(new_n652), .ZN(new_n924));
  OAI211_X1 g738(.A(new_n693), .B(new_n923), .C1(new_n886), .C2(new_n924), .ZN(new_n925));
  NOR2_X1   g739(.A1(new_n921), .A2(new_n925), .ZN(new_n926));
  AND3_X1   g740(.A1(new_n745), .A2(new_n465), .A3(new_n748), .ZN(new_n927));
  AOI21_X1  g741(.A(new_n748), .B1(new_n745), .B2(new_n465), .ZN(new_n928));
  OAI21_X1  g742(.A(new_n743), .B1(new_n927), .B2(new_n928), .ZN(new_n929));
  NAND2_X1  g743(.A1(new_n740), .A2(new_n765), .ZN(new_n930));
  NOR2_X1   g744(.A1(new_n929), .A2(new_n930), .ZN(new_n931));
  AOI21_X1  g745(.A(new_n894), .B1(new_n788), .B2(new_n796), .ZN(new_n932));
  NAND4_X1  g746(.A1(new_n926), .A2(new_n931), .A3(new_n932), .A4(new_n910), .ZN(new_n933));
  OAI21_X1  g747(.A(new_n918), .B1(new_n933), .B2(new_n915), .ZN(new_n934));
  NAND3_X1  g748(.A1(new_n913), .A2(KEYINPUT53), .A3(new_n916), .ZN(new_n935));
  NAND3_X1  g749(.A1(new_n934), .A2(new_n935), .A3(KEYINPUT54), .ZN(new_n936));
  AOI21_X1  g750(.A(new_n879), .B1(new_n920), .B2(new_n936), .ZN(new_n937));
  NAND2_X1  g751(.A1(new_n569), .A2(new_n207), .ZN(new_n938));
  XNOR2_X1  g752(.A(new_n938), .B(KEYINPUT123), .ZN(new_n939));
  OAI21_X1  g753(.A(new_n841), .B1(new_n937), .B2(new_n939), .ZN(new_n940));
  INV_X1    g754(.A(KEYINPUT124), .ZN(new_n941));
  NAND2_X1  g755(.A1(new_n940), .A2(new_n941), .ZN(new_n942));
  OAI211_X1 g756(.A(KEYINPUT124), .B(new_n841), .C1(new_n937), .C2(new_n939), .ZN(new_n943));
  NAND2_X1  g757(.A1(new_n942), .A2(new_n943), .ZN(G75));
  NAND2_X1  g758(.A1(new_n934), .A2(new_n935), .ZN(new_n945));
  NAND3_X1  g759(.A1(new_n945), .A2(G210), .A3(G902), .ZN(new_n946));
  INV_X1    g760(.A(KEYINPUT56), .ZN(new_n947));
  NOR3_X1   g761(.A1(new_n301), .A2(new_n305), .A3(new_n300), .ZN(new_n948));
  NOR2_X1   g762(.A1(new_n948), .A2(new_n274), .ZN(new_n949));
  XNOR2_X1  g763(.A(new_n949), .B(KEYINPUT55), .ZN(new_n950));
  AND3_X1   g764(.A1(new_n946), .A2(new_n947), .A3(new_n950), .ZN(new_n951));
  AOI21_X1  g765(.A(new_n950), .B1(new_n946), .B2(new_n947), .ZN(new_n952));
  NOR2_X1   g766(.A1(new_n317), .A2(G952), .ZN(new_n953));
  NOR3_X1   g767(.A1(new_n951), .A2(new_n952), .A3(new_n953), .ZN(G51));
  XNOR2_X1  g768(.A(new_n388), .B(KEYINPUT57), .ZN(new_n955));
  NAND3_X1  g769(.A1(new_n920), .A2(new_n936), .A3(new_n955), .ZN(new_n956));
  OAI21_X1  g770(.A(new_n956), .B1(new_n386), .B2(new_n379), .ZN(new_n957));
  NAND2_X1  g771(.A1(new_n945), .A2(G902), .ZN(new_n958));
  OR2_X1    g772(.A1(new_n958), .A2(new_n805), .ZN(new_n959));
  AOI21_X1  g773(.A(new_n953), .B1(new_n957), .B2(new_n959), .ZN(G54));
  NAND2_X1  g774(.A1(KEYINPUT58), .A2(G475), .ZN(new_n961));
  OAI21_X1  g775(.A(new_n647), .B1(new_n958), .B2(new_n961), .ZN(new_n962));
  INV_X1    g776(.A(new_n953), .ZN(new_n963));
  NAND2_X1  g777(.A1(new_n962), .A2(new_n963), .ZN(new_n964));
  NOR3_X1   g778(.A1(new_n958), .A2(new_n647), .A3(new_n961), .ZN(new_n965));
  NOR2_X1   g779(.A1(new_n964), .A2(new_n965), .ZN(G60));
  XNOR2_X1  g780(.A(new_n673), .B(KEYINPUT59), .ZN(new_n967));
  NAND3_X1  g781(.A1(new_n920), .A2(new_n936), .A3(new_n967), .ZN(new_n968));
  AND2_X1   g782(.A1(new_n669), .A2(new_n670), .ZN(new_n969));
  AND3_X1   g783(.A1(new_n968), .A2(KEYINPUT125), .A3(new_n969), .ZN(new_n970));
  OAI21_X1  g784(.A(new_n963), .B1(new_n968), .B2(new_n969), .ZN(new_n971));
  AOI21_X1  g785(.A(KEYINPUT125), .B1(new_n968), .B2(new_n969), .ZN(new_n972));
  NOR3_X1   g786(.A1(new_n970), .A2(new_n971), .A3(new_n972), .ZN(G63));
  NOR2_X1   g787(.A1(new_n917), .A2(new_n919), .ZN(new_n974));
  NAND2_X1  g788(.A1(G217), .A2(G902), .ZN(new_n975));
  XNOR2_X1  g789(.A(new_n975), .B(KEYINPUT60), .ZN(new_n976));
  OAI21_X1  g790(.A(new_n509), .B1(new_n974), .B2(new_n976), .ZN(new_n977));
  INV_X1    g791(.A(new_n976), .ZN(new_n978));
  NAND3_X1  g792(.A1(new_n945), .A2(new_n690), .A3(new_n978), .ZN(new_n979));
  NAND3_X1  g793(.A1(new_n977), .A2(new_n963), .A3(new_n979), .ZN(new_n980));
  INV_X1    g794(.A(KEYINPUT61), .ZN(new_n981));
  NAND2_X1  g795(.A1(new_n980), .A2(new_n981), .ZN(new_n982));
  NAND4_X1  g796(.A1(new_n977), .A2(new_n979), .A3(KEYINPUT61), .A4(new_n963), .ZN(new_n983));
  NAND2_X1  g797(.A1(new_n982), .A2(new_n983), .ZN(G66));
  INV_X1    g798(.A(new_n578), .ZN(new_n985));
  AOI21_X1  g799(.A(new_n207), .B1(new_n985), .B2(G224), .ZN(new_n986));
  NAND2_X1  g800(.A1(new_n931), .A2(new_n890), .ZN(new_n987));
  AOI21_X1  g801(.A(new_n986), .B1(new_n987), .B2(new_n317), .ZN(new_n988));
  OAI211_X1 g802(.A(new_n267), .B(new_n273), .C1(G898), .C2(new_n317), .ZN(new_n989));
  XOR2_X1   g803(.A(new_n988), .B(new_n989), .Z(G69));
  OAI22_X1  g804(.A1(new_n411), .A2(new_n412), .B1(KEYINPUT30), .B2(new_n406), .ZN(new_n991));
  XOR2_X1   g805(.A(new_n991), .B(new_n643), .Z(new_n992));
  AOI21_X1  g806(.A(new_n992), .B1(G900), .B2(new_n575), .ZN(new_n993));
  OR3_X1    g807(.A1(new_n832), .A2(new_n532), .A3(new_n763), .ZN(new_n994));
  OAI21_X1  g808(.A(new_n799), .B1(new_n994), .B2(new_n809), .ZN(new_n995));
  AOI21_X1  g809(.A(new_n995), .B1(new_n788), .B2(new_n796), .ZN(new_n996));
  AND2_X1   g810(.A1(new_n906), .A2(new_n773), .ZN(new_n997));
  NAND4_X1  g811(.A1(new_n996), .A2(new_n820), .A3(new_n834), .A4(new_n997), .ZN(new_n998));
  OAI21_X1  g812(.A(new_n993), .B1(new_n998), .B2(new_n575), .ZN(new_n999));
  NAND2_X1  g813(.A1(new_n676), .A2(new_n883), .ZN(new_n1000));
  NOR2_X1   g814(.A1(new_n713), .A2(new_n784), .ZN(new_n1001));
  NAND3_X1  g815(.A1(new_n870), .A2(new_n1000), .A3(new_n1001), .ZN(new_n1002));
  NAND3_X1  g816(.A1(new_n820), .A2(new_n834), .A3(new_n1002), .ZN(new_n1003));
  NAND2_X1  g817(.A1(new_n729), .A2(new_n997), .ZN(new_n1004));
  NOR2_X1   g818(.A1(new_n1004), .A2(KEYINPUT62), .ZN(new_n1005));
  NOR2_X1   g819(.A1(new_n1003), .A2(new_n1005), .ZN(new_n1006));
  NAND2_X1  g820(.A1(new_n1004), .A2(KEYINPUT62), .ZN(new_n1007));
  AOI21_X1  g821(.A(new_n575), .B1(new_n1006), .B2(new_n1007), .ZN(new_n1008));
  INV_X1    g822(.A(new_n992), .ZN(new_n1009));
  OAI21_X1  g823(.A(new_n999), .B1(new_n1008), .B2(new_n1009), .ZN(new_n1010));
  AOI21_X1  g824(.A(new_n317), .B1(G227), .B2(G900), .ZN(new_n1011));
  XNOR2_X1  g825(.A(new_n1011), .B(KEYINPUT127), .ZN(new_n1012));
  AOI21_X1  g826(.A(new_n1012), .B1(new_n999), .B2(KEYINPUT126), .ZN(new_n1013));
  XOR2_X1   g827(.A(new_n1010), .B(new_n1013), .Z(G72));
  NAND2_X1  g828(.A1(G472), .A2(G902), .ZN(new_n1015));
  XOR2_X1   g829(.A(new_n1015), .B(KEYINPUT63), .Z(new_n1016));
  NAND2_X1  g830(.A1(new_n413), .A2(new_n424), .ZN(new_n1017));
  OAI21_X1  g831(.A(new_n1016), .B1(new_n1017), .B2(new_n431), .ZN(new_n1018));
  NOR3_X1   g832(.A1(new_n974), .A2(new_n724), .A3(new_n1018), .ZN(new_n1019));
  OAI21_X1  g833(.A(new_n1016), .B1(new_n998), .B2(new_n987), .ZN(new_n1020));
  NAND4_X1  g834(.A1(new_n1020), .A2(new_n424), .A3(new_n432), .A4(new_n413), .ZN(new_n1021));
  NAND2_X1  g835(.A1(new_n1021), .A2(new_n963), .ZN(new_n1022));
  NAND2_X1  g836(.A1(new_n1006), .A2(new_n1007), .ZN(new_n1023));
  OAI21_X1  g837(.A(new_n1016), .B1(new_n1023), .B2(new_n987), .ZN(new_n1024));
  AOI211_X1 g838(.A(new_n1019), .B(new_n1022), .C1(new_n724), .C2(new_n1024), .ZN(G57));
endmodule


