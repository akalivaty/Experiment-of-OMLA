//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 0 0 0 0 1 0 0 1 1 0 0 1 1 0 1 0 1 0 0 1 1 1 1 1 1 0 0 0 0 0 0 0 1 0 0 0 1 0 0 1 1 0 0 1 0 1 1 0 1 0 0 0 1 0 1 1 1 0 1 1 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:41:44 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n983,
    new_n984, new_n985, new_n986, new_n987, new_n988, new_n989, new_n990,
    new_n991, new_n992, new_n993, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1025, new_n1026, new_n1027, new_n1028,
    new_n1029, new_n1030, new_n1031, new_n1032, new_n1033, new_n1034,
    new_n1035, new_n1036, new_n1037, new_n1038, new_n1039, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1053,
    new_n1054, new_n1055, new_n1056, new_n1057, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1192, new_n1193,
    new_n1194, new_n1195, new_n1196, new_n1197, new_n1198, new_n1199,
    new_n1200, new_n1201, new_n1202, new_n1203, new_n1204, new_n1205,
    new_n1206, new_n1207, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1217, new_n1218,
    new_n1219, new_n1220, new_n1221, new_n1222, new_n1223, new_n1224,
    new_n1225, new_n1226, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1288, new_n1289, new_n1290;
  INV_X1    g0000(.A(G50), .ZN(new_n201));
  INV_X1    g0001(.A(G58), .ZN(new_n202));
  INV_X1    g0002(.A(G68), .ZN(new_n203));
  NAND3_X1  g0003(.A1(new_n201), .A2(new_n202), .A3(new_n203), .ZN(new_n204));
  NOR2_X1   g0004(.A1(new_n204), .A2(G77), .ZN(G353));
  OAI21_X1  g0005(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0006(.A1(G1), .A2(G20), .ZN(new_n207));
  INV_X1    g0007(.A(G232), .ZN(new_n208));
  INV_X1    g0008(.A(G87), .ZN(new_n209));
  INV_X1    g0009(.A(G250), .ZN(new_n210));
  OAI22_X1  g0010(.A1(new_n202), .A2(new_n208), .B1(new_n209), .B2(new_n210), .ZN(new_n211));
  AOI21_X1  g0011(.A(new_n211), .B1(G97), .B2(G257), .ZN(new_n212));
  INV_X1    g0012(.A(G226), .ZN(new_n213));
  INV_X1    g0013(.A(G107), .ZN(new_n214));
  INV_X1    g0014(.A(G264), .ZN(new_n215));
  OAI22_X1  g0015(.A1(new_n201), .A2(new_n213), .B1(new_n214), .B2(new_n215), .ZN(new_n216));
  AOI21_X1  g0016(.A(new_n216), .B1(G116), .B2(G270), .ZN(new_n217));
  XNOR2_X1  g0017(.A(KEYINPUT65), .B(G244), .ZN(new_n218));
  NAND2_X1  g0018(.A1(new_n218), .A2(G77), .ZN(new_n219));
  NAND3_X1  g0019(.A1(new_n212), .A2(new_n217), .A3(new_n219), .ZN(new_n220));
  INV_X1    g0020(.A(G238), .ZN(new_n221));
  NOR2_X1   g0021(.A1(new_n203), .A2(new_n221), .ZN(new_n222));
  OAI21_X1  g0022(.A(new_n207), .B1(new_n220), .B2(new_n222), .ZN(new_n223));
  XOR2_X1   g0023(.A(new_n223), .B(KEYINPUT1), .Z(new_n224));
  NOR2_X1   g0024(.A1(new_n207), .A2(G13), .ZN(new_n225));
  INV_X1    g0025(.A(new_n225), .ZN(new_n226));
  INV_X1    g0026(.A(G257), .ZN(new_n227));
  AOI211_X1 g0027(.A(new_n210), .B(new_n226), .C1(new_n227), .C2(new_n215), .ZN(new_n228));
  NAND2_X1  g0028(.A1(G1), .A2(G13), .ZN(new_n229));
  INV_X1    g0029(.A(G20), .ZN(new_n230));
  NOR2_X1   g0030(.A1(new_n229), .A2(new_n230), .ZN(new_n231));
  OAI21_X1  g0031(.A(G50), .B1(G58), .B2(G68), .ZN(new_n232));
  XOR2_X1   g0032(.A(new_n232), .B(KEYINPUT64), .Z(new_n233));
  AOI22_X1  g0033(.A1(new_n228), .A2(KEYINPUT0), .B1(new_n231), .B2(new_n233), .ZN(new_n234));
  OAI211_X1 g0034(.A(new_n224), .B(new_n234), .C1(KEYINPUT0), .C2(new_n228), .ZN(new_n235));
  INV_X1    g0035(.A(new_n235), .ZN(G361));
  XNOR2_X1  g0036(.A(G238), .B(G244), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n237), .B(G232), .ZN(new_n238));
  XNOR2_X1  g0038(.A(KEYINPUT2), .B(G226), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XOR2_X1   g0040(.A(G250), .B(G257), .Z(new_n241));
  XNOR2_X1  g0041(.A(G264), .B(G270), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n240), .B(new_n243), .ZN(G358));
  XOR2_X1   g0044(.A(G68), .B(G77), .Z(new_n245));
  XNOR2_X1  g0045(.A(G50), .B(G58), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n245), .B(new_n246), .ZN(new_n247));
  XOR2_X1   g0047(.A(G87), .B(G97), .Z(new_n248));
  XNOR2_X1  g0048(.A(G107), .B(G116), .ZN(new_n249));
  XNOR2_X1  g0049(.A(new_n248), .B(new_n249), .ZN(new_n250));
  XNOR2_X1  g0050(.A(new_n247), .B(new_n250), .ZN(G351));
  INV_X1    g0051(.A(G13), .ZN(new_n252));
  NOR3_X1   g0052(.A1(new_n252), .A2(new_n230), .A3(G1), .ZN(new_n253));
  NAND2_X1  g0053(.A1(new_n253), .A2(new_n201), .ZN(new_n254));
  OAI21_X1  g0054(.A(G50), .B1(new_n230), .B2(G1), .ZN(new_n255));
  XNOR2_X1  g0055(.A(new_n255), .B(KEYINPUT68), .ZN(new_n256));
  NAND3_X1  g0056(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n257));
  NAND2_X1  g0057(.A1(new_n257), .A2(new_n229), .ZN(new_n258));
  NOR2_X1   g0058(.A1(new_n253), .A2(new_n258), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n256), .A2(new_n259), .ZN(new_n260));
  INV_X1    g0060(.A(KEYINPUT67), .ZN(new_n261));
  INV_X1    g0061(.A(G33), .ZN(new_n262));
  NAND3_X1  g0062(.A1(new_n261), .A2(new_n230), .A3(new_n262), .ZN(new_n263));
  OAI21_X1  g0063(.A(KEYINPUT67), .B1(G20), .B2(G33), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n263), .A2(new_n264), .ZN(new_n265));
  INV_X1    g0065(.A(new_n265), .ZN(new_n266));
  INV_X1    g0066(.A(G150), .ZN(new_n267));
  XNOR2_X1  g0067(.A(KEYINPUT8), .B(G58), .ZN(new_n268));
  NAND2_X1  g0068(.A1(new_n230), .A2(G33), .ZN(new_n269));
  OAI22_X1  g0069(.A1(new_n266), .A2(new_n267), .B1(new_n268), .B2(new_n269), .ZN(new_n270));
  AOI21_X1  g0070(.A(new_n270), .B1(G20), .B2(new_n204), .ZN(new_n271));
  INV_X1    g0071(.A(new_n258), .ZN(new_n272));
  OAI211_X1 g0072(.A(new_n254), .B(new_n260), .C1(new_n271), .C2(new_n272), .ZN(new_n273));
  XNOR2_X1  g0073(.A(KEYINPUT3), .B(G33), .ZN(new_n274));
  NAND2_X1  g0074(.A1(G223), .A2(G1698), .ZN(new_n275));
  INV_X1    g0075(.A(G1698), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n276), .A2(G222), .ZN(new_n277));
  NAND3_X1  g0077(.A1(new_n274), .A2(new_n275), .A3(new_n277), .ZN(new_n278));
  AOI21_X1  g0078(.A(new_n229), .B1(G33), .B2(G41), .ZN(new_n279));
  OAI211_X1 g0079(.A(new_n278), .B(new_n279), .C1(G77), .C2(new_n274), .ZN(new_n280));
  INV_X1    g0080(.A(G1), .ZN(new_n281));
  OAI211_X1 g0081(.A(new_n281), .B(G274), .C1(G41), .C2(G45), .ZN(new_n282));
  INV_X1    g0082(.A(KEYINPUT66), .ZN(new_n283));
  XNOR2_X1  g0083(.A(new_n282), .B(new_n283), .ZN(new_n284));
  INV_X1    g0084(.A(G41), .ZN(new_n285));
  INV_X1    g0085(.A(G45), .ZN(new_n286));
  AOI21_X1  g0086(.A(G1), .B1(new_n285), .B2(new_n286), .ZN(new_n287));
  NOR2_X1   g0087(.A1(new_n279), .A2(new_n287), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n288), .A2(G226), .ZN(new_n289));
  NAND3_X1  g0089(.A1(new_n280), .A2(new_n284), .A3(new_n289), .ZN(new_n290));
  INV_X1    g0090(.A(new_n290), .ZN(new_n291));
  INV_X1    g0091(.A(G179), .ZN(new_n292));
  AND3_X1   g0092(.A1(new_n291), .A2(KEYINPUT69), .A3(new_n292), .ZN(new_n293));
  AOI21_X1  g0093(.A(KEYINPUT69), .B1(new_n291), .B2(new_n292), .ZN(new_n294));
  OAI221_X1 g0094(.A(new_n273), .B1(G169), .B2(new_n291), .C1(new_n293), .C2(new_n294), .ZN(new_n295));
  INV_X1    g0095(.A(new_n295), .ZN(new_n296));
  INV_X1    g0096(.A(KEYINPUT9), .ZN(new_n297));
  OR2_X1    g0097(.A1(new_n273), .A2(new_n297), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n290), .A2(G200), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n291), .A2(G190), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n273), .A2(new_n297), .ZN(new_n301));
  NAND4_X1  g0101(.A1(new_n298), .A2(new_n299), .A3(new_n300), .A4(new_n301), .ZN(new_n302));
  OR2_X1    g0102(.A1(new_n302), .A2(KEYINPUT10), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n302), .A2(KEYINPUT10), .ZN(new_n304));
  AOI21_X1  g0104(.A(new_n296), .B1(new_n303), .B2(new_n304), .ZN(new_n305));
  NAND2_X1  g0105(.A1(G33), .A2(G97), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n208), .A2(G1698), .ZN(new_n307));
  OAI21_X1  g0107(.A(new_n307), .B1(G226), .B2(G1698), .ZN(new_n308));
  INV_X1    g0108(.A(KEYINPUT3), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n309), .A2(G33), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n262), .A2(KEYINPUT3), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n310), .A2(new_n311), .ZN(new_n312));
  OAI21_X1  g0112(.A(new_n306), .B1(new_n308), .B2(new_n312), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n313), .A2(new_n279), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n288), .A2(G238), .ZN(new_n315));
  NAND3_X1  g0115(.A1(new_n314), .A2(new_n284), .A3(new_n315), .ZN(new_n316));
  OR2_X1    g0116(.A1(new_n316), .A2(KEYINPUT13), .ZN(new_n317));
  INV_X1    g0117(.A(KEYINPUT71), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n316), .A2(KEYINPUT13), .ZN(new_n319));
  NAND3_X1  g0119(.A1(new_n317), .A2(new_n318), .A3(new_n319), .ZN(new_n320));
  OR3_X1    g0120(.A1(new_n316), .A2(new_n318), .A3(KEYINPUT13), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n320), .A2(new_n321), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n322), .A2(G179), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n317), .A2(new_n319), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n324), .A2(G169), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n325), .A2(KEYINPUT14), .ZN(new_n326));
  INV_X1    g0126(.A(KEYINPUT14), .ZN(new_n327));
  NAND3_X1  g0127(.A1(new_n324), .A2(new_n327), .A3(G169), .ZN(new_n328));
  NAND3_X1  g0128(.A1(new_n323), .A2(new_n326), .A3(new_n328), .ZN(new_n329));
  OAI21_X1  g0129(.A(new_n272), .B1(G1), .B2(new_n230), .ZN(new_n330));
  OR2_X1    g0130(.A1(new_n330), .A2(new_n203), .ZN(new_n331));
  XOR2_X1   g0131(.A(new_n331), .B(KEYINPUT73), .Z(new_n332));
  INV_X1    g0132(.A(new_n332), .ZN(new_n333));
  NOR2_X1   g0133(.A1(new_n252), .A2(G1), .ZN(new_n334));
  NAND3_X1  g0134(.A1(new_n334), .A2(G20), .A3(new_n203), .ZN(new_n335));
  XOR2_X1   g0135(.A(new_n335), .B(KEYINPUT12), .Z(new_n336));
  INV_X1    g0136(.A(new_n336), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n265), .A2(G50), .ZN(new_n338));
  AOI22_X1  g0138(.A1(new_n338), .A2(KEYINPUT72), .B1(G20), .B2(new_n203), .ZN(new_n339));
  INV_X1    g0139(.A(G77), .ZN(new_n340));
  OAI221_X1 g0140(.A(new_n339), .B1(KEYINPUT72), .B2(new_n338), .C1(new_n340), .C2(new_n269), .ZN(new_n341));
  INV_X1    g0141(.A(KEYINPUT11), .ZN(new_n342));
  NAND3_X1  g0142(.A1(new_n341), .A2(new_n342), .A3(new_n258), .ZN(new_n343));
  INV_X1    g0143(.A(new_n343), .ZN(new_n344));
  AOI21_X1  g0144(.A(new_n342), .B1(new_n341), .B2(new_n258), .ZN(new_n345));
  OAI211_X1 g0145(.A(new_n333), .B(new_n337), .C1(new_n344), .C2(new_n345), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n329), .A2(new_n346), .ZN(new_n347));
  INV_X1    g0147(.A(G190), .ZN(new_n348));
  AOI21_X1  g0148(.A(new_n348), .B1(new_n320), .B2(new_n321), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n324), .A2(G200), .ZN(new_n350));
  INV_X1    g0150(.A(new_n350), .ZN(new_n351));
  NOR3_X1   g0151(.A1(new_n346), .A2(new_n349), .A3(new_n351), .ZN(new_n352));
  INV_X1    g0152(.A(new_n352), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n288), .A2(new_n218), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n354), .A2(new_n284), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n355), .A2(KEYINPUT70), .ZN(new_n356));
  NAND2_X1  g0156(.A1(G238), .A2(G1698), .ZN(new_n357));
  OAI211_X1 g0157(.A(new_n274), .B(new_n357), .C1(new_n208), .C2(G1698), .ZN(new_n358));
  OAI211_X1 g0158(.A(new_n358), .B(new_n279), .C1(G107), .C2(new_n274), .ZN(new_n359));
  INV_X1    g0159(.A(KEYINPUT70), .ZN(new_n360));
  NAND3_X1  g0160(.A1(new_n354), .A2(new_n284), .A3(new_n360), .ZN(new_n361));
  AND3_X1   g0161(.A1(new_n356), .A2(new_n359), .A3(new_n361), .ZN(new_n362));
  OR2_X1    g0162(.A1(new_n362), .A2(G169), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n334), .A2(G20), .ZN(new_n364));
  NOR2_X1   g0164(.A1(new_n364), .A2(G77), .ZN(new_n365));
  NOR2_X1   g0165(.A1(new_n330), .A2(new_n340), .ZN(new_n366));
  INV_X1    g0166(.A(new_n268), .ZN(new_n367));
  AOI22_X1  g0167(.A1(new_n367), .A2(new_n265), .B1(G20), .B2(G77), .ZN(new_n368));
  XOR2_X1   g0168(.A(KEYINPUT15), .B(G87), .Z(new_n369));
  INV_X1    g0169(.A(new_n369), .ZN(new_n370));
  OAI21_X1  g0170(.A(new_n368), .B1(new_n269), .B2(new_n370), .ZN(new_n371));
  AOI211_X1 g0171(.A(new_n365), .B(new_n366), .C1(new_n371), .C2(new_n258), .ZN(new_n372));
  AOI21_X1  g0172(.A(new_n372), .B1(new_n362), .B2(new_n292), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n363), .A2(new_n373), .ZN(new_n374));
  NAND4_X1  g0174(.A1(new_n305), .A2(new_n347), .A3(new_n353), .A4(new_n374), .ZN(new_n375));
  INV_X1    g0175(.A(KEYINPUT18), .ZN(new_n376));
  NOR2_X1   g0176(.A1(new_n367), .A2(new_n253), .ZN(new_n377));
  AOI21_X1  g0177(.A(new_n377), .B1(new_n367), .B2(new_n330), .ZN(new_n378));
  NAND3_X1  g0178(.A1(new_n309), .A2(KEYINPUT74), .A3(G33), .ZN(new_n379));
  INV_X1    g0179(.A(KEYINPUT74), .ZN(new_n380));
  AOI21_X1  g0180(.A(new_n380), .B1(KEYINPUT3), .B2(new_n262), .ZN(new_n381));
  NOR2_X1   g0181(.A1(new_n262), .A2(KEYINPUT3), .ZN(new_n382));
  OAI21_X1  g0182(.A(new_n379), .B1(new_n381), .B2(new_n382), .ZN(new_n383));
  XNOR2_X1  g0183(.A(KEYINPUT75), .B(KEYINPUT7), .ZN(new_n384));
  NAND3_X1  g0184(.A1(new_n383), .A2(new_n230), .A3(new_n384), .ZN(new_n385));
  INV_X1    g0185(.A(KEYINPUT7), .ZN(new_n386));
  OAI21_X1  g0186(.A(KEYINPUT74), .B1(new_n309), .B2(G33), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n387), .A2(new_n310), .ZN(new_n388));
  AOI21_X1  g0188(.A(G20), .B1(new_n388), .B2(new_n379), .ZN(new_n389));
  OAI211_X1 g0189(.A(new_n385), .B(G68), .C1(new_n386), .C2(new_n389), .ZN(new_n390));
  XNOR2_X1  g0190(.A(G58), .B(G68), .ZN(new_n391));
  AOI22_X1  g0191(.A1(new_n265), .A2(G159), .B1(new_n391), .B2(G20), .ZN(new_n392));
  NAND3_X1  g0192(.A1(new_n390), .A2(KEYINPUT16), .A3(new_n392), .ZN(new_n393));
  AND2_X1   g0193(.A1(new_n393), .A2(new_n258), .ZN(new_n394));
  OAI21_X1  g0194(.A(new_n384), .B1(new_n274), .B2(G20), .ZN(new_n395));
  NOR2_X1   g0195(.A1(new_n309), .A2(G33), .ZN(new_n396));
  OAI211_X1 g0196(.A(KEYINPUT7), .B(new_n230), .C1(new_n382), .C2(new_n396), .ZN(new_n397));
  NAND2_X1  g0197(.A1(new_n395), .A2(new_n397), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n398), .A2(G68), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n399), .A2(KEYINPUT76), .ZN(new_n400));
  INV_X1    g0200(.A(KEYINPUT76), .ZN(new_n401));
  NAND3_X1  g0201(.A1(new_n398), .A2(new_n401), .A3(G68), .ZN(new_n402));
  NAND3_X1  g0202(.A1(new_n400), .A2(new_n392), .A3(new_n402), .ZN(new_n403));
  INV_X1    g0203(.A(KEYINPUT16), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n403), .A2(new_n404), .ZN(new_n405));
  AOI21_X1  g0205(.A(new_n378), .B1(new_n394), .B2(new_n405), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n213), .A2(G1698), .ZN(new_n407));
  OR2_X1    g0207(.A1(G223), .A2(G1698), .ZN(new_n408));
  NAND4_X1  g0208(.A1(new_n388), .A2(new_n379), .A3(new_n407), .A4(new_n408), .ZN(new_n409));
  OAI21_X1  g0209(.A(new_n409), .B1(new_n262), .B2(new_n209), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n410), .A2(new_n279), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n288), .A2(G232), .ZN(new_n412));
  NAND3_X1  g0212(.A1(new_n411), .A2(new_n412), .A3(new_n284), .ZN(new_n413));
  NAND2_X1  g0213(.A1(new_n413), .A2(G169), .ZN(new_n414));
  NAND4_X1  g0214(.A1(new_n411), .A2(G179), .A3(new_n412), .A4(new_n284), .ZN(new_n415));
  AND2_X1   g0215(.A1(new_n414), .A2(new_n415), .ZN(new_n416));
  OAI21_X1  g0216(.A(new_n376), .B1(new_n406), .B2(new_n416), .ZN(new_n417));
  INV_X1    g0217(.A(new_n378), .ZN(new_n418));
  AOI21_X1  g0218(.A(new_n401), .B1(new_n398), .B2(G68), .ZN(new_n419));
  AOI211_X1 g0219(.A(KEYINPUT76), .B(new_n203), .C1(new_n395), .C2(new_n397), .ZN(new_n420));
  NOR2_X1   g0220(.A1(new_n419), .A2(new_n420), .ZN(new_n421));
  AOI21_X1  g0221(.A(KEYINPUT16), .B1(new_n421), .B2(new_n392), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n393), .A2(new_n258), .ZN(new_n423));
  OAI21_X1  g0223(.A(new_n418), .B1(new_n422), .B2(new_n423), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n414), .A2(new_n415), .ZN(new_n425));
  NAND3_X1  g0225(.A1(new_n424), .A2(KEYINPUT18), .A3(new_n425), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n417), .A2(new_n426), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n413), .A2(G200), .ZN(new_n428));
  OAI211_X1 g0228(.A(new_n418), .B(new_n428), .C1(new_n422), .C2(new_n423), .ZN(new_n429));
  INV_X1    g0229(.A(new_n429), .ZN(new_n430));
  INV_X1    g0230(.A(KEYINPUT17), .ZN(new_n431));
  OR2_X1    g0231(.A1(new_n431), .A2(KEYINPUT77), .ZN(new_n432));
  NOR2_X1   g0232(.A1(new_n413), .A2(new_n348), .ZN(new_n433));
  INV_X1    g0233(.A(new_n433), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n431), .A2(KEYINPUT77), .ZN(new_n435));
  NAND4_X1  g0235(.A1(new_n430), .A2(new_n432), .A3(new_n434), .A4(new_n435), .ZN(new_n436));
  OAI211_X1 g0236(.A(KEYINPUT77), .B(new_n431), .C1(new_n429), .C2(new_n433), .ZN(new_n437));
  NAND2_X1  g0237(.A1(new_n362), .A2(G190), .ZN(new_n438));
  INV_X1    g0238(.A(G200), .ZN(new_n439));
  OAI211_X1 g0239(.A(new_n438), .B(new_n372), .C1(new_n362), .C2(new_n439), .ZN(new_n440));
  NAND4_X1  g0240(.A1(new_n427), .A2(new_n436), .A3(new_n437), .A4(new_n440), .ZN(new_n441));
  NOR2_X1   g0241(.A1(new_n209), .A2(G20), .ZN(new_n442));
  NAND4_X1  g0242(.A1(new_n388), .A2(KEYINPUT22), .A3(new_n379), .A4(new_n442), .ZN(new_n443));
  INV_X1    g0243(.A(G116), .ZN(new_n444));
  NOR3_X1   g0244(.A1(new_n262), .A2(new_n444), .A3(G20), .ZN(new_n445));
  NAND3_X1  g0245(.A1(new_n442), .A2(new_n310), .A3(new_n311), .ZN(new_n446));
  INV_X1    g0246(.A(KEYINPUT22), .ZN(new_n447));
  AOI21_X1  g0247(.A(new_n445), .B1(new_n446), .B2(new_n447), .ZN(new_n448));
  NOR2_X1   g0248(.A1(new_n230), .A2(G107), .ZN(new_n449));
  INV_X1    g0249(.A(KEYINPUT23), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n450), .A2(KEYINPUT88), .ZN(new_n451));
  INV_X1    g0251(.A(KEYINPUT88), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n452), .A2(KEYINPUT23), .ZN(new_n453));
  NAND3_X1  g0253(.A1(new_n449), .A2(new_n451), .A3(new_n453), .ZN(new_n454));
  OAI211_X1 g0254(.A(KEYINPUT88), .B(new_n450), .C1(new_n230), .C2(G107), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n454), .A2(new_n455), .ZN(new_n456));
  NAND3_X1  g0256(.A1(new_n443), .A2(new_n448), .A3(new_n456), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n457), .A2(KEYINPUT24), .ZN(new_n458));
  INV_X1    g0258(.A(KEYINPUT24), .ZN(new_n459));
  NAND4_X1  g0259(.A1(new_n443), .A2(new_n448), .A3(new_n459), .A4(new_n456), .ZN(new_n460));
  AOI21_X1  g0260(.A(new_n272), .B1(new_n458), .B2(new_n460), .ZN(new_n461));
  NAND2_X1  g0261(.A1(new_n334), .A2(new_n449), .ZN(new_n462));
  INV_X1    g0262(.A(new_n462), .ZN(new_n463));
  INV_X1    g0263(.A(KEYINPUT25), .ZN(new_n464));
  NOR2_X1   g0264(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n281), .A2(G33), .ZN(new_n466));
  NAND3_X1  g0266(.A1(new_n272), .A2(new_n364), .A3(new_n466), .ZN(new_n467));
  INV_X1    g0267(.A(new_n467), .ZN(new_n468));
  AOI22_X1  g0268(.A1(new_n468), .A2(G107), .B1(new_n464), .B2(new_n463), .ZN(new_n469));
  INV_X1    g0269(.A(new_n469), .ZN(new_n470));
  NOR3_X1   g0270(.A1(new_n461), .A2(new_n465), .A3(new_n470), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n227), .A2(G1698), .ZN(new_n472));
  NAND2_X1  g0272(.A1(new_n210), .A2(new_n276), .ZN(new_n473));
  NAND4_X1  g0273(.A1(new_n388), .A2(new_n379), .A3(new_n472), .A4(new_n473), .ZN(new_n474));
  INV_X1    g0274(.A(G294), .ZN(new_n475));
  OAI21_X1  g0275(.A(new_n474), .B1(new_n262), .B2(new_n475), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n476), .A2(new_n279), .ZN(new_n477));
  INV_X1    g0277(.A(KEYINPUT81), .ZN(new_n478));
  NOR2_X1   g0278(.A1(new_n285), .A2(KEYINPUT5), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n281), .A2(G45), .ZN(new_n480));
  OAI21_X1  g0280(.A(new_n478), .B1(new_n479), .B2(new_n480), .ZN(new_n481));
  NOR2_X1   g0281(.A1(new_n286), .A2(G1), .ZN(new_n482));
  INV_X1    g0282(.A(KEYINPUT5), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n483), .A2(G41), .ZN(new_n484));
  NAND3_X1  g0284(.A1(new_n482), .A2(KEYINPUT81), .A3(new_n484), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n285), .A2(KEYINPUT5), .ZN(new_n486));
  NAND4_X1  g0286(.A1(new_n481), .A2(new_n485), .A3(G274), .A4(new_n486), .ZN(new_n487));
  NOR2_X1   g0287(.A1(new_n487), .A2(new_n279), .ZN(new_n488));
  INV_X1    g0288(.A(new_n488), .ZN(new_n489));
  NAND3_X1  g0289(.A1(new_n481), .A2(new_n486), .A3(new_n485), .ZN(new_n490));
  INV_X1    g0290(.A(new_n279), .ZN(new_n491));
  NAND3_X1  g0291(.A1(new_n490), .A2(G264), .A3(new_n491), .ZN(new_n492));
  NAND3_X1  g0292(.A1(new_n477), .A2(new_n489), .A3(new_n492), .ZN(new_n493));
  INV_X1    g0293(.A(G169), .ZN(new_n494));
  AND2_X1   g0294(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  NOR2_X1   g0295(.A1(new_n493), .A2(G179), .ZN(new_n496));
  NOR3_X1   g0296(.A1(new_n471), .A2(new_n495), .A3(new_n496), .ZN(new_n497));
  NAND3_X1  g0297(.A1(new_n490), .A2(G270), .A3(new_n491), .ZN(new_n498));
  OAI21_X1  g0298(.A(new_n498), .B1(new_n279), .B2(new_n487), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n215), .A2(G1698), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n227), .A2(new_n276), .ZN(new_n501));
  NAND4_X1  g0301(.A1(new_n388), .A2(new_n379), .A3(new_n500), .A4(new_n501), .ZN(new_n502));
  XNOR2_X1  g0302(.A(KEYINPUT87), .B(G303), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n312), .A2(new_n503), .ZN(new_n504));
  AOI21_X1  g0304(.A(new_n491), .B1(new_n502), .B2(new_n504), .ZN(new_n505));
  OAI21_X1  g0305(.A(G200), .B1(new_n499), .B2(new_n505), .ZN(new_n506));
  INV_X1    g0306(.A(new_n505), .ZN(new_n507));
  NAND4_X1  g0307(.A1(new_n507), .A2(new_n489), .A3(G190), .A4(new_n498), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n253), .A2(new_n444), .ZN(new_n509));
  NAND3_X1  g0309(.A1(new_n259), .A2(G116), .A3(new_n466), .ZN(new_n510));
  AOI21_X1  g0310(.A(G20), .B1(new_n262), .B2(G97), .ZN(new_n511));
  NAND3_X1  g0311(.A1(KEYINPUT79), .A2(G33), .A3(G283), .ZN(new_n512));
  INV_X1    g0312(.A(new_n512), .ZN(new_n513));
  AOI21_X1  g0313(.A(KEYINPUT79), .B1(G33), .B2(G283), .ZN(new_n514));
  OAI21_X1  g0314(.A(new_n511), .B1(new_n513), .B2(new_n514), .ZN(new_n515));
  AOI22_X1  g0315(.A1(new_n257), .A2(new_n229), .B1(G20), .B2(new_n444), .ZN(new_n516));
  AND3_X1   g0316(.A1(new_n515), .A2(KEYINPUT20), .A3(new_n516), .ZN(new_n517));
  AOI21_X1  g0317(.A(KEYINPUT20), .B1(new_n515), .B2(new_n516), .ZN(new_n518));
  OAI211_X1 g0318(.A(new_n509), .B(new_n510), .C1(new_n517), .C2(new_n518), .ZN(new_n519));
  INV_X1    g0319(.A(new_n519), .ZN(new_n520));
  NAND3_X1  g0320(.A1(new_n506), .A2(new_n508), .A3(new_n520), .ZN(new_n521));
  OAI211_X1 g0321(.A(new_n519), .B(G169), .C1(new_n499), .C2(new_n505), .ZN(new_n522));
  INV_X1    g0322(.A(KEYINPUT21), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  NOR2_X1   g0324(.A1(new_n499), .A2(new_n505), .ZN(new_n525));
  NAND3_X1  g0325(.A1(new_n525), .A2(G179), .A3(new_n519), .ZN(new_n526));
  NAND3_X1  g0326(.A1(new_n507), .A2(new_n489), .A3(new_n498), .ZN(new_n527));
  NAND4_X1  g0327(.A1(new_n527), .A2(KEYINPUT21), .A3(G169), .A4(new_n519), .ZN(new_n528));
  NAND4_X1  g0328(.A1(new_n521), .A2(new_n524), .A3(new_n526), .A4(new_n528), .ZN(new_n529));
  NOR2_X1   g0329(.A1(new_n497), .A2(new_n529), .ZN(new_n530));
  NOR2_X1   g0330(.A1(new_n369), .A2(new_n364), .ZN(new_n531));
  NOR2_X1   g0331(.A1(new_n467), .A2(new_n209), .ZN(new_n532));
  NAND4_X1  g0332(.A1(new_n388), .A2(new_n230), .A3(G68), .A4(new_n379), .ZN(new_n533));
  INV_X1    g0333(.A(KEYINPUT19), .ZN(new_n534));
  OAI21_X1  g0334(.A(new_n230), .B1(new_n306), .B2(new_n534), .ZN(new_n535));
  NOR4_X1   g0335(.A1(KEYINPUT86), .A2(G87), .A3(G97), .A4(G107), .ZN(new_n536));
  INV_X1    g0336(.A(KEYINPUT86), .ZN(new_n537));
  NOR2_X1   g0337(.A1(G87), .A2(G97), .ZN(new_n538));
  AOI21_X1  g0338(.A(new_n537), .B1(new_n538), .B2(new_n214), .ZN(new_n539));
  OAI21_X1  g0339(.A(new_n535), .B1(new_n536), .B2(new_n539), .ZN(new_n540));
  INV_X1    g0340(.A(G97), .ZN(new_n541));
  OAI21_X1  g0341(.A(new_n534), .B1(new_n269), .B2(new_n541), .ZN(new_n542));
  NAND3_X1  g0342(.A1(new_n533), .A2(new_n540), .A3(new_n542), .ZN(new_n543));
  AOI211_X1 g0343(.A(new_n531), .B(new_n532), .C1(new_n543), .C2(new_n258), .ZN(new_n544));
  AOI21_X1  g0344(.A(new_n210), .B1(new_n482), .B2(KEYINPUT85), .ZN(new_n545));
  OAI211_X1 g0345(.A(new_n491), .B(new_n545), .C1(KEYINPUT85), .C2(new_n482), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n482), .A2(G274), .ZN(new_n547));
  INV_X1    g0347(.A(KEYINPUT84), .ZN(new_n548));
  XNOR2_X1  g0348(.A(new_n547), .B(new_n548), .ZN(new_n549));
  NOR2_X1   g0349(.A1(new_n262), .A2(new_n444), .ZN(new_n550));
  AND3_X1   g0350(.A1(new_n309), .A2(KEYINPUT74), .A3(G33), .ZN(new_n551));
  AOI21_X1  g0351(.A(new_n551), .B1(new_n310), .B2(new_n387), .ZN(new_n552));
  NOR2_X1   g0352(.A1(G238), .A2(G1698), .ZN(new_n553));
  INV_X1    g0353(.A(G244), .ZN(new_n554));
  AOI21_X1  g0354(.A(new_n553), .B1(new_n554), .B2(G1698), .ZN(new_n555));
  AOI21_X1  g0355(.A(new_n550), .B1(new_n552), .B2(new_n555), .ZN(new_n556));
  OAI211_X1 g0356(.A(new_n546), .B(new_n549), .C1(new_n556), .C2(new_n491), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n557), .A2(G200), .ZN(new_n558));
  AND3_X1   g0358(.A1(new_n388), .A2(new_n555), .A3(new_n379), .ZN(new_n559));
  OAI21_X1  g0359(.A(new_n279), .B1(new_n559), .B2(new_n550), .ZN(new_n560));
  NAND4_X1  g0360(.A1(new_n560), .A2(G190), .A3(new_n546), .A4(new_n549), .ZN(new_n561));
  NAND3_X1  g0361(.A1(new_n544), .A2(new_n558), .A3(new_n561), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n557), .A2(new_n494), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n543), .A2(new_n258), .ZN(new_n564));
  INV_X1    g0364(.A(new_n531), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n468), .A2(new_n369), .ZN(new_n566));
  NAND3_X1  g0366(.A1(new_n564), .A2(new_n565), .A3(new_n566), .ZN(new_n567));
  NAND4_X1  g0367(.A1(new_n560), .A2(new_n292), .A3(new_n546), .A4(new_n549), .ZN(new_n568));
  NAND3_X1  g0368(.A1(new_n563), .A2(new_n567), .A3(new_n568), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n562), .A2(new_n569), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n493), .A2(G200), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n458), .A2(new_n460), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n572), .A2(new_n258), .ZN(new_n573));
  INV_X1    g0373(.A(new_n465), .ZN(new_n574));
  AND4_X1   g0374(.A1(new_n571), .A2(new_n573), .A3(new_n574), .A4(new_n469), .ZN(new_n575));
  INV_X1    g0375(.A(new_n493), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n576), .A2(G190), .ZN(new_n577));
  AOI21_X1  g0377(.A(new_n570), .B1(new_n575), .B2(new_n577), .ZN(new_n578));
  NOR2_X1   g0378(.A1(new_n364), .A2(G97), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n579), .A2(KEYINPUT78), .ZN(new_n580));
  OAI22_X1  g0380(.A1(new_n467), .A2(new_n541), .B1(new_n579), .B2(KEYINPUT78), .ZN(new_n581));
  INV_X1    g0381(.A(new_n581), .ZN(new_n582));
  AOI21_X1  g0382(.A(new_n214), .B1(new_n395), .B2(new_n397), .ZN(new_n583));
  INV_X1    g0383(.A(KEYINPUT6), .ZN(new_n584));
  NOR2_X1   g0384(.A1(new_n541), .A2(new_n214), .ZN(new_n585));
  NOR2_X1   g0385(.A1(G97), .A2(G107), .ZN(new_n586));
  OAI21_X1  g0386(.A(new_n584), .B1(new_n585), .B2(new_n586), .ZN(new_n587));
  NAND3_X1  g0387(.A1(new_n214), .A2(KEYINPUT6), .A3(G97), .ZN(new_n588));
  AOI21_X1  g0388(.A(new_n230), .B1(new_n587), .B2(new_n588), .ZN(new_n589));
  NOR2_X1   g0389(.A1(new_n266), .A2(new_n340), .ZN(new_n590));
  NOR3_X1   g0390(.A1(new_n583), .A2(new_n589), .A3(new_n590), .ZN(new_n591));
  OAI211_X1 g0391(.A(new_n580), .B(new_n582), .C1(new_n591), .C2(new_n272), .ZN(new_n592));
  NOR3_X1   g0392(.A1(new_n554), .A2(KEYINPUT4), .A3(G1698), .ZN(new_n593));
  OAI211_X1 g0393(.A(new_n379), .B(new_n593), .C1(new_n381), .C2(new_n382), .ZN(new_n594));
  NOR2_X1   g0394(.A1(new_n554), .A2(G1698), .ZN(new_n595));
  NAND3_X1  g0395(.A1(new_n595), .A2(new_n310), .A3(new_n311), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n596), .A2(KEYINPUT4), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n594), .A2(new_n597), .ZN(new_n598));
  NOR2_X1   g0398(.A1(new_n210), .A2(new_n276), .ZN(new_n599));
  INV_X1    g0399(.A(new_n514), .ZN(new_n600));
  AOI22_X1  g0400(.A1(new_n274), .A2(new_n599), .B1(new_n600), .B2(new_n512), .ZN(new_n601));
  AND3_X1   g0401(.A1(new_n598), .A2(KEYINPUT80), .A3(new_n601), .ZN(new_n602));
  AOI21_X1  g0402(.A(KEYINPUT80), .B1(new_n598), .B2(new_n601), .ZN(new_n603));
  NOR3_X1   g0403(.A1(new_n602), .A2(new_n603), .A3(new_n491), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n490), .A2(new_n491), .ZN(new_n605));
  OAI21_X1  g0405(.A(new_n489), .B1(new_n227), .B2(new_n605), .ZN(new_n606));
  NOR2_X1   g0406(.A1(new_n604), .A2(new_n606), .ZN(new_n607));
  AOI21_X1  g0407(.A(new_n592), .B1(new_n607), .B2(G190), .ZN(new_n608));
  OAI21_X1  g0408(.A(G200), .B1(new_n604), .B2(new_n606), .ZN(new_n609));
  INV_X1    g0409(.A(KEYINPUT82), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n609), .A2(new_n610), .ZN(new_n611));
  INV_X1    g0411(.A(new_n603), .ZN(new_n612));
  NAND3_X1  g0412(.A1(new_n598), .A2(KEYINPUT80), .A3(new_n601), .ZN(new_n613));
  NAND3_X1  g0413(.A1(new_n612), .A2(new_n279), .A3(new_n613), .ZN(new_n614));
  INV_X1    g0414(.A(new_n605), .ZN(new_n615));
  AOI21_X1  g0415(.A(new_n488), .B1(new_n615), .B2(G257), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n614), .A2(new_n616), .ZN(new_n617));
  NAND3_X1  g0417(.A1(new_n617), .A2(KEYINPUT82), .A3(G200), .ZN(new_n618));
  NAND3_X1  g0418(.A1(new_n608), .A2(new_n611), .A3(new_n618), .ZN(new_n619));
  OAI21_X1  g0419(.A(G169), .B1(new_n604), .B2(new_n606), .ZN(new_n620));
  NAND3_X1  g0420(.A1(new_n614), .A2(G179), .A3(new_n616), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  INV_X1    g0422(.A(KEYINPUT83), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n592), .A2(new_n623), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n398), .A2(G107), .ZN(new_n625));
  INV_X1    g0425(.A(new_n589), .ZN(new_n626));
  INV_X1    g0426(.A(new_n590), .ZN(new_n627));
  NAND3_X1  g0427(.A1(new_n625), .A2(new_n626), .A3(new_n627), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n628), .A2(new_n258), .ZN(new_n629));
  NAND4_X1  g0429(.A1(new_n629), .A2(KEYINPUT83), .A3(new_n580), .A4(new_n582), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n624), .A2(new_n630), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n622), .A2(new_n631), .ZN(new_n632));
  NAND4_X1  g0432(.A1(new_n530), .A2(new_n578), .A3(new_n619), .A4(new_n632), .ZN(new_n633));
  NOR3_X1   g0433(.A1(new_n375), .A2(new_n441), .A3(new_n633), .ZN(G372));
  NOR2_X1   g0434(.A1(new_n375), .A2(new_n441), .ZN(new_n635));
  NAND3_X1  g0435(.A1(new_n573), .A2(new_n574), .A3(new_n469), .ZN(new_n636));
  INV_X1    g0436(.A(new_n496), .ZN(new_n637));
  OAI211_X1 g0437(.A(new_n636), .B(new_n637), .C1(G169), .C2(new_n576), .ZN(new_n638));
  AND3_X1   g0438(.A1(new_n524), .A2(new_n526), .A3(new_n528), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  NAND4_X1  g0440(.A1(new_n640), .A2(new_n578), .A3(new_n619), .A4(new_n632), .ZN(new_n641));
  INV_X1    g0441(.A(new_n592), .ZN(new_n642));
  AOI21_X1  g0442(.A(new_n642), .B1(new_n620), .B2(new_n621), .ZN(new_n643));
  INV_X1    g0443(.A(KEYINPUT26), .ZN(new_n644));
  AND2_X1   g0444(.A1(new_n562), .A2(new_n569), .ZN(new_n645));
  NAND3_X1  g0445(.A1(new_n643), .A2(new_n644), .A3(new_n645), .ZN(new_n646));
  NAND3_X1  g0446(.A1(new_n645), .A2(new_n622), .A3(new_n631), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n647), .A2(KEYINPUT26), .ZN(new_n648));
  NAND4_X1  g0448(.A1(new_n641), .A2(new_n569), .A3(new_n646), .A4(new_n648), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n635), .A2(new_n649), .ZN(new_n650));
  INV_X1    g0450(.A(new_n374), .ZN(new_n651));
  AOI22_X1  g0451(.A1(new_n353), .A2(new_n651), .B1(new_n329), .B2(new_n346), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n436), .A2(new_n437), .ZN(new_n653));
  OAI21_X1  g0453(.A(new_n427), .B1(new_n652), .B2(new_n653), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n303), .A2(new_n304), .ZN(new_n655));
  AOI21_X1  g0455(.A(new_n296), .B1(new_n654), .B2(new_n655), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n650), .A2(new_n656), .ZN(G369));
  NOR2_X1   g0457(.A1(new_n252), .A2(G20), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n658), .A2(new_n281), .ZN(new_n659));
  OR2_X1    g0459(.A1(new_n659), .A2(KEYINPUT27), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n659), .A2(KEYINPUT27), .ZN(new_n661));
  NAND3_X1  g0461(.A1(new_n660), .A2(G213), .A3(new_n661), .ZN(new_n662));
  INV_X1    g0462(.A(G343), .ZN(new_n663));
  NOR2_X1   g0463(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  NOR2_X1   g0464(.A1(new_n638), .A2(new_n664), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n636), .A2(new_n664), .ZN(new_n666));
  XNOR2_X1  g0466(.A(new_n666), .B(KEYINPUT89), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n575), .A2(new_n577), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  AOI21_X1  g0469(.A(new_n665), .B1(new_n669), .B2(new_n638), .ZN(new_n670));
  NOR2_X1   g0470(.A1(new_n639), .A2(new_n664), .ZN(new_n671));
  AND2_X1   g0471(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  NOR2_X1   g0472(.A1(new_n672), .A2(new_n665), .ZN(new_n673));
  INV_X1    g0473(.A(new_n664), .ZN(new_n674));
  NOR2_X1   g0474(.A1(new_n520), .A2(new_n674), .ZN(new_n675));
  INV_X1    g0475(.A(new_n675), .ZN(new_n676));
  NAND3_X1  g0476(.A1(new_n639), .A2(new_n521), .A3(new_n676), .ZN(new_n677));
  OAI21_X1  g0477(.A(new_n677), .B1(new_n639), .B2(new_n676), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n678), .A2(G330), .ZN(new_n679));
  INV_X1    g0479(.A(new_n679), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n670), .A2(new_n680), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n673), .A2(new_n681), .ZN(G399));
  NOR2_X1   g0482(.A1(new_n226), .A2(G41), .ZN(new_n683));
  INV_X1    g0483(.A(new_n683), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n684), .A2(G1), .ZN(new_n685));
  OR3_X1    g0485(.A1(new_n536), .A2(new_n539), .A3(G116), .ZN(new_n686));
  INV_X1    g0486(.A(new_n233), .ZN(new_n687));
  OAI22_X1  g0487(.A1(new_n685), .A2(new_n686), .B1(new_n687), .B2(new_n684), .ZN(new_n688));
  XNOR2_X1  g0488(.A(new_n688), .B(KEYINPUT28), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n649), .A2(new_n674), .ZN(new_n690));
  INV_X1    g0490(.A(KEYINPUT90), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  INV_X1    g0492(.A(KEYINPUT29), .ZN(new_n693));
  NAND3_X1  g0493(.A1(new_n649), .A2(KEYINPUT90), .A3(new_n674), .ZN(new_n694));
  NAND3_X1  g0494(.A1(new_n692), .A2(new_n693), .A3(new_n694), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n695), .A2(KEYINPUT91), .ZN(new_n696));
  NAND2_X1  g0496(.A1(new_n647), .A2(new_n644), .ZN(new_n697));
  INV_X1    g0497(.A(KEYINPUT92), .ZN(new_n698));
  NAND4_X1  g0498(.A1(new_n645), .A2(new_n622), .A3(KEYINPUT26), .A4(new_n592), .ZN(new_n699));
  NAND3_X1  g0499(.A1(new_n697), .A2(new_n698), .A3(new_n699), .ZN(new_n700));
  OR2_X1    g0500(.A1(new_n699), .A2(new_n698), .ZN(new_n701));
  NAND3_X1  g0501(.A1(new_n700), .A2(new_n569), .A3(new_n701), .ZN(new_n702));
  INV_X1    g0502(.A(KEYINPUT93), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  NAND4_X1  g0504(.A1(new_n700), .A2(new_n701), .A3(KEYINPUT93), .A4(new_n569), .ZN(new_n705));
  NAND3_X1  g0505(.A1(new_n704), .A2(new_n641), .A3(new_n705), .ZN(new_n706));
  NAND3_X1  g0506(.A1(new_n706), .A2(KEYINPUT29), .A3(new_n674), .ZN(new_n707));
  INV_X1    g0507(.A(KEYINPUT91), .ZN(new_n708));
  NAND4_X1  g0508(.A1(new_n692), .A2(new_n708), .A3(new_n693), .A4(new_n694), .ZN(new_n709));
  NAND3_X1  g0509(.A1(new_n696), .A2(new_n707), .A3(new_n709), .ZN(new_n710));
  NOR2_X1   g0510(.A1(new_n527), .A2(new_n292), .ZN(new_n711));
  NAND2_X1  g0511(.A1(new_n477), .A2(new_n492), .ZN(new_n712));
  NOR2_X1   g0512(.A1(new_n712), .A2(new_n557), .ZN(new_n713));
  NAND3_X1  g0513(.A1(new_n607), .A2(new_n711), .A3(new_n713), .ZN(new_n714));
  INV_X1    g0514(.A(KEYINPUT30), .ZN(new_n715));
  NAND2_X1  g0515(.A1(new_n714), .A2(new_n715), .ZN(new_n716));
  NOR2_X1   g0516(.A1(new_n525), .A2(G179), .ZN(new_n717));
  NAND4_X1  g0517(.A1(new_n617), .A2(new_n717), .A3(new_n493), .A4(new_n557), .ZN(new_n718));
  NAND4_X1  g0518(.A1(new_n607), .A2(KEYINPUT30), .A3(new_n711), .A4(new_n713), .ZN(new_n719));
  NAND3_X1  g0519(.A1(new_n716), .A2(new_n718), .A3(new_n719), .ZN(new_n720));
  NAND2_X1  g0520(.A1(new_n720), .A2(new_n664), .ZN(new_n721));
  OAI211_X1 g0521(.A(KEYINPUT31), .B(new_n721), .C1(new_n633), .C2(new_n664), .ZN(new_n722));
  INV_X1    g0522(.A(KEYINPUT31), .ZN(new_n723));
  NAND3_X1  g0523(.A1(new_n720), .A2(new_n723), .A3(new_n664), .ZN(new_n724));
  NAND2_X1  g0524(.A1(new_n722), .A2(new_n724), .ZN(new_n725));
  INV_X1    g0525(.A(G330), .ZN(new_n726));
  NOR2_X1   g0526(.A1(new_n725), .A2(new_n726), .ZN(new_n727));
  INV_X1    g0527(.A(new_n727), .ZN(new_n728));
  NAND2_X1  g0528(.A1(new_n710), .A2(new_n728), .ZN(new_n729));
  INV_X1    g0529(.A(new_n729), .ZN(new_n730));
  OAI21_X1  g0530(.A(new_n689), .B1(new_n730), .B2(G1), .ZN(G364));
  AOI21_X1  g0531(.A(new_n685), .B1(G45), .B2(new_n658), .ZN(new_n732));
  NOR2_X1   g0532(.A1(new_n680), .A2(new_n732), .ZN(new_n733));
  OAI21_X1  g0533(.A(new_n733), .B1(G330), .B2(new_n678), .ZN(new_n734));
  NOR2_X1   g0534(.A1(new_n230), .A2(G190), .ZN(new_n735));
  NOR2_X1   g0535(.A1(new_n292), .A2(G200), .ZN(new_n736));
  AND2_X1   g0536(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  INV_X1    g0537(.A(new_n737), .ZN(new_n738));
  NAND3_X1  g0538(.A1(G20), .A2(G179), .A3(G200), .ZN(new_n739));
  NOR2_X1   g0539(.A1(new_n739), .A2(new_n348), .ZN(new_n740));
  INV_X1    g0540(.A(new_n740), .ZN(new_n741));
  OAI22_X1  g0541(.A1(new_n738), .A2(new_n340), .B1(new_n201), .B2(new_n741), .ZN(new_n742));
  NOR2_X1   g0542(.A1(new_n230), .A2(new_n348), .ZN(new_n743));
  NAND2_X1  g0543(.A1(new_n743), .A2(new_n736), .ZN(new_n744));
  INV_X1    g0544(.A(new_n744), .ZN(new_n745));
  AOI21_X1  g0545(.A(new_n742), .B1(G58), .B2(new_n745), .ZN(new_n746));
  XNOR2_X1  g0546(.A(new_n746), .B(KEYINPUT95), .ZN(new_n747));
  NOR2_X1   g0547(.A1(new_n739), .A2(G190), .ZN(new_n748));
  INV_X1    g0548(.A(new_n748), .ZN(new_n749));
  NOR2_X1   g0549(.A1(G179), .A2(G200), .ZN(new_n750));
  AOI21_X1  g0550(.A(new_n230), .B1(new_n750), .B2(G190), .ZN(new_n751));
  OAI22_X1  g0551(.A1(new_n749), .A2(new_n203), .B1(new_n751), .B2(new_n541), .ZN(new_n752));
  NOR2_X1   g0552(.A1(new_n439), .A2(G179), .ZN(new_n753));
  NAND2_X1  g0553(.A1(new_n735), .A2(new_n753), .ZN(new_n754));
  NAND2_X1  g0554(.A1(new_n743), .A2(new_n753), .ZN(new_n755));
  OAI221_X1 g0555(.A(new_n274), .B1(new_n754), .B2(new_n214), .C1(new_n209), .C2(new_n755), .ZN(new_n756));
  OR3_X1    g0556(.A1(new_n747), .A2(new_n752), .A3(new_n756), .ZN(new_n757));
  NAND2_X1  g0557(.A1(new_n735), .A2(new_n750), .ZN(new_n758));
  INV_X1    g0558(.A(new_n758), .ZN(new_n759));
  NAND2_X1  g0559(.A1(new_n759), .A2(G159), .ZN(new_n760));
  XNOR2_X1  g0560(.A(new_n760), .B(KEYINPUT32), .ZN(new_n761));
  AND2_X1   g0561(.A1(new_n737), .A2(G311), .ZN(new_n762));
  INV_X1    g0562(.A(G322), .ZN(new_n763));
  OAI21_X1  g0563(.A(new_n312), .B1(new_n744), .B2(new_n763), .ZN(new_n764));
  XNOR2_X1  g0564(.A(KEYINPUT96), .B(G326), .ZN(new_n765));
  OAI22_X1  g0565(.A1(new_n741), .A2(new_n765), .B1(new_n475), .B2(new_n751), .ZN(new_n766));
  INV_X1    g0566(.A(new_n755), .ZN(new_n767));
  AOI211_X1 g0567(.A(new_n764), .B(new_n766), .C1(G303), .C2(new_n767), .ZN(new_n768));
  INV_X1    g0568(.A(new_n754), .ZN(new_n769));
  AOI22_X1  g0569(.A1(G283), .A2(new_n769), .B1(new_n759), .B2(G329), .ZN(new_n770));
  XOR2_X1   g0570(.A(new_n770), .B(KEYINPUT97), .Z(new_n771));
  XNOR2_X1  g0571(.A(KEYINPUT98), .B(G317), .ZN(new_n772));
  XOR2_X1   g0572(.A(new_n772), .B(KEYINPUT33), .Z(new_n773));
  OAI211_X1 g0573(.A(new_n768), .B(new_n771), .C1(new_n749), .C2(new_n773), .ZN(new_n774));
  OAI22_X1  g0574(.A1(new_n757), .A2(new_n761), .B1(new_n762), .B2(new_n774), .ZN(new_n775));
  OAI211_X1 g0575(.A(G1), .B(G13), .C1(new_n230), .C2(G169), .ZN(new_n776));
  XOR2_X1   g0576(.A(new_n776), .B(KEYINPUT94), .Z(new_n777));
  INV_X1    g0577(.A(new_n777), .ZN(new_n778));
  NOR2_X1   g0578(.A1(G13), .A2(G33), .ZN(new_n779));
  INV_X1    g0579(.A(new_n779), .ZN(new_n780));
  NOR2_X1   g0580(.A1(new_n780), .A2(G20), .ZN(new_n781));
  NOR2_X1   g0581(.A1(new_n778), .A2(new_n781), .ZN(new_n782));
  NAND3_X1  g0582(.A1(new_n274), .A2(G355), .A3(new_n225), .ZN(new_n783));
  NOR2_X1   g0583(.A1(new_n552), .A2(new_n226), .ZN(new_n784));
  OAI21_X1  g0584(.A(new_n784), .B1(new_n687), .B2(G45), .ZN(new_n785));
  NOR2_X1   g0585(.A1(new_n247), .A2(new_n286), .ZN(new_n786));
  OAI221_X1 g0586(.A(new_n783), .B1(G116), .B2(new_n225), .C1(new_n785), .C2(new_n786), .ZN(new_n787));
  AOI22_X1  g0587(.A1(new_n775), .A2(new_n778), .B1(new_n782), .B2(new_n787), .ZN(new_n788));
  INV_X1    g0588(.A(new_n781), .ZN(new_n789));
  OAI211_X1 g0589(.A(new_n788), .B(new_n732), .C1(new_n678), .C2(new_n789), .ZN(new_n790));
  AND2_X1   g0590(.A1(new_n734), .A2(new_n790), .ZN(new_n791));
  INV_X1    g0591(.A(new_n791), .ZN(G396));
  OR2_X1    g0592(.A1(new_n372), .A2(new_n674), .ZN(new_n793));
  NAND2_X1  g0593(.A1(new_n440), .A2(new_n793), .ZN(new_n794));
  NAND2_X1  g0594(.A1(new_n794), .A2(new_n374), .ZN(new_n795));
  NAND2_X1  g0595(.A1(new_n651), .A2(new_n674), .ZN(new_n796));
  INV_X1    g0596(.A(KEYINPUT99), .ZN(new_n797));
  NAND3_X1  g0597(.A1(new_n795), .A2(new_n796), .A3(new_n797), .ZN(new_n798));
  AOI22_X1  g0598(.A1(new_n440), .A2(new_n793), .B1(new_n373), .B2(new_n363), .ZN(new_n799));
  NOR2_X1   g0599(.A1(new_n374), .A2(new_n664), .ZN(new_n800));
  OAI21_X1  g0600(.A(KEYINPUT99), .B1(new_n799), .B2(new_n800), .ZN(new_n801));
  NAND2_X1  g0601(.A1(new_n798), .A2(new_n801), .ZN(new_n802));
  INV_X1    g0602(.A(new_n802), .ZN(new_n803));
  NAND3_X1  g0603(.A1(new_n692), .A2(new_n694), .A3(new_n803), .ZN(new_n804));
  NAND3_X1  g0604(.A1(new_n649), .A2(new_n802), .A3(new_n674), .ZN(new_n805));
  NAND2_X1  g0605(.A1(new_n804), .A2(new_n805), .ZN(new_n806));
  XNOR2_X1  g0606(.A(new_n806), .B(new_n727), .ZN(new_n807));
  INV_X1    g0607(.A(new_n732), .ZN(new_n808));
  NAND2_X1  g0608(.A1(new_n807), .A2(new_n808), .ZN(new_n809));
  AOI22_X1  g0609(.A1(new_n745), .A2(G143), .B1(G150), .B2(new_n748), .ZN(new_n810));
  INV_X1    g0610(.A(G137), .ZN(new_n811));
  INV_X1    g0611(.A(G159), .ZN(new_n812));
  OAI221_X1 g0612(.A(new_n810), .B1(new_n811), .B2(new_n741), .C1(new_n812), .C2(new_n738), .ZN(new_n813));
  XNOR2_X1  g0613(.A(new_n813), .B(KEYINPUT34), .ZN(new_n814));
  NAND2_X1  g0614(.A1(new_n769), .A2(G68), .ZN(new_n815));
  INV_X1    g0615(.A(G132), .ZN(new_n816));
  OAI22_X1  g0616(.A1(new_n755), .A2(new_n201), .B1(new_n758), .B2(new_n816), .ZN(new_n817));
  INV_X1    g0617(.A(new_n751), .ZN(new_n818));
  AOI211_X1 g0618(.A(new_n383), .B(new_n817), .C1(G58), .C2(new_n818), .ZN(new_n819));
  NAND3_X1  g0619(.A1(new_n814), .A2(new_n815), .A3(new_n819), .ZN(new_n820));
  NOR2_X1   g0620(.A1(new_n754), .A2(new_n209), .ZN(new_n821));
  OAI22_X1  g0621(.A1(new_n738), .A2(new_n444), .B1(new_n755), .B2(new_n214), .ZN(new_n822));
  AOI211_X1 g0622(.A(new_n821), .B(new_n822), .C1(G311), .C2(new_n759), .ZN(new_n823));
  INV_X1    g0623(.A(G283), .ZN(new_n824));
  INV_X1    g0624(.A(G303), .ZN(new_n825));
  OAI22_X1  g0625(.A1(new_n749), .A2(new_n824), .B1(new_n741), .B2(new_n825), .ZN(new_n826));
  AOI211_X1 g0626(.A(new_n274), .B(new_n826), .C1(G294), .C2(new_n745), .ZN(new_n827));
  OAI211_X1 g0627(.A(new_n823), .B(new_n827), .C1(new_n541), .C2(new_n751), .ZN(new_n828));
  AOI21_X1  g0628(.A(new_n777), .B1(new_n820), .B2(new_n828), .ZN(new_n829));
  NOR2_X1   g0629(.A1(new_n778), .A2(new_n779), .ZN(new_n830));
  AOI21_X1  g0630(.A(new_n829), .B1(new_n340), .B2(new_n830), .ZN(new_n831));
  OAI211_X1 g0631(.A(new_n732), .B(new_n831), .C1(new_n802), .C2(new_n780), .ZN(new_n832));
  NAND2_X1  g0632(.A1(new_n809), .A2(new_n832), .ZN(G384));
  NOR2_X1   g0633(.A1(new_n347), .A2(new_n664), .ZN(new_n834));
  INV_X1    g0634(.A(KEYINPUT102), .ZN(new_n835));
  NAND3_X1  g0635(.A1(new_n427), .A2(new_n436), .A3(new_n437), .ZN(new_n836));
  INV_X1    g0636(.A(new_n662), .ZN(new_n837));
  AOI21_X1  g0637(.A(KEYINPUT16), .B1(new_n390), .B2(new_n392), .ZN(new_n838));
  OAI21_X1  g0638(.A(new_n418), .B1(new_n423), .B2(new_n838), .ZN(new_n839));
  NAND3_X1  g0639(.A1(new_n836), .A2(new_n837), .A3(new_n839), .ZN(new_n840));
  NAND3_X1  g0640(.A1(new_n406), .A2(new_n434), .A3(new_n428), .ZN(new_n841));
  NAND3_X1  g0641(.A1(new_n414), .A2(new_n415), .A3(new_n662), .ZN(new_n842));
  NAND2_X1  g0642(.A1(new_n839), .A2(new_n842), .ZN(new_n843));
  NAND2_X1  g0643(.A1(new_n841), .A2(new_n843), .ZN(new_n844));
  NAND2_X1  g0644(.A1(new_n844), .A2(KEYINPUT37), .ZN(new_n845));
  NAND2_X1  g0645(.A1(new_n424), .A2(new_n842), .ZN(new_n846));
  NAND2_X1  g0646(.A1(new_n841), .A2(new_n846), .ZN(new_n847));
  OAI21_X1  g0647(.A(new_n845), .B1(KEYINPUT37), .B2(new_n847), .ZN(new_n848));
  AND3_X1   g0648(.A1(new_n840), .A2(KEYINPUT38), .A3(new_n848), .ZN(new_n849));
  AOI21_X1  g0649(.A(KEYINPUT38), .B1(new_n840), .B2(new_n848), .ZN(new_n850));
  OAI21_X1  g0650(.A(KEYINPUT39), .B1(new_n849), .B2(new_n850), .ZN(new_n851));
  NAND3_X1  g0651(.A1(new_n836), .A2(new_n424), .A3(new_n837), .ZN(new_n852));
  XNOR2_X1  g0652(.A(new_n847), .B(KEYINPUT37), .ZN(new_n853));
  NAND2_X1  g0653(.A1(new_n852), .A2(new_n853), .ZN(new_n854));
  INV_X1    g0654(.A(KEYINPUT38), .ZN(new_n855));
  NAND2_X1  g0655(.A1(new_n854), .A2(new_n855), .ZN(new_n856));
  INV_X1    g0656(.A(KEYINPUT39), .ZN(new_n857));
  NAND3_X1  g0657(.A1(new_n840), .A2(KEYINPUT38), .A3(new_n848), .ZN(new_n858));
  NAND3_X1  g0658(.A1(new_n856), .A2(new_n857), .A3(new_n858), .ZN(new_n859));
  AOI21_X1  g0659(.A(new_n835), .B1(new_n851), .B2(new_n859), .ZN(new_n860));
  AOI21_X1  g0660(.A(KEYINPUT38), .B1(new_n852), .B2(new_n853), .ZN(new_n861));
  NOR3_X1   g0661(.A1(new_n849), .A2(new_n861), .A3(KEYINPUT39), .ZN(new_n862));
  NOR2_X1   g0662(.A1(new_n862), .A2(KEYINPUT102), .ZN(new_n863));
  OAI21_X1  g0663(.A(new_n834), .B1(new_n860), .B2(new_n863), .ZN(new_n864));
  NAND2_X1  g0664(.A1(new_n346), .A2(new_n664), .ZN(new_n865));
  NAND3_X1  g0665(.A1(new_n353), .A2(new_n347), .A3(new_n865), .ZN(new_n866));
  OAI211_X1 g0666(.A(new_n346), .B(new_n664), .C1(new_n352), .C2(new_n329), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n866), .A2(new_n867), .ZN(new_n868));
  INV_X1    g0668(.A(new_n868), .ZN(new_n869));
  AOI21_X1  g0669(.A(new_n869), .B1(new_n796), .B2(new_n805), .ZN(new_n870));
  OAI21_X1  g0670(.A(new_n870), .B1(new_n850), .B2(new_n849), .ZN(new_n871));
  NAND3_X1  g0671(.A1(new_n417), .A2(new_n426), .A3(new_n662), .ZN(new_n872));
  NAND3_X1  g0672(.A1(new_n864), .A2(new_n871), .A3(new_n872), .ZN(new_n873));
  NAND4_X1  g0673(.A1(new_n696), .A2(new_n635), .A3(new_n707), .A4(new_n709), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n874), .A2(new_n656), .ZN(new_n875));
  XNOR2_X1  g0675(.A(new_n873), .B(new_n875), .ZN(new_n876));
  INV_X1    g0676(.A(KEYINPUT40), .ZN(new_n877));
  NOR2_X1   g0677(.A1(new_n869), .A2(new_n803), .ZN(new_n878));
  INV_X1    g0678(.A(KEYINPUT103), .ZN(new_n879));
  AND3_X1   g0679(.A1(new_n722), .A2(new_n879), .A3(new_n724), .ZN(new_n880));
  AOI21_X1  g0680(.A(new_n879), .B1(new_n722), .B2(new_n724), .ZN(new_n881));
  OAI21_X1  g0681(.A(new_n878), .B1(new_n880), .B2(new_n881), .ZN(new_n882));
  NOR2_X1   g0682(.A1(new_n849), .A2(new_n850), .ZN(new_n883));
  OAI21_X1  g0683(.A(new_n877), .B1(new_n882), .B2(new_n883), .ZN(new_n884));
  AOI21_X1  g0684(.A(new_n877), .B1(new_n856), .B2(new_n858), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n725), .A2(KEYINPUT103), .ZN(new_n886));
  NAND3_X1  g0686(.A1(new_n722), .A2(new_n879), .A3(new_n724), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n886), .A2(new_n887), .ZN(new_n888));
  NAND3_X1  g0688(.A1(new_n885), .A2(new_n888), .A3(new_n878), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n884), .A2(new_n889), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n888), .A2(new_n635), .ZN(new_n891));
  XNOR2_X1  g0691(.A(new_n890), .B(new_n891), .ZN(new_n892));
  NOR2_X1   g0692(.A1(new_n892), .A2(new_n726), .ZN(new_n893));
  XNOR2_X1  g0693(.A(new_n876), .B(new_n893), .ZN(new_n894));
  OAI21_X1  g0694(.A(new_n894), .B1(new_n281), .B2(new_n658), .ZN(new_n895));
  OAI211_X1 g0695(.A(new_n233), .B(G77), .C1(new_n202), .C2(new_n203), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n201), .A2(G68), .ZN(new_n897));
  AOI211_X1 g0697(.A(new_n281), .B(G13), .C1(new_n896), .C2(new_n897), .ZN(new_n898));
  XNOR2_X1  g0698(.A(new_n898), .B(KEYINPUT101), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n587), .A2(new_n588), .ZN(new_n900));
  AOI21_X1  g0700(.A(new_n444), .B1(new_n900), .B2(KEYINPUT35), .ZN(new_n901));
  OAI211_X1 g0701(.A(new_n901), .B(new_n231), .C1(KEYINPUT35), .C2(new_n900), .ZN(new_n902));
  XOR2_X1   g0702(.A(KEYINPUT100), .B(KEYINPUT36), .Z(new_n903));
  XNOR2_X1  g0703(.A(new_n902), .B(new_n903), .ZN(new_n904));
  NAND3_X1  g0704(.A1(new_n895), .A2(new_n899), .A3(new_n904), .ZN(G367));
  OAI211_X1 g0705(.A(new_n619), .B(new_n632), .C1(new_n642), .C2(new_n674), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n643), .A2(new_n664), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n672), .A2(new_n908), .ZN(new_n909));
  INV_X1    g0709(.A(KEYINPUT42), .ZN(new_n910));
  XNOR2_X1  g0710(.A(new_n909), .B(new_n910), .ZN(new_n911));
  INV_X1    g0711(.A(new_n908), .ZN(new_n912));
  OAI21_X1  g0712(.A(new_n632), .B1(new_n912), .B2(new_n638), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n913), .A2(new_n674), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n911), .A2(new_n914), .ZN(new_n915));
  INV_X1    g0715(.A(KEYINPUT104), .ZN(new_n916));
  XNOR2_X1  g0716(.A(new_n915), .B(new_n916), .ZN(new_n917));
  OR2_X1    g0717(.A1(new_n544), .A2(new_n674), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n645), .A2(new_n918), .ZN(new_n919));
  OAI21_X1  g0719(.A(new_n919), .B1(new_n569), .B2(new_n918), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n920), .A2(KEYINPUT43), .ZN(new_n921));
  OR2_X1    g0721(.A1(new_n920), .A2(KEYINPUT43), .ZN(new_n922));
  NAND3_X1  g0722(.A1(new_n917), .A2(new_n921), .A3(new_n922), .ZN(new_n923));
  OAI21_X1  g0723(.A(new_n923), .B1(new_n917), .B2(new_n922), .ZN(new_n924));
  NOR2_X1   g0724(.A1(new_n681), .A2(new_n912), .ZN(new_n925));
  INV_X1    g0725(.A(new_n925), .ZN(new_n926));
  NAND2_X1  g0726(.A1(new_n924), .A2(new_n926), .ZN(new_n927));
  OAI211_X1 g0727(.A(new_n923), .B(new_n925), .C1(new_n917), .C2(new_n922), .ZN(new_n928));
  XNOR2_X1  g0728(.A(new_n683), .B(KEYINPUT41), .ZN(new_n929));
  INV_X1    g0729(.A(new_n929), .ZN(new_n930));
  XNOR2_X1  g0730(.A(new_n670), .B(new_n671), .ZN(new_n931));
  XNOR2_X1  g0731(.A(new_n931), .B(new_n680), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n730), .A2(new_n932), .ZN(new_n933));
  OR2_X1    g0733(.A1(new_n933), .A2(KEYINPUT105), .ZN(new_n934));
  NOR2_X1   g0734(.A1(new_n673), .A2(new_n908), .ZN(new_n935));
  NOR2_X1   g0735(.A1(new_n935), .A2(KEYINPUT44), .ZN(new_n936));
  INV_X1    g0736(.A(KEYINPUT44), .ZN(new_n937));
  NOR3_X1   g0737(.A1(new_n673), .A2(new_n937), .A3(new_n908), .ZN(new_n938));
  AND3_X1   g0738(.A1(new_n673), .A2(KEYINPUT45), .A3(new_n908), .ZN(new_n939));
  AOI21_X1  g0739(.A(KEYINPUT45), .B1(new_n673), .B2(new_n908), .ZN(new_n940));
  OAI22_X1  g0740(.A1(new_n936), .A2(new_n938), .B1(new_n939), .B2(new_n940), .ZN(new_n941));
  NAND3_X1  g0741(.A1(new_n941), .A2(KEYINPUT106), .A3(new_n681), .ZN(new_n942));
  XNOR2_X1  g0742(.A(new_n935), .B(KEYINPUT44), .ZN(new_n943));
  OR2_X1    g0743(.A1(new_n939), .A2(new_n940), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n681), .A2(KEYINPUT106), .ZN(new_n945));
  OR2_X1    g0745(.A1(new_n681), .A2(KEYINPUT106), .ZN(new_n946));
  NAND4_X1  g0746(.A1(new_n943), .A2(new_n944), .A3(new_n945), .A4(new_n946), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n942), .A2(new_n947), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n933), .A2(KEYINPUT105), .ZN(new_n949));
  NAND3_X1  g0749(.A1(new_n934), .A2(new_n948), .A3(new_n949), .ZN(new_n950));
  AOI21_X1  g0750(.A(new_n930), .B1(new_n950), .B2(new_n730), .ZN(new_n951));
  AOI21_X1  g0751(.A(new_n281), .B1(new_n658), .B2(G45), .ZN(new_n952));
  INV_X1    g0752(.A(new_n952), .ZN(new_n953));
  OAI211_X1 g0753(.A(new_n927), .B(new_n928), .C1(new_n951), .C2(new_n953), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n769), .A2(G77), .ZN(new_n955));
  OAI221_X1 g0755(.A(new_n955), .B1(new_n267), .B2(new_n744), .C1(new_n201), .C2(new_n738), .ZN(new_n956));
  AOI21_X1  g0756(.A(new_n956), .B1(G137), .B2(new_n759), .ZN(new_n957));
  NOR2_X1   g0757(.A1(new_n751), .A2(new_n203), .ZN(new_n958));
  OAI21_X1  g0758(.A(new_n274), .B1(new_n749), .B2(new_n812), .ZN(new_n959));
  AOI211_X1 g0759(.A(new_n958), .B(new_n959), .C1(G143), .C2(new_n740), .ZN(new_n960));
  OAI211_X1 g0760(.A(new_n957), .B(new_n960), .C1(new_n202), .C2(new_n755), .ZN(new_n961));
  XNOR2_X1  g0761(.A(KEYINPUT107), .B(G311), .ZN(new_n962));
  OAI22_X1  g0762(.A1(new_n475), .A2(new_n749), .B1(new_n741), .B2(new_n962), .ZN(new_n963));
  NAND2_X1  g0763(.A1(new_n767), .A2(G116), .ZN(new_n964));
  INV_X1    g0764(.A(KEYINPUT46), .ZN(new_n965));
  NOR2_X1   g0765(.A1(new_n964), .A2(new_n965), .ZN(new_n966));
  AOI211_X1 g0766(.A(new_n963), .B(new_n966), .C1(G107), .C2(new_n818), .ZN(new_n967));
  AOI21_X1  g0767(.A(new_n552), .B1(new_n964), .B2(new_n965), .ZN(new_n968));
  NOR2_X1   g0768(.A1(new_n754), .A2(new_n541), .ZN(new_n969));
  INV_X1    g0769(.A(new_n503), .ZN(new_n970));
  NOR2_X1   g0770(.A1(new_n970), .A2(new_n744), .ZN(new_n971));
  AOI211_X1 g0771(.A(new_n969), .B(new_n971), .C1(G283), .C2(new_n737), .ZN(new_n972));
  NAND3_X1  g0772(.A1(new_n967), .A2(new_n968), .A3(new_n972), .ZN(new_n973));
  INV_X1    g0773(.A(G317), .ZN(new_n974));
  NOR2_X1   g0774(.A1(new_n758), .A2(new_n974), .ZN(new_n975));
  OAI21_X1  g0775(.A(new_n961), .B1(new_n973), .B2(new_n975), .ZN(new_n976));
  XNOR2_X1  g0776(.A(new_n976), .B(KEYINPUT47), .ZN(new_n977));
  AOI21_X1  g0777(.A(new_n808), .B1(new_n977), .B2(new_n778), .ZN(new_n978));
  INV_X1    g0778(.A(new_n784), .ZN(new_n979));
  OAI221_X1 g0779(.A(new_n782), .B1(new_n225), .B2(new_n370), .C1(new_n243), .C2(new_n979), .ZN(new_n980));
  OAI211_X1 g0780(.A(new_n978), .B(new_n980), .C1(new_n789), .C2(new_n920), .ZN(new_n981));
  NAND2_X1  g0781(.A1(new_n954), .A2(new_n981), .ZN(G387));
  OR2_X1    g0782(.A1(new_n730), .A2(new_n932), .ZN(new_n983));
  NAND3_X1  g0783(.A1(new_n983), .A2(new_n683), .A3(new_n933), .ZN(new_n984));
  OAI21_X1  g0784(.A(new_n383), .B1(new_n758), .B2(new_n765), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n818), .A2(G283), .ZN(new_n986));
  AOI22_X1  g0786(.A1(new_n737), .A2(new_n503), .B1(G322), .B2(new_n740), .ZN(new_n987));
  OAI221_X1 g0787(.A(new_n987), .B1(new_n974), .B2(new_n744), .C1(new_n749), .C2(new_n962), .ZN(new_n988));
  INV_X1    g0788(.A(KEYINPUT48), .ZN(new_n989));
  OAI221_X1 g0789(.A(new_n986), .B1(new_n475), .B2(new_n755), .C1(new_n988), .C2(new_n989), .ZN(new_n990));
  XOR2_X1   g0790(.A(new_n990), .B(KEYINPUT110), .Z(new_n991));
  AOI21_X1  g0791(.A(new_n991), .B1(new_n989), .B2(new_n988), .ZN(new_n992));
  AOI21_X1  g0792(.A(new_n985), .B1(new_n992), .B2(KEYINPUT49), .ZN(new_n993));
  OAI221_X1 g0793(.A(new_n993), .B1(KEYINPUT49), .B2(new_n992), .C1(new_n444), .C2(new_n754), .ZN(new_n994));
  NOR2_X1   g0794(.A1(new_n744), .A2(new_n201), .ZN(new_n995));
  AOI22_X1  g0795(.A1(G150), .A2(new_n759), .B1(new_n737), .B2(G68), .ZN(new_n996));
  NAND2_X1  g0796(.A1(new_n740), .A2(G159), .ZN(new_n997));
  INV_X1    g0797(.A(KEYINPUT109), .ZN(new_n998));
  OAI21_X1  g0798(.A(new_n996), .B1(new_n997), .B2(new_n998), .ZN(new_n999));
  AOI21_X1  g0799(.A(new_n999), .B1(new_n998), .B2(new_n997), .ZN(new_n1000));
  NOR2_X1   g0800(.A1(new_n755), .A2(new_n340), .ZN(new_n1001));
  NOR2_X1   g0801(.A1(new_n1001), .A2(new_n383), .ZN(new_n1002));
  NOR2_X1   g0802(.A1(new_n370), .A2(new_n751), .ZN(new_n1003));
  AOI211_X1 g0803(.A(new_n969), .B(new_n1003), .C1(new_n367), .C2(new_n748), .ZN(new_n1004));
  NAND3_X1  g0804(.A1(new_n1000), .A2(new_n1002), .A3(new_n1004), .ZN(new_n1005));
  OAI21_X1  g0805(.A(new_n994), .B1(new_n995), .B2(new_n1005), .ZN(new_n1006));
  OR3_X1    g0806(.A1(new_n268), .A2(KEYINPUT50), .A3(G50), .ZN(new_n1007));
  OAI21_X1  g0807(.A(KEYINPUT50), .B1(new_n268), .B2(G50), .ZN(new_n1008));
  NAND2_X1  g0808(.A1(G68), .A2(G77), .ZN(new_n1009));
  NAND4_X1  g0809(.A1(new_n1007), .A2(new_n1008), .A3(new_n286), .A4(new_n1009), .ZN(new_n1010));
  OAI21_X1  g0810(.A(new_n784), .B1(new_n1010), .B2(new_n686), .ZN(new_n1011));
  XNOR2_X1  g0811(.A(new_n1011), .B(KEYINPUT108), .ZN(new_n1012));
  OAI21_X1  g0812(.A(new_n1012), .B1(new_n286), .B2(new_n240), .ZN(new_n1013));
  NAND3_X1  g0813(.A1(new_n686), .A2(new_n225), .A3(new_n274), .ZN(new_n1014));
  OAI211_X1 g0814(.A(new_n1013), .B(new_n1014), .C1(G107), .C2(new_n225), .ZN(new_n1015));
  AOI22_X1  g0815(.A1(new_n1006), .A2(new_n778), .B1(new_n782), .B2(new_n1015), .ZN(new_n1016));
  OAI211_X1 g0816(.A(new_n1016), .B(new_n732), .C1(new_n670), .C2(new_n789), .ZN(new_n1017));
  INV_X1    g0817(.A(new_n1017), .ZN(new_n1018));
  AOI21_X1  g0818(.A(new_n1018), .B1(new_n953), .B2(new_n932), .ZN(new_n1019));
  NAND2_X1  g0819(.A1(new_n984), .A2(new_n1019), .ZN(new_n1020));
  NAND2_X1  g0820(.A1(new_n1020), .A2(KEYINPUT111), .ZN(new_n1021));
  INV_X1    g0821(.A(KEYINPUT111), .ZN(new_n1022));
  NAND3_X1  g0822(.A1(new_n984), .A2(new_n1019), .A3(new_n1022), .ZN(new_n1023));
  NAND2_X1  g0823(.A1(new_n1021), .A2(new_n1023), .ZN(G393));
  INV_X1    g0824(.A(new_n933), .ZN(new_n1025));
  OAI211_X1 g0825(.A(new_n950), .B(new_n683), .C1(new_n948), .C2(new_n1025), .ZN(new_n1026));
  NAND2_X1  g0826(.A1(new_n912), .A2(new_n781), .ZN(new_n1027));
  OAI221_X1 g0827(.A(new_n782), .B1(new_n541), .B2(new_n225), .C1(new_n250), .C2(new_n979), .ZN(new_n1028));
  NOR2_X1   g0828(.A1(new_n751), .A2(new_n340), .ZN(new_n1029));
  AOI21_X1  g0829(.A(new_n821), .B1(new_n367), .B2(new_n737), .ZN(new_n1030));
  OAI21_X1  g0830(.A(new_n1030), .B1(new_n203), .B2(new_n755), .ZN(new_n1031));
  AOI211_X1 g0831(.A(new_n1029), .B(new_n1031), .C1(G143), .C2(new_n759), .ZN(new_n1032));
  AOI21_X1  g0832(.A(new_n383), .B1(new_n748), .B2(G50), .ZN(new_n1033));
  OAI22_X1  g0833(.A1(new_n741), .A2(new_n267), .B1(new_n744), .B2(new_n812), .ZN(new_n1034));
  XNOR2_X1  g0834(.A(KEYINPUT112), .B(KEYINPUT51), .ZN(new_n1035));
  XNOR2_X1  g0835(.A(new_n1034), .B(new_n1035), .ZN(new_n1036));
  NAND3_X1  g0836(.A1(new_n1032), .A2(new_n1033), .A3(new_n1036), .ZN(new_n1037));
  NOR2_X1   g0837(.A1(new_n738), .A2(new_n475), .ZN(new_n1038));
  AOI22_X1  g0838(.A1(new_n745), .A2(G311), .B1(G317), .B2(new_n740), .ZN(new_n1039));
  XOR2_X1   g0839(.A(new_n1039), .B(KEYINPUT52), .Z(new_n1040));
  OAI22_X1  g0840(.A1(new_n970), .A2(new_n749), .B1(new_n444), .B2(new_n751), .ZN(new_n1041));
  AOI21_X1  g0841(.A(new_n274), .B1(new_n769), .B2(G107), .ZN(new_n1042));
  OAI221_X1 g0842(.A(new_n1042), .B1(new_n824), .B2(new_n755), .C1(new_n763), .C2(new_n758), .ZN(new_n1043));
  INV_X1    g0843(.A(KEYINPUT113), .ZN(new_n1044));
  AOI21_X1  g0844(.A(new_n1041), .B1(new_n1043), .B2(new_n1044), .ZN(new_n1045));
  OAI211_X1 g0845(.A(new_n1040), .B(new_n1045), .C1(new_n1044), .C2(new_n1043), .ZN(new_n1046));
  OAI21_X1  g0846(.A(new_n1037), .B1(new_n1038), .B2(new_n1046), .ZN(new_n1047));
  AOI21_X1  g0847(.A(new_n808), .B1(new_n1047), .B2(new_n778), .ZN(new_n1048));
  AND3_X1   g0848(.A1(new_n1027), .A2(new_n1028), .A3(new_n1048), .ZN(new_n1049));
  AOI21_X1  g0849(.A(new_n1049), .B1(new_n948), .B2(new_n953), .ZN(new_n1050));
  AND2_X1   g0850(.A1(new_n1026), .A2(new_n1050), .ZN(new_n1051));
  INV_X1    g0851(.A(new_n1051), .ZN(G390));
  OAI211_X1 g0852(.A(G330), .B(new_n635), .C1(new_n880), .C2(new_n881), .ZN(new_n1053));
  INV_X1    g0853(.A(KEYINPUT115), .ZN(new_n1054));
  NAND2_X1  g0854(.A1(new_n1053), .A2(new_n1054), .ZN(new_n1055));
  NAND4_X1  g0855(.A1(new_n888), .A2(KEYINPUT115), .A3(G330), .A4(new_n635), .ZN(new_n1056));
  NAND2_X1  g0856(.A1(new_n1055), .A2(new_n1056), .ZN(new_n1057));
  AND3_X1   g0857(.A1(new_n1057), .A2(new_n874), .A3(new_n656), .ZN(new_n1058));
  NAND2_X1  g0858(.A1(new_n802), .A2(G330), .ZN(new_n1059));
  INV_X1    g0859(.A(new_n1059), .ZN(new_n1060));
  OAI21_X1  g0860(.A(new_n1060), .B1(new_n880), .B2(new_n881), .ZN(new_n1061));
  NAND2_X1  g0861(.A1(new_n1061), .A2(new_n869), .ZN(new_n1062));
  NAND3_X1  g0862(.A1(new_n706), .A2(new_n674), .A3(new_n802), .ZN(new_n1063));
  NOR2_X1   g0863(.A1(new_n725), .A2(new_n1059), .ZN(new_n1064));
  NAND2_X1  g0864(.A1(new_n1064), .A2(new_n868), .ZN(new_n1065));
  NAND4_X1  g0865(.A1(new_n1062), .A2(new_n796), .A3(new_n1063), .A4(new_n1065), .ZN(new_n1066));
  OAI211_X1 g0866(.A(new_n868), .B(new_n1060), .C1(new_n880), .C2(new_n881), .ZN(new_n1067));
  OAI21_X1  g0867(.A(new_n869), .B1(new_n725), .B2(new_n1059), .ZN(new_n1068));
  NAND2_X1  g0868(.A1(new_n1067), .A2(new_n1068), .ZN(new_n1069));
  NAND2_X1  g0869(.A1(new_n805), .A2(new_n796), .ZN(new_n1070));
  AOI21_X1  g0870(.A(KEYINPUT116), .B1(new_n1069), .B2(new_n1070), .ZN(new_n1071));
  INV_X1    g0871(.A(KEYINPUT116), .ZN(new_n1072));
  INV_X1    g0872(.A(new_n1070), .ZN(new_n1073));
  AOI211_X1 g0873(.A(new_n1072), .B(new_n1073), .C1(new_n1067), .C2(new_n1068), .ZN(new_n1074));
  OAI21_X1  g0874(.A(new_n1066), .B1(new_n1071), .B2(new_n1074), .ZN(new_n1075));
  NAND2_X1  g0875(.A1(new_n840), .A2(new_n848), .ZN(new_n1076));
  NAND2_X1  g0876(.A1(new_n1076), .A2(new_n855), .ZN(new_n1077));
  AOI21_X1  g0877(.A(new_n857), .B1(new_n1077), .B2(new_n858), .ZN(new_n1078));
  OAI21_X1  g0878(.A(KEYINPUT102), .B1(new_n862), .B2(new_n1078), .ZN(new_n1079));
  NAND2_X1  g0879(.A1(new_n859), .A2(new_n835), .ZN(new_n1080));
  INV_X1    g0880(.A(KEYINPUT114), .ZN(new_n1081));
  OAI21_X1  g0881(.A(new_n1081), .B1(new_n870), .B2(new_n834), .ZN(new_n1082));
  NAND2_X1  g0882(.A1(new_n1070), .A2(new_n868), .ZN(new_n1083));
  INV_X1    g0883(.A(new_n834), .ZN(new_n1084));
  NAND3_X1  g0884(.A1(new_n1083), .A2(KEYINPUT114), .A3(new_n1084), .ZN(new_n1085));
  NAND4_X1  g0885(.A1(new_n1079), .A2(new_n1080), .A3(new_n1082), .A4(new_n1085), .ZN(new_n1086));
  NAND2_X1  g0886(.A1(new_n1063), .A2(new_n796), .ZN(new_n1087));
  NAND2_X1  g0887(.A1(new_n1087), .A2(new_n868), .ZN(new_n1088));
  AOI21_X1  g0888(.A(new_n834), .B1(new_n856), .B2(new_n858), .ZN(new_n1089));
  NAND2_X1  g0889(.A1(new_n1088), .A2(new_n1089), .ZN(new_n1090));
  INV_X1    g0890(.A(new_n1065), .ZN(new_n1091));
  AND3_X1   g0891(.A1(new_n1086), .A2(new_n1090), .A3(new_n1091), .ZN(new_n1092));
  INV_X1    g0892(.A(new_n1067), .ZN(new_n1093));
  AOI21_X1  g0893(.A(new_n1093), .B1(new_n1086), .B2(new_n1090), .ZN(new_n1094));
  OAI211_X1 g0894(.A(new_n1058), .B(new_n1075), .C1(new_n1092), .C2(new_n1094), .ZN(new_n1095));
  NAND2_X1  g0895(.A1(new_n1075), .A2(new_n1058), .ZN(new_n1096));
  NAND2_X1  g0896(.A1(new_n1086), .A2(new_n1090), .ZN(new_n1097));
  NAND2_X1  g0897(.A1(new_n1097), .A2(new_n1067), .ZN(new_n1098));
  NAND3_X1  g0898(.A1(new_n1086), .A2(new_n1090), .A3(new_n1091), .ZN(new_n1099));
  NAND3_X1  g0899(.A1(new_n1096), .A2(new_n1098), .A3(new_n1099), .ZN(new_n1100));
  NAND3_X1  g0900(.A1(new_n1095), .A2(new_n1100), .A3(new_n683), .ZN(new_n1101));
  NOR2_X1   g0901(.A1(new_n860), .A2(new_n863), .ZN(new_n1102));
  AND2_X1   g0902(.A1(new_n1085), .A2(new_n1082), .ZN(new_n1103));
  AOI22_X1  g0903(.A1(new_n1102), .A2(new_n1103), .B1(new_n1088), .B2(new_n1089), .ZN(new_n1104));
  OAI21_X1  g0904(.A(new_n1099), .B1(new_n1104), .B2(new_n1093), .ZN(new_n1105));
  NAND2_X1  g0905(.A1(new_n830), .A2(new_n268), .ZN(new_n1106));
  NAND2_X1  g0906(.A1(new_n740), .A2(G128), .ZN(new_n1107));
  OAI21_X1  g0907(.A(new_n1107), .B1(new_n749), .B2(new_n811), .ZN(new_n1108));
  NAND3_X1  g0908(.A1(new_n767), .A2(KEYINPUT53), .A3(G150), .ZN(new_n1109));
  INV_X1    g0909(.A(KEYINPUT53), .ZN(new_n1110));
  OAI21_X1  g0910(.A(new_n1110), .B1(new_n755), .B2(new_n267), .ZN(new_n1111));
  AOI21_X1  g0911(.A(new_n1108), .B1(new_n1109), .B2(new_n1111), .ZN(new_n1112));
  INV_X1    g0912(.A(G125), .ZN(new_n1113));
  OAI22_X1  g0913(.A1(new_n744), .A2(new_n816), .B1(new_n758), .B2(new_n1113), .ZN(new_n1114));
  XOR2_X1   g0914(.A(KEYINPUT54), .B(G143), .Z(new_n1115));
  AOI21_X1  g0915(.A(new_n1114), .B1(new_n737), .B2(new_n1115), .ZN(new_n1116));
  NAND2_X1  g0916(.A1(new_n769), .A2(G50), .ZN(new_n1117));
  AOI21_X1  g0917(.A(new_n312), .B1(new_n818), .B2(G159), .ZN(new_n1118));
  NAND4_X1  g0918(.A1(new_n1112), .A2(new_n1116), .A3(new_n1117), .A4(new_n1118), .ZN(new_n1119));
  OAI221_X1 g0919(.A(new_n815), .B1(new_n444), .B2(new_n744), .C1(new_n475), .C2(new_n758), .ZN(new_n1120));
  INV_X1    g0920(.A(KEYINPUT117), .ZN(new_n1121));
  OAI21_X1  g0921(.A(new_n312), .B1(new_n755), .B2(new_n209), .ZN(new_n1122));
  AOI21_X1  g0922(.A(new_n1120), .B1(new_n1121), .B2(new_n1122), .ZN(new_n1123));
  NOR2_X1   g0923(.A1(new_n741), .A2(new_n824), .ZN(new_n1124));
  AOI211_X1 g0924(.A(new_n1029), .B(new_n1124), .C1(G107), .C2(new_n748), .ZN(new_n1125));
  OAI211_X1 g0925(.A(new_n1123), .B(new_n1125), .C1(new_n1121), .C2(new_n1122), .ZN(new_n1126));
  NOR2_X1   g0926(.A1(new_n738), .A2(new_n541), .ZN(new_n1127));
  OAI21_X1  g0927(.A(new_n1119), .B1(new_n1126), .B2(new_n1127), .ZN(new_n1128));
  XOR2_X1   g0928(.A(new_n1128), .B(KEYINPUT118), .Z(new_n1129));
  OAI21_X1  g0929(.A(new_n732), .B1(new_n1129), .B2(new_n777), .ZN(new_n1130));
  AOI21_X1  g0930(.A(new_n1130), .B1(new_n1102), .B2(new_n779), .ZN(new_n1131));
  AOI22_X1  g0931(.A1(new_n1105), .A2(new_n953), .B1(new_n1106), .B2(new_n1131), .ZN(new_n1132));
  AOI21_X1  g0932(.A(KEYINPUT119), .B1(new_n1101), .B2(new_n1132), .ZN(new_n1133));
  INV_X1    g0933(.A(new_n1133), .ZN(new_n1134));
  NAND3_X1  g0934(.A1(new_n1101), .A2(KEYINPUT119), .A3(new_n1132), .ZN(new_n1135));
  NAND2_X1  g0935(.A1(new_n1134), .A2(new_n1135), .ZN(G378));
  NAND3_X1  g0936(.A1(new_n884), .A2(new_n889), .A3(G330), .ZN(new_n1137));
  XNOR2_X1  g0937(.A(KEYINPUT123), .B(KEYINPUT55), .ZN(new_n1138));
  INV_X1    g0938(.A(new_n1138), .ZN(new_n1139));
  XNOR2_X1  g0939(.A(new_n305), .B(new_n1139), .ZN(new_n1140));
  NAND2_X1  g0940(.A1(new_n273), .A2(new_n837), .ZN(new_n1141));
  XNOR2_X1  g0941(.A(new_n1141), .B(KEYINPUT56), .ZN(new_n1142));
  XOR2_X1   g0942(.A(KEYINPUT121), .B(KEYINPUT122), .Z(new_n1143));
  XNOR2_X1  g0943(.A(new_n1142), .B(new_n1143), .ZN(new_n1144));
  XNOR2_X1  g0944(.A(new_n1140), .B(new_n1144), .ZN(new_n1145));
  NAND2_X1  g0945(.A1(new_n1137), .A2(new_n1145), .ZN(new_n1146));
  INV_X1    g0946(.A(new_n1145), .ZN(new_n1147));
  NAND4_X1  g0947(.A1(new_n1147), .A2(new_n884), .A3(G330), .A4(new_n889), .ZN(new_n1148));
  NAND2_X1  g0948(.A1(new_n1146), .A2(new_n1148), .ZN(new_n1149));
  AND3_X1   g0949(.A1(new_n864), .A2(new_n871), .A3(new_n872), .ZN(new_n1150));
  NAND2_X1  g0950(.A1(new_n1149), .A2(new_n1150), .ZN(new_n1151));
  NAND3_X1  g0951(.A1(new_n873), .A2(new_n1148), .A3(new_n1146), .ZN(new_n1152));
  NAND2_X1  g0952(.A1(new_n1151), .A2(new_n1152), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n1153), .A2(new_n953), .ZN(new_n1154));
  AOI21_X1  g0954(.A(new_n808), .B1(new_n830), .B2(new_n201), .ZN(new_n1155));
  XNOR2_X1  g0955(.A(new_n1155), .B(KEYINPUT120), .ZN(new_n1156));
  NAND2_X1  g0956(.A1(new_n552), .A2(G33), .ZN(new_n1157));
  INV_X1    g0957(.A(new_n1157), .ZN(new_n1158));
  OAI21_X1  g0958(.A(new_n201), .B1(new_n1158), .B2(G41), .ZN(new_n1159));
  AOI22_X1  g0959(.A1(new_n818), .A2(G150), .B1(G125), .B2(new_n740), .ZN(new_n1160));
  INV_X1    g0960(.A(new_n1160), .ZN(new_n1161));
  AOI22_X1  g0961(.A1(G128), .A2(new_n745), .B1(new_n767), .B2(new_n1115), .ZN(new_n1162));
  OAI21_X1  g0962(.A(new_n1162), .B1(new_n811), .B2(new_n738), .ZN(new_n1163));
  AOI211_X1 g0963(.A(new_n1161), .B(new_n1163), .C1(G132), .C2(new_n748), .ZN(new_n1164));
  INV_X1    g0964(.A(KEYINPUT59), .ZN(new_n1165));
  OAI221_X1 g0965(.A(new_n262), .B1(new_n812), .B2(new_n754), .C1(new_n1164), .C2(new_n1165), .ZN(new_n1166));
  AOI21_X1  g0966(.A(G41), .B1(new_n759), .B2(G124), .ZN(new_n1167));
  INV_X1    g0967(.A(new_n1164), .ZN(new_n1168));
  OAI21_X1  g0968(.A(new_n1167), .B1(new_n1168), .B2(KEYINPUT59), .ZN(new_n1169));
  OAI21_X1  g0969(.A(new_n1159), .B1(new_n1166), .B2(new_n1169), .ZN(new_n1170));
  AOI22_X1  g0970(.A1(G107), .A2(new_n745), .B1(new_n759), .B2(G283), .ZN(new_n1171));
  OAI221_X1 g0971(.A(new_n1171), .B1(new_n202), .B2(new_n754), .C1(new_n370), .C2(new_n738), .ZN(new_n1172));
  AOI21_X1  g0972(.A(new_n958), .B1(new_n740), .B2(G116), .ZN(new_n1173));
  OAI211_X1 g0973(.A(new_n1173), .B(new_n383), .C1(new_n541), .C2(new_n749), .ZN(new_n1174));
  NOR4_X1   g0974(.A1(new_n1172), .A2(new_n1174), .A3(G41), .A4(new_n1001), .ZN(new_n1175));
  XNOR2_X1  g0975(.A(new_n1175), .B(KEYINPUT58), .ZN(new_n1176));
  OAI21_X1  g0976(.A(new_n778), .B1(new_n1170), .B2(new_n1176), .ZN(new_n1177));
  OAI211_X1 g0977(.A(new_n1156), .B(new_n1177), .C1(new_n1145), .C2(new_n780), .ZN(new_n1178));
  NAND2_X1  g0978(.A1(new_n1154), .A2(new_n1178), .ZN(new_n1179));
  AOI21_X1  g0979(.A(new_n1096), .B1(new_n1098), .B2(new_n1099), .ZN(new_n1180));
  NAND3_X1  g0980(.A1(new_n1057), .A2(new_n874), .A3(new_n656), .ZN(new_n1181));
  OAI21_X1  g0981(.A(new_n1153), .B1(new_n1180), .B2(new_n1181), .ZN(new_n1182));
  INV_X1    g0982(.A(KEYINPUT57), .ZN(new_n1183));
  AOI21_X1  g0983(.A(new_n684), .B1(new_n1182), .B2(new_n1183), .ZN(new_n1184));
  NOR2_X1   g0984(.A1(new_n1092), .A2(new_n1094), .ZN(new_n1185));
  OAI21_X1  g0985(.A(new_n1058), .B1(new_n1185), .B2(new_n1096), .ZN(new_n1186));
  OR2_X1    g0986(.A1(new_n1152), .A2(KEYINPUT124), .ZN(new_n1187));
  NAND3_X1  g0987(.A1(new_n1151), .A2(KEYINPUT124), .A3(new_n1152), .ZN(new_n1188));
  NAND4_X1  g0988(.A1(new_n1186), .A2(KEYINPUT57), .A3(new_n1187), .A4(new_n1188), .ZN(new_n1189));
  AOI21_X1  g0989(.A(new_n1179), .B1(new_n1184), .B2(new_n1189), .ZN(new_n1190));
  INV_X1    g0990(.A(new_n1190), .ZN(G375));
  NAND2_X1  g0991(.A1(new_n1075), .A2(new_n953), .ZN(new_n1192));
  INV_X1    g0992(.A(KEYINPUT125), .ZN(new_n1193));
  NAND2_X1  g0993(.A1(new_n1192), .A2(new_n1193), .ZN(new_n1194));
  NAND3_X1  g0994(.A1(new_n1075), .A2(KEYINPUT125), .A3(new_n953), .ZN(new_n1195));
  AND2_X1   g0995(.A1(new_n1194), .A2(new_n1195), .ZN(new_n1196));
  OAI22_X1  g0996(.A1(new_n749), .A2(new_n444), .B1(new_n741), .B2(new_n475), .ZN(new_n1197));
  NOR3_X1   g0997(.A1(new_n1197), .A2(new_n1003), .A3(new_n274), .ZN(new_n1198));
  NAND2_X1  g0998(.A1(new_n767), .A2(G97), .ZN(new_n1199));
  OAI22_X1  g0999(.A1(new_n744), .A2(new_n824), .B1(new_n758), .B2(new_n825), .ZN(new_n1200));
  AOI21_X1  g1000(.A(new_n1200), .B1(G107), .B2(new_n737), .ZN(new_n1201));
  NAND4_X1  g1001(.A1(new_n1198), .A2(new_n955), .A3(new_n1199), .A4(new_n1201), .ZN(new_n1202));
  NOR2_X1   g1002(.A1(new_n754), .A2(new_n202), .ZN(new_n1203));
  OAI22_X1  g1003(.A1(new_n738), .A2(new_n267), .B1(new_n755), .B2(new_n812), .ZN(new_n1204));
  AOI211_X1 g1004(.A(new_n1203), .B(new_n1204), .C1(G128), .C2(new_n759), .ZN(new_n1205));
  AOI22_X1  g1005(.A1(new_n818), .A2(G50), .B1(new_n1115), .B2(new_n748), .ZN(new_n1206));
  AOI21_X1  g1006(.A(new_n383), .B1(G137), .B2(new_n745), .ZN(new_n1207));
  NAND3_X1  g1007(.A1(new_n1205), .A2(new_n1206), .A3(new_n1207), .ZN(new_n1208));
  NOR2_X1   g1008(.A1(new_n741), .A2(new_n816), .ZN(new_n1209));
  OAI21_X1  g1009(.A(new_n1202), .B1(new_n1208), .B2(new_n1209), .ZN(new_n1210));
  AOI22_X1  g1010(.A1(new_n1210), .A2(new_n778), .B1(new_n203), .B2(new_n830), .ZN(new_n1211));
  OAI211_X1 g1011(.A(new_n732), .B(new_n1211), .C1(new_n868), .C2(new_n780), .ZN(new_n1212));
  NOR2_X1   g1012(.A1(new_n1075), .A2(new_n1058), .ZN(new_n1213));
  INV_X1    g1013(.A(new_n1213), .ZN(new_n1214));
  NAND3_X1  g1014(.A1(new_n1214), .A2(new_n929), .A3(new_n1096), .ZN(new_n1215));
  NAND3_X1  g1015(.A1(new_n1196), .A2(new_n1212), .A3(new_n1215), .ZN(G381));
  NAND2_X1  g1016(.A1(new_n1101), .A2(new_n1132), .ZN(new_n1217));
  NAND2_X1  g1017(.A1(new_n1217), .A2(KEYINPUT126), .ZN(new_n1218));
  INV_X1    g1018(.A(KEYINPUT126), .ZN(new_n1219));
  NAND3_X1  g1019(.A1(new_n1101), .A2(new_n1219), .A3(new_n1132), .ZN(new_n1220));
  NAND2_X1  g1020(.A1(new_n1218), .A2(new_n1220), .ZN(new_n1221));
  NAND2_X1  g1021(.A1(new_n1190), .A2(new_n1221), .ZN(new_n1222));
  NOR3_X1   g1022(.A1(new_n1222), .A2(G384), .A3(G381), .ZN(new_n1223));
  AND3_X1   g1023(.A1(new_n954), .A2(new_n1051), .A3(new_n981), .ZN(new_n1224));
  NAND3_X1  g1024(.A1(new_n1021), .A2(new_n791), .A3(new_n1023), .ZN(new_n1225));
  INV_X1    g1025(.A(new_n1225), .ZN(new_n1226));
  NAND3_X1  g1026(.A1(new_n1223), .A2(new_n1224), .A3(new_n1226), .ZN(G407));
  OAI211_X1 g1027(.A(G407), .B(G213), .C1(G343), .C2(new_n1222), .ZN(G409));
  NAND2_X1  g1028(.A1(G393), .A2(G396), .ZN(new_n1229));
  NAND2_X1  g1029(.A1(new_n1229), .A2(new_n1225), .ZN(new_n1230));
  AOI21_X1  g1030(.A(new_n1051), .B1(new_n981), .B2(new_n954), .ZN(new_n1231));
  OAI21_X1  g1031(.A(new_n1230), .B1(new_n1224), .B2(new_n1231), .ZN(new_n1232));
  NAND2_X1  g1032(.A1(G387), .A2(G390), .ZN(new_n1233));
  NAND3_X1  g1033(.A1(new_n954), .A2(new_n1051), .A3(new_n981), .ZN(new_n1234));
  INV_X1    g1034(.A(new_n1230), .ZN(new_n1235));
  NAND3_X1  g1035(.A1(new_n1233), .A2(new_n1234), .A3(new_n1235), .ZN(new_n1236));
  AND2_X1   g1036(.A1(new_n1232), .A2(new_n1236), .ZN(new_n1237));
  OR2_X1    g1037(.A1(new_n1071), .A2(new_n1074), .ZN(new_n1238));
  NAND4_X1  g1038(.A1(new_n1238), .A2(KEYINPUT60), .A3(new_n1181), .A4(new_n1066), .ZN(new_n1239));
  INV_X1    g1039(.A(KEYINPUT60), .ZN(new_n1240));
  OAI21_X1  g1040(.A(new_n1240), .B1(new_n1075), .B2(new_n1058), .ZN(new_n1241));
  NAND4_X1  g1041(.A1(new_n1239), .A2(new_n1241), .A3(new_n683), .A4(new_n1096), .ZN(new_n1242));
  NAND3_X1  g1042(.A1(new_n1196), .A2(new_n1212), .A3(new_n1242), .ZN(new_n1243));
  INV_X1    g1043(.A(G384), .ZN(new_n1244));
  NAND2_X1  g1044(.A1(new_n1243), .A2(new_n1244), .ZN(new_n1245));
  NAND4_X1  g1045(.A1(new_n1196), .A2(G384), .A3(new_n1212), .A4(new_n1242), .ZN(new_n1246));
  INV_X1    g1046(.A(G213), .ZN(new_n1247));
  NOR2_X1   g1047(.A1(new_n1247), .A2(G343), .ZN(new_n1248));
  NAND2_X1  g1048(.A1(new_n1248), .A2(KEYINPUT127), .ZN(new_n1249));
  NAND3_X1  g1049(.A1(new_n1245), .A2(new_n1246), .A3(new_n1249), .ZN(new_n1250));
  NAND2_X1  g1050(.A1(new_n1248), .A2(G2897), .ZN(new_n1251));
  NAND2_X1  g1051(.A1(new_n1250), .A2(new_n1251), .ZN(new_n1252));
  INV_X1    g1052(.A(new_n1251), .ZN(new_n1253));
  NAND4_X1  g1053(.A1(new_n1245), .A2(new_n1246), .A3(new_n1253), .A4(new_n1249), .ZN(new_n1254));
  NAND2_X1  g1054(.A1(new_n1252), .A2(new_n1254), .ZN(new_n1255));
  NAND3_X1  g1055(.A1(new_n1187), .A2(new_n1188), .A3(new_n953), .ZN(new_n1256));
  OAI211_X1 g1056(.A(new_n1256), .B(new_n1178), .C1(new_n1182), .C2(new_n930), .ZN(new_n1257));
  AOI22_X1  g1057(.A1(new_n1190), .A2(G378), .B1(new_n1221), .B2(new_n1257), .ZN(new_n1258));
  OAI21_X1  g1058(.A(new_n1255), .B1(new_n1258), .B2(new_n1248), .ZN(new_n1259));
  AND2_X1   g1059(.A1(new_n1151), .A2(new_n1152), .ZN(new_n1260));
  AOI21_X1  g1060(.A(new_n1181), .B1(new_n1105), .B2(new_n1075), .ZN(new_n1261));
  OAI21_X1  g1061(.A(new_n1183), .B1(new_n1260), .B2(new_n1261), .ZN(new_n1262));
  NAND3_X1  g1062(.A1(new_n1189), .A2(new_n1262), .A3(new_n683), .ZN(new_n1263));
  INV_X1    g1063(.A(new_n1179), .ZN(new_n1264));
  INV_X1    g1064(.A(new_n1135), .ZN(new_n1265));
  OAI211_X1 g1065(.A(new_n1263), .B(new_n1264), .C1(new_n1133), .C2(new_n1265), .ZN(new_n1266));
  INV_X1    g1066(.A(new_n1220), .ZN(new_n1267));
  AOI21_X1  g1067(.A(new_n1219), .B1(new_n1101), .B2(new_n1132), .ZN(new_n1268));
  OAI21_X1  g1068(.A(new_n1257), .B1(new_n1267), .B2(new_n1268), .ZN(new_n1269));
  NAND2_X1  g1069(.A1(new_n1266), .A2(new_n1269), .ZN(new_n1270));
  NAND2_X1  g1070(.A1(new_n1245), .A2(new_n1246), .ZN(new_n1271));
  INV_X1    g1071(.A(new_n1271), .ZN(new_n1272));
  INV_X1    g1072(.A(new_n1248), .ZN(new_n1273));
  NAND3_X1  g1073(.A1(new_n1270), .A2(new_n1272), .A3(new_n1273), .ZN(new_n1274));
  AOI21_X1  g1074(.A(KEYINPUT62), .B1(new_n1259), .B2(new_n1274), .ZN(new_n1275));
  INV_X1    g1075(.A(KEYINPUT61), .ZN(new_n1276));
  AOI211_X1 g1076(.A(new_n1271), .B(new_n1248), .C1(new_n1266), .C2(new_n1269), .ZN(new_n1277));
  INV_X1    g1077(.A(KEYINPUT62), .ZN(new_n1278));
  OAI21_X1  g1078(.A(new_n1276), .B1(new_n1277), .B2(new_n1278), .ZN(new_n1279));
  OAI21_X1  g1079(.A(new_n1237), .B1(new_n1275), .B2(new_n1279), .ZN(new_n1280));
  AOI21_X1  g1080(.A(KEYINPUT61), .B1(new_n1232), .B2(new_n1236), .ZN(new_n1281));
  NAND2_X1  g1081(.A1(new_n1277), .A2(KEYINPUT63), .ZN(new_n1282));
  INV_X1    g1082(.A(KEYINPUT63), .ZN(new_n1283));
  NAND2_X1  g1083(.A1(new_n1270), .A2(new_n1273), .ZN(new_n1284));
  AOI21_X1  g1084(.A(new_n1283), .B1(new_n1284), .B2(new_n1255), .ZN(new_n1285));
  OAI211_X1 g1085(.A(new_n1281), .B(new_n1282), .C1(new_n1285), .C2(new_n1277), .ZN(new_n1286));
  NAND2_X1  g1086(.A1(new_n1280), .A2(new_n1286), .ZN(G405));
  INV_X1    g1087(.A(new_n1221), .ZN(new_n1288));
  OAI21_X1  g1088(.A(new_n1266), .B1(new_n1288), .B2(new_n1190), .ZN(new_n1289));
  XNOR2_X1  g1089(.A(new_n1289), .B(new_n1272), .ZN(new_n1290));
  XNOR2_X1  g1090(.A(new_n1290), .B(new_n1237), .ZN(G402));
endmodule


