

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n513, n514, n515, n516,
         n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527,
         n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538,
         n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549,
         n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560,
         n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571,
         n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582,
         n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593,
         n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604,
         n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615,
         n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626,
         n627, n628, n629, n630, n631, n632, n633, n634, n635, n636, n637,
         n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, n648,
         n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659,
         n660, n661, n662, n663, n664, n665, n666, n667, n668, n669, n670,
         n671, n672, n673, n674, n675, n676, n677, n678, n679, n680, n681,
         n682, n683, n684, n685, n686, n687, n688, n689, n690, n691, n692,
         n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, n703,
         n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, n714,
         n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, n725,
         n726, n727, n728, n729, n730, n731, n732, n733, n734, n735, n736,
         n737, n738, n739, n740, n741, n742, n743, n744, n745, n746, n747,
         n748, n749, n750, n751, n752, n753, n754, n755, n756, n757, n758,
         n759, n760, n761, n762, n763, n764, n765, n766, n767, n768, n769,
         n770, n771, n772, n773, n774, n775, n776, n777, n778, n779, n780,
         n781, n782, n783, n784, n785, n786, n787, n788, n789, n790, n791,
         n792, n793, n794, n795, n796, n797, n798, n799, n800, n801, n802,
         n803, n804, n805, n806, n807, n808, n809, n810, n811, n812, n813,
         n814, n815, n816, n817, n818, n819, n820, n821, n822, n823, n824,
         n825, n826, n827, n828, n829, n830, n831, n832, n833, n834, n835,
         n836, n837, n838, n839, n840, n841, n842, n843, n844, n845, n846,
         n847, n848, n849, n850, n851, n852, n853, n854, n855, n856, n857,
         n858, n859, n860, n861, n862, n863, n864, n865, n866, n867, n868,
         n869, n870, n871, n872, n873, n874, n875, n876, n877, n878, n879,
         n880, n881, n882, n883, n884, n885, n886, n887, n888, n889, n890,
         n891, n892, n893, n894, n895, n896, n897, n898, n899, n900, n901,
         n902, n903, n904, n905, n906, n907, n908, n909, n910, n911, n912,
         n913, n914, n915, n916, n917, n918, n919, n920, n921, n922, n923,
         n924, n925, n926, n927, n928, n929, n930, n931, n932, n933, n934,
         n935, n936, n937, n938, n939, n940, n941, n942, n943, n944, n945,
         n946, n947, n948, n949, n950, n951, n952, n953, n954, n955, n956,
         n957, n958, n959, n960, n961, n962, n963, n964, n965, n966, n967,
         n968, n969, n970, n971, n972, n973, n974, n975, n976, n977, n978,
         n979, n980, n981, n982, n983, n984, n985, n986, n987, n988, n989,
         n990, n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000,
         n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010,
         n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  AND2_X2 U547 ( .A1(n683), .A2(n682), .ZN(n684) );
  XNOR2_X2 U548 ( .A(n589), .B(n588), .ZN(n753) );
  XNOR2_X2 U549 ( .A(KEYINPUT93), .B(n622), .ZN(n624) );
  NOR2_X2 U550 ( .A1(G1966), .A2(n656), .ZN(n671) );
  NAND2_X2 U551 ( .A1(G8), .A2(n658), .ZN(n656) );
  NOR2_X2 U552 ( .A1(n624), .A2(n623), .ZN(n633) );
  AND2_X1 U553 ( .A1(n704), .A2(n591), .ZN(n640) );
  BUF_X1 U554 ( .A(n583), .Z(n982) );
  NOR2_X1 U555 ( .A1(G2105), .A2(n520), .ZN(n577) );
  NOR2_X1 U556 ( .A1(n604), .A2(n997), .ZN(n606) );
  NAND2_X1 U557 ( .A1(n700), .A2(n514), .ZN(n701) );
  NOR2_X1 U558 ( .A1(G2104), .A2(G2105), .ZN(n517) );
  XNOR2_X1 U559 ( .A(n579), .B(n578), .ZN(n580) );
  XOR2_X1 U560 ( .A(KEYINPUT26), .B(KEYINPUT95), .Z(n513) );
  OR2_X1 U561 ( .A1(n656), .A2(n699), .ZN(n514) );
  XOR2_X1 U562 ( .A(KEYINPUT87), .B(n518), .Z(n515) );
  XNOR2_X1 U563 ( .A(n590), .B(n513), .ZN(n593) );
  INV_X1 U564 ( .A(KEYINPUT64), .ZN(n605) );
  XNOR2_X1 U565 ( .A(n606), .B(n605), .ZN(n618) );
  INV_X1 U566 ( .A(KEYINPUT29), .ZN(n638) );
  NOR2_X1 U567 ( .A1(n652), .A2(n651), .ZN(n653) );
  INV_X1 U568 ( .A(KEYINPUT23), .ZN(n578) );
  NOR2_X1 U569 ( .A1(G164), .A2(G1384), .ZN(n704) );
  INV_X1 U570 ( .A(KEYINPUT17), .ZN(n516) );
  NAND2_X1 U571 ( .A1(n583), .A2(G138), .ZN(n518) );
  XNOR2_X1 U572 ( .A(n517), .B(n516), .ZN(n583) );
  NOR2_X1 U573 ( .A1(G651), .A2(n567), .ZN(n783) );
  NOR2_X1 U574 ( .A1(n524), .A2(n523), .ZN(G164) );
  INV_X1 U575 ( .A(G2104), .ZN(n520) );
  BUF_X1 U576 ( .A(n577), .Z(n983) );
  NAND2_X1 U577 ( .A1(n983), .A2(G102), .ZN(n519) );
  NAND2_X1 U578 ( .A1(n519), .A2(n515), .ZN(n524) );
  AND2_X1 U579 ( .A1(G2104), .A2(G2105), .ZN(n978) );
  NAND2_X1 U580 ( .A1(G114), .A2(n978), .ZN(n522) );
  AND2_X1 U581 ( .A1(n520), .A2(G2105), .ZN(n979) );
  NAND2_X1 U582 ( .A1(G126), .A2(n979), .ZN(n521) );
  NAND2_X1 U583 ( .A1(n522), .A2(n521), .ZN(n523) );
  XOR2_X1 U584 ( .A(KEYINPUT0), .B(G543), .Z(n567) );
  INV_X1 U585 ( .A(G651), .ZN(n526) );
  NOR2_X1 U586 ( .A1(n567), .A2(n526), .ZN(n785) );
  NAND2_X1 U587 ( .A1(n785), .A2(G73), .ZN(n525) );
  XNOR2_X1 U588 ( .A(KEYINPUT2), .B(n525), .ZN(n532) );
  NOR2_X1 U589 ( .A1(G651), .A2(G543), .ZN(n788) );
  NAND2_X1 U590 ( .A1(G86), .A2(n788), .ZN(n529) );
  NOR2_X1 U591 ( .A1(G543), .A2(n526), .ZN(n527) );
  XOR2_X1 U592 ( .A(KEYINPUT1), .B(n527), .Z(n789) );
  NAND2_X1 U593 ( .A1(G61), .A2(n789), .ZN(n528) );
  NAND2_X1 U594 ( .A1(n529), .A2(n528), .ZN(n530) );
  XOR2_X1 U595 ( .A(KEYINPUT82), .B(n530), .Z(n531) );
  NAND2_X1 U596 ( .A1(n532), .A2(n531), .ZN(n533) );
  XNOR2_X1 U597 ( .A(n533), .B(KEYINPUT83), .ZN(n535) );
  NAND2_X1 U598 ( .A1(G48), .A2(n783), .ZN(n534) );
  NAND2_X1 U599 ( .A1(n535), .A2(n534), .ZN(G305) );
  NAND2_X1 U600 ( .A1(G64), .A2(n789), .ZN(n536) );
  XOR2_X1 U601 ( .A(KEYINPUT68), .B(n536), .Z(n543) );
  NAND2_X1 U602 ( .A1(G90), .A2(n788), .ZN(n538) );
  NAND2_X1 U603 ( .A1(G77), .A2(n785), .ZN(n537) );
  NAND2_X1 U604 ( .A1(n538), .A2(n537), .ZN(n539) );
  XNOR2_X1 U605 ( .A(n539), .B(KEYINPUT9), .ZN(n541) );
  NAND2_X1 U606 ( .A1(G52), .A2(n783), .ZN(n540) );
  NAND2_X1 U607 ( .A1(n541), .A2(n540), .ZN(n542) );
  NOR2_X1 U608 ( .A1(n543), .A2(n542), .ZN(G171) );
  NAND2_X1 U609 ( .A1(G63), .A2(n789), .ZN(n545) );
  NAND2_X1 U610 ( .A1(G51), .A2(n783), .ZN(n544) );
  NAND2_X1 U611 ( .A1(n545), .A2(n544), .ZN(n546) );
  XNOR2_X1 U612 ( .A(KEYINPUT6), .B(n546), .ZN(n554) );
  NAND2_X1 U613 ( .A1(G89), .A2(n788), .ZN(n547) );
  XNOR2_X1 U614 ( .A(n547), .B(KEYINPUT4), .ZN(n548) );
  XNOR2_X1 U615 ( .A(n548), .B(KEYINPUT74), .ZN(n550) );
  NAND2_X1 U616 ( .A1(G76), .A2(n785), .ZN(n549) );
  NAND2_X1 U617 ( .A1(n550), .A2(n549), .ZN(n551) );
  XNOR2_X1 U618 ( .A(KEYINPUT75), .B(n551), .ZN(n552) );
  XNOR2_X1 U619 ( .A(KEYINPUT5), .B(n552), .ZN(n553) );
  NOR2_X1 U620 ( .A1(n554), .A2(n553), .ZN(n555) );
  XOR2_X1 U621 ( .A(KEYINPUT7), .B(n555), .Z(G168) );
  XOR2_X1 U622 ( .A(G168), .B(KEYINPUT8), .Z(n556) );
  XNOR2_X1 U623 ( .A(KEYINPUT76), .B(n556), .ZN(G286) );
  NAND2_X1 U624 ( .A1(G88), .A2(n788), .ZN(n558) );
  NAND2_X1 U625 ( .A1(G75), .A2(n785), .ZN(n557) );
  NAND2_X1 U626 ( .A1(n558), .A2(n557), .ZN(n562) );
  NAND2_X1 U627 ( .A1(G62), .A2(n789), .ZN(n560) );
  NAND2_X1 U628 ( .A1(G50), .A2(n783), .ZN(n559) );
  NAND2_X1 U629 ( .A1(n560), .A2(n559), .ZN(n561) );
  NOR2_X1 U630 ( .A1(n562), .A2(n561), .ZN(G166) );
  INV_X1 U631 ( .A(G166), .ZN(G303) );
  NAND2_X1 U632 ( .A1(G49), .A2(n783), .ZN(n564) );
  NAND2_X1 U633 ( .A1(G74), .A2(G651), .ZN(n563) );
  NAND2_X1 U634 ( .A1(n564), .A2(n563), .ZN(n565) );
  XOR2_X1 U635 ( .A(KEYINPUT81), .B(n565), .Z(n566) );
  NOR2_X1 U636 ( .A1(n789), .A2(n566), .ZN(n569) );
  NAND2_X1 U637 ( .A1(n567), .A2(G87), .ZN(n568) );
  NAND2_X1 U638 ( .A1(n569), .A2(n568), .ZN(G288) );
  NAND2_X1 U639 ( .A1(G60), .A2(n789), .ZN(n571) );
  NAND2_X1 U640 ( .A1(G47), .A2(n783), .ZN(n570) );
  NAND2_X1 U641 ( .A1(n571), .A2(n570), .ZN(n575) );
  NAND2_X1 U642 ( .A1(G85), .A2(n788), .ZN(n573) );
  NAND2_X1 U643 ( .A1(G72), .A2(n785), .ZN(n572) );
  NAND2_X1 U644 ( .A1(n573), .A2(n572), .ZN(n574) );
  NOR2_X1 U645 ( .A1(n575), .A2(n574), .ZN(n576) );
  XNOR2_X1 U646 ( .A(n576), .B(KEYINPUT67), .ZN(G290) );
  XNOR2_X1 U647 ( .A(G1981), .B(G305), .ZN(n871) );
  NAND2_X1 U648 ( .A1(n979), .A2(G125), .ZN(n581) );
  NAND2_X1 U649 ( .A1(n577), .A2(G101), .ZN(n579) );
  NAND2_X1 U650 ( .A1(n581), .A2(n580), .ZN(n582) );
  XNOR2_X1 U651 ( .A(n582), .B(KEYINPUT66), .ZN(n587) );
  NAND2_X1 U652 ( .A1(G137), .A2(n982), .ZN(n585) );
  NAND2_X1 U653 ( .A1(G113), .A2(n978), .ZN(n584) );
  NAND2_X1 U654 ( .A1(n585), .A2(n584), .ZN(n586) );
  NOR2_X1 U655 ( .A1(n587), .A2(n586), .ZN(n589) );
  INV_X1 U656 ( .A(KEYINPUT65), .ZN(n588) );
  NAND2_X1 U657 ( .A1(n753), .A2(G40), .ZN(n703) );
  INV_X1 U658 ( .A(n703), .ZN(n591) );
  NAND2_X1 U659 ( .A1(n640), .A2(G1996), .ZN(n590) );
  NAND2_X1 U660 ( .A1(n704), .A2(n591), .ZN(n658) );
  NAND2_X1 U661 ( .A1(n658), .A2(G1341), .ZN(n592) );
  NAND2_X1 U662 ( .A1(n593), .A2(n592), .ZN(n604) );
  NAND2_X1 U663 ( .A1(n788), .A2(G81), .ZN(n594) );
  XNOR2_X1 U664 ( .A(n594), .B(KEYINPUT12), .ZN(n596) );
  NAND2_X1 U665 ( .A1(G68), .A2(n785), .ZN(n595) );
  NAND2_X1 U666 ( .A1(n596), .A2(n595), .ZN(n598) );
  XOR2_X1 U667 ( .A(KEYINPUT13), .B(KEYINPUT72), .Z(n597) );
  XNOR2_X1 U668 ( .A(n598), .B(n597), .ZN(n601) );
  NAND2_X1 U669 ( .A1(n789), .A2(G56), .ZN(n599) );
  XOR2_X1 U670 ( .A(KEYINPUT14), .B(n599), .Z(n600) );
  NOR2_X1 U671 ( .A1(n601), .A2(n600), .ZN(n603) );
  NAND2_X1 U672 ( .A1(n783), .A2(G43), .ZN(n602) );
  NAND2_X1 U673 ( .A1(n603), .A2(n602), .ZN(n997) );
  NAND2_X1 U674 ( .A1(G92), .A2(n788), .ZN(n608) );
  NAND2_X1 U675 ( .A1(G79), .A2(n785), .ZN(n607) );
  NAND2_X1 U676 ( .A1(n608), .A2(n607), .ZN(n612) );
  NAND2_X1 U677 ( .A1(G66), .A2(n789), .ZN(n610) );
  NAND2_X1 U678 ( .A1(G54), .A2(n783), .ZN(n609) );
  NAND2_X1 U679 ( .A1(n610), .A2(n609), .ZN(n611) );
  NOR2_X1 U680 ( .A1(n612), .A2(n611), .ZN(n613) );
  XOR2_X1 U681 ( .A(KEYINPUT15), .B(n613), .Z(n998) );
  INV_X1 U682 ( .A(n998), .ZN(n768) );
  OR2_X1 U683 ( .A1(n618), .A2(n768), .ZN(n617) );
  NOR2_X1 U684 ( .A1(n640), .A2(G1348), .ZN(n615) );
  NOR2_X1 U685 ( .A1(G2067), .A2(n658), .ZN(n614) );
  NOR2_X1 U686 ( .A1(n615), .A2(n614), .ZN(n616) );
  NAND2_X1 U687 ( .A1(n617), .A2(n616), .ZN(n620) );
  NAND2_X1 U688 ( .A1(n618), .A2(n768), .ZN(n619) );
  NAND2_X1 U689 ( .A1(n620), .A2(n619), .ZN(n632) );
  NAND2_X1 U690 ( .A1(G2072), .A2(n640), .ZN(n621) );
  XOR2_X1 U691 ( .A(KEYINPUT27), .B(n621), .Z(n622) );
  INV_X1 U692 ( .A(G1956), .ZN(n903) );
  NOR2_X1 U693 ( .A1(n640), .A2(n903), .ZN(n623) );
  NAND2_X1 U694 ( .A1(G65), .A2(n789), .ZN(n626) );
  NAND2_X1 U695 ( .A1(G53), .A2(n783), .ZN(n625) );
  NAND2_X1 U696 ( .A1(n626), .A2(n625), .ZN(n630) );
  NAND2_X1 U697 ( .A1(G91), .A2(n788), .ZN(n628) );
  NAND2_X1 U698 ( .A1(G78), .A2(n785), .ZN(n627) );
  NAND2_X1 U699 ( .A1(n628), .A2(n627), .ZN(n629) );
  NOR2_X1 U700 ( .A1(n630), .A2(n629), .ZN(n797) );
  NAND2_X1 U701 ( .A1(n633), .A2(n797), .ZN(n631) );
  NAND2_X1 U702 ( .A1(n632), .A2(n631), .ZN(n637) );
  NOR2_X1 U703 ( .A1(n633), .A2(n797), .ZN(n635) );
  XOR2_X1 U704 ( .A(KEYINPUT28), .B(KEYINPUT94), .Z(n634) );
  XNOR2_X1 U705 ( .A(n635), .B(n634), .ZN(n636) );
  NAND2_X1 U706 ( .A1(n637), .A2(n636), .ZN(n639) );
  XNOR2_X1 U707 ( .A(n639), .B(n638), .ZN(n645) );
  XOR2_X1 U708 ( .A(G2078), .B(KEYINPUT25), .Z(n927) );
  NAND2_X1 U709 ( .A1(n640), .A2(n927), .ZN(n642) );
  NAND2_X1 U710 ( .A1(G1961), .A2(n658), .ZN(n641) );
  NAND2_X1 U711 ( .A1(n642), .A2(n641), .ZN(n643) );
  XOR2_X1 U712 ( .A(KEYINPUT92), .B(n643), .Z(n650) );
  NAND2_X1 U713 ( .A1(n650), .A2(G171), .ZN(n644) );
  NAND2_X1 U714 ( .A1(n645), .A2(n644), .ZN(n655) );
  NOR2_X1 U715 ( .A1(G2084), .A2(n658), .ZN(n669) );
  NOR2_X1 U716 ( .A1(n671), .A2(n669), .ZN(n646) );
  NAND2_X1 U717 ( .A1(G8), .A2(n646), .ZN(n647) );
  XNOR2_X1 U718 ( .A(KEYINPUT30), .B(n647), .ZN(n648) );
  NOR2_X1 U719 ( .A1(G168), .A2(n648), .ZN(n649) );
  XNOR2_X1 U720 ( .A(n649), .B(KEYINPUT96), .ZN(n652) );
  NOR2_X1 U721 ( .A1(n650), .A2(G171), .ZN(n651) );
  XOR2_X1 U722 ( .A(KEYINPUT31), .B(n653), .Z(n654) );
  NAND2_X1 U723 ( .A1(n655), .A2(n654), .ZN(n673) );
  NAND2_X1 U724 ( .A1(n673), .A2(G286), .ZN(n663) );
  NOR2_X1 U725 ( .A1(G1971), .A2(n656), .ZN(n657) );
  XNOR2_X1 U726 ( .A(n657), .B(KEYINPUT98), .ZN(n660) );
  NOR2_X1 U727 ( .A1(n658), .A2(G2090), .ZN(n659) );
  NOR2_X1 U728 ( .A1(n660), .A2(n659), .ZN(n661) );
  NAND2_X1 U729 ( .A1(n661), .A2(G303), .ZN(n662) );
  NAND2_X1 U730 ( .A1(n663), .A2(n662), .ZN(n664) );
  NAND2_X1 U731 ( .A1(n664), .A2(G8), .ZN(n666) );
  XOR2_X1 U732 ( .A(KEYINPUT32), .B(KEYINPUT99), .Z(n665) );
  XNOR2_X1 U733 ( .A(n666), .B(n665), .ZN(n691) );
  NAND2_X1 U734 ( .A1(G1976), .A2(G288), .ZN(n878) );
  INV_X1 U735 ( .A(n656), .ZN(n667) );
  NAND2_X1 U736 ( .A1(n878), .A2(n667), .ZN(n679) );
  INV_X1 U737 ( .A(n679), .ZN(n668) );
  AND2_X1 U738 ( .A1(n691), .A2(n668), .ZN(n677) );
  NAND2_X1 U739 ( .A1(G8), .A2(n669), .ZN(n670) );
  XNOR2_X1 U740 ( .A(KEYINPUT91), .B(n670), .ZN(n675) );
  INV_X1 U741 ( .A(n671), .ZN(n672) );
  NAND2_X1 U742 ( .A1(n673), .A2(n672), .ZN(n674) );
  NOR2_X1 U743 ( .A1(n675), .A2(n674), .ZN(n676) );
  XNOR2_X1 U744 ( .A(KEYINPUT97), .B(n676), .ZN(n692) );
  NAND2_X1 U745 ( .A1(n677), .A2(n692), .ZN(n683) );
  INV_X1 U746 ( .A(KEYINPUT33), .ZN(n681) );
  NOR2_X1 U747 ( .A1(G1976), .A2(G288), .ZN(n685) );
  NOR2_X1 U748 ( .A1(G1971), .A2(G303), .ZN(n678) );
  NOR2_X1 U749 ( .A1(n685), .A2(n678), .ZN(n879) );
  OR2_X1 U750 ( .A1(n679), .A2(n879), .ZN(n680) );
  AND2_X1 U751 ( .A1(n681), .A2(n680), .ZN(n682) );
  XNOR2_X1 U752 ( .A(n684), .B(KEYINPUT100), .ZN(n688) );
  NAND2_X1 U753 ( .A1(n685), .A2(KEYINPUT33), .ZN(n686) );
  NOR2_X1 U754 ( .A1(n656), .A2(n686), .ZN(n687) );
  NOR2_X1 U755 ( .A1(n688), .A2(n687), .ZN(n689) );
  XNOR2_X1 U756 ( .A(n689), .B(KEYINPUT101), .ZN(n690) );
  NOR2_X1 U757 ( .A1(n871), .A2(n690), .ZN(n702) );
  NAND2_X1 U758 ( .A1(n692), .A2(n691), .ZN(n695) );
  NOR2_X1 U759 ( .A1(G2090), .A2(G303), .ZN(n693) );
  NAND2_X1 U760 ( .A1(G8), .A2(n693), .ZN(n694) );
  NAND2_X1 U761 ( .A1(n695), .A2(n694), .ZN(n696) );
  XNOR2_X1 U762 ( .A(KEYINPUT102), .B(n696), .ZN(n697) );
  NAND2_X1 U763 ( .A1(n656), .A2(n697), .ZN(n700) );
  NOR2_X1 U764 ( .A1(G1981), .A2(G305), .ZN(n698) );
  XOR2_X1 U765 ( .A(n698), .B(KEYINPUT24), .Z(n699) );
  NOR2_X1 U766 ( .A1(n702), .A2(n701), .ZN(n734) );
  NOR2_X1 U767 ( .A1(n704), .A2(n703), .ZN(n747) );
  NAND2_X1 U768 ( .A1(G140), .A2(n982), .ZN(n706) );
  NAND2_X1 U769 ( .A1(G104), .A2(n983), .ZN(n705) );
  NAND2_X1 U770 ( .A1(n706), .A2(n705), .ZN(n707) );
  XNOR2_X1 U771 ( .A(KEYINPUT34), .B(n707), .ZN(n712) );
  NAND2_X1 U772 ( .A1(G116), .A2(n978), .ZN(n709) );
  NAND2_X1 U773 ( .A1(G128), .A2(n979), .ZN(n708) );
  NAND2_X1 U774 ( .A1(n709), .A2(n708), .ZN(n710) );
  XOR2_X1 U775 ( .A(KEYINPUT35), .B(n710), .Z(n711) );
  NOR2_X1 U776 ( .A1(n712), .A2(n711), .ZN(n713) );
  XNOR2_X1 U777 ( .A(KEYINPUT36), .B(n713), .ZN(n992) );
  XNOR2_X1 U778 ( .A(G2067), .B(KEYINPUT37), .ZN(n745) );
  NOR2_X1 U779 ( .A1(n992), .A2(n745), .ZN(n856) );
  NAND2_X1 U780 ( .A1(n747), .A2(n856), .ZN(n744) );
  NAND2_X1 U781 ( .A1(G131), .A2(n982), .ZN(n715) );
  NAND2_X1 U782 ( .A1(G95), .A2(n983), .ZN(n714) );
  NAND2_X1 U783 ( .A1(n715), .A2(n714), .ZN(n719) );
  NAND2_X1 U784 ( .A1(G107), .A2(n978), .ZN(n717) );
  NAND2_X1 U785 ( .A1(G119), .A2(n979), .ZN(n716) );
  NAND2_X1 U786 ( .A1(n717), .A2(n716), .ZN(n718) );
  OR2_X1 U787 ( .A1(n719), .A2(n718), .ZN(n970) );
  NAND2_X1 U788 ( .A1(G1991), .A2(n970), .ZN(n730) );
  NAND2_X1 U789 ( .A1(G105), .A2(n983), .ZN(n720) );
  XNOR2_X1 U790 ( .A(n720), .B(KEYINPUT38), .ZN(n728) );
  NAND2_X1 U791 ( .A1(n978), .A2(G117), .ZN(n721) );
  XNOR2_X1 U792 ( .A(n721), .B(KEYINPUT88), .ZN(n723) );
  NAND2_X1 U793 ( .A1(G129), .A2(n979), .ZN(n722) );
  NAND2_X1 U794 ( .A1(n723), .A2(n722), .ZN(n726) );
  NAND2_X1 U795 ( .A1(G141), .A2(n982), .ZN(n724) );
  XNOR2_X1 U796 ( .A(KEYINPUT89), .B(n724), .ZN(n725) );
  NOR2_X1 U797 ( .A1(n726), .A2(n725), .ZN(n727) );
  NAND2_X1 U798 ( .A1(n728), .A2(n727), .ZN(n974) );
  NAND2_X1 U799 ( .A1(G1996), .A2(n974), .ZN(n729) );
  NAND2_X1 U800 ( .A1(n730), .A2(n729), .ZN(n843) );
  NAND2_X1 U801 ( .A1(n843), .A2(n747), .ZN(n731) );
  XOR2_X1 U802 ( .A(KEYINPUT90), .B(n731), .Z(n739) );
  INV_X1 U803 ( .A(n739), .ZN(n732) );
  NAND2_X1 U804 ( .A1(n744), .A2(n732), .ZN(n733) );
  NOR2_X1 U805 ( .A1(n734), .A2(n733), .ZN(n736) );
  XNOR2_X1 U806 ( .A(G1986), .B(G290), .ZN(n875) );
  NAND2_X1 U807 ( .A1(n875), .A2(n747), .ZN(n735) );
  NAND2_X1 U808 ( .A1(n736), .A2(n735), .ZN(n751) );
  NOR2_X1 U809 ( .A1(G1996), .A2(n974), .ZN(n850) );
  NOR2_X1 U810 ( .A1(G1986), .A2(G290), .ZN(n737) );
  NOR2_X1 U811 ( .A1(G1991), .A2(n970), .ZN(n844) );
  NOR2_X1 U812 ( .A1(n737), .A2(n844), .ZN(n738) );
  NOR2_X1 U813 ( .A1(n739), .A2(n738), .ZN(n740) );
  NOR2_X1 U814 ( .A1(n850), .A2(n740), .ZN(n741) );
  XOR2_X1 U815 ( .A(n741), .B(KEYINPUT103), .Z(n742) );
  XNOR2_X1 U816 ( .A(KEYINPUT39), .B(n742), .ZN(n743) );
  NAND2_X1 U817 ( .A1(n744), .A2(n743), .ZN(n746) );
  NAND2_X1 U818 ( .A1(n992), .A2(n745), .ZN(n860) );
  NAND2_X1 U819 ( .A1(n746), .A2(n860), .ZN(n748) );
  NAND2_X1 U820 ( .A1(n748), .A2(n747), .ZN(n749) );
  XNOR2_X1 U821 ( .A(KEYINPUT104), .B(n749), .ZN(n750) );
  NAND2_X1 U822 ( .A1(n751), .A2(n750), .ZN(n752) );
  XNOR2_X1 U823 ( .A(n752), .B(KEYINPUT40), .ZN(G329) );
  BUF_X1 U824 ( .A(n753), .Z(G160) );
  NAND2_X1 U825 ( .A1(G111), .A2(n978), .ZN(n760) );
  NAND2_X1 U826 ( .A1(G135), .A2(n982), .ZN(n755) );
  NAND2_X1 U827 ( .A1(G99), .A2(n983), .ZN(n754) );
  NAND2_X1 U828 ( .A1(n755), .A2(n754), .ZN(n758) );
  NAND2_X1 U829 ( .A1(n979), .A2(G123), .ZN(n756) );
  XOR2_X1 U830 ( .A(KEYINPUT18), .B(n756), .Z(n757) );
  NOR2_X1 U831 ( .A1(n758), .A2(n757), .ZN(n759) );
  NAND2_X1 U832 ( .A1(n760), .A2(n759), .ZN(n761) );
  XNOR2_X1 U833 ( .A(n761), .B(KEYINPUT78), .ZN(n972) );
  XNOR2_X1 U834 ( .A(n972), .B(G2096), .ZN(n762) );
  OR2_X1 U835 ( .A1(G2100), .A2(n762), .ZN(G156) );
  INV_X1 U836 ( .A(G57), .ZN(G237) );
  INV_X1 U837 ( .A(n797), .ZN(G299) );
  NAND2_X1 U838 ( .A1(G94), .A2(G452), .ZN(n763) );
  XNOR2_X1 U839 ( .A(n763), .B(KEYINPUT69), .ZN(G173) );
  NAND2_X1 U840 ( .A1(G7), .A2(G661), .ZN(n764) );
  XNOR2_X1 U841 ( .A(n764), .B(KEYINPUT10), .ZN(n765) );
  XNOR2_X1 U842 ( .A(KEYINPUT70), .B(n765), .ZN(G223) );
  INV_X1 U843 ( .A(G223), .ZN(n821) );
  NAND2_X1 U844 ( .A1(n821), .A2(G567), .ZN(n766) );
  XNOR2_X1 U845 ( .A(n766), .B(KEYINPUT11), .ZN(n767) );
  XNOR2_X1 U846 ( .A(KEYINPUT71), .B(n767), .ZN(G234) );
  XNOR2_X1 U847 ( .A(G860), .B(KEYINPUT73), .ZN(n774) );
  OR2_X1 U848 ( .A1(n997), .A2(n774), .ZN(G153) );
  INV_X1 U849 ( .A(G171), .ZN(G301) );
  NAND2_X1 U850 ( .A1(G868), .A2(G301), .ZN(n770) );
  INV_X1 U851 ( .A(G868), .ZN(n771) );
  NAND2_X1 U852 ( .A1(n768), .A2(n771), .ZN(n769) );
  NAND2_X1 U853 ( .A1(n770), .A2(n769), .ZN(G284) );
  NAND2_X1 U854 ( .A1(G868), .A2(G286), .ZN(n773) );
  NAND2_X1 U855 ( .A1(G299), .A2(n771), .ZN(n772) );
  NAND2_X1 U856 ( .A1(n773), .A2(n772), .ZN(G297) );
  NAND2_X1 U857 ( .A1(n774), .A2(G559), .ZN(n775) );
  NAND2_X1 U858 ( .A1(n775), .A2(n998), .ZN(n776) );
  XNOR2_X1 U859 ( .A(n776), .B(KEYINPUT77), .ZN(n777) );
  XOR2_X1 U860 ( .A(KEYINPUT16), .B(n777), .Z(G148) );
  NOR2_X1 U861 ( .A1(G868), .A2(n997), .ZN(n780) );
  NAND2_X1 U862 ( .A1(n998), .A2(G868), .ZN(n778) );
  NOR2_X1 U863 ( .A1(G559), .A2(n778), .ZN(n779) );
  NOR2_X1 U864 ( .A1(n780), .A2(n779), .ZN(G282) );
  XNOR2_X1 U865 ( .A(n997), .B(KEYINPUT79), .ZN(n782) );
  NAND2_X1 U866 ( .A1(n998), .A2(G559), .ZN(n781) );
  XOR2_X1 U867 ( .A(n782), .B(n781), .Z(n804) );
  NOR2_X1 U868 ( .A1(n804), .A2(G860), .ZN(n794) );
  NAND2_X1 U869 ( .A1(G55), .A2(n783), .ZN(n784) );
  XNOR2_X1 U870 ( .A(n784), .B(KEYINPUT80), .ZN(n787) );
  NAND2_X1 U871 ( .A1(n785), .A2(G80), .ZN(n786) );
  NAND2_X1 U872 ( .A1(n787), .A2(n786), .ZN(n793) );
  NAND2_X1 U873 ( .A1(G93), .A2(n788), .ZN(n791) );
  NAND2_X1 U874 ( .A1(G67), .A2(n789), .ZN(n790) );
  NAND2_X1 U875 ( .A1(n791), .A2(n790), .ZN(n792) );
  NOR2_X1 U876 ( .A1(n793), .A2(n792), .ZN(n796) );
  XNOR2_X1 U877 ( .A(n794), .B(n796), .ZN(G145) );
  NOR2_X1 U878 ( .A1(G868), .A2(n796), .ZN(n795) );
  XNOR2_X1 U879 ( .A(n795), .B(KEYINPUT85), .ZN(n807) );
  XNOR2_X1 U880 ( .A(n797), .B(n796), .ZN(n801) );
  XNOR2_X1 U881 ( .A(KEYINPUT84), .B(KEYINPUT19), .ZN(n799) );
  XNOR2_X1 U882 ( .A(G290), .B(G166), .ZN(n798) );
  XNOR2_X1 U883 ( .A(n799), .B(n798), .ZN(n800) );
  XNOR2_X1 U884 ( .A(n801), .B(n800), .ZN(n802) );
  XOR2_X1 U885 ( .A(n802), .B(G305), .Z(n803) );
  XNOR2_X1 U886 ( .A(G288), .B(n803), .ZN(n999) );
  XOR2_X1 U887 ( .A(n804), .B(n999), .Z(n805) );
  NAND2_X1 U888 ( .A1(G868), .A2(n805), .ZN(n806) );
  NAND2_X1 U889 ( .A1(n807), .A2(n806), .ZN(G295) );
  NAND2_X1 U890 ( .A1(G2078), .A2(G2084), .ZN(n808) );
  XOR2_X1 U891 ( .A(KEYINPUT20), .B(n808), .Z(n809) );
  NAND2_X1 U892 ( .A1(G2090), .A2(n809), .ZN(n810) );
  XNOR2_X1 U893 ( .A(KEYINPUT21), .B(n810), .ZN(n811) );
  NAND2_X1 U894 ( .A1(n811), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U895 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NAND2_X1 U896 ( .A1(G132), .A2(G82), .ZN(n812) );
  XNOR2_X1 U897 ( .A(n812), .B(KEYINPUT22), .ZN(n813) );
  XNOR2_X1 U898 ( .A(n813), .B(KEYINPUT86), .ZN(n814) );
  NOR2_X1 U899 ( .A1(G218), .A2(n814), .ZN(n815) );
  NAND2_X1 U900 ( .A1(G96), .A2(n815), .ZN(n947) );
  NAND2_X1 U901 ( .A1(G2106), .A2(n947), .ZN(n819) );
  NAND2_X1 U902 ( .A1(G120), .A2(G108), .ZN(n816) );
  NOR2_X1 U903 ( .A1(G237), .A2(n816), .ZN(n817) );
  NAND2_X1 U904 ( .A1(G69), .A2(n817), .ZN(n948) );
  NAND2_X1 U905 ( .A1(G567), .A2(n948), .ZN(n818) );
  NAND2_X1 U906 ( .A1(n819), .A2(n818), .ZN(n949) );
  NAND2_X1 U907 ( .A1(G661), .A2(G483), .ZN(n820) );
  NOR2_X1 U908 ( .A1(n949), .A2(n820), .ZN(n824) );
  NAND2_X1 U909 ( .A1(n824), .A2(G36), .ZN(G176) );
  NAND2_X1 U910 ( .A1(G2106), .A2(n821), .ZN(G217) );
  AND2_X1 U911 ( .A1(G15), .A2(G2), .ZN(n822) );
  NAND2_X1 U912 ( .A1(G661), .A2(n822), .ZN(G259) );
  NAND2_X1 U913 ( .A1(G3), .A2(G1), .ZN(n823) );
  NAND2_X1 U914 ( .A1(n824), .A2(n823), .ZN(G188) );
  XOR2_X1 U915 ( .A(G108), .B(KEYINPUT112), .Z(G238) );
  NAND2_X1 U917 ( .A1(G124), .A2(n979), .ZN(n825) );
  XNOR2_X1 U918 ( .A(n825), .B(KEYINPUT44), .ZN(n826) );
  XNOR2_X1 U919 ( .A(n826), .B(KEYINPUT108), .ZN(n828) );
  NAND2_X1 U920 ( .A1(G100), .A2(n983), .ZN(n827) );
  NAND2_X1 U921 ( .A1(n828), .A2(n827), .ZN(n832) );
  NAND2_X1 U922 ( .A1(G136), .A2(n982), .ZN(n830) );
  NAND2_X1 U923 ( .A1(G112), .A2(n978), .ZN(n829) );
  NAND2_X1 U924 ( .A1(n830), .A2(n829), .ZN(n831) );
  NOR2_X1 U925 ( .A1(n832), .A2(n831), .ZN(G162) );
  INV_X1 U926 ( .A(KEYINPUT55), .ZN(n940) );
  XOR2_X1 U927 ( .A(KEYINPUT116), .B(KEYINPUT52), .Z(n863) );
  NAND2_X1 U928 ( .A1(G139), .A2(n982), .ZN(n834) );
  NAND2_X1 U929 ( .A1(G103), .A2(n983), .ZN(n833) );
  NAND2_X1 U930 ( .A1(n834), .A2(n833), .ZN(n839) );
  NAND2_X1 U931 ( .A1(G115), .A2(n978), .ZN(n836) );
  NAND2_X1 U932 ( .A1(G127), .A2(n979), .ZN(n835) );
  NAND2_X1 U933 ( .A1(n836), .A2(n835), .ZN(n837) );
  XOR2_X1 U934 ( .A(KEYINPUT47), .B(n837), .Z(n838) );
  NOR2_X1 U935 ( .A1(n839), .A2(n838), .ZN(n977) );
  XOR2_X1 U936 ( .A(G2072), .B(n977), .Z(n841) );
  XOR2_X1 U937 ( .A(G164), .B(G2078), .Z(n840) );
  NOR2_X1 U938 ( .A1(n841), .A2(n840), .ZN(n842) );
  XOR2_X1 U939 ( .A(KEYINPUT50), .B(n842), .Z(n859) );
  NOR2_X1 U940 ( .A1(n844), .A2(n843), .ZN(n845) );
  NAND2_X1 U941 ( .A1(n972), .A2(n845), .ZN(n847) );
  XOR2_X1 U942 ( .A(G160), .B(G2084), .Z(n846) );
  NOR2_X1 U943 ( .A1(n847), .A2(n846), .ZN(n854) );
  XNOR2_X1 U944 ( .A(KEYINPUT51), .B(KEYINPUT114), .ZN(n852) );
  XNOR2_X1 U945 ( .A(G2090), .B(G162), .ZN(n848) );
  XNOR2_X1 U946 ( .A(n848), .B(KEYINPUT113), .ZN(n849) );
  NOR2_X1 U947 ( .A1(n850), .A2(n849), .ZN(n851) );
  XOR2_X1 U948 ( .A(n852), .B(n851), .Z(n853) );
  NAND2_X1 U949 ( .A1(n854), .A2(n853), .ZN(n855) );
  NOR2_X1 U950 ( .A1(n856), .A2(n855), .ZN(n857) );
  XNOR2_X1 U951 ( .A(KEYINPUT115), .B(n857), .ZN(n858) );
  NOR2_X1 U952 ( .A1(n859), .A2(n858), .ZN(n861) );
  NAND2_X1 U953 ( .A1(n861), .A2(n860), .ZN(n862) );
  XNOR2_X1 U954 ( .A(n863), .B(n862), .ZN(n864) );
  NAND2_X1 U955 ( .A1(n940), .A2(n864), .ZN(n865) );
  NAND2_X1 U956 ( .A1(n865), .A2(G29), .ZN(n920) );
  XOR2_X1 U957 ( .A(KEYINPUT56), .B(G16), .Z(n891) );
  XOR2_X1 U958 ( .A(G1341), .B(KEYINPUT122), .Z(n866) );
  XNOR2_X1 U959 ( .A(n997), .B(n866), .ZN(n869) );
  XNOR2_X1 U960 ( .A(G171), .B(G1961), .ZN(n867) );
  XNOR2_X1 U961 ( .A(n867), .B(KEYINPUT120), .ZN(n868) );
  NAND2_X1 U962 ( .A1(n869), .A2(n868), .ZN(n888) );
  XOR2_X1 U963 ( .A(G168), .B(G1966), .Z(n870) );
  NOR2_X1 U964 ( .A1(n871), .A2(n870), .ZN(n872) );
  XNOR2_X1 U965 ( .A(KEYINPUT57), .B(n872), .ZN(n873) );
  XNOR2_X1 U966 ( .A(n873), .B(KEYINPUT119), .ZN(n886) );
  XNOR2_X1 U967 ( .A(n998), .B(G1348), .ZN(n877) );
  XNOR2_X1 U968 ( .A(G1956), .B(G299), .ZN(n874) );
  NOR2_X1 U969 ( .A1(n875), .A2(n874), .ZN(n876) );
  NAND2_X1 U970 ( .A1(n877), .A2(n876), .ZN(n884) );
  AND2_X1 U971 ( .A1(G303), .A2(G1971), .ZN(n881) );
  NAND2_X1 U972 ( .A1(n879), .A2(n878), .ZN(n880) );
  NOR2_X1 U973 ( .A1(n881), .A2(n880), .ZN(n882) );
  XNOR2_X1 U974 ( .A(KEYINPUT121), .B(n882), .ZN(n883) );
  NOR2_X1 U975 ( .A1(n884), .A2(n883), .ZN(n885) );
  NAND2_X1 U976 ( .A1(n886), .A2(n885), .ZN(n887) );
  NOR2_X1 U977 ( .A1(n888), .A2(n887), .ZN(n889) );
  XOR2_X1 U978 ( .A(KEYINPUT123), .B(n889), .Z(n890) );
  NOR2_X1 U979 ( .A1(n891), .A2(n890), .ZN(n918) );
  XNOR2_X1 U980 ( .A(G1986), .B(G24), .ZN(n893) );
  XNOR2_X1 U981 ( .A(G1971), .B(G22), .ZN(n892) );
  NOR2_X1 U982 ( .A1(n893), .A2(n892), .ZN(n895) );
  XOR2_X1 U983 ( .A(G1976), .B(G23), .Z(n894) );
  NAND2_X1 U984 ( .A1(n895), .A2(n894), .ZN(n897) );
  XOR2_X1 U985 ( .A(KEYINPUT126), .B(KEYINPUT58), .Z(n896) );
  XNOR2_X1 U986 ( .A(n897), .B(n896), .ZN(n901) );
  XNOR2_X1 U987 ( .A(G1961), .B(G5), .ZN(n899) );
  XNOR2_X1 U988 ( .A(G21), .B(G1966), .ZN(n898) );
  NOR2_X1 U989 ( .A1(n899), .A2(n898), .ZN(n900) );
  NAND2_X1 U990 ( .A1(n901), .A2(n900), .ZN(n913) );
  XOR2_X1 U991 ( .A(G1348), .B(KEYINPUT59), .Z(n902) );
  XNOR2_X1 U992 ( .A(G4), .B(n902), .ZN(n910) );
  XNOR2_X1 U993 ( .A(G20), .B(n903), .ZN(n907) );
  XNOR2_X1 U994 ( .A(G1341), .B(G19), .ZN(n905) );
  XNOR2_X1 U995 ( .A(G6), .B(G1981), .ZN(n904) );
  NOR2_X1 U996 ( .A1(n905), .A2(n904), .ZN(n906) );
  NAND2_X1 U997 ( .A1(n907), .A2(n906), .ZN(n908) );
  XOR2_X1 U998 ( .A(KEYINPUT125), .B(n908), .Z(n909) );
  NOR2_X1 U999 ( .A1(n910), .A2(n909), .ZN(n911) );
  XOR2_X1 U1000 ( .A(KEYINPUT60), .B(n911), .Z(n912) );
  NOR2_X1 U1001 ( .A1(n913), .A2(n912), .ZN(n914) );
  XOR2_X1 U1002 ( .A(KEYINPUT61), .B(n914), .Z(n916) );
  XNOR2_X1 U1003 ( .A(G16), .B(KEYINPUT124), .ZN(n915) );
  NOR2_X1 U1004 ( .A1(n916), .A2(n915), .ZN(n917) );
  NOR2_X1 U1005 ( .A1(n918), .A2(n917), .ZN(n919) );
  NAND2_X1 U1006 ( .A1(n920), .A2(n919), .ZN(n945) );
  XNOR2_X1 U1007 ( .A(G2090), .B(G35), .ZN(n935) );
  XOR2_X1 U1008 ( .A(G1991), .B(G25), .Z(n921) );
  NAND2_X1 U1009 ( .A1(G28), .A2(n921), .ZN(n922) );
  XNOR2_X1 U1010 ( .A(n922), .B(KEYINPUT117), .ZN(n926) );
  XNOR2_X1 U1011 ( .A(G1996), .B(G32), .ZN(n924) );
  XNOR2_X1 U1012 ( .A(G2067), .B(G26), .ZN(n923) );
  NOR2_X1 U1013 ( .A1(n924), .A2(n923), .ZN(n925) );
  NAND2_X1 U1014 ( .A1(n926), .A2(n925), .ZN(n932) );
  XOR2_X1 U1015 ( .A(n927), .B(G27), .Z(n930) );
  XOR2_X1 U1016 ( .A(G33), .B(KEYINPUT118), .Z(n928) );
  XNOR2_X1 U1017 ( .A(G2072), .B(n928), .ZN(n929) );
  NAND2_X1 U1018 ( .A1(n930), .A2(n929), .ZN(n931) );
  NOR2_X1 U1019 ( .A1(n932), .A2(n931), .ZN(n933) );
  XNOR2_X1 U1020 ( .A(KEYINPUT53), .B(n933), .ZN(n934) );
  NOR2_X1 U1021 ( .A1(n935), .A2(n934), .ZN(n938) );
  XOR2_X1 U1022 ( .A(G2084), .B(KEYINPUT54), .Z(n936) );
  XNOR2_X1 U1023 ( .A(G34), .B(n936), .ZN(n937) );
  NAND2_X1 U1024 ( .A1(n938), .A2(n937), .ZN(n939) );
  XNOR2_X1 U1025 ( .A(n940), .B(n939), .ZN(n942) );
  INV_X1 U1026 ( .A(G29), .ZN(n941) );
  NAND2_X1 U1027 ( .A1(n942), .A2(n941), .ZN(n943) );
  NAND2_X1 U1028 ( .A1(G11), .A2(n943), .ZN(n944) );
  NOR2_X1 U1029 ( .A1(n945), .A2(n944), .ZN(n946) );
  XNOR2_X1 U1030 ( .A(n946), .B(KEYINPUT62), .ZN(G311) );
  XNOR2_X1 U1031 ( .A(KEYINPUT127), .B(G311), .ZN(G150) );
  INV_X1 U1032 ( .A(G132), .ZN(G219) );
  INV_X1 U1033 ( .A(G120), .ZN(G236) );
  INV_X1 U1034 ( .A(G82), .ZN(G220) );
  NOR2_X1 U1035 ( .A1(n948), .A2(n947), .ZN(G325) );
  INV_X1 U1036 ( .A(G325), .ZN(G261) );
  XOR2_X1 U1037 ( .A(KEYINPUT106), .B(n949), .Z(G319) );
  XOR2_X1 U1038 ( .A(KEYINPUT107), .B(G2084), .Z(n951) );
  XNOR2_X1 U1039 ( .A(G2067), .B(G2078), .ZN(n950) );
  XNOR2_X1 U1040 ( .A(n951), .B(n950), .ZN(n952) );
  XOR2_X1 U1041 ( .A(n952), .B(G2678), .Z(n954) );
  XNOR2_X1 U1042 ( .A(G2072), .B(KEYINPUT42), .ZN(n953) );
  XNOR2_X1 U1043 ( .A(n954), .B(n953), .ZN(n958) );
  XOR2_X1 U1044 ( .A(G2100), .B(G2096), .Z(n956) );
  XNOR2_X1 U1045 ( .A(G2090), .B(KEYINPUT43), .ZN(n955) );
  XNOR2_X1 U1046 ( .A(n956), .B(n955), .ZN(n957) );
  XOR2_X1 U1047 ( .A(n958), .B(n957), .Z(G227) );
  XOR2_X1 U1048 ( .A(G1981), .B(G1966), .Z(n960) );
  XNOR2_X1 U1049 ( .A(G1986), .B(G1961), .ZN(n959) );
  XNOR2_X1 U1050 ( .A(n960), .B(n959), .ZN(n961) );
  XOR2_X1 U1051 ( .A(n961), .B(KEYINPUT41), .Z(n963) );
  XNOR2_X1 U1052 ( .A(G1991), .B(G1956), .ZN(n962) );
  XNOR2_X1 U1053 ( .A(n963), .B(n962), .ZN(n967) );
  XOR2_X1 U1054 ( .A(G2474), .B(G1976), .Z(n965) );
  XNOR2_X1 U1055 ( .A(G1996), .B(G1971), .ZN(n964) );
  XNOR2_X1 U1056 ( .A(n965), .B(n964), .ZN(n966) );
  XNOR2_X1 U1057 ( .A(n967), .B(n966), .ZN(G229) );
  XOR2_X1 U1058 ( .A(KEYINPUT109), .B(KEYINPUT46), .Z(n969) );
  XNOR2_X1 U1059 ( .A(KEYINPUT48), .B(KEYINPUT110), .ZN(n968) );
  XNOR2_X1 U1060 ( .A(n969), .B(n968), .ZN(n971) );
  XNOR2_X1 U1061 ( .A(n971), .B(n970), .ZN(n976) );
  XOR2_X1 U1062 ( .A(G164), .B(n972), .Z(n973) );
  XNOR2_X1 U1063 ( .A(n974), .B(n973), .ZN(n975) );
  XNOR2_X1 U1064 ( .A(n976), .B(n975), .ZN(n994) );
  XNOR2_X1 U1065 ( .A(n977), .B(G162), .ZN(n990) );
  NAND2_X1 U1066 ( .A1(G118), .A2(n978), .ZN(n981) );
  NAND2_X1 U1067 ( .A1(G130), .A2(n979), .ZN(n980) );
  NAND2_X1 U1068 ( .A1(n981), .A2(n980), .ZN(n988) );
  NAND2_X1 U1069 ( .A1(G142), .A2(n982), .ZN(n985) );
  NAND2_X1 U1070 ( .A1(G106), .A2(n983), .ZN(n984) );
  NAND2_X1 U1071 ( .A1(n985), .A2(n984), .ZN(n986) );
  XOR2_X1 U1072 ( .A(KEYINPUT45), .B(n986), .Z(n987) );
  NOR2_X1 U1073 ( .A1(n988), .A2(n987), .ZN(n989) );
  XNOR2_X1 U1074 ( .A(n990), .B(n989), .ZN(n991) );
  XNOR2_X1 U1075 ( .A(n992), .B(n991), .ZN(n993) );
  XNOR2_X1 U1076 ( .A(n994), .B(n993), .ZN(n995) );
  XNOR2_X1 U1077 ( .A(n995), .B(G160), .ZN(n996) );
  NOR2_X1 U1078 ( .A1(G37), .A2(n996), .ZN(G395) );
  XNOR2_X1 U1079 ( .A(G286), .B(n997), .ZN(n1002) );
  XNOR2_X1 U1080 ( .A(G171), .B(n998), .ZN(n1000) );
  XNOR2_X1 U1081 ( .A(n1000), .B(n999), .ZN(n1001) );
  XNOR2_X1 U1082 ( .A(n1002), .B(n1001), .ZN(n1003) );
  NOR2_X1 U1083 ( .A1(G37), .A2(n1003), .ZN(G397) );
  XOR2_X1 U1084 ( .A(G2443), .B(G2430), .Z(n1005) );
  XNOR2_X1 U1085 ( .A(G1348), .B(G2451), .ZN(n1004) );
  XNOR2_X1 U1086 ( .A(n1005), .B(n1004), .ZN(n1012) );
  XOR2_X1 U1087 ( .A(G2438), .B(KEYINPUT105), .Z(n1007) );
  XNOR2_X1 U1088 ( .A(G1341), .B(G2454), .ZN(n1006) );
  XNOR2_X1 U1089 ( .A(n1007), .B(n1006), .ZN(n1008) );
  XOR2_X1 U1090 ( .A(n1008), .B(G2435), .Z(n1010) );
  XNOR2_X1 U1091 ( .A(G2446), .B(G2427), .ZN(n1009) );
  XNOR2_X1 U1092 ( .A(n1010), .B(n1009), .ZN(n1011) );
  XNOR2_X1 U1093 ( .A(n1012), .B(n1011), .ZN(n1013) );
  NAND2_X1 U1094 ( .A1(n1013), .A2(G14), .ZN(n1020) );
  NAND2_X1 U1095 ( .A1(n1020), .A2(G319), .ZN(n1017) );
  NOR2_X1 U1096 ( .A1(G227), .A2(G229), .ZN(n1014) );
  XOR2_X1 U1097 ( .A(KEYINPUT111), .B(n1014), .Z(n1015) );
  XNOR2_X1 U1098 ( .A(n1015), .B(KEYINPUT49), .ZN(n1016) );
  NOR2_X1 U1099 ( .A1(n1017), .A2(n1016), .ZN(n1019) );
  NOR2_X1 U1100 ( .A1(G395), .A2(G397), .ZN(n1018) );
  NAND2_X1 U1101 ( .A1(n1019), .A2(n1018), .ZN(G225) );
  INV_X1 U1102 ( .A(G225), .ZN(G308) );
  INV_X1 U1103 ( .A(G96), .ZN(G221) );
  INV_X1 U1104 ( .A(G69), .ZN(G235) );
  INV_X1 U1105 ( .A(n1020), .ZN(G401) );
endmodule

