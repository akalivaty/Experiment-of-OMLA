

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n294, n295, n296, n297, n298, n299, n300, n301, n302, n303, n304,
         n305, n306, n307, n308, n309, n310, n311, n312, n313, n314, n315,
         n316, n317, n318, n319, n320, n321, n322, n323, n324, n325, n326,
         n327, n328, n329, n330, n331, n332, n333, n334, n335, n336, n337,
         n338, n339, n340, n341, n342, n343, n344, n345, n346, n347, n348,
         n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359,
         n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370,
         n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381,
         n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392,
         n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403,
         n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414,
         n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425,
         n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436,
         n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447,
         n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458,
         n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469,
         n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480,
         n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491,
         n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502,
         n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n513,
         n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
         n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
         n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590,
         n591, n592, n593, n594, n595, n596, n597, n598, n599, n600;

  XNOR2_X1 U326 ( .A(KEYINPUT46), .B(KEYINPUT107), .ZN(n395) );
  XNOR2_X1 U327 ( .A(n377), .B(n376), .ZN(n380) );
  XNOR2_X1 U328 ( .A(n375), .B(n374), .ZN(n376) );
  XNOR2_X1 U329 ( .A(KEYINPUT72), .B(KEYINPUT32), .ZN(n367) );
  XNOR2_X1 U330 ( .A(n445), .B(n367), .ZN(n370) );
  XNOR2_X1 U331 ( .A(n396), .B(n395), .ZN(n398) );
  INV_X1 U332 ( .A(KEYINPUT54), .ZN(n423) );
  XNOR2_X1 U333 ( .A(n423), .B(KEYINPUT118), .ZN(n424) );
  XNOR2_X1 U334 ( .A(n356), .B(n355), .ZN(n357) );
  XNOR2_X1 U335 ( .A(n358), .B(n357), .ZN(n361) );
  XNOR2_X1 U336 ( .A(n363), .B(n362), .ZN(n585) );
  XNOR2_X1 U337 ( .A(n585), .B(KEYINPUT36), .ZN(n516) );
  XNOR2_X1 U338 ( .A(n462), .B(KEYINPUT123), .ZN(n598) );
  XNOR2_X1 U339 ( .A(n468), .B(n467), .ZN(n469) );
  XNOR2_X1 U340 ( .A(n472), .B(n471), .ZN(n473) );
  XNOR2_X1 U341 ( .A(n470), .B(n469), .ZN(G1355GAT) );
  XNOR2_X1 U342 ( .A(n474), .B(n473), .ZN(G1353GAT) );
  XOR2_X1 U343 ( .A(G148GAT), .B(KEYINPUT6), .Z(n295) );
  XNOR2_X1 U344 ( .A(KEYINPUT5), .B(KEYINPUT4), .ZN(n294) );
  XNOR2_X1 U345 ( .A(n295), .B(n294), .ZN(n309) );
  XOR2_X1 U346 ( .A(KEYINPUT1), .B(G85GAT), .Z(n297) );
  XNOR2_X1 U347 ( .A(G29GAT), .B(G1GAT), .ZN(n296) );
  XNOR2_X1 U348 ( .A(n297), .B(n296), .ZN(n301) );
  XOR2_X1 U349 ( .A(KEYINPUT85), .B(G57GAT), .Z(n299) );
  XNOR2_X1 U350 ( .A(G141GAT), .B(G120GAT), .ZN(n298) );
  XNOR2_X1 U351 ( .A(n299), .B(n298), .ZN(n300) );
  XOR2_X1 U352 ( .A(n301), .B(n300), .Z(n307) );
  XNOR2_X1 U353 ( .A(G155GAT), .B(KEYINPUT3), .ZN(n302) );
  XNOR2_X1 U354 ( .A(n302), .B(KEYINPUT2), .ZN(n432) );
  XOR2_X1 U355 ( .A(n432), .B(G162GAT), .Z(n304) );
  NAND2_X1 U356 ( .A1(G225GAT), .A2(G233GAT), .ZN(n303) );
  XNOR2_X1 U357 ( .A(n304), .B(n303), .ZN(n305) );
  XNOR2_X1 U358 ( .A(G134GAT), .B(n305), .ZN(n306) );
  XNOR2_X1 U359 ( .A(n307), .B(n306), .ZN(n308) );
  XNOR2_X1 U360 ( .A(n309), .B(n308), .ZN(n313) );
  XOR2_X1 U361 ( .A(KEYINPUT77), .B(KEYINPUT0), .Z(n311) );
  XNOR2_X1 U362 ( .A(KEYINPUT78), .B(G127GAT), .ZN(n310) );
  XNOR2_X1 U363 ( .A(n311), .B(n310), .ZN(n312) );
  XNOR2_X1 U364 ( .A(G113GAT), .B(n312), .ZN(n459) );
  XNOR2_X1 U365 ( .A(n313), .B(n459), .ZN(n572) );
  XOR2_X1 U366 ( .A(KEYINPUT30), .B(KEYINPUT69), .Z(n315) );
  XNOR2_X1 U367 ( .A(G50GAT), .B(G113GAT), .ZN(n314) );
  XNOR2_X1 U368 ( .A(n315), .B(n314), .ZN(n319) );
  XOR2_X1 U369 ( .A(KEYINPUT29), .B(KEYINPUT68), .Z(n317) );
  XNOR2_X1 U370 ( .A(KEYINPUT67), .B(G197GAT), .ZN(n316) );
  XNOR2_X1 U371 ( .A(n317), .B(n316), .ZN(n318) );
  XNOR2_X1 U372 ( .A(n319), .B(n318), .ZN(n329) );
  XNOR2_X1 U373 ( .A(G29GAT), .B(KEYINPUT7), .ZN(n320) );
  XNOR2_X1 U374 ( .A(n320), .B(KEYINPUT8), .ZN(n348) );
  XOR2_X1 U375 ( .A(n348), .B(KEYINPUT70), .Z(n322) );
  NAND2_X1 U376 ( .A1(G229GAT), .A2(G233GAT), .ZN(n321) );
  XNOR2_X1 U377 ( .A(n322), .B(n321), .ZN(n323) );
  XOR2_X1 U378 ( .A(G169GAT), .B(G8GAT), .Z(n413) );
  XNOR2_X1 U379 ( .A(n323), .B(n413), .ZN(n327) );
  XOR2_X1 U380 ( .A(G43GAT), .B(G36GAT), .Z(n325) );
  XOR2_X1 U381 ( .A(G141GAT), .B(G22GAT), .Z(n438) );
  XOR2_X1 U382 ( .A(G1GAT), .B(G15GAT), .Z(n332) );
  XNOR2_X1 U383 ( .A(n438), .B(n332), .ZN(n324) );
  XNOR2_X1 U384 ( .A(n325), .B(n324), .ZN(n326) );
  XNOR2_X1 U385 ( .A(n327), .B(n326), .ZN(n328) );
  XNOR2_X1 U386 ( .A(n329), .B(n328), .ZN(n588) );
  XOR2_X1 U387 ( .A(KEYINPUT75), .B(KEYINPUT12), .Z(n331) );
  XNOR2_X1 U388 ( .A(KEYINPUT15), .B(KEYINPUT14), .ZN(n330) );
  XNOR2_X1 U389 ( .A(n331), .B(n330), .ZN(n336) );
  XOR2_X1 U390 ( .A(G57GAT), .B(KEYINPUT13), .Z(n369) );
  XOR2_X1 U391 ( .A(n369), .B(G155GAT), .Z(n334) );
  XNOR2_X1 U392 ( .A(n332), .B(G127GAT), .ZN(n333) );
  XNOR2_X1 U393 ( .A(n334), .B(n333), .ZN(n335) );
  XOR2_X1 U394 ( .A(n336), .B(n335), .Z(n338) );
  NAND2_X1 U395 ( .A1(G231GAT), .A2(G233GAT), .ZN(n337) );
  XNOR2_X1 U396 ( .A(n338), .B(n337), .ZN(n346) );
  XOR2_X1 U397 ( .A(G78GAT), .B(G64GAT), .Z(n340) );
  XNOR2_X1 U398 ( .A(G8GAT), .B(G71GAT), .ZN(n339) );
  XNOR2_X1 U399 ( .A(n340), .B(n339), .ZN(n344) );
  XOR2_X1 U400 ( .A(G211GAT), .B(KEYINPUT76), .Z(n342) );
  XNOR2_X1 U401 ( .A(G22GAT), .B(G183GAT), .ZN(n341) );
  XNOR2_X1 U402 ( .A(n342), .B(n341), .ZN(n343) );
  XOR2_X1 U403 ( .A(n344), .B(n343), .Z(n345) );
  XNOR2_X1 U404 ( .A(n346), .B(n345), .ZN(n599) );
  XNOR2_X1 U405 ( .A(G99GAT), .B(G85GAT), .ZN(n347) );
  XNOR2_X1 U406 ( .A(n347), .B(KEYINPUT71), .ZN(n378) );
  XNOR2_X1 U407 ( .A(n348), .B(n378), .ZN(n363) );
  XOR2_X1 U408 ( .A(KEYINPUT73), .B(KEYINPUT11), .Z(n350) );
  XNOR2_X1 U409 ( .A(G106GAT), .B(G92GAT), .ZN(n349) );
  XNOR2_X1 U410 ( .A(n350), .B(n349), .ZN(n354) );
  XOR2_X1 U411 ( .A(KEYINPUT9), .B(G218GAT), .Z(n352) );
  XOR2_X1 U412 ( .A(G43GAT), .B(G134GAT), .Z(n446) );
  XOR2_X1 U413 ( .A(G50GAT), .B(G162GAT), .Z(n437) );
  XNOR2_X1 U414 ( .A(n446), .B(n437), .ZN(n351) );
  XNOR2_X1 U415 ( .A(n352), .B(n351), .ZN(n353) );
  XOR2_X1 U416 ( .A(n354), .B(n353), .Z(n358) );
  NAND2_X1 U417 ( .A1(G232GAT), .A2(G233GAT), .ZN(n356) );
  INV_X1 U418 ( .A(KEYINPUT10), .ZN(n355) );
  XNOR2_X1 U419 ( .A(G36GAT), .B(G190GAT), .ZN(n359) );
  XNOR2_X1 U420 ( .A(n359), .B(KEYINPUT74), .ZN(n407) );
  XNOR2_X1 U421 ( .A(n407), .B(KEYINPUT66), .ZN(n360) );
  XNOR2_X1 U422 ( .A(n361), .B(n360), .ZN(n362) );
  NAND2_X1 U423 ( .A1(n599), .A2(n516), .ZN(n366) );
  XNOR2_X1 U424 ( .A(KEYINPUT108), .B(KEYINPUT45), .ZN(n364) );
  XNOR2_X1 U425 ( .A(n364), .B(KEYINPUT65), .ZN(n365) );
  XNOR2_X1 U426 ( .A(n366), .B(n365), .ZN(n391) );
  XOR2_X1 U427 ( .A(G120GAT), .B(G71GAT), .Z(n445) );
  INV_X1 U428 ( .A(n370), .ZN(n368) );
  NAND2_X1 U429 ( .A1(n368), .A2(n369), .ZN(n373) );
  INV_X1 U430 ( .A(n369), .ZN(n371) );
  NAND2_X1 U431 ( .A1(n371), .A2(n370), .ZN(n372) );
  NAND2_X1 U432 ( .A1(n373), .A2(n372), .ZN(n377) );
  NAND2_X1 U433 ( .A1(G230GAT), .A2(G233GAT), .ZN(n375) );
  INV_X1 U434 ( .A(KEYINPUT31), .ZN(n374) );
  XNOR2_X1 U435 ( .A(n378), .B(KEYINPUT33), .ZN(n379) );
  XNOR2_X1 U436 ( .A(n380), .B(n379), .ZN(n384) );
  INV_X1 U437 ( .A(n384), .ZN(n383) );
  XOR2_X1 U438 ( .A(G64GAT), .B(G204GAT), .Z(n382) );
  XNOR2_X1 U439 ( .A(G176GAT), .B(G92GAT), .ZN(n381) );
  XNOR2_X1 U440 ( .A(n382), .B(n381), .ZN(n406) );
  NAND2_X1 U441 ( .A1(n383), .A2(n406), .ZN(n387) );
  INV_X1 U442 ( .A(n406), .ZN(n385) );
  NAND2_X1 U443 ( .A1(n385), .A2(n384), .ZN(n386) );
  NAND2_X1 U444 ( .A1(n387), .A2(n386), .ZN(n390) );
  XNOR2_X1 U445 ( .A(G148GAT), .B(G106GAT), .ZN(n388) );
  XNOR2_X1 U446 ( .A(n388), .B(G78GAT), .ZN(n435) );
  INV_X1 U447 ( .A(n435), .ZN(n389) );
  XNOR2_X1 U448 ( .A(n390), .B(n389), .ZN(n394) );
  INV_X1 U449 ( .A(n394), .ZN(n487) );
  NAND2_X1 U450 ( .A1(n391), .A2(n487), .ZN(n392) );
  NOR2_X1 U451 ( .A1(n588), .A2(n392), .ZN(n393) );
  XOR2_X1 U452 ( .A(KEYINPUT109), .B(n393), .Z(n402) );
  XNOR2_X1 U453 ( .A(KEYINPUT41), .B(n394), .ZN(n578) );
  INV_X1 U454 ( .A(n588), .ZN(n574) );
  NOR2_X1 U455 ( .A1(n578), .A2(n574), .ZN(n396) );
  NOR2_X1 U456 ( .A1(n585), .A2(n599), .ZN(n397) );
  AND2_X1 U457 ( .A1(n398), .A2(n397), .ZN(n400) );
  INV_X1 U458 ( .A(KEYINPUT47), .ZN(n399) );
  XNOR2_X1 U459 ( .A(n400), .B(n399), .ZN(n401) );
  NOR2_X1 U460 ( .A1(n402), .A2(n401), .ZN(n403) );
  XNOR2_X1 U461 ( .A(n403), .B(KEYINPUT48), .ZN(n555) );
  XOR2_X1 U462 ( .A(KEYINPUT18), .B(KEYINPUT17), .Z(n405) );
  XNOR2_X1 U463 ( .A(G183GAT), .B(KEYINPUT19), .ZN(n404) );
  XNOR2_X1 U464 ( .A(n405), .B(n404), .ZN(n450) );
  XNOR2_X1 U465 ( .A(n450), .B(n406), .ZN(n411) );
  XOR2_X1 U466 ( .A(n407), .B(KEYINPUT86), .Z(n409) );
  NAND2_X1 U467 ( .A1(G226GAT), .A2(G233GAT), .ZN(n408) );
  XNOR2_X1 U468 ( .A(n409), .B(n408), .ZN(n410) );
  XNOR2_X1 U469 ( .A(n411), .B(n410), .ZN(n412) );
  XOR2_X1 U470 ( .A(n412), .B(KEYINPUT87), .Z(n415) );
  XNOR2_X1 U471 ( .A(n413), .B(KEYINPUT75), .ZN(n414) );
  XNOR2_X1 U472 ( .A(n415), .B(n414), .ZN(n421) );
  XNOR2_X1 U473 ( .A(G211GAT), .B(KEYINPUT21), .ZN(n416) );
  XNOR2_X1 U474 ( .A(n416), .B(KEYINPUT83), .ZN(n417) );
  XOR2_X1 U475 ( .A(n417), .B(KEYINPUT82), .Z(n419) );
  XNOR2_X1 U476 ( .A(G197GAT), .B(G218GAT), .ZN(n418) );
  XNOR2_X1 U477 ( .A(n419), .B(n418), .ZN(n431) );
  INV_X1 U478 ( .A(n431), .ZN(n420) );
  XNOR2_X1 U479 ( .A(n421), .B(n420), .ZN(n546) );
  XNOR2_X1 U480 ( .A(n546), .B(KEYINPUT117), .ZN(n422) );
  NOR2_X1 U481 ( .A1(n555), .A2(n422), .ZN(n425) );
  XNOR2_X1 U482 ( .A(n425), .B(n424), .ZN(n426) );
  NOR2_X1 U483 ( .A1(n572), .A2(n426), .ZN(n427) );
  XNOR2_X1 U484 ( .A(KEYINPUT64), .B(n427), .ZN(n480) );
  XOR2_X1 U485 ( .A(KEYINPUT22), .B(KEYINPUT23), .Z(n429) );
  XNOR2_X1 U486 ( .A(G204GAT), .B(KEYINPUT84), .ZN(n428) );
  XNOR2_X1 U487 ( .A(n429), .B(n428), .ZN(n430) );
  XNOR2_X1 U488 ( .A(n431), .B(n430), .ZN(n442) );
  XOR2_X1 U489 ( .A(n432), .B(KEYINPUT24), .Z(n434) );
  NAND2_X1 U490 ( .A1(G228GAT), .A2(G233GAT), .ZN(n433) );
  XNOR2_X1 U491 ( .A(n434), .B(n433), .ZN(n436) );
  XOR2_X1 U492 ( .A(n436), .B(n435), .Z(n440) );
  XNOR2_X1 U493 ( .A(n438), .B(n437), .ZN(n439) );
  XNOR2_X1 U494 ( .A(n440), .B(n439), .ZN(n441) );
  XNOR2_X1 U495 ( .A(n442), .B(n441), .ZN(n497) );
  XOR2_X1 U496 ( .A(KEYINPUT80), .B(KEYINPUT81), .Z(n444) );
  XNOR2_X1 U497 ( .A(G15GAT), .B(KEYINPUT79), .ZN(n443) );
  XNOR2_X1 U498 ( .A(n444), .B(n443), .ZN(n457) );
  XOR2_X1 U499 ( .A(G99GAT), .B(G190GAT), .Z(n448) );
  XNOR2_X1 U500 ( .A(n446), .B(n445), .ZN(n447) );
  XNOR2_X1 U501 ( .A(n448), .B(n447), .ZN(n449) );
  XOR2_X1 U502 ( .A(n449), .B(G176GAT), .Z(n455) );
  XOR2_X1 U503 ( .A(n450), .B(KEYINPUT20), .Z(n452) );
  NAND2_X1 U504 ( .A1(G227GAT), .A2(G233GAT), .ZN(n451) );
  XNOR2_X1 U505 ( .A(n452), .B(n451), .ZN(n453) );
  XNOR2_X1 U506 ( .A(G169GAT), .B(n453), .ZN(n454) );
  XNOR2_X1 U507 ( .A(n455), .B(n454), .ZN(n456) );
  XOR2_X1 U508 ( .A(n457), .B(n456), .Z(n458) );
  XNOR2_X1 U509 ( .A(n459), .B(n458), .ZN(n482) );
  INV_X1 U510 ( .A(n482), .ZN(n594) );
  NOR2_X1 U511 ( .A1(n497), .A2(n594), .ZN(n461) );
  XNOR2_X1 U512 ( .A(KEYINPUT90), .B(KEYINPUT26), .ZN(n460) );
  XNOR2_X1 U513 ( .A(n461), .B(n460), .ZN(n491) );
  NAND2_X1 U514 ( .A1(n480), .A2(n491), .ZN(n462) );
  NAND2_X1 U515 ( .A1(n598), .A2(n588), .ZN(n466) );
  XOR2_X1 U516 ( .A(G197GAT), .B(KEYINPUT124), .Z(n464) );
  XNOR2_X1 U517 ( .A(KEYINPUT60), .B(KEYINPUT59), .ZN(n463) );
  XNOR2_X1 U518 ( .A(n464), .B(n463), .ZN(n465) );
  XNOR2_X1 U519 ( .A(n466), .B(n465), .ZN(G1352GAT) );
  NAND2_X1 U520 ( .A1(n598), .A2(n516), .ZN(n470) );
  XOR2_X1 U521 ( .A(KEYINPUT62), .B(KEYINPUT127), .Z(n468) );
  XNOR2_X1 U522 ( .A(G218GAT), .B(KEYINPUT126), .ZN(n467) );
  NAND2_X1 U523 ( .A1(n598), .A2(n394), .ZN(n474) );
  XOR2_X1 U524 ( .A(KEYINPUT61), .B(KEYINPUT125), .Z(n472) );
  INV_X1 U525 ( .A(G204GAT), .ZN(n471) );
  XOR2_X1 U526 ( .A(KEYINPUT56), .B(KEYINPUT121), .Z(n476) );
  XNOR2_X1 U527 ( .A(KEYINPUT119), .B(KEYINPUT120), .ZN(n475) );
  XNOR2_X1 U528 ( .A(n476), .B(n475), .ZN(n477) );
  XOR2_X1 U529 ( .A(n477), .B(KEYINPUT122), .Z(n479) );
  XNOR2_X1 U530 ( .A(G176GAT), .B(KEYINPUT57), .ZN(n478) );
  XOR2_X1 U531 ( .A(n479), .B(n478), .Z(n484) );
  XOR2_X1 U532 ( .A(KEYINPUT100), .B(n578), .Z(n560) );
  AND2_X1 U533 ( .A1(n497), .A2(n480), .ZN(n481) );
  XNOR2_X1 U534 ( .A(KEYINPUT55), .B(n481), .ZN(n593) );
  NOR2_X1 U535 ( .A1(n482), .A2(n593), .ZN(n590) );
  NAND2_X1 U536 ( .A1(n560), .A2(n590), .ZN(n483) );
  XNOR2_X1 U537 ( .A(n484), .B(n483), .ZN(G1349GAT) );
  XNOR2_X1 U538 ( .A(G1GAT), .B(KEYINPUT34), .ZN(n485) );
  XNOR2_X1 U539 ( .A(n485), .B(KEYINPUT94), .ZN(n486) );
  XOR2_X1 U540 ( .A(KEYINPUT95), .B(n486), .Z(n507) );
  NAND2_X1 U541 ( .A1(n588), .A2(n487), .ZN(n520) );
  INV_X1 U542 ( .A(n599), .ZN(n581) );
  NOR2_X1 U543 ( .A1(n585), .A2(n581), .ZN(n488) );
  XNOR2_X1 U544 ( .A(n488), .B(KEYINPUT16), .ZN(n504) );
  NAND2_X1 U545 ( .A1(n546), .A2(n594), .ZN(n489) );
  NAND2_X1 U546 ( .A1(n497), .A2(n489), .ZN(n490) );
  XNOR2_X1 U547 ( .A(KEYINPUT25), .B(n490), .ZN(n493) );
  XNOR2_X1 U548 ( .A(n546), .B(KEYINPUT27), .ZN(n496) );
  NAND2_X1 U549 ( .A1(n491), .A2(n496), .ZN(n571) );
  XNOR2_X1 U550 ( .A(KEYINPUT91), .B(n571), .ZN(n492) );
  NOR2_X1 U551 ( .A1(n493), .A2(n492), .ZN(n494) );
  NOR2_X1 U552 ( .A1(n494), .A2(n572), .ZN(n495) );
  XOR2_X1 U553 ( .A(KEYINPUT92), .B(n495), .Z(n503) );
  INV_X1 U554 ( .A(n496), .ZN(n499) );
  XNOR2_X1 U555 ( .A(n497), .B(KEYINPUT28), .ZN(n512) );
  NAND2_X1 U556 ( .A1(n572), .A2(n512), .ZN(n498) );
  NOR2_X1 U557 ( .A1(n499), .A2(n498), .ZN(n556) );
  XOR2_X1 U558 ( .A(n556), .B(KEYINPUT88), .Z(n500) );
  NOR2_X1 U559 ( .A1(n594), .A2(n500), .ZN(n501) );
  XNOR2_X1 U560 ( .A(KEYINPUT89), .B(n501), .ZN(n502) );
  NAND2_X1 U561 ( .A1(n503), .A2(n502), .ZN(n515) );
  NAND2_X1 U562 ( .A1(n504), .A2(n515), .ZN(n505) );
  XOR2_X1 U563 ( .A(KEYINPUT93), .B(n505), .Z(n531) );
  NOR2_X1 U564 ( .A1(n520), .A2(n531), .ZN(n513) );
  NAND2_X1 U565 ( .A1(n513), .A2(n572), .ZN(n506) );
  XNOR2_X1 U566 ( .A(n507), .B(n506), .ZN(G1324GAT) );
  NAND2_X1 U567 ( .A1(n513), .A2(n546), .ZN(n508) );
  XNOR2_X1 U568 ( .A(n508), .B(G8GAT), .ZN(G1325GAT) );
  XOR2_X1 U569 ( .A(KEYINPUT35), .B(KEYINPUT96), .Z(n510) );
  NAND2_X1 U570 ( .A1(n513), .A2(n594), .ZN(n509) );
  XNOR2_X1 U571 ( .A(n510), .B(n509), .ZN(n511) );
  XNOR2_X1 U572 ( .A(G15GAT), .B(n511), .ZN(G1326GAT) );
  INV_X1 U573 ( .A(n512), .ZN(n551) );
  NAND2_X1 U574 ( .A1(n513), .A2(n551), .ZN(n514) );
  XNOR2_X1 U575 ( .A(n514), .B(G22GAT), .ZN(G1327GAT) );
  XOR2_X1 U576 ( .A(G29GAT), .B(KEYINPUT39), .Z(n524) );
  NAND2_X1 U577 ( .A1(n516), .A2(n515), .ZN(n517) );
  NOR2_X1 U578 ( .A1(n599), .A2(n517), .ZN(n519) );
  XOR2_X1 U579 ( .A(KEYINPUT97), .B(KEYINPUT37), .Z(n518) );
  XNOR2_X1 U580 ( .A(n519), .B(n518), .ZN(n542) );
  NOR2_X1 U581 ( .A1(n542), .A2(n520), .ZN(n522) );
  XNOR2_X1 U582 ( .A(KEYINPUT38), .B(KEYINPUT98), .ZN(n521) );
  XNOR2_X1 U583 ( .A(n522), .B(n521), .ZN(n529) );
  NAND2_X1 U584 ( .A1(n529), .A2(n572), .ZN(n523) );
  XNOR2_X1 U585 ( .A(n524), .B(n523), .ZN(G1328GAT) );
  XOR2_X1 U586 ( .A(G36GAT), .B(KEYINPUT99), .Z(n526) );
  NAND2_X1 U587 ( .A1(n529), .A2(n546), .ZN(n525) );
  XNOR2_X1 U588 ( .A(n526), .B(n525), .ZN(G1329GAT) );
  NAND2_X1 U589 ( .A1(n594), .A2(n529), .ZN(n527) );
  XNOR2_X1 U590 ( .A(n527), .B(KEYINPUT40), .ZN(n528) );
  XNOR2_X1 U591 ( .A(G43GAT), .B(n528), .ZN(G1330GAT) );
  NAND2_X1 U592 ( .A1(n529), .A2(n551), .ZN(n530) );
  XNOR2_X1 U593 ( .A(n530), .B(G50GAT), .ZN(G1331GAT) );
  XOR2_X1 U594 ( .A(KEYINPUT42), .B(KEYINPUT101), .Z(n533) );
  NAND2_X1 U595 ( .A1(n574), .A2(n560), .ZN(n541) );
  NOR2_X1 U596 ( .A1(n531), .A2(n541), .ZN(n538) );
  NAND2_X1 U597 ( .A1(n538), .A2(n572), .ZN(n532) );
  XNOR2_X1 U598 ( .A(n533), .B(n532), .ZN(n534) );
  XNOR2_X1 U599 ( .A(G57GAT), .B(n534), .ZN(G1332GAT) );
  NAND2_X1 U600 ( .A1(n538), .A2(n546), .ZN(n535) );
  XNOR2_X1 U601 ( .A(n535), .B(G64GAT), .ZN(G1333GAT) );
  NAND2_X1 U602 ( .A1(n594), .A2(n538), .ZN(n536) );
  XNOR2_X1 U603 ( .A(n536), .B(KEYINPUT102), .ZN(n537) );
  XNOR2_X1 U604 ( .A(G71GAT), .B(n537), .ZN(G1334GAT) );
  XOR2_X1 U605 ( .A(G78GAT), .B(KEYINPUT43), .Z(n540) );
  NAND2_X1 U606 ( .A1(n538), .A2(n551), .ZN(n539) );
  XNOR2_X1 U607 ( .A(n540), .B(n539), .ZN(G1335GAT) );
  XOR2_X1 U608 ( .A(KEYINPUT103), .B(KEYINPUT104), .Z(n544) );
  NOR2_X1 U609 ( .A1(n542), .A2(n541), .ZN(n552) );
  NAND2_X1 U610 ( .A1(n552), .A2(n572), .ZN(n543) );
  XNOR2_X1 U611 ( .A(n544), .B(n543), .ZN(n545) );
  XNOR2_X1 U612 ( .A(G85GAT), .B(n545), .ZN(G1336GAT) );
  XOR2_X1 U613 ( .A(KEYINPUT105), .B(KEYINPUT106), .Z(n548) );
  NAND2_X1 U614 ( .A1(n552), .A2(n546), .ZN(n547) );
  XNOR2_X1 U615 ( .A(n548), .B(n547), .ZN(n549) );
  XNOR2_X1 U616 ( .A(G92GAT), .B(n549), .ZN(G1337GAT) );
  NAND2_X1 U617 ( .A1(n594), .A2(n552), .ZN(n550) );
  XNOR2_X1 U618 ( .A(n550), .B(G99GAT), .ZN(G1338GAT) );
  NAND2_X1 U619 ( .A1(n552), .A2(n551), .ZN(n553) );
  XNOR2_X1 U620 ( .A(n553), .B(KEYINPUT44), .ZN(n554) );
  XNOR2_X1 U621 ( .A(G106GAT), .B(n554), .ZN(G1339GAT) );
  NAND2_X1 U622 ( .A1(n556), .A2(n594), .ZN(n557) );
  NOR2_X1 U623 ( .A1(n555), .A2(n557), .ZN(n566) );
  NAND2_X1 U624 ( .A1(n566), .A2(n588), .ZN(n558) );
  XNOR2_X1 U625 ( .A(n558), .B(KEYINPUT110), .ZN(n559) );
  XNOR2_X1 U626 ( .A(G113GAT), .B(n559), .ZN(G1340GAT) );
  XOR2_X1 U627 ( .A(KEYINPUT49), .B(KEYINPUT111), .Z(n562) );
  NAND2_X1 U628 ( .A1(n566), .A2(n560), .ZN(n561) );
  XNOR2_X1 U629 ( .A(n562), .B(n561), .ZN(n563) );
  XOR2_X1 U630 ( .A(G120GAT), .B(n563), .Z(G1341GAT) );
  NAND2_X1 U631 ( .A1(n599), .A2(n566), .ZN(n564) );
  XNOR2_X1 U632 ( .A(n564), .B(KEYINPUT50), .ZN(n565) );
  XNOR2_X1 U633 ( .A(G127GAT), .B(n565), .ZN(G1342GAT) );
  XOR2_X1 U634 ( .A(KEYINPUT112), .B(KEYINPUT51), .Z(n568) );
  NAND2_X1 U635 ( .A1(n566), .A2(n585), .ZN(n567) );
  XNOR2_X1 U636 ( .A(n568), .B(n567), .ZN(n570) );
  XOR2_X1 U637 ( .A(G134GAT), .B(KEYINPUT113), .Z(n569) );
  XNOR2_X1 U638 ( .A(n570), .B(n569), .ZN(G1343GAT) );
  NOR2_X1 U639 ( .A1(n555), .A2(n571), .ZN(n573) );
  NAND2_X1 U640 ( .A1(n573), .A2(n572), .ZN(n586) );
  NOR2_X1 U641 ( .A1(n574), .A2(n586), .ZN(n575) );
  XOR2_X1 U642 ( .A(G141GAT), .B(n575), .Z(G1344GAT) );
  XOR2_X1 U643 ( .A(KEYINPUT53), .B(KEYINPUT52), .Z(n577) );
  XNOR2_X1 U644 ( .A(G148GAT), .B(KEYINPUT114), .ZN(n576) );
  XNOR2_X1 U645 ( .A(n577), .B(n576), .ZN(n580) );
  NOR2_X1 U646 ( .A1(n578), .A2(n586), .ZN(n579) );
  XOR2_X1 U647 ( .A(n580), .B(n579), .Z(G1345GAT) );
  NOR2_X1 U648 ( .A1(n581), .A2(n586), .ZN(n583) );
  XNOR2_X1 U649 ( .A(KEYINPUT115), .B(KEYINPUT116), .ZN(n582) );
  XNOR2_X1 U650 ( .A(n583), .B(n582), .ZN(n584) );
  XNOR2_X1 U651 ( .A(G155GAT), .B(n584), .ZN(G1346GAT) );
  INV_X1 U652 ( .A(n585), .ZN(n592) );
  NOR2_X1 U653 ( .A1(n592), .A2(n586), .ZN(n587) );
  XOR2_X1 U654 ( .A(G162GAT), .B(n587), .Z(G1347GAT) );
  NAND2_X1 U655 ( .A1(n590), .A2(n588), .ZN(n589) );
  XNOR2_X1 U656 ( .A(n589), .B(G169GAT), .ZN(G1348GAT) );
  NAND2_X1 U657 ( .A1(n599), .A2(n590), .ZN(n591) );
  XNOR2_X1 U658 ( .A(n591), .B(G183GAT), .ZN(G1350GAT) );
  NOR2_X1 U659 ( .A1(n593), .A2(n592), .ZN(n595) );
  NAND2_X1 U660 ( .A1(n595), .A2(n594), .ZN(n596) );
  XNOR2_X1 U661 ( .A(n596), .B(KEYINPUT58), .ZN(n597) );
  XNOR2_X1 U662 ( .A(G190GAT), .B(n597), .ZN(G1351GAT) );
  NAND2_X1 U663 ( .A1(n599), .A2(n598), .ZN(n600) );
  XNOR2_X1 U664 ( .A(n600), .B(G211GAT), .ZN(G1354GAT) );
endmodule

