//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 1 0 1 1 1 1 0 1 1 0 1 1 1 0 0 1 1 1 0 1 0 1 1 1 1 1 1 0 0 0 0 1 0 1 0 0 0 0 0 0 0 1 1 1 0 1 1 0 1 1 0 0 1 0 1 0 1 0 0 0 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:28:02 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n703, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n712, new_n713, new_n714,
    new_n715, new_n716, new_n717, new_n718, new_n719, new_n720, new_n721,
    new_n722, new_n723, new_n724, new_n725, new_n726, new_n727, new_n729,
    new_n730, new_n731, new_n732, new_n733, new_n734, new_n735, new_n736,
    new_n737, new_n738, new_n739, new_n740, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n758, new_n759,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n799, new_n800, new_n801, new_n802, new_n803,
    new_n804, new_n805, new_n806, new_n807, new_n808, new_n809, new_n810,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n935, new_n936, new_n937, new_n938,
    new_n939, new_n940, new_n941, new_n942, new_n943, new_n944, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n976,
    new_n977, new_n978, new_n979, new_n980, new_n981, new_n982, new_n983,
    new_n984, new_n985, new_n986, new_n988, new_n989, new_n990, new_n991,
    new_n992, new_n993, new_n994, new_n995, new_n996, new_n997, new_n998,
    new_n999, new_n1000, new_n1001, new_n1002, new_n1004, new_n1005,
    new_n1006, new_n1007, new_n1008, new_n1009, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1017, new_n1018,
    new_n1019, new_n1020, new_n1021, new_n1022, new_n1023, new_n1024,
    new_n1025, new_n1026, new_n1027, new_n1028, new_n1029, new_n1030,
    new_n1031, new_n1032, new_n1033, new_n1034, new_n1035, new_n1036,
    new_n1037, new_n1038, new_n1039, new_n1040, new_n1042, new_n1043,
    new_n1044, new_n1045, new_n1046, new_n1047, new_n1048, new_n1049,
    new_n1050, new_n1051, new_n1052, new_n1053, new_n1054, new_n1055,
    new_n1056, new_n1057;
  INV_X1    g000(.A(G217), .ZN(new_n187));
  XOR2_X1   g001(.A(KEYINPUT77), .B(G902), .Z(new_n188));
  AOI21_X1  g002(.A(new_n187), .B1(new_n188), .B2(G234), .ZN(new_n189));
  XNOR2_X1  g003(.A(KEYINPUT78), .B(G125), .ZN(new_n190));
  INV_X1    g004(.A(KEYINPUT16), .ZN(new_n191));
  INV_X1    g005(.A(G140), .ZN(new_n192));
  NAND3_X1  g006(.A1(new_n190), .A2(new_n191), .A3(new_n192), .ZN(new_n193));
  NOR2_X1   g007(.A1(G125), .A2(G140), .ZN(new_n194));
  AOI21_X1  g008(.A(new_n194), .B1(new_n190), .B2(G140), .ZN(new_n195));
  OAI21_X1  g009(.A(new_n193), .B1(new_n195), .B2(new_n191), .ZN(new_n196));
  INV_X1    g010(.A(G146), .ZN(new_n197));
  OR2_X1    g011(.A1(new_n196), .A2(new_n197), .ZN(new_n198));
  XNOR2_X1  g012(.A(G125), .B(G140), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n199), .A2(new_n197), .ZN(new_n200));
  INV_X1    g014(.A(G128), .ZN(new_n201));
  NOR2_X1   g015(.A1(new_n201), .A2(G119), .ZN(new_n202));
  INV_X1    g016(.A(KEYINPUT70), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n203), .A2(new_n201), .ZN(new_n204));
  NAND2_X1  g018(.A1(KEYINPUT70), .A2(G128), .ZN(new_n205));
  AND2_X1   g019(.A1(new_n204), .A2(new_n205), .ZN(new_n206));
  AOI21_X1  g020(.A(new_n202), .B1(new_n206), .B2(G119), .ZN(new_n207));
  INV_X1    g021(.A(new_n207), .ZN(new_n208));
  INV_X1    g022(.A(KEYINPUT79), .ZN(new_n209));
  XNOR2_X1  g023(.A(KEYINPUT24), .B(G110), .ZN(new_n210));
  NAND3_X1  g024(.A1(new_n208), .A2(new_n209), .A3(new_n210), .ZN(new_n211));
  INV_X1    g025(.A(G110), .ZN(new_n212));
  AOI21_X1  g026(.A(KEYINPUT23), .B1(new_n201), .B2(G119), .ZN(new_n213));
  NOR2_X1   g027(.A1(new_n213), .A2(new_n202), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n206), .A2(G119), .ZN(new_n215));
  INV_X1    g029(.A(KEYINPUT23), .ZN(new_n216));
  OAI211_X1 g030(.A(new_n212), .B(new_n214), .C1(new_n215), .C2(new_n216), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n211), .A2(new_n217), .ZN(new_n218));
  AOI21_X1  g032(.A(new_n209), .B1(new_n208), .B2(new_n210), .ZN(new_n219));
  OAI211_X1 g033(.A(new_n198), .B(new_n200), .C1(new_n218), .C2(new_n219), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n196), .A2(new_n197), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n198), .A2(new_n221), .ZN(new_n222));
  OAI21_X1  g036(.A(new_n214), .B1(new_n215), .B2(new_n216), .ZN(new_n223));
  INV_X1    g037(.A(new_n210), .ZN(new_n224));
  AOI22_X1  g038(.A1(new_n223), .A2(G110), .B1(new_n207), .B2(new_n224), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n222), .A2(new_n225), .ZN(new_n226));
  INV_X1    g040(.A(KEYINPUT80), .ZN(new_n227));
  NAND3_X1  g041(.A1(new_n220), .A2(new_n226), .A3(new_n227), .ZN(new_n228));
  XNOR2_X1  g042(.A(KEYINPUT22), .B(G137), .ZN(new_n229));
  INV_X1    g043(.A(G953), .ZN(new_n230));
  AND3_X1   g044(.A1(new_n230), .A2(G221), .A3(G234), .ZN(new_n231));
  XOR2_X1   g045(.A(new_n229), .B(new_n231), .Z(new_n232));
  INV_X1    g046(.A(new_n232), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n228), .A2(new_n233), .ZN(new_n234));
  INV_X1    g048(.A(new_n234), .ZN(new_n235));
  AOI21_X1  g049(.A(new_n227), .B1(new_n220), .B2(new_n226), .ZN(new_n236));
  INV_X1    g050(.A(new_n236), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n237), .A2(new_n228), .ZN(new_n238));
  AOI21_X1  g052(.A(new_n235), .B1(new_n238), .B2(new_n232), .ZN(new_n239));
  AOI21_X1  g053(.A(KEYINPUT25), .B1(new_n239), .B2(new_n188), .ZN(new_n240));
  INV_X1    g054(.A(new_n228), .ZN(new_n241));
  OAI21_X1  g055(.A(new_n232), .B1(new_n241), .B2(new_n236), .ZN(new_n242));
  AND4_X1   g056(.A1(KEYINPUT25), .A2(new_n242), .A3(new_n188), .A4(new_n234), .ZN(new_n243));
  OAI21_X1  g057(.A(new_n189), .B1(new_n240), .B2(new_n243), .ZN(new_n244));
  NOR2_X1   g058(.A1(new_n189), .A2(G902), .ZN(new_n245));
  INV_X1    g059(.A(new_n245), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n242), .A2(new_n234), .ZN(new_n247));
  XNOR2_X1  g061(.A(new_n247), .B(KEYINPUT81), .ZN(new_n248));
  OAI21_X1  g062(.A(new_n244), .B1(new_n246), .B2(new_n248), .ZN(new_n249));
  XOR2_X1   g063(.A(KEYINPUT66), .B(G137), .Z(new_n250));
  NAND3_X1  g064(.A1(new_n250), .A2(KEYINPUT11), .A3(G134), .ZN(new_n251));
  XNOR2_X1  g065(.A(KEYINPUT67), .B(G131), .ZN(new_n252));
  INV_X1    g066(.A(G137), .ZN(new_n253));
  OAI21_X1  g067(.A(KEYINPUT11), .B1(new_n253), .B2(G134), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n253), .A2(G134), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n254), .A2(new_n255), .ZN(new_n256));
  AND3_X1   g070(.A1(new_n251), .A2(new_n252), .A3(new_n256), .ZN(new_n257));
  INV_X1    g071(.A(G131), .ZN(new_n258));
  XNOR2_X1  g072(.A(KEYINPUT66), .B(G137), .ZN(new_n259));
  INV_X1    g073(.A(G134), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n259), .A2(new_n260), .ZN(new_n261));
  AOI21_X1  g075(.A(new_n258), .B1(new_n261), .B2(new_n255), .ZN(new_n262));
  OAI21_X1  g076(.A(KEYINPUT68), .B1(new_n257), .B2(new_n262), .ZN(new_n263));
  OAI21_X1  g077(.A(KEYINPUT65), .B1(new_n197), .B2(G143), .ZN(new_n264));
  INV_X1    g078(.A(KEYINPUT65), .ZN(new_n265));
  INV_X1    g079(.A(G143), .ZN(new_n266));
  NAND3_X1  g080(.A1(new_n265), .A2(new_n266), .A3(G146), .ZN(new_n267));
  AOI22_X1  g081(.A1(new_n264), .A2(new_n267), .B1(G143), .B2(new_n197), .ZN(new_n268));
  INV_X1    g082(.A(KEYINPUT1), .ZN(new_n269));
  NAND3_X1  g083(.A1(new_n268), .A2(new_n269), .A3(G128), .ZN(new_n270));
  XNOR2_X1  g084(.A(G143), .B(G146), .ZN(new_n271));
  OAI21_X1  g085(.A(KEYINPUT1), .B1(new_n266), .B2(G146), .ZN(new_n272));
  INV_X1    g086(.A(KEYINPUT69), .ZN(new_n273));
  AOI22_X1  g087(.A1(new_n272), .A2(new_n273), .B1(new_n204), .B2(new_n205), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n197), .A2(G143), .ZN(new_n275));
  NAND3_X1  g089(.A1(new_n275), .A2(KEYINPUT69), .A3(KEYINPUT1), .ZN(new_n276));
  AOI211_X1 g090(.A(KEYINPUT71), .B(new_n271), .C1(new_n274), .C2(new_n276), .ZN(new_n277));
  INV_X1    g091(.A(KEYINPUT71), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n272), .A2(new_n273), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n204), .A2(new_n205), .ZN(new_n280));
  NAND3_X1  g094(.A1(new_n279), .A2(new_n276), .A3(new_n280), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n266), .A2(G146), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n275), .A2(new_n282), .ZN(new_n283));
  AOI21_X1  g097(.A(new_n278), .B1(new_n281), .B2(new_n283), .ZN(new_n284));
  OAI21_X1  g098(.A(new_n270), .B1(new_n277), .B2(new_n284), .ZN(new_n285));
  NAND3_X1  g099(.A1(new_n251), .A2(new_n252), .A3(new_n256), .ZN(new_n286));
  INV_X1    g100(.A(KEYINPUT68), .ZN(new_n287));
  AND2_X1   g101(.A1(new_n261), .A2(new_n255), .ZN(new_n288));
  OAI211_X1 g102(.A(new_n286), .B(new_n287), .C1(new_n258), .C2(new_n288), .ZN(new_n289));
  NAND3_X1  g103(.A1(new_n263), .A2(new_n285), .A3(new_n289), .ZN(new_n290));
  AOI21_X1  g104(.A(new_n258), .B1(new_n251), .B2(new_n256), .ZN(new_n291));
  OR2_X1    g105(.A1(new_n257), .A2(new_n291), .ZN(new_n292));
  NAND2_X1  g106(.A1(KEYINPUT0), .A2(G128), .ZN(new_n293));
  INV_X1    g107(.A(new_n293), .ZN(new_n294));
  NOR2_X1   g108(.A1(KEYINPUT0), .A2(G128), .ZN(new_n295));
  NOR2_X1   g109(.A1(new_n294), .A2(new_n295), .ZN(new_n296));
  AOI22_X1  g110(.A1(new_n268), .A2(new_n294), .B1(new_n296), .B2(new_n283), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n292), .A2(new_n297), .ZN(new_n298));
  NAND2_X1  g112(.A1(new_n290), .A2(new_n298), .ZN(new_n299));
  XOR2_X1   g113(.A(KEYINPUT64), .B(KEYINPUT30), .Z(new_n300));
  NAND2_X1  g114(.A1(new_n299), .A2(new_n300), .ZN(new_n301));
  INV_X1    g115(.A(G119), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n302), .A2(G116), .ZN(new_n303));
  INV_X1    g117(.A(G116), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n304), .A2(G119), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n303), .A2(new_n305), .ZN(new_n306));
  XNOR2_X1  g120(.A(KEYINPUT2), .B(G113), .ZN(new_n307));
  NOR2_X1   g121(.A1(new_n306), .A2(new_n307), .ZN(new_n308));
  INV_X1    g122(.A(new_n308), .ZN(new_n309));
  INV_X1    g123(.A(KEYINPUT72), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n306), .A2(new_n307), .ZN(new_n311));
  NAND3_X1  g125(.A1(new_n309), .A2(new_n310), .A3(new_n311), .ZN(new_n312));
  NAND3_X1  g126(.A1(new_n306), .A2(new_n307), .A3(KEYINPUT72), .ZN(new_n313));
  NAND2_X1  g127(.A1(new_n312), .A2(new_n313), .ZN(new_n314));
  INV_X1    g128(.A(new_n314), .ZN(new_n315));
  INV_X1    g129(.A(KEYINPUT73), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n285), .A2(new_n316), .ZN(new_n317));
  NOR2_X1   g131(.A1(new_n257), .A2(new_n262), .ZN(new_n318));
  OAI211_X1 g132(.A(KEYINPUT73), .B(new_n270), .C1(new_n277), .C2(new_n284), .ZN(new_n319));
  NAND3_X1  g133(.A1(new_n317), .A2(new_n318), .A3(new_n319), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n320), .A2(new_n298), .ZN(new_n321));
  INV_X1    g135(.A(KEYINPUT30), .ZN(new_n322));
  OAI211_X1 g136(.A(new_n301), .B(new_n315), .C1(new_n321), .C2(new_n322), .ZN(new_n323));
  NAND3_X1  g137(.A1(new_n320), .A2(new_n314), .A3(new_n298), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n323), .A2(new_n324), .ZN(new_n325));
  NOR2_X1   g139(.A1(G237), .A2(G953), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n326), .A2(G210), .ZN(new_n327));
  XOR2_X1   g141(.A(new_n327), .B(KEYINPUT27), .Z(new_n328));
  XNOR2_X1  g142(.A(KEYINPUT26), .B(G101), .ZN(new_n329));
  XNOR2_X1  g143(.A(new_n328), .B(new_n329), .ZN(new_n330));
  AOI21_X1  g144(.A(KEYINPUT29), .B1(new_n325), .B2(new_n330), .ZN(new_n331));
  INV_X1    g145(.A(new_n324), .ZN(new_n332));
  AOI22_X1  g146(.A1(new_n332), .A2(KEYINPUT28), .B1(new_n315), .B2(new_n299), .ZN(new_n333));
  OAI21_X1  g147(.A(new_n333), .B1(KEYINPUT28), .B2(new_n332), .ZN(new_n334));
  XNOR2_X1  g148(.A(new_n330), .B(KEYINPUT74), .ZN(new_n335));
  OAI21_X1  g149(.A(new_n331), .B1(new_n334), .B2(new_n335), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n336), .A2(KEYINPUT75), .ZN(new_n337));
  INV_X1    g151(.A(KEYINPUT75), .ZN(new_n338));
  OAI211_X1 g152(.A(new_n331), .B(new_n338), .C1(new_n334), .C2(new_n335), .ZN(new_n339));
  INV_X1    g153(.A(new_n188), .ZN(new_n340));
  AOI21_X1  g154(.A(new_n314), .B1(new_n320), .B2(new_n298), .ZN(new_n341));
  OAI21_X1  g155(.A(KEYINPUT28), .B1(new_n332), .B2(new_n341), .ZN(new_n342));
  INV_X1    g156(.A(KEYINPUT76), .ZN(new_n343));
  INV_X1    g157(.A(KEYINPUT28), .ZN(new_n344));
  AOI21_X1  g158(.A(new_n343), .B1(new_n324), .B2(new_n344), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n342), .A2(new_n345), .ZN(new_n346));
  NAND3_X1  g160(.A1(new_n324), .A2(new_n343), .A3(new_n344), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n346), .A2(new_n347), .ZN(new_n348));
  INV_X1    g162(.A(new_n330), .ZN(new_n349));
  AND2_X1   g163(.A1(new_n349), .A2(KEYINPUT29), .ZN(new_n350));
  AOI21_X1  g164(.A(new_n340), .B1(new_n348), .B2(new_n350), .ZN(new_n351));
  NAND3_X1  g165(.A1(new_n337), .A2(new_n339), .A3(new_n351), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n352), .A2(G472), .ZN(new_n353));
  NAND3_X1  g167(.A1(new_n323), .A2(new_n324), .A3(new_n349), .ZN(new_n354));
  INV_X1    g168(.A(KEYINPUT31), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n354), .A2(new_n355), .ZN(new_n356));
  NAND4_X1  g170(.A1(new_n323), .A2(KEYINPUT31), .A3(new_n324), .A4(new_n349), .ZN(new_n357));
  AOI22_X1  g171(.A1(new_n356), .A2(new_n357), .B1(new_n334), .B2(new_n335), .ZN(new_n358));
  NOR2_X1   g172(.A1(G472), .A2(G902), .ZN(new_n359));
  INV_X1    g173(.A(new_n359), .ZN(new_n360));
  OAI21_X1  g174(.A(KEYINPUT32), .B1(new_n358), .B2(new_n360), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n356), .A2(new_n357), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n334), .A2(new_n335), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n362), .A2(new_n363), .ZN(new_n364));
  INV_X1    g178(.A(KEYINPUT32), .ZN(new_n365));
  NAND3_X1  g179(.A1(new_n364), .A2(new_n365), .A3(new_n359), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n361), .A2(new_n366), .ZN(new_n367));
  AOI21_X1  g181(.A(new_n249), .B1(new_n353), .B2(new_n367), .ZN(new_n368));
  INV_X1    g182(.A(KEYINPUT89), .ZN(new_n369));
  INV_X1    g183(.A(new_n190), .ZN(new_n370));
  OAI21_X1  g184(.A(new_n369), .B1(new_n297), .B2(new_n370), .ZN(new_n371));
  INV_X1    g185(.A(new_n371), .ZN(new_n372));
  NOR3_X1   g186(.A1(new_n297), .A2(new_n369), .A3(new_n370), .ZN(new_n373));
  OAI21_X1  g187(.A(KEYINPUT90), .B1(new_n372), .B2(new_n373), .ZN(new_n374));
  INV_X1    g188(.A(new_n373), .ZN(new_n375));
  INV_X1    g189(.A(KEYINPUT90), .ZN(new_n376));
  NAND3_X1  g190(.A1(new_n375), .A2(new_n376), .A3(new_n371), .ZN(new_n377));
  INV_X1    g191(.A(new_n270), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n281), .A2(new_n283), .ZN(new_n379));
  NAND2_X1  g193(.A1(new_n379), .A2(KEYINPUT71), .ZN(new_n380));
  NAND3_X1  g194(.A1(new_n281), .A2(new_n278), .A3(new_n283), .ZN(new_n381));
  AOI21_X1  g195(.A(new_n378), .B1(new_n380), .B2(new_n381), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n382), .A2(new_n370), .ZN(new_n383));
  NAND3_X1  g197(.A1(new_n374), .A2(new_n377), .A3(new_n383), .ZN(new_n384));
  INV_X1    g198(.A(G224), .ZN(new_n385));
  NOR2_X1   g199(.A1(new_n385), .A2(G953), .ZN(new_n386));
  NAND2_X1  g200(.A1(new_n384), .A2(new_n386), .ZN(new_n387));
  INV_X1    g201(.A(new_n386), .ZN(new_n388));
  NAND4_X1  g202(.A1(new_n374), .A2(new_n377), .A3(new_n388), .A4(new_n383), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n387), .A2(new_n389), .ZN(new_n390));
  INV_X1    g204(.A(G104), .ZN(new_n391));
  OAI21_X1  g205(.A(KEYINPUT3), .B1(new_n391), .B2(G107), .ZN(new_n392));
  INV_X1    g206(.A(KEYINPUT3), .ZN(new_n393));
  INV_X1    g207(.A(G107), .ZN(new_n394));
  NAND3_X1  g208(.A1(new_n393), .A2(new_n394), .A3(G104), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n391), .A2(G107), .ZN(new_n396));
  NAND3_X1  g210(.A1(new_n392), .A2(new_n395), .A3(new_n396), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n397), .A2(G101), .ZN(new_n398));
  INV_X1    g212(.A(G101), .ZN(new_n399));
  NAND4_X1  g213(.A1(new_n392), .A2(new_n395), .A3(new_n399), .A4(new_n396), .ZN(new_n400));
  NAND3_X1  g214(.A1(new_n398), .A2(KEYINPUT4), .A3(new_n400), .ZN(new_n401));
  INV_X1    g215(.A(KEYINPUT4), .ZN(new_n402));
  NAND3_X1  g216(.A1(new_n397), .A2(new_n402), .A3(G101), .ZN(new_n403));
  NAND4_X1  g217(.A1(new_n312), .A2(new_n401), .A3(new_n313), .A4(new_n403), .ZN(new_n404));
  NOR2_X1   g218(.A1(new_n303), .A2(KEYINPUT5), .ZN(new_n405));
  INV_X1    g219(.A(G113), .ZN(new_n406));
  NOR2_X1   g220(.A1(new_n405), .A2(new_n406), .ZN(new_n407));
  NAND3_X1  g221(.A1(new_n303), .A2(new_n305), .A3(KEYINPUT5), .ZN(new_n408));
  NAND2_X1  g222(.A1(new_n407), .A2(new_n408), .ZN(new_n409));
  INV_X1    g223(.A(KEYINPUT87), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n409), .A2(new_n410), .ZN(new_n411));
  INV_X1    g225(.A(new_n396), .ZN(new_n412));
  NOR2_X1   g226(.A1(new_n391), .A2(G107), .ZN(new_n413));
  OAI21_X1  g227(.A(G101), .B1(new_n412), .B2(new_n413), .ZN(new_n414));
  NAND2_X1  g228(.A1(new_n414), .A2(new_n400), .ZN(new_n415));
  INV_X1    g229(.A(new_n415), .ZN(new_n416));
  NAND3_X1  g230(.A1(new_n407), .A2(KEYINPUT87), .A3(new_n408), .ZN(new_n417));
  NAND4_X1  g231(.A1(new_n411), .A2(new_n309), .A3(new_n416), .A4(new_n417), .ZN(new_n418));
  XNOR2_X1  g232(.A(G110), .B(G122), .ZN(new_n419));
  XNOR2_X1  g233(.A(new_n419), .B(KEYINPUT88), .ZN(new_n420));
  NAND3_X1  g234(.A1(new_n404), .A2(new_n418), .A3(new_n420), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n421), .A2(KEYINPUT6), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n404), .A2(new_n418), .ZN(new_n423));
  INV_X1    g237(.A(new_n420), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n423), .A2(new_n424), .ZN(new_n425));
  XNOR2_X1  g239(.A(new_n422), .B(new_n425), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n390), .A2(new_n426), .ZN(new_n427));
  AND2_X1   g241(.A1(new_n388), .A2(KEYINPUT7), .ZN(new_n428));
  NOR2_X1   g242(.A1(new_n372), .A2(new_n373), .ZN(new_n429));
  AOI21_X1  g243(.A(new_n428), .B1(new_n429), .B2(new_n383), .ZN(new_n430));
  XNOR2_X1  g244(.A(new_n420), .B(KEYINPUT8), .ZN(new_n431));
  NAND4_X1  g245(.A1(new_n411), .A2(new_n309), .A3(new_n415), .A4(new_n417), .ZN(new_n432));
  AOI21_X1  g246(.A(new_n308), .B1(new_n407), .B2(new_n408), .ZN(new_n433));
  AND2_X1   g247(.A1(new_n433), .A2(KEYINPUT91), .ZN(new_n434));
  OAI21_X1  g248(.A(new_n416), .B1(new_n433), .B2(KEYINPUT91), .ZN(new_n435));
  OAI211_X1 g249(.A(new_n431), .B(new_n432), .C1(new_n434), .C2(new_n435), .ZN(new_n436));
  NAND2_X1  g250(.A1(new_n436), .A2(new_n421), .ZN(new_n437));
  NOR2_X1   g251(.A1(new_n430), .A2(new_n437), .ZN(new_n438));
  NAND4_X1  g252(.A1(new_n374), .A2(new_n377), .A3(new_n383), .A4(new_n428), .ZN(new_n439));
  AOI21_X1  g253(.A(G902), .B1(new_n438), .B2(new_n439), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n427), .A2(new_n440), .ZN(new_n441));
  OAI21_X1  g255(.A(G210), .B1(G237), .B2(G902), .ZN(new_n442));
  INV_X1    g256(.A(new_n442), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n441), .A2(new_n443), .ZN(new_n444));
  NAND3_X1  g258(.A1(new_n427), .A2(new_n440), .A3(new_n442), .ZN(new_n445));
  NAND3_X1  g259(.A1(new_n444), .A2(KEYINPUT92), .A3(new_n445), .ZN(new_n446));
  OR2_X1    g260(.A1(new_n445), .A2(KEYINPUT92), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n446), .A2(new_n447), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n206), .A2(G143), .ZN(new_n449));
  INV_X1    g263(.A(KEYINPUT97), .ZN(new_n450));
  NOR2_X1   g264(.A1(new_n201), .A2(G143), .ZN(new_n451));
  AOI21_X1  g265(.A(new_n450), .B1(new_n451), .B2(KEYINPUT13), .ZN(new_n452));
  OAI211_X1 g266(.A(new_n449), .B(new_n452), .C1(KEYINPUT13), .C2(new_n451), .ZN(new_n453));
  NOR2_X1   g267(.A1(new_n280), .A2(new_n266), .ZN(new_n454));
  NOR2_X1   g268(.A1(new_n451), .A2(KEYINPUT13), .ZN(new_n455));
  OAI21_X1  g269(.A(new_n450), .B1(new_n454), .B2(new_n455), .ZN(new_n456));
  AND3_X1   g270(.A1(new_n453), .A2(G134), .A3(new_n456), .ZN(new_n457));
  INV_X1    g271(.A(new_n451), .ZN(new_n458));
  NAND3_X1  g272(.A1(new_n449), .A2(new_n260), .A3(new_n458), .ZN(new_n459));
  INV_X1    g273(.A(KEYINPUT96), .ZN(new_n460));
  INV_X1    g274(.A(G122), .ZN(new_n461));
  OAI21_X1  g275(.A(new_n460), .B1(new_n461), .B2(G116), .ZN(new_n462));
  NAND3_X1  g276(.A1(new_n304), .A2(KEYINPUT96), .A3(G122), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n461), .A2(G116), .ZN(new_n465));
  NAND2_X1  g279(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  NOR2_X1   g280(.A1(new_n466), .A2(G107), .ZN(new_n467));
  AOI21_X1  g281(.A(new_n394), .B1(new_n464), .B2(new_n465), .ZN(new_n468));
  OAI21_X1  g282(.A(new_n459), .B1(new_n467), .B2(new_n468), .ZN(new_n469));
  AOI21_X1  g283(.A(new_n260), .B1(new_n449), .B2(new_n458), .ZN(new_n470));
  NOR3_X1   g284(.A1(new_n454), .A2(G134), .A3(new_n451), .ZN(new_n471));
  OAI22_X1  g285(.A1(new_n470), .A2(new_n471), .B1(G107), .B2(new_n466), .ZN(new_n472));
  OR2_X1    g286(.A1(new_n464), .A2(KEYINPUT14), .ZN(new_n473));
  AOI22_X1  g287(.A1(new_n464), .A2(KEYINPUT14), .B1(G116), .B2(new_n461), .ZN(new_n474));
  AOI21_X1  g288(.A(new_n394), .B1(new_n473), .B2(new_n474), .ZN(new_n475));
  OAI22_X1  g289(.A1(new_n457), .A2(new_n469), .B1(new_n472), .B2(new_n475), .ZN(new_n476));
  XNOR2_X1  g290(.A(KEYINPUT9), .B(G234), .ZN(new_n477));
  NOR3_X1   g291(.A1(new_n477), .A2(new_n187), .A3(G953), .ZN(new_n478));
  INV_X1    g292(.A(new_n478), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n476), .A2(new_n479), .ZN(new_n480));
  OAI221_X1 g294(.A(new_n478), .B1(new_n472), .B2(new_n475), .C1(new_n457), .C2(new_n469), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n480), .A2(new_n481), .ZN(new_n482));
  NAND2_X1  g296(.A1(new_n482), .A2(new_n188), .ZN(new_n483));
  INV_X1    g297(.A(G478), .ZN(new_n484));
  NOR2_X1   g298(.A1(new_n484), .A2(KEYINPUT15), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n483), .A2(new_n485), .ZN(new_n486));
  INV_X1    g300(.A(new_n485), .ZN(new_n487));
  NAND3_X1  g301(.A1(new_n482), .A2(new_n188), .A3(new_n487), .ZN(new_n488));
  NAND3_X1  g302(.A1(new_n486), .A2(KEYINPUT98), .A3(new_n488), .ZN(new_n489));
  INV_X1    g303(.A(KEYINPUT98), .ZN(new_n490));
  AOI21_X1  g304(.A(new_n487), .B1(new_n482), .B2(new_n188), .ZN(new_n491));
  AOI211_X1 g305(.A(new_n340), .B(new_n485), .C1(new_n480), .C2(new_n481), .ZN(new_n492));
  OAI21_X1  g306(.A(new_n490), .B1(new_n491), .B2(new_n492), .ZN(new_n493));
  AND2_X1   g307(.A1(new_n489), .A2(new_n493), .ZN(new_n494));
  INV_X1    g308(.A(G952), .ZN(new_n495));
  AOI211_X1 g309(.A(G953), .B(new_n495), .C1(G234), .C2(G237), .ZN(new_n496));
  AOI211_X1 g310(.A(new_n230), .B(new_n188), .C1(G234), .C2(G237), .ZN(new_n497));
  XNOR2_X1  g311(.A(KEYINPUT21), .B(G898), .ZN(new_n498));
  AOI21_X1  g312(.A(new_n496), .B1(new_n497), .B2(new_n498), .ZN(new_n499));
  INV_X1    g313(.A(new_n499), .ZN(new_n500));
  INV_X1    g314(.A(KEYINPUT20), .ZN(new_n501));
  NOR2_X1   g315(.A1(G475), .A2(G902), .ZN(new_n502));
  OR2_X1    g316(.A1(new_n266), .A2(KEYINPUT94), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n326), .A2(G214), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  XNOR2_X1  g319(.A(KEYINPUT94), .B(G143), .ZN(new_n506));
  OAI21_X1  g320(.A(new_n505), .B1(new_n504), .B2(new_n506), .ZN(new_n507));
  INV_X1    g321(.A(new_n252), .ZN(new_n508));
  OR2_X1    g322(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  INV_X1    g323(.A(KEYINPUT17), .ZN(new_n510));
  NAND2_X1  g324(.A1(new_n507), .A2(new_n508), .ZN(new_n511));
  NAND3_X1  g325(.A1(new_n509), .A2(new_n510), .A3(new_n511), .ZN(new_n512));
  NAND3_X1  g326(.A1(new_n507), .A2(KEYINPUT17), .A3(new_n508), .ZN(new_n513));
  NAND4_X1  g327(.A1(new_n512), .A2(new_n198), .A3(new_n221), .A4(new_n513), .ZN(new_n514));
  NAND2_X1  g328(.A1(KEYINPUT18), .A2(G131), .ZN(new_n515));
  XNOR2_X1  g329(.A(new_n507), .B(new_n515), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n195), .A2(G146), .ZN(new_n517));
  AOI21_X1  g331(.A(KEYINPUT95), .B1(new_n517), .B2(new_n200), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n517), .A2(new_n200), .ZN(new_n519));
  INV_X1    g333(.A(KEYINPUT95), .ZN(new_n520));
  NOR2_X1   g334(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  OAI21_X1  g335(.A(new_n516), .B1(new_n518), .B2(new_n521), .ZN(new_n522));
  XNOR2_X1  g336(.A(G113), .B(G122), .ZN(new_n523));
  XNOR2_X1  g337(.A(new_n523), .B(new_n391), .ZN(new_n524));
  AND3_X1   g338(.A1(new_n514), .A2(new_n522), .A3(new_n524), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n509), .A2(new_n511), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n195), .A2(KEYINPUT19), .ZN(new_n527));
  INV_X1    g341(.A(KEYINPUT19), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n199), .A2(new_n528), .ZN(new_n529));
  NAND3_X1  g343(.A1(new_n527), .A2(new_n197), .A3(new_n529), .ZN(new_n530));
  NAND3_X1  g344(.A1(new_n526), .A2(new_n198), .A3(new_n530), .ZN(new_n531));
  AOI21_X1  g345(.A(new_n524), .B1(new_n522), .B2(new_n531), .ZN(new_n532));
  OAI211_X1 g346(.A(new_n501), .B(new_n502), .C1(new_n525), .C2(new_n532), .ZN(new_n533));
  INV_X1    g347(.A(new_n502), .ZN(new_n534));
  INV_X1    g348(.A(new_n532), .ZN(new_n535));
  NAND3_X1  g349(.A1(new_n514), .A2(new_n522), .A3(new_n524), .ZN(new_n536));
  AOI21_X1  g350(.A(new_n534), .B1(new_n535), .B2(new_n536), .ZN(new_n537));
  XNOR2_X1  g351(.A(KEYINPUT93), .B(KEYINPUT20), .ZN(new_n538));
  OAI21_X1  g352(.A(new_n533), .B1(new_n537), .B2(new_n538), .ZN(new_n539));
  INV_X1    g353(.A(G902), .ZN(new_n540));
  AOI21_X1  g354(.A(new_n524), .B1(new_n514), .B2(new_n522), .ZN(new_n541));
  OAI21_X1  g355(.A(new_n540), .B1(new_n525), .B2(new_n541), .ZN(new_n542));
  NAND2_X1  g356(.A1(new_n542), .A2(G475), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n539), .A2(new_n543), .ZN(new_n544));
  INV_X1    g358(.A(new_n544), .ZN(new_n545));
  NAND3_X1  g359(.A1(new_n494), .A2(new_n500), .A3(new_n545), .ZN(new_n546));
  OAI21_X1  g360(.A(G214), .B1(G237), .B2(G902), .ZN(new_n547));
  INV_X1    g361(.A(new_n547), .ZN(new_n548));
  NOR3_X1   g362(.A1(new_n448), .A2(new_n546), .A3(new_n548), .ZN(new_n549));
  INV_X1    g363(.A(G221), .ZN(new_n550));
  INV_X1    g364(.A(new_n477), .ZN(new_n551));
  AOI21_X1  g365(.A(new_n550), .B1(new_n551), .B2(new_n540), .ZN(new_n552));
  INV_X1    g366(.A(KEYINPUT86), .ZN(new_n553));
  NOR2_X1   g367(.A1(new_n257), .A2(new_n291), .ZN(new_n554));
  AND2_X1   g368(.A1(new_n416), .A2(KEYINPUT10), .ZN(new_n555));
  NAND3_X1  g369(.A1(new_n317), .A2(new_n319), .A3(new_n555), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n556), .A2(KEYINPUT83), .ZN(new_n557));
  INV_X1    g371(.A(KEYINPUT83), .ZN(new_n558));
  NAND4_X1  g372(.A1(new_n317), .A2(new_n558), .A3(new_n319), .A4(new_n555), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n557), .A2(new_n559), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n401), .A2(new_n403), .ZN(new_n561));
  INV_X1    g375(.A(new_n561), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n562), .A2(new_n297), .ZN(new_n563));
  AOI21_X1  g377(.A(new_n201), .B1(new_n275), .B2(KEYINPUT1), .ZN(new_n564));
  OR2_X1    g378(.A1(new_n268), .A2(new_n564), .ZN(new_n565));
  AOI21_X1  g379(.A(new_n415), .B1(new_n565), .B2(new_n270), .ZN(new_n566));
  XNOR2_X1  g380(.A(KEYINPUT82), .B(KEYINPUT10), .ZN(new_n567));
  OAI21_X1  g381(.A(new_n563), .B1(new_n566), .B2(new_n567), .ZN(new_n568));
  INV_X1    g382(.A(new_n568), .ZN(new_n569));
  AOI21_X1  g383(.A(new_n554), .B1(new_n560), .B2(new_n569), .ZN(new_n570));
  AOI211_X1 g384(.A(new_n292), .B(new_n568), .C1(new_n557), .C2(new_n559), .ZN(new_n571));
  XNOR2_X1  g385(.A(G110), .B(G140), .ZN(new_n572));
  NAND2_X1  g386(.A1(new_n230), .A2(G227), .ZN(new_n573));
  XOR2_X1   g387(.A(new_n572), .B(new_n573), .Z(new_n574));
  NOR3_X1   g388(.A1(new_n570), .A2(new_n571), .A3(new_n574), .ZN(new_n575));
  INV_X1    g389(.A(new_n574), .ZN(new_n576));
  AOI21_X1  g390(.A(new_n568), .B1(new_n557), .B2(new_n559), .ZN(new_n577));
  NAND2_X1  g391(.A1(new_n577), .A2(new_n554), .ZN(new_n578));
  OAI211_X1 g392(.A(new_n270), .B(new_n415), .C1(new_n277), .C2(new_n284), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n565), .A2(new_n270), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n580), .A2(new_n416), .ZN(new_n581));
  AOI21_X1  g395(.A(new_n554), .B1(new_n579), .B2(new_n581), .ZN(new_n582));
  NAND2_X1  g396(.A1(new_n582), .A2(KEYINPUT12), .ZN(new_n583));
  INV_X1    g397(.A(KEYINPUT84), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  NAND3_X1  g399(.A1(new_n582), .A2(KEYINPUT84), .A3(KEYINPUT12), .ZN(new_n586));
  NAND2_X1  g400(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  INV_X1    g401(.A(KEYINPUT85), .ZN(new_n588));
  INV_X1    g402(.A(KEYINPUT12), .ZN(new_n589));
  AOI21_X1  g403(.A(new_n566), .B1(new_n382), .B2(new_n415), .ZN(new_n590));
  OAI211_X1 g404(.A(new_n588), .B(new_n589), .C1(new_n590), .C2(new_n554), .ZN(new_n591));
  OAI21_X1  g405(.A(KEYINPUT85), .B1(new_n582), .B2(KEYINPUT12), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  NAND2_X1  g407(.A1(new_n587), .A2(new_n593), .ZN(new_n594));
  AOI21_X1  g408(.A(new_n576), .B1(new_n578), .B2(new_n594), .ZN(new_n595));
  OAI21_X1  g409(.A(new_n553), .B1(new_n575), .B2(new_n595), .ZN(new_n596));
  NAND2_X1  g410(.A1(new_n560), .A2(new_n569), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n597), .A2(new_n292), .ZN(new_n598));
  AOI21_X1  g412(.A(new_n574), .B1(new_n577), .B2(new_n554), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  AOI22_X1  g414(.A1(new_n585), .A2(new_n586), .B1(new_n591), .B2(new_n592), .ZN(new_n601));
  OAI21_X1  g415(.A(new_n574), .B1(new_n571), .B2(new_n601), .ZN(new_n602));
  NAND3_X1  g416(.A1(new_n600), .A2(new_n602), .A3(KEYINPUT86), .ZN(new_n603));
  NAND3_X1  g417(.A1(new_n596), .A2(G469), .A3(new_n603), .ZN(new_n604));
  INV_X1    g418(.A(G469), .ZN(new_n605));
  NOR2_X1   g419(.A1(new_n605), .A2(new_n540), .ZN(new_n606));
  OAI21_X1  g420(.A(new_n574), .B1(new_n570), .B2(new_n571), .ZN(new_n607));
  NAND3_X1  g421(.A1(new_n578), .A2(new_n594), .A3(new_n576), .ZN(new_n608));
  AOI21_X1  g422(.A(new_n340), .B1(new_n607), .B2(new_n608), .ZN(new_n609));
  AOI21_X1  g423(.A(new_n606), .B1(new_n609), .B2(new_n605), .ZN(new_n610));
  AOI21_X1  g424(.A(new_n552), .B1(new_n604), .B2(new_n610), .ZN(new_n611));
  AND2_X1   g425(.A1(new_n549), .A2(new_n611), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n368), .A2(new_n612), .ZN(new_n613));
  XNOR2_X1  g427(.A(new_n613), .B(G101), .ZN(G3));
  INV_X1    g428(.A(new_n611), .ZN(new_n615));
  OAI21_X1  g429(.A(G472), .B1(new_n358), .B2(new_n340), .ZN(new_n616));
  NAND2_X1  g430(.A1(new_n364), .A2(new_n359), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  NOR3_X1   g432(.A1(new_n615), .A2(new_n249), .A3(new_n618), .ZN(new_n619));
  AOI21_X1  g433(.A(new_n548), .B1(new_n444), .B2(new_n445), .ZN(new_n620));
  INV_X1    g434(.A(new_n620), .ZN(new_n621));
  NOR2_X1   g435(.A1(new_n340), .A2(new_n484), .ZN(new_n622));
  NOR2_X1   g436(.A1(new_n482), .A2(KEYINPUT33), .ZN(new_n623));
  INV_X1    g437(.A(KEYINPUT33), .ZN(new_n624));
  AOI21_X1  g438(.A(new_n624), .B1(new_n480), .B2(new_n481), .ZN(new_n625));
  OAI21_X1  g439(.A(new_n622), .B1(new_n623), .B2(new_n625), .ZN(new_n626));
  NAND2_X1  g440(.A1(new_n483), .A2(new_n484), .ZN(new_n627));
  NAND2_X1  g441(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  NAND2_X1  g442(.A1(new_n544), .A2(new_n628), .ZN(new_n629));
  NOR3_X1   g443(.A1(new_n621), .A2(new_n499), .A3(new_n629), .ZN(new_n630));
  NAND2_X1  g444(.A1(new_n619), .A2(new_n630), .ZN(new_n631));
  XOR2_X1   g445(.A(KEYINPUT34), .B(G104), .Z(new_n632));
  XNOR2_X1  g446(.A(new_n631), .B(new_n632), .ZN(G6));
  XOR2_X1   g447(.A(new_n499), .B(KEYINPUT99), .Z(new_n634));
  INV_X1    g448(.A(new_n634), .ZN(new_n635));
  NOR2_X1   g449(.A1(new_n494), .A2(new_n635), .ZN(new_n636));
  XNOR2_X1  g450(.A(new_n537), .B(new_n538), .ZN(new_n637));
  AND2_X1   g451(.A1(new_n637), .A2(new_n543), .ZN(new_n638));
  AND3_X1   g452(.A1(new_n636), .A2(KEYINPUT100), .A3(new_n638), .ZN(new_n639));
  AOI21_X1  g453(.A(KEYINPUT100), .B1(new_n636), .B2(new_n638), .ZN(new_n640));
  NOR3_X1   g454(.A1(new_n639), .A2(new_n640), .A3(new_n621), .ZN(new_n641));
  NAND2_X1  g455(.A1(new_n619), .A2(new_n641), .ZN(new_n642));
  XOR2_X1   g456(.A(KEYINPUT35), .B(G107), .Z(new_n643));
  XNOR2_X1  g457(.A(new_n642), .B(new_n643), .ZN(G9));
  NAND3_X1  g458(.A1(new_n239), .A2(KEYINPUT25), .A3(new_n188), .ZN(new_n645));
  INV_X1    g459(.A(KEYINPUT25), .ZN(new_n646));
  OAI21_X1  g460(.A(new_n646), .B1(new_n247), .B2(new_n340), .ZN(new_n647));
  NAND2_X1  g461(.A1(new_n645), .A2(new_n647), .ZN(new_n648));
  NAND2_X1  g462(.A1(new_n220), .A2(new_n226), .ZN(new_n649));
  NOR2_X1   g463(.A1(new_n233), .A2(KEYINPUT36), .ZN(new_n650));
  XNOR2_X1  g464(.A(new_n649), .B(new_n650), .ZN(new_n651));
  AOI22_X1  g465(.A1(new_n648), .A2(new_n189), .B1(new_n245), .B2(new_n651), .ZN(new_n652));
  NOR2_X1   g466(.A1(new_n618), .A2(new_n652), .ZN(new_n653));
  NAND2_X1  g467(.A1(new_n612), .A2(new_n653), .ZN(new_n654));
  XNOR2_X1  g468(.A(new_n654), .B(KEYINPUT101), .ZN(new_n655));
  XNOR2_X1  g469(.A(KEYINPUT37), .B(G110), .ZN(new_n656));
  XNOR2_X1  g470(.A(new_n655), .B(new_n656), .ZN(G12));
  NAND2_X1  g471(.A1(new_n651), .A2(new_n245), .ZN(new_n658));
  NAND2_X1  g472(.A1(new_n244), .A2(new_n658), .ZN(new_n659));
  NAND2_X1  g473(.A1(new_n659), .A2(new_n620), .ZN(new_n660));
  INV_X1    g474(.A(new_n496), .ZN(new_n661));
  INV_X1    g475(.A(new_n497), .ZN(new_n662));
  OAI21_X1  g476(.A(new_n661), .B1(new_n662), .B2(G900), .ZN(new_n663));
  NAND2_X1  g477(.A1(new_n638), .A2(new_n663), .ZN(new_n664));
  NOR3_X1   g478(.A1(new_n660), .A2(new_n494), .A3(new_n664), .ZN(new_n665));
  NAND2_X1  g479(.A1(new_n353), .A2(new_n367), .ZN(new_n666));
  AND3_X1   g480(.A1(new_n665), .A2(new_n666), .A3(new_n611), .ZN(new_n667));
  XNOR2_X1  g481(.A(new_n667), .B(new_n201), .ZN(G30));
  INV_X1    g482(.A(G472), .ZN(new_n669));
  OAI21_X1  g483(.A(new_n335), .B1(new_n332), .B2(new_n341), .ZN(new_n670));
  NAND2_X1  g484(.A1(new_n354), .A2(new_n670), .ZN(new_n671));
  AOI21_X1  g485(.A(new_n669), .B1(new_n671), .B2(new_n540), .ZN(new_n672));
  AOI21_X1  g486(.A(new_n672), .B1(new_n361), .B2(new_n366), .ZN(new_n673));
  INV_X1    g487(.A(new_n673), .ZN(new_n674));
  XOR2_X1   g488(.A(KEYINPUT102), .B(KEYINPUT38), .Z(new_n675));
  XNOR2_X1  g489(.A(new_n675), .B(KEYINPUT103), .ZN(new_n676));
  XNOR2_X1  g490(.A(new_n448), .B(new_n676), .ZN(new_n677));
  AOI22_X1  g491(.A1(new_n489), .A2(new_n493), .B1(new_n539), .B2(new_n543), .ZN(new_n678));
  AND3_X1   g492(.A1(new_n652), .A2(new_n547), .A3(new_n678), .ZN(new_n679));
  AND3_X1   g493(.A1(new_n674), .A2(new_n677), .A3(new_n679), .ZN(new_n680));
  XNOR2_X1  g494(.A(new_n663), .B(KEYINPUT39), .ZN(new_n681));
  NAND2_X1  g495(.A1(new_n611), .A2(new_n681), .ZN(new_n682));
  OR2_X1    g496(.A1(new_n682), .A2(KEYINPUT40), .ZN(new_n683));
  NAND2_X1  g497(.A1(new_n682), .A2(KEYINPUT40), .ZN(new_n684));
  NAND3_X1  g498(.A1(new_n680), .A2(new_n683), .A3(new_n684), .ZN(new_n685));
  XNOR2_X1  g499(.A(new_n685), .B(G143), .ZN(G45));
  NAND3_X1  g500(.A1(new_n544), .A2(new_n628), .A3(new_n663), .ZN(new_n687));
  INV_X1    g501(.A(KEYINPUT104), .ZN(new_n688));
  XNOR2_X1  g502(.A(new_n687), .B(new_n688), .ZN(new_n689));
  NOR2_X1   g503(.A1(new_n660), .A2(new_n689), .ZN(new_n690));
  NAND3_X1  g504(.A1(new_n666), .A2(new_n611), .A3(new_n690), .ZN(new_n691));
  XNOR2_X1  g505(.A(new_n691), .B(G146), .ZN(G48));
  NAND2_X1  g506(.A1(new_n609), .A2(new_n605), .ZN(new_n693));
  INV_X1    g507(.A(new_n552), .ZN(new_n694));
  NAND2_X1  g508(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  INV_X1    g509(.A(KEYINPUT105), .ZN(new_n696));
  OR3_X1    g510(.A1(new_n609), .A2(new_n696), .A3(new_n605), .ZN(new_n697));
  OAI21_X1  g511(.A(new_n696), .B1(new_n609), .B2(new_n605), .ZN(new_n698));
  AOI21_X1  g512(.A(new_n695), .B1(new_n697), .B2(new_n698), .ZN(new_n699));
  NAND3_X1  g513(.A1(new_n368), .A2(new_n630), .A3(new_n699), .ZN(new_n700));
  XNOR2_X1  g514(.A(KEYINPUT41), .B(G113), .ZN(new_n701));
  XNOR2_X1  g515(.A(new_n700), .B(new_n701), .ZN(G15));
  NAND3_X1  g516(.A1(new_n368), .A2(new_n641), .A3(new_n699), .ZN(new_n703));
  XNOR2_X1  g517(.A(new_n703), .B(G116), .ZN(G18));
  NAND2_X1  g518(.A1(new_n697), .A2(new_n698), .ZN(new_n705));
  INV_X1    g519(.A(new_n695), .ZN(new_n706));
  NAND3_X1  g520(.A1(new_n705), .A2(new_n706), .A3(new_n620), .ZN(new_n707));
  INV_X1    g521(.A(new_n707), .ZN(new_n708));
  AOI21_X1  g522(.A(new_n546), .B1(new_n353), .B2(new_n367), .ZN(new_n709));
  NAND3_X1  g523(.A1(new_n708), .A2(new_n659), .A3(new_n709), .ZN(new_n710));
  XNOR2_X1  g524(.A(new_n710), .B(G119), .ZN(G21));
  INV_X1    g525(.A(KEYINPUT107), .ZN(new_n712));
  INV_X1    g526(.A(new_n678), .ZN(new_n713));
  OAI21_X1  g527(.A(new_n712), .B1(new_n621), .B2(new_n713), .ZN(new_n714));
  NAND3_X1  g528(.A1(new_n620), .A2(KEYINPUT107), .A3(new_n678), .ZN(new_n715));
  AOI21_X1  g529(.A(new_n635), .B1(new_n714), .B2(new_n715), .ZN(new_n716));
  INV_X1    g530(.A(new_n249), .ZN(new_n717));
  INV_X1    g531(.A(new_n335), .ZN(new_n718));
  INV_X1    g532(.A(KEYINPUT106), .ZN(new_n719));
  AOI21_X1  g533(.A(new_n718), .B1(new_n348), .B2(new_n719), .ZN(new_n720));
  NAND3_X1  g534(.A1(new_n346), .A2(KEYINPUT106), .A3(new_n347), .ZN(new_n721));
  NAND2_X1  g535(.A1(new_n720), .A2(new_n721), .ZN(new_n722));
  AOI21_X1  g536(.A(new_n360), .B1(new_n722), .B2(new_n362), .ZN(new_n723));
  AOI21_X1  g537(.A(new_n669), .B1(new_n364), .B2(new_n188), .ZN(new_n724));
  NOR2_X1   g538(.A1(new_n723), .A2(new_n724), .ZN(new_n725));
  NAND4_X1  g539(.A1(new_n716), .A2(new_n717), .A3(new_n725), .A4(new_n699), .ZN(new_n726));
  XNOR2_X1  g540(.A(KEYINPUT108), .B(G122), .ZN(new_n727));
  XNOR2_X1  g541(.A(new_n726), .B(new_n727), .ZN(G24));
  INV_X1    g542(.A(KEYINPUT109), .ZN(new_n729));
  NOR3_X1   g543(.A1(new_n723), .A2(new_n689), .A3(new_n724), .ZN(new_n730));
  NAND4_X1  g544(.A1(new_n708), .A2(new_n729), .A3(new_n659), .A4(new_n730), .ZN(new_n731));
  NAND3_X1  g545(.A1(new_n699), .A2(new_n620), .A3(new_n659), .ZN(new_n732));
  AOI22_X1  g546(.A1(new_n539), .A2(new_n543), .B1(new_n626), .B2(new_n627), .ZN(new_n733));
  AOI21_X1  g547(.A(KEYINPUT104), .B1(new_n733), .B2(new_n663), .ZN(new_n734));
  AND4_X1   g548(.A1(KEYINPUT104), .A2(new_n544), .A3(new_n628), .A4(new_n663), .ZN(new_n735));
  NOR2_X1   g549(.A1(new_n734), .A2(new_n735), .ZN(new_n736));
  AOI22_X1  g550(.A1(new_n720), .A2(new_n721), .B1(new_n356), .B2(new_n357), .ZN(new_n737));
  OAI211_X1 g551(.A(new_n736), .B(new_n616), .C1(new_n737), .C2(new_n360), .ZN(new_n738));
  OAI21_X1  g552(.A(KEYINPUT109), .B1(new_n732), .B2(new_n738), .ZN(new_n739));
  NAND2_X1  g553(.A1(new_n731), .A2(new_n739), .ZN(new_n740));
  XNOR2_X1  g554(.A(new_n740), .B(G125), .ZN(G27));
  INV_X1    g555(.A(KEYINPUT42), .ZN(new_n742));
  NOR2_X1   g556(.A1(new_n575), .A2(new_n595), .ZN(new_n743));
  NAND2_X1  g557(.A1(new_n743), .A2(G469), .ZN(new_n744));
  INV_X1    g558(.A(new_n606), .ZN(new_n745));
  NAND3_X1  g559(.A1(new_n744), .A2(new_n693), .A3(new_n745), .ZN(new_n746));
  NOR2_X1   g560(.A1(new_n552), .A2(new_n548), .ZN(new_n747));
  AND3_X1   g561(.A1(new_n746), .A2(new_n448), .A3(new_n747), .ZN(new_n748));
  NAND3_X1  g562(.A1(new_n368), .A2(new_n736), .A3(new_n748), .ZN(new_n749));
  AOI22_X1  g563(.A1(new_n367), .A2(KEYINPUT110), .B1(new_n352), .B2(G472), .ZN(new_n750));
  INV_X1    g564(.A(KEYINPUT110), .ZN(new_n751));
  NAND3_X1  g565(.A1(new_n361), .A2(new_n366), .A3(new_n751), .ZN(new_n752));
  AOI21_X1  g566(.A(new_n249), .B1(new_n750), .B2(new_n752), .ZN(new_n753));
  NAND4_X1  g567(.A1(new_n736), .A2(new_n746), .A3(new_n448), .A4(new_n747), .ZN(new_n754));
  NOR2_X1   g568(.A1(new_n754), .A2(new_n742), .ZN(new_n755));
  AOI22_X1  g569(.A1(new_n742), .A2(new_n749), .B1(new_n753), .B2(new_n755), .ZN(new_n756));
  XNOR2_X1  g570(.A(new_n756), .B(new_n258), .ZN(G33));
  NOR2_X1   g571(.A1(new_n664), .A2(new_n494), .ZN(new_n758));
  NAND4_X1  g572(.A1(new_n666), .A2(new_n748), .A3(new_n717), .A4(new_n758), .ZN(new_n759));
  XNOR2_X1  g573(.A(new_n759), .B(G134), .ZN(G36));
  OAI211_X1 g574(.A(new_n545), .B(new_n628), .C1(KEYINPUT113), .C2(KEYINPUT43), .ZN(new_n761));
  INV_X1    g575(.A(KEYINPUT43), .ZN(new_n762));
  NAND3_X1  g576(.A1(new_n539), .A2(KEYINPUT113), .A3(new_n543), .ZN(new_n763));
  INV_X1    g577(.A(new_n628), .ZN(new_n764));
  OAI211_X1 g578(.A(new_n762), .B(new_n763), .C1(new_n764), .C2(new_n544), .ZN(new_n765));
  INV_X1    g579(.A(KEYINPUT114), .ZN(new_n766));
  AND3_X1   g580(.A1(new_n761), .A2(new_n765), .A3(new_n766), .ZN(new_n767));
  AOI21_X1  g581(.A(new_n766), .B1(new_n761), .B2(new_n765), .ZN(new_n768));
  OR2_X1    g582(.A1(new_n767), .A2(new_n768), .ZN(new_n769));
  NAND4_X1  g583(.A1(new_n769), .A2(KEYINPUT44), .A3(new_n618), .A4(new_n659), .ZN(new_n770));
  INV_X1    g584(.A(KEYINPUT44), .ZN(new_n771));
  OAI21_X1  g585(.A(new_n659), .B1(new_n767), .B2(new_n768), .ZN(new_n772));
  INV_X1    g586(.A(new_n618), .ZN(new_n773));
  OAI21_X1  g587(.A(new_n771), .B1(new_n772), .B2(new_n773), .ZN(new_n774));
  NAND2_X1  g588(.A1(new_n448), .A2(new_n547), .ZN(new_n775));
  INV_X1    g589(.A(new_n775), .ZN(new_n776));
  AND3_X1   g590(.A1(new_n770), .A2(new_n774), .A3(new_n776), .ZN(new_n777));
  AOI21_X1  g591(.A(KEYINPUT45), .B1(new_n596), .B2(new_n603), .ZN(new_n778));
  OAI21_X1  g592(.A(KEYINPUT111), .B1(new_n778), .B2(new_n605), .ZN(new_n779));
  INV_X1    g593(.A(KEYINPUT45), .ZN(new_n780));
  AND3_X1   g594(.A1(new_n600), .A2(new_n602), .A3(KEYINPUT86), .ZN(new_n781));
  AOI21_X1  g595(.A(KEYINPUT86), .B1(new_n600), .B2(new_n602), .ZN(new_n782));
  OAI21_X1  g596(.A(new_n780), .B1(new_n781), .B2(new_n782), .ZN(new_n783));
  INV_X1    g597(.A(KEYINPUT111), .ZN(new_n784));
  NAND3_X1  g598(.A1(new_n783), .A2(new_n784), .A3(G469), .ZN(new_n785));
  NAND2_X1  g599(.A1(new_n743), .A2(KEYINPUT45), .ZN(new_n786));
  NAND3_X1  g600(.A1(new_n779), .A2(new_n785), .A3(new_n786), .ZN(new_n787));
  NAND2_X1  g601(.A1(new_n787), .A2(new_n745), .ZN(new_n788));
  INV_X1    g602(.A(KEYINPUT46), .ZN(new_n789));
  NAND2_X1  g603(.A1(new_n788), .A2(new_n789), .ZN(new_n790));
  INV_X1    g604(.A(KEYINPUT112), .ZN(new_n791));
  NOR2_X1   g605(.A1(new_n606), .A2(new_n789), .ZN(new_n792));
  AND3_X1   g606(.A1(new_n787), .A2(new_n791), .A3(new_n792), .ZN(new_n793));
  AOI21_X1  g607(.A(new_n791), .B1(new_n787), .B2(new_n792), .ZN(new_n794));
  OAI211_X1 g608(.A(new_n790), .B(new_n693), .C1(new_n793), .C2(new_n794), .ZN(new_n795));
  AND2_X1   g609(.A1(new_n681), .A2(new_n694), .ZN(new_n796));
  NAND3_X1  g610(.A1(new_n777), .A2(new_n795), .A3(new_n796), .ZN(new_n797));
  XNOR2_X1  g611(.A(new_n797), .B(G137), .ZN(G39));
  NOR2_X1   g612(.A1(new_n793), .A2(new_n794), .ZN(new_n799));
  NAND2_X1  g613(.A1(new_n596), .A2(new_n603), .ZN(new_n800));
  AOI21_X1  g614(.A(new_n605), .B1(new_n800), .B2(new_n780), .ZN(new_n801));
  AOI22_X1  g615(.A1(new_n801), .A2(new_n784), .B1(KEYINPUT45), .B2(new_n743), .ZN(new_n802));
  AOI21_X1  g616(.A(new_n606), .B1(new_n802), .B2(new_n779), .ZN(new_n803));
  OAI21_X1  g617(.A(new_n693), .B1(new_n803), .B2(KEYINPUT46), .ZN(new_n804));
  OAI21_X1  g618(.A(new_n694), .B1(new_n799), .B2(new_n804), .ZN(new_n805));
  NAND2_X1  g619(.A1(new_n805), .A2(KEYINPUT47), .ZN(new_n806));
  INV_X1    g620(.A(KEYINPUT47), .ZN(new_n807));
  NAND3_X1  g621(.A1(new_n795), .A2(new_n807), .A3(new_n694), .ZN(new_n808));
  NOR4_X1   g622(.A1(new_n666), .A2(new_n717), .A3(new_n689), .A4(new_n775), .ZN(new_n809));
  NAND3_X1  g623(.A1(new_n806), .A2(new_n808), .A3(new_n809), .ZN(new_n810));
  XNOR2_X1  g624(.A(new_n810), .B(G140), .ZN(G42));
  INV_X1    g625(.A(KEYINPUT119), .ZN(new_n812));
  INV_X1    g626(.A(KEYINPUT48), .ZN(new_n813));
  AOI21_X1  g627(.A(new_n661), .B1(new_n761), .B2(new_n765), .ZN(new_n814));
  NAND3_X1  g628(.A1(new_n699), .A2(new_n776), .A3(new_n814), .ZN(new_n815));
  INV_X1    g629(.A(new_n815), .ZN(new_n816));
  AOI21_X1  g630(.A(new_n813), .B1(new_n753), .B2(new_n816), .ZN(new_n817));
  INV_X1    g631(.A(new_n817), .ZN(new_n818));
  NAND3_X1  g632(.A1(new_n753), .A2(new_n813), .A3(new_n816), .ZN(new_n819));
  NAND2_X1  g633(.A1(new_n818), .A2(new_n819), .ZN(new_n820));
  NAND3_X1  g634(.A1(new_n725), .A2(new_n717), .A3(new_n814), .ZN(new_n821));
  OAI211_X1 g635(.A(G952), .B(new_n230), .C1(new_n821), .C2(new_n707), .ZN(new_n822));
  NAND3_X1  g636(.A1(new_n699), .A2(new_n496), .A3(new_n776), .ZN(new_n823));
  NAND2_X1  g637(.A1(new_n673), .A2(new_n717), .ZN(new_n824));
  NOR3_X1   g638(.A1(new_n823), .A2(new_n824), .A3(new_n629), .ZN(new_n825));
  NOR2_X1   g639(.A1(new_n822), .A2(new_n825), .ZN(new_n826));
  AOI21_X1  g640(.A(KEYINPUT118), .B1(new_n820), .B2(new_n826), .ZN(new_n827));
  INV_X1    g641(.A(new_n819), .ZN(new_n828));
  OAI211_X1 g642(.A(new_n826), .B(KEYINPUT118), .C1(new_n828), .C2(new_n817), .ZN(new_n829));
  INV_X1    g643(.A(new_n829), .ZN(new_n830));
  OR2_X1    g644(.A1(new_n827), .A2(new_n830), .ZN(new_n831));
  NOR2_X1   g645(.A1(new_n821), .A2(new_n775), .ZN(new_n832));
  INV_X1    g646(.A(new_n832), .ZN(new_n833));
  NAND2_X1  g647(.A1(new_n806), .A2(new_n808), .ZN(new_n834));
  NAND3_X1  g648(.A1(new_n705), .A2(new_n552), .A3(new_n693), .ZN(new_n835));
  AOI21_X1  g649(.A(new_n833), .B1(new_n834), .B2(new_n835), .ZN(new_n836));
  OR2_X1    g650(.A1(new_n823), .A2(new_n824), .ZN(new_n837));
  NAND2_X1  g651(.A1(new_n545), .A2(new_n764), .ZN(new_n838));
  OAI211_X1 g652(.A(new_n616), .B(new_n659), .C1(new_n737), .C2(new_n360), .ZN(new_n839));
  OAI22_X1  g653(.A1(new_n837), .A2(new_n838), .B1(new_n815), .B2(new_n839), .ZN(new_n840));
  INV_X1    g654(.A(KEYINPUT117), .ZN(new_n841));
  OR2_X1    g655(.A1(new_n840), .A2(new_n841), .ZN(new_n842));
  INV_X1    g656(.A(KEYINPUT51), .ZN(new_n843));
  NOR2_X1   g657(.A1(new_n677), .A2(new_n547), .ZN(new_n844));
  NAND2_X1  g658(.A1(new_n844), .A2(new_n699), .ZN(new_n845));
  INV_X1    g659(.A(KEYINPUT50), .ZN(new_n846));
  OR3_X1    g660(.A1(new_n845), .A2(new_n846), .A3(new_n821), .ZN(new_n847));
  OAI21_X1  g661(.A(new_n846), .B1(new_n845), .B2(new_n821), .ZN(new_n848));
  AOI21_X1  g662(.A(new_n843), .B1(new_n847), .B2(new_n848), .ZN(new_n849));
  NAND2_X1  g663(.A1(new_n840), .A2(new_n841), .ZN(new_n850));
  NAND3_X1  g664(.A1(new_n842), .A2(new_n849), .A3(new_n850), .ZN(new_n851));
  OAI21_X1  g665(.A(new_n831), .B1(new_n836), .B2(new_n851), .ZN(new_n852));
  NAND2_X1  g666(.A1(new_n787), .A2(new_n792), .ZN(new_n853));
  NAND2_X1  g667(.A1(new_n853), .A2(KEYINPUT112), .ZN(new_n854));
  NAND3_X1  g668(.A1(new_n787), .A2(new_n791), .A3(new_n792), .ZN(new_n855));
  NAND2_X1  g669(.A1(new_n854), .A2(new_n855), .ZN(new_n856));
  AOI22_X1  g670(.A1(new_n788), .A2(new_n789), .B1(new_n605), .B2(new_n609), .ZN(new_n857));
  AOI211_X1 g671(.A(KEYINPUT47), .B(new_n552), .C1(new_n856), .C2(new_n857), .ZN(new_n858));
  AOI21_X1  g672(.A(new_n807), .B1(new_n795), .B2(new_n694), .ZN(new_n859));
  OAI21_X1  g673(.A(new_n835), .B1(new_n858), .B2(new_n859), .ZN(new_n860));
  NAND2_X1  g674(.A1(new_n860), .A2(new_n832), .ZN(new_n861));
  AND2_X1   g675(.A1(new_n847), .A2(new_n848), .ZN(new_n862));
  NOR2_X1   g676(.A1(new_n862), .A2(new_n840), .ZN(new_n863));
  AOI21_X1  g677(.A(KEYINPUT51), .B1(new_n861), .B2(new_n863), .ZN(new_n864));
  OAI21_X1  g678(.A(new_n812), .B1(new_n852), .B2(new_n864), .ZN(new_n865));
  INV_X1    g679(.A(new_n863), .ZN(new_n866));
  OAI21_X1  g680(.A(new_n843), .B1(new_n836), .B2(new_n866), .ZN(new_n867));
  NOR2_X1   g681(.A1(new_n827), .A2(new_n830), .ZN(new_n868));
  INV_X1    g682(.A(new_n851), .ZN(new_n869));
  AOI21_X1  g683(.A(new_n868), .B1(new_n861), .B2(new_n869), .ZN(new_n870));
  NAND3_X1  g684(.A1(new_n867), .A2(new_n870), .A3(KEYINPUT119), .ZN(new_n871));
  INV_X1    g685(.A(new_n667), .ZN(new_n872));
  NAND4_X1  g686(.A1(new_n244), .A2(new_n694), .A3(new_n658), .A4(new_n663), .ZN(new_n873));
  AOI21_X1  g687(.A(new_n873), .B1(new_n714), .B2(new_n715), .ZN(new_n874));
  NAND3_X1  g688(.A1(new_n874), .A2(new_n674), .A3(new_n746), .ZN(new_n875));
  AND2_X1   g689(.A1(new_n875), .A2(new_n691), .ZN(new_n876));
  NAND3_X1  g690(.A1(new_n740), .A2(new_n872), .A3(new_n876), .ZN(new_n877));
  INV_X1    g691(.A(KEYINPUT52), .ZN(new_n878));
  NAND2_X1  g692(.A1(new_n877), .A2(new_n878), .ZN(new_n879));
  AOI21_X1  g693(.A(new_n667), .B1(new_n731), .B2(new_n739), .ZN(new_n880));
  NAND3_X1  g694(.A1(new_n880), .A2(KEYINPUT52), .A3(new_n876), .ZN(new_n881));
  NAND2_X1  g695(.A1(new_n879), .A2(new_n881), .ZN(new_n882));
  NAND4_X1  g696(.A1(new_n710), .A2(new_n700), .A3(new_n703), .A4(new_n726), .ZN(new_n883));
  INV_X1    g697(.A(KEYINPUT53), .ZN(new_n884));
  NOR3_X1   g698(.A1(new_n756), .A2(new_n883), .A3(new_n884), .ZN(new_n885));
  NOR2_X1   g699(.A1(new_n491), .A2(new_n492), .ZN(new_n886));
  OAI21_X1  g700(.A(new_n629), .B1(new_n886), .B2(new_n544), .ZN(new_n887));
  NAND2_X1  g701(.A1(new_n887), .A2(new_n634), .ZN(new_n888));
  NOR3_X1   g702(.A1(new_n888), .A2(new_n548), .A3(new_n448), .ZN(new_n889));
  NAND4_X1  g703(.A1(new_n889), .A2(new_n773), .A3(new_n717), .A4(new_n611), .ZN(new_n890));
  NAND3_X1  g704(.A1(new_n613), .A2(new_n654), .A3(new_n890), .ZN(new_n891));
  INV_X1    g705(.A(new_n891), .ZN(new_n892));
  OR2_X1    g706(.A1(new_n754), .A2(new_n839), .ZN(new_n893));
  NAND3_X1  g707(.A1(new_n638), .A2(new_n886), .A3(new_n663), .ZN(new_n894));
  NOR3_X1   g708(.A1(new_n775), .A2(new_n652), .A3(new_n894), .ZN(new_n895));
  NAND3_X1  g709(.A1(new_n666), .A2(new_n895), .A3(new_n611), .ZN(new_n896));
  AND3_X1   g710(.A1(new_n759), .A2(new_n893), .A3(new_n896), .ZN(new_n897));
  AOI21_X1  g711(.A(KEYINPUT116), .B1(new_n892), .B2(new_n897), .ZN(new_n898));
  NAND3_X1  g712(.A1(new_n759), .A2(new_n893), .A3(new_n896), .ZN(new_n899));
  INV_X1    g713(.A(KEYINPUT116), .ZN(new_n900));
  NOR3_X1   g714(.A1(new_n899), .A2(new_n891), .A3(new_n900), .ZN(new_n901));
  NOR2_X1   g715(.A1(new_n898), .A2(new_n901), .ZN(new_n902));
  NAND3_X1  g716(.A1(new_n882), .A2(new_n885), .A3(new_n902), .ZN(new_n903));
  INV_X1    g717(.A(KEYINPUT54), .ZN(new_n904));
  INV_X1    g718(.A(new_n883), .ZN(new_n905));
  NAND2_X1  g719(.A1(new_n749), .A2(new_n742), .ZN(new_n906));
  NAND2_X1  g720(.A1(new_n753), .A2(new_n755), .ZN(new_n907));
  NAND2_X1  g721(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  NAND4_X1  g722(.A1(new_n905), .A2(new_n908), .A3(new_n892), .A4(new_n897), .ZN(new_n909));
  AOI21_X1  g723(.A(new_n909), .B1(new_n879), .B2(new_n881), .ZN(new_n910));
  XOR2_X1   g724(.A(KEYINPUT115), .B(KEYINPUT53), .Z(new_n911));
  INV_X1    g725(.A(new_n911), .ZN(new_n912));
  OAI211_X1 g726(.A(new_n903), .B(new_n904), .C1(new_n910), .C2(new_n912), .ZN(new_n913));
  NOR2_X1   g727(.A1(new_n754), .A2(new_n839), .ZN(new_n914));
  AOI21_X1  g728(.A(new_n615), .B1(new_n367), .B2(new_n353), .ZN(new_n915));
  AOI21_X1  g729(.A(new_n914), .B1(new_n915), .B2(new_n895), .ZN(new_n916));
  OAI21_X1  g730(.A(new_n612), .B1(new_n368), .B2(new_n653), .ZN(new_n917));
  NAND4_X1  g731(.A1(new_n916), .A2(new_n759), .A3(new_n890), .A4(new_n917), .ZN(new_n918));
  NOR3_X1   g732(.A1(new_n918), .A2(new_n756), .A3(new_n883), .ZN(new_n919));
  AOI21_X1  g733(.A(KEYINPUT52), .B1(new_n880), .B2(new_n876), .ZN(new_n920));
  AND4_X1   g734(.A1(KEYINPUT52), .A2(new_n740), .A3(new_n872), .A4(new_n876), .ZN(new_n921));
  OAI211_X1 g735(.A(new_n919), .B(new_n911), .C1(new_n920), .C2(new_n921), .ZN(new_n922));
  OAI211_X1 g736(.A(new_n922), .B(KEYINPUT54), .C1(new_n910), .C2(new_n884), .ZN(new_n923));
  AND2_X1   g737(.A1(new_n913), .A2(new_n923), .ZN(new_n924));
  NAND3_X1  g738(.A1(new_n865), .A2(new_n871), .A3(new_n924), .ZN(new_n925));
  NAND2_X1  g739(.A1(new_n495), .A2(new_n230), .ZN(new_n926));
  NAND2_X1  g740(.A1(new_n925), .A2(new_n926), .ZN(new_n927));
  NAND2_X1  g741(.A1(new_n705), .A2(new_n693), .ZN(new_n928));
  AND2_X1   g742(.A1(new_n928), .A2(KEYINPUT49), .ZN(new_n929));
  NAND3_X1  g743(.A1(new_n545), .A2(new_n628), .A3(new_n747), .ZN(new_n930));
  NOR3_X1   g744(.A1(new_n929), .A2(new_n677), .A3(new_n930), .ZN(new_n931));
  NOR2_X1   g745(.A1(new_n674), .A2(new_n249), .ZN(new_n932));
  OAI211_X1 g746(.A(new_n931), .B(new_n932), .C1(KEYINPUT49), .C2(new_n928), .ZN(new_n933));
  NAND2_X1  g747(.A1(new_n927), .A2(new_n933), .ZN(G75));
  NOR2_X1   g748(.A1(new_n921), .A2(new_n920), .ZN(new_n935));
  OAI21_X1  g749(.A(new_n911), .B1(new_n935), .B2(new_n909), .ZN(new_n936));
  AOI21_X1  g750(.A(new_n188), .B1(new_n936), .B2(new_n903), .ZN(new_n937));
  NAND2_X1  g751(.A1(new_n937), .A2(new_n443), .ZN(new_n938));
  INV_X1    g752(.A(KEYINPUT56), .ZN(new_n939));
  XOR2_X1   g753(.A(new_n390), .B(new_n426), .Z(new_n940));
  XNOR2_X1  g754(.A(new_n940), .B(KEYINPUT55), .ZN(new_n941));
  AND3_X1   g755(.A1(new_n938), .A2(new_n939), .A3(new_n941), .ZN(new_n942));
  AOI21_X1  g756(.A(new_n941), .B1(new_n938), .B2(new_n939), .ZN(new_n943));
  NOR2_X1   g757(.A1(new_n230), .A2(G952), .ZN(new_n944));
  NOR3_X1   g758(.A1(new_n942), .A2(new_n943), .A3(new_n944), .ZN(G51));
  INV_X1    g759(.A(KEYINPUT121), .ZN(new_n946));
  INV_X1    g760(.A(new_n787), .ZN(new_n947));
  AND3_X1   g761(.A1(new_n937), .A2(new_n946), .A3(new_n947), .ZN(new_n948));
  AOI21_X1  g762(.A(new_n946), .B1(new_n937), .B2(new_n947), .ZN(new_n949));
  NOR2_X1   g763(.A1(new_n948), .A2(new_n949), .ZN(new_n950));
  AOI21_X1  g764(.A(new_n912), .B1(new_n882), .B2(new_n919), .ZN(new_n951));
  NOR2_X1   g765(.A1(new_n756), .A2(new_n883), .ZN(new_n952));
  NAND3_X1  g766(.A1(new_n892), .A2(new_n897), .A3(KEYINPUT116), .ZN(new_n953));
  OAI21_X1  g767(.A(new_n900), .B1(new_n899), .B2(new_n891), .ZN(new_n954));
  NAND4_X1  g768(.A1(new_n952), .A2(new_n953), .A3(KEYINPUT53), .A4(new_n954), .ZN(new_n955));
  NOR2_X1   g769(.A1(new_n935), .A2(new_n955), .ZN(new_n956));
  OAI21_X1  g770(.A(KEYINPUT54), .B1(new_n951), .B2(new_n956), .ZN(new_n957));
  NAND2_X1  g771(.A1(new_n957), .A2(new_n913), .ZN(new_n958));
  XNOR2_X1  g772(.A(KEYINPUT120), .B(KEYINPUT57), .ZN(new_n959));
  XNOR2_X1  g773(.A(new_n959), .B(new_n606), .ZN(new_n960));
  NAND2_X1  g774(.A1(new_n958), .A2(new_n960), .ZN(new_n961));
  NAND2_X1  g775(.A1(new_n607), .A2(new_n608), .ZN(new_n962));
  NAND2_X1  g776(.A1(new_n961), .A2(new_n962), .ZN(new_n963));
  AOI21_X1  g777(.A(new_n944), .B1(new_n950), .B2(new_n963), .ZN(G54));
  AND2_X1   g778(.A1(KEYINPUT58), .A2(G475), .ZN(new_n965));
  OAI211_X1 g779(.A(new_n340), .B(new_n965), .C1(new_n951), .C2(new_n956), .ZN(new_n966));
  NAND3_X1  g780(.A1(new_n966), .A2(new_n535), .A3(new_n536), .ZN(new_n967));
  INV_X1    g781(.A(new_n944), .ZN(new_n968));
  NAND2_X1  g782(.A1(new_n535), .A2(new_n536), .ZN(new_n969));
  NAND3_X1  g783(.A1(new_n937), .A2(new_n969), .A3(new_n965), .ZN(new_n970));
  NAND3_X1  g784(.A1(new_n967), .A2(new_n968), .A3(new_n970), .ZN(new_n971));
  INV_X1    g785(.A(KEYINPUT122), .ZN(new_n972));
  NAND2_X1  g786(.A1(new_n971), .A2(new_n972), .ZN(new_n973));
  NAND4_X1  g787(.A1(new_n967), .A2(new_n970), .A3(KEYINPUT122), .A4(new_n968), .ZN(new_n974));
  NAND2_X1  g788(.A1(new_n973), .A2(new_n974), .ZN(G60));
  NAND2_X1  g789(.A1(G478), .A2(G902), .ZN(new_n976));
  XOR2_X1   g790(.A(new_n976), .B(KEYINPUT59), .Z(new_n977));
  AOI21_X1  g791(.A(new_n977), .B1(new_n913), .B2(new_n923), .ZN(new_n978));
  OR2_X1    g792(.A1(new_n623), .A2(new_n625), .ZN(new_n979));
  OAI21_X1  g793(.A(new_n968), .B1(new_n978), .B2(new_n979), .ZN(new_n980));
  INV_X1    g794(.A(KEYINPUT123), .ZN(new_n981));
  INV_X1    g795(.A(new_n979), .ZN(new_n982));
  NOR2_X1   g796(.A1(new_n982), .A2(new_n977), .ZN(new_n983));
  AOI21_X1  g797(.A(new_n981), .B1(new_n958), .B2(new_n983), .ZN(new_n984));
  INV_X1    g798(.A(new_n983), .ZN(new_n985));
  AOI211_X1 g799(.A(KEYINPUT123), .B(new_n985), .C1(new_n957), .C2(new_n913), .ZN(new_n986));
  NOR3_X1   g800(.A1(new_n980), .A2(new_n984), .A3(new_n986), .ZN(G63));
  NAND2_X1  g801(.A1(G217), .A2(G902), .ZN(new_n988));
  XNOR2_X1  g802(.A(new_n988), .B(KEYINPUT60), .ZN(new_n989));
  INV_X1    g803(.A(new_n989), .ZN(new_n990));
  OAI211_X1 g804(.A(new_n651), .B(new_n990), .C1(new_n951), .C2(new_n956), .ZN(new_n991));
  AOI21_X1  g805(.A(new_n989), .B1(new_n936), .B2(new_n903), .ZN(new_n992));
  INV_X1    g806(.A(new_n248), .ZN(new_n993));
  OAI211_X1 g807(.A(new_n991), .B(new_n968), .C1(new_n992), .C2(new_n993), .ZN(new_n994));
  NAND2_X1  g808(.A1(KEYINPUT124), .A2(KEYINPUT61), .ZN(new_n995));
  INV_X1    g809(.A(KEYINPUT124), .ZN(new_n996));
  INV_X1    g810(.A(KEYINPUT61), .ZN(new_n997));
  NAND2_X1  g811(.A1(new_n996), .A2(new_n997), .ZN(new_n998));
  NAND3_X1  g812(.A1(new_n994), .A2(new_n995), .A3(new_n998), .ZN(new_n999));
  OAI21_X1  g813(.A(new_n990), .B1(new_n951), .B2(new_n956), .ZN(new_n1000));
  AOI21_X1  g814(.A(new_n944), .B1(new_n1000), .B2(new_n248), .ZN(new_n1001));
  NAND4_X1  g815(.A1(new_n1001), .A2(new_n996), .A3(new_n997), .A4(new_n991), .ZN(new_n1002));
  AND2_X1   g816(.A1(new_n999), .A2(new_n1002), .ZN(G66));
  NAND2_X1  g817(.A1(new_n905), .A2(new_n892), .ZN(new_n1004));
  NAND2_X1  g818(.A1(new_n1004), .A2(new_n230), .ZN(new_n1005));
  OAI21_X1  g819(.A(G953), .B1(new_n498), .B2(new_n385), .ZN(new_n1006));
  NAND2_X1  g820(.A1(new_n1005), .A2(new_n1006), .ZN(new_n1007));
  INV_X1    g821(.A(G898), .ZN(new_n1008));
  AOI21_X1  g822(.A(new_n426), .B1(new_n1008), .B2(G953), .ZN(new_n1009));
  XOR2_X1   g823(.A(new_n1007), .B(new_n1009), .Z(G69));
  INV_X1    g824(.A(new_n691), .ZN(new_n1011));
  AOI211_X1 g825(.A(new_n667), .B(new_n1011), .C1(new_n739), .C2(new_n731), .ZN(new_n1012));
  NAND3_X1  g826(.A1(new_n1012), .A2(KEYINPUT62), .A3(new_n685), .ZN(new_n1013));
  NAND3_X1  g827(.A1(new_n880), .A2(new_n685), .A3(new_n691), .ZN(new_n1014));
  INV_X1    g828(.A(KEYINPUT62), .ZN(new_n1015));
  NAND2_X1  g829(.A1(new_n1014), .A2(new_n1015), .ZN(new_n1016));
  NAND2_X1  g830(.A1(new_n1013), .A2(new_n1016), .ZN(new_n1017));
  AND2_X1   g831(.A1(new_n795), .A2(new_n796), .ZN(new_n1018));
  XNOR2_X1  g832(.A(new_n887), .B(KEYINPUT125), .ZN(new_n1019));
  NOR3_X1   g833(.A1(new_n682), .A2(new_n1019), .A3(new_n775), .ZN(new_n1020));
  AOI22_X1  g834(.A1(new_n1018), .A2(new_n777), .B1(new_n368), .B2(new_n1020), .ZN(new_n1021));
  NAND3_X1  g835(.A1(new_n1017), .A2(new_n1021), .A3(new_n810), .ZN(new_n1022));
  NAND2_X1  g836(.A1(new_n1022), .A2(new_n230), .ZN(new_n1023));
  OAI21_X1  g837(.A(new_n301), .B1(new_n321), .B2(new_n322), .ZN(new_n1024));
  NAND2_X1  g838(.A1(new_n527), .A2(new_n529), .ZN(new_n1025));
  XOR2_X1   g839(.A(new_n1024), .B(new_n1025), .Z(new_n1026));
  NAND2_X1  g840(.A1(new_n1023), .A2(new_n1026), .ZN(new_n1027));
  AOI21_X1  g841(.A(new_n1026), .B1(G900), .B2(G953), .ZN(new_n1028));
  NAND2_X1  g842(.A1(new_n797), .A2(new_n1012), .ZN(new_n1029));
  INV_X1    g843(.A(KEYINPUT126), .ZN(new_n1030));
  NAND2_X1  g844(.A1(new_n1029), .A2(new_n1030), .ZN(new_n1031));
  NAND2_X1  g845(.A1(new_n908), .A2(new_n759), .ZN(new_n1032));
  INV_X1    g846(.A(new_n753), .ZN(new_n1033));
  AOI21_X1  g847(.A(new_n1033), .B1(new_n715), .B2(new_n714), .ZN(new_n1034));
  AOI21_X1  g848(.A(new_n1032), .B1(new_n1018), .B2(new_n1034), .ZN(new_n1035));
  NAND3_X1  g849(.A1(new_n797), .A2(new_n1012), .A3(KEYINPUT126), .ZN(new_n1036));
  NAND4_X1  g850(.A1(new_n1031), .A2(new_n810), .A3(new_n1035), .A4(new_n1036), .ZN(new_n1037));
  OAI21_X1  g851(.A(new_n1028), .B1(new_n1037), .B2(G953), .ZN(new_n1038));
  NAND2_X1  g852(.A1(new_n1027), .A2(new_n1038), .ZN(new_n1039));
  AOI21_X1  g853(.A(new_n230), .B1(G227), .B2(G900), .ZN(new_n1040));
  XNOR2_X1  g854(.A(new_n1039), .B(new_n1040), .ZN(G72));
  NAND2_X1  g855(.A1(G472), .A2(G902), .ZN(new_n1042));
  XOR2_X1   g856(.A(new_n1042), .B(KEYINPUT63), .Z(new_n1043));
  OAI21_X1  g857(.A(new_n1043), .B1(new_n1037), .B2(new_n1004), .ZN(new_n1044));
  NOR2_X1   g858(.A1(new_n325), .A2(new_n349), .ZN(new_n1045));
  NAND2_X1  g859(.A1(new_n1044), .A2(new_n1045), .ZN(new_n1046));
  OAI21_X1  g860(.A(new_n1043), .B1(new_n1022), .B2(new_n1004), .ZN(new_n1047));
  AOI21_X1  g861(.A(new_n330), .B1(new_n323), .B2(new_n324), .ZN(new_n1048));
  NAND2_X1  g862(.A1(new_n1047), .A2(new_n1048), .ZN(new_n1049));
  INV_X1    g863(.A(new_n1043), .ZN(new_n1050));
  NOR3_X1   g864(.A1(new_n1045), .A2(new_n1050), .A3(new_n1048), .ZN(new_n1051));
  OAI211_X1 g865(.A(new_n922), .B(new_n1051), .C1(new_n910), .C2(new_n884), .ZN(new_n1052));
  AND2_X1   g866(.A1(new_n1052), .A2(new_n968), .ZN(new_n1053));
  NAND3_X1  g867(.A1(new_n1046), .A2(new_n1049), .A3(new_n1053), .ZN(new_n1054));
  NAND2_X1  g868(.A1(new_n1054), .A2(KEYINPUT127), .ZN(new_n1055));
  INV_X1    g869(.A(KEYINPUT127), .ZN(new_n1056));
  NAND4_X1  g870(.A1(new_n1046), .A2(new_n1049), .A3(new_n1053), .A4(new_n1056), .ZN(new_n1057));
  NAND2_X1  g871(.A1(new_n1055), .A2(new_n1057), .ZN(G57));
endmodule


