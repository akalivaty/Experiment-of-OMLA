//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 1 0 0 1 1 0 0 1 0 0 0 1 1 0 1 1 1 0 0 1 1 1 1 1 0 1 1 1 1 1 1 1 1 0 1 1 1 1 0 1 1 0 1 1 1 1 1 1 1 1 1 0 1 1 0 0 0 0 1 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:35:25 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n228, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n237, new_n238, new_n239,
    new_n240, new_n241, new_n242, new_n244, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n595, new_n596, new_n597, new_n598,
    new_n599, new_n600, new_n601, new_n602, new_n603, new_n604, new_n605,
    new_n606, new_n607, new_n608, new_n609, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n687, new_n688, new_n689, new_n690, new_n691, new_n692,
    new_n693, new_n694, new_n695, new_n696, new_n697, new_n698, new_n699,
    new_n700, new_n701, new_n702, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n798, new_n799,
    new_n800, new_n801, new_n802, new_n803, new_n804, new_n805, new_n806,
    new_n807, new_n808, new_n809, new_n810, new_n811, new_n812, new_n813,
    new_n814, new_n815, new_n816, new_n817, new_n818, new_n819, new_n820,
    new_n821, new_n822, new_n823, new_n824, new_n825, new_n826, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n977, new_n978, new_n979, new_n980, new_n981, new_n982, new_n983,
    new_n984, new_n985, new_n986, new_n987, new_n988, new_n989, new_n990,
    new_n991, new_n992, new_n993, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1013, new_n1014, new_n1015, new_n1016,
    new_n1017, new_n1018, new_n1019, new_n1020, new_n1021, new_n1022,
    new_n1023, new_n1024, new_n1025, new_n1026, new_n1027, new_n1028,
    new_n1029, new_n1030, new_n1031, new_n1032, new_n1033, new_n1034,
    new_n1035, new_n1036, new_n1037, new_n1038, new_n1040, new_n1041,
    new_n1042, new_n1043, new_n1044, new_n1045, new_n1046, new_n1047,
    new_n1048, new_n1049, new_n1050, new_n1051, new_n1052, new_n1053,
    new_n1054, new_n1055, new_n1056, new_n1057, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1119, new_n1120,
    new_n1121, new_n1122, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1177, new_n1178, new_n1179, new_n1180, new_n1181,
    new_n1182, new_n1183, new_n1184, new_n1185, new_n1186, new_n1187,
    new_n1188, new_n1189, new_n1190, new_n1191, new_n1192, new_n1193,
    new_n1194, new_n1195, new_n1196, new_n1198, new_n1199, new_n1200,
    new_n1202, new_n1203, new_n1205, new_n1206, new_n1207, new_n1208,
    new_n1209, new_n1210, new_n1211, new_n1212, new_n1213, new_n1214,
    new_n1215, new_n1216, new_n1217, new_n1218, new_n1219, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1264, new_n1265, new_n1266, new_n1267, new_n1268, new_n1269,
    new_n1270, new_n1271, new_n1272;
  INV_X1    g0000(.A(G50), .ZN(new_n201));
  INV_X1    g0001(.A(G58), .ZN(new_n202));
  INV_X1    g0002(.A(G68), .ZN(new_n203));
  NAND3_X1  g0003(.A1(new_n201), .A2(new_n202), .A3(new_n203), .ZN(new_n204));
  NOR2_X1   g0004(.A1(new_n204), .A2(G77), .ZN(G353));
  OAI21_X1  g0005(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0006(.A1(G1), .A2(G20), .ZN(new_n207));
  NOR2_X1   g0007(.A1(new_n207), .A2(G13), .ZN(new_n208));
  OAI211_X1 g0008(.A(new_n208), .B(G250), .C1(G257), .C2(G264), .ZN(new_n209));
  XNOR2_X1  g0009(.A(new_n209), .B(KEYINPUT0), .ZN(new_n210));
  NAND2_X1  g0010(.A1(new_n202), .A2(new_n203), .ZN(new_n211));
  NAND2_X1  g0011(.A1(new_n211), .A2(G50), .ZN(new_n212));
  INV_X1    g0012(.A(new_n212), .ZN(new_n213));
  NAND2_X1  g0013(.A1(G1), .A2(G13), .ZN(new_n214));
  INV_X1    g0014(.A(G20), .ZN(new_n215));
  NOR2_X1   g0015(.A1(new_n214), .A2(new_n215), .ZN(new_n216));
  NAND2_X1  g0016(.A1(new_n213), .A2(new_n216), .ZN(new_n217));
  AOI22_X1  g0017(.A1(G50), .A2(G226), .B1(G97), .B2(G257), .ZN(new_n218));
  INV_X1    g0018(.A(G232), .ZN(new_n219));
  INV_X1    g0019(.A(G238), .ZN(new_n220));
  OAI221_X1 g0020(.A(new_n218), .B1(new_n202), .B2(new_n219), .C1(new_n203), .C2(new_n220), .ZN(new_n221));
  AOI22_X1  g0021(.A1(G107), .A2(G264), .B1(G116), .B2(G270), .ZN(new_n222));
  AOI22_X1  g0022(.A1(G77), .A2(G244), .B1(G87), .B2(G250), .ZN(new_n223));
  NAND2_X1  g0023(.A1(new_n222), .A2(new_n223), .ZN(new_n224));
  OAI21_X1  g0024(.A(new_n207), .B1(new_n221), .B2(new_n224), .ZN(new_n225));
  OAI211_X1 g0025(.A(new_n210), .B(new_n217), .C1(KEYINPUT1), .C2(new_n225), .ZN(new_n226));
  AOI21_X1  g0026(.A(new_n226), .B1(KEYINPUT1), .B2(new_n225), .ZN(G361));
  XNOR2_X1  g0027(.A(G226), .B(G232), .ZN(new_n228));
  XNOR2_X1  g0028(.A(G238), .B(G244), .ZN(new_n229));
  XNOR2_X1  g0029(.A(new_n228), .B(new_n229), .ZN(new_n230));
  XNOR2_X1  g0030(.A(KEYINPUT64), .B(KEYINPUT2), .ZN(new_n231));
  XNOR2_X1  g0031(.A(new_n230), .B(new_n231), .ZN(new_n232));
  XNOR2_X1  g0032(.A(G250), .B(G257), .ZN(new_n233));
  XNOR2_X1  g0033(.A(G264), .B(G270), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n233), .B(new_n234), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n232), .B(new_n235), .ZN(G358));
  XOR2_X1   g0036(.A(G68), .B(G77), .Z(new_n237));
  XOR2_X1   g0037(.A(G50), .B(G58), .Z(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XOR2_X1   g0039(.A(G87), .B(G97), .Z(new_n240));
  XNOR2_X1  g0040(.A(G107), .B(G116), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XOR2_X1   g0042(.A(new_n239), .B(new_n242), .Z(G351));
  INV_X1    g0043(.A(G33), .ZN(new_n244));
  NAND2_X1  g0044(.A1(new_n244), .A2(KEYINPUT3), .ZN(new_n245));
  INV_X1    g0045(.A(KEYINPUT3), .ZN(new_n246));
  NAND2_X1  g0046(.A1(new_n246), .A2(G33), .ZN(new_n247));
  NAND2_X1  g0047(.A1(new_n245), .A2(new_n247), .ZN(new_n248));
  NAND2_X1  g0048(.A1(new_n248), .A2(G77), .ZN(new_n249));
  XNOR2_X1  g0049(.A(KEYINPUT3), .B(G33), .ZN(new_n250));
  INV_X1    g0050(.A(G1698), .ZN(new_n251));
  NAND3_X1  g0051(.A1(new_n250), .A2(G222), .A3(new_n251), .ZN(new_n252));
  NAND2_X1  g0052(.A1(new_n250), .A2(G1698), .ZN(new_n253));
  XNOR2_X1  g0053(.A(new_n253), .B(KEYINPUT66), .ZN(new_n254));
  INV_X1    g0054(.A(G223), .ZN(new_n255));
  OAI211_X1 g0055(.A(new_n249), .B(new_n252), .C1(new_n254), .C2(new_n255), .ZN(new_n256));
  NAND2_X1  g0056(.A1(G33), .A2(G41), .ZN(new_n257));
  NAND3_X1  g0057(.A1(new_n257), .A2(G1), .A3(G13), .ZN(new_n258));
  INV_X1    g0058(.A(new_n258), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n256), .A2(new_n259), .ZN(new_n260));
  INV_X1    g0060(.A(G1), .ZN(new_n261));
  OAI21_X1  g0061(.A(new_n261), .B1(G41), .B2(G45), .ZN(new_n262));
  INV_X1    g0062(.A(new_n262), .ZN(new_n263));
  NAND3_X1  g0063(.A1(new_n263), .A2(new_n258), .A3(G274), .ZN(new_n264));
  INV_X1    g0064(.A(G226), .ZN(new_n265));
  NAND2_X1  g0065(.A1(new_n258), .A2(new_n262), .ZN(new_n266));
  OAI21_X1  g0066(.A(new_n264), .B1(new_n265), .B2(new_n266), .ZN(new_n267));
  XOR2_X1   g0067(.A(new_n267), .B(KEYINPUT65), .Z(new_n268));
  NAND2_X1  g0068(.A1(new_n260), .A2(new_n268), .ZN(new_n269));
  INV_X1    g0069(.A(new_n269), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n270), .A2(G190), .ZN(new_n271));
  NOR2_X1   g0071(.A1(G20), .A2(G33), .ZN(new_n272));
  AOI22_X1  g0072(.A1(new_n204), .A2(G20), .B1(G150), .B2(new_n272), .ZN(new_n273));
  XNOR2_X1  g0073(.A(KEYINPUT8), .B(G58), .ZN(new_n274));
  INV_X1    g0074(.A(KEYINPUT68), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n274), .A2(new_n275), .ZN(new_n276));
  OR3_X1    g0076(.A1(new_n275), .A2(new_n202), .A3(KEYINPUT8), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n276), .A2(new_n277), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n215), .A2(G33), .ZN(new_n279));
  OAI21_X1  g0079(.A(new_n273), .B1(new_n278), .B2(new_n279), .ZN(new_n280));
  OAI21_X1  g0080(.A(new_n214), .B1(new_n207), .B2(new_n244), .ZN(new_n281));
  NAND2_X1  g0081(.A1(new_n281), .A2(KEYINPUT67), .ZN(new_n282));
  INV_X1    g0082(.A(KEYINPUT67), .ZN(new_n283));
  OAI211_X1 g0083(.A(new_n283), .B(new_n214), .C1(new_n207), .C2(new_n244), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n282), .A2(new_n284), .ZN(new_n285));
  INV_X1    g0085(.A(new_n285), .ZN(new_n286));
  INV_X1    g0086(.A(G13), .ZN(new_n287));
  NOR3_X1   g0087(.A1(new_n287), .A2(new_n215), .A3(G1), .ZN(new_n288));
  AOI22_X1  g0088(.A1(new_n280), .A2(new_n286), .B1(new_n201), .B2(new_n288), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n261), .A2(G20), .ZN(new_n290));
  AND2_X1   g0090(.A1(new_n285), .A2(new_n290), .ZN(new_n291));
  INV_X1    g0091(.A(new_n291), .ZN(new_n292));
  OAI21_X1  g0092(.A(new_n289), .B1(new_n201), .B2(new_n292), .ZN(new_n293));
  INV_X1    g0093(.A(KEYINPUT9), .ZN(new_n294));
  OR2_X1    g0094(.A1(new_n293), .A2(new_n294), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n269), .A2(G200), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n293), .A2(new_n294), .ZN(new_n297));
  NAND4_X1  g0097(.A1(new_n271), .A2(new_n295), .A3(new_n296), .A4(new_n297), .ZN(new_n298));
  INV_X1    g0098(.A(KEYINPUT10), .ZN(new_n299));
  INV_X1    g0099(.A(KEYINPUT70), .ZN(new_n300));
  AOI21_X1  g0100(.A(new_n299), .B1(new_n296), .B2(new_n300), .ZN(new_n301));
  XNOR2_X1  g0101(.A(new_n298), .B(new_n301), .ZN(new_n302));
  INV_X1    g0102(.A(G179), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n270), .A2(new_n303), .ZN(new_n304));
  INV_X1    g0104(.A(G169), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n269), .A2(new_n305), .ZN(new_n306));
  NAND3_X1  g0106(.A1(new_n304), .A2(new_n293), .A3(new_n306), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n302), .A2(new_n307), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n203), .A2(G20), .ZN(new_n309));
  INV_X1    g0109(.A(G77), .ZN(new_n310));
  INV_X1    g0110(.A(new_n272), .ZN(new_n311));
  OAI221_X1 g0111(.A(new_n309), .B1(new_n279), .B2(new_n310), .C1(new_n311), .C2(new_n201), .ZN(new_n312));
  NAND3_X1  g0112(.A1(new_n286), .A2(KEYINPUT11), .A3(new_n312), .ZN(new_n313));
  NOR2_X1   g0113(.A1(new_n287), .A2(G1), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n314), .A2(KEYINPUT12), .ZN(new_n315));
  OAI221_X1 g0115(.A(new_n313), .B1(KEYINPUT12), .B2(new_n288), .C1(new_n309), .C2(new_n315), .ZN(new_n316));
  AOI21_X1  g0116(.A(new_n203), .B1(new_n292), .B2(KEYINPUT12), .ZN(new_n317));
  AOI21_X1  g0117(.A(KEYINPUT11), .B1(new_n286), .B2(new_n312), .ZN(new_n318));
  NOR3_X1   g0118(.A1(new_n316), .A2(new_n317), .A3(new_n318), .ZN(new_n319));
  INV_X1    g0119(.A(new_n319), .ZN(new_n320));
  NAND2_X1  g0120(.A1(new_n219), .A2(G1698), .ZN(new_n321));
  OAI211_X1 g0121(.A(new_n250), .B(new_n321), .C1(G226), .C2(G1698), .ZN(new_n322));
  NAND2_X1  g0122(.A1(G33), .A2(G97), .ZN(new_n323));
  AOI21_X1  g0123(.A(new_n258), .B1(new_n322), .B2(new_n323), .ZN(new_n324));
  OAI21_X1  g0124(.A(new_n264), .B1(new_n220), .B2(new_n266), .ZN(new_n325));
  NOR2_X1   g0125(.A1(new_n324), .A2(new_n325), .ZN(new_n326));
  XOR2_X1   g0126(.A(new_n326), .B(KEYINPUT13), .Z(new_n327));
  INV_X1    g0127(.A(KEYINPUT14), .ZN(new_n328));
  NAND3_X1  g0128(.A1(new_n327), .A2(new_n328), .A3(G169), .ZN(new_n329));
  OAI21_X1  g0129(.A(new_n329), .B1(new_n303), .B2(new_n327), .ZN(new_n330));
  AOI21_X1  g0130(.A(new_n328), .B1(new_n327), .B2(G169), .ZN(new_n331));
  OAI21_X1  g0131(.A(new_n320), .B1(new_n330), .B2(new_n331), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n291), .A2(G77), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n288), .A2(new_n310), .ZN(new_n334));
  NOR2_X1   g0134(.A1(new_n274), .A2(new_n311), .ZN(new_n335));
  XNOR2_X1  g0135(.A(KEYINPUT15), .B(G87), .ZN(new_n336));
  OAI22_X1  g0136(.A1(new_n336), .A2(new_n279), .B1(new_n215), .B2(new_n310), .ZN(new_n337));
  OAI21_X1  g0137(.A(new_n286), .B1(new_n335), .B2(new_n337), .ZN(new_n338));
  NAND3_X1  g0138(.A1(new_n333), .A2(new_n334), .A3(new_n338), .ZN(new_n339));
  NAND3_X1  g0139(.A1(new_n250), .A2(G232), .A3(new_n251), .ZN(new_n340));
  INV_X1    g0140(.A(KEYINPUT69), .ZN(new_n341));
  AOI22_X1  g0141(.A1(new_n340), .A2(new_n341), .B1(G107), .B2(new_n248), .ZN(new_n342));
  OAI221_X1 g0142(.A(new_n342), .B1(new_n341), .B2(new_n340), .C1(new_n254), .C2(new_n220), .ZN(new_n343));
  AND2_X1   g0143(.A1(new_n343), .A2(new_n259), .ZN(new_n344));
  INV_X1    g0144(.A(G244), .ZN(new_n345));
  OAI21_X1  g0145(.A(new_n264), .B1(new_n345), .B2(new_n266), .ZN(new_n346));
  NOR2_X1   g0146(.A1(new_n344), .A2(new_n346), .ZN(new_n347));
  AOI21_X1  g0147(.A(new_n339), .B1(new_n347), .B2(G190), .ZN(new_n348));
  INV_X1    g0148(.A(G200), .ZN(new_n349));
  OAI21_X1  g0149(.A(new_n348), .B1(new_n349), .B2(new_n347), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n327), .A2(G200), .ZN(new_n351));
  INV_X1    g0151(.A(G190), .ZN(new_n352));
  OAI211_X1 g0152(.A(new_n351), .B(new_n319), .C1(new_n352), .C2(new_n327), .ZN(new_n353));
  INV_X1    g0153(.A(new_n339), .ZN(new_n354));
  AOI21_X1  g0154(.A(new_n354), .B1(new_n347), .B2(new_n303), .ZN(new_n355));
  OAI21_X1  g0155(.A(new_n305), .B1(new_n344), .B2(new_n346), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n355), .A2(new_n356), .ZN(new_n357));
  NAND4_X1  g0157(.A1(new_n332), .A2(new_n350), .A3(new_n353), .A4(new_n357), .ZN(new_n358));
  INV_X1    g0158(.A(KEYINPUT16), .ZN(new_n359));
  NAND2_X1  g0159(.A1(G58), .A2(G68), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n360), .A2(KEYINPUT72), .ZN(new_n361));
  INV_X1    g0161(.A(KEYINPUT72), .ZN(new_n362));
  NAND3_X1  g0162(.A1(new_n362), .A2(G58), .A3(G68), .ZN(new_n363));
  NAND3_X1  g0163(.A1(new_n361), .A2(new_n363), .A3(new_n211), .ZN(new_n364));
  AOI22_X1  g0164(.A1(new_n364), .A2(G20), .B1(G159), .B2(new_n272), .ZN(new_n365));
  INV_X1    g0165(.A(KEYINPUT7), .ZN(new_n366));
  OAI21_X1  g0166(.A(new_n366), .B1(new_n250), .B2(G20), .ZN(new_n367));
  NAND3_X1  g0167(.A1(new_n248), .A2(KEYINPUT7), .A3(new_n215), .ZN(new_n368));
  AOI21_X1  g0168(.A(new_n203), .B1(new_n367), .B2(new_n368), .ZN(new_n369));
  OAI21_X1  g0169(.A(new_n365), .B1(new_n369), .B2(KEYINPUT73), .ZN(new_n370));
  INV_X1    g0170(.A(KEYINPUT73), .ZN(new_n371));
  AOI211_X1 g0171(.A(new_n371), .B(new_n203), .C1(new_n367), .C2(new_n368), .ZN(new_n372));
  OAI21_X1  g0172(.A(new_n359), .B1(new_n370), .B2(new_n372), .ZN(new_n373));
  OAI21_X1  g0173(.A(KEYINPUT71), .B1(new_n246), .B2(G33), .ZN(new_n374));
  INV_X1    g0174(.A(KEYINPUT71), .ZN(new_n375));
  NAND3_X1  g0175(.A1(new_n375), .A2(new_n244), .A3(KEYINPUT3), .ZN(new_n376));
  AND3_X1   g0176(.A1(new_n374), .A2(new_n376), .A3(new_n247), .ZN(new_n377));
  OAI21_X1  g0177(.A(KEYINPUT7), .B1(new_n377), .B2(G20), .ZN(new_n378));
  NAND3_X1  g0178(.A1(new_n374), .A2(new_n376), .A3(new_n247), .ZN(new_n379));
  NAND3_X1  g0179(.A1(new_n379), .A2(new_n366), .A3(new_n215), .ZN(new_n380));
  NAND3_X1  g0180(.A1(new_n378), .A2(G68), .A3(new_n380), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n365), .A2(KEYINPUT16), .ZN(new_n382));
  INV_X1    g0182(.A(new_n382), .ZN(new_n383));
  AOI21_X1  g0183(.A(new_n285), .B1(new_n381), .B2(new_n383), .ZN(new_n384));
  INV_X1    g0184(.A(KEYINPUT74), .ZN(new_n385));
  AOI21_X1  g0185(.A(new_n278), .B1(new_n285), .B2(new_n290), .ZN(new_n386));
  AOI21_X1  g0186(.A(new_n288), .B1(new_n276), .B2(new_n277), .ZN(new_n387));
  OAI21_X1  g0187(.A(new_n385), .B1(new_n386), .B2(new_n387), .ZN(new_n388));
  INV_X1    g0188(.A(new_n387), .ZN(new_n389));
  OAI211_X1 g0189(.A(KEYINPUT74), .B(new_n389), .C1(new_n291), .C2(new_n278), .ZN(new_n390));
  AOI22_X1  g0190(.A1(new_n373), .A2(new_n384), .B1(new_n388), .B2(new_n390), .ZN(new_n391));
  INV_X1    g0191(.A(new_n264), .ZN(new_n392));
  NAND3_X1  g0192(.A1(new_n258), .A2(G232), .A3(new_n262), .ZN(new_n393));
  INV_X1    g0193(.A(KEYINPUT75), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n393), .A2(new_n394), .ZN(new_n395));
  NAND4_X1  g0195(.A1(new_n258), .A2(new_n262), .A3(KEYINPUT75), .A4(G232), .ZN(new_n396));
  AOI21_X1  g0196(.A(new_n392), .B1(new_n395), .B2(new_n396), .ZN(new_n397));
  NAND2_X1  g0197(.A1(G33), .A2(G87), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n265), .A2(G1698), .ZN(new_n399));
  OAI21_X1  g0199(.A(new_n399), .B1(G223), .B2(G1698), .ZN(new_n400));
  OAI21_X1  g0200(.A(new_n398), .B1(new_n379), .B2(new_n400), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n401), .A2(new_n259), .ZN(new_n402));
  AOI21_X1  g0202(.A(new_n305), .B1(new_n397), .B2(new_n402), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n395), .A2(new_n396), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n404), .A2(new_n264), .ZN(new_n405));
  NOR2_X1   g0205(.A1(G223), .A2(G1698), .ZN(new_n406));
  AOI21_X1  g0206(.A(new_n406), .B1(new_n265), .B2(G1698), .ZN(new_n407));
  NAND4_X1  g0207(.A1(new_n407), .A2(new_n374), .A3(new_n247), .A4(new_n376), .ZN(new_n408));
  AOI21_X1  g0208(.A(new_n258), .B1(new_n408), .B2(new_n398), .ZN(new_n409));
  NOR2_X1   g0209(.A1(new_n405), .A2(new_n409), .ZN(new_n410));
  AOI21_X1  g0210(.A(new_n403), .B1(G179), .B2(new_n410), .ZN(new_n411));
  OAI21_X1  g0211(.A(KEYINPUT18), .B1(new_n391), .B2(new_n411), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n388), .A2(new_n390), .ZN(new_n413));
  NAND2_X1  g0213(.A1(new_n364), .A2(G20), .ZN(new_n414));
  INV_X1    g0214(.A(G159), .ZN(new_n415));
  OAI21_X1  g0215(.A(new_n414), .B1(new_n415), .B2(new_n311), .ZN(new_n416));
  AOI21_X1  g0216(.A(KEYINPUT7), .B1(new_n248), .B2(new_n215), .ZN(new_n417));
  AOI211_X1 g0217(.A(new_n366), .B(G20), .C1(new_n245), .C2(new_n247), .ZN(new_n418));
  OAI21_X1  g0218(.A(G68), .B1(new_n417), .B2(new_n418), .ZN(new_n419));
  AOI21_X1  g0219(.A(new_n416), .B1(new_n419), .B2(new_n371), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n369), .A2(KEYINPUT73), .ZN(new_n421));
  AOI21_X1  g0221(.A(KEYINPUT16), .B1(new_n420), .B2(new_n421), .ZN(new_n422));
  AND3_X1   g0222(.A1(new_n379), .A2(new_n366), .A3(new_n215), .ZN(new_n423));
  AOI21_X1  g0223(.A(new_n366), .B1(new_n379), .B2(new_n215), .ZN(new_n424));
  NOR3_X1   g0224(.A1(new_n423), .A2(new_n424), .A3(new_n203), .ZN(new_n425));
  OAI21_X1  g0225(.A(new_n286), .B1(new_n425), .B2(new_n382), .ZN(new_n426));
  OAI21_X1  g0226(.A(new_n413), .B1(new_n422), .B2(new_n426), .ZN(new_n427));
  INV_X1    g0227(.A(KEYINPUT18), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n410), .A2(G179), .ZN(new_n429));
  OAI21_X1  g0229(.A(new_n429), .B1(new_n305), .B2(new_n410), .ZN(new_n430));
  NAND3_X1  g0230(.A1(new_n427), .A2(new_n428), .A3(new_n430), .ZN(new_n431));
  AND2_X1   g0231(.A1(new_n412), .A2(new_n431), .ZN(new_n432));
  OAI21_X1  g0232(.A(new_n349), .B1(new_n405), .B2(new_n409), .ZN(new_n433));
  NAND3_X1  g0233(.A1(new_n397), .A2(new_n402), .A3(new_n352), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n433), .A2(new_n434), .ZN(new_n435));
  OAI211_X1 g0235(.A(new_n435), .B(new_n413), .C1(new_n422), .C2(new_n426), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n436), .A2(KEYINPUT17), .ZN(new_n437));
  INV_X1    g0237(.A(KEYINPUT17), .ZN(new_n438));
  NAND3_X1  g0238(.A1(new_n391), .A2(new_n438), .A3(new_n435), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n437), .A2(new_n439), .ZN(new_n440));
  NAND2_X1  g0240(.A1(new_n432), .A2(new_n440), .ZN(new_n441));
  NOR3_X1   g0241(.A1(new_n308), .A2(new_n358), .A3(new_n441), .ZN(new_n442));
  NAND3_X1  g0242(.A1(new_n377), .A2(new_n215), .A3(G68), .ZN(new_n443));
  INV_X1    g0243(.A(G87), .ZN(new_n444));
  INV_X1    g0244(.A(G97), .ZN(new_n445));
  INV_X1    g0245(.A(G107), .ZN(new_n446));
  NAND3_X1  g0246(.A1(new_n444), .A2(new_n445), .A3(new_n446), .ZN(new_n447));
  NAND2_X1  g0247(.A1(new_n323), .A2(new_n215), .ZN(new_n448));
  NAND3_X1  g0248(.A1(new_n447), .A2(new_n448), .A3(KEYINPUT19), .ZN(new_n449));
  NOR2_X1   g0249(.A1(new_n279), .A2(new_n445), .ZN(new_n450));
  OAI211_X1 g0250(.A(new_n443), .B(new_n449), .C1(KEYINPUT19), .C2(new_n450), .ZN(new_n451));
  AOI22_X1  g0251(.A1(new_n451), .A2(new_n286), .B1(new_n288), .B2(new_n336), .ZN(new_n452));
  INV_X1    g0252(.A(new_n452), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n345), .A2(G1698), .ZN(new_n454));
  OAI21_X1  g0254(.A(new_n454), .B1(G238), .B2(G1698), .ZN(new_n455));
  INV_X1    g0255(.A(G116), .ZN(new_n456));
  OAI22_X1  g0256(.A1(new_n379), .A2(new_n455), .B1(new_n244), .B2(new_n456), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n457), .A2(new_n259), .ZN(new_n458));
  AND2_X1   g0258(.A1(new_n261), .A2(G45), .ZN(new_n459));
  INV_X1    g0259(.A(G274), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  OAI211_X1 g0261(.A(new_n461), .B(new_n258), .C1(G250), .C2(new_n459), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n458), .A2(new_n462), .ZN(new_n463));
  INV_X1    g0263(.A(KEYINPUT78), .ZN(new_n464));
  XNOR2_X1  g0264(.A(new_n463), .B(new_n464), .ZN(new_n465));
  AOI21_X1  g0265(.A(new_n453), .B1(new_n465), .B2(G190), .ZN(new_n466));
  AOI21_X1  g0266(.A(new_n288), .B1(new_n261), .B2(G33), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n285), .A2(new_n467), .ZN(new_n468));
  NOR2_X1   g0268(.A1(new_n468), .A2(new_n444), .ZN(new_n469));
  INV_X1    g0269(.A(new_n469), .ZN(new_n470));
  XNOR2_X1  g0270(.A(new_n463), .B(KEYINPUT78), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n471), .A2(G200), .ZN(new_n472));
  AND3_X1   g0272(.A1(new_n466), .A2(new_n470), .A3(new_n472), .ZN(new_n473));
  INV_X1    g0273(.A(new_n468), .ZN(new_n474));
  INV_X1    g0274(.A(new_n336), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n474), .A2(new_n475), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n452), .A2(new_n476), .ZN(new_n477));
  INV_X1    g0277(.A(new_n477), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n465), .A2(new_n303), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n471), .A2(new_n305), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n479), .A2(new_n480), .ZN(new_n481));
  INV_X1    g0281(.A(KEYINPUT79), .ZN(new_n482));
  AOI21_X1  g0282(.A(new_n478), .B1(new_n481), .B2(new_n482), .ZN(new_n483));
  NAND3_X1  g0283(.A1(new_n479), .A2(new_n480), .A3(KEYINPUT79), .ZN(new_n484));
  AOI21_X1  g0284(.A(new_n473), .B1(new_n483), .B2(new_n484), .ZN(new_n485));
  NOR2_X1   g0285(.A1(new_n468), .A2(new_n446), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n288), .A2(new_n446), .ZN(new_n487));
  XNOR2_X1  g0287(.A(new_n487), .B(KEYINPUT25), .ZN(new_n488));
  NOR2_X1   g0288(.A1(new_n486), .A2(new_n488), .ZN(new_n489));
  INV_X1    g0289(.A(new_n489), .ZN(new_n490));
  NOR3_X1   g0290(.A1(new_n244), .A2(new_n456), .A3(G20), .ZN(new_n491));
  INV_X1    g0291(.A(KEYINPUT23), .ZN(new_n492));
  OAI21_X1  g0292(.A(new_n492), .B1(new_n215), .B2(G107), .ZN(new_n493));
  NAND3_X1  g0293(.A1(new_n446), .A2(KEYINPUT23), .A3(G20), .ZN(new_n494));
  AOI21_X1  g0294(.A(new_n491), .B1(new_n493), .B2(new_n494), .ZN(new_n495));
  NAND3_X1  g0295(.A1(new_n215), .A2(KEYINPUT22), .A3(G87), .ZN(new_n496));
  NOR3_X1   g0296(.A1(new_n248), .A2(G20), .A3(new_n444), .ZN(new_n497));
  OAI221_X1 g0297(.A(new_n495), .B1(new_n379), .B2(new_n496), .C1(new_n497), .C2(KEYINPUT22), .ZN(new_n498));
  XNOR2_X1  g0298(.A(new_n498), .B(KEYINPUT24), .ZN(new_n499));
  AOI21_X1  g0299(.A(new_n490), .B1(new_n499), .B2(new_n286), .ZN(new_n500));
  INV_X1    g0300(.A(G257), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n501), .A2(G1698), .ZN(new_n502));
  OAI21_X1  g0302(.A(new_n502), .B1(G250), .B2(G1698), .ZN(new_n503));
  INV_X1    g0303(.A(G294), .ZN(new_n504));
  OAI22_X1  g0304(.A1(new_n379), .A2(new_n503), .B1(new_n244), .B2(new_n504), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n505), .A2(new_n259), .ZN(new_n506));
  INV_X1    g0306(.A(KEYINPUT5), .ZN(new_n507));
  OAI211_X1 g0307(.A(new_n261), .B(G45), .C1(new_n507), .C2(G41), .ZN(new_n508));
  INV_X1    g0308(.A(G41), .ZN(new_n509));
  NOR2_X1   g0309(.A1(new_n509), .A2(KEYINPUT5), .ZN(new_n510));
  NOR2_X1   g0310(.A1(new_n508), .A2(new_n510), .ZN(new_n511));
  NAND3_X1  g0311(.A1(new_n511), .A2(G274), .A3(new_n258), .ZN(new_n512));
  OAI21_X1  g0312(.A(new_n258), .B1(new_n508), .B2(new_n510), .ZN(new_n513));
  INV_X1    g0313(.A(new_n513), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n514), .A2(G264), .ZN(new_n515));
  AND3_X1   g0315(.A1(new_n506), .A2(new_n512), .A3(new_n515), .ZN(new_n516));
  OR2_X1    g0316(.A1(new_n516), .A2(KEYINPUT81), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n516), .A2(KEYINPUT81), .ZN(new_n518));
  NAND3_X1  g0318(.A1(new_n517), .A2(G169), .A3(new_n518), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n516), .A2(G179), .ZN(new_n520));
  AOI21_X1  g0320(.A(new_n500), .B1(new_n519), .B2(new_n520), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n517), .A2(new_n518), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n522), .A2(new_n352), .ZN(new_n523));
  NOR2_X1   g0323(.A1(new_n516), .A2(G200), .ZN(new_n524));
  INV_X1    g0324(.A(new_n524), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n523), .A2(new_n525), .ZN(new_n526));
  AOI21_X1  g0326(.A(new_n521), .B1(new_n526), .B2(new_n500), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n474), .A2(G116), .ZN(new_n528));
  AOI21_X1  g0328(.A(G20), .B1(G33), .B2(G283), .ZN(new_n529));
  OAI21_X1  g0329(.A(new_n529), .B1(G33), .B2(new_n445), .ZN(new_n530));
  OAI211_X1 g0330(.A(new_n530), .B(new_n281), .C1(new_n215), .C2(G116), .ZN(new_n531));
  INV_X1    g0331(.A(KEYINPUT20), .ZN(new_n532));
  XNOR2_X1  g0332(.A(new_n531), .B(new_n532), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n288), .A2(new_n456), .ZN(new_n534));
  NAND3_X1  g0334(.A1(new_n528), .A2(new_n533), .A3(new_n534), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n514), .A2(G270), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n536), .A2(new_n512), .ZN(new_n537));
  MUX2_X1   g0337(.A(G257), .B(G264), .S(G1698), .Z(new_n538));
  NAND2_X1  g0338(.A1(new_n377), .A2(new_n538), .ZN(new_n539));
  XOR2_X1   g0339(.A(KEYINPUT80), .B(G303), .Z(new_n540));
  INV_X1    g0340(.A(new_n540), .ZN(new_n541));
  NAND2_X1  g0341(.A1(new_n541), .A2(new_n248), .ZN(new_n542));
  AOI21_X1  g0342(.A(new_n258), .B1(new_n539), .B2(new_n542), .ZN(new_n543));
  OR2_X1    g0343(.A1(new_n537), .A2(new_n543), .ZN(new_n544));
  NAND4_X1  g0344(.A1(new_n535), .A2(new_n544), .A3(KEYINPUT21), .A4(G169), .ZN(new_n545));
  NOR3_X1   g0345(.A1(new_n537), .A2(new_n543), .A3(new_n303), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n535), .A2(new_n546), .ZN(new_n547));
  AND2_X1   g0347(.A1(new_n545), .A2(new_n547), .ZN(new_n548));
  AOI21_X1  g0348(.A(new_n535), .B1(new_n544), .B2(G200), .ZN(new_n549));
  OAI21_X1  g0349(.A(new_n549), .B1(new_n352), .B2(new_n544), .ZN(new_n550));
  NAND3_X1  g0350(.A1(new_n535), .A2(new_n544), .A3(G169), .ZN(new_n551));
  INV_X1    g0351(.A(KEYINPUT21), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  NAND3_X1  g0353(.A1(new_n548), .A2(new_n550), .A3(new_n553), .ZN(new_n554));
  INV_X1    g0354(.A(KEYINPUT6), .ZN(new_n555));
  NOR2_X1   g0355(.A1(new_n445), .A2(new_n446), .ZN(new_n556));
  NOR2_X1   g0356(.A1(G97), .A2(G107), .ZN(new_n557));
  OAI21_X1  g0357(.A(new_n555), .B1(new_n556), .B2(new_n557), .ZN(new_n558));
  NAND3_X1  g0358(.A1(new_n446), .A2(KEYINPUT6), .A3(G97), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n560), .A2(G20), .ZN(new_n561));
  OAI21_X1  g0361(.A(new_n561), .B1(new_n310), .B2(new_n311), .ZN(new_n562));
  AOI21_X1  g0362(.A(new_n446), .B1(new_n367), .B2(new_n368), .ZN(new_n563));
  OAI21_X1  g0363(.A(new_n286), .B1(new_n562), .B2(new_n563), .ZN(new_n564));
  INV_X1    g0364(.A(new_n288), .ZN(new_n565));
  NOR2_X1   g0365(.A1(new_n565), .A2(G97), .ZN(new_n566));
  AOI21_X1  g0366(.A(new_n566), .B1(new_n474), .B2(G97), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n564), .A2(new_n567), .ZN(new_n568));
  INV_X1    g0368(.A(KEYINPUT77), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n568), .A2(new_n569), .ZN(new_n570));
  OAI21_X1  g0370(.A(new_n512), .B1(new_n513), .B2(new_n501), .ZN(new_n571));
  INV_X1    g0371(.A(KEYINPUT4), .ZN(new_n572));
  OAI21_X1  g0372(.A(new_n572), .B1(new_n379), .B2(new_n345), .ZN(new_n573));
  NOR3_X1   g0373(.A1(new_n572), .A2(new_n345), .A3(G1698), .ZN(new_n574));
  AOI22_X1  g0374(.A1(new_n250), .A2(new_n574), .B1(G33), .B2(G283), .ZN(new_n575));
  AOI21_X1  g0375(.A(new_n572), .B1(new_n250), .B2(G250), .ZN(new_n576));
  OAI211_X1 g0376(.A(new_n573), .B(new_n575), .C1(new_n251), .C2(new_n576), .ZN(new_n577));
  AOI21_X1  g0377(.A(new_n571), .B1(new_n577), .B2(new_n259), .ZN(new_n578));
  INV_X1    g0378(.A(new_n578), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n579), .A2(new_n305), .ZN(new_n580));
  INV_X1    g0380(.A(KEYINPUT76), .ZN(new_n581));
  OR2_X1    g0381(.A1(new_n571), .A2(new_n581), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n577), .A2(new_n259), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n571), .A2(new_n581), .ZN(new_n584));
  NAND4_X1  g0384(.A1(new_n582), .A2(new_n303), .A3(new_n583), .A4(new_n584), .ZN(new_n585));
  NAND3_X1  g0385(.A1(new_n564), .A2(KEYINPUT77), .A3(new_n567), .ZN(new_n586));
  NAND4_X1  g0386(.A1(new_n570), .A2(new_n580), .A3(new_n585), .A4(new_n586), .ZN(new_n587));
  NAND3_X1  g0387(.A1(new_n582), .A2(new_n583), .A3(new_n584), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n588), .A2(G200), .ZN(new_n589));
  INV_X1    g0389(.A(new_n568), .ZN(new_n590));
  OAI211_X1 g0390(.A(new_n589), .B(new_n590), .C1(new_n352), .C2(new_n579), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n587), .A2(new_n591), .ZN(new_n592));
  NOR2_X1   g0392(.A1(new_n554), .A2(new_n592), .ZN(new_n593));
  AND4_X1   g0393(.A1(new_n442), .A2(new_n485), .A3(new_n527), .A4(new_n593), .ZN(G372));
  NAND2_X1  g0394(.A1(new_n463), .A2(new_n305), .ZN(new_n595));
  OAI211_X1 g0395(.A(new_n477), .B(new_n595), .C1(new_n471), .C2(G179), .ZN(new_n596));
  AOI21_X1  g0396(.A(new_n469), .B1(new_n463), .B2(G200), .ZN(new_n597));
  OAI211_X1 g0397(.A(new_n452), .B(new_n597), .C1(new_n471), .C2(new_n352), .ZN(new_n598));
  AND2_X1   g0398(.A1(new_n596), .A2(new_n598), .ZN(new_n599));
  AOI21_X1  g0399(.A(G190), .B1(new_n517), .B2(new_n518), .ZN(new_n600));
  OAI21_X1  g0400(.A(new_n500), .B1(new_n600), .B2(new_n524), .ZN(new_n601));
  NAND4_X1  g0401(.A1(new_n599), .A2(new_n601), .A3(new_n587), .A4(new_n591), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n548), .A2(new_n553), .ZN(new_n603));
  NOR2_X1   g0403(.A1(new_n603), .A2(new_n521), .ZN(new_n604));
  OAI21_X1  g0404(.A(new_n596), .B1(new_n602), .B2(new_n604), .ZN(new_n605));
  INV_X1    g0405(.A(new_n605), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n596), .A2(new_n598), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n580), .A2(new_n585), .ZN(new_n608));
  NOR4_X1   g0408(.A1(new_n607), .A2(KEYINPUT26), .A3(new_n608), .A4(new_n590), .ZN(new_n609));
  NOR2_X1   g0409(.A1(new_n471), .A2(G179), .ZN(new_n610));
  NOR2_X1   g0410(.A1(new_n465), .A2(G169), .ZN(new_n611));
  OAI21_X1  g0411(.A(new_n482), .B1(new_n610), .B2(new_n611), .ZN(new_n612));
  NAND3_X1  g0412(.A1(new_n612), .A2(new_n484), .A3(new_n477), .ZN(new_n613));
  INV_X1    g0413(.A(new_n473), .ZN(new_n614));
  INV_X1    g0414(.A(new_n587), .ZN(new_n615));
  NAND3_X1  g0415(.A1(new_n613), .A2(new_n614), .A3(new_n615), .ZN(new_n616));
  AOI21_X1  g0416(.A(new_n609), .B1(new_n616), .B2(KEYINPUT26), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n606), .A2(new_n617), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n442), .A2(new_n618), .ZN(new_n619));
  INV_X1    g0419(.A(new_n307), .ZN(new_n620));
  NAND3_X1  g0420(.A1(new_n353), .A2(new_n355), .A3(new_n356), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n332), .A2(new_n621), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n622), .A2(new_n440), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n412), .A2(new_n431), .ZN(new_n624));
  INV_X1    g0424(.A(KEYINPUT82), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  NAND3_X1  g0426(.A1(new_n412), .A2(new_n431), .A3(KEYINPUT82), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n623), .A2(new_n628), .ZN(new_n629));
  AOI21_X1  g0429(.A(new_n620), .B1(new_n629), .B2(new_n302), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n619), .A2(new_n630), .ZN(G369));
  NAND2_X1  g0431(.A1(new_n314), .A2(new_n215), .ZN(new_n632));
  OR2_X1    g0432(.A1(new_n632), .A2(KEYINPUT27), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n632), .A2(KEYINPUT27), .ZN(new_n634));
  NAND3_X1  g0434(.A1(new_n633), .A2(new_n634), .A3(G213), .ZN(new_n635));
  INV_X1    g0435(.A(G343), .ZN(new_n636));
  NOR2_X1   g0436(.A1(new_n635), .A2(new_n636), .ZN(new_n637));
  AND2_X1   g0437(.A1(new_n535), .A2(new_n637), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n603), .A2(new_n638), .ZN(new_n639));
  OAI21_X1  g0439(.A(new_n639), .B1(new_n554), .B2(new_n638), .ZN(new_n640));
  XOR2_X1   g0440(.A(new_n640), .B(KEYINPUT83), .Z(new_n641));
  AND2_X1   g0441(.A1(new_n641), .A2(G330), .ZN(new_n642));
  INV_X1    g0442(.A(new_n637), .ZN(new_n643));
  OAI21_X1  g0443(.A(new_n527), .B1(new_n500), .B2(new_n643), .ZN(new_n644));
  INV_X1    g0444(.A(new_n521), .ZN(new_n645));
  OAI21_X1  g0445(.A(new_n644), .B1(new_n645), .B2(new_n643), .ZN(new_n646));
  INV_X1    g0446(.A(KEYINPUT84), .ZN(new_n647));
  XNOR2_X1  g0447(.A(new_n646), .B(new_n647), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n642), .A2(new_n648), .ZN(new_n649));
  XOR2_X1   g0449(.A(new_n649), .B(KEYINPUT85), .Z(new_n650));
  INV_X1    g0450(.A(new_n650), .ZN(new_n651));
  AOI21_X1  g0451(.A(new_n637), .B1(new_n548), .B2(new_n553), .ZN(new_n652));
  AOI22_X1  g0452(.A1(new_n648), .A2(new_n652), .B1(new_n521), .B2(new_n643), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n651), .A2(new_n653), .ZN(G399));
  INV_X1    g0454(.A(new_n208), .ZN(new_n655));
  NOR2_X1   g0455(.A1(new_n655), .A2(G41), .ZN(new_n656));
  INV_X1    g0456(.A(new_n656), .ZN(new_n657));
  NOR2_X1   g0457(.A1(new_n447), .A2(G116), .ZN(new_n658));
  NAND3_X1  g0458(.A1(new_n657), .A2(G1), .A3(new_n658), .ZN(new_n659));
  OAI21_X1  g0459(.A(new_n659), .B1(new_n212), .B2(new_n657), .ZN(new_n660));
  XNOR2_X1  g0460(.A(new_n660), .B(KEYINPUT28), .ZN(new_n661));
  INV_X1    g0461(.A(KEYINPUT26), .ZN(new_n662));
  NOR4_X1   g0462(.A1(new_n607), .A2(new_n662), .A3(new_n608), .A4(new_n590), .ZN(new_n663));
  AOI21_X1  g0463(.A(new_n663), .B1(new_n616), .B2(new_n662), .ZN(new_n664));
  OAI211_X1 g0464(.A(KEYINPUT29), .B(new_n643), .C1(new_n664), .C2(new_n605), .ZN(new_n665));
  AOI21_X1  g0465(.A(new_n637), .B1(new_n606), .B2(new_n617), .ZN(new_n666));
  OAI21_X1  g0466(.A(new_n665), .B1(new_n666), .B2(KEYINPUT29), .ZN(new_n667));
  NAND4_X1  g0467(.A1(new_n485), .A2(new_n593), .A3(new_n527), .A4(new_n643), .ZN(new_n668));
  AND2_X1   g0468(.A1(new_n506), .A2(new_n515), .ZN(new_n669));
  NAND3_X1  g0469(.A1(new_n546), .A2(new_n669), .A3(new_n578), .ZN(new_n670));
  INV_X1    g0470(.A(KEYINPUT30), .ZN(new_n671));
  OR3_X1    g0471(.A1(new_n670), .A2(new_n471), .A3(new_n671), .ZN(new_n672));
  INV_X1    g0472(.A(new_n516), .ZN(new_n673));
  AOI21_X1  g0473(.A(G179), .B1(new_n458), .B2(new_n462), .ZN(new_n674));
  NAND4_X1  g0474(.A1(new_n588), .A2(new_n673), .A3(new_n544), .A4(new_n674), .ZN(new_n675));
  OAI21_X1  g0475(.A(new_n671), .B1(new_n670), .B2(new_n471), .ZN(new_n676));
  NAND3_X1  g0476(.A1(new_n672), .A2(new_n675), .A3(new_n676), .ZN(new_n677));
  AOI21_X1  g0477(.A(KEYINPUT31), .B1(new_n677), .B2(new_n637), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n678), .A2(KEYINPUT86), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n668), .A2(new_n679), .ZN(new_n680));
  NAND3_X1  g0480(.A1(new_n677), .A2(KEYINPUT31), .A3(new_n637), .ZN(new_n681));
  AOI21_X1  g0481(.A(new_n678), .B1(KEYINPUT86), .B2(new_n681), .ZN(new_n682));
  OAI21_X1  g0482(.A(G330), .B1(new_n680), .B2(new_n682), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n667), .A2(new_n683), .ZN(new_n684));
  INV_X1    g0484(.A(new_n684), .ZN(new_n685));
  OAI21_X1  g0485(.A(new_n661), .B1(new_n685), .B2(G1), .ZN(G364));
  NOR2_X1   g0486(.A1(new_n287), .A2(G20), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n687), .A2(G45), .ZN(new_n688));
  NAND3_X1  g0488(.A1(new_n657), .A2(G1), .A3(new_n688), .ZN(new_n689));
  INV_X1    g0489(.A(new_n689), .ZN(new_n690));
  NOR2_X1   g0490(.A1(new_n642), .A2(new_n690), .ZN(new_n691));
  OAI21_X1  g0491(.A(new_n691), .B1(G330), .B2(new_n641), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n379), .A2(new_n208), .ZN(new_n693));
  XOR2_X1   g0493(.A(new_n693), .B(KEYINPUT87), .Z(new_n694));
  NAND2_X1  g0494(.A1(new_n239), .A2(G45), .ZN(new_n695));
  OAI211_X1 g0495(.A(new_n694), .B(new_n695), .C1(G45), .C2(new_n212), .ZN(new_n696));
  INV_X1    g0496(.A(G355), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n250), .A2(new_n208), .ZN(new_n698));
  OAI221_X1 g0498(.A(new_n696), .B1(G116), .B2(new_n208), .C1(new_n697), .C2(new_n698), .ZN(new_n699));
  NOR2_X1   g0499(.A1(G13), .A2(G33), .ZN(new_n700));
  INV_X1    g0500(.A(new_n700), .ZN(new_n701));
  NOR2_X1   g0501(.A1(new_n701), .A2(G20), .ZN(new_n702));
  AOI21_X1  g0502(.A(new_n214), .B1(G20), .B2(new_n305), .ZN(new_n703));
  NOR2_X1   g0503(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  AOI21_X1  g0504(.A(new_n689), .B1(new_n699), .B2(new_n704), .ZN(new_n705));
  INV_X1    g0505(.A(new_n703), .ZN(new_n706));
  NOR2_X1   g0506(.A1(new_n215), .A2(new_n303), .ZN(new_n707));
  XNOR2_X1  g0507(.A(new_n707), .B(KEYINPUT88), .ZN(new_n708));
  NOR2_X1   g0508(.A1(G190), .A2(G200), .ZN(new_n709));
  NAND2_X1  g0509(.A1(new_n708), .A2(new_n709), .ZN(new_n710));
  INV_X1    g0510(.A(new_n710), .ZN(new_n711));
  NOR2_X1   g0511(.A1(new_n352), .A2(G200), .ZN(new_n712));
  NAND2_X1  g0512(.A1(new_n708), .A2(new_n712), .ZN(new_n713));
  INV_X1    g0513(.A(new_n713), .ZN(new_n714));
  AOI22_X1  g0514(.A1(G311), .A2(new_n711), .B1(new_n714), .B2(G322), .ZN(new_n715));
  NOR2_X1   g0515(.A1(new_n349), .A2(G179), .ZN(new_n716));
  NAND3_X1  g0516(.A1(new_n716), .A2(G20), .A3(new_n352), .ZN(new_n717));
  INV_X1    g0517(.A(KEYINPUT90), .ZN(new_n718));
  OR2_X1    g0518(.A1(new_n717), .A2(new_n718), .ZN(new_n719));
  NAND2_X1  g0519(.A1(new_n717), .A2(new_n718), .ZN(new_n720));
  NAND2_X1  g0520(.A1(new_n719), .A2(new_n720), .ZN(new_n721));
  INV_X1    g0521(.A(new_n721), .ZN(new_n722));
  NAND3_X1  g0522(.A1(new_n709), .A2(G20), .A3(new_n303), .ZN(new_n723));
  OR2_X1    g0523(.A1(new_n723), .A2(KEYINPUT89), .ZN(new_n724));
  NAND2_X1  g0524(.A1(new_n723), .A2(KEYINPUT89), .ZN(new_n725));
  NAND2_X1  g0525(.A1(new_n724), .A2(new_n725), .ZN(new_n726));
  INV_X1    g0526(.A(new_n726), .ZN(new_n727));
  AOI22_X1  g0527(.A1(new_n722), .A2(G283), .B1(new_n727), .B2(G329), .ZN(new_n728));
  NAND2_X1  g0528(.A1(new_n715), .A2(new_n728), .ZN(new_n729));
  INV_X1    g0529(.A(G303), .ZN(new_n730));
  NAND3_X1  g0530(.A1(new_n716), .A2(G20), .A3(G190), .ZN(new_n731));
  NAND2_X1  g0531(.A1(new_n707), .A2(G200), .ZN(new_n732));
  NOR2_X1   g0532(.A1(new_n732), .A2(new_n352), .ZN(new_n733));
  INV_X1    g0533(.A(new_n733), .ZN(new_n734));
  INV_X1    g0534(.A(G326), .ZN(new_n735));
  OAI221_X1 g0535(.A(new_n248), .B1(new_n730), .B2(new_n731), .C1(new_n734), .C2(new_n735), .ZN(new_n736));
  NOR2_X1   g0536(.A1(new_n732), .A2(G190), .ZN(new_n737));
  INV_X1    g0537(.A(G317), .ZN(new_n738));
  NAND2_X1  g0538(.A1(new_n738), .A2(KEYINPUT33), .ZN(new_n739));
  OR2_X1    g0539(.A1(new_n738), .A2(KEYINPUT33), .ZN(new_n740));
  NAND3_X1  g0540(.A1(new_n737), .A2(new_n739), .A3(new_n740), .ZN(new_n741));
  AOI21_X1  g0541(.A(new_n215), .B1(new_n712), .B2(new_n303), .ZN(new_n742));
  OAI21_X1  g0542(.A(new_n741), .B1(new_n504), .B2(new_n742), .ZN(new_n743));
  NOR3_X1   g0543(.A1(new_n729), .A2(new_n736), .A3(new_n743), .ZN(new_n744));
  XOR2_X1   g0544(.A(new_n742), .B(KEYINPUT92), .Z(new_n745));
  INV_X1    g0545(.A(new_n745), .ZN(new_n746));
  NOR2_X1   g0546(.A1(new_n746), .A2(new_n445), .ZN(new_n747));
  AOI22_X1  g0547(.A1(new_n737), .A2(G68), .B1(new_n733), .B2(G50), .ZN(new_n748));
  OAI221_X1 g0548(.A(new_n748), .B1(new_n713), .B2(new_n202), .C1(new_n310), .C2(new_n710), .ZN(new_n749));
  INV_X1    g0549(.A(KEYINPUT32), .ZN(new_n750));
  OAI21_X1  g0550(.A(new_n750), .B1(new_n726), .B2(new_n415), .ZN(new_n751));
  NAND3_X1  g0551(.A1(new_n727), .A2(KEYINPUT32), .A3(G159), .ZN(new_n752));
  AOI211_X1 g0552(.A(new_n747), .B(new_n749), .C1(new_n751), .C2(new_n752), .ZN(new_n753));
  NOR2_X1   g0553(.A1(new_n721), .A2(new_n446), .ZN(new_n754));
  NOR2_X1   g0554(.A1(new_n731), .A2(new_n444), .ZN(new_n755));
  NOR3_X1   g0555(.A1(new_n754), .A2(new_n248), .A3(new_n755), .ZN(new_n756));
  XNOR2_X1  g0556(.A(new_n756), .B(KEYINPUT91), .ZN(new_n757));
  AOI21_X1  g0557(.A(new_n744), .B1(new_n753), .B2(new_n757), .ZN(new_n758));
  INV_X1    g0558(.A(new_n702), .ZN(new_n759));
  OAI221_X1 g0559(.A(new_n705), .B1(new_n706), .B2(new_n758), .C1(new_n641), .C2(new_n759), .ZN(new_n760));
  NAND2_X1  g0560(.A1(new_n692), .A2(new_n760), .ZN(G396));
  AOI22_X1  g0561(.A1(new_n737), .A2(G150), .B1(new_n733), .B2(G137), .ZN(new_n762));
  INV_X1    g0562(.A(G143), .ZN(new_n763));
  OAI221_X1 g0563(.A(new_n762), .B1(new_n713), .B2(new_n763), .C1(new_n415), .C2(new_n710), .ZN(new_n764));
  XNOR2_X1  g0564(.A(new_n764), .B(KEYINPUT94), .ZN(new_n765));
  INV_X1    g0565(.A(KEYINPUT34), .ZN(new_n766));
  AND2_X1   g0566(.A1(new_n765), .A2(new_n766), .ZN(new_n767));
  NOR2_X1   g0567(.A1(new_n765), .A2(new_n766), .ZN(new_n768));
  OAI221_X1 g0568(.A(new_n377), .B1(new_n731), .B2(new_n201), .C1(new_n202), .C2(new_n742), .ZN(new_n769));
  INV_X1    g0569(.A(G132), .ZN(new_n770));
  OAI22_X1  g0570(.A1(new_n721), .A2(new_n203), .B1(new_n770), .B2(new_n726), .ZN(new_n771));
  NOR4_X1   g0571(.A1(new_n767), .A2(new_n768), .A3(new_n769), .A4(new_n771), .ZN(new_n772));
  OAI221_X1 g0572(.A(new_n248), .B1(new_n446), .B2(new_n731), .C1(new_n734), .C2(new_n730), .ZN(new_n773));
  AOI211_X1 g0573(.A(new_n773), .B(new_n747), .C1(G283), .C2(new_n737), .ZN(new_n774));
  NOR2_X1   g0574(.A1(new_n721), .A2(new_n444), .ZN(new_n775));
  AOI21_X1  g0575(.A(new_n775), .B1(G294), .B2(new_n714), .ZN(new_n776));
  AOI22_X1  g0576(.A1(new_n711), .A2(G116), .B1(new_n727), .B2(G311), .ZN(new_n777));
  AND3_X1   g0577(.A1(new_n774), .A2(new_n776), .A3(new_n777), .ZN(new_n778));
  OAI21_X1  g0578(.A(new_n703), .B1(new_n772), .B2(new_n778), .ZN(new_n779));
  NOR2_X1   g0579(.A1(new_n703), .A2(new_n700), .ZN(new_n780));
  AOI21_X1  g0580(.A(new_n689), .B1(new_n310), .B2(new_n780), .ZN(new_n781));
  XNOR2_X1  g0581(.A(new_n781), .B(KEYINPUT93), .ZN(new_n782));
  NAND2_X1  g0582(.A1(new_n779), .A2(new_n782), .ZN(new_n783));
  XOR2_X1   g0583(.A(new_n783), .B(KEYINPUT95), .Z(new_n784));
  NAND2_X1  g0584(.A1(new_n339), .A2(new_n637), .ZN(new_n785));
  XNOR2_X1  g0585(.A(new_n785), .B(KEYINPUT96), .ZN(new_n786));
  AOI22_X1  g0586(.A1(new_n350), .A2(new_n786), .B1(new_n356), .B2(new_n355), .ZN(new_n787));
  NOR2_X1   g0587(.A1(new_n357), .A2(new_n637), .ZN(new_n788));
  NOR2_X1   g0588(.A1(new_n787), .A2(new_n788), .ZN(new_n789));
  OAI21_X1  g0589(.A(new_n784), .B1(new_n701), .B2(new_n789), .ZN(new_n790));
  XOR2_X1   g0590(.A(new_n790), .B(KEYINPUT97), .Z(new_n791));
  XNOR2_X1  g0591(.A(new_n666), .B(new_n789), .ZN(new_n792));
  OR2_X1    g0592(.A1(new_n792), .A2(new_n683), .ZN(new_n793));
  AOI21_X1  g0593(.A(new_n690), .B1(new_n792), .B2(new_n683), .ZN(new_n794));
  AND2_X1   g0594(.A1(new_n793), .A2(new_n794), .ZN(new_n795));
  NOR2_X1   g0595(.A1(new_n791), .A2(new_n795), .ZN(new_n796));
  INV_X1    g0596(.A(new_n796), .ZN(G384));
  NOR2_X1   g0597(.A1(new_n687), .A2(new_n261), .ZN(new_n798));
  INV_X1    g0598(.A(KEYINPUT102), .ZN(new_n799));
  OR2_X1    g0599(.A1(new_n332), .A2(new_n637), .ZN(new_n800));
  INV_X1    g0600(.A(KEYINPUT100), .ZN(new_n801));
  NOR2_X1   g0601(.A1(new_n391), .A2(new_n635), .ZN(new_n802));
  AND3_X1   g0602(.A1(new_n412), .A2(new_n431), .A3(KEYINPUT82), .ZN(new_n803));
  AOI21_X1  g0603(.A(KEYINPUT82), .B1(new_n412), .B2(new_n431), .ZN(new_n804));
  NOR2_X1   g0604(.A1(new_n803), .A2(new_n804), .ZN(new_n805));
  NAND2_X1  g0605(.A1(new_n440), .A2(KEYINPUT99), .ZN(new_n806));
  INV_X1    g0606(.A(KEYINPUT99), .ZN(new_n807));
  NAND3_X1  g0607(.A1(new_n437), .A2(new_n439), .A3(new_n807), .ZN(new_n808));
  NAND2_X1  g0608(.A1(new_n806), .A2(new_n808), .ZN(new_n809));
  OAI21_X1  g0609(.A(new_n802), .B1(new_n805), .B2(new_n809), .ZN(new_n810));
  OAI21_X1  g0610(.A(new_n436), .B1(new_n391), .B2(new_n411), .ZN(new_n811));
  OAI21_X1  g0611(.A(KEYINPUT37), .B1(new_n811), .B2(new_n802), .ZN(new_n812));
  NAND2_X1  g0612(.A1(new_n427), .A2(new_n430), .ZN(new_n813));
  INV_X1    g0613(.A(new_n635), .ZN(new_n814));
  NAND2_X1  g0614(.A1(new_n427), .A2(new_n814), .ZN(new_n815));
  INV_X1    g0615(.A(KEYINPUT37), .ZN(new_n816));
  NAND4_X1  g0616(.A1(new_n813), .A2(new_n815), .A3(new_n816), .A4(new_n436), .ZN(new_n817));
  NAND3_X1  g0617(.A1(new_n812), .A2(KEYINPUT98), .A3(new_n817), .ZN(new_n818));
  INV_X1    g0618(.A(KEYINPUT98), .ZN(new_n819));
  OAI211_X1 g0619(.A(new_n819), .B(KEYINPUT37), .C1(new_n811), .C2(new_n802), .ZN(new_n820));
  AND2_X1   g0620(.A1(new_n818), .A2(new_n820), .ZN(new_n821));
  AOI21_X1  g0621(.A(KEYINPUT38), .B1(new_n810), .B2(new_n821), .ZN(new_n822));
  AOI21_X1  g0622(.A(KEYINPUT16), .B1(new_n381), .B2(new_n365), .ZN(new_n823));
  OAI22_X1  g0623(.A1(new_n426), .A2(new_n823), .B1(new_n386), .B2(new_n387), .ZN(new_n824));
  NAND2_X1  g0624(.A1(new_n824), .A2(new_n430), .ZN(new_n825));
  NAND2_X1  g0625(.A1(new_n824), .A2(new_n814), .ZN(new_n826));
  NAND3_X1  g0626(.A1(new_n825), .A2(new_n826), .A3(new_n436), .ZN(new_n827));
  NAND2_X1  g0627(.A1(new_n827), .A2(KEYINPUT37), .ZN(new_n828));
  NAND2_X1  g0628(.A1(new_n828), .A2(new_n817), .ZN(new_n829));
  AOI21_X1  g0629(.A(new_n624), .B1(new_n437), .B2(new_n439), .ZN(new_n830));
  OAI211_X1 g0630(.A(KEYINPUT38), .B(new_n829), .C1(new_n830), .C2(new_n826), .ZN(new_n831));
  INV_X1    g0631(.A(KEYINPUT39), .ZN(new_n832));
  NAND2_X1  g0632(.A1(new_n831), .A2(new_n832), .ZN(new_n833));
  OAI21_X1  g0633(.A(new_n801), .B1(new_n822), .B2(new_n833), .ZN(new_n834));
  INV_X1    g0634(.A(KEYINPUT38), .ZN(new_n835));
  AND3_X1   g0635(.A1(new_n437), .A2(new_n439), .A3(new_n807), .ZN(new_n836));
  AOI21_X1  g0636(.A(new_n807), .B1(new_n437), .B2(new_n439), .ZN(new_n837));
  NOR2_X1   g0637(.A1(new_n836), .A2(new_n837), .ZN(new_n838));
  AOI21_X1  g0638(.A(new_n815), .B1(new_n628), .B2(new_n838), .ZN(new_n839));
  NAND2_X1  g0639(.A1(new_n818), .A2(new_n820), .ZN(new_n840));
  OAI21_X1  g0640(.A(new_n835), .B1(new_n839), .B2(new_n840), .ZN(new_n841));
  AND2_X1   g0641(.A1(new_n828), .A2(new_n817), .ZN(new_n842));
  AOI21_X1  g0642(.A(new_n826), .B1(new_n432), .B2(new_n440), .ZN(new_n843));
  NOR2_X1   g0643(.A1(new_n842), .A2(new_n843), .ZN(new_n844));
  AOI21_X1  g0644(.A(KEYINPUT39), .B1(new_n844), .B2(KEYINPUT38), .ZN(new_n845));
  NAND3_X1  g0645(.A1(new_n841), .A2(new_n845), .A3(KEYINPUT100), .ZN(new_n846));
  OAI21_X1  g0646(.A(new_n835), .B1(new_n842), .B2(new_n843), .ZN(new_n847));
  AOI21_X1  g0647(.A(new_n832), .B1(new_n847), .B2(new_n831), .ZN(new_n848));
  INV_X1    g0648(.A(new_n848), .ZN(new_n849));
  NAND3_X1  g0649(.A1(new_n834), .A2(new_n846), .A3(new_n849), .ZN(new_n850));
  NAND2_X1  g0650(.A1(new_n850), .A2(KEYINPUT101), .ZN(new_n851));
  INV_X1    g0651(.A(KEYINPUT101), .ZN(new_n852));
  NAND4_X1  g0652(.A1(new_n834), .A2(new_n846), .A3(new_n852), .A4(new_n849), .ZN(new_n853));
  AOI21_X1  g0653(.A(new_n800), .B1(new_n851), .B2(new_n853), .ZN(new_n854));
  AOI21_X1  g0654(.A(new_n788), .B1(new_n666), .B2(new_n789), .ZN(new_n855));
  NOR2_X1   g0655(.A1(new_n319), .A2(new_n643), .ZN(new_n856));
  INV_X1    g0656(.A(new_n856), .ZN(new_n857));
  NAND3_X1  g0657(.A1(new_n332), .A2(new_n353), .A3(new_n857), .ZN(new_n858));
  OAI21_X1  g0658(.A(new_n856), .B1(new_n330), .B2(new_n331), .ZN(new_n859));
  NAND2_X1  g0659(.A1(new_n858), .A2(new_n859), .ZN(new_n860));
  INV_X1    g0660(.A(new_n860), .ZN(new_n861));
  NOR2_X1   g0661(.A1(new_n855), .A2(new_n861), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n847), .A2(new_n831), .ZN(new_n863));
  NAND2_X1  g0663(.A1(new_n862), .A2(new_n863), .ZN(new_n864));
  NOR2_X1   g0664(.A1(new_n628), .A2(new_n814), .ZN(new_n865));
  INV_X1    g0665(.A(new_n865), .ZN(new_n866));
  NAND2_X1  g0666(.A1(new_n864), .A2(new_n866), .ZN(new_n867));
  OAI21_X1  g0667(.A(new_n799), .B1(new_n854), .B2(new_n867), .ZN(new_n868));
  INV_X1    g0668(.A(new_n800), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n841), .A2(new_n845), .ZN(new_n870));
  AOI21_X1  g0670(.A(new_n848), .B1(new_n870), .B2(new_n801), .ZN(new_n871));
  AOI21_X1  g0671(.A(new_n852), .B1(new_n871), .B2(new_n846), .ZN(new_n872));
  AND4_X1   g0672(.A1(new_n852), .A2(new_n834), .A3(new_n846), .A4(new_n849), .ZN(new_n873));
  OAI21_X1  g0673(.A(new_n869), .B1(new_n872), .B2(new_n873), .ZN(new_n874));
  AOI21_X1  g0674(.A(new_n865), .B1(new_n862), .B2(new_n863), .ZN(new_n875));
  NAND3_X1  g0675(.A1(new_n874), .A2(KEYINPUT102), .A3(new_n875), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n868), .A2(new_n876), .ZN(new_n877));
  OAI211_X1 g0677(.A(new_n442), .B(new_n665), .C1(new_n666), .C2(KEYINPUT29), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n878), .A2(new_n630), .ZN(new_n879));
  XOR2_X1   g0679(.A(new_n877), .B(new_n879), .Z(new_n880));
  NAND2_X1  g0680(.A1(new_n678), .A2(KEYINPUT103), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n668), .A2(new_n881), .ZN(new_n882));
  INV_X1    g0682(.A(new_n882), .ZN(new_n883));
  AOI21_X1  g0683(.A(new_n678), .B1(KEYINPUT103), .B2(new_n681), .ZN(new_n884));
  INV_X1    g0684(.A(new_n884), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n883), .A2(new_n885), .ZN(new_n886));
  INV_X1    g0686(.A(new_n787), .ZN(new_n887));
  INV_X1    g0687(.A(new_n788), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n887), .A2(new_n888), .ZN(new_n889));
  NOR2_X1   g0689(.A1(new_n889), .A2(new_n861), .ZN(new_n890));
  AND2_X1   g0690(.A1(new_n886), .A2(new_n890), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n891), .A2(KEYINPUT40), .ZN(new_n892));
  AND2_X1   g0692(.A1(new_n841), .A2(new_n831), .ZN(new_n893));
  NOR2_X1   g0693(.A1(new_n892), .A2(new_n893), .ZN(new_n894));
  AOI21_X1  g0694(.A(KEYINPUT40), .B1(new_n891), .B2(new_n863), .ZN(new_n895));
  NOR2_X1   g0695(.A1(new_n894), .A2(new_n895), .ZN(new_n896));
  INV_X1    g0696(.A(new_n896), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n886), .A2(new_n442), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n897), .A2(new_n898), .ZN(new_n899));
  NAND3_X1  g0699(.A1(new_n896), .A2(new_n442), .A3(new_n886), .ZN(new_n900));
  NAND3_X1  g0700(.A1(new_n899), .A2(G330), .A3(new_n900), .ZN(new_n901));
  AOI21_X1  g0701(.A(new_n798), .B1(new_n880), .B2(new_n901), .ZN(new_n902));
  OAI21_X1  g0702(.A(new_n902), .B1(new_n880), .B2(new_n901), .ZN(new_n903));
  OR2_X1    g0703(.A1(new_n560), .A2(KEYINPUT35), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n560), .A2(KEYINPUT35), .ZN(new_n905));
  NAND4_X1  g0705(.A1(new_n904), .A2(G116), .A3(new_n216), .A4(new_n905), .ZN(new_n906));
  XNOR2_X1  g0706(.A(new_n906), .B(KEYINPUT36), .ZN(new_n907));
  NAND4_X1  g0707(.A1(new_n213), .A2(G77), .A3(new_n363), .A4(new_n361), .ZN(new_n908));
  OAI21_X1  g0708(.A(new_n908), .B1(G50), .B2(new_n203), .ZN(new_n909));
  NAND3_X1  g0709(.A1(new_n909), .A2(G1), .A3(new_n287), .ZN(new_n910));
  NAND3_X1  g0710(.A1(new_n903), .A2(new_n907), .A3(new_n910), .ZN(G367));
  NAND2_X1  g0711(.A1(new_n688), .A2(G1), .ZN(new_n912));
  INV_X1    g0712(.A(new_n912), .ZN(new_n913));
  XNOR2_X1  g0713(.A(new_n648), .B(new_n652), .ZN(new_n914));
  XNOR2_X1  g0714(.A(new_n914), .B(new_n642), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n915), .A2(new_n685), .ZN(new_n916));
  NOR2_X1   g0716(.A1(new_n590), .A2(new_n643), .ZN(new_n917));
  OR2_X1    g0717(.A1(new_n592), .A2(new_n917), .ZN(new_n918));
  NAND3_X1  g0718(.A1(new_n917), .A2(new_n580), .A3(new_n585), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n918), .A2(new_n919), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n653), .A2(new_n920), .ZN(new_n921));
  XOR2_X1   g0721(.A(new_n921), .B(KEYINPUT45), .Z(new_n922));
  NOR2_X1   g0722(.A1(new_n653), .A2(new_n920), .ZN(new_n923));
  XNOR2_X1  g0723(.A(new_n923), .B(KEYINPUT44), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n922), .A2(new_n924), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n925), .A2(new_n651), .ZN(new_n926));
  NAND3_X1  g0726(.A1(new_n922), .A2(new_n650), .A3(new_n924), .ZN(new_n927));
  AOI21_X1  g0727(.A(new_n916), .B1(new_n926), .B2(new_n927), .ZN(new_n928));
  NOR2_X1   g0728(.A1(new_n928), .A2(new_n684), .ZN(new_n929));
  XOR2_X1   g0729(.A(new_n656), .B(KEYINPUT41), .Z(new_n930));
  OAI21_X1  g0730(.A(new_n913), .B1(new_n929), .B2(new_n930), .ZN(new_n931));
  NAND3_X1  g0731(.A1(new_n648), .A2(new_n652), .A3(new_n920), .ZN(new_n932));
  OR2_X1    g0732(.A1(new_n932), .A2(KEYINPUT42), .ZN(new_n933));
  INV_X1    g0733(.A(new_n920), .ZN(new_n934));
  OAI21_X1  g0734(.A(new_n587), .B1(new_n934), .B2(new_n645), .ZN(new_n935));
  AOI22_X1  g0735(.A1(new_n932), .A2(KEYINPUT42), .B1(new_n643), .B2(new_n935), .ZN(new_n936));
  AOI21_X1  g0736(.A(new_n643), .B1(new_n452), .B2(new_n470), .ZN(new_n937));
  NAND4_X1  g0737(.A1(new_n479), .A2(new_n477), .A3(new_n595), .A4(new_n937), .ZN(new_n938));
  OAI21_X1  g0738(.A(new_n938), .B1(new_n607), .B2(new_n937), .ZN(new_n939));
  AOI22_X1  g0739(.A1(new_n933), .A2(new_n936), .B1(KEYINPUT43), .B2(new_n939), .ZN(new_n940));
  OR2_X1    g0740(.A1(new_n939), .A2(KEYINPUT43), .ZN(new_n941));
  XNOR2_X1  g0741(.A(new_n940), .B(new_n941), .ZN(new_n942));
  NOR2_X1   g0742(.A1(new_n651), .A2(new_n934), .ZN(new_n943));
  XNOR2_X1  g0743(.A(new_n942), .B(new_n943), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n931), .A2(new_n944), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n694), .A2(new_n235), .ZN(new_n946));
  INV_X1    g0746(.A(new_n704), .ZN(new_n947));
  AOI21_X1  g0747(.A(new_n947), .B1(new_n655), .B2(new_n475), .ZN(new_n948));
  AOI21_X1  g0748(.A(new_n689), .B1(new_n946), .B2(new_n948), .ZN(new_n949));
  NAND2_X1  g0749(.A1(new_n745), .A2(G68), .ZN(new_n950));
  INV_X1    g0750(.A(G150), .ZN(new_n951));
  OAI21_X1  g0751(.A(new_n950), .B1(new_n951), .B2(new_n713), .ZN(new_n952));
  XNOR2_X1  g0752(.A(new_n952), .B(KEYINPUT105), .ZN(new_n953));
  INV_X1    g0753(.A(new_n731), .ZN(new_n954));
  AOI21_X1  g0754(.A(new_n248), .B1(new_n954), .B2(G58), .ZN(new_n955));
  INV_X1    g0755(.A(new_n737), .ZN(new_n956));
  OAI221_X1 g0756(.A(new_n955), .B1(new_n956), .B2(new_n415), .C1(new_n763), .C2(new_n734), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n722), .A2(G77), .ZN(new_n958));
  INV_X1    g0758(.A(G137), .ZN(new_n959));
  OAI221_X1 g0759(.A(new_n958), .B1(new_n959), .B2(new_n726), .C1(new_n710), .C2(new_n201), .ZN(new_n960));
  NOR3_X1   g0760(.A1(new_n953), .A2(new_n957), .A3(new_n960), .ZN(new_n961));
  OAI221_X1 g0761(.A(new_n379), .B1(new_n726), .B2(new_n738), .C1(new_n721), .C2(new_n445), .ZN(new_n962));
  INV_X1    g0762(.A(KEYINPUT104), .ZN(new_n963));
  NAND2_X1  g0763(.A1(new_n962), .A2(new_n963), .ZN(new_n964));
  NOR2_X1   g0764(.A1(new_n962), .A2(new_n963), .ZN(new_n965));
  NAND2_X1  g0765(.A1(new_n737), .A2(G294), .ZN(new_n966));
  NOR2_X1   g0766(.A1(new_n731), .A2(new_n456), .ZN(new_n967));
  OAI221_X1 g0767(.A(new_n966), .B1(KEYINPUT46), .B2(new_n967), .C1(new_n446), .C2(new_n742), .ZN(new_n968));
  AOI22_X1  g0768(.A1(new_n967), .A2(KEYINPUT46), .B1(new_n733), .B2(G311), .ZN(new_n969));
  INV_X1    g0769(.A(G283), .ZN(new_n970));
  OAI221_X1 g0770(.A(new_n969), .B1(new_n713), .B2(new_n540), .C1(new_n970), .C2(new_n710), .ZN(new_n971));
  NOR3_X1   g0771(.A1(new_n965), .A2(new_n968), .A3(new_n971), .ZN(new_n972));
  AOI21_X1  g0772(.A(new_n961), .B1(new_n964), .B2(new_n972), .ZN(new_n973));
  XNOR2_X1  g0773(.A(new_n973), .B(KEYINPUT47), .ZN(new_n974));
  OAI221_X1 g0774(.A(new_n949), .B1(new_n759), .B2(new_n939), .C1(new_n974), .C2(new_n706), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n945), .A2(new_n975), .ZN(G387));
  OR2_X1    g0776(.A1(new_n648), .A2(new_n759), .ZN(new_n977));
  OAI22_X1  g0777(.A1(new_n698), .A2(new_n658), .B1(G107), .B2(new_n208), .ZN(new_n978));
  XNOR2_X1  g0778(.A(KEYINPUT106), .B(KEYINPUT50), .ZN(new_n979));
  OR3_X1    g0779(.A1(new_n274), .A2(new_n979), .A3(G50), .ZN(new_n980));
  OAI21_X1  g0780(.A(new_n979), .B1(new_n274), .B2(G50), .ZN(new_n981));
  AOI21_X1  g0781(.A(G45), .B1(G68), .B2(G77), .ZN(new_n982));
  NAND4_X1  g0782(.A1(new_n980), .A2(new_n658), .A3(new_n981), .A4(new_n982), .ZN(new_n983));
  AND2_X1   g0783(.A1(new_n694), .A2(new_n983), .ZN(new_n984));
  NAND2_X1  g0784(.A1(new_n232), .A2(G45), .ZN(new_n985));
  AOI21_X1  g0785(.A(new_n978), .B1(new_n984), .B2(new_n985), .ZN(new_n986));
  OAI21_X1  g0786(.A(new_n690), .B1(new_n986), .B2(new_n947), .ZN(new_n987));
  XOR2_X1   g0787(.A(KEYINPUT107), .B(G322), .Z(new_n988));
  AOI22_X1  g0788(.A1(G311), .A2(new_n737), .B1(new_n733), .B2(new_n988), .ZN(new_n989));
  OAI221_X1 g0789(.A(new_n989), .B1(new_n713), .B2(new_n738), .C1(new_n540), .C2(new_n710), .ZN(new_n990));
  INV_X1    g0790(.A(KEYINPUT48), .ZN(new_n991));
  OR2_X1    g0791(.A1(new_n990), .A2(new_n991), .ZN(new_n992));
  OAI22_X1  g0792(.A1(new_n742), .A2(new_n970), .B1(new_n731), .B2(new_n504), .ZN(new_n993));
  AOI21_X1  g0793(.A(new_n993), .B1(new_n990), .B2(new_n991), .ZN(new_n994));
  NAND3_X1  g0794(.A1(new_n992), .A2(KEYINPUT49), .A3(new_n994), .ZN(new_n995));
  OAI221_X1 g0795(.A(new_n379), .B1(new_n726), .B2(new_n735), .C1(new_n721), .C2(new_n456), .ZN(new_n996));
  XOR2_X1   g0796(.A(new_n996), .B(KEYINPUT108), .Z(new_n997));
  NAND2_X1  g0797(.A1(new_n995), .A2(new_n997), .ZN(new_n998));
  AOI21_X1  g0798(.A(KEYINPUT49), .B1(new_n992), .B2(new_n994), .ZN(new_n999));
  AOI22_X1  g0799(.A1(G50), .A2(new_n714), .B1(new_n711), .B2(G68), .ZN(new_n1000));
  OAI21_X1  g0800(.A(new_n1000), .B1(new_n278), .B2(new_n956), .ZN(new_n1001));
  AOI22_X1  g0801(.A1(new_n722), .A2(G97), .B1(new_n727), .B2(G150), .ZN(new_n1002));
  NAND2_X1  g0802(.A1(new_n745), .A2(new_n475), .ZN(new_n1003));
  NOR2_X1   g0803(.A1(new_n731), .A2(new_n310), .ZN(new_n1004));
  AOI211_X1 g0804(.A(new_n379), .B(new_n1004), .C1(G159), .C2(new_n733), .ZN(new_n1005));
  NAND3_X1  g0805(.A1(new_n1002), .A2(new_n1003), .A3(new_n1005), .ZN(new_n1006));
  OAI22_X1  g0806(.A1(new_n998), .A2(new_n999), .B1(new_n1001), .B2(new_n1006), .ZN(new_n1007));
  AOI21_X1  g0807(.A(new_n987), .B1(new_n1007), .B2(new_n703), .ZN(new_n1008));
  AOI22_X1  g0808(.A1(new_n915), .A2(new_n912), .B1(new_n977), .B2(new_n1008), .ZN(new_n1009));
  NAND2_X1  g0809(.A1(new_n916), .A2(new_n656), .ZN(new_n1010));
  NOR2_X1   g0810(.A1(new_n915), .A2(new_n685), .ZN(new_n1011));
  OAI21_X1  g0811(.A(new_n1009), .B1(new_n1010), .B2(new_n1011), .ZN(G393));
  NOR2_X1   g0812(.A1(new_n928), .A2(new_n657), .ZN(new_n1013));
  INV_X1    g0813(.A(new_n916), .ZN(new_n1014));
  NAND2_X1  g0814(.A1(new_n926), .A2(new_n927), .ZN(new_n1015));
  OAI21_X1  g0815(.A(new_n1013), .B1(new_n1014), .B2(new_n1015), .ZN(new_n1016));
  NAND2_X1  g0816(.A1(new_n934), .A2(new_n702), .ZN(new_n1017));
  AOI22_X1  g0817(.A1(new_n714), .A2(G311), .B1(G317), .B2(new_n733), .ZN(new_n1018));
  XOR2_X1   g0818(.A(new_n1018), .B(KEYINPUT52), .Z(new_n1019));
  NOR2_X1   g0819(.A1(new_n742), .A2(new_n456), .ZN(new_n1020));
  OAI21_X1  g0820(.A(new_n248), .B1(new_n731), .B2(new_n970), .ZN(new_n1021));
  AOI211_X1 g0821(.A(new_n1020), .B(new_n1021), .C1(new_n541), .C2(new_n737), .ZN(new_n1022));
  NAND2_X1  g0822(.A1(new_n711), .A2(G294), .ZN(new_n1023));
  AOI21_X1  g0823(.A(new_n754), .B1(new_n727), .B2(new_n988), .ZN(new_n1024));
  NAND4_X1  g0824(.A1(new_n1019), .A2(new_n1022), .A3(new_n1023), .A4(new_n1024), .ZN(new_n1025));
  NOR2_X1   g0825(.A1(new_n710), .A2(new_n274), .ZN(new_n1026));
  AOI211_X1 g0826(.A(new_n1026), .B(new_n775), .C1(G143), .C2(new_n727), .ZN(new_n1027));
  OAI22_X1  g0827(.A1(new_n713), .A2(new_n415), .B1(new_n951), .B2(new_n734), .ZN(new_n1028));
  XNOR2_X1  g0828(.A(new_n1028), .B(KEYINPUT51), .ZN(new_n1029));
  OAI221_X1 g0829(.A(new_n377), .B1(new_n203), .B2(new_n731), .C1(new_n956), .C2(new_n201), .ZN(new_n1030));
  AOI21_X1  g0830(.A(new_n1030), .B1(G77), .B2(new_n745), .ZN(new_n1031));
  NAND3_X1  g0831(.A1(new_n1027), .A2(new_n1029), .A3(new_n1031), .ZN(new_n1032));
  AOI21_X1  g0832(.A(new_n706), .B1(new_n1025), .B2(new_n1032), .ZN(new_n1033));
  INV_X1    g0833(.A(new_n694), .ZN(new_n1034));
  OR2_X1    g0834(.A1(new_n1034), .A2(new_n242), .ZN(new_n1035));
  AOI21_X1  g0835(.A(new_n947), .B1(G97), .B2(new_n655), .ZN(new_n1036));
  AOI211_X1 g0836(.A(new_n689), .B(new_n1033), .C1(new_n1035), .C2(new_n1036), .ZN(new_n1037));
  AOI22_X1  g0837(.A1(new_n1015), .A2(new_n912), .B1(new_n1017), .B2(new_n1037), .ZN(new_n1038));
  NAND2_X1  g0838(.A1(new_n1016), .A2(new_n1038), .ZN(G390));
  NAND3_X1  g0839(.A1(new_n851), .A2(new_n700), .A3(new_n853), .ZN(new_n1040));
  AOI21_X1  g0840(.A(new_n689), .B1(new_n278), .B2(new_n780), .ZN(new_n1041));
  XOR2_X1   g0841(.A(new_n1041), .B(KEYINPUT114), .Z(new_n1042));
  AOI22_X1  g0842(.A1(new_n714), .A2(G116), .B1(new_n727), .B2(G294), .ZN(new_n1043));
  OAI221_X1 g0843(.A(new_n1043), .B1(new_n203), .B2(new_n721), .C1(new_n445), .C2(new_n710), .ZN(new_n1044));
  AOI211_X1 g0844(.A(new_n250), .B(new_n755), .C1(G107), .C2(new_n737), .ZN(new_n1045));
  OAI221_X1 g0845(.A(new_n1045), .B1(new_n970), .B2(new_n734), .C1(new_n746), .C2(new_n310), .ZN(new_n1046));
  INV_X1    g0846(.A(G128), .ZN(new_n1047));
  INV_X1    g0847(.A(KEYINPUT53), .ZN(new_n1048));
  NOR2_X1   g0848(.A1(new_n731), .A2(new_n951), .ZN(new_n1049));
  OAI22_X1  g0849(.A1(new_n734), .A2(new_n1047), .B1(new_n1048), .B2(new_n1049), .ZN(new_n1050));
  AOI21_X1  g0850(.A(new_n1050), .B1(new_n1048), .B2(new_n1049), .ZN(new_n1051));
  OAI21_X1  g0851(.A(new_n250), .B1(new_n956), .B2(new_n959), .ZN(new_n1052));
  XNOR2_X1  g0852(.A(KEYINPUT54), .B(G143), .ZN(new_n1053));
  INV_X1    g0853(.A(new_n1053), .ZN(new_n1054));
  AOI21_X1  g0854(.A(new_n1052), .B1(new_n711), .B2(new_n1054), .ZN(new_n1055));
  OAI211_X1 g0855(.A(new_n1051), .B(new_n1055), .C1(new_n415), .C2(new_n746), .ZN(new_n1056));
  AOI22_X1  g0856(.A1(new_n722), .A2(G50), .B1(new_n727), .B2(G125), .ZN(new_n1057));
  OAI21_X1  g0857(.A(new_n1057), .B1(new_n770), .B2(new_n713), .ZN(new_n1058));
  OAI22_X1  g0858(.A1(new_n1044), .A2(new_n1046), .B1(new_n1056), .B2(new_n1058), .ZN(new_n1059));
  AOI21_X1  g0859(.A(new_n1042), .B1(new_n1059), .B2(new_n703), .ZN(new_n1060));
  NAND2_X1  g0860(.A1(new_n1040), .A2(new_n1060), .ZN(new_n1061));
  XOR2_X1   g0861(.A(new_n1061), .B(KEYINPUT115), .Z(new_n1062));
  OAI21_X1  g0862(.A(new_n800), .B1(new_n855), .B2(new_n861), .ZN(new_n1063));
  NAND3_X1  g0863(.A1(new_n851), .A2(new_n853), .A3(new_n1063), .ZN(new_n1064));
  NOR2_X1   g0864(.A1(new_n893), .A2(new_n869), .ZN(new_n1065));
  OAI211_X1 g0865(.A(new_n643), .B(new_n887), .C1(new_n664), .C2(new_n605), .ZN(new_n1066));
  NAND2_X1  g0866(.A1(new_n1066), .A2(new_n888), .ZN(new_n1067));
  INV_X1    g0867(.A(KEYINPUT109), .ZN(new_n1068));
  NAND2_X1  g0868(.A1(new_n1067), .A2(new_n1068), .ZN(new_n1069));
  NAND3_X1  g0869(.A1(new_n1066), .A2(KEYINPUT109), .A3(new_n888), .ZN(new_n1070));
  NAND2_X1  g0870(.A1(new_n1069), .A2(new_n1070), .ZN(new_n1071));
  OAI21_X1  g0871(.A(new_n1065), .B1(new_n1071), .B2(new_n861), .ZN(new_n1072));
  NAND2_X1  g0872(.A1(new_n681), .A2(KEYINPUT86), .ZN(new_n1073));
  INV_X1    g0873(.A(new_n678), .ZN(new_n1074));
  NAND2_X1  g0874(.A1(new_n1073), .A2(new_n1074), .ZN(new_n1075));
  NAND3_X1  g0875(.A1(new_n1075), .A2(new_n668), .A3(new_n679), .ZN(new_n1076));
  NAND3_X1  g0876(.A1(new_n1076), .A2(G330), .A3(new_n789), .ZN(new_n1077));
  NOR2_X1   g0877(.A1(new_n1077), .A2(new_n861), .ZN(new_n1078));
  NAND3_X1  g0878(.A1(new_n886), .A2(new_n890), .A3(G330), .ZN(new_n1079));
  OAI21_X1  g0879(.A(new_n1078), .B1(new_n1079), .B2(KEYINPUT110), .ZN(new_n1080));
  AND3_X1   g0880(.A1(new_n1064), .A2(new_n1072), .A3(new_n1080), .ZN(new_n1081));
  INV_X1    g0881(.A(G330), .ZN(new_n1082));
  AOI21_X1  g0882(.A(new_n1082), .B1(new_n883), .B2(new_n885), .ZN(new_n1083));
  NAND3_X1  g0883(.A1(new_n1083), .A2(KEYINPUT110), .A3(new_n890), .ZN(new_n1084));
  AOI21_X1  g0884(.A(new_n1084), .B1(new_n1064), .B2(new_n1072), .ZN(new_n1085));
  NOR2_X1   g0885(.A1(new_n1081), .A2(new_n1085), .ZN(new_n1086));
  AOI21_X1  g0886(.A(new_n1062), .B1(new_n912), .B2(new_n1086), .ZN(new_n1087));
  INV_X1    g0887(.A(new_n1086), .ZN(new_n1088));
  NAND3_X1  g0888(.A1(new_n886), .A2(G330), .A3(new_n442), .ZN(new_n1089));
  NAND3_X1  g0889(.A1(new_n1089), .A2(new_n878), .A3(new_n630), .ZN(new_n1090));
  NAND2_X1  g0890(.A1(new_n1090), .A2(KEYINPUT111), .ZN(new_n1091));
  INV_X1    g0891(.A(KEYINPUT111), .ZN(new_n1092));
  NAND4_X1  g0892(.A1(new_n1089), .A2(new_n878), .A3(new_n1092), .A4(new_n630), .ZN(new_n1093));
  NAND2_X1  g0893(.A1(new_n1091), .A2(new_n1093), .ZN(new_n1094));
  OAI211_X1 g0894(.A(G330), .B(new_n789), .C1(new_n882), .C2(new_n884), .ZN(new_n1095));
  NAND2_X1  g0895(.A1(new_n1095), .A2(new_n861), .ZN(new_n1096));
  NAND4_X1  g0896(.A1(new_n1076), .A2(G330), .A3(new_n789), .A4(new_n860), .ZN(new_n1097));
  AND2_X1   g0897(.A1(new_n1096), .A2(new_n1097), .ZN(new_n1098));
  OAI21_X1  g0898(.A(new_n861), .B1(new_n683), .B2(new_n889), .ZN(new_n1099));
  NAND2_X1  g0899(.A1(new_n1079), .A2(new_n1099), .ZN(new_n1100));
  INV_X1    g0900(.A(new_n855), .ZN(new_n1101));
  AOI22_X1  g0901(.A1(new_n1071), .A2(new_n1098), .B1(new_n1100), .B2(new_n1101), .ZN(new_n1102));
  NOR2_X1   g0902(.A1(new_n1094), .A2(new_n1102), .ZN(new_n1103));
  INV_X1    g0903(.A(new_n1103), .ZN(new_n1104));
  NAND2_X1  g0904(.A1(new_n1088), .A2(new_n1104), .ZN(new_n1105));
  NAND2_X1  g0905(.A1(new_n1064), .A2(new_n1072), .ZN(new_n1106));
  INV_X1    g0906(.A(new_n1084), .ZN(new_n1107));
  NAND2_X1  g0907(.A1(new_n1106), .A2(new_n1107), .ZN(new_n1108));
  NAND3_X1  g0908(.A1(new_n1064), .A2(new_n1072), .A3(new_n1080), .ZN(new_n1109));
  NAND3_X1  g0909(.A1(new_n1108), .A2(new_n1103), .A3(new_n1109), .ZN(new_n1110));
  NAND2_X1  g0910(.A1(new_n1110), .A2(KEYINPUT112), .ZN(new_n1111));
  INV_X1    g0911(.A(KEYINPUT112), .ZN(new_n1112));
  NAND4_X1  g0912(.A1(new_n1108), .A2(new_n1103), .A3(new_n1112), .A4(new_n1109), .ZN(new_n1113));
  AOI21_X1  g0913(.A(new_n657), .B1(new_n1111), .B2(new_n1113), .ZN(new_n1114));
  INV_X1    g0914(.A(KEYINPUT113), .ZN(new_n1115));
  OAI21_X1  g0915(.A(new_n1105), .B1(new_n1114), .B2(new_n1115), .ZN(new_n1116));
  AOI211_X1 g0916(.A(KEYINPUT113), .B(new_n657), .C1(new_n1111), .C2(new_n1113), .ZN(new_n1117));
  OAI21_X1  g0917(.A(new_n1087), .B1(new_n1116), .B2(new_n1117), .ZN(G378));
  INV_X1    g0918(.A(KEYINPUT57), .ZN(new_n1119));
  NOR2_X1   g0919(.A1(new_n897), .A2(new_n1082), .ZN(new_n1120));
  INV_X1    g0920(.A(new_n1120), .ZN(new_n1121));
  XNOR2_X1  g0921(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1122));
  XOR2_X1   g0922(.A(new_n308), .B(new_n1122), .Z(new_n1123));
  NAND2_X1  g0923(.A1(new_n293), .A2(new_n814), .ZN(new_n1124));
  XNOR2_X1  g0924(.A(new_n1123), .B(new_n1124), .ZN(new_n1125));
  INV_X1    g0925(.A(KEYINPUT117), .ZN(new_n1126));
  NAND2_X1  g0926(.A1(new_n1125), .A2(new_n1126), .ZN(new_n1127));
  AND3_X1   g0927(.A1(new_n868), .A2(new_n876), .A3(new_n1127), .ZN(new_n1128));
  AOI21_X1  g0928(.A(new_n1127), .B1(new_n868), .B2(new_n876), .ZN(new_n1129));
  OAI21_X1  g0929(.A(new_n1121), .B1(new_n1128), .B2(new_n1129), .ZN(new_n1130));
  INV_X1    g0930(.A(new_n1127), .ZN(new_n1131));
  NOR3_X1   g0931(.A1(new_n854), .A2(new_n867), .A3(new_n799), .ZN(new_n1132));
  AOI21_X1  g0932(.A(KEYINPUT102), .B1(new_n874), .B2(new_n875), .ZN(new_n1133));
  OAI21_X1  g0933(.A(new_n1131), .B1(new_n1132), .B2(new_n1133), .ZN(new_n1134));
  NAND3_X1  g0934(.A1(new_n868), .A2(new_n876), .A3(new_n1127), .ZN(new_n1135));
  NAND3_X1  g0935(.A1(new_n1134), .A2(new_n1120), .A3(new_n1135), .ZN(new_n1136));
  NAND2_X1  g0936(.A1(new_n1130), .A2(new_n1136), .ZN(new_n1137));
  AOI21_X1  g0937(.A(new_n1094), .B1(new_n1111), .B2(new_n1113), .ZN(new_n1138));
  OAI21_X1  g0938(.A(new_n1119), .B1(new_n1137), .B2(new_n1138), .ZN(new_n1139));
  INV_X1    g0939(.A(new_n1094), .ZN(new_n1140));
  AOI21_X1  g0940(.A(new_n1112), .B1(new_n1086), .B2(new_n1103), .ZN(new_n1141));
  INV_X1    g0941(.A(new_n1113), .ZN(new_n1142));
  OAI21_X1  g0942(.A(new_n1140), .B1(new_n1141), .B2(new_n1142), .ZN(new_n1143));
  NAND4_X1  g0943(.A1(new_n1143), .A2(KEYINPUT57), .A3(new_n1136), .A4(new_n1130), .ZN(new_n1144));
  NAND3_X1  g0944(.A1(new_n1139), .A2(new_n1144), .A3(new_n656), .ZN(new_n1145));
  NAND3_X1  g0945(.A1(new_n1130), .A2(new_n1136), .A3(new_n912), .ZN(new_n1146));
  INV_X1    g0946(.A(new_n780), .ZN(new_n1147));
  OAI21_X1  g0947(.A(new_n690), .B1(G50), .B2(new_n1147), .ZN(new_n1148));
  NOR2_X1   g0948(.A1(new_n710), .A2(new_n336), .ZN(new_n1149));
  NOR2_X1   g0949(.A1(new_n721), .A2(new_n202), .ZN(new_n1150));
  AOI211_X1 g0950(.A(new_n1149), .B(new_n1150), .C1(G283), .C2(new_n727), .ZN(new_n1151));
  NAND2_X1  g0951(.A1(new_n714), .A2(G107), .ZN(new_n1152));
  XNOR2_X1  g0952(.A(new_n1152), .B(KEYINPUT116), .ZN(new_n1153));
  OAI22_X1  g0953(.A1(new_n956), .A2(new_n445), .B1(new_n734), .B2(new_n456), .ZN(new_n1154));
  NOR4_X1   g0954(.A1(new_n1154), .A2(new_n1004), .A3(G41), .A4(new_n377), .ZN(new_n1155));
  NAND4_X1  g0955(.A1(new_n1151), .A2(new_n1153), .A3(new_n950), .A4(new_n1155), .ZN(new_n1156));
  INV_X1    g0956(.A(KEYINPUT58), .ZN(new_n1157));
  OAI21_X1  g0957(.A(new_n509), .B1(new_n379), .B2(new_n244), .ZN(new_n1158));
  AOI22_X1  g0958(.A1(new_n1156), .A2(new_n1157), .B1(new_n201), .B2(new_n1158), .ZN(new_n1159));
  AOI22_X1  g0959(.A1(G128), .A2(new_n714), .B1(new_n711), .B2(G137), .ZN(new_n1160));
  NAND2_X1  g0960(.A1(new_n745), .A2(G150), .ZN(new_n1161));
  NAND2_X1  g0961(.A1(new_n733), .A2(G125), .ZN(new_n1162));
  AOI22_X1  g0962(.A1(new_n737), .A2(G132), .B1(new_n954), .B2(new_n1054), .ZN(new_n1163));
  NAND4_X1  g0963(.A1(new_n1160), .A2(new_n1161), .A3(new_n1162), .A4(new_n1163), .ZN(new_n1164));
  NOR2_X1   g0964(.A1(new_n1164), .A2(KEYINPUT59), .ZN(new_n1165));
  NAND2_X1  g0965(.A1(new_n1164), .A2(KEYINPUT59), .ZN(new_n1166));
  OAI211_X1 g0966(.A(new_n244), .B(new_n509), .C1(new_n721), .C2(new_n415), .ZN(new_n1167));
  AOI21_X1  g0967(.A(new_n1167), .B1(G124), .B2(new_n727), .ZN(new_n1168));
  NAND2_X1  g0968(.A1(new_n1166), .A2(new_n1168), .ZN(new_n1169));
  OAI221_X1 g0969(.A(new_n1159), .B1(new_n1157), .B2(new_n1156), .C1(new_n1165), .C2(new_n1169), .ZN(new_n1170));
  AOI21_X1  g0970(.A(new_n1148), .B1(new_n1170), .B2(new_n703), .ZN(new_n1171));
  INV_X1    g0971(.A(new_n1125), .ZN(new_n1172));
  OAI21_X1  g0972(.A(new_n1171), .B1(new_n1172), .B2(new_n701), .ZN(new_n1173));
  NAND2_X1  g0973(.A1(new_n1146), .A2(new_n1173), .ZN(new_n1174));
  INV_X1    g0974(.A(new_n1174), .ZN(new_n1175));
  NAND2_X1  g0975(.A1(new_n1145), .A2(new_n1175), .ZN(G375));
  OAI21_X1  g0976(.A(new_n690), .B1(G68), .B2(new_n1147), .ZN(new_n1177));
  AOI21_X1  g0977(.A(new_n1150), .B1(G137), .B2(new_n714), .ZN(new_n1178));
  OAI221_X1 g0978(.A(new_n1178), .B1(new_n1047), .B2(new_n726), .C1(new_n951), .C2(new_n710), .ZN(new_n1179));
  AOI21_X1  g0979(.A(new_n379), .B1(new_n954), .B2(G159), .ZN(new_n1180));
  AOI22_X1  g0980(.A1(G132), .A2(new_n733), .B1(new_n737), .B2(new_n1054), .ZN(new_n1181));
  OAI211_X1 g0981(.A(new_n1180), .B(new_n1181), .C1(new_n746), .C2(new_n201), .ZN(new_n1182));
  AOI22_X1  g0982(.A1(new_n714), .A2(G283), .B1(new_n727), .B2(G303), .ZN(new_n1183));
  OAI211_X1 g0983(.A(new_n1183), .B(new_n958), .C1(new_n446), .C2(new_n710), .ZN(new_n1184));
  OAI21_X1  g0984(.A(new_n248), .B1(new_n731), .B2(new_n445), .ZN(new_n1185));
  AOI21_X1  g0985(.A(new_n1185), .B1(G116), .B2(new_n737), .ZN(new_n1186));
  OAI211_X1 g0986(.A(new_n1003), .B(new_n1186), .C1(new_n504), .C2(new_n734), .ZN(new_n1187));
  OAI22_X1  g0987(.A1(new_n1179), .A2(new_n1182), .B1(new_n1184), .B2(new_n1187), .ZN(new_n1188));
  AOI21_X1  g0988(.A(new_n1177), .B1(new_n1188), .B2(new_n703), .ZN(new_n1189));
  OAI21_X1  g0989(.A(new_n1189), .B1(new_n860), .B2(new_n701), .ZN(new_n1190));
  NOR2_X1   g0990(.A1(new_n1102), .A2(new_n913), .ZN(new_n1191));
  OAI21_X1  g0991(.A(new_n1190), .B1(new_n1191), .B2(KEYINPUT119), .ZN(new_n1192));
  AOI21_X1  g0992(.A(new_n1192), .B1(KEYINPUT119), .B2(new_n1191), .ZN(new_n1193));
  NAND2_X1  g0993(.A1(new_n1094), .A2(new_n1102), .ZN(new_n1194));
  XOR2_X1   g0994(.A(new_n930), .B(KEYINPUT118), .Z(new_n1195));
  NAND3_X1  g0995(.A1(new_n1104), .A2(new_n1194), .A3(new_n1195), .ZN(new_n1196));
  NAND2_X1  g0996(.A1(new_n1193), .A2(new_n1196), .ZN(G381));
  OR3_X1    g0997(.A1(G393), .A2(G396), .A3(G384), .ZN(new_n1198));
  NOR4_X1   g0998(.A1(G387), .A2(G390), .A3(G381), .A4(new_n1198), .ZN(new_n1199));
  INV_X1    g0999(.A(G378), .ZN(new_n1200));
  NAND4_X1  g1000(.A1(new_n1199), .A2(new_n1200), .A3(new_n1175), .A4(new_n1145), .ZN(G407));
  NAND2_X1  g1001(.A1(new_n636), .A2(G213), .ZN(new_n1202));
  OR3_X1    g1002(.A1(G375), .A2(G378), .A3(new_n1202), .ZN(new_n1203));
  NAND3_X1  g1003(.A1(G407), .A2(G213), .A3(new_n1203), .ZN(G409));
  INV_X1    g1004(.A(KEYINPUT125), .ZN(new_n1205));
  INV_X1    g1005(.A(new_n1195), .ZN(new_n1206));
  NOR3_X1   g1006(.A1(new_n1137), .A2(new_n1138), .A3(new_n1206), .ZN(new_n1207));
  NOR2_X1   g1007(.A1(new_n1207), .A2(new_n1174), .ZN(new_n1208));
  OAI21_X1  g1008(.A(KEYINPUT120), .B1(new_n1208), .B2(G378), .ZN(new_n1209));
  NAND4_X1  g1009(.A1(new_n1143), .A2(new_n1136), .A3(new_n1130), .A4(new_n1195), .ZN(new_n1210));
  NAND3_X1  g1010(.A1(new_n1210), .A2(new_n1146), .A3(new_n1173), .ZN(new_n1211));
  OAI21_X1  g1011(.A(new_n656), .B1(new_n1141), .B2(new_n1142), .ZN(new_n1212));
  NAND2_X1  g1012(.A1(new_n1212), .A2(KEYINPUT113), .ZN(new_n1213));
  NAND2_X1  g1013(.A1(new_n1114), .A2(new_n1115), .ZN(new_n1214));
  NAND3_X1  g1014(.A1(new_n1213), .A2(new_n1214), .A3(new_n1105), .ZN(new_n1215));
  INV_X1    g1015(.A(KEYINPUT120), .ZN(new_n1216));
  NAND4_X1  g1016(.A1(new_n1211), .A2(new_n1215), .A3(new_n1216), .A4(new_n1087), .ZN(new_n1217));
  NAND3_X1  g1017(.A1(new_n1145), .A2(G378), .A3(new_n1175), .ZN(new_n1218));
  NAND3_X1  g1018(.A1(new_n1209), .A2(new_n1217), .A3(new_n1218), .ZN(new_n1219));
  AOI21_X1  g1019(.A(KEYINPUT121), .B1(new_n1094), .B2(new_n1102), .ZN(new_n1220));
  INV_X1    g1020(.A(KEYINPUT60), .ZN(new_n1221));
  AND2_X1   g1021(.A1(new_n1220), .A2(new_n1221), .ZN(new_n1222));
  OAI211_X1 g1022(.A(new_n1104), .B(new_n656), .C1(new_n1220), .C2(new_n1221), .ZN(new_n1223));
  OAI21_X1  g1023(.A(new_n1193), .B1(new_n1222), .B2(new_n1223), .ZN(new_n1224));
  XNOR2_X1  g1024(.A(new_n1224), .B(G384), .ZN(new_n1225));
  NAND3_X1  g1025(.A1(new_n1219), .A2(new_n1202), .A3(new_n1225), .ZN(new_n1226));
  INV_X1    g1026(.A(KEYINPUT122), .ZN(new_n1227));
  NAND2_X1  g1027(.A1(new_n1226), .A2(new_n1227), .ZN(new_n1228));
  INV_X1    g1028(.A(KEYINPUT62), .ZN(new_n1229));
  NAND4_X1  g1029(.A1(new_n1219), .A2(KEYINPUT122), .A3(new_n1202), .A4(new_n1225), .ZN(new_n1230));
  AND3_X1   g1030(.A1(new_n1228), .A2(new_n1229), .A3(new_n1230), .ZN(new_n1231));
  NAND2_X1  g1031(.A1(new_n1219), .A2(new_n1202), .ZN(new_n1232));
  OR2_X1    g1032(.A1(new_n1224), .A2(new_n796), .ZN(new_n1233));
  NAND2_X1  g1033(.A1(new_n1224), .A2(new_n796), .ZN(new_n1234));
  AOI21_X1  g1034(.A(KEYINPUT123), .B1(new_n1233), .B2(new_n1234), .ZN(new_n1235));
  NAND2_X1  g1035(.A1(new_n1225), .A2(KEYINPUT123), .ZN(new_n1236));
  INV_X1    g1036(.A(G2897), .ZN(new_n1237));
  NOR2_X1   g1037(.A1(new_n1202), .A2(new_n1237), .ZN(new_n1238));
  AOI21_X1  g1038(.A(new_n1235), .B1(new_n1236), .B2(new_n1238), .ZN(new_n1239));
  NOR4_X1   g1039(.A1(new_n1225), .A2(KEYINPUT123), .A3(new_n1237), .A4(new_n1202), .ZN(new_n1240));
  NOR2_X1   g1040(.A1(new_n1239), .A2(new_n1240), .ZN(new_n1241));
  AOI21_X1  g1041(.A(KEYINPUT61), .B1(new_n1232), .B2(new_n1241), .ZN(new_n1242));
  NAND2_X1  g1042(.A1(new_n1226), .A2(KEYINPUT62), .ZN(new_n1243));
  NAND2_X1  g1043(.A1(new_n1242), .A2(new_n1243), .ZN(new_n1244));
  OAI21_X1  g1044(.A(new_n1205), .B1(new_n1231), .B2(new_n1244), .ZN(new_n1245));
  AOI21_X1  g1045(.A(G390), .B1(new_n945), .B2(new_n975), .ZN(new_n1246));
  INV_X1    g1046(.A(new_n1246), .ZN(new_n1247));
  NAND3_X1  g1047(.A1(new_n945), .A2(G390), .A3(new_n975), .ZN(new_n1248));
  NAND2_X1  g1048(.A1(new_n1247), .A2(new_n1248), .ZN(new_n1249));
  XNOR2_X1  g1049(.A(G393), .B(G396), .ZN(new_n1250));
  OAI21_X1  g1050(.A(new_n1250), .B1(new_n1246), .B2(KEYINPUT124), .ZN(new_n1251));
  NAND2_X1  g1051(.A1(new_n1249), .A2(new_n1251), .ZN(new_n1252));
  NAND4_X1  g1052(.A1(new_n1247), .A2(new_n1248), .A3(KEYINPUT124), .A4(new_n1250), .ZN(new_n1253));
  NAND2_X1  g1053(.A1(new_n1252), .A2(new_n1253), .ZN(new_n1254));
  INV_X1    g1054(.A(new_n1254), .ZN(new_n1255));
  NAND3_X1  g1055(.A1(new_n1228), .A2(new_n1229), .A3(new_n1230), .ZN(new_n1256));
  NAND4_X1  g1056(.A1(new_n1256), .A2(KEYINPUT125), .A3(new_n1242), .A4(new_n1243), .ZN(new_n1257));
  NAND3_X1  g1057(.A1(new_n1245), .A2(new_n1255), .A3(new_n1257), .ZN(new_n1258));
  NAND4_X1  g1058(.A1(new_n1219), .A2(KEYINPUT63), .A3(new_n1202), .A4(new_n1225), .ZN(new_n1259));
  AND3_X1   g1059(.A1(new_n1254), .A2(new_n1259), .A3(new_n1242), .ZN(new_n1260));
  AND2_X1   g1060(.A1(new_n1228), .A2(new_n1230), .ZN(new_n1261));
  OAI21_X1  g1061(.A(new_n1260), .B1(new_n1261), .B2(KEYINPUT63), .ZN(new_n1262));
  NAND2_X1  g1062(.A1(new_n1258), .A2(new_n1262), .ZN(G405));
  OR2_X1    g1063(.A1(new_n1254), .A2(KEYINPUT126), .ZN(new_n1264));
  NAND2_X1  g1064(.A1(new_n1254), .A2(KEYINPUT126), .ZN(new_n1265));
  INV_X1    g1065(.A(new_n1225), .ZN(new_n1266));
  NAND2_X1  g1066(.A1(G375), .A2(new_n1200), .ZN(new_n1267));
  AOI21_X1  g1067(.A(new_n1266), .B1(new_n1267), .B2(new_n1218), .ZN(new_n1268));
  NAND3_X1  g1068(.A1(new_n1267), .A2(new_n1218), .A3(new_n1266), .ZN(new_n1269));
  INV_X1    g1069(.A(new_n1269), .ZN(new_n1270));
  OAI211_X1 g1070(.A(new_n1264), .B(new_n1265), .C1(new_n1268), .C2(new_n1270), .ZN(new_n1271));
  OR3_X1    g1071(.A1(new_n1265), .A2(new_n1268), .A3(new_n1270), .ZN(new_n1272));
  NAND2_X1  g1072(.A1(new_n1271), .A2(new_n1272), .ZN(G402));
endmodule


