//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 0 1 1 1 1 1 0 1 0 0 1 1 1 0 0 0 0 0 1 1 1 1 1 0 1 0 1 0 1 1 1 0 1 1 1 0 0 1 1 1 0 1 0 1 0 0 1 1 1 1 0 1 1 1 1 0 1 0 1 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:18:36 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n672, new_n673,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n705, new_n706, new_n707, new_n708, new_n709, new_n710,
    new_n711, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n730, new_n731, new_n732, new_n734,
    new_n735, new_n736, new_n737, new_n739, new_n740, new_n741, new_n743,
    new_n744, new_n745, new_n746, new_n747, new_n748, new_n749, new_n750,
    new_n751, new_n752, new_n754, new_n756, new_n757, new_n758, new_n759,
    new_n760, new_n761, new_n762, new_n763, new_n764, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n773, new_n774, new_n775,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n835, new_n836, new_n837, new_n839, new_n840, new_n842, new_n843,
    new_n844, new_n845, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n909,
    new_n910, new_n912, new_n913, new_n914, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n925, new_n926,
    new_n928, new_n929, new_n930, new_n931, new_n932, new_n933, new_n934,
    new_n935, new_n937, new_n938, new_n939, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n948, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n956, new_n957, new_n958, new_n959,
    new_n960, new_n961, new_n962, new_n963, new_n964, new_n965, new_n966,
    new_n968, new_n969, new_n970, new_n971;
  XNOR2_X1  g000(.A(G113gat), .B(G141gat), .ZN(new_n202));
  XNOR2_X1  g001(.A(new_n202), .B(G197gat), .ZN(new_n203));
  XOR2_X1   g002(.A(KEYINPUT11), .B(G169gat), .Z(new_n204));
  XNOR2_X1  g003(.A(new_n203), .B(new_n204), .ZN(new_n205));
  XNOR2_X1  g004(.A(new_n205), .B(KEYINPUT12), .ZN(new_n206));
  XOR2_X1   g005(.A(new_n206), .B(KEYINPUT86), .Z(new_n207));
  INV_X1    g006(.A(KEYINPUT87), .ZN(new_n208));
  INV_X1    g007(.A(G50gat), .ZN(new_n209));
  OAI21_X1  g008(.A(new_n208), .B1(new_n209), .B2(G43gat), .ZN(new_n210));
  NAND2_X1  g009(.A1(new_n209), .A2(G43gat), .ZN(new_n211));
  INV_X1    g010(.A(G43gat), .ZN(new_n212));
  NAND3_X1  g011(.A1(new_n212), .A2(KEYINPUT87), .A3(G50gat), .ZN(new_n213));
  NAND3_X1  g012(.A1(new_n210), .A2(new_n211), .A3(new_n213), .ZN(new_n214));
  INV_X1    g013(.A(KEYINPUT15), .ZN(new_n215));
  NAND2_X1  g014(.A1(new_n214), .A2(new_n215), .ZN(new_n216));
  INV_X1    g015(.A(KEYINPUT88), .ZN(new_n217));
  NAND2_X1  g016(.A1(new_n216), .A2(new_n217), .ZN(new_n218));
  NAND2_X1  g017(.A1(new_n212), .A2(G50gat), .ZN(new_n219));
  NAND3_X1  g018(.A1(new_n211), .A2(new_n219), .A3(KEYINPUT15), .ZN(new_n220));
  INV_X1    g019(.A(KEYINPUT14), .ZN(new_n221));
  INV_X1    g020(.A(G36gat), .ZN(new_n222));
  NOR3_X1   g021(.A1(new_n221), .A2(new_n222), .A3(G29gat), .ZN(new_n223));
  INV_X1    g022(.A(new_n223), .ZN(new_n224));
  NAND2_X1  g023(.A1(KEYINPUT14), .A2(G29gat), .ZN(new_n225));
  INV_X1    g024(.A(new_n225), .ZN(new_n226));
  NOR2_X1   g025(.A1(KEYINPUT14), .A2(G29gat), .ZN(new_n227));
  OAI21_X1  g026(.A(new_n222), .B1(new_n226), .B2(new_n227), .ZN(new_n228));
  NAND2_X1  g027(.A1(new_n224), .A2(new_n228), .ZN(new_n229));
  NAND3_X1  g028(.A1(new_n214), .A2(KEYINPUT88), .A3(new_n215), .ZN(new_n230));
  NAND4_X1  g029(.A1(new_n218), .A2(new_n220), .A3(new_n229), .A4(new_n230), .ZN(new_n231));
  INV_X1    g030(.A(KEYINPUT89), .ZN(new_n232));
  OAI21_X1  g031(.A(new_n232), .B1(new_n229), .B2(new_n220), .ZN(new_n233));
  INV_X1    g032(.A(new_n233), .ZN(new_n234));
  NOR2_X1   g033(.A1(new_n231), .A2(new_n234), .ZN(new_n235));
  INV_X1    g034(.A(G29gat), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n221), .A2(new_n236), .ZN(new_n237));
  AOI21_X1  g036(.A(G36gat), .B1(new_n237), .B2(new_n225), .ZN(new_n238));
  OAI21_X1  g037(.A(new_n220), .B1(new_n238), .B2(new_n223), .ZN(new_n239));
  AOI21_X1  g038(.A(new_n239), .B1(new_n217), .B2(new_n216), .ZN(new_n240));
  AOI21_X1  g039(.A(new_n233), .B1(new_n240), .B2(new_n230), .ZN(new_n241));
  NOR2_X1   g040(.A1(new_n235), .A2(new_n241), .ZN(new_n242));
  INV_X1    g041(.A(KEYINPUT92), .ZN(new_n243));
  XNOR2_X1  g042(.A(G15gat), .B(G22gat), .ZN(new_n244));
  NAND2_X1  g043(.A1(new_n244), .A2(KEYINPUT90), .ZN(new_n245));
  INV_X1    g044(.A(G1gat), .ZN(new_n246));
  NAND2_X1  g045(.A1(new_n245), .A2(new_n246), .ZN(new_n247));
  NAND3_X1  g046(.A1(new_n244), .A2(KEYINPUT90), .A3(G1gat), .ZN(new_n248));
  INV_X1    g047(.A(KEYINPUT16), .ZN(new_n249));
  NAND2_X1  g048(.A1(new_n244), .A2(new_n249), .ZN(new_n250));
  NAND3_X1  g049(.A1(new_n247), .A2(new_n248), .A3(new_n250), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n251), .A2(G8gat), .ZN(new_n252));
  INV_X1    g051(.A(new_n252), .ZN(new_n253));
  NOR2_X1   g052(.A1(new_n251), .A2(G8gat), .ZN(new_n254));
  OAI21_X1  g053(.A(new_n243), .B1(new_n253), .B2(new_n254), .ZN(new_n255));
  INV_X1    g054(.A(new_n254), .ZN(new_n256));
  NAND3_X1  g055(.A1(new_n256), .A2(KEYINPUT92), .A3(new_n252), .ZN(new_n257));
  NAND3_X1  g056(.A1(new_n242), .A2(new_n255), .A3(new_n257), .ZN(new_n258));
  NAND2_X1  g057(.A1(G229gat), .A2(G233gat), .ZN(new_n259));
  AND3_X1   g058(.A1(new_n258), .A2(KEYINPUT18), .A3(new_n259), .ZN(new_n260));
  INV_X1    g059(.A(KEYINPUT17), .ZN(new_n261));
  OAI21_X1  g060(.A(new_n261), .B1(new_n235), .B2(new_n241), .ZN(new_n262));
  NAND2_X1  g061(.A1(new_n231), .A2(new_n234), .ZN(new_n263));
  NAND3_X1  g062(.A1(new_n240), .A2(new_n233), .A3(new_n230), .ZN(new_n264));
  NAND3_X1  g063(.A1(new_n263), .A2(new_n264), .A3(KEYINPUT17), .ZN(new_n265));
  NAND2_X1  g064(.A1(new_n262), .A2(new_n265), .ZN(new_n266));
  NAND2_X1  g065(.A1(new_n256), .A2(new_n252), .ZN(new_n267));
  INV_X1    g066(.A(new_n267), .ZN(new_n268));
  AOI21_X1  g067(.A(KEYINPUT91), .B1(new_n266), .B2(new_n268), .ZN(new_n269));
  INV_X1    g068(.A(KEYINPUT91), .ZN(new_n270));
  AOI211_X1 g069(.A(new_n270), .B(new_n267), .C1(new_n262), .C2(new_n265), .ZN(new_n271));
  OAI21_X1  g070(.A(new_n260), .B1(new_n269), .B2(new_n271), .ZN(new_n272));
  NAND2_X1  g071(.A1(new_n255), .A2(new_n257), .ZN(new_n273));
  NAND2_X1  g072(.A1(new_n263), .A2(new_n264), .ZN(new_n274));
  NAND2_X1  g073(.A1(new_n273), .A2(new_n274), .ZN(new_n275));
  NAND2_X1  g074(.A1(new_n275), .A2(new_n258), .ZN(new_n276));
  XOR2_X1   g075(.A(new_n259), .B(KEYINPUT13), .Z(new_n277));
  NAND2_X1  g076(.A1(new_n276), .A2(new_n277), .ZN(new_n278));
  NAND2_X1  g077(.A1(new_n272), .A2(new_n278), .ZN(new_n279));
  XNOR2_X1  g078(.A(KEYINPUT93), .B(KEYINPUT18), .ZN(new_n280));
  INV_X1    g079(.A(new_n280), .ZN(new_n281));
  AND3_X1   g080(.A1(new_n263), .A2(new_n264), .A3(KEYINPUT17), .ZN(new_n282));
  AOI21_X1  g081(.A(KEYINPUT17), .B1(new_n263), .B2(new_n264), .ZN(new_n283));
  OAI21_X1  g082(.A(new_n268), .B1(new_n282), .B2(new_n283), .ZN(new_n284));
  NAND2_X1  g083(.A1(new_n284), .A2(new_n270), .ZN(new_n285));
  NAND3_X1  g084(.A1(new_n266), .A2(KEYINPUT91), .A3(new_n268), .ZN(new_n286));
  NAND2_X1  g085(.A1(new_n285), .A2(new_n286), .ZN(new_n287));
  AND2_X1   g086(.A1(new_n258), .A2(new_n259), .ZN(new_n288));
  AOI21_X1  g087(.A(new_n281), .B1(new_n287), .B2(new_n288), .ZN(new_n289));
  OAI21_X1  g088(.A(new_n207), .B1(new_n279), .B2(new_n289), .ZN(new_n290));
  AOI22_X1  g089(.A1(new_n287), .A2(new_n260), .B1(new_n276), .B2(new_n277), .ZN(new_n291));
  OAI21_X1  g090(.A(new_n288), .B1(new_n269), .B2(new_n271), .ZN(new_n292));
  NAND2_X1  g091(.A1(new_n292), .A2(new_n280), .ZN(new_n293));
  NAND3_X1  g092(.A1(new_n291), .A2(new_n293), .A3(new_n206), .ZN(new_n294));
  NAND2_X1  g093(.A1(new_n290), .A2(new_n294), .ZN(new_n295));
  INV_X1    g094(.A(new_n295), .ZN(new_n296));
  XOR2_X1   g095(.A(G141gat), .B(G148gat), .Z(new_n297));
  INV_X1    g096(.A(G155gat), .ZN(new_n298));
  INV_X1    g097(.A(G162gat), .ZN(new_n299));
  OAI21_X1  g098(.A(KEYINPUT2), .B1(new_n298), .B2(new_n299), .ZN(new_n300));
  NAND2_X1  g099(.A1(new_n297), .A2(new_n300), .ZN(new_n301));
  XNOR2_X1  g100(.A(G155gat), .B(G162gat), .ZN(new_n302));
  INV_X1    g101(.A(new_n302), .ZN(new_n303));
  NAND2_X1  g102(.A1(new_n301), .A2(new_n303), .ZN(new_n304));
  NAND3_X1  g103(.A1(new_n297), .A2(new_n302), .A3(new_n300), .ZN(new_n305));
  NAND2_X1  g104(.A1(new_n304), .A2(new_n305), .ZN(new_n306));
  XNOR2_X1  g105(.A(G197gat), .B(G204gat), .ZN(new_n307));
  INV_X1    g106(.A(KEYINPUT22), .ZN(new_n308));
  INV_X1    g107(.A(G211gat), .ZN(new_n309));
  INV_X1    g108(.A(G218gat), .ZN(new_n310));
  OAI21_X1  g109(.A(new_n308), .B1(new_n309), .B2(new_n310), .ZN(new_n311));
  NAND2_X1  g110(.A1(new_n307), .A2(new_n311), .ZN(new_n312));
  XNOR2_X1  g111(.A(G211gat), .B(G218gat), .ZN(new_n313));
  INV_X1    g112(.A(new_n313), .ZN(new_n314));
  NAND2_X1  g113(.A1(new_n312), .A2(new_n314), .ZN(new_n315));
  NAND3_X1  g114(.A1(new_n313), .A2(new_n307), .A3(new_n311), .ZN(new_n316));
  AOI21_X1  g115(.A(KEYINPUT29), .B1(new_n315), .B2(new_n316), .ZN(new_n317));
  INV_X1    g116(.A(KEYINPUT80), .ZN(new_n318));
  AND2_X1   g117(.A1(new_n317), .A2(new_n318), .ZN(new_n319));
  INV_X1    g118(.A(KEYINPUT3), .ZN(new_n320));
  OAI21_X1  g119(.A(new_n320), .B1(new_n317), .B2(new_n318), .ZN(new_n321));
  OAI21_X1  g120(.A(new_n306), .B1(new_n319), .B2(new_n321), .ZN(new_n322));
  INV_X1    g121(.A(G228gat), .ZN(new_n323));
  INV_X1    g122(.A(G233gat), .ZN(new_n324));
  NOR2_X1   g123(.A1(new_n323), .A2(new_n324), .ZN(new_n325));
  INV_X1    g124(.A(new_n325), .ZN(new_n326));
  NAND3_X1  g125(.A1(new_n304), .A2(new_n320), .A3(new_n305), .ZN(new_n327));
  XOR2_X1   g126(.A(KEYINPUT78), .B(KEYINPUT29), .Z(new_n328));
  NAND2_X1  g127(.A1(new_n327), .A2(new_n328), .ZN(new_n329));
  NAND2_X1  g128(.A1(new_n315), .A2(new_n316), .ZN(new_n330));
  INV_X1    g129(.A(new_n330), .ZN(new_n331));
  AOI21_X1  g130(.A(new_n326), .B1(new_n329), .B2(new_n331), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n322), .A2(new_n332), .ZN(new_n333));
  INV_X1    g132(.A(KEYINPUT81), .ZN(new_n334));
  NAND2_X1  g133(.A1(new_n333), .A2(new_n334), .ZN(new_n335));
  NAND3_X1  g134(.A1(new_n322), .A2(KEYINPUT81), .A3(new_n332), .ZN(new_n336));
  NAND2_X1  g135(.A1(new_n335), .A2(new_n336), .ZN(new_n337));
  AND2_X1   g136(.A1(new_n330), .A2(new_n328), .ZN(new_n338));
  OAI21_X1  g137(.A(new_n306), .B1(new_n338), .B2(KEYINPUT3), .ZN(new_n339));
  NAND2_X1  g138(.A1(new_n329), .A2(new_n331), .ZN(new_n340));
  AOI21_X1  g139(.A(new_n325), .B1(new_n339), .B2(new_n340), .ZN(new_n341));
  INV_X1    g140(.A(new_n341), .ZN(new_n342));
  NAND2_X1  g141(.A1(new_n337), .A2(new_n342), .ZN(new_n343));
  XOR2_X1   g142(.A(KEYINPUT31), .B(G50gat), .Z(new_n344));
  NAND2_X1  g143(.A1(new_n343), .A2(new_n344), .ZN(new_n345));
  XNOR2_X1  g144(.A(G78gat), .B(G106gat), .ZN(new_n346));
  XNOR2_X1  g145(.A(new_n346), .B(G22gat), .ZN(new_n347));
  INV_X1    g146(.A(new_n344), .ZN(new_n348));
  NAND3_X1  g147(.A1(new_n337), .A2(new_n348), .A3(new_n342), .ZN(new_n349));
  NAND3_X1  g148(.A1(new_n345), .A2(new_n347), .A3(new_n349), .ZN(new_n350));
  INV_X1    g149(.A(new_n347), .ZN(new_n351));
  AOI21_X1  g150(.A(new_n348), .B1(new_n337), .B2(new_n342), .ZN(new_n352));
  AOI211_X1 g151(.A(new_n344), .B(new_n341), .C1(new_n335), .C2(new_n336), .ZN(new_n353));
  OAI21_X1  g152(.A(new_n351), .B1(new_n352), .B2(new_n353), .ZN(new_n354));
  NAND2_X1  g153(.A1(new_n350), .A2(new_n354), .ZN(new_n355));
  INV_X1    g154(.A(KEYINPUT73), .ZN(new_n356));
  INV_X1    g155(.A(G227gat), .ZN(new_n357));
  NOR2_X1   g156(.A1(new_n357), .A2(new_n324), .ZN(new_n358));
  INV_X1    g157(.A(new_n358), .ZN(new_n359));
  INV_X1    g158(.A(KEYINPUT70), .ZN(new_n360));
  NAND2_X1  g159(.A1(G183gat), .A2(G190gat), .ZN(new_n361));
  NAND2_X1  g160(.A1(new_n361), .A2(KEYINPUT24), .ZN(new_n362));
  INV_X1    g161(.A(KEYINPUT24), .ZN(new_n363));
  NAND3_X1  g162(.A1(new_n363), .A2(G183gat), .A3(G190gat), .ZN(new_n364));
  AND2_X1   g163(.A1(new_n362), .A2(new_n364), .ZN(new_n365));
  AND2_X1   g164(.A1(KEYINPUT69), .A2(G183gat), .ZN(new_n366));
  NOR2_X1   g165(.A1(KEYINPUT69), .A2(G183gat), .ZN(new_n367));
  NOR3_X1   g166(.A1(new_n366), .A2(new_n367), .A3(G190gat), .ZN(new_n368));
  OAI21_X1  g167(.A(new_n360), .B1(new_n365), .B2(new_n368), .ZN(new_n369));
  NOR2_X1   g168(.A1(G169gat), .A2(G176gat), .ZN(new_n370));
  INV_X1    g169(.A(KEYINPUT68), .ZN(new_n371));
  NAND2_X1  g170(.A1(new_n370), .A2(new_n371), .ZN(new_n372));
  OAI21_X1  g171(.A(KEYINPUT68), .B1(G169gat), .B2(G176gat), .ZN(new_n373));
  NAND3_X1  g172(.A1(new_n372), .A2(KEYINPUT23), .A3(new_n373), .ZN(new_n374));
  INV_X1    g173(.A(KEYINPUT66), .ZN(new_n375));
  OAI21_X1  g174(.A(new_n375), .B1(new_n370), .B2(KEYINPUT23), .ZN(new_n376));
  INV_X1    g175(.A(KEYINPUT23), .ZN(new_n377));
  OAI211_X1 g176(.A(new_n377), .B(KEYINPUT66), .C1(G169gat), .C2(G176gat), .ZN(new_n378));
  NAND2_X1  g177(.A1(G169gat), .A2(G176gat), .ZN(new_n379));
  NAND2_X1  g178(.A1(new_n379), .A2(KEYINPUT67), .ZN(new_n380));
  INV_X1    g179(.A(KEYINPUT67), .ZN(new_n381));
  NAND3_X1  g180(.A1(new_n381), .A2(G169gat), .A3(G176gat), .ZN(new_n382));
  AOI22_X1  g181(.A1(new_n376), .A2(new_n378), .B1(new_n380), .B2(new_n382), .ZN(new_n383));
  NAND2_X1  g182(.A1(new_n362), .A2(new_n364), .ZN(new_n384));
  XNOR2_X1  g183(.A(KEYINPUT69), .B(G183gat), .ZN(new_n385));
  OAI211_X1 g184(.A(new_n384), .B(KEYINPUT70), .C1(G190gat), .C2(new_n385), .ZN(new_n386));
  NAND4_X1  g185(.A1(new_n369), .A2(new_n374), .A3(new_n383), .A4(new_n386), .ZN(new_n387));
  NAND2_X1  g186(.A1(new_n387), .A2(KEYINPUT25), .ZN(new_n388));
  INV_X1    g187(.A(KEYINPUT26), .ZN(new_n389));
  NAND3_X1  g188(.A1(new_n372), .A2(new_n389), .A3(new_n373), .ZN(new_n390));
  OAI211_X1 g189(.A(KEYINPUT71), .B(KEYINPUT26), .C1(G169gat), .C2(G176gat), .ZN(new_n391));
  NAND2_X1  g190(.A1(new_n380), .A2(new_n382), .ZN(new_n392));
  INV_X1    g191(.A(KEYINPUT71), .ZN(new_n393));
  OAI21_X1  g192(.A(new_n393), .B1(new_n370), .B2(new_n389), .ZN(new_n394));
  NAND4_X1  g193(.A1(new_n390), .A2(new_n391), .A3(new_n392), .A4(new_n394), .ZN(new_n395));
  OAI21_X1  g194(.A(KEYINPUT27), .B1(new_n366), .B2(new_n367), .ZN(new_n396));
  OR2_X1    g195(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n397));
  NAND2_X1  g196(.A1(new_n396), .A2(new_n397), .ZN(new_n398));
  INV_X1    g197(.A(G190gat), .ZN(new_n399));
  AOI21_X1  g198(.A(KEYINPUT28), .B1(new_n398), .B2(new_n399), .ZN(new_n400));
  XOR2_X1   g199(.A(KEYINPUT27), .B(G183gat), .Z(new_n401));
  INV_X1    g200(.A(KEYINPUT28), .ZN(new_n402));
  NOR3_X1   g201(.A1(new_n401), .A2(new_n402), .A3(G190gat), .ZN(new_n403));
  OAI211_X1 g202(.A(new_n361), .B(new_n395), .C1(new_n400), .C2(new_n403), .ZN(new_n404));
  INV_X1    g203(.A(KEYINPUT64), .ZN(new_n405));
  OR3_X1    g204(.A1(new_n405), .A2(G183gat), .A3(G190gat), .ZN(new_n406));
  OAI21_X1  g205(.A(new_n405), .B1(G183gat), .B2(G190gat), .ZN(new_n407));
  NAND3_X1  g206(.A1(new_n384), .A2(new_n406), .A3(new_n407), .ZN(new_n408));
  AND2_X1   g207(.A1(KEYINPUT65), .A2(G169gat), .ZN(new_n409));
  NOR2_X1   g208(.A1(KEYINPUT65), .A2(G169gat), .ZN(new_n410));
  NOR2_X1   g209(.A1(new_n409), .A2(new_n410), .ZN(new_n411));
  NOR2_X1   g210(.A1(new_n377), .A2(G176gat), .ZN(new_n412));
  AOI21_X1  g211(.A(KEYINPUT25), .B1(new_n411), .B2(new_n412), .ZN(new_n413));
  AND3_X1   g212(.A1(new_n383), .A2(new_n408), .A3(new_n413), .ZN(new_n414));
  INV_X1    g213(.A(new_n414), .ZN(new_n415));
  NAND3_X1  g214(.A1(new_n388), .A2(new_n404), .A3(new_n415), .ZN(new_n416));
  XNOR2_X1  g215(.A(G113gat), .B(G120gat), .ZN(new_n417));
  INV_X1    g216(.A(KEYINPUT72), .ZN(new_n418));
  INV_X1    g217(.A(KEYINPUT1), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n418), .A2(new_n419), .ZN(new_n420));
  NOR2_X1   g219(.A1(new_n417), .A2(new_n420), .ZN(new_n421));
  XNOR2_X1  g220(.A(G127gat), .B(G134gat), .ZN(new_n422));
  NAND2_X1  g221(.A1(new_n421), .A2(new_n422), .ZN(new_n423));
  INV_X1    g222(.A(new_n422), .ZN(new_n424));
  OAI21_X1  g223(.A(new_n424), .B1(new_n417), .B2(new_n420), .ZN(new_n425));
  NAND2_X1  g224(.A1(new_n423), .A2(new_n425), .ZN(new_n426));
  NAND2_X1  g225(.A1(new_n416), .A2(new_n426), .ZN(new_n427));
  AOI21_X1  g226(.A(new_n414), .B1(new_n387), .B2(KEYINPUT25), .ZN(new_n428));
  INV_X1    g227(.A(new_n426), .ZN(new_n429));
  NAND3_X1  g228(.A1(new_n428), .A2(new_n429), .A3(new_n404), .ZN(new_n430));
  AOI21_X1  g229(.A(new_n359), .B1(new_n427), .B2(new_n430), .ZN(new_n431));
  OAI21_X1  g230(.A(new_n356), .B1(new_n431), .B2(KEYINPUT33), .ZN(new_n432));
  XOR2_X1   g231(.A(G15gat), .B(G43gat), .Z(new_n433));
  XNOR2_X1  g232(.A(new_n433), .B(KEYINPUT74), .ZN(new_n434));
  XNOR2_X1  g233(.A(G71gat), .B(G99gat), .ZN(new_n435));
  XNOR2_X1  g234(.A(new_n434), .B(new_n435), .ZN(new_n436));
  AND4_X1   g235(.A1(new_n429), .A2(new_n388), .A3(new_n404), .A4(new_n415), .ZN(new_n437));
  AOI21_X1  g236(.A(new_n429), .B1(new_n428), .B2(new_n404), .ZN(new_n438));
  OAI21_X1  g237(.A(new_n358), .B1(new_n437), .B2(new_n438), .ZN(new_n439));
  AOI21_X1  g238(.A(new_n436), .B1(new_n439), .B2(KEYINPUT32), .ZN(new_n440));
  INV_X1    g239(.A(KEYINPUT33), .ZN(new_n441));
  NAND3_X1  g240(.A1(new_n439), .A2(KEYINPUT73), .A3(new_n441), .ZN(new_n442));
  NAND3_X1  g241(.A1(new_n432), .A2(new_n440), .A3(new_n442), .ZN(new_n443));
  INV_X1    g242(.A(KEYINPUT75), .ZN(new_n444));
  AOI21_X1  g243(.A(new_n441), .B1(new_n436), .B2(new_n444), .ZN(new_n445));
  OAI21_X1  g244(.A(new_n445), .B1(new_n444), .B2(new_n436), .ZN(new_n446));
  NAND3_X1  g245(.A1(new_n439), .A2(new_n446), .A3(KEYINPUT32), .ZN(new_n447));
  NAND2_X1  g246(.A1(new_n443), .A2(new_n447), .ZN(new_n448));
  INV_X1    g247(.A(KEYINPUT77), .ZN(new_n449));
  NAND2_X1  g248(.A1(new_n448), .A2(new_n449), .ZN(new_n450));
  NAND3_X1  g249(.A1(new_n443), .A2(KEYINPUT77), .A3(new_n447), .ZN(new_n451));
  INV_X1    g250(.A(KEYINPUT34), .ZN(new_n452));
  NAND4_X1  g251(.A1(new_n427), .A2(new_n452), .A3(new_n359), .A4(new_n430), .ZN(new_n453));
  XNOR2_X1  g252(.A(new_n453), .B(KEYINPUT76), .ZN(new_n454));
  NAND3_X1  g253(.A1(new_n427), .A2(new_n359), .A3(new_n430), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n455), .A2(KEYINPUT34), .ZN(new_n456));
  NAND2_X1  g255(.A1(new_n454), .A2(new_n456), .ZN(new_n457));
  INV_X1    g256(.A(new_n457), .ZN(new_n458));
  NAND3_X1  g257(.A1(new_n450), .A2(new_n451), .A3(new_n458), .ZN(new_n459));
  NAND4_X1  g258(.A1(new_n457), .A2(KEYINPUT77), .A3(new_n443), .A4(new_n447), .ZN(new_n460));
  NAND2_X1  g259(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  INV_X1    g260(.A(KEYINPUT83), .ZN(new_n462));
  NAND2_X1  g261(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  NAND3_X1  g262(.A1(new_n459), .A2(KEYINPUT83), .A3(new_n460), .ZN(new_n464));
  AOI21_X1  g263(.A(new_n355), .B1(new_n463), .B2(new_n464), .ZN(new_n465));
  XNOR2_X1  g264(.A(KEYINPUT84), .B(KEYINPUT35), .ZN(new_n466));
  XNOR2_X1  g265(.A(G8gat), .B(G36gat), .ZN(new_n467));
  XNOR2_X1  g266(.A(G64gat), .B(G92gat), .ZN(new_n468));
  XOR2_X1   g267(.A(new_n467), .B(new_n468), .Z(new_n469));
  AND2_X1   g268(.A1(G226gat), .A2(G233gat), .ZN(new_n470));
  NAND2_X1  g269(.A1(new_n416), .A2(new_n470), .ZN(new_n471));
  INV_X1    g270(.A(new_n471), .ZN(new_n472));
  AOI21_X1  g271(.A(new_n470), .B1(new_n416), .B2(new_n328), .ZN(new_n473));
  OAI21_X1  g272(.A(new_n331), .B1(new_n472), .B2(new_n473), .ZN(new_n474));
  AOI21_X1  g273(.A(KEYINPUT29), .B1(new_n428), .B2(new_n404), .ZN(new_n475));
  OAI211_X1 g274(.A(new_n471), .B(new_n330), .C1(new_n475), .C2(new_n470), .ZN(new_n476));
  AOI21_X1  g275(.A(new_n469), .B1(new_n474), .B2(new_n476), .ZN(new_n477));
  INV_X1    g276(.A(new_n477), .ZN(new_n478));
  NAND2_X1  g277(.A1(new_n478), .A2(KEYINPUT30), .ZN(new_n479));
  NAND3_X1  g278(.A1(new_n474), .A2(new_n476), .A3(new_n469), .ZN(new_n480));
  INV_X1    g279(.A(new_n480), .ZN(new_n481));
  NAND2_X1  g280(.A1(new_n479), .A2(new_n481), .ZN(new_n482));
  NAND3_X1  g281(.A1(new_n478), .A2(KEYINPUT30), .A3(new_n480), .ZN(new_n483));
  AND2_X1   g282(.A1(new_n482), .A2(new_n483), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n306), .A2(new_n426), .ZN(new_n485));
  NAND4_X1  g284(.A1(new_n304), .A2(new_n423), .A3(new_n305), .A4(new_n425), .ZN(new_n486));
  AND2_X1   g285(.A1(new_n485), .A2(new_n486), .ZN(new_n487));
  NAND2_X1  g286(.A1(G225gat), .A2(G233gat), .ZN(new_n488));
  OAI21_X1  g287(.A(KEYINPUT5), .B1(new_n487), .B2(new_n488), .ZN(new_n489));
  NAND2_X1  g288(.A1(new_n306), .A2(KEYINPUT3), .ZN(new_n490));
  NAND3_X1  g289(.A1(new_n490), .A2(new_n327), .A3(new_n426), .ZN(new_n491));
  INV_X1    g290(.A(new_n486), .ZN(new_n492));
  NAND2_X1  g291(.A1(new_n492), .A2(KEYINPUT4), .ZN(new_n493));
  INV_X1    g292(.A(KEYINPUT4), .ZN(new_n494));
  NAND2_X1  g293(.A1(new_n486), .A2(new_n494), .ZN(new_n495));
  NAND4_X1  g294(.A1(new_n491), .A2(new_n493), .A3(new_n488), .A4(new_n495), .ZN(new_n496));
  NAND2_X1  g295(.A1(new_n489), .A2(new_n496), .ZN(new_n497));
  XNOR2_X1  g296(.A(new_n486), .B(KEYINPUT4), .ZN(new_n498));
  NAND4_X1  g297(.A1(new_n498), .A2(KEYINPUT5), .A3(new_n488), .A4(new_n491), .ZN(new_n499));
  NAND2_X1  g298(.A1(new_n497), .A2(new_n499), .ZN(new_n500));
  XNOR2_X1  g299(.A(G1gat), .B(G29gat), .ZN(new_n501));
  XNOR2_X1  g300(.A(new_n501), .B(KEYINPUT0), .ZN(new_n502));
  XNOR2_X1  g301(.A(G57gat), .B(G85gat), .ZN(new_n503));
  XOR2_X1   g302(.A(new_n502), .B(new_n503), .Z(new_n504));
  AOI21_X1  g303(.A(KEYINPUT6), .B1(new_n500), .B2(new_n504), .ZN(new_n505));
  INV_X1    g304(.A(new_n504), .ZN(new_n506));
  NAND3_X1  g305(.A1(new_n497), .A2(new_n499), .A3(new_n506), .ZN(new_n507));
  NAND2_X1  g306(.A1(new_n505), .A2(new_n507), .ZN(new_n508));
  NAND2_X1  g307(.A1(new_n508), .A2(KEYINPUT82), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n500), .A2(new_n504), .ZN(new_n510));
  INV_X1    g309(.A(KEYINPUT82), .ZN(new_n511));
  INV_X1    g310(.A(KEYINPUT6), .ZN(new_n512));
  NAND4_X1  g311(.A1(new_n510), .A2(new_n511), .A3(new_n512), .A4(new_n507), .ZN(new_n513));
  INV_X1    g312(.A(new_n507), .ZN(new_n514));
  NAND2_X1  g313(.A1(new_n514), .A2(KEYINPUT6), .ZN(new_n515));
  AND2_X1   g314(.A1(new_n513), .A2(new_n515), .ZN(new_n516));
  AOI211_X1 g315(.A(new_n466), .B(new_n484), .C1(new_n509), .C2(new_n516), .ZN(new_n517));
  NAND2_X1  g316(.A1(new_n465), .A2(new_n517), .ZN(new_n518));
  INV_X1    g317(.A(KEYINPUT85), .ZN(new_n519));
  INV_X1    g318(.A(new_n355), .ZN(new_n520));
  AOI21_X1  g319(.A(new_n519), .B1(new_n461), .B2(new_n520), .ZN(new_n521));
  AOI211_X1 g320(.A(KEYINPUT85), .B(new_n355), .C1(new_n459), .C2(new_n460), .ZN(new_n522));
  NAND2_X1  g321(.A1(new_n482), .A2(new_n483), .ZN(new_n523));
  AND2_X1   g322(.A1(new_n505), .A2(KEYINPUT79), .ZN(new_n524));
  OAI21_X1  g323(.A(new_n507), .B1(new_n505), .B2(KEYINPUT79), .ZN(new_n525));
  OAI21_X1  g324(.A(new_n515), .B1(new_n524), .B2(new_n525), .ZN(new_n526));
  NAND2_X1  g325(.A1(new_n523), .A2(new_n526), .ZN(new_n527));
  NOR3_X1   g326(.A1(new_n521), .A2(new_n522), .A3(new_n527), .ZN(new_n528));
  INV_X1    g327(.A(KEYINPUT35), .ZN(new_n529));
  OAI21_X1  g328(.A(new_n518), .B1(new_n528), .B2(new_n529), .ZN(new_n530));
  NAND2_X1  g329(.A1(new_n498), .A2(new_n491), .ZN(new_n531));
  INV_X1    g330(.A(new_n488), .ZN(new_n532));
  NAND2_X1  g331(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  INV_X1    g332(.A(KEYINPUT39), .ZN(new_n534));
  AOI21_X1  g333(.A(new_n534), .B1(new_n487), .B2(new_n488), .ZN(new_n535));
  NAND2_X1  g334(.A1(new_n533), .A2(new_n535), .ZN(new_n536));
  NAND3_X1  g335(.A1(new_n531), .A2(new_n534), .A3(new_n532), .ZN(new_n537));
  NAND3_X1  g336(.A1(new_n536), .A2(new_n504), .A3(new_n537), .ZN(new_n538));
  INV_X1    g337(.A(KEYINPUT40), .ZN(new_n539));
  NOR2_X1   g338(.A1(new_n538), .A2(new_n539), .ZN(new_n540));
  NOR2_X1   g339(.A1(new_n540), .A2(new_n514), .ZN(new_n541));
  NAND2_X1  g340(.A1(new_n538), .A2(new_n539), .ZN(new_n542));
  NAND4_X1  g341(.A1(new_n482), .A2(new_n483), .A3(new_n541), .A4(new_n542), .ZN(new_n543));
  OAI21_X1  g342(.A(new_n330), .B1(new_n472), .B2(new_n473), .ZN(new_n544));
  OAI211_X1 g343(.A(new_n471), .B(new_n331), .C1(new_n475), .C2(new_n470), .ZN(new_n545));
  NAND3_X1  g344(.A1(new_n544), .A2(KEYINPUT37), .A3(new_n545), .ZN(new_n546));
  INV_X1    g345(.A(KEYINPUT38), .ZN(new_n547));
  INV_X1    g346(.A(KEYINPUT37), .ZN(new_n548));
  NOR2_X1   g347(.A1(new_n469), .A2(new_n548), .ZN(new_n549));
  OAI211_X1 g348(.A(new_n546), .B(new_n547), .C1(new_n477), .C2(new_n549), .ZN(new_n550));
  NAND4_X1  g349(.A1(new_n516), .A2(new_n480), .A3(new_n550), .A4(new_n509), .ZN(new_n551));
  OR2_X1    g350(.A1(new_n477), .A2(new_n549), .ZN(new_n552));
  NAND2_X1  g351(.A1(new_n474), .A2(new_n476), .ZN(new_n553));
  NAND2_X1  g352(.A1(new_n553), .A2(KEYINPUT37), .ZN(new_n554));
  AOI21_X1  g353(.A(new_n547), .B1(new_n552), .B2(new_n554), .ZN(new_n555));
  OAI211_X1 g354(.A(new_n520), .B(new_n543), .C1(new_n551), .C2(new_n555), .ZN(new_n556));
  NAND2_X1  g355(.A1(new_n527), .A2(new_n355), .ZN(new_n557));
  NAND2_X1  g356(.A1(new_n556), .A2(new_n557), .ZN(new_n558));
  AND3_X1   g357(.A1(new_n459), .A2(KEYINPUT36), .A3(new_n460), .ZN(new_n559));
  AOI21_X1  g358(.A(KEYINPUT36), .B1(new_n459), .B2(new_n460), .ZN(new_n560));
  NOR3_X1   g359(.A1(new_n558), .A2(new_n559), .A3(new_n560), .ZN(new_n561));
  INV_X1    g360(.A(new_n561), .ZN(new_n562));
  AOI21_X1  g361(.A(new_n296), .B1(new_n530), .B2(new_n562), .ZN(new_n563));
  INV_X1    g362(.A(KEYINPUT9), .ZN(new_n564));
  INV_X1    g363(.A(G71gat), .ZN(new_n565));
  INV_X1    g364(.A(G78gat), .ZN(new_n566));
  OAI21_X1  g365(.A(new_n564), .B1(new_n565), .B2(new_n566), .ZN(new_n567));
  OR2_X1    g366(.A1(G57gat), .A2(G64gat), .ZN(new_n568));
  NAND2_X1  g367(.A1(G57gat), .A2(G64gat), .ZN(new_n569));
  AND2_X1   g368(.A1(new_n568), .A2(new_n569), .ZN(new_n570));
  XNOR2_X1  g369(.A(G71gat), .B(G78gat), .ZN(new_n571));
  INV_X1    g370(.A(new_n571), .ZN(new_n572));
  INV_X1    g371(.A(KEYINPUT94), .ZN(new_n573));
  OAI211_X1 g372(.A(new_n567), .B(new_n570), .C1(new_n572), .C2(new_n573), .ZN(new_n574));
  NAND3_X1  g373(.A1(new_n567), .A2(new_n568), .A3(new_n569), .ZN(new_n575));
  NAND3_X1  g374(.A1(new_n568), .A2(new_n573), .A3(new_n569), .ZN(new_n576));
  NAND3_X1  g375(.A1(new_n575), .A2(new_n576), .A3(new_n571), .ZN(new_n577));
  NAND2_X1  g376(.A1(new_n574), .A2(new_n577), .ZN(new_n578));
  AOI22_X1  g377(.A1(new_n255), .A2(new_n257), .B1(KEYINPUT21), .B2(new_n578), .ZN(new_n579));
  NOR2_X1   g378(.A1(new_n578), .A2(KEYINPUT21), .ZN(new_n580));
  XNOR2_X1  g379(.A(G127gat), .B(G155gat), .ZN(new_n581));
  XNOR2_X1  g380(.A(new_n580), .B(new_n581), .ZN(new_n582));
  XNOR2_X1  g381(.A(new_n579), .B(new_n582), .ZN(new_n583));
  NAND2_X1  g382(.A1(G231gat), .A2(G233gat), .ZN(new_n584));
  XNOR2_X1  g383(.A(new_n584), .B(KEYINPUT95), .ZN(new_n585));
  XOR2_X1   g384(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n586));
  XNOR2_X1  g385(.A(new_n585), .B(new_n586), .ZN(new_n587));
  XNOR2_X1  g386(.A(G183gat), .B(G211gat), .ZN(new_n588));
  XNOR2_X1  g387(.A(new_n587), .B(new_n588), .ZN(new_n589));
  OR2_X1    g388(.A1(new_n583), .A2(new_n589), .ZN(new_n590));
  NAND2_X1  g389(.A1(new_n583), .A2(new_n589), .ZN(new_n591));
  NAND2_X1  g390(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  INV_X1    g391(.A(new_n592), .ZN(new_n593));
  NAND2_X1  g392(.A1(G85gat), .A2(G92gat), .ZN(new_n594));
  XNOR2_X1  g393(.A(new_n594), .B(KEYINPUT7), .ZN(new_n595));
  OR2_X1    g394(.A1(G99gat), .A2(G106gat), .ZN(new_n596));
  NAND2_X1  g395(.A1(G99gat), .A2(G106gat), .ZN(new_n597));
  NAND2_X1  g396(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  INV_X1    g397(.A(G85gat), .ZN(new_n599));
  INV_X1    g398(.A(G92gat), .ZN(new_n600));
  AOI22_X1  g399(.A1(KEYINPUT8), .A2(new_n597), .B1(new_n599), .B2(new_n600), .ZN(new_n601));
  NAND3_X1  g400(.A1(new_n595), .A2(new_n598), .A3(new_n601), .ZN(new_n602));
  INV_X1    g401(.A(new_n602), .ZN(new_n603));
  AOI21_X1  g402(.A(new_n598), .B1(new_n595), .B2(new_n601), .ZN(new_n604));
  NOR2_X1   g403(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  AOI21_X1  g404(.A(new_n605), .B1(new_n262), .B2(new_n265), .ZN(new_n606));
  INV_X1    g405(.A(new_n606), .ZN(new_n607));
  XNOR2_X1  g406(.A(G190gat), .B(G218gat), .ZN(new_n608));
  INV_X1    g407(.A(new_n608), .ZN(new_n609));
  AND2_X1   g408(.A1(G232gat), .A2(G233gat), .ZN(new_n610));
  NAND2_X1  g409(.A1(new_n610), .A2(KEYINPUT41), .ZN(new_n611));
  INV_X1    g410(.A(new_n605), .ZN(new_n612));
  OAI21_X1  g411(.A(new_n611), .B1(new_n274), .B2(new_n612), .ZN(new_n613));
  INV_X1    g412(.A(new_n613), .ZN(new_n614));
  NAND3_X1  g413(.A1(new_n607), .A2(new_n609), .A3(new_n614), .ZN(new_n615));
  OAI21_X1  g414(.A(new_n608), .B1(new_n606), .B2(new_n613), .ZN(new_n616));
  NOR2_X1   g415(.A1(new_n610), .A2(KEYINPUT41), .ZN(new_n617));
  XNOR2_X1  g416(.A(new_n617), .B(G134gat), .ZN(new_n618));
  XNOR2_X1  g417(.A(new_n618), .B(new_n299), .ZN(new_n619));
  NAND4_X1  g418(.A1(new_n615), .A2(new_n616), .A3(KEYINPUT96), .A4(new_n619), .ZN(new_n620));
  INV_X1    g419(.A(new_n620), .ZN(new_n621));
  INV_X1    g420(.A(KEYINPUT96), .ZN(new_n622));
  NAND2_X1  g421(.A1(new_n616), .A2(new_n622), .ZN(new_n623));
  AOI22_X1  g422(.A1(new_n623), .A2(new_n619), .B1(new_n615), .B2(new_n616), .ZN(new_n624));
  NOR2_X1   g423(.A1(new_n621), .A2(new_n624), .ZN(new_n625));
  NOR2_X1   g424(.A1(new_n593), .A2(new_n625), .ZN(new_n626));
  INV_X1    g425(.A(new_n626), .ZN(new_n627));
  INV_X1    g426(.A(new_n604), .ZN(new_n628));
  NAND3_X1  g427(.A1(new_n578), .A2(new_n628), .A3(new_n602), .ZN(new_n629));
  OAI211_X1 g428(.A(new_n574), .B(new_n577), .C1(new_n603), .C2(new_n604), .ZN(new_n630));
  NAND2_X1  g429(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  NAND2_X1  g430(.A1(G230gat), .A2(G233gat), .ZN(new_n632));
  INV_X1    g431(.A(new_n632), .ZN(new_n633));
  NAND2_X1  g432(.A1(new_n631), .A2(new_n633), .ZN(new_n634));
  OR2_X1    g433(.A1(new_n634), .A2(KEYINPUT97), .ZN(new_n635));
  INV_X1    g434(.A(KEYINPUT10), .ZN(new_n636));
  NAND3_X1  g435(.A1(new_n629), .A2(new_n630), .A3(new_n636), .ZN(new_n637));
  NAND3_X1  g436(.A1(new_n605), .A2(KEYINPUT10), .A3(new_n578), .ZN(new_n638));
  NAND2_X1  g437(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  NAND2_X1  g438(.A1(new_n639), .A2(new_n632), .ZN(new_n640));
  NAND2_X1  g439(.A1(new_n634), .A2(KEYINPUT97), .ZN(new_n641));
  NAND3_X1  g440(.A1(new_n635), .A2(new_n640), .A3(new_n641), .ZN(new_n642));
  XNOR2_X1  g441(.A(G120gat), .B(G148gat), .ZN(new_n643));
  XNOR2_X1  g442(.A(G176gat), .B(G204gat), .ZN(new_n644));
  XOR2_X1   g443(.A(new_n643), .B(new_n644), .Z(new_n645));
  INV_X1    g444(.A(new_n645), .ZN(new_n646));
  NAND2_X1  g445(.A1(new_n642), .A2(new_n646), .ZN(new_n647));
  NAND4_X1  g446(.A1(new_n635), .A2(new_n645), .A3(new_n640), .A4(new_n641), .ZN(new_n648));
  NAND2_X1  g447(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  NOR2_X1   g448(.A1(new_n627), .A2(new_n649), .ZN(new_n650));
  NAND2_X1  g449(.A1(new_n563), .A2(new_n650), .ZN(new_n651));
  NOR2_X1   g450(.A1(new_n651), .A2(new_n526), .ZN(new_n652));
  XNOR2_X1  g451(.A(new_n652), .B(new_n246), .ZN(G1324gat));
  NOR2_X1   g452(.A1(new_n651), .A2(new_n523), .ZN(new_n654));
  XOR2_X1   g453(.A(KEYINPUT16), .B(G8gat), .Z(new_n655));
  NAND2_X1  g454(.A1(new_n654), .A2(new_n655), .ZN(new_n656));
  INV_X1    g455(.A(G8gat), .ZN(new_n657));
  OAI21_X1  g456(.A(new_n656), .B1(new_n654), .B2(new_n657), .ZN(new_n658));
  MUX2_X1   g457(.A(new_n656), .B(new_n658), .S(KEYINPUT42), .Z(G1325gat));
  INV_X1    g458(.A(KEYINPUT98), .ZN(new_n660));
  OAI21_X1  g459(.A(new_n660), .B1(new_n559), .B2(new_n560), .ZN(new_n661));
  INV_X1    g460(.A(KEYINPUT36), .ZN(new_n662));
  NAND2_X1  g461(.A1(new_n461), .A2(new_n662), .ZN(new_n663));
  NAND3_X1  g462(.A1(new_n459), .A2(KEYINPUT36), .A3(new_n460), .ZN(new_n664));
  NAND3_X1  g463(.A1(new_n663), .A2(KEYINPUT98), .A3(new_n664), .ZN(new_n665));
  NAND2_X1  g464(.A1(new_n661), .A2(new_n665), .ZN(new_n666));
  OAI21_X1  g465(.A(G15gat), .B1(new_n651), .B2(new_n666), .ZN(new_n667));
  NAND2_X1  g466(.A1(new_n463), .A2(new_n464), .ZN(new_n668));
  INV_X1    g467(.A(new_n668), .ZN(new_n669));
  OR2_X1    g468(.A1(new_n669), .A2(G15gat), .ZN(new_n670));
  OAI21_X1  g469(.A(new_n667), .B1(new_n651), .B2(new_n670), .ZN(G1326gat));
  NOR2_X1   g470(.A1(new_n651), .A2(new_n520), .ZN(new_n672));
  XOR2_X1   g471(.A(KEYINPUT43), .B(G22gat), .Z(new_n673));
  XNOR2_X1  g472(.A(new_n672), .B(new_n673), .ZN(G1327gat));
  INV_X1    g473(.A(KEYINPUT44), .ZN(new_n675));
  AOI21_X1  g474(.A(new_n558), .B1(new_n661), .B2(new_n665), .ZN(new_n676));
  AND3_X1   g475(.A1(new_n443), .A2(KEYINPUT77), .A3(new_n447), .ZN(new_n677));
  AOI21_X1  g476(.A(KEYINPUT77), .B1(new_n443), .B2(new_n447), .ZN(new_n678));
  NOR3_X1   g477(.A1(new_n677), .A2(new_n678), .A3(new_n457), .ZN(new_n679));
  INV_X1    g478(.A(new_n460), .ZN(new_n680));
  OAI21_X1  g479(.A(new_n520), .B1(new_n679), .B2(new_n680), .ZN(new_n681));
  NAND2_X1  g480(.A1(new_n681), .A2(KEYINPUT85), .ZN(new_n682));
  INV_X1    g481(.A(new_n527), .ZN(new_n683));
  NAND3_X1  g482(.A1(new_n461), .A2(new_n519), .A3(new_n520), .ZN(new_n684));
  NAND3_X1  g483(.A1(new_n682), .A2(new_n683), .A3(new_n684), .ZN(new_n685));
  NAND2_X1  g484(.A1(new_n685), .A2(KEYINPUT35), .ZN(new_n686));
  AOI21_X1  g485(.A(new_n676), .B1(new_n686), .B2(new_n518), .ZN(new_n687));
  INV_X1    g486(.A(new_n625), .ZN(new_n688));
  OAI21_X1  g487(.A(new_n675), .B1(new_n687), .B2(new_n688), .ZN(new_n689));
  AOI22_X1  g488(.A1(new_n685), .A2(KEYINPUT35), .B1(new_n465), .B2(new_n517), .ZN(new_n690));
  OAI211_X1 g489(.A(KEYINPUT44), .B(new_n625), .C1(new_n690), .C2(new_n561), .ZN(new_n691));
  AND2_X1   g490(.A1(new_n689), .A2(new_n691), .ZN(new_n692));
  NOR2_X1   g491(.A1(new_n592), .A2(new_n649), .ZN(new_n693));
  AND2_X1   g492(.A1(new_n693), .A2(new_n295), .ZN(new_n694));
  NAND2_X1  g493(.A1(new_n692), .A2(new_n694), .ZN(new_n695));
  OAI21_X1  g494(.A(G29gat), .B1(new_n695), .B2(new_n526), .ZN(new_n696));
  NAND2_X1  g495(.A1(new_n693), .A2(new_n625), .ZN(new_n697));
  XOR2_X1   g496(.A(new_n697), .B(KEYINPUT99), .Z(new_n698));
  OAI211_X1 g497(.A(new_n295), .B(new_n698), .C1(new_n690), .C2(new_n561), .ZN(new_n699));
  INV_X1    g498(.A(new_n699), .ZN(new_n700));
  INV_X1    g499(.A(new_n526), .ZN(new_n701));
  NAND3_X1  g500(.A1(new_n700), .A2(new_n236), .A3(new_n701), .ZN(new_n702));
  XNOR2_X1  g501(.A(new_n702), .B(KEYINPUT45), .ZN(new_n703));
  NAND2_X1  g502(.A1(new_n696), .A2(new_n703), .ZN(G1328gat));
  NAND3_X1  g503(.A1(new_n700), .A2(new_n222), .A3(new_n484), .ZN(new_n705));
  AND2_X1   g504(.A1(KEYINPUT100), .A2(KEYINPUT46), .ZN(new_n706));
  NOR2_X1   g505(.A1(KEYINPUT100), .A2(KEYINPUT46), .ZN(new_n707));
  OAI21_X1  g506(.A(new_n705), .B1(new_n706), .B2(new_n707), .ZN(new_n708));
  OAI21_X1  g507(.A(KEYINPUT101), .B1(new_n695), .B2(new_n523), .ZN(new_n709));
  NAND2_X1  g508(.A1(new_n709), .A2(G36gat), .ZN(new_n710));
  NOR3_X1   g509(.A1(new_n695), .A2(KEYINPUT101), .A3(new_n523), .ZN(new_n711));
  OAI221_X1 g510(.A(new_n708), .B1(new_n706), .B2(new_n705), .C1(new_n710), .C2(new_n711), .ZN(G1329gat));
  INV_X1    g511(.A(new_n666), .ZN(new_n713));
  NAND4_X1  g512(.A1(new_n689), .A2(new_n713), .A3(new_n691), .A4(new_n694), .ZN(new_n714));
  NAND2_X1  g513(.A1(new_n714), .A2(G43gat), .ZN(new_n715));
  INV_X1    g514(.A(KEYINPUT103), .ZN(new_n716));
  NOR2_X1   g515(.A1(new_n669), .A2(G43gat), .ZN(new_n717));
  INV_X1    g516(.A(new_n717), .ZN(new_n718));
  OAI21_X1  g517(.A(new_n716), .B1(new_n699), .B2(new_n718), .ZN(new_n719));
  NAND4_X1  g518(.A1(new_n563), .A2(KEYINPUT103), .A3(new_n698), .A4(new_n717), .ZN(new_n720));
  AND2_X1   g519(.A1(new_n719), .A2(new_n720), .ZN(new_n721));
  AOI21_X1  g520(.A(KEYINPUT102), .B1(new_n715), .B2(new_n721), .ZN(new_n722));
  INV_X1    g521(.A(KEYINPUT104), .ZN(new_n723));
  NOR3_X1   g522(.A1(new_n722), .A2(new_n723), .A3(KEYINPUT47), .ZN(new_n724));
  OR2_X1    g523(.A1(new_n722), .A2(new_n723), .ZN(new_n725));
  INV_X1    g524(.A(KEYINPUT47), .ZN(new_n726));
  NAND2_X1  g525(.A1(new_n715), .A2(new_n721), .ZN(new_n727));
  AOI21_X1  g526(.A(new_n726), .B1(new_n727), .B2(new_n723), .ZN(new_n728));
  AOI21_X1  g527(.A(new_n724), .B1(new_n725), .B2(new_n728), .ZN(G1330gat));
  OAI21_X1  g528(.A(new_n209), .B1(new_n699), .B2(new_n520), .ZN(new_n730));
  NAND2_X1  g529(.A1(new_n355), .A2(G50gat), .ZN(new_n731));
  OAI21_X1  g530(.A(new_n730), .B1(new_n695), .B2(new_n731), .ZN(new_n732));
  XNOR2_X1  g531(.A(new_n732), .B(KEYINPUT48), .ZN(G1331gat));
  INV_X1    g532(.A(new_n649), .ZN(new_n734));
  NOR4_X1   g533(.A1(new_n687), .A2(new_n295), .A3(new_n627), .A4(new_n734), .ZN(new_n735));
  XOR2_X1   g534(.A(new_n526), .B(KEYINPUT105), .Z(new_n736));
  NAND2_X1  g535(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  XNOR2_X1  g536(.A(new_n737), .B(G57gat), .ZN(G1332gat));
  NAND2_X1  g537(.A1(new_n735), .A2(new_n484), .ZN(new_n739));
  OAI21_X1  g538(.A(new_n739), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n740));
  XOR2_X1   g539(.A(KEYINPUT49), .B(G64gat), .Z(new_n741));
  OAI21_X1  g540(.A(new_n740), .B1(new_n739), .B2(new_n741), .ZN(G1333gat));
  NAND2_X1  g541(.A1(new_n735), .A2(new_n668), .ZN(new_n743));
  NAND2_X1  g542(.A1(new_n743), .A2(new_n565), .ZN(new_n744));
  NAND3_X1  g543(.A1(new_n735), .A2(G71gat), .A3(new_n713), .ZN(new_n745));
  INV_X1    g544(.A(KEYINPUT106), .ZN(new_n746));
  AND2_X1   g545(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  NOR2_X1   g546(.A1(new_n745), .A2(new_n746), .ZN(new_n748));
  OAI21_X1  g547(.A(new_n744), .B1(new_n747), .B2(new_n748), .ZN(new_n749));
  NAND2_X1  g548(.A1(new_n749), .A2(KEYINPUT50), .ZN(new_n750));
  INV_X1    g549(.A(KEYINPUT50), .ZN(new_n751));
  OAI211_X1 g550(.A(new_n751), .B(new_n744), .C1(new_n747), .C2(new_n748), .ZN(new_n752));
  NAND2_X1  g551(.A1(new_n750), .A2(new_n752), .ZN(G1334gat));
  NAND2_X1  g552(.A1(new_n735), .A2(new_n355), .ZN(new_n754));
  XNOR2_X1  g553(.A(new_n754), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g554(.A1(new_n295), .A2(new_n592), .ZN(new_n756));
  NAND2_X1  g555(.A1(new_n756), .A2(new_n649), .ZN(new_n757));
  XOR2_X1   g556(.A(new_n757), .B(KEYINPUT107), .Z(new_n758));
  NAND2_X1  g557(.A1(new_n692), .A2(new_n758), .ZN(new_n759));
  OAI21_X1  g558(.A(G85gat), .B1(new_n759), .B2(new_n526), .ZN(new_n760));
  OAI211_X1 g559(.A(new_n625), .B(new_n756), .C1(new_n690), .C2(new_n676), .ZN(new_n761));
  INV_X1    g560(.A(KEYINPUT51), .ZN(new_n762));
  XNOR2_X1  g561(.A(new_n761), .B(new_n762), .ZN(new_n763));
  NAND4_X1  g562(.A1(new_n763), .A2(new_n599), .A3(new_n701), .A4(new_n649), .ZN(new_n764));
  NAND2_X1  g563(.A1(new_n760), .A2(new_n764), .ZN(G1336gat));
  OAI21_X1  g564(.A(G92gat), .B1(new_n759), .B2(new_n523), .ZN(new_n766));
  NAND4_X1  g565(.A1(new_n763), .A2(new_n600), .A3(new_n484), .A4(new_n649), .ZN(new_n767));
  NAND2_X1  g566(.A1(new_n766), .A2(new_n767), .ZN(new_n768));
  NAND2_X1  g567(.A1(new_n768), .A2(KEYINPUT52), .ZN(new_n769));
  INV_X1    g568(.A(KEYINPUT52), .ZN(new_n770));
  NAND3_X1  g569(.A1(new_n766), .A2(new_n770), .A3(new_n767), .ZN(new_n771));
  NAND2_X1  g570(.A1(new_n769), .A2(new_n771), .ZN(G1337gat));
  XNOR2_X1  g571(.A(KEYINPUT108), .B(G99gat), .ZN(new_n773));
  NAND4_X1  g572(.A1(new_n763), .A2(new_n668), .A3(new_n649), .A4(new_n773), .ZN(new_n774));
  NOR2_X1   g573(.A1(new_n759), .A2(new_n666), .ZN(new_n775));
  OAI21_X1  g574(.A(new_n774), .B1(new_n775), .B2(new_n773), .ZN(G1338gat));
  INV_X1    g575(.A(KEYINPUT111), .ZN(new_n777));
  NOR3_X1   g576(.A1(new_n520), .A2(G106gat), .A3(new_n734), .ZN(new_n778));
  XOR2_X1   g577(.A(new_n778), .B(KEYINPUT110), .Z(new_n779));
  AND3_X1   g578(.A1(new_n763), .A2(new_n777), .A3(new_n779), .ZN(new_n780));
  AOI21_X1  g579(.A(new_n777), .B1(new_n763), .B2(new_n779), .ZN(new_n781));
  NAND4_X1  g580(.A1(new_n689), .A2(new_n355), .A3(new_n691), .A4(new_n758), .ZN(new_n782));
  XOR2_X1   g581(.A(KEYINPUT109), .B(G106gat), .Z(new_n783));
  INV_X1    g582(.A(new_n783), .ZN(new_n784));
  AND2_X1   g583(.A1(new_n782), .A2(new_n784), .ZN(new_n785));
  NOR3_X1   g584(.A1(new_n780), .A2(new_n781), .A3(new_n785), .ZN(new_n786));
  INV_X1    g585(.A(KEYINPUT53), .ZN(new_n787));
  NAND2_X1  g586(.A1(new_n763), .A2(new_n778), .ZN(new_n788));
  INV_X1    g587(.A(KEYINPUT112), .ZN(new_n789));
  NAND2_X1  g588(.A1(new_n788), .A2(new_n789), .ZN(new_n790));
  NAND3_X1  g589(.A1(new_n763), .A2(KEYINPUT112), .A3(new_n778), .ZN(new_n791));
  NAND3_X1  g590(.A1(new_n790), .A2(new_n787), .A3(new_n791), .ZN(new_n792));
  OR2_X1    g591(.A1(new_n782), .A2(KEYINPUT113), .ZN(new_n793));
  NAND2_X1  g592(.A1(new_n782), .A2(KEYINPUT113), .ZN(new_n794));
  AOI21_X1  g593(.A(new_n783), .B1(new_n793), .B2(new_n794), .ZN(new_n795));
  OAI22_X1  g594(.A1(new_n786), .A2(new_n787), .B1(new_n792), .B2(new_n795), .ZN(G1339gat));
  NOR3_X1   g595(.A1(new_n627), .A2(new_n295), .A3(new_n649), .ZN(new_n797));
  INV_X1    g596(.A(KEYINPUT114), .ZN(new_n798));
  AOI21_X1  g597(.A(new_n259), .B1(new_n287), .B2(new_n258), .ZN(new_n799));
  NOR2_X1   g598(.A1(new_n276), .A2(new_n277), .ZN(new_n800));
  OAI21_X1  g599(.A(new_n205), .B1(new_n799), .B2(new_n800), .ZN(new_n801));
  AND3_X1   g600(.A1(new_n294), .A2(new_n801), .A3(new_n649), .ZN(new_n802));
  NAND3_X1  g601(.A1(new_n637), .A2(new_n633), .A3(new_n638), .ZN(new_n803));
  NAND3_X1  g602(.A1(new_n640), .A2(KEYINPUT54), .A3(new_n803), .ZN(new_n804));
  AOI21_X1  g603(.A(new_n633), .B1(new_n637), .B2(new_n638), .ZN(new_n805));
  INV_X1    g604(.A(KEYINPUT54), .ZN(new_n806));
  AOI21_X1  g605(.A(new_n645), .B1(new_n805), .B2(new_n806), .ZN(new_n807));
  NAND3_X1  g606(.A1(new_n804), .A2(KEYINPUT55), .A3(new_n807), .ZN(new_n808));
  NAND2_X1  g607(.A1(new_n808), .A2(new_n648), .ZN(new_n809));
  AOI21_X1  g608(.A(KEYINPUT55), .B1(new_n804), .B2(new_n807), .ZN(new_n810));
  OR2_X1    g609(.A1(new_n809), .A2(new_n810), .ZN(new_n811));
  AOI21_X1  g610(.A(new_n811), .B1(new_n290), .B2(new_n294), .ZN(new_n812));
  OAI21_X1  g611(.A(new_n798), .B1(new_n802), .B2(new_n812), .ZN(new_n813));
  NOR2_X1   g612(.A1(new_n809), .A2(new_n810), .ZN(new_n814));
  AND3_X1   g613(.A1(new_n291), .A2(new_n293), .A3(new_n206), .ZN(new_n815));
  INV_X1    g614(.A(new_n207), .ZN(new_n816));
  AOI21_X1  g615(.A(new_n816), .B1(new_n291), .B2(new_n293), .ZN(new_n817));
  OAI21_X1  g616(.A(new_n814), .B1(new_n815), .B2(new_n817), .ZN(new_n818));
  NAND3_X1  g617(.A1(new_n294), .A2(new_n801), .A3(new_n649), .ZN(new_n819));
  NAND3_X1  g618(.A1(new_n818), .A2(KEYINPUT114), .A3(new_n819), .ZN(new_n820));
  NAND3_X1  g619(.A1(new_n813), .A2(new_n820), .A3(new_n688), .ZN(new_n821));
  NAND4_X1  g620(.A1(new_n625), .A2(new_n294), .A3(new_n801), .A4(new_n814), .ZN(new_n822));
  NAND2_X1  g621(.A1(new_n821), .A2(new_n822), .ZN(new_n823));
  AOI21_X1  g622(.A(new_n797), .B1(new_n823), .B2(new_n593), .ZN(new_n824));
  NOR3_X1   g623(.A1(new_n824), .A2(new_n355), .A3(new_n669), .ZN(new_n825));
  NOR2_X1   g624(.A1(new_n484), .A2(new_n526), .ZN(new_n826));
  NAND2_X1  g625(.A1(new_n825), .A2(new_n826), .ZN(new_n827));
  OAI21_X1  g626(.A(G113gat), .B1(new_n827), .B2(new_n296), .ZN(new_n828));
  INV_X1    g627(.A(new_n824), .ZN(new_n829));
  AND2_X1   g628(.A1(new_n829), .A2(new_n736), .ZN(new_n830));
  NAND4_X1  g629(.A1(new_n830), .A2(new_n523), .A3(new_n682), .A4(new_n684), .ZN(new_n831));
  OR2_X1    g630(.A1(new_n296), .A2(G113gat), .ZN(new_n832));
  OAI21_X1  g631(.A(new_n828), .B1(new_n831), .B2(new_n832), .ZN(new_n833));
  XNOR2_X1  g632(.A(new_n833), .B(KEYINPUT115), .ZN(G1340gat));
  OAI21_X1  g633(.A(G120gat), .B1(new_n827), .B2(new_n734), .ZN(new_n835));
  NOR2_X1   g634(.A1(new_n734), .A2(G120gat), .ZN(new_n836));
  XNOR2_X1  g635(.A(new_n836), .B(KEYINPUT116), .ZN(new_n837));
  OAI21_X1  g636(.A(new_n835), .B1(new_n831), .B2(new_n837), .ZN(G1341gat));
  OAI21_X1  g637(.A(G127gat), .B1(new_n827), .B2(new_n593), .ZN(new_n839));
  OR2_X1    g638(.A1(new_n593), .A2(G127gat), .ZN(new_n840));
  OAI21_X1  g639(.A(new_n839), .B1(new_n831), .B2(new_n840), .ZN(G1342gat));
  OR3_X1    g640(.A1(new_n831), .A2(G134gat), .A3(new_n688), .ZN(new_n842));
  OR2_X1    g641(.A1(new_n842), .A2(KEYINPUT56), .ZN(new_n843));
  OAI21_X1  g642(.A(G134gat), .B1(new_n827), .B2(new_n688), .ZN(new_n844));
  NAND2_X1  g643(.A1(new_n842), .A2(KEYINPUT56), .ZN(new_n845));
  NAND3_X1  g644(.A1(new_n843), .A2(new_n844), .A3(new_n845), .ZN(G1343gat));
  NAND2_X1  g645(.A1(new_n666), .A2(new_n826), .ZN(new_n847));
  INV_X1    g646(.A(new_n847), .ZN(new_n848));
  AOI21_X1  g647(.A(KEYINPUT57), .B1(new_n829), .B2(new_n355), .ZN(new_n849));
  AOI21_X1  g648(.A(KEYINPUT117), .B1(new_n804), .B2(new_n807), .ZN(new_n850));
  NOR2_X1   g649(.A1(new_n850), .A2(KEYINPUT55), .ZN(new_n851));
  NAND3_X1  g650(.A1(new_n804), .A2(KEYINPUT117), .A3(new_n807), .ZN(new_n852));
  AOI21_X1  g651(.A(new_n809), .B1(new_n851), .B2(new_n852), .ZN(new_n853));
  NAND2_X1  g652(.A1(new_n295), .A2(new_n853), .ZN(new_n854));
  AOI21_X1  g653(.A(new_n625), .B1(new_n854), .B2(new_n819), .ZN(new_n855));
  INV_X1    g654(.A(new_n855), .ZN(new_n856));
  NAND2_X1  g655(.A1(new_n856), .A2(new_n822), .ZN(new_n857));
  AOI21_X1  g656(.A(new_n797), .B1(new_n857), .B2(new_n593), .ZN(new_n858));
  INV_X1    g657(.A(KEYINPUT57), .ZN(new_n859));
  NOR3_X1   g658(.A1(new_n858), .A2(new_n859), .A3(new_n520), .ZN(new_n860));
  OAI21_X1  g659(.A(new_n848), .B1(new_n849), .B2(new_n860), .ZN(new_n861));
  OAI21_X1  g660(.A(G141gat), .B1(new_n861), .B2(new_n296), .ZN(new_n862));
  NAND2_X1  g661(.A1(new_n829), .A2(new_n736), .ZN(new_n863));
  NAND2_X1  g662(.A1(new_n666), .A2(new_n355), .ZN(new_n864));
  NOR3_X1   g663(.A1(new_n863), .A2(new_n484), .A3(new_n864), .ZN(new_n865));
  NOR2_X1   g664(.A1(new_n296), .A2(G141gat), .ZN(new_n866));
  AOI21_X1  g665(.A(KEYINPUT58), .B1(new_n865), .B2(new_n866), .ZN(new_n867));
  NAND2_X1  g666(.A1(new_n862), .A2(new_n867), .ZN(new_n868));
  NAND2_X1  g667(.A1(new_n861), .A2(KEYINPUT118), .ZN(new_n869));
  INV_X1    g668(.A(KEYINPUT118), .ZN(new_n870));
  OAI211_X1 g669(.A(new_n870), .B(new_n848), .C1(new_n849), .C2(new_n860), .ZN(new_n871));
  NAND3_X1  g670(.A1(new_n869), .A2(new_n295), .A3(new_n871), .ZN(new_n872));
  AOI22_X1  g671(.A1(new_n872), .A2(G141gat), .B1(new_n865), .B2(new_n866), .ZN(new_n873));
  INV_X1    g672(.A(KEYINPUT58), .ZN(new_n874));
  OAI21_X1  g673(.A(new_n868), .B1(new_n873), .B2(new_n874), .ZN(G1344gat));
  NAND3_X1  g674(.A1(new_n869), .A2(new_n649), .A3(new_n871), .ZN(new_n876));
  INV_X1    g675(.A(KEYINPUT59), .ZN(new_n877));
  NAND3_X1  g676(.A1(new_n876), .A2(new_n877), .A3(G148gat), .ZN(new_n878));
  INV_X1    g677(.A(G148gat), .ZN(new_n879));
  NOR2_X1   g678(.A1(new_n520), .A2(new_n859), .ZN(new_n880));
  AOI21_X1  g679(.A(new_n592), .B1(new_n821), .B2(new_n822), .ZN(new_n881));
  OAI21_X1  g680(.A(new_n880), .B1(new_n881), .B2(new_n797), .ZN(new_n882));
  INV_X1    g681(.A(KEYINPUT119), .ZN(new_n883));
  NAND2_X1  g682(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  OAI211_X1 g683(.A(KEYINPUT119), .B(new_n880), .C1(new_n881), .C2(new_n797), .ZN(new_n885));
  INV_X1    g684(.A(new_n797), .ZN(new_n886));
  NAND2_X1  g685(.A1(new_n623), .A2(new_n619), .ZN(new_n887));
  NAND2_X1  g686(.A1(new_n615), .A2(new_n616), .ZN(new_n888));
  NAND2_X1  g687(.A1(new_n887), .A2(new_n888), .ZN(new_n889));
  INV_X1    g688(.A(KEYINPUT120), .ZN(new_n890));
  NAND4_X1  g689(.A1(new_n889), .A2(new_n814), .A3(new_n890), .A4(new_n620), .ZN(new_n891));
  NAND3_X1  g690(.A1(new_n891), .A2(new_n294), .A3(new_n801), .ZN(new_n892));
  AOI21_X1  g691(.A(new_n890), .B1(new_n625), .B2(new_n814), .ZN(new_n893));
  NOR2_X1   g692(.A1(new_n892), .A2(new_n893), .ZN(new_n894));
  OAI21_X1  g693(.A(new_n593), .B1(new_n855), .B2(new_n894), .ZN(new_n895));
  NAND2_X1  g694(.A1(new_n886), .A2(new_n895), .ZN(new_n896));
  NAND2_X1  g695(.A1(new_n896), .A2(new_n355), .ZN(new_n897));
  NAND2_X1  g696(.A1(new_n897), .A2(new_n859), .ZN(new_n898));
  NAND3_X1  g697(.A1(new_n884), .A2(new_n885), .A3(new_n898), .ZN(new_n899));
  NOR2_X1   g698(.A1(new_n847), .A2(new_n734), .ZN(new_n900));
  AOI21_X1  g699(.A(new_n879), .B1(new_n899), .B2(new_n900), .ZN(new_n901));
  NOR2_X1   g700(.A1(new_n901), .A2(new_n877), .ZN(new_n902));
  NOR2_X1   g701(.A1(new_n902), .A2(KEYINPUT121), .ZN(new_n903));
  INV_X1    g702(.A(KEYINPUT121), .ZN(new_n904));
  NOR3_X1   g703(.A1(new_n901), .A2(new_n904), .A3(new_n877), .ZN(new_n905));
  OAI21_X1  g704(.A(new_n878), .B1(new_n903), .B2(new_n905), .ZN(new_n906));
  NAND3_X1  g705(.A1(new_n865), .A2(new_n879), .A3(new_n649), .ZN(new_n907));
  NAND2_X1  g706(.A1(new_n906), .A2(new_n907), .ZN(G1345gat));
  NAND3_X1  g707(.A1(new_n865), .A2(new_n298), .A3(new_n592), .ZN(new_n909));
  AND3_X1   g708(.A1(new_n869), .A2(new_n592), .A3(new_n871), .ZN(new_n910));
  OAI21_X1  g709(.A(new_n909), .B1(new_n910), .B2(new_n298), .ZN(G1346gat));
  NAND3_X1  g710(.A1(new_n865), .A2(new_n299), .A3(new_n625), .ZN(new_n912));
  XNOR2_X1  g711(.A(new_n912), .B(KEYINPUT122), .ZN(new_n913));
  AND3_X1   g712(.A1(new_n869), .A2(new_n625), .A3(new_n871), .ZN(new_n914));
  OAI21_X1  g713(.A(new_n913), .B1(new_n299), .B2(new_n914), .ZN(G1347gat));
  NOR2_X1   g714(.A1(new_n736), .A2(new_n523), .ZN(new_n916));
  NAND2_X1  g715(.A1(new_n825), .A2(new_n916), .ZN(new_n917));
  OAI21_X1  g716(.A(G169gat), .B1(new_n917), .B2(new_n296), .ZN(new_n918));
  NOR2_X1   g717(.A1(new_n824), .A2(new_n701), .ZN(new_n919));
  NOR3_X1   g718(.A1(new_n521), .A2(new_n522), .A3(new_n523), .ZN(new_n920));
  NAND2_X1  g719(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  XOR2_X1   g720(.A(new_n921), .B(KEYINPUT123), .Z(new_n922));
  NAND2_X1  g721(.A1(new_n295), .A2(new_n411), .ZN(new_n923));
  OAI21_X1  g722(.A(new_n918), .B1(new_n922), .B2(new_n923), .ZN(G1348gat));
  OAI21_X1  g723(.A(G176gat), .B1(new_n917), .B2(new_n734), .ZN(new_n925));
  OR2_X1    g724(.A1(new_n734), .A2(G176gat), .ZN(new_n926));
  OAI21_X1  g725(.A(new_n925), .B1(new_n922), .B2(new_n926), .ZN(G1349gat));
  NOR3_X1   g726(.A1(new_n921), .A2(new_n401), .A3(new_n593), .ZN(new_n928));
  INV_X1    g727(.A(KEYINPUT124), .ZN(new_n929));
  XNOR2_X1  g728(.A(new_n928), .B(new_n929), .ZN(new_n930));
  OAI21_X1  g729(.A(new_n385), .B1(new_n917), .B2(new_n593), .ZN(new_n931));
  NAND2_X1  g730(.A1(new_n930), .A2(new_n931), .ZN(new_n932));
  NAND2_X1  g731(.A1(new_n932), .A2(KEYINPUT60), .ZN(new_n933));
  INV_X1    g732(.A(KEYINPUT60), .ZN(new_n934));
  NAND3_X1  g733(.A1(new_n930), .A2(new_n934), .A3(new_n931), .ZN(new_n935));
  NAND2_X1  g734(.A1(new_n933), .A2(new_n935), .ZN(G1350gat));
  OAI21_X1  g735(.A(G190gat), .B1(new_n917), .B2(new_n688), .ZN(new_n937));
  XNOR2_X1  g736(.A(new_n937), .B(KEYINPUT61), .ZN(new_n938));
  NAND2_X1  g737(.A1(new_n625), .A2(new_n399), .ZN(new_n939));
  OAI21_X1  g738(.A(new_n938), .B1(new_n922), .B2(new_n939), .ZN(G1351gat));
  NOR2_X1   g739(.A1(new_n864), .A2(new_n523), .ZN(new_n941));
  NAND2_X1  g740(.A1(new_n919), .A2(new_n941), .ZN(new_n942));
  INV_X1    g741(.A(new_n942), .ZN(new_n943));
  AOI21_X1  g742(.A(G197gat), .B1(new_n943), .B2(new_n295), .ZN(new_n944));
  NAND2_X1  g743(.A1(new_n666), .A2(new_n916), .ZN(new_n945));
  AOI22_X1  g744(.A1(new_n882), .A2(new_n883), .B1(new_n897), .B2(new_n859), .ZN(new_n946));
  AOI21_X1  g745(.A(new_n945), .B1(new_n946), .B2(new_n885), .ZN(new_n947));
  AND2_X1   g746(.A1(new_n295), .A2(G197gat), .ZN(new_n948));
  AOI21_X1  g747(.A(new_n944), .B1(new_n947), .B2(new_n948), .ZN(G1352gat));
  NOR3_X1   g748(.A1(new_n942), .A2(G204gat), .A3(new_n734), .ZN(new_n950));
  XNOR2_X1  g749(.A(new_n950), .B(KEYINPUT62), .ZN(new_n951));
  INV_X1    g750(.A(new_n945), .ZN(new_n952));
  NAND2_X1  g751(.A1(new_n899), .A2(new_n952), .ZN(new_n953));
  OAI21_X1  g752(.A(G204gat), .B1(new_n953), .B2(new_n734), .ZN(new_n954));
  NAND2_X1  g753(.A1(new_n951), .A2(new_n954), .ZN(G1353gat));
  NAND3_X1  g754(.A1(new_n943), .A2(new_n309), .A3(new_n592), .ZN(new_n956));
  OAI21_X1  g755(.A(G211gat), .B1(KEYINPUT125), .B2(KEYINPUT63), .ZN(new_n957));
  NAND2_X1  g756(.A1(KEYINPUT125), .A2(KEYINPUT63), .ZN(new_n958));
  AOI211_X1 g757(.A(new_n957), .B(new_n958), .C1(new_n947), .C2(new_n592), .ZN(new_n959));
  NAND3_X1  g758(.A1(new_n899), .A2(new_n592), .A3(new_n952), .ZN(new_n960));
  INV_X1    g759(.A(new_n957), .ZN(new_n961));
  AOI22_X1  g760(.A1(new_n960), .A2(new_n961), .B1(KEYINPUT125), .B2(KEYINPUT63), .ZN(new_n962));
  OAI21_X1  g761(.A(new_n956), .B1(new_n959), .B2(new_n962), .ZN(new_n963));
  NAND2_X1  g762(.A1(new_n963), .A2(KEYINPUT126), .ZN(new_n964));
  INV_X1    g763(.A(KEYINPUT126), .ZN(new_n965));
  OAI211_X1 g764(.A(new_n965), .B(new_n956), .C1(new_n959), .C2(new_n962), .ZN(new_n966));
  NAND2_X1  g765(.A1(new_n964), .A2(new_n966), .ZN(G1354gat));
  OAI21_X1  g766(.A(G218gat), .B1(new_n953), .B2(new_n688), .ZN(new_n968));
  NAND2_X1  g767(.A1(new_n625), .A2(new_n310), .ZN(new_n969));
  OAI21_X1  g768(.A(new_n968), .B1(new_n942), .B2(new_n969), .ZN(new_n970));
  INV_X1    g769(.A(KEYINPUT127), .ZN(new_n971));
  XNOR2_X1  g770(.A(new_n970), .B(new_n971), .ZN(G1355gat));
endmodule


