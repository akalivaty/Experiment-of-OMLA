//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 1 1 1 1 0 1 1 0 1 0 0 1 0 1 1 1 0 0 0 0 0 1 1 1 0 0 0 1 0 0 1 0 1 0 1 1 0 0 0 0 0 1 1 1 0 0 0 1 0 1 0 1 0 1 0 1 0 1 0 0 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:34:34 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n447, new_n451, new_n452, new_n453, new_n454, new_n455,
    new_n458, new_n459, new_n460, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n483, new_n484, new_n485, new_n486,
    new_n487, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n532, new_n533, new_n534, new_n535, new_n536, new_n537, new_n538,
    new_n539, new_n540, new_n541, new_n544, new_n545, new_n546, new_n547,
    new_n548, new_n549, new_n550, new_n551, new_n552, new_n553, new_n554,
    new_n555, new_n556, new_n557, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n567, new_n568, new_n569, new_n570, new_n573,
    new_n574, new_n576, new_n577, new_n578, new_n579, new_n580, new_n581,
    new_n582, new_n583, new_n584, new_n585, new_n586, new_n587, new_n588,
    new_n589, new_n590, new_n591, new_n592, new_n593, new_n594, new_n595,
    new_n596, new_n597, new_n600, new_n601, new_n602, new_n603, new_n605,
    new_n606, new_n607, new_n608, new_n609, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n638, new_n641, new_n643, new_n644, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n677, new_n678,
    new_n679, new_n680, new_n681, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n692, new_n693,
    new_n694, new_n695, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n713, new_n714, new_n715,
    new_n716, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n851, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1194, new_n1195;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  XNOR2_X1  g007(.A(KEYINPUT64), .B(G2066), .ZN(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(new_n436));
  XNOR2_X1  g011(.A(new_n436), .B(KEYINPUT65), .ZN(G220));
  XOR2_X1   g012(.A(KEYINPUT66), .B(G96), .Z(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  INV_X1    g015(.A(G57), .ZN(G237));
  XOR2_X1   g016(.A(KEYINPUT67), .B(G108), .Z(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g025(.A1(G220), .A2(G218), .A3(G219), .A4(G221), .ZN(new_n451));
  XNOR2_X1  g026(.A(new_n451), .B(KEYINPUT2), .ZN(new_n452));
  INV_X1    g027(.A(new_n452), .ZN(new_n453));
  NOR4_X1   g028(.A1(G238), .A2(G237), .A3(G235), .A4(G236), .ZN(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(new_n455));
  NOR2_X1   g030(.A1(new_n453), .A2(new_n455), .ZN(G325));
  INV_X1    g031(.A(G325), .ZN(G261));
  NAND2_X1  g032(.A1(new_n453), .A2(G2106), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n455), .A2(G567), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  INV_X1    g035(.A(new_n460), .ZN(G319));
  AND2_X1   g036(.A1(KEYINPUT68), .A2(G2105), .ZN(new_n462));
  NOR2_X1   g037(.A1(KEYINPUT68), .A2(G2105), .ZN(new_n463));
  NOR2_X1   g038(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  XNOR2_X1  g039(.A(KEYINPUT3), .B(G2104), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n465), .A2(G125), .ZN(new_n466));
  NAND2_X1  g041(.A1(G113), .A2(G2104), .ZN(new_n467));
  AOI21_X1  g042(.A(new_n464), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  INV_X1    g043(.A(KEYINPUT69), .ZN(new_n469));
  INV_X1    g044(.A(G2104), .ZN(new_n470));
  NOR2_X1   g045(.A1(new_n470), .A2(G2105), .ZN(new_n471));
  AOI21_X1  g046(.A(new_n469), .B1(new_n471), .B2(G101), .ZN(new_n472));
  INV_X1    g047(.A(G2105), .ZN(new_n473));
  NAND4_X1  g048(.A1(new_n469), .A2(new_n473), .A3(G101), .A4(G2104), .ZN(new_n474));
  INV_X1    g049(.A(new_n474), .ZN(new_n475));
  AND2_X1   g050(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n476));
  NOR2_X1   g051(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n477));
  OAI21_X1  g052(.A(G137), .B1(new_n476), .B2(new_n477), .ZN(new_n478));
  XNOR2_X1  g053(.A(KEYINPUT68), .B(G2105), .ZN(new_n479));
  OAI22_X1  g054(.A1(new_n472), .A2(new_n475), .B1(new_n478), .B2(new_n479), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n480), .A2(KEYINPUT70), .ZN(new_n481));
  NAND3_X1  g056(.A1(new_n464), .A2(new_n465), .A3(G137), .ZN(new_n482));
  NAND3_X1  g057(.A1(new_n473), .A2(G101), .A3(G2104), .ZN(new_n483));
  NAND2_X1  g058(.A1(new_n483), .A2(KEYINPUT69), .ZN(new_n484));
  NAND2_X1  g059(.A1(new_n484), .A2(new_n474), .ZN(new_n485));
  INV_X1    g060(.A(KEYINPUT70), .ZN(new_n486));
  NAND3_X1  g061(.A1(new_n482), .A2(new_n485), .A3(new_n486), .ZN(new_n487));
  AOI21_X1  g062(.A(new_n468), .B1(new_n481), .B2(new_n487), .ZN(G160));
  NOR2_X1   g063(.A1(new_n476), .A2(new_n477), .ZN(new_n489));
  NOR2_X1   g064(.A1(new_n489), .A2(new_n464), .ZN(new_n490));
  NAND2_X1  g065(.A1(new_n490), .A2(G124), .ZN(new_n491));
  NOR2_X1   g066(.A1(new_n464), .A2(G112), .ZN(new_n492));
  OAI21_X1  g067(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n493));
  OAI21_X1  g068(.A(new_n491), .B1(new_n492), .B2(new_n493), .ZN(new_n494));
  NOR2_X1   g069(.A1(new_n489), .A2(G2105), .ZN(new_n495));
  INV_X1    g070(.A(new_n495), .ZN(new_n496));
  INV_X1    g071(.A(G136), .ZN(new_n497));
  OR3_X1    g072(.A1(new_n496), .A2(KEYINPUT71), .A3(new_n497), .ZN(new_n498));
  OAI21_X1  g073(.A(KEYINPUT71), .B1(new_n496), .B2(new_n497), .ZN(new_n499));
  AOI21_X1  g074(.A(new_n494), .B1(new_n498), .B2(new_n499), .ZN(G162));
  AND3_X1   g075(.A1(new_n473), .A2(G102), .A3(G2104), .ZN(new_n501));
  INV_X1    g076(.A(KEYINPUT4), .ZN(new_n502));
  NOR3_X1   g077(.A1(new_n462), .A2(new_n463), .A3(new_n502), .ZN(new_n503));
  INV_X1    g078(.A(G138), .ZN(new_n504));
  INV_X1    g079(.A(KEYINPUT3), .ZN(new_n505));
  NAND2_X1  g080(.A1(new_n505), .A2(new_n470), .ZN(new_n506));
  NAND2_X1  g081(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n507));
  AOI21_X1  g082(.A(new_n504), .B1(new_n506), .B2(new_n507), .ZN(new_n508));
  AOI21_X1  g083(.A(new_n501), .B1(new_n503), .B2(new_n508), .ZN(new_n509));
  INV_X1    g084(.A(G126), .ZN(new_n510));
  AOI21_X1  g085(.A(new_n510), .B1(new_n506), .B2(new_n507), .ZN(new_n511));
  AND2_X1   g086(.A1(G114), .A2(G2104), .ZN(new_n512));
  OAI21_X1  g087(.A(G2105), .B1(new_n511), .B2(new_n512), .ZN(new_n513));
  OAI21_X1  g088(.A(G138), .B1(new_n476), .B2(new_n477), .ZN(new_n514));
  OAI21_X1  g089(.A(new_n502), .B1(new_n514), .B2(new_n479), .ZN(new_n515));
  NAND3_X1  g090(.A1(new_n509), .A2(new_n513), .A3(new_n515), .ZN(new_n516));
  INV_X1    g091(.A(new_n516), .ZN(G164));
  NOR2_X1   g092(.A1(KEYINPUT6), .A2(G651), .ZN(new_n518));
  XNOR2_X1  g093(.A(KEYINPUT72), .B(G651), .ZN(new_n519));
  AOI21_X1  g094(.A(new_n518), .B1(new_n519), .B2(KEYINPUT6), .ZN(new_n520));
  INV_X1    g095(.A(KEYINPUT5), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n521), .A2(G543), .ZN(new_n522));
  INV_X1    g097(.A(G543), .ZN(new_n523));
  AND3_X1   g098(.A1(new_n523), .A2(KEYINPUT73), .A3(KEYINPUT5), .ZN(new_n524));
  AOI21_X1  g099(.A(KEYINPUT73), .B1(new_n523), .B2(KEYINPUT5), .ZN(new_n525));
  OAI21_X1  g100(.A(new_n522), .B1(new_n524), .B2(new_n525), .ZN(new_n526));
  NOR2_X1   g101(.A1(new_n520), .A2(new_n526), .ZN(new_n527));
  XNOR2_X1  g102(.A(KEYINPUT74), .B(G88), .ZN(new_n528));
  NAND2_X1  g103(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  AND2_X1   g104(.A1(KEYINPUT72), .A2(G651), .ZN(new_n530));
  NOR2_X1   g105(.A1(KEYINPUT72), .A2(G651), .ZN(new_n531));
  OAI21_X1  g106(.A(KEYINPUT6), .B1(new_n530), .B2(new_n531), .ZN(new_n532));
  INV_X1    g107(.A(new_n518), .ZN(new_n533));
  AOI21_X1  g108(.A(new_n523), .B1(new_n532), .B2(new_n533), .ZN(new_n534));
  NAND2_X1  g109(.A1(new_n534), .A2(G50), .ZN(new_n535));
  INV_X1    g110(.A(new_n519), .ZN(new_n536));
  INV_X1    g111(.A(KEYINPUT73), .ZN(new_n537));
  OAI21_X1  g112(.A(new_n537), .B1(new_n521), .B2(G543), .ZN(new_n538));
  NAND3_X1  g113(.A1(new_n523), .A2(KEYINPUT73), .A3(KEYINPUT5), .ZN(new_n539));
  AOI22_X1  g114(.A1(new_n538), .A2(new_n539), .B1(new_n521), .B2(G543), .ZN(new_n540));
  AOI22_X1  g115(.A1(new_n540), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n541));
  OAI211_X1 g116(.A(new_n529), .B(new_n535), .C1(new_n536), .C2(new_n541), .ZN(G303));
  INV_X1    g117(.A(G303), .ZN(G166));
  NAND2_X1  g118(.A1(new_n532), .A2(new_n533), .ZN(new_n544));
  NAND3_X1  g119(.A1(new_n544), .A2(G89), .A3(new_n540), .ZN(new_n545));
  NAND3_X1  g120(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n546));
  INV_X1    g121(.A(KEYINPUT7), .ZN(new_n547));
  NAND2_X1  g122(.A1(new_n546), .A2(new_n547), .ZN(new_n548));
  INV_X1    g123(.A(new_n534), .ZN(new_n549));
  XNOR2_X1  g124(.A(KEYINPUT75), .B(G51), .ZN(new_n550));
  OAI211_X1 g125(.A(new_n545), .B(new_n548), .C1(new_n549), .C2(new_n550), .ZN(new_n551));
  INV_X1    g126(.A(G651), .ZN(new_n552));
  NAND2_X1  g127(.A1(new_n540), .A2(G63), .ZN(new_n553));
  NAND3_X1  g128(.A1(KEYINPUT7), .A2(G76), .A3(G543), .ZN(new_n554));
  AOI21_X1  g129(.A(new_n552), .B1(new_n553), .B2(new_n554), .ZN(new_n555));
  OR3_X1    g130(.A1(new_n551), .A2(KEYINPUT76), .A3(new_n555), .ZN(new_n556));
  OAI21_X1  g131(.A(KEYINPUT76), .B1(new_n551), .B2(new_n555), .ZN(new_n557));
  NAND2_X1  g132(.A1(new_n556), .A2(new_n557), .ZN(G168));
  NAND2_X1  g133(.A1(new_n534), .A2(G52), .ZN(new_n559));
  INV_X1    g134(.A(new_n527), .ZN(new_n560));
  INV_X1    g135(.A(G90), .ZN(new_n561));
  OAI21_X1  g136(.A(new_n559), .B1(new_n560), .B2(new_n561), .ZN(new_n562));
  AOI22_X1  g137(.A1(new_n540), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n563));
  NOR2_X1   g138(.A1(new_n563), .A2(new_n536), .ZN(new_n564));
  OR2_X1    g139(.A1(new_n562), .A2(new_n564), .ZN(G301));
  INV_X1    g140(.A(G301), .ZN(G171));
  AOI22_X1  g141(.A1(new_n540), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n567));
  OR2_X1    g142(.A1(new_n567), .A2(new_n536), .ZN(new_n568));
  AOI22_X1  g143(.A1(new_n527), .A2(G81), .B1(G43), .B2(new_n534), .ZN(new_n569));
  AND2_X1   g144(.A1(new_n568), .A2(new_n569), .ZN(new_n570));
  NAND2_X1  g145(.A1(new_n570), .A2(G860), .ZN(G153));
  NAND4_X1  g146(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g147(.A1(G1), .A2(G3), .ZN(new_n573));
  XNOR2_X1  g148(.A(new_n573), .B(KEYINPUT8), .ZN(new_n574));
  NAND4_X1  g149(.A1(G319), .A2(G483), .A3(G661), .A4(new_n574), .ZN(G188));
  NAND3_X1  g150(.A1(new_n544), .A2(G91), .A3(new_n540), .ZN(new_n576));
  NAND2_X1  g151(.A1(new_n576), .A2(KEYINPUT79), .ZN(new_n577));
  INV_X1    g152(.A(KEYINPUT79), .ZN(new_n578));
  NAND4_X1  g153(.A1(new_n544), .A2(new_n540), .A3(new_n578), .A4(G91), .ZN(new_n579));
  NAND2_X1  g154(.A1(G78), .A2(G543), .ZN(new_n580));
  INV_X1    g155(.A(G65), .ZN(new_n581));
  OAI21_X1  g156(.A(new_n580), .B1(new_n526), .B2(new_n581), .ZN(new_n582));
  AOI22_X1  g157(.A1(new_n577), .A2(new_n579), .B1(G651), .B2(new_n582), .ZN(new_n583));
  INV_X1    g158(.A(KEYINPUT78), .ZN(new_n584));
  AND2_X1   g159(.A1(KEYINPUT77), .A2(G53), .ZN(new_n585));
  INV_X1    g160(.A(KEYINPUT6), .ZN(new_n586));
  OR2_X1    g161(.A1(KEYINPUT72), .A2(G651), .ZN(new_n587));
  NAND2_X1  g162(.A1(KEYINPUT72), .A2(G651), .ZN(new_n588));
  AOI21_X1  g163(.A(new_n586), .B1(new_n587), .B2(new_n588), .ZN(new_n589));
  OAI211_X1 g164(.A(G543), .B(new_n585), .C1(new_n589), .C2(new_n518), .ZN(new_n590));
  INV_X1    g165(.A(KEYINPUT9), .ZN(new_n591));
  NOR2_X1   g166(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  AOI21_X1  g167(.A(KEYINPUT9), .B1(new_n534), .B2(new_n585), .ZN(new_n593));
  OAI21_X1  g168(.A(new_n584), .B1(new_n592), .B2(new_n593), .ZN(new_n594));
  NAND2_X1  g169(.A1(new_n590), .A2(new_n591), .ZN(new_n595));
  NAND3_X1  g170(.A1(new_n534), .A2(KEYINPUT9), .A3(new_n585), .ZN(new_n596));
  NAND3_X1  g171(.A1(new_n595), .A2(KEYINPUT78), .A3(new_n596), .ZN(new_n597));
  NAND3_X1  g172(.A1(new_n583), .A2(new_n594), .A3(new_n597), .ZN(G299));
  INV_X1    g173(.A(G168), .ZN(G286));
  NAND2_X1  g174(.A1(new_n527), .A2(G87), .ZN(new_n600));
  XNOR2_X1  g175(.A(new_n600), .B(KEYINPUT80), .ZN(new_n601));
  OR2_X1    g176(.A1(new_n540), .A2(G74), .ZN(new_n602));
  AOI22_X1  g177(.A1(new_n602), .A2(G651), .B1(new_n534), .B2(G49), .ZN(new_n603));
  NAND2_X1  g178(.A1(new_n601), .A2(new_n603), .ZN(G288));
  OAI211_X1 g179(.A(G61), .B(new_n522), .C1(new_n524), .C2(new_n525), .ZN(new_n605));
  INV_X1    g180(.A(KEYINPUT81), .ZN(new_n606));
  NAND2_X1  g181(.A1(new_n605), .A2(new_n606), .ZN(new_n607));
  NAND3_X1  g182(.A1(new_n540), .A2(KEYINPUT81), .A3(G61), .ZN(new_n608));
  NAND2_X1  g183(.A1(G73), .A2(G543), .ZN(new_n609));
  NAND3_X1  g184(.A1(new_n607), .A2(new_n608), .A3(new_n609), .ZN(new_n610));
  NAND2_X1  g185(.A1(new_n610), .A2(new_n519), .ZN(new_n611));
  INV_X1    g186(.A(KEYINPUT82), .ZN(new_n612));
  NAND2_X1  g187(.A1(G48), .A2(G543), .ZN(new_n613));
  OAI21_X1  g188(.A(new_n612), .B1(new_n520), .B2(new_n613), .ZN(new_n614));
  INV_X1    g189(.A(new_n613), .ZN(new_n615));
  NAND3_X1  g190(.A1(new_n544), .A2(KEYINPUT82), .A3(new_n615), .ZN(new_n616));
  AOI22_X1  g191(.A1(new_n614), .A2(new_n616), .B1(new_n527), .B2(G86), .ZN(new_n617));
  NAND2_X1  g192(.A1(new_n611), .A2(new_n617), .ZN(G305));
  NAND2_X1  g193(.A1(new_n534), .A2(G47), .ZN(new_n619));
  INV_X1    g194(.A(G85), .ZN(new_n620));
  OAI21_X1  g195(.A(new_n619), .B1(new_n560), .B2(new_n620), .ZN(new_n621));
  XNOR2_X1  g196(.A(new_n621), .B(KEYINPUT83), .ZN(new_n622));
  AOI22_X1  g197(.A1(new_n540), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n623));
  OR2_X1    g198(.A1(new_n623), .A2(new_n536), .ZN(new_n624));
  NAND2_X1  g199(.A1(new_n622), .A2(new_n624), .ZN(G290));
  NAND2_X1  g200(.A1(G301), .A2(G868), .ZN(new_n626));
  NAND2_X1  g201(.A1(new_n527), .A2(G92), .ZN(new_n627));
  INV_X1    g202(.A(KEYINPUT10), .ZN(new_n628));
  XNOR2_X1  g203(.A(new_n627), .B(new_n628), .ZN(new_n629));
  NAND2_X1  g204(.A1(G79), .A2(G543), .ZN(new_n630));
  INV_X1    g205(.A(G66), .ZN(new_n631));
  OAI21_X1  g206(.A(new_n630), .B1(new_n526), .B2(new_n631), .ZN(new_n632));
  AOI22_X1  g207(.A1(new_n632), .A2(G651), .B1(G54), .B2(new_n534), .ZN(new_n633));
  NAND2_X1  g208(.A1(new_n629), .A2(new_n633), .ZN(new_n634));
  INV_X1    g209(.A(new_n634), .ZN(new_n635));
  OAI21_X1  g210(.A(new_n626), .B1(new_n635), .B2(G868), .ZN(G284));
  OAI21_X1  g211(.A(new_n626), .B1(new_n635), .B2(G868), .ZN(G321));
  NOR2_X1   g212(.A1(G299), .A2(G868), .ZN(new_n638));
  AOI21_X1  g213(.A(new_n638), .B1(G868), .B2(G168), .ZN(G297));
  AOI21_X1  g214(.A(new_n638), .B1(G868), .B2(G168), .ZN(G280));
  INV_X1    g215(.A(G559), .ZN(new_n641));
  OAI21_X1  g216(.A(new_n635), .B1(new_n641), .B2(G860), .ZN(G148));
  NAND2_X1  g217(.A1(new_n635), .A2(new_n641), .ZN(new_n643));
  NAND2_X1  g218(.A1(new_n643), .A2(G868), .ZN(new_n644));
  OAI21_X1  g219(.A(new_n644), .B1(G868), .B2(new_n570), .ZN(G323));
  XNOR2_X1  g220(.A(G323), .B(KEYINPUT11), .ZN(G282));
  INV_X1    g221(.A(G111), .ZN(new_n647));
  INV_X1    g222(.A(KEYINPUT85), .ZN(new_n648));
  OAI21_X1  g223(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n649));
  AOI22_X1  g224(.A1(new_n479), .A2(new_n647), .B1(new_n648), .B2(new_n649), .ZN(new_n650));
  OAI21_X1  g225(.A(new_n650), .B1(new_n648), .B2(new_n649), .ZN(new_n651));
  NAND2_X1  g226(.A1(new_n495), .A2(G135), .ZN(new_n652));
  NAND2_X1  g227(.A1(new_n490), .A2(G123), .ZN(new_n653));
  NAND3_X1  g228(.A1(new_n651), .A2(new_n652), .A3(new_n653), .ZN(new_n654));
  INV_X1    g229(.A(new_n654), .ZN(new_n655));
  XNOR2_X1  g230(.A(KEYINPUT86), .B(G2096), .ZN(new_n656));
  OR2_X1    g231(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  NAND2_X1  g232(.A1(new_n655), .A2(new_n656), .ZN(new_n658));
  NAND2_X1  g233(.A1(new_n465), .A2(new_n471), .ZN(new_n659));
  XOR2_X1   g234(.A(KEYINPUT84), .B(KEYINPUT12), .Z(new_n660));
  XNOR2_X1  g235(.A(new_n659), .B(new_n660), .ZN(new_n661));
  XNOR2_X1  g236(.A(KEYINPUT13), .B(G2100), .ZN(new_n662));
  XNOR2_X1  g237(.A(new_n661), .B(new_n662), .ZN(new_n663));
  NAND3_X1  g238(.A1(new_n657), .A2(new_n658), .A3(new_n663), .ZN(G156));
  XNOR2_X1  g239(.A(KEYINPUT15), .B(G2435), .ZN(new_n665));
  XNOR2_X1  g240(.A(new_n665), .B(G2438), .ZN(new_n666));
  XNOR2_X1  g241(.A(G2427), .B(G2430), .ZN(new_n667));
  NAND2_X1  g242(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  NAND2_X1  g243(.A1(new_n668), .A2(KEYINPUT14), .ZN(new_n669));
  XOR2_X1   g244(.A(new_n669), .B(KEYINPUT87), .Z(new_n670));
  OAI21_X1  g245(.A(new_n670), .B1(new_n666), .B2(new_n667), .ZN(new_n671));
  XOR2_X1   g246(.A(G1341), .B(G1348), .Z(new_n672));
  XNOR2_X1  g247(.A(new_n671), .B(new_n672), .ZN(new_n673));
  XNOR2_X1  g248(.A(G2443), .B(G2446), .ZN(new_n674));
  XNOR2_X1  g249(.A(new_n673), .B(new_n674), .ZN(new_n675));
  INV_X1    g250(.A(new_n675), .ZN(new_n676));
  XOR2_X1   g251(.A(G2451), .B(G2454), .Z(new_n677));
  XNOR2_X1  g252(.A(new_n677), .B(KEYINPUT16), .ZN(new_n678));
  XNOR2_X1  g253(.A(new_n678), .B(KEYINPUT88), .ZN(new_n679));
  INV_X1    g254(.A(new_n679), .ZN(new_n680));
  OAI21_X1  g255(.A(G14), .B1(new_n676), .B2(new_n680), .ZN(new_n681));
  AOI21_X1  g256(.A(new_n681), .B1(new_n680), .B2(new_n676), .ZN(G401));
  XOR2_X1   g257(.A(G2072), .B(G2078), .Z(new_n683));
  XOR2_X1   g258(.A(new_n683), .B(KEYINPUT17), .Z(new_n684));
  XOR2_X1   g259(.A(G2084), .B(G2090), .Z(new_n685));
  XNOR2_X1  g260(.A(G2067), .B(G2678), .ZN(new_n686));
  OAI21_X1  g261(.A(new_n684), .B1(new_n685), .B2(new_n686), .ZN(new_n687));
  NAND2_X1  g262(.A1(new_n685), .A2(new_n686), .ZN(new_n688));
  INV_X1    g263(.A(new_n685), .ZN(new_n689));
  NAND2_X1  g264(.A1(new_n689), .A2(new_n683), .ZN(new_n690));
  OAI211_X1 g265(.A(new_n687), .B(new_n688), .C1(new_n686), .C2(new_n690), .ZN(new_n691));
  NOR2_X1   g266(.A1(new_n688), .A2(new_n683), .ZN(new_n692));
  XNOR2_X1  g267(.A(new_n692), .B(KEYINPUT18), .ZN(new_n693));
  NAND2_X1  g268(.A1(new_n691), .A2(new_n693), .ZN(new_n694));
  XOR2_X1   g269(.A(new_n694), .B(G2096), .Z(new_n695));
  XNOR2_X1  g270(.A(new_n695), .B(G2100), .ZN(G227));
  XOR2_X1   g271(.A(G1956), .B(G2474), .Z(new_n697));
  XNOR2_X1  g272(.A(new_n697), .B(KEYINPUT89), .ZN(new_n698));
  XNOR2_X1  g273(.A(G1961), .B(G1966), .ZN(new_n699));
  INV_X1    g274(.A(new_n699), .ZN(new_n700));
  NAND2_X1  g275(.A1(new_n698), .A2(new_n700), .ZN(new_n701));
  XNOR2_X1  g276(.A(G1971), .B(G1976), .ZN(new_n702));
  XNOR2_X1  g277(.A(new_n702), .B(KEYINPUT19), .ZN(new_n703));
  NOR2_X1   g278(.A1(new_n701), .A2(new_n703), .ZN(new_n704));
  XOR2_X1   g279(.A(new_n704), .B(KEYINPUT20), .Z(new_n705));
  NOR2_X1   g280(.A1(new_n698), .A2(new_n700), .ZN(new_n706));
  INV_X1    g281(.A(new_n706), .ZN(new_n707));
  NAND3_X1  g282(.A1(new_n707), .A2(new_n703), .A3(new_n701), .ZN(new_n708));
  OAI211_X1 g283(.A(new_n705), .B(new_n708), .C1(new_n703), .C2(new_n707), .ZN(new_n709));
  XNOR2_X1  g284(.A(new_n709), .B(G1986), .ZN(new_n710));
  XNOR2_X1  g285(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n711));
  XNOR2_X1  g286(.A(new_n710), .B(new_n711), .ZN(new_n712));
  XNOR2_X1  g287(.A(G1991), .B(G1996), .ZN(new_n713));
  INV_X1    g288(.A(G1981), .ZN(new_n714));
  XNOR2_X1  g289(.A(new_n713), .B(new_n714), .ZN(new_n715));
  XNOR2_X1  g290(.A(new_n712), .B(new_n715), .ZN(new_n716));
  INV_X1    g291(.A(new_n716), .ZN(G229));
  INV_X1    g292(.A(new_n603), .ZN(new_n718));
  OR2_X1    g293(.A1(new_n600), .A2(KEYINPUT80), .ZN(new_n719));
  NAND2_X1  g294(.A1(new_n600), .A2(KEYINPUT80), .ZN(new_n720));
  AOI21_X1  g295(.A(new_n718), .B1(new_n719), .B2(new_n720), .ZN(new_n721));
  INV_X1    g296(.A(G16), .ZN(new_n722));
  NOR2_X1   g297(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  AOI21_X1  g298(.A(new_n723), .B1(new_n722), .B2(G23), .ZN(new_n724));
  XOR2_X1   g299(.A(KEYINPUT33), .B(G1976), .Z(new_n725));
  INV_X1    g300(.A(new_n725), .ZN(new_n726));
  OR2_X1    g301(.A1(new_n724), .A2(new_n726), .ZN(new_n727));
  NAND2_X1  g302(.A1(new_n724), .A2(new_n726), .ZN(new_n728));
  NAND2_X1  g303(.A1(new_n722), .A2(G22), .ZN(new_n729));
  OAI21_X1  g304(.A(new_n729), .B1(G166), .B2(new_n722), .ZN(new_n730));
  XOR2_X1   g305(.A(new_n730), .B(G1971), .Z(new_n731));
  NOR2_X1   g306(.A1(G6), .A2(G16), .ZN(new_n732));
  AOI22_X1  g307(.A1(new_n605), .A2(new_n606), .B1(G73), .B2(G543), .ZN(new_n733));
  AOI21_X1  g308(.A(new_n536), .B1(new_n733), .B2(new_n608), .ZN(new_n734));
  NAND3_X1  g309(.A1(new_n544), .A2(G86), .A3(new_n540), .ZN(new_n735));
  AOI21_X1  g310(.A(KEYINPUT82), .B1(new_n544), .B2(new_n615), .ZN(new_n736));
  AOI211_X1 g311(.A(new_n612), .B(new_n613), .C1(new_n532), .C2(new_n533), .ZN(new_n737));
  OAI21_X1  g312(.A(new_n735), .B1(new_n736), .B2(new_n737), .ZN(new_n738));
  NOR2_X1   g313(.A1(new_n734), .A2(new_n738), .ZN(new_n739));
  AOI21_X1  g314(.A(new_n732), .B1(new_n739), .B2(G16), .ZN(new_n740));
  XOR2_X1   g315(.A(KEYINPUT32), .B(G1981), .Z(new_n741));
  XNOR2_X1  g316(.A(new_n740), .B(new_n741), .ZN(new_n742));
  NAND4_X1  g317(.A1(new_n727), .A2(new_n728), .A3(new_n731), .A4(new_n742), .ZN(new_n743));
  XOR2_X1   g318(.A(new_n743), .B(KEYINPUT34), .Z(new_n744));
  NAND2_X1  g319(.A1(new_n722), .A2(G24), .ZN(new_n745));
  INV_X1    g320(.A(G290), .ZN(new_n746));
  OAI21_X1  g321(.A(new_n745), .B1(new_n746), .B2(new_n722), .ZN(new_n747));
  INV_X1    g322(.A(G1986), .ZN(new_n748));
  XNOR2_X1  g323(.A(new_n747), .B(new_n748), .ZN(new_n749));
  AND2_X1   g324(.A1(new_n749), .A2(KEYINPUT90), .ZN(new_n750));
  INV_X1    g325(.A(G29), .ZN(new_n751));
  NAND2_X1  g326(.A1(new_n751), .A2(G25), .ZN(new_n752));
  AOI22_X1  g327(.A1(G119), .A2(new_n490), .B1(new_n495), .B2(G131), .ZN(new_n753));
  OAI221_X1 g328(.A(G2104), .B1(G95), .B2(G2105), .C1(new_n464), .C2(G107), .ZN(new_n754));
  NAND2_X1  g329(.A1(new_n753), .A2(new_n754), .ZN(new_n755));
  INV_X1    g330(.A(new_n755), .ZN(new_n756));
  OAI21_X1  g331(.A(new_n752), .B1(new_n756), .B2(new_n751), .ZN(new_n757));
  XOR2_X1   g332(.A(KEYINPUT35), .B(G1991), .Z(new_n758));
  XOR2_X1   g333(.A(new_n757), .B(new_n758), .Z(new_n759));
  NOR3_X1   g334(.A1(new_n750), .A2(KEYINPUT91), .A3(new_n759), .ZN(new_n760));
  OAI211_X1 g335(.A(new_n744), .B(new_n760), .C1(KEYINPUT90), .C2(new_n749), .ZN(new_n761));
  INV_X1    g336(.A(KEYINPUT36), .ZN(new_n762));
  OR2_X1    g337(.A1(new_n761), .A2(new_n762), .ZN(new_n763));
  NAND2_X1  g338(.A1(new_n761), .A2(new_n762), .ZN(new_n764));
  NAND2_X1  g339(.A1(new_n751), .A2(G32), .ZN(new_n765));
  NAND2_X1  g340(.A1(new_n471), .A2(G105), .ZN(new_n766));
  INV_X1    g341(.A(G141), .ZN(new_n767));
  OAI21_X1  g342(.A(new_n766), .B1(new_n496), .B2(new_n767), .ZN(new_n768));
  NAND2_X1  g343(.A1(new_n490), .A2(G129), .ZN(new_n769));
  NAND3_X1  g344(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n770));
  XOR2_X1   g345(.A(new_n770), .B(KEYINPUT26), .Z(new_n771));
  NAND2_X1  g346(.A1(new_n769), .A2(new_n771), .ZN(new_n772));
  OR2_X1    g347(.A1(new_n768), .A2(new_n772), .ZN(new_n773));
  INV_X1    g348(.A(new_n773), .ZN(new_n774));
  OAI21_X1  g349(.A(new_n765), .B1(new_n774), .B2(new_n751), .ZN(new_n775));
  XOR2_X1   g350(.A(KEYINPUT27), .B(G1996), .Z(new_n776));
  OR2_X1    g351(.A1(new_n775), .A2(new_n776), .ZN(new_n777));
  INV_X1    g352(.A(G28), .ZN(new_n778));
  OR2_X1    g353(.A1(new_n778), .A2(KEYINPUT30), .ZN(new_n779));
  AOI21_X1  g354(.A(G29), .B1(new_n778), .B2(KEYINPUT30), .ZN(new_n780));
  OR2_X1    g355(.A1(KEYINPUT31), .A2(G11), .ZN(new_n781));
  NAND2_X1  g356(.A1(KEYINPUT31), .A2(G11), .ZN(new_n782));
  AOI22_X1  g357(.A1(new_n779), .A2(new_n780), .B1(new_n781), .B2(new_n782), .ZN(new_n783));
  OAI21_X1  g358(.A(new_n783), .B1(new_n654), .B2(new_n751), .ZN(new_n784));
  AOI21_X1  g359(.A(new_n784), .B1(new_n775), .B2(new_n776), .ZN(new_n785));
  AND2_X1   g360(.A1(new_n751), .A2(G33), .ZN(new_n786));
  NAND3_X1  g361(.A1(new_n464), .A2(G103), .A3(G2104), .ZN(new_n787));
  XOR2_X1   g362(.A(new_n787), .B(KEYINPUT25), .Z(new_n788));
  NAND2_X1  g363(.A1(new_n495), .A2(G139), .ZN(new_n789));
  AOI22_X1  g364(.A1(new_n465), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n790));
  OAI211_X1 g365(.A(new_n788), .B(new_n789), .C1(new_n464), .C2(new_n790), .ZN(new_n791));
  AOI21_X1  g366(.A(new_n786), .B1(new_n791), .B2(G29), .ZN(new_n792));
  INV_X1    g367(.A(G2072), .ZN(new_n793));
  NAND2_X1  g368(.A1(new_n792), .A2(new_n793), .ZN(new_n794));
  NOR2_X1   g369(.A1(G164), .A2(new_n751), .ZN(new_n795));
  AOI21_X1  g370(.A(new_n795), .B1(G27), .B2(new_n751), .ZN(new_n796));
  INV_X1    g371(.A(G2078), .ZN(new_n797));
  NAND2_X1  g372(.A1(new_n796), .A2(new_n797), .ZN(new_n798));
  NAND4_X1  g373(.A1(new_n777), .A2(new_n785), .A3(new_n794), .A4(new_n798), .ZN(new_n799));
  NOR2_X1   g374(.A1(new_n796), .A2(new_n797), .ZN(new_n800));
  INV_X1    g375(.A(G35), .ZN(new_n801));
  OR3_X1    g376(.A1(new_n801), .A2(KEYINPUT95), .A3(G29), .ZN(new_n802));
  OAI21_X1  g377(.A(KEYINPUT95), .B1(new_n801), .B2(G29), .ZN(new_n803));
  OAI211_X1 g378(.A(new_n802), .B(new_n803), .C1(G162), .C2(new_n751), .ZN(new_n804));
  XNOR2_X1  g379(.A(KEYINPUT96), .B(KEYINPUT29), .ZN(new_n805));
  XNOR2_X1  g380(.A(new_n805), .B(G2090), .ZN(new_n806));
  XNOR2_X1  g381(.A(new_n804), .B(new_n806), .ZN(new_n807));
  NOR3_X1   g382(.A1(new_n799), .A2(new_n800), .A3(new_n807), .ZN(new_n808));
  NAND2_X1  g383(.A1(new_n751), .A2(G26), .ZN(new_n809));
  XOR2_X1   g384(.A(new_n809), .B(KEYINPUT28), .Z(new_n810));
  NAND2_X1  g385(.A1(new_n490), .A2(G128), .ZN(new_n811));
  XNOR2_X1  g386(.A(new_n811), .B(KEYINPUT93), .ZN(new_n812));
  OR2_X1    g387(.A1(new_n464), .A2(G116), .ZN(new_n813));
  OAI21_X1  g388(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n814));
  INV_X1    g389(.A(new_n814), .ZN(new_n815));
  AOI22_X1  g390(.A1(new_n813), .A2(new_n815), .B1(new_n495), .B2(G140), .ZN(new_n816));
  NAND2_X1  g391(.A1(new_n812), .A2(new_n816), .ZN(new_n817));
  AOI21_X1  g392(.A(new_n810), .B1(new_n817), .B2(G29), .ZN(new_n818));
  XNOR2_X1  g393(.A(new_n818), .B(G2067), .ZN(new_n819));
  INV_X1    g394(.A(KEYINPUT24), .ZN(new_n820));
  INV_X1    g395(.A(G34), .ZN(new_n821));
  AOI21_X1  g396(.A(G29), .B1(new_n820), .B2(new_n821), .ZN(new_n822));
  OAI21_X1  g397(.A(new_n822), .B1(new_n820), .B2(new_n821), .ZN(new_n823));
  OAI21_X1  g398(.A(new_n823), .B1(G160), .B2(new_n751), .ZN(new_n824));
  AND2_X1   g399(.A1(new_n824), .A2(G2084), .ZN(new_n825));
  NAND2_X1  g400(.A1(new_n722), .A2(G5), .ZN(new_n826));
  OAI21_X1  g401(.A(new_n826), .B1(G171), .B2(new_n722), .ZN(new_n827));
  AOI21_X1  g402(.A(new_n825), .B1(new_n827), .B2(G1961), .ZN(new_n828));
  NOR2_X1   g403(.A1(new_n827), .A2(G1961), .ZN(new_n829));
  NAND2_X1  g404(.A1(new_n722), .A2(G19), .ZN(new_n830));
  OAI21_X1  g405(.A(new_n830), .B1(new_n570), .B2(new_n722), .ZN(new_n831));
  XNOR2_X1  g406(.A(new_n831), .B(G1341), .ZN(new_n832));
  NOR2_X1   g407(.A1(new_n824), .A2(G2084), .ZN(new_n833));
  NOR3_X1   g408(.A1(new_n829), .A2(new_n832), .A3(new_n833), .ZN(new_n834));
  NAND4_X1  g409(.A1(new_n808), .A2(new_n819), .A3(new_n828), .A4(new_n834), .ZN(new_n835));
  NAND2_X1  g410(.A1(new_n722), .A2(G4), .ZN(new_n836));
  OAI21_X1  g411(.A(new_n836), .B1(new_n635), .B2(new_n722), .ZN(new_n837));
  XNOR2_X1  g412(.A(KEYINPUT92), .B(G1348), .ZN(new_n838));
  XNOR2_X1  g413(.A(new_n837), .B(new_n838), .ZN(new_n839));
  NOR2_X1   g414(.A1(new_n792), .A2(new_n793), .ZN(new_n840));
  XNOR2_X1  g415(.A(new_n840), .B(KEYINPUT94), .ZN(new_n841));
  NAND2_X1  g416(.A1(new_n839), .A2(new_n841), .ZN(new_n842));
  NAND2_X1  g417(.A1(new_n722), .A2(G20), .ZN(new_n843));
  XOR2_X1   g418(.A(new_n843), .B(KEYINPUT23), .Z(new_n844));
  AOI21_X1  g419(.A(new_n844), .B1(G299), .B2(G16), .ZN(new_n845));
  INV_X1    g420(.A(G1956), .ZN(new_n846));
  XNOR2_X1  g421(.A(new_n845), .B(new_n846), .ZN(new_n847));
  NOR2_X1   g422(.A1(G16), .A2(G21), .ZN(new_n848));
  AOI21_X1  g423(.A(new_n848), .B1(G168), .B2(G16), .ZN(new_n849));
  XNOR2_X1  g424(.A(new_n849), .B(G1966), .ZN(new_n850));
  NOR4_X1   g425(.A1(new_n835), .A2(new_n842), .A3(new_n847), .A4(new_n850), .ZN(new_n851));
  NAND3_X1  g426(.A1(new_n763), .A2(new_n764), .A3(new_n851), .ZN(G150));
  INV_X1    g427(.A(G150), .ZN(G311));
  AOI22_X1  g428(.A1(new_n527), .A2(G93), .B1(G55), .B2(new_n534), .ZN(new_n854));
  AOI22_X1  g429(.A1(new_n540), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n855));
  OAI21_X1  g430(.A(new_n854), .B1(new_n536), .B2(new_n855), .ZN(new_n856));
  XOR2_X1   g431(.A(new_n570), .B(new_n856), .Z(new_n857));
  XOR2_X1   g432(.A(new_n857), .B(KEYINPUT38), .Z(new_n858));
  NAND2_X1  g433(.A1(new_n635), .A2(G559), .ZN(new_n859));
  XNOR2_X1  g434(.A(new_n858), .B(new_n859), .ZN(new_n860));
  AND2_X1   g435(.A1(new_n860), .A2(KEYINPUT39), .ZN(new_n861));
  NOR2_X1   g436(.A1(new_n860), .A2(KEYINPUT39), .ZN(new_n862));
  NOR3_X1   g437(.A1(new_n861), .A2(new_n862), .A3(G860), .ZN(new_n863));
  NAND2_X1  g438(.A1(new_n856), .A2(G860), .ZN(new_n864));
  XNOR2_X1  g439(.A(new_n864), .B(KEYINPUT37), .ZN(new_n865));
  OR2_X1    g440(.A1(new_n863), .A2(new_n865), .ZN(G145));
  XNOR2_X1  g441(.A(new_n516), .B(KEYINPUT97), .ZN(new_n867));
  XNOR2_X1  g442(.A(new_n791), .B(new_n867), .ZN(new_n868));
  XNOR2_X1  g443(.A(new_n868), .B(new_n661), .ZN(new_n869));
  XNOR2_X1  g444(.A(new_n817), .B(new_n773), .ZN(new_n870));
  AOI22_X1  g445(.A1(G130), .A2(new_n490), .B1(new_n495), .B2(G142), .ZN(new_n871));
  OAI221_X1 g446(.A(G2104), .B1(G106), .B2(G2105), .C1(new_n464), .C2(G118), .ZN(new_n872));
  NAND2_X1  g447(.A1(new_n871), .A2(new_n872), .ZN(new_n873));
  XOR2_X1   g448(.A(new_n873), .B(new_n755), .Z(new_n874));
  XNOR2_X1  g449(.A(new_n870), .B(new_n874), .ZN(new_n875));
  XNOR2_X1  g450(.A(new_n869), .B(new_n875), .ZN(new_n876));
  XNOR2_X1  g451(.A(G162), .B(G160), .ZN(new_n877));
  XNOR2_X1  g452(.A(new_n877), .B(new_n654), .ZN(new_n878));
  AOI21_X1  g453(.A(G37), .B1(new_n876), .B2(new_n878), .ZN(new_n879));
  OAI21_X1  g454(.A(new_n879), .B1(new_n878), .B2(new_n876), .ZN(new_n880));
  XNOR2_X1  g455(.A(new_n880), .B(KEYINPUT40), .ZN(G395));
  XNOR2_X1  g456(.A(new_n721), .B(KEYINPUT100), .ZN(new_n882));
  XNOR2_X1  g457(.A(new_n882), .B(new_n739), .ZN(new_n883));
  XNOR2_X1  g458(.A(G290), .B(G166), .ZN(new_n884));
  XNOR2_X1  g459(.A(new_n883), .B(new_n884), .ZN(new_n885));
  XNOR2_X1  g460(.A(new_n885), .B(KEYINPUT42), .ZN(new_n886));
  XOR2_X1   g461(.A(new_n634), .B(G299), .Z(new_n887));
  INV_X1    g462(.A(KEYINPUT41), .ZN(new_n888));
  XNOR2_X1  g463(.A(new_n887), .B(new_n888), .ZN(new_n889));
  XNOR2_X1  g464(.A(new_n857), .B(new_n643), .ZN(new_n890));
  INV_X1    g465(.A(new_n890), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n889), .A2(new_n891), .ZN(new_n892));
  XNOR2_X1  g467(.A(new_n887), .B(KEYINPUT98), .ZN(new_n893));
  AOI22_X1  g468(.A1(new_n892), .A2(KEYINPUT99), .B1(new_n890), .B2(new_n893), .ZN(new_n894));
  OAI21_X1  g469(.A(new_n894), .B1(KEYINPUT99), .B2(new_n892), .ZN(new_n895));
  XNOR2_X1  g470(.A(new_n886), .B(new_n895), .ZN(new_n896));
  MUX2_X1   g471(.A(new_n856), .B(new_n896), .S(G868), .Z(G295));
  MUX2_X1   g472(.A(new_n856), .B(new_n896), .S(G868), .Z(G331));
  XNOR2_X1  g473(.A(G168), .B(G171), .ZN(new_n899));
  XOR2_X1   g474(.A(new_n899), .B(new_n857), .Z(new_n900));
  NAND2_X1  g475(.A1(new_n900), .A2(new_n887), .ZN(new_n901));
  XNOR2_X1  g476(.A(new_n899), .B(new_n857), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n889), .A2(new_n902), .ZN(new_n903));
  AND2_X1   g478(.A1(new_n901), .A2(new_n903), .ZN(new_n904));
  INV_X1    g479(.A(new_n885), .ZN(new_n905));
  AOI21_X1  g480(.A(G37), .B1(new_n904), .B2(new_n905), .ZN(new_n906));
  OAI21_X1  g481(.A(new_n906), .B1(new_n905), .B2(new_n904), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n903), .A2(KEYINPUT102), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n900), .A2(new_n893), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  NOR2_X1   g485(.A1(new_n903), .A2(KEYINPUT102), .ZN(new_n911));
  OAI21_X1  g486(.A(new_n885), .B1(new_n910), .B2(new_n911), .ZN(new_n912));
  AND2_X1   g487(.A1(new_n912), .A2(new_n906), .ZN(new_n913));
  MUX2_X1   g488(.A(new_n907), .B(new_n913), .S(KEYINPUT43), .Z(new_n914));
  NAND2_X1  g489(.A1(new_n914), .A2(KEYINPUT44), .ZN(new_n915));
  INV_X1    g490(.A(KEYINPUT43), .ZN(new_n916));
  NOR2_X1   g491(.A1(new_n904), .A2(new_n905), .ZN(new_n917));
  INV_X1    g492(.A(G37), .ZN(new_n918));
  NAND2_X1  g493(.A1(new_n901), .A2(new_n903), .ZN(new_n919));
  OAI21_X1  g494(.A(new_n918), .B1(new_n919), .B2(new_n885), .ZN(new_n920));
  OAI21_X1  g495(.A(KEYINPUT43), .B1(new_n917), .B2(new_n920), .ZN(new_n921));
  INV_X1    g496(.A(KEYINPUT101), .ZN(new_n922));
  AOI22_X1  g497(.A1(new_n913), .A2(new_n916), .B1(new_n921), .B2(new_n922), .ZN(new_n923));
  NAND3_X1  g498(.A1(new_n907), .A2(KEYINPUT101), .A3(KEYINPUT43), .ZN(new_n924));
  AND2_X1   g499(.A1(new_n923), .A2(new_n924), .ZN(new_n925));
  OAI21_X1  g500(.A(new_n915), .B1(new_n925), .B2(KEYINPUT44), .ZN(G397));
  INV_X1    g501(.A(G40), .ZN(new_n927));
  AOI211_X1 g502(.A(new_n927), .B(new_n468), .C1(new_n481), .C2(new_n487), .ZN(new_n928));
  INV_X1    g503(.A(G1384), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n516), .A2(new_n929), .ZN(new_n930));
  INV_X1    g505(.A(KEYINPUT45), .ZN(new_n931));
  NAND2_X1  g506(.A1(new_n930), .A2(new_n931), .ZN(new_n932));
  NAND3_X1  g507(.A1(new_n928), .A2(new_n932), .A3(KEYINPUT111), .ZN(new_n933));
  XNOR2_X1  g508(.A(KEYINPUT103), .B(KEYINPUT45), .ZN(new_n934));
  INV_X1    g509(.A(new_n934), .ZN(new_n935));
  NAND3_X1  g510(.A1(new_n516), .A2(new_n929), .A3(new_n935), .ZN(new_n936));
  INV_X1    g511(.A(KEYINPUT112), .ZN(new_n937));
  NAND2_X1  g512(.A1(new_n936), .A2(new_n937), .ZN(new_n938));
  NAND4_X1  g513(.A1(new_n516), .A2(KEYINPUT112), .A3(new_n929), .A4(new_n935), .ZN(new_n939));
  NAND2_X1  g514(.A1(new_n938), .A2(new_n939), .ZN(new_n940));
  INV_X1    g515(.A(KEYINPUT111), .ZN(new_n941));
  AOI21_X1  g516(.A(KEYINPUT45), .B1(new_n516), .B2(new_n929), .ZN(new_n942));
  INV_X1    g517(.A(new_n468), .ZN(new_n943));
  AND3_X1   g518(.A1(new_n482), .A2(new_n486), .A3(new_n485), .ZN(new_n944));
  AOI21_X1  g519(.A(new_n486), .B1(new_n482), .B2(new_n485), .ZN(new_n945));
  OAI211_X1 g520(.A(G40), .B(new_n943), .C1(new_n944), .C2(new_n945), .ZN(new_n946));
  OAI21_X1  g521(.A(new_n941), .B1(new_n942), .B2(new_n946), .ZN(new_n947));
  NAND3_X1  g522(.A1(new_n933), .A2(new_n940), .A3(new_n947), .ZN(new_n948));
  INV_X1    g523(.A(G1966), .ZN(new_n949));
  NAND2_X1  g524(.A1(new_n948), .A2(new_n949), .ZN(new_n950));
  NAND2_X1  g525(.A1(new_n930), .A2(KEYINPUT50), .ZN(new_n951));
  INV_X1    g526(.A(KEYINPUT105), .ZN(new_n952));
  INV_X1    g527(.A(KEYINPUT50), .ZN(new_n953));
  NAND3_X1  g528(.A1(new_n516), .A2(new_n953), .A3(new_n929), .ZN(new_n954));
  NAND3_X1  g529(.A1(new_n951), .A2(new_n952), .A3(new_n954), .ZN(new_n955));
  NAND3_X1  g530(.A1(new_n930), .A2(KEYINPUT105), .A3(KEYINPUT50), .ZN(new_n956));
  NAND2_X1  g531(.A1(new_n955), .A2(new_n956), .ZN(new_n957));
  INV_X1    g532(.A(G2084), .ZN(new_n958));
  NAND3_X1  g533(.A1(new_n957), .A2(new_n958), .A3(new_n928), .ZN(new_n959));
  NAND2_X1  g534(.A1(new_n950), .A2(new_n959), .ZN(new_n960));
  NAND2_X1  g535(.A1(new_n960), .A2(G8), .ZN(new_n961));
  NOR2_X1   g536(.A1(new_n961), .A2(G286), .ZN(new_n962));
  INV_X1    g537(.A(G8), .ZN(new_n963));
  INV_X1    g538(.A(G2090), .ZN(new_n964));
  NAND3_X1  g539(.A1(G160), .A2(G40), .A3(new_n964), .ZN(new_n965));
  INV_X1    g540(.A(new_n965), .ZN(new_n966));
  AND3_X1   g541(.A1(new_n516), .A2(new_n953), .A3(new_n929), .ZN(new_n967));
  AOI21_X1  g542(.A(new_n953), .B1(new_n516), .B2(new_n929), .ZN(new_n968));
  NOR3_X1   g543(.A1(new_n967), .A2(new_n968), .A3(KEYINPUT105), .ZN(new_n969));
  INV_X1    g544(.A(new_n956), .ZN(new_n970));
  OAI21_X1  g545(.A(new_n966), .B1(new_n969), .B2(new_n970), .ZN(new_n971));
  NAND2_X1  g546(.A1(new_n930), .A2(new_n934), .ZN(new_n972));
  NAND3_X1  g547(.A1(new_n516), .A2(KEYINPUT45), .A3(new_n929), .ZN(new_n973));
  NAND3_X1  g548(.A1(new_n928), .A2(new_n972), .A3(new_n973), .ZN(new_n974));
  XOR2_X1   g549(.A(KEYINPUT104), .B(G1971), .Z(new_n975));
  INV_X1    g550(.A(new_n975), .ZN(new_n976));
  NAND2_X1  g551(.A1(new_n974), .A2(new_n976), .ZN(new_n977));
  AOI21_X1  g552(.A(new_n963), .B1(new_n971), .B2(new_n977), .ZN(new_n978));
  INV_X1    g553(.A(KEYINPUT55), .ZN(new_n979));
  AND3_X1   g554(.A1(G303), .A2(new_n979), .A3(G8), .ZN(new_n980));
  AOI21_X1  g555(.A(new_n979), .B1(G303), .B2(G8), .ZN(new_n981));
  NOR2_X1   g556(.A1(new_n980), .A2(new_n981), .ZN(new_n982));
  OAI21_X1  g557(.A(new_n962), .B1(new_n978), .B2(new_n982), .ZN(new_n983));
  NOR2_X1   g558(.A1(new_n946), .A2(new_n930), .ZN(new_n984));
  NOR2_X1   g559(.A1(new_n984), .A2(new_n963), .ZN(new_n985));
  INV_X1    g560(.A(new_n985), .ZN(new_n986));
  AOI21_X1  g561(.A(new_n714), .B1(new_n611), .B2(new_n617), .ZN(new_n987));
  INV_X1    g562(.A(new_n987), .ZN(new_n988));
  INV_X1    g563(.A(KEYINPUT108), .ZN(new_n989));
  XOR2_X1   g564(.A(KEYINPUT107), .B(G1981), .Z(new_n990));
  AOI21_X1  g565(.A(new_n989), .B1(new_n739), .B2(new_n990), .ZN(new_n991));
  AND4_X1   g566(.A1(new_n989), .A2(new_n611), .A3(new_n617), .A4(new_n990), .ZN(new_n992));
  OAI21_X1  g567(.A(new_n988), .B1(new_n991), .B2(new_n992), .ZN(new_n993));
  INV_X1    g568(.A(KEYINPUT49), .ZN(new_n994));
  AOI21_X1  g569(.A(new_n986), .B1(new_n993), .B2(new_n994), .ZN(new_n995));
  OAI211_X1 g570(.A(KEYINPUT49), .B(new_n988), .C1(new_n991), .C2(new_n992), .ZN(new_n996));
  NOR2_X1   g571(.A1(new_n996), .A2(KEYINPUT109), .ZN(new_n997));
  INV_X1    g572(.A(KEYINPUT109), .ZN(new_n998));
  NAND3_X1  g573(.A1(new_n611), .A2(new_n617), .A3(new_n990), .ZN(new_n999));
  NAND2_X1  g574(.A1(new_n999), .A2(KEYINPUT108), .ZN(new_n1000));
  NAND4_X1  g575(.A1(new_n611), .A2(new_n617), .A3(new_n989), .A4(new_n990), .ZN(new_n1001));
  AOI21_X1  g576(.A(new_n987), .B1(new_n1000), .B2(new_n1001), .ZN(new_n1002));
  AOI21_X1  g577(.A(new_n998), .B1(new_n1002), .B2(KEYINPUT49), .ZN(new_n1003));
  OAI21_X1  g578(.A(new_n995), .B1(new_n997), .B2(new_n1003), .ZN(new_n1004));
  INV_X1    g579(.A(G1976), .ZN(new_n1005));
  OAI21_X1  g580(.A(new_n985), .B1(G288), .B2(new_n1005), .ZN(new_n1006));
  AND2_X1   g581(.A1(new_n1006), .A2(KEYINPUT52), .ZN(new_n1007));
  INV_X1    g582(.A(KEYINPUT52), .ZN(new_n1008));
  OAI21_X1  g583(.A(new_n1008), .B1(new_n721), .B2(G1976), .ZN(new_n1009));
  NOR2_X1   g584(.A1(new_n1006), .A2(new_n1009), .ZN(new_n1010));
  NOR2_X1   g585(.A1(new_n1007), .A2(new_n1010), .ZN(new_n1011));
  NAND2_X1  g586(.A1(new_n1004), .A2(new_n1011), .ZN(new_n1012));
  OAI21_X1  g587(.A(KEYINPUT63), .B1(new_n983), .B2(new_n1012), .ZN(new_n1013));
  NAND2_X1  g588(.A1(new_n996), .A2(KEYINPUT109), .ZN(new_n1014));
  NAND3_X1  g589(.A1(new_n1002), .A2(new_n998), .A3(KEYINPUT49), .ZN(new_n1015));
  NAND2_X1  g590(.A1(new_n1014), .A2(new_n1015), .ZN(new_n1016));
  AOI211_X1 g591(.A(G1976), .B(G288), .C1(new_n1016), .C2(new_n995), .ZN(new_n1017));
  NAND2_X1  g592(.A1(new_n1000), .A2(new_n1001), .ZN(new_n1018));
  INV_X1    g593(.A(new_n1018), .ZN(new_n1019));
  OAI21_X1  g594(.A(new_n985), .B1(new_n1017), .B2(new_n1019), .ZN(new_n1020));
  INV_X1    g595(.A(KEYINPUT110), .ZN(new_n1021));
  NAND4_X1  g596(.A1(new_n928), .A2(new_n951), .A3(new_n964), .A4(new_n954), .ZN(new_n1022));
  AOI21_X1  g597(.A(new_n963), .B1(new_n977), .B2(new_n1022), .ZN(new_n1023));
  OAI21_X1  g598(.A(new_n1021), .B1(new_n1023), .B2(new_n982), .ZN(new_n1024));
  OR2_X1    g599(.A1(new_n980), .A2(new_n981), .ZN(new_n1025));
  NOR3_X1   g600(.A1(new_n967), .A2(new_n968), .A3(new_n946), .ZN(new_n1026));
  AOI22_X1  g601(.A1(new_n1026), .A2(new_n964), .B1(new_n974), .B2(new_n976), .ZN(new_n1027));
  OAI211_X1 g602(.A(KEYINPUT110), .B(new_n1025), .C1(new_n1027), .C2(new_n963), .ZN(new_n1028));
  AOI21_X1  g603(.A(KEYINPUT63), .B1(new_n1024), .B2(new_n1028), .ZN(new_n1029));
  AOI21_X1  g604(.A(new_n965), .B1(new_n955), .B2(new_n956), .ZN(new_n1030));
  AOI21_X1  g605(.A(new_n935), .B1(new_n516), .B2(new_n929), .ZN(new_n1031));
  NOR2_X1   g606(.A1(new_n1031), .A2(new_n946), .ZN(new_n1032));
  AOI21_X1  g607(.A(new_n975), .B1(new_n1032), .B2(new_n973), .ZN(new_n1033));
  OAI211_X1 g608(.A(new_n982), .B(G8), .C1(new_n1030), .C2(new_n1033), .ZN(new_n1034));
  INV_X1    g609(.A(KEYINPUT106), .ZN(new_n1035));
  NAND2_X1  g610(.A1(new_n1034), .A2(new_n1035), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n971), .A2(new_n977), .ZN(new_n1037));
  NAND4_X1  g612(.A1(new_n1037), .A2(KEYINPUT106), .A3(G8), .A4(new_n982), .ZN(new_n1038));
  AOI22_X1  g613(.A1(new_n962), .A2(new_n1029), .B1(new_n1036), .B2(new_n1038), .ZN(new_n1039));
  OAI211_X1 g614(.A(new_n1013), .B(new_n1020), .C1(new_n1012), .C2(new_n1039), .ZN(new_n1040));
  XOR2_X1   g615(.A(KEYINPUT119), .B(KEYINPUT54), .Z(new_n1041));
  XNOR2_X1  g616(.A(KEYINPUT120), .B(KEYINPUT53), .ZN(new_n1042));
  OAI21_X1  g617(.A(new_n1042), .B1(new_n974), .B2(G2078), .ZN(new_n1043));
  INV_X1    g618(.A(new_n1043), .ZN(new_n1044));
  OAI21_X1  g619(.A(new_n928), .B1(new_n969), .B2(new_n970), .ZN(new_n1045));
  INV_X1    g620(.A(KEYINPUT114), .ZN(new_n1046));
  NAND2_X1  g621(.A1(new_n1045), .A2(new_n1046), .ZN(new_n1047));
  AOI21_X1  g622(.A(new_n946), .B1(new_n955), .B2(new_n956), .ZN(new_n1048));
  NAND2_X1  g623(.A1(new_n1048), .A2(KEYINPUT114), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n1047), .A2(new_n1049), .ZN(new_n1050));
  INV_X1    g625(.A(G1961), .ZN(new_n1051));
  AOI21_X1  g626(.A(new_n1044), .B1(new_n1050), .B2(new_n1051), .ZN(new_n1052));
  NAND2_X1  g627(.A1(new_n797), .A2(KEYINPUT53), .ZN(new_n1053));
  OR2_X1    g628(.A1(new_n948), .A2(new_n1053), .ZN(new_n1054));
  AOI21_X1  g629(.A(G301), .B1(new_n1052), .B2(new_n1054), .ZN(new_n1055));
  AOI21_X1  g630(.A(KEYINPUT114), .B1(new_n957), .B2(new_n928), .ZN(new_n1056));
  AOI211_X1 g631(.A(new_n1046), .B(new_n946), .C1(new_n955), .C2(new_n956), .ZN(new_n1057));
  OAI21_X1  g632(.A(new_n1051), .B1(new_n1056), .B2(new_n1057), .ZN(new_n1058));
  OR2_X1    g633(.A1(new_n974), .A2(new_n1053), .ZN(new_n1059));
  AND4_X1   g634(.A1(G301), .A2(new_n1058), .A3(new_n1043), .A4(new_n1059), .ZN(new_n1060));
  OAI21_X1  g635(.A(new_n1041), .B1(new_n1055), .B2(new_n1060), .ZN(new_n1061));
  NAND3_X1  g636(.A1(new_n1052), .A2(G301), .A3(new_n1054), .ZN(new_n1062));
  NAND3_X1  g637(.A1(new_n1058), .A2(new_n1043), .A3(new_n1059), .ZN(new_n1063));
  NAND2_X1  g638(.A1(new_n1063), .A2(G171), .ZN(new_n1064));
  NAND3_X1  g639(.A1(new_n1062), .A2(new_n1064), .A3(KEYINPUT54), .ZN(new_n1065));
  NAND2_X1  g640(.A1(new_n1061), .A2(new_n1065), .ZN(new_n1066));
  NOR3_X1   g641(.A1(new_n592), .A2(new_n593), .A3(KEYINPUT57), .ZN(new_n1067));
  AOI22_X1  g642(.A1(G299), .A2(KEYINPUT57), .B1(new_n583), .B2(new_n1067), .ZN(new_n1068));
  NAND3_X1  g643(.A1(new_n928), .A2(new_n951), .A3(new_n954), .ZN(new_n1069));
  NAND2_X1  g644(.A1(new_n1069), .A2(new_n846), .ZN(new_n1070));
  XNOR2_X1  g645(.A(KEYINPUT56), .B(G2072), .ZN(new_n1071));
  NAND3_X1  g646(.A1(new_n1032), .A2(new_n973), .A3(new_n1071), .ZN(new_n1072));
  NAND3_X1  g647(.A1(new_n1068), .A2(new_n1070), .A3(new_n1072), .ZN(new_n1073));
  INV_X1    g648(.A(new_n1073), .ZN(new_n1074));
  AOI21_X1  g649(.A(G1348), .B1(new_n1047), .B2(new_n1049), .ZN(new_n1075));
  INV_X1    g650(.A(G2067), .ZN(new_n1076));
  NAND2_X1  g651(.A1(new_n984), .A2(new_n1076), .ZN(new_n1077));
  XNOR2_X1  g652(.A(new_n1077), .B(KEYINPUT113), .ZN(new_n1078));
  INV_X1    g653(.A(new_n1078), .ZN(new_n1079));
  OAI21_X1  g654(.A(new_n635), .B1(new_n1075), .B2(new_n1079), .ZN(new_n1080));
  INV_X1    g655(.A(new_n1071), .ZN(new_n1081));
  OAI22_X1  g656(.A1(new_n1026), .A2(G1956), .B1(new_n974), .B2(new_n1081), .ZN(new_n1082));
  NAND2_X1  g657(.A1(G299), .A2(KEYINPUT57), .ZN(new_n1083));
  NAND2_X1  g658(.A1(new_n1067), .A2(new_n583), .ZN(new_n1084));
  NAND2_X1  g659(.A1(new_n1083), .A2(new_n1084), .ZN(new_n1085));
  NAND2_X1  g660(.A1(new_n1082), .A2(new_n1085), .ZN(new_n1086));
  AOI21_X1  g661(.A(new_n1074), .B1(new_n1080), .B2(new_n1086), .ZN(new_n1087));
  NAND4_X1  g662(.A1(new_n1068), .A2(new_n1070), .A3(KEYINPUT115), .A4(new_n1072), .ZN(new_n1088));
  NAND2_X1  g663(.A1(new_n1088), .A2(KEYINPUT61), .ZN(new_n1089));
  XNOR2_X1  g664(.A(KEYINPUT58), .B(G1341), .ZN(new_n1090));
  OAI22_X1  g665(.A1(new_n974), .A2(G1996), .B1(new_n984), .B2(new_n1090), .ZN(new_n1091));
  NAND2_X1  g666(.A1(new_n1091), .A2(new_n570), .ZN(new_n1092));
  INV_X1    g667(.A(KEYINPUT59), .ZN(new_n1093));
  NAND2_X1  g668(.A1(new_n1092), .A2(new_n1093), .ZN(new_n1094));
  NAND3_X1  g669(.A1(new_n1091), .A2(KEYINPUT59), .A3(new_n570), .ZN(new_n1095));
  AND3_X1   g670(.A1(new_n1089), .A2(new_n1094), .A3(new_n1095), .ZN(new_n1096));
  INV_X1    g671(.A(KEYINPUT116), .ZN(new_n1097));
  NAND3_X1  g672(.A1(new_n1086), .A2(new_n1097), .A3(new_n1073), .ZN(new_n1098));
  NAND3_X1  g673(.A1(new_n1082), .A2(KEYINPUT116), .A3(new_n1085), .ZN(new_n1099));
  INV_X1    g674(.A(KEYINPUT115), .ZN(new_n1100));
  NOR2_X1   g675(.A1(new_n1100), .A2(KEYINPUT61), .ZN(new_n1101));
  NAND3_X1  g676(.A1(new_n1098), .A2(new_n1099), .A3(new_n1101), .ZN(new_n1102));
  INV_X1    g677(.A(G1348), .ZN(new_n1103));
  OAI21_X1  g678(.A(new_n1103), .B1(new_n1056), .B2(new_n1057), .ZN(new_n1104));
  NAND4_X1  g679(.A1(new_n1104), .A2(KEYINPUT60), .A3(new_n634), .A4(new_n1078), .ZN(new_n1105));
  AND3_X1   g680(.A1(new_n1096), .A2(new_n1102), .A3(new_n1105), .ZN(new_n1106));
  INV_X1    g681(.A(KEYINPUT60), .ZN(new_n1107));
  OAI21_X1  g682(.A(new_n1107), .B1(new_n1075), .B2(new_n1079), .ZN(new_n1108));
  NAND3_X1  g683(.A1(new_n1104), .A2(KEYINPUT60), .A3(new_n1078), .ZN(new_n1109));
  NAND3_X1  g684(.A1(new_n1108), .A2(new_n635), .A3(new_n1109), .ZN(new_n1110));
  AOI21_X1  g685(.A(new_n1087), .B1(new_n1106), .B2(new_n1110), .ZN(new_n1111));
  NOR2_X1   g686(.A1(new_n1066), .A2(new_n1111), .ZN(new_n1112));
  INV_X1    g687(.A(KEYINPUT118), .ZN(new_n1113));
  NAND3_X1  g688(.A1(new_n556), .A2(G8), .A3(new_n557), .ZN(new_n1114));
  XNOR2_X1  g689(.A(new_n1114), .B(KEYINPUT117), .ZN(new_n1115));
  AOI22_X1  g690(.A1(new_n958), .A2(new_n1048), .B1(new_n948), .B2(new_n949), .ZN(new_n1116));
  OAI21_X1  g691(.A(new_n1115), .B1(new_n1116), .B2(new_n963), .ZN(new_n1117));
  INV_X1    g692(.A(new_n1114), .ZN(new_n1118));
  NOR2_X1   g693(.A1(new_n1118), .A2(KEYINPUT51), .ZN(new_n1119));
  AOI22_X1  g694(.A1(new_n1117), .A2(KEYINPUT51), .B1(new_n961), .B2(new_n1119), .ZN(new_n1120));
  NOR2_X1   g695(.A1(new_n1116), .A2(new_n1114), .ZN(new_n1121));
  OAI21_X1  g696(.A(new_n1113), .B1(new_n1120), .B2(new_n1121), .ZN(new_n1122));
  AOI21_X1  g697(.A(new_n963), .B1(new_n950), .B2(new_n959), .ZN(new_n1123));
  INV_X1    g698(.A(KEYINPUT117), .ZN(new_n1124));
  XNOR2_X1  g699(.A(new_n1114), .B(new_n1124), .ZN(new_n1125));
  OAI21_X1  g700(.A(KEYINPUT51), .B1(new_n1123), .B2(new_n1125), .ZN(new_n1126));
  OAI21_X1  g701(.A(new_n1119), .B1(new_n1116), .B2(new_n963), .ZN(new_n1127));
  NAND2_X1  g702(.A1(new_n1126), .A2(new_n1127), .ZN(new_n1128));
  INV_X1    g703(.A(new_n1121), .ZN(new_n1129));
  NAND3_X1  g704(.A1(new_n1128), .A2(KEYINPUT118), .A3(new_n1129), .ZN(new_n1130));
  INV_X1    g705(.A(KEYINPUT121), .ZN(new_n1131));
  NAND2_X1  g706(.A1(new_n1036), .A2(new_n1038), .ZN(new_n1132));
  NAND2_X1  g707(.A1(new_n1024), .A2(new_n1028), .ZN(new_n1133));
  NAND2_X1  g708(.A1(new_n1132), .A2(new_n1133), .ZN(new_n1134));
  OAI21_X1  g709(.A(new_n1131), .B1(new_n1134), .B2(new_n1012), .ZN(new_n1135));
  NAND2_X1  g710(.A1(new_n1006), .A2(KEYINPUT52), .ZN(new_n1136));
  OAI21_X1  g711(.A(new_n1136), .B1(new_n1006), .B2(new_n1009), .ZN(new_n1137));
  AOI21_X1  g712(.A(new_n1137), .B1(new_n1016), .B2(new_n995), .ZN(new_n1138));
  NAND4_X1  g713(.A1(new_n1138), .A2(KEYINPUT121), .A3(new_n1132), .A4(new_n1133), .ZN(new_n1139));
  AOI22_X1  g714(.A1(new_n1122), .A2(new_n1130), .B1(new_n1135), .B2(new_n1139), .ZN(new_n1140));
  AOI21_X1  g715(.A(new_n1040), .B1(new_n1112), .B2(new_n1140), .ZN(new_n1141));
  AOI21_X1  g716(.A(KEYINPUT118), .B1(new_n1128), .B2(new_n1129), .ZN(new_n1142));
  AOI211_X1 g717(.A(new_n1113), .B(new_n1121), .C1(new_n1126), .C2(new_n1127), .ZN(new_n1143));
  OAI21_X1  g718(.A(KEYINPUT62), .B1(new_n1142), .B2(new_n1143), .ZN(new_n1144));
  INV_X1    g719(.A(KEYINPUT62), .ZN(new_n1145));
  NAND3_X1  g720(.A1(new_n1122), .A2(new_n1145), .A3(new_n1130), .ZN(new_n1146));
  INV_X1    g721(.A(new_n1055), .ZN(new_n1147));
  AOI21_X1  g722(.A(new_n1147), .B1(new_n1135), .B2(new_n1139), .ZN(new_n1148));
  NAND3_X1  g723(.A1(new_n1144), .A2(new_n1146), .A3(new_n1148), .ZN(new_n1149));
  NAND2_X1  g724(.A1(new_n1149), .A2(KEYINPUT122), .ZN(new_n1150));
  INV_X1    g725(.A(KEYINPUT122), .ZN(new_n1151));
  NAND4_X1  g726(.A1(new_n1144), .A2(new_n1146), .A3(new_n1148), .A4(new_n1151), .ZN(new_n1152));
  NAND3_X1  g727(.A1(new_n1141), .A2(new_n1150), .A3(new_n1152), .ZN(new_n1153));
  NOR2_X1   g728(.A1(new_n972), .A2(new_n946), .ZN(new_n1154));
  XNOR2_X1  g729(.A(new_n817), .B(new_n1076), .ZN(new_n1155));
  XOR2_X1   g730(.A(new_n773), .B(G1996), .Z(new_n1156));
  AND2_X1   g731(.A1(new_n1155), .A2(new_n1156), .ZN(new_n1157));
  NAND2_X1  g732(.A1(new_n756), .A2(new_n758), .ZN(new_n1158));
  OR2_X1    g733(.A1(new_n756), .A2(new_n758), .ZN(new_n1159));
  NAND3_X1  g734(.A1(new_n1157), .A2(new_n1158), .A3(new_n1159), .ZN(new_n1160));
  NAND2_X1  g735(.A1(new_n746), .A2(new_n748), .ZN(new_n1161));
  INV_X1    g736(.A(new_n1161), .ZN(new_n1162));
  OR2_X1    g737(.A1(new_n1160), .A2(new_n1162), .ZN(new_n1163));
  NOR2_X1   g738(.A1(new_n746), .A2(new_n748), .ZN(new_n1164));
  OAI21_X1  g739(.A(new_n1154), .B1(new_n1163), .B2(new_n1164), .ZN(new_n1165));
  NAND2_X1  g740(.A1(new_n1153), .A2(new_n1165), .ZN(new_n1166));
  NAND2_X1  g741(.A1(new_n1155), .A2(new_n774), .ZN(new_n1167));
  NAND2_X1  g742(.A1(new_n1167), .A2(new_n1154), .ZN(new_n1168));
  INV_X1    g743(.A(KEYINPUT124), .ZN(new_n1169));
  XNOR2_X1  g744(.A(new_n1168), .B(new_n1169), .ZN(new_n1170));
  NOR3_X1   g745(.A1(new_n972), .A2(G1996), .A3(new_n946), .ZN(new_n1171));
  OR2_X1    g746(.A1(new_n1171), .A2(KEYINPUT46), .ZN(new_n1172));
  NAND2_X1  g747(.A1(new_n1171), .A2(KEYINPUT46), .ZN(new_n1173));
  NAND3_X1  g748(.A1(new_n1170), .A2(new_n1172), .A3(new_n1173), .ZN(new_n1174));
  INV_X1    g749(.A(KEYINPUT47), .ZN(new_n1175));
  INV_X1    g750(.A(new_n1157), .ZN(new_n1176));
  XNOR2_X1  g751(.A(new_n1158), .B(KEYINPUT123), .ZN(new_n1177));
  OAI22_X1  g752(.A1(new_n1176), .A2(new_n1177), .B1(G2067), .B2(new_n817), .ZN(new_n1178));
  AOI22_X1  g753(.A1(new_n1174), .A2(new_n1175), .B1(new_n1154), .B2(new_n1178), .ZN(new_n1179));
  NAND2_X1  g754(.A1(new_n1160), .A2(new_n1154), .ZN(new_n1180));
  INV_X1    g755(.A(KEYINPUT125), .ZN(new_n1181));
  XNOR2_X1  g756(.A(new_n1180), .B(new_n1181), .ZN(new_n1182));
  NAND2_X1  g757(.A1(new_n1162), .A2(new_n1154), .ZN(new_n1183));
  XNOR2_X1  g758(.A(new_n1183), .B(KEYINPUT48), .ZN(new_n1184));
  NAND2_X1  g759(.A1(new_n1182), .A2(new_n1184), .ZN(new_n1185));
  OAI211_X1 g760(.A(new_n1179), .B(new_n1185), .C1(new_n1175), .C2(new_n1174), .ZN(new_n1186));
  XNOR2_X1  g761(.A(new_n1186), .B(KEYINPUT126), .ZN(new_n1187));
  NAND2_X1  g762(.A1(new_n1166), .A2(new_n1187), .ZN(new_n1188));
  INV_X1    g763(.A(KEYINPUT127), .ZN(new_n1189));
  NAND2_X1  g764(.A1(new_n1188), .A2(new_n1189), .ZN(new_n1190));
  NAND3_X1  g765(.A1(new_n1166), .A2(KEYINPUT127), .A3(new_n1187), .ZN(new_n1191));
  NAND2_X1  g766(.A1(new_n1190), .A2(new_n1191), .ZN(G329));
  assign    G231 = 1'b0;
  NAND2_X1  g767(.A1(new_n923), .A2(new_n924), .ZN(new_n1194));
  NOR4_X1   g768(.A1(G229), .A2(G401), .A3(new_n460), .A4(G227), .ZN(new_n1195));
  NAND3_X1  g769(.A1(new_n1194), .A2(new_n880), .A3(new_n1195), .ZN(G225));
  INV_X1    g770(.A(G225), .ZN(G308));
endmodule


