//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 0 0 0 0 0 0 0 1 0 0 1 1 0 0 1 0 1 1 1 0 1 1 1 1 1 0 0 1 0 0 0 0 1 1 1 0 1 1 0 1 1 1 0 0 1 1 1 1 0 0 1 0 1 0 0 1 0 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:26:02 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n710,
    new_n711, new_n712, new_n713, new_n714, new_n715, new_n716, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n731, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n748, new_n749,
    new_n750, new_n751, new_n752, new_n753, new_n754, new_n755, new_n756,
    new_n757, new_n758, new_n759, new_n760, new_n761, new_n762, new_n763,
    new_n764, new_n766, new_n767, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n786, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n817,
    new_n818, new_n819, new_n820, new_n821, new_n822, new_n823, new_n824,
    new_n825, new_n826, new_n827, new_n828, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n942, new_n943, new_n944, new_n945,
    new_n946, new_n947, new_n948, new_n949, new_n950, new_n951, new_n952,
    new_n953, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n974, new_n975, new_n976,
    new_n977, new_n978, new_n979, new_n980, new_n981, new_n982, new_n983,
    new_n984, new_n985, new_n987, new_n988, new_n989, new_n990, new_n991,
    new_n992, new_n993, new_n994, new_n995, new_n996, new_n998, new_n999,
    new_n1000, new_n1001, new_n1002, new_n1003, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1017, new_n1018,
    new_n1019, new_n1020, new_n1021, new_n1022, new_n1023, new_n1024,
    new_n1025, new_n1026, new_n1027, new_n1028, new_n1029, new_n1030,
    new_n1031, new_n1032, new_n1033, new_n1034, new_n1035, new_n1037,
    new_n1038, new_n1039, new_n1040, new_n1041, new_n1042, new_n1043,
    new_n1044, new_n1045, new_n1046, new_n1047, new_n1048, new_n1049,
    new_n1050, new_n1051, new_n1052, new_n1053, new_n1054;
  NOR2_X1   g000(.A1(G237), .A2(G953), .ZN(new_n187));
  NAND2_X1  g001(.A1(new_n187), .A2(G210), .ZN(new_n188));
  XNOR2_X1  g002(.A(new_n188), .B(KEYINPUT27), .ZN(new_n189));
  XNOR2_X1  g003(.A(KEYINPUT26), .B(G101), .ZN(new_n190));
  XNOR2_X1  g004(.A(new_n189), .B(new_n190), .ZN(new_n191));
  INV_X1    g005(.A(new_n191), .ZN(new_n192));
  INV_X1    g006(.A(KEYINPUT70), .ZN(new_n193));
  INV_X1    g007(.A(G131), .ZN(new_n194));
  INV_X1    g008(.A(KEYINPUT66), .ZN(new_n195));
  INV_X1    g009(.A(G137), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n195), .A2(new_n196), .ZN(new_n197));
  NAND2_X1  g011(.A1(KEYINPUT66), .A2(G137), .ZN(new_n198));
  AOI21_X1  g012(.A(G134), .B1(new_n197), .B2(new_n198), .ZN(new_n199));
  INV_X1    g013(.A(KEYINPUT67), .ZN(new_n200));
  INV_X1    g014(.A(G134), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n201), .A2(KEYINPUT65), .ZN(new_n202));
  INV_X1    g016(.A(KEYINPUT65), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n203), .A2(G134), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n202), .A2(new_n204), .ZN(new_n205));
  AOI22_X1  g019(.A1(new_n199), .A2(new_n200), .B1(new_n205), .B2(new_n196), .ZN(new_n206));
  AND2_X1   g020(.A1(KEYINPUT66), .A2(G137), .ZN(new_n207));
  NOR2_X1   g021(.A1(KEYINPUT66), .A2(G137), .ZN(new_n208));
  OAI21_X1  g022(.A(new_n201), .B1(new_n207), .B2(new_n208), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n209), .A2(KEYINPUT67), .ZN(new_n210));
  AOI21_X1  g024(.A(new_n194), .B1(new_n206), .B2(new_n210), .ZN(new_n211));
  AOI21_X1  g025(.A(KEYINPUT11), .B1(new_n205), .B2(new_n196), .ZN(new_n212));
  NAND3_X1  g026(.A1(new_n202), .A2(new_n204), .A3(G137), .ZN(new_n213));
  AND2_X1   g027(.A1(KEYINPUT11), .A2(G134), .ZN(new_n214));
  NAND3_X1  g028(.A1(new_n197), .A2(new_n198), .A3(new_n214), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n213), .A2(new_n215), .ZN(new_n216));
  NOR3_X1   g030(.A1(new_n212), .A2(new_n216), .A3(G131), .ZN(new_n217));
  OAI21_X1  g031(.A(new_n193), .B1(new_n211), .B2(new_n217), .ZN(new_n218));
  XNOR2_X1  g032(.A(KEYINPUT65), .B(G134), .ZN(new_n219));
  OAI22_X1  g033(.A1(new_n209), .A2(KEYINPUT67), .B1(new_n219), .B2(G137), .ZN(new_n220));
  NOR2_X1   g034(.A1(new_n199), .A2(new_n200), .ZN(new_n221));
  OAI21_X1  g035(.A(G131), .B1(new_n220), .B2(new_n221), .ZN(new_n222));
  INV_X1    g036(.A(KEYINPUT11), .ZN(new_n223));
  OAI21_X1  g037(.A(new_n223), .B1(new_n219), .B2(G137), .ZN(new_n224));
  NAND4_X1  g038(.A1(new_n224), .A2(new_n194), .A3(new_n213), .A4(new_n215), .ZN(new_n225));
  NAND3_X1  g039(.A1(new_n222), .A2(KEYINPUT70), .A3(new_n225), .ZN(new_n226));
  INV_X1    g040(.A(G146), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n227), .A2(G143), .ZN(new_n228));
  INV_X1    g042(.A(G143), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n229), .A2(G146), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n228), .A2(new_n230), .ZN(new_n231));
  OAI21_X1  g045(.A(KEYINPUT1), .B1(new_n229), .B2(G146), .ZN(new_n232));
  NAND3_X1  g046(.A1(new_n231), .A2(G128), .A3(new_n232), .ZN(new_n233));
  INV_X1    g047(.A(G128), .ZN(new_n234));
  OAI211_X1 g048(.A(new_n228), .B(new_n230), .C1(KEYINPUT1), .C2(new_n234), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n233), .A2(new_n235), .ZN(new_n236));
  INV_X1    g050(.A(new_n236), .ZN(new_n237));
  NAND3_X1  g051(.A1(new_n218), .A2(new_n226), .A3(new_n237), .ZN(new_n238));
  INV_X1    g052(.A(G119), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n239), .A2(G116), .ZN(new_n240));
  INV_X1    g054(.A(G116), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n241), .A2(G119), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n240), .A2(new_n242), .ZN(new_n243));
  INV_X1    g057(.A(KEYINPUT68), .ZN(new_n244));
  INV_X1    g058(.A(KEYINPUT2), .ZN(new_n245));
  INV_X1    g059(.A(G113), .ZN(new_n246));
  NAND3_X1  g060(.A1(new_n244), .A2(new_n245), .A3(new_n246), .ZN(new_n247));
  OAI21_X1  g061(.A(KEYINPUT68), .B1(KEYINPUT2), .B2(G113), .ZN(new_n248));
  AND2_X1   g062(.A1(new_n247), .A2(new_n248), .ZN(new_n249));
  NOR2_X1   g063(.A1(new_n245), .A2(new_n246), .ZN(new_n250));
  OAI21_X1  g064(.A(new_n243), .B1(new_n249), .B2(new_n250), .ZN(new_n251));
  AOI22_X1  g065(.A1(new_n247), .A2(new_n248), .B1(KEYINPUT2), .B2(G113), .ZN(new_n252));
  INV_X1    g066(.A(new_n243), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n252), .A2(new_n253), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n251), .A2(new_n254), .ZN(new_n255));
  NAND2_X1  g069(.A1(KEYINPUT0), .A2(G128), .ZN(new_n256));
  INV_X1    g070(.A(new_n256), .ZN(new_n257));
  OR3_X1    g071(.A1(KEYINPUT64), .A2(KEYINPUT0), .A3(G128), .ZN(new_n258));
  AOI21_X1  g072(.A(new_n257), .B1(new_n231), .B2(new_n258), .ZN(new_n259));
  OAI21_X1  g073(.A(KEYINPUT64), .B1(KEYINPUT0), .B2(G128), .ZN(new_n260));
  AOI22_X1  g074(.A1(new_n228), .A2(new_n230), .B1(new_n260), .B2(new_n256), .ZN(new_n261));
  NOR3_X1   g075(.A1(new_n259), .A2(KEYINPUT69), .A3(new_n261), .ZN(new_n262));
  INV_X1    g076(.A(KEYINPUT69), .ZN(new_n263));
  XNOR2_X1  g077(.A(G143), .B(G146), .ZN(new_n264));
  NOR3_X1   g078(.A1(KEYINPUT64), .A2(KEYINPUT0), .A3(G128), .ZN(new_n265));
  OAI21_X1  g079(.A(new_n256), .B1(new_n264), .B2(new_n265), .ZN(new_n266));
  NAND2_X1  g080(.A1(new_n260), .A2(new_n256), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n231), .A2(new_n267), .ZN(new_n268));
  AOI21_X1  g082(.A(new_n263), .B1(new_n266), .B2(new_n268), .ZN(new_n269));
  NOR2_X1   g083(.A1(new_n262), .A2(new_n269), .ZN(new_n270));
  OAI21_X1  g084(.A(G131), .B1(new_n212), .B2(new_n216), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n271), .A2(new_n225), .ZN(new_n272));
  AOI21_X1  g086(.A(new_n255), .B1(new_n270), .B2(new_n272), .ZN(new_n273));
  AOI21_X1  g087(.A(new_n192), .B1(new_n238), .B2(new_n273), .ZN(new_n274));
  INV_X1    g088(.A(KEYINPUT30), .ZN(new_n275));
  AOI21_X1  g089(.A(new_n275), .B1(new_n270), .B2(new_n272), .ZN(new_n276));
  AND2_X1   g090(.A1(new_n238), .A2(new_n276), .ZN(new_n277));
  AND3_X1   g091(.A1(new_n222), .A2(new_n225), .A3(new_n237), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n266), .A2(new_n268), .ZN(new_n279));
  INV_X1    g093(.A(new_n279), .ZN(new_n280));
  AOI21_X1  g094(.A(new_n280), .B1(new_n271), .B2(new_n225), .ZN(new_n281));
  OAI21_X1  g095(.A(new_n275), .B1(new_n278), .B2(new_n281), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n282), .A2(new_n255), .ZN(new_n283));
  OAI21_X1  g097(.A(new_n274), .B1(new_n277), .B2(new_n283), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n284), .A2(KEYINPUT31), .ZN(new_n285));
  XNOR2_X1  g099(.A(KEYINPUT72), .B(KEYINPUT28), .ZN(new_n286));
  NAND2_X1  g100(.A1(new_n238), .A2(new_n273), .ZN(new_n287));
  OAI21_X1  g101(.A(new_n255), .B1(new_n278), .B2(new_n281), .ZN(new_n288));
  AOI21_X1  g102(.A(new_n286), .B1(new_n287), .B2(new_n288), .ZN(new_n289));
  AOI21_X1  g103(.A(KEYINPUT28), .B1(new_n238), .B2(new_n273), .ZN(new_n290));
  OAI21_X1  g104(.A(new_n192), .B1(new_n289), .B2(new_n290), .ZN(new_n291));
  XNOR2_X1  g105(.A(KEYINPUT71), .B(KEYINPUT31), .ZN(new_n292));
  OAI211_X1 g106(.A(new_n274), .B(new_n292), .C1(new_n277), .C2(new_n283), .ZN(new_n293));
  NAND3_X1  g107(.A1(new_n285), .A2(new_n291), .A3(new_n293), .ZN(new_n294));
  NOR2_X1   g108(.A1(G472), .A2(G902), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n294), .A2(new_n295), .ZN(new_n296));
  INV_X1    g110(.A(KEYINPUT32), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n296), .A2(new_n297), .ZN(new_n298));
  NOR3_X1   g112(.A1(new_n297), .A2(G472), .A3(G902), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n294), .A2(new_n299), .ZN(new_n300));
  NAND2_X1  g114(.A1(new_n300), .A2(KEYINPUT73), .ZN(new_n301));
  INV_X1    g115(.A(new_n287), .ZN(new_n302));
  INV_X1    g116(.A(new_n255), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n270), .A2(new_n272), .ZN(new_n304));
  AOI21_X1  g118(.A(new_n303), .B1(new_n238), .B2(new_n304), .ZN(new_n305));
  OAI21_X1  g119(.A(KEYINPUT28), .B1(new_n302), .B2(new_n305), .ZN(new_n306));
  INV_X1    g120(.A(KEYINPUT29), .ZN(new_n307));
  NOR3_X1   g121(.A1(new_n290), .A2(new_n307), .A3(new_n192), .ZN(new_n308));
  AOI21_X1  g122(.A(G902), .B1(new_n306), .B2(new_n308), .ZN(new_n309));
  AND2_X1   g123(.A1(new_n271), .A2(new_n225), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n222), .A2(new_n225), .ZN(new_n311));
  OAI22_X1  g125(.A1(new_n310), .A2(new_n280), .B1(new_n311), .B2(new_n236), .ZN(new_n312));
  AOI21_X1  g126(.A(new_n303), .B1(new_n312), .B2(new_n275), .ZN(new_n313));
  NAND3_X1  g127(.A1(new_n238), .A2(KEYINPUT30), .A3(new_n304), .ZN(new_n314));
  AOI22_X1  g128(.A1(new_n313), .A2(new_n314), .B1(new_n238), .B2(new_n273), .ZN(new_n315));
  OAI21_X1  g129(.A(new_n307), .B1(new_n315), .B2(new_n191), .ZN(new_n316));
  NOR3_X1   g130(.A1(new_n289), .A2(new_n192), .A3(new_n290), .ZN(new_n317));
  OAI21_X1  g131(.A(new_n309), .B1(new_n316), .B2(new_n317), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n318), .A2(G472), .ZN(new_n319));
  INV_X1    g133(.A(KEYINPUT73), .ZN(new_n320));
  NAND3_X1  g134(.A1(new_n294), .A2(new_n320), .A3(new_n299), .ZN(new_n321));
  NAND4_X1  g135(.A1(new_n298), .A2(new_n301), .A3(new_n319), .A4(new_n321), .ZN(new_n322));
  INV_X1    g136(.A(G217), .ZN(new_n323));
  INV_X1    g137(.A(G902), .ZN(new_n324));
  AOI21_X1  g138(.A(new_n323), .B1(G234), .B2(new_n324), .ZN(new_n325));
  INV_X1    g139(.A(KEYINPUT74), .ZN(new_n326));
  OAI21_X1  g140(.A(new_n326), .B1(new_n239), .B2(G128), .ZN(new_n327));
  AOI22_X1  g141(.A1(new_n327), .A2(KEYINPUT23), .B1(new_n239), .B2(G128), .ZN(new_n328));
  INV_X1    g142(.A(KEYINPUT23), .ZN(new_n329));
  OAI211_X1 g143(.A(new_n326), .B(new_n329), .C1(new_n239), .C2(G128), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n328), .A2(new_n330), .ZN(new_n331));
  XNOR2_X1  g145(.A(G119), .B(G128), .ZN(new_n332));
  XOR2_X1   g146(.A(KEYINPUT24), .B(G110), .Z(new_n333));
  OAI22_X1  g147(.A1(new_n331), .A2(G110), .B1(new_n332), .B2(new_n333), .ZN(new_n334));
  INV_X1    g148(.A(G140), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n335), .A2(G125), .ZN(new_n336));
  INV_X1    g150(.A(G125), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n337), .A2(G140), .ZN(new_n338));
  NAND3_X1  g152(.A1(new_n336), .A2(new_n338), .A3(KEYINPUT16), .ZN(new_n339));
  OR3_X1    g153(.A1(new_n337), .A2(KEYINPUT16), .A3(G140), .ZN(new_n340));
  NAND3_X1  g154(.A1(new_n339), .A2(new_n340), .A3(G146), .ZN(new_n341));
  XNOR2_X1  g155(.A(G125), .B(G140), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n342), .A2(new_n227), .ZN(new_n343));
  NAND3_X1  g157(.A1(new_n334), .A2(new_n341), .A3(new_n343), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n339), .A2(new_n340), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n345), .A2(new_n227), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n346), .A2(new_n341), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n331), .A2(G110), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n333), .A2(new_n332), .ZN(new_n349));
  NAND3_X1  g163(.A1(new_n347), .A2(new_n348), .A3(new_n349), .ZN(new_n350));
  XNOR2_X1  g164(.A(KEYINPUT22), .B(G137), .ZN(new_n351));
  INV_X1    g165(.A(G953), .ZN(new_n352));
  NAND3_X1  g166(.A1(new_n352), .A2(G221), .A3(G234), .ZN(new_n353));
  XNOR2_X1  g167(.A(new_n351), .B(new_n353), .ZN(new_n354));
  AND3_X1   g168(.A1(new_n344), .A2(new_n350), .A3(new_n354), .ZN(new_n355));
  AOI21_X1  g169(.A(new_n354), .B1(new_n344), .B2(new_n350), .ZN(new_n356));
  NOR2_X1   g170(.A1(new_n355), .A2(new_n356), .ZN(new_n357));
  AOI21_X1  g171(.A(KEYINPUT25), .B1(new_n357), .B2(new_n324), .ZN(new_n358));
  INV_X1    g172(.A(KEYINPUT25), .ZN(new_n359));
  NOR4_X1   g173(.A1(new_n355), .A2(new_n356), .A3(new_n359), .A4(G902), .ZN(new_n360));
  OAI21_X1  g174(.A(new_n325), .B1(new_n358), .B2(new_n360), .ZN(new_n361));
  NOR2_X1   g175(.A1(new_n325), .A2(G902), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n357), .A2(new_n362), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n361), .A2(new_n363), .ZN(new_n364));
  INV_X1    g178(.A(new_n364), .ZN(new_n365));
  INV_X1    g179(.A(KEYINPUT77), .ZN(new_n366));
  INV_X1    g180(.A(G104), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n367), .A2(G107), .ZN(new_n368));
  INV_X1    g182(.A(G107), .ZN(new_n369));
  AND3_X1   g183(.A1(new_n369), .A2(KEYINPUT3), .A3(G104), .ZN(new_n370));
  AOI21_X1  g184(.A(KEYINPUT3), .B1(new_n369), .B2(G104), .ZN(new_n371));
  OAI21_X1  g185(.A(new_n368), .B1(new_n370), .B2(new_n371), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n372), .A2(KEYINPUT75), .ZN(new_n373));
  INV_X1    g187(.A(KEYINPUT3), .ZN(new_n374));
  OAI21_X1  g188(.A(new_n374), .B1(new_n367), .B2(G107), .ZN(new_n375));
  NAND3_X1  g189(.A1(new_n369), .A2(KEYINPUT3), .A3(G104), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n375), .A2(new_n376), .ZN(new_n377));
  INV_X1    g191(.A(KEYINPUT75), .ZN(new_n378));
  NAND3_X1  g192(.A1(new_n377), .A2(new_n378), .A3(new_n368), .ZN(new_n379));
  NAND3_X1  g193(.A1(new_n373), .A2(new_n379), .A3(G101), .ZN(new_n380));
  INV_X1    g194(.A(G101), .ZN(new_n381));
  OAI211_X1 g195(.A(new_n381), .B(new_n368), .C1(new_n370), .C2(new_n371), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n382), .A2(KEYINPUT4), .ZN(new_n383));
  INV_X1    g197(.A(new_n383), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n380), .A2(new_n384), .ZN(new_n385));
  NOR2_X1   g199(.A1(new_n381), .A2(KEYINPUT4), .ZN(new_n386));
  NAND3_X1  g200(.A1(new_n373), .A2(new_n379), .A3(new_n386), .ZN(new_n387));
  NAND3_X1  g201(.A1(new_n385), .A2(new_n270), .A3(new_n387), .ZN(new_n388));
  INV_X1    g202(.A(KEYINPUT76), .ZN(new_n389));
  OAI21_X1  g203(.A(new_n389), .B1(new_n369), .B2(G104), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n369), .A2(G104), .ZN(new_n391));
  NAND3_X1  g205(.A1(new_n367), .A2(KEYINPUT76), .A3(G107), .ZN(new_n392));
  NAND3_X1  g206(.A1(new_n390), .A2(new_n391), .A3(new_n392), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n393), .A2(G101), .ZN(new_n394));
  NAND4_X1  g208(.A1(new_n394), .A2(new_n382), .A3(new_n235), .A4(new_n233), .ZN(new_n395));
  XNOR2_X1  g209(.A(new_n395), .B(KEYINPUT10), .ZN(new_n396));
  AND3_X1   g210(.A1(new_n388), .A2(new_n396), .A3(new_n310), .ZN(new_n397));
  AOI21_X1  g211(.A(new_n310), .B1(new_n388), .B2(new_n396), .ZN(new_n398));
  XNOR2_X1  g212(.A(G110), .B(G140), .ZN(new_n399));
  INV_X1    g213(.A(G227), .ZN(new_n400));
  NOR2_X1   g214(.A1(new_n400), .A2(G953), .ZN(new_n401));
  XNOR2_X1  g215(.A(new_n399), .B(new_n401), .ZN(new_n402));
  NOR3_X1   g216(.A1(new_n397), .A2(new_n398), .A3(new_n402), .ZN(new_n403));
  INV_X1    g217(.A(new_n402), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n394), .A2(new_n382), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n405), .A2(new_n236), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n406), .A2(new_n395), .ZN(new_n407));
  NAND2_X1  g221(.A1(new_n407), .A2(new_n272), .ZN(new_n408));
  INV_X1    g222(.A(KEYINPUT12), .ZN(new_n409));
  NAND2_X1  g223(.A1(new_n408), .A2(new_n409), .ZN(new_n410));
  NAND3_X1  g224(.A1(new_n407), .A2(KEYINPUT12), .A3(new_n272), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n410), .A2(new_n411), .ZN(new_n412));
  NAND3_X1  g226(.A1(new_n388), .A2(new_n396), .A3(new_n310), .ZN(new_n413));
  AOI21_X1  g227(.A(new_n404), .B1(new_n412), .B2(new_n413), .ZN(new_n414));
  OAI21_X1  g228(.A(new_n366), .B1(new_n403), .B2(new_n414), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n279), .A2(KEYINPUT69), .ZN(new_n416));
  NAND3_X1  g230(.A1(new_n266), .A2(new_n263), .A3(new_n268), .ZN(new_n417));
  NAND3_X1  g231(.A1(new_n387), .A2(new_n416), .A3(new_n417), .ZN(new_n418));
  NOR2_X1   g232(.A1(new_n369), .A2(G104), .ZN(new_n419));
  AOI211_X1 g233(.A(KEYINPUT75), .B(new_n419), .C1(new_n375), .C2(new_n376), .ZN(new_n420));
  AOI21_X1  g234(.A(new_n378), .B1(new_n377), .B2(new_n368), .ZN(new_n421));
  NOR2_X1   g235(.A1(new_n420), .A2(new_n421), .ZN(new_n422));
  AOI21_X1  g236(.A(new_n383), .B1(new_n422), .B2(G101), .ZN(new_n423));
  NOR2_X1   g237(.A1(new_n418), .A2(new_n423), .ZN(new_n424));
  INV_X1    g238(.A(KEYINPUT10), .ZN(new_n425));
  XNOR2_X1  g239(.A(new_n395), .B(new_n425), .ZN(new_n426));
  OAI21_X1  g240(.A(new_n272), .B1(new_n424), .B2(new_n426), .ZN(new_n427));
  NAND3_X1  g241(.A1(new_n427), .A2(new_n413), .A3(new_n404), .ZN(new_n428));
  NOR2_X1   g242(.A1(new_n424), .A2(new_n426), .ZN(new_n429));
  AOI22_X1  g243(.A1(new_n429), .A2(new_n310), .B1(new_n411), .B2(new_n410), .ZN(new_n430));
  OAI211_X1 g244(.A(new_n428), .B(KEYINPUT77), .C1(new_n430), .C2(new_n404), .ZN(new_n431));
  NAND3_X1  g245(.A1(new_n415), .A2(new_n431), .A3(G469), .ZN(new_n432));
  INV_X1    g246(.A(G469), .ZN(new_n433));
  NOR2_X1   g247(.A1(new_n433), .A2(new_n324), .ZN(new_n434));
  OAI21_X1  g248(.A(new_n402), .B1(new_n397), .B2(new_n398), .ZN(new_n435));
  NAND3_X1  g249(.A1(new_n412), .A2(new_n413), .A3(new_n404), .ZN(new_n436));
  AOI21_X1  g250(.A(G902), .B1(new_n435), .B2(new_n436), .ZN(new_n437));
  AOI21_X1  g251(.A(new_n434), .B1(new_n437), .B2(new_n433), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n432), .A2(new_n438), .ZN(new_n439));
  INV_X1    g253(.A(KEYINPUT20), .ZN(new_n440));
  XNOR2_X1  g254(.A(G113), .B(G122), .ZN(new_n441));
  XNOR2_X1  g255(.A(new_n441), .B(new_n367), .ZN(new_n442));
  NAND3_X1  g256(.A1(new_n187), .A2(G143), .A3(G214), .ZN(new_n443));
  INV_X1    g257(.A(new_n443), .ZN(new_n444));
  AOI21_X1  g258(.A(G143), .B1(new_n187), .B2(G214), .ZN(new_n445));
  OAI21_X1  g259(.A(G131), .B1(new_n444), .B2(new_n445), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n187), .A2(G214), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n447), .A2(new_n229), .ZN(new_n448));
  NAND3_X1  g262(.A1(new_n448), .A2(new_n194), .A3(new_n443), .ZN(new_n449));
  AND2_X1   g263(.A1(new_n339), .A2(new_n340), .ZN(new_n450));
  AOI22_X1  g264(.A1(new_n446), .A2(new_n449), .B1(new_n450), .B2(G146), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n336), .A2(new_n338), .ZN(new_n452));
  INV_X1    g266(.A(KEYINPUT19), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n452), .A2(new_n453), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n342), .A2(KEYINPUT19), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n454), .A2(new_n455), .ZN(new_n456));
  AOI21_X1  g270(.A(KEYINPUT84), .B1(new_n456), .B2(new_n227), .ZN(new_n457));
  INV_X1    g271(.A(KEYINPUT84), .ZN(new_n458));
  AOI211_X1 g272(.A(new_n458), .B(G146), .C1(new_n454), .C2(new_n455), .ZN(new_n459));
  OAI21_X1  g273(.A(new_n451), .B1(new_n457), .B2(new_n459), .ZN(new_n460));
  INV_X1    g274(.A(KEYINPUT83), .ZN(new_n461));
  AOI21_X1  g275(.A(new_n461), .B1(new_n342), .B2(new_n227), .ZN(new_n462));
  NOR2_X1   g276(.A1(new_n342), .A2(new_n227), .ZN(new_n463));
  OR2_X1    g277(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n462), .A2(new_n463), .ZN(new_n465));
  NAND2_X1  g279(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  NAND2_X1  g280(.A1(KEYINPUT18), .A2(G131), .ZN(new_n467));
  OAI21_X1  g281(.A(new_n467), .B1(new_n444), .B2(new_n445), .ZN(new_n468));
  NAND4_X1  g282(.A1(new_n448), .A2(KEYINPUT18), .A3(G131), .A4(new_n443), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  NAND2_X1  g284(.A1(new_n466), .A2(new_n470), .ZN(new_n471));
  AOI21_X1  g285(.A(new_n442), .B1(new_n460), .B2(new_n471), .ZN(new_n472));
  AOI22_X1  g286(.A1(new_n464), .A2(new_n465), .B1(new_n469), .B2(new_n468), .ZN(new_n473));
  OAI211_X1 g287(.A(KEYINPUT17), .B(G131), .C1(new_n444), .C2(new_n445), .ZN(new_n474));
  NAND3_X1  g288(.A1(new_n474), .A2(new_n346), .A3(new_n341), .ZN(new_n475));
  NOR3_X1   g289(.A1(new_n444), .A2(new_n445), .A3(G131), .ZN(new_n476));
  AOI21_X1  g290(.A(new_n194), .B1(new_n448), .B2(new_n443), .ZN(new_n477));
  NOR2_X1   g291(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  INV_X1    g292(.A(KEYINPUT17), .ZN(new_n479));
  AOI22_X1  g293(.A1(KEYINPUT85), .A2(new_n475), .B1(new_n478), .B2(new_n479), .ZN(new_n480));
  INV_X1    g294(.A(KEYINPUT85), .ZN(new_n481));
  NAND4_X1  g295(.A1(new_n474), .A2(new_n346), .A3(new_n481), .A4(new_n341), .ZN(new_n482));
  AOI21_X1  g296(.A(new_n473), .B1(new_n480), .B2(new_n482), .ZN(new_n483));
  AOI21_X1  g297(.A(new_n472), .B1(new_n483), .B2(new_n442), .ZN(new_n484));
  NOR2_X1   g298(.A1(G475), .A2(G902), .ZN(new_n485));
  INV_X1    g299(.A(new_n485), .ZN(new_n486));
  OAI211_X1 g300(.A(KEYINPUT86), .B(new_n440), .C1(new_n484), .C2(new_n486), .ZN(new_n487));
  NAND2_X1  g301(.A1(new_n475), .A2(KEYINPUT85), .ZN(new_n488));
  NAND2_X1  g302(.A1(new_n478), .A2(new_n479), .ZN(new_n489));
  NAND3_X1  g303(.A1(new_n488), .A2(new_n482), .A3(new_n489), .ZN(new_n490));
  AND3_X1   g304(.A1(new_n490), .A2(new_n442), .A3(new_n471), .ZN(new_n491));
  AOI21_X1  g305(.A(new_n442), .B1(new_n490), .B2(new_n471), .ZN(new_n492));
  OAI21_X1  g306(.A(new_n324), .B1(new_n491), .B2(new_n492), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n493), .A2(G475), .ZN(new_n494));
  NAND3_X1  g308(.A1(new_n490), .A2(new_n442), .A3(new_n471), .ZN(new_n495));
  INV_X1    g309(.A(new_n442), .ZN(new_n496));
  OAI21_X1  g310(.A(new_n341), .B1(new_n476), .B2(new_n477), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n456), .A2(new_n227), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n498), .A2(new_n458), .ZN(new_n499));
  NAND3_X1  g313(.A1(new_n456), .A2(KEYINPUT84), .A3(new_n227), .ZN(new_n500));
  AOI21_X1  g314(.A(new_n497), .B1(new_n499), .B2(new_n500), .ZN(new_n501));
  OAI21_X1  g315(.A(new_n496), .B1(new_n501), .B2(new_n473), .ZN(new_n502));
  AOI21_X1  g316(.A(new_n486), .B1(new_n495), .B2(new_n502), .ZN(new_n503));
  INV_X1    g317(.A(KEYINPUT86), .ZN(new_n504));
  OAI21_X1  g318(.A(KEYINPUT20), .B1(new_n503), .B2(new_n504), .ZN(new_n505));
  AOI211_X1 g319(.A(KEYINPUT86), .B(new_n486), .C1(new_n495), .C2(new_n502), .ZN(new_n506));
  OAI211_X1 g320(.A(new_n487), .B(new_n494), .C1(new_n505), .C2(new_n506), .ZN(new_n507));
  NOR2_X1   g321(.A1(new_n241), .A2(G122), .ZN(new_n508));
  INV_X1    g322(.A(G122), .ZN(new_n509));
  NOR2_X1   g323(.A1(new_n509), .A2(G116), .ZN(new_n510));
  NOR2_X1   g324(.A1(new_n508), .A2(new_n510), .ZN(new_n511));
  XNOR2_X1  g325(.A(new_n511), .B(new_n369), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n229), .A2(G128), .ZN(new_n513));
  INV_X1    g327(.A(KEYINPUT13), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n234), .A2(G143), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  NOR2_X1   g331(.A1(new_n513), .A2(new_n514), .ZN(new_n518));
  OAI21_X1  g332(.A(G134), .B1(new_n517), .B2(new_n518), .ZN(new_n519));
  NAND3_X1  g333(.A1(new_n219), .A2(new_n513), .A3(new_n516), .ZN(new_n520));
  NAND3_X1  g334(.A1(new_n512), .A2(new_n519), .A3(new_n520), .ZN(new_n521));
  XNOR2_X1  g335(.A(KEYINPUT9), .B(G234), .ZN(new_n522));
  NOR3_X1   g336(.A1(new_n522), .A2(new_n323), .A3(G953), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n513), .A2(new_n516), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n205), .A2(new_n524), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n520), .A2(new_n525), .ZN(new_n526));
  INV_X1    g340(.A(KEYINPUT87), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n511), .A2(new_n369), .ZN(new_n529));
  NAND3_X1  g343(.A1(new_n520), .A2(new_n525), .A3(KEYINPUT87), .ZN(new_n530));
  NAND3_X1  g344(.A1(new_n528), .A2(new_n529), .A3(new_n530), .ZN(new_n531));
  OAI21_X1  g345(.A(KEYINPUT14), .B1(new_n509), .B2(G116), .ZN(new_n532));
  INV_X1    g346(.A(KEYINPUT88), .ZN(new_n533));
  XNOR2_X1  g347(.A(new_n532), .B(new_n533), .ZN(new_n534));
  INV_X1    g348(.A(KEYINPUT14), .ZN(new_n535));
  AOI21_X1  g349(.A(new_n508), .B1(new_n535), .B2(new_n510), .ZN(new_n536));
  AOI21_X1  g350(.A(new_n369), .B1(new_n534), .B2(new_n536), .ZN(new_n537));
  OAI211_X1 g351(.A(new_n521), .B(new_n523), .C1(new_n531), .C2(new_n537), .ZN(new_n538));
  INV_X1    g352(.A(KEYINPUT89), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n538), .A2(new_n539), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n534), .A2(new_n536), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n541), .A2(G107), .ZN(new_n542));
  NAND4_X1  g356(.A1(new_n542), .A2(new_n529), .A3(new_n530), .A4(new_n528), .ZN(new_n543));
  NAND4_X1  g357(.A1(new_n543), .A2(KEYINPUT89), .A3(new_n521), .A4(new_n523), .ZN(new_n544));
  OAI21_X1  g358(.A(new_n521), .B1(new_n531), .B2(new_n537), .ZN(new_n545));
  INV_X1    g359(.A(new_n523), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n545), .A2(new_n546), .ZN(new_n547));
  NAND3_X1  g361(.A1(new_n540), .A2(new_n544), .A3(new_n547), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n548), .A2(new_n324), .ZN(new_n549));
  INV_X1    g363(.A(G478), .ZN(new_n550));
  NOR2_X1   g364(.A1(new_n550), .A2(KEYINPUT15), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n549), .A2(new_n551), .ZN(new_n552));
  NOR2_X1   g366(.A1(KEYINPUT90), .A2(G952), .ZN(new_n553));
  INV_X1    g367(.A(new_n553), .ZN(new_n554));
  NAND2_X1  g368(.A1(KEYINPUT90), .A2(G952), .ZN(new_n555));
  AOI21_X1  g369(.A(G953), .B1(new_n554), .B2(new_n555), .ZN(new_n556));
  INV_X1    g370(.A(G234), .ZN(new_n557));
  INV_X1    g371(.A(G237), .ZN(new_n558));
  OAI21_X1  g372(.A(new_n556), .B1(new_n557), .B2(new_n558), .ZN(new_n559));
  INV_X1    g373(.A(new_n559), .ZN(new_n560));
  XNOR2_X1  g374(.A(KEYINPUT21), .B(G898), .ZN(new_n561));
  AOI211_X1 g375(.A(new_n324), .B(new_n352), .C1(G234), .C2(G237), .ZN(new_n562));
  AOI21_X1  g376(.A(new_n560), .B1(new_n561), .B2(new_n562), .ZN(new_n563));
  INV_X1    g377(.A(new_n563), .ZN(new_n564));
  INV_X1    g378(.A(new_n551), .ZN(new_n565));
  NAND3_X1  g379(.A1(new_n548), .A2(new_n324), .A3(new_n565), .ZN(new_n566));
  NAND3_X1  g380(.A1(new_n552), .A2(new_n564), .A3(new_n566), .ZN(new_n567));
  NOR2_X1   g381(.A1(new_n507), .A2(new_n567), .ZN(new_n568));
  OAI21_X1  g382(.A(G221), .B1(new_n522), .B2(G902), .ZN(new_n569));
  AND3_X1   g383(.A1(new_n439), .A2(new_n568), .A3(new_n569), .ZN(new_n570));
  INV_X1    g384(.A(new_n405), .ZN(new_n571));
  NOR2_X1   g385(.A1(new_n241), .A2(G119), .ZN(new_n572));
  INV_X1    g386(.A(KEYINPUT5), .ZN(new_n573));
  AOI21_X1  g387(.A(new_n246), .B1(new_n572), .B2(new_n573), .ZN(new_n574));
  INV_X1    g388(.A(KEYINPUT78), .ZN(new_n575));
  NAND3_X1  g389(.A1(new_n240), .A2(new_n242), .A3(KEYINPUT5), .ZN(new_n576));
  NAND3_X1  g390(.A1(new_n574), .A2(new_n575), .A3(new_n576), .ZN(new_n577));
  AND3_X1   g391(.A1(new_n240), .A2(new_n242), .A3(KEYINPUT5), .ZN(new_n578));
  OAI21_X1  g392(.A(G113), .B1(new_n240), .B2(KEYINPUT5), .ZN(new_n579));
  OAI21_X1  g393(.A(KEYINPUT78), .B1(new_n578), .B2(new_n579), .ZN(new_n580));
  NAND4_X1  g394(.A1(new_n571), .A2(new_n254), .A3(new_n577), .A4(new_n580), .ZN(new_n581));
  NAND2_X1  g395(.A1(new_n387), .A2(new_n255), .ZN(new_n582));
  OAI21_X1  g396(.A(new_n581), .B1(new_n423), .B2(new_n582), .ZN(new_n583));
  XNOR2_X1  g397(.A(G110), .B(G122), .ZN(new_n584));
  INV_X1    g398(.A(new_n584), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n583), .A2(new_n585), .ZN(new_n586));
  OAI211_X1 g400(.A(new_n581), .B(new_n584), .C1(new_n423), .C2(new_n582), .ZN(new_n587));
  NAND3_X1  g401(.A1(new_n586), .A2(KEYINPUT6), .A3(new_n587), .ZN(new_n588));
  NAND2_X1  g402(.A1(new_n279), .A2(G125), .ZN(new_n589));
  OAI21_X1  g403(.A(new_n589), .B1(G125), .B2(new_n236), .ZN(new_n590));
  AND2_X1   g404(.A1(new_n352), .A2(G224), .ZN(new_n591));
  INV_X1    g405(.A(new_n591), .ZN(new_n592));
  XNOR2_X1  g406(.A(new_n590), .B(new_n592), .ZN(new_n593));
  INV_X1    g407(.A(KEYINPUT6), .ZN(new_n594));
  NAND3_X1  g408(.A1(new_n583), .A2(new_n594), .A3(new_n585), .ZN(new_n595));
  NAND3_X1  g409(.A1(new_n588), .A2(new_n593), .A3(new_n595), .ZN(new_n596));
  INV_X1    g410(.A(KEYINPUT7), .ZN(new_n597));
  AOI21_X1  g411(.A(new_n591), .B1(KEYINPUT80), .B2(new_n597), .ZN(new_n598));
  OAI21_X1  g412(.A(new_n598), .B1(KEYINPUT80), .B2(new_n597), .ZN(new_n599));
  OAI211_X1 g413(.A(new_n589), .B(new_n599), .C1(G125), .C2(new_n236), .ZN(new_n600));
  NAND3_X1  g414(.A1(new_n580), .A2(new_n254), .A3(new_n577), .ZN(new_n601));
  NOR2_X1   g415(.A1(new_n601), .A2(new_n571), .ZN(new_n602));
  XNOR2_X1  g416(.A(KEYINPUT79), .B(KEYINPUT8), .ZN(new_n603));
  XNOR2_X1  g417(.A(new_n584), .B(new_n603), .ZN(new_n604));
  AOI22_X1  g418(.A1(new_n252), .A2(new_n253), .B1(new_n574), .B2(new_n576), .ZN(new_n605));
  OAI21_X1  g419(.A(new_n604), .B1(new_n405), .B2(new_n605), .ZN(new_n606));
  OAI21_X1  g420(.A(new_n600), .B1(new_n602), .B2(new_n606), .ZN(new_n607));
  NOR2_X1   g421(.A1(new_n601), .A2(new_n405), .ZN(new_n608));
  AND2_X1   g422(.A1(new_n387), .A2(new_n255), .ZN(new_n609));
  AOI21_X1  g423(.A(new_n608), .B1(new_n609), .B2(new_n385), .ZN(new_n610));
  AOI21_X1  g424(.A(new_n607), .B1(new_n610), .B2(new_n584), .ZN(new_n611));
  NAND3_X1  g425(.A1(new_n590), .A2(KEYINPUT7), .A3(new_n592), .ZN(new_n612));
  INV_X1    g426(.A(KEYINPUT81), .ZN(new_n613));
  NAND2_X1  g427(.A1(new_n612), .A2(new_n613), .ZN(new_n614));
  NAND4_X1  g428(.A1(new_n590), .A2(KEYINPUT81), .A3(KEYINPUT7), .A4(new_n592), .ZN(new_n615));
  NAND2_X1  g429(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  AOI21_X1  g430(.A(G902), .B1(new_n611), .B2(new_n616), .ZN(new_n617));
  OAI21_X1  g431(.A(G210), .B1(G237), .B2(G902), .ZN(new_n618));
  AND3_X1   g432(.A1(new_n596), .A2(new_n617), .A3(new_n618), .ZN(new_n619));
  AOI21_X1  g433(.A(new_n618), .B1(new_n596), .B2(new_n617), .ZN(new_n620));
  NOR3_X1   g434(.A1(new_n619), .A2(new_n620), .A3(KEYINPUT82), .ZN(new_n621));
  OAI21_X1  g435(.A(G214), .B1(G237), .B2(G902), .ZN(new_n622));
  INV_X1    g436(.A(new_n622), .ZN(new_n623));
  NAND3_X1  g437(.A1(new_n596), .A2(new_n617), .A3(new_n618), .ZN(new_n624));
  INV_X1    g438(.A(KEYINPUT82), .ZN(new_n625));
  NOR2_X1   g439(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  NOR3_X1   g440(.A1(new_n621), .A2(new_n623), .A3(new_n626), .ZN(new_n627));
  NAND4_X1  g441(.A1(new_n322), .A2(new_n365), .A3(new_n570), .A4(new_n627), .ZN(new_n628));
  XNOR2_X1  g442(.A(new_n628), .B(G101), .ZN(G3));
  OAI21_X1  g443(.A(new_n622), .B1(new_n619), .B2(new_n620), .ZN(new_n630));
  NAND2_X1  g444(.A1(new_n630), .A2(KEYINPUT92), .ZN(new_n631));
  XOR2_X1   g445(.A(KEYINPUT93), .B(G478), .Z(new_n632));
  NAND2_X1  g446(.A1(new_n549), .A2(new_n632), .ZN(new_n633));
  INV_X1    g447(.A(KEYINPUT33), .ZN(new_n634));
  NAND2_X1  g448(.A1(new_n548), .A2(new_n634), .ZN(new_n635));
  NAND3_X1  g449(.A1(new_n547), .A2(KEYINPUT33), .A3(new_n538), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n635), .A2(new_n636), .ZN(new_n637));
  NAND2_X1  g451(.A1(new_n324), .A2(G478), .ZN(new_n638));
  OAI21_X1  g452(.A(new_n633), .B1(new_n637), .B2(new_n638), .ZN(new_n639));
  NAND2_X1  g453(.A1(new_n639), .A2(new_n507), .ZN(new_n640));
  INV_X1    g454(.A(new_n640), .ZN(new_n641));
  INV_X1    g455(.A(KEYINPUT92), .ZN(new_n642));
  OAI211_X1 g456(.A(new_n642), .B(new_n622), .C1(new_n619), .C2(new_n620), .ZN(new_n643));
  AND4_X1   g457(.A1(new_n564), .A2(new_n631), .A3(new_n641), .A4(new_n643), .ZN(new_n644));
  NAND2_X1  g458(.A1(KEYINPUT91), .A2(G472), .ZN(new_n645));
  AND3_X1   g459(.A1(new_n294), .A2(new_n324), .A3(new_n645), .ZN(new_n646));
  AOI21_X1  g460(.A(new_n645), .B1(new_n294), .B2(new_n324), .ZN(new_n647));
  NOR2_X1   g461(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  INV_X1    g462(.A(new_n569), .ZN(new_n649));
  AOI211_X1 g463(.A(new_n649), .B(new_n364), .C1(new_n432), .C2(new_n438), .ZN(new_n650));
  NAND3_X1  g464(.A1(new_n644), .A2(new_n648), .A3(new_n650), .ZN(new_n651));
  XOR2_X1   g465(.A(KEYINPUT34), .B(G104), .Z(new_n652));
  XNOR2_X1  g466(.A(new_n651), .B(new_n652), .ZN(G6));
  OR2_X1    g467(.A1(new_n505), .A2(new_n506), .ZN(new_n654));
  AND2_X1   g468(.A1(new_n487), .A2(new_n494), .ZN(new_n655));
  NAND2_X1  g469(.A1(new_n552), .A2(new_n566), .ZN(new_n656));
  NAND3_X1  g470(.A1(new_n654), .A2(new_n655), .A3(new_n656), .ZN(new_n657));
  INV_X1    g471(.A(new_n657), .ZN(new_n658));
  AND4_X1   g472(.A1(new_n564), .A2(new_n631), .A3(new_n658), .A4(new_n643), .ZN(new_n659));
  NAND3_X1  g473(.A1(new_n659), .A2(new_n648), .A3(new_n650), .ZN(new_n660));
  XOR2_X1   g474(.A(KEYINPUT35), .B(G107), .Z(new_n661));
  XNOR2_X1  g475(.A(new_n660), .B(new_n661), .ZN(G9));
  INV_X1    g476(.A(new_n325), .ZN(new_n663));
  NAND2_X1  g477(.A1(new_n357), .A2(new_n324), .ZN(new_n664));
  NAND2_X1  g478(.A1(new_n664), .A2(new_n359), .ZN(new_n665));
  INV_X1    g479(.A(new_n360), .ZN(new_n666));
  AOI21_X1  g480(.A(new_n663), .B1(new_n665), .B2(new_n666), .ZN(new_n667));
  NAND2_X1  g481(.A1(new_n344), .A2(new_n350), .ZN(new_n668));
  INV_X1    g482(.A(new_n354), .ZN(new_n669));
  NOR2_X1   g483(.A1(new_n669), .A2(KEYINPUT36), .ZN(new_n670));
  XNOR2_X1  g484(.A(new_n668), .B(new_n670), .ZN(new_n671));
  AND2_X1   g485(.A1(new_n671), .A2(new_n362), .ZN(new_n672));
  NOR2_X1   g486(.A1(new_n667), .A2(new_n672), .ZN(new_n673));
  NOR3_X1   g487(.A1(new_n646), .A2(new_n647), .A3(new_n673), .ZN(new_n674));
  NAND3_X1  g488(.A1(new_n674), .A2(new_n570), .A3(new_n627), .ZN(new_n675));
  XOR2_X1   g489(.A(KEYINPUT37), .B(G110), .Z(new_n676));
  XNOR2_X1  g490(.A(new_n675), .B(new_n676), .ZN(G12));
  AND3_X1   g491(.A1(new_n294), .A2(new_n320), .A3(new_n299), .ZN(new_n678));
  AOI21_X1  g492(.A(new_n320), .B1(new_n294), .B2(new_n299), .ZN(new_n679));
  NOR2_X1   g493(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  AOI22_X1  g494(.A1(new_n297), .A2(new_n296), .B1(new_n318), .B2(G472), .ZN(new_n681));
  AOI21_X1  g495(.A(new_n673), .B1(new_n680), .B2(new_n681), .ZN(new_n682));
  AOI21_X1  g496(.A(new_n649), .B1(new_n432), .B2(new_n438), .ZN(new_n683));
  AND2_X1   g497(.A1(new_n631), .A2(new_n643), .ZN(new_n684));
  INV_X1    g498(.A(new_n562), .ZN(new_n685));
  OAI21_X1  g499(.A(new_n559), .B1(G900), .B2(new_n685), .ZN(new_n686));
  XNOR2_X1  g500(.A(new_n686), .B(KEYINPUT94), .ZN(new_n687));
  NOR2_X1   g501(.A1(new_n657), .A2(new_n687), .ZN(new_n688));
  NAND4_X1  g502(.A1(new_n682), .A2(new_n683), .A3(new_n684), .A4(new_n688), .ZN(new_n689));
  XNOR2_X1  g503(.A(new_n689), .B(G128), .ZN(G30));
  XOR2_X1   g504(.A(new_n687), .B(KEYINPUT39), .Z(new_n691));
  NAND2_X1  g505(.A1(new_n683), .A2(new_n691), .ZN(new_n692));
  XNOR2_X1  g506(.A(new_n692), .B(KEYINPUT40), .ZN(new_n693));
  OR2_X1    g507(.A1(new_n302), .A2(new_n305), .ZN(new_n694));
  OAI21_X1  g508(.A(new_n324), .B1(new_n694), .B2(new_n191), .ZN(new_n695));
  NOR2_X1   g509(.A1(new_n315), .A2(new_n192), .ZN(new_n696));
  OAI21_X1  g510(.A(G472), .B1(new_n695), .B2(new_n696), .ZN(new_n697));
  NAND4_X1  g511(.A1(new_n298), .A2(new_n301), .A3(new_n321), .A4(new_n697), .ZN(new_n698));
  AND2_X1   g512(.A1(new_n507), .A2(new_n656), .ZN(new_n699));
  NAND4_X1  g513(.A1(new_n698), .A2(new_n622), .A3(new_n673), .A4(new_n699), .ZN(new_n700));
  INV_X1    g514(.A(new_n626), .ZN(new_n701));
  NAND2_X1  g515(.A1(new_n596), .A2(new_n617), .ZN(new_n702));
  INV_X1    g516(.A(new_n618), .ZN(new_n703));
  NAND2_X1  g517(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  NAND3_X1  g518(.A1(new_n704), .A2(new_n625), .A3(new_n624), .ZN(new_n705));
  NAND2_X1  g519(.A1(new_n701), .A2(new_n705), .ZN(new_n706));
  XNOR2_X1  g520(.A(new_n706), .B(KEYINPUT38), .ZN(new_n707));
  OR3_X1    g521(.A1(new_n693), .A2(new_n700), .A3(new_n707), .ZN(new_n708));
  XNOR2_X1  g522(.A(new_n708), .B(G143), .ZN(G45));
  INV_X1    g523(.A(new_n687), .ZN(new_n710));
  AND3_X1   g524(.A1(new_n639), .A2(new_n507), .A3(new_n710), .ZN(new_n711));
  NAND3_X1  g525(.A1(new_n631), .A2(new_n711), .A3(new_n643), .ZN(new_n712));
  INV_X1    g526(.A(KEYINPUT95), .ZN(new_n713));
  NAND2_X1  g527(.A1(new_n712), .A2(new_n713), .ZN(new_n714));
  NAND4_X1  g528(.A1(new_n631), .A2(new_n711), .A3(KEYINPUT95), .A4(new_n643), .ZN(new_n715));
  NAND4_X1  g529(.A1(new_n714), .A2(new_n682), .A3(new_n683), .A4(new_n715), .ZN(new_n716));
  XNOR2_X1  g530(.A(new_n716), .B(G146), .ZN(G48));
  AOI21_X1  g531(.A(new_n364), .B1(new_n680), .B2(new_n681), .ZN(new_n718));
  INV_X1    g532(.A(KEYINPUT96), .ZN(new_n719));
  NAND2_X1  g533(.A1(new_n435), .A2(new_n436), .ZN(new_n720));
  AOI21_X1  g534(.A(new_n433), .B1(new_n720), .B2(new_n324), .ZN(new_n721));
  AOI211_X1 g535(.A(G469), .B(G902), .C1(new_n435), .C2(new_n436), .ZN(new_n722));
  NOR2_X1   g536(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  AOI21_X1  g537(.A(new_n719), .B1(new_n723), .B2(new_n569), .ZN(new_n724));
  NOR4_X1   g538(.A1(new_n721), .A2(new_n722), .A3(KEYINPUT96), .A4(new_n649), .ZN(new_n725));
  NOR2_X1   g539(.A1(new_n724), .A2(new_n725), .ZN(new_n726));
  NAND3_X1  g540(.A1(new_n718), .A2(new_n644), .A3(new_n726), .ZN(new_n727));
  XOR2_X1   g541(.A(KEYINPUT41), .B(G113), .Z(new_n728));
  XNOR2_X1  g542(.A(new_n728), .B(KEYINPUT97), .ZN(new_n729));
  XNOR2_X1  g543(.A(new_n727), .B(new_n729), .ZN(G15));
  NAND3_X1  g544(.A1(new_n659), .A2(new_n718), .A3(new_n726), .ZN(new_n731));
  XNOR2_X1  g545(.A(new_n731), .B(G116), .ZN(G18));
  INV_X1    g546(.A(KEYINPUT98), .ZN(new_n733));
  INV_X1    g547(.A(new_n673), .ZN(new_n734));
  NAND3_X1  g548(.A1(new_n322), .A2(new_n568), .A3(new_n734), .ZN(new_n735));
  NAND2_X1  g549(.A1(new_n720), .A2(new_n324), .ZN(new_n736));
  NAND2_X1  g550(.A1(new_n736), .A2(G469), .ZN(new_n737));
  NAND2_X1  g551(.A1(new_n437), .A2(new_n433), .ZN(new_n738));
  NAND3_X1  g552(.A1(new_n737), .A2(new_n569), .A3(new_n738), .ZN(new_n739));
  INV_X1    g553(.A(new_n739), .ZN(new_n740));
  NAND3_X1  g554(.A1(new_n740), .A2(new_n631), .A3(new_n643), .ZN(new_n741));
  OAI21_X1  g555(.A(new_n733), .B1(new_n735), .B2(new_n741), .ZN(new_n742));
  INV_X1    g556(.A(new_n741), .ZN(new_n743));
  NAND4_X1  g557(.A1(new_n682), .A2(new_n743), .A3(KEYINPUT98), .A4(new_n568), .ZN(new_n744));
  NAND2_X1  g558(.A1(new_n742), .A2(new_n744), .ZN(new_n745));
  XOR2_X1   g559(.A(KEYINPUT99), .B(G119), .Z(new_n746));
  XNOR2_X1  g560(.A(new_n745), .B(new_n746), .ZN(G21));
  NAND2_X1  g561(.A1(new_n739), .A2(KEYINPUT96), .ZN(new_n748));
  NAND4_X1  g562(.A1(new_n737), .A2(new_n719), .A3(new_n738), .A4(new_n569), .ZN(new_n749));
  NAND3_X1  g563(.A1(new_n748), .A2(new_n564), .A3(new_n749), .ZN(new_n750));
  NAND2_X1  g564(.A1(new_n364), .A2(KEYINPUT100), .ZN(new_n751));
  INV_X1    g565(.A(KEYINPUT100), .ZN(new_n752));
  NAND3_X1  g566(.A1(new_n361), .A2(new_n363), .A3(new_n752), .ZN(new_n753));
  NAND2_X1  g567(.A1(new_n751), .A2(new_n753), .ZN(new_n754));
  NAND2_X1  g568(.A1(new_n294), .A2(new_n324), .ZN(new_n755));
  NAND2_X1  g569(.A1(new_n755), .A2(G472), .ZN(new_n756));
  NAND2_X1  g570(.A1(new_n285), .A2(new_n293), .ZN(new_n757));
  INV_X1    g571(.A(new_n290), .ZN(new_n758));
  AOI21_X1  g572(.A(new_n191), .B1(new_n306), .B2(new_n758), .ZN(new_n759));
  OAI21_X1  g573(.A(new_n295), .B1(new_n757), .B2(new_n759), .ZN(new_n760));
  NAND3_X1  g574(.A1(new_n754), .A2(new_n756), .A3(new_n760), .ZN(new_n761));
  NOR2_X1   g575(.A1(new_n750), .A2(new_n761), .ZN(new_n762));
  AND3_X1   g576(.A1(new_n631), .A2(new_n699), .A3(new_n643), .ZN(new_n763));
  NAND2_X1  g577(.A1(new_n762), .A2(new_n763), .ZN(new_n764));
  XNOR2_X1  g578(.A(new_n764), .B(G122), .ZN(G24));
  NAND4_X1  g579(.A1(new_n711), .A2(new_n756), .A3(new_n734), .A4(new_n760), .ZN(new_n766));
  NOR2_X1   g580(.A1(new_n741), .A2(new_n766), .ZN(new_n767));
  XNOR2_X1  g581(.A(new_n767), .B(new_n337), .ZN(G27));
  NAND3_X1  g582(.A1(new_n298), .A2(new_n319), .A3(new_n300), .ZN(new_n769));
  NAND2_X1  g583(.A1(new_n769), .A2(new_n754), .ZN(new_n770));
  AOI21_X1  g584(.A(new_n623), .B1(new_n701), .B2(new_n705), .ZN(new_n771));
  XOR2_X1   g585(.A(new_n434), .B(KEYINPUT101), .Z(new_n772));
  INV_X1    g586(.A(new_n772), .ZN(new_n773));
  NOR2_X1   g587(.A1(new_n403), .A2(new_n414), .ZN(new_n774));
  AOI21_X1  g588(.A(new_n773), .B1(new_n774), .B2(G469), .ZN(new_n775));
  AOI21_X1  g589(.A(new_n649), .B1(new_n775), .B2(new_n738), .ZN(new_n776));
  NAND3_X1  g590(.A1(new_n771), .A2(new_n711), .A3(new_n776), .ZN(new_n777));
  OAI21_X1  g591(.A(KEYINPUT42), .B1(new_n770), .B2(new_n777), .ZN(new_n778));
  OAI211_X1 g592(.A(new_n776), .B(new_n622), .C1(new_n621), .C2(new_n626), .ZN(new_n779));
  INV_X1    g593(.A(new_n779), .ZN(new_n780));
  NOR3_X1   g594(.A1(new_n640), .A2(KEYINPUT42), .A3(new_n687), .ZN(new_n781));
  NAND4_X1  g595(.A1(new_n780), .A2(new_n322), .A3(new_n365), .A4(new_n781), .ZN(new_n782));
  NAND2_X1  g596(.A1(new_n778), .A2(new_n782), .ZN(new_n783));
  XOR2_X1   g597(.A(KEYINPUT102), .B(G131), .Z(new_n784));
  XNOR2_X1  g598(.A(new_n783), .B(new_n784), .ZN(G33));
  NAND4_X1  g599(.A1(new_n780), .A2(new_n322), .A3(new_n365), .A4(new_n688), .ZN(new_n786));
  XNOR2_X1  g600(.A(new_n786), .B(G134), .ZN(G36));
  AOI21_X1  g601(.A(new_n433), .B1(new_n774), .B2(KEYINPUT45), .ZN(new_n788));
  INV_X1    g602(.A(new_n788), .ZN(new_n789));
  AOI21_X1  g603(.A(KEYINPUT45), .B1(new_n415), .B2(new_n431), .ZN(new_n790));
  OR3_X1    g604(.A1(new_n789), .A2(new_n790), .A3(KEYINPUT103), .ZN(new_n791));
  OAI21_X1  g605(.A(KEYINPUT103), .B1(new_n789), .B2(new_n790), .ZN(new_n792));
  NAND2_X1  g606(.A1(new_n791), .A2(new_n792), .ZN(new_n793));
  INV_X1    g607(.A(new_n793), .ZN(new_n794));
  NAND2_X1  g608(.A1(new_n772), .A2(KEYINPUT46), .ZN(new_n795));
  OAI211_X1 g609(.A(KEYINPUT104), .B(new_n738), .C1(new_n794), .C2(new_n795), .ZN(new_n796));
  INV_X1    g610(.A(KEYINPUT104), .ZN(new_n797));
  AOI21_X1  g611(.A(new_n795), .B1(new_n791), .B2(new_n792), .ZN(new_n798));
  OAI21_X1  g612(.A(new_n797), .B1(new_n798), .B2(new_n722), .ZN(new_n799));
  NOR2_X1   g613(.A1(new_n794), .A2(new_n773), .ZN(new_n800));
  OAI211_X1 g614(.A(new_n796), .B(new_n799), .C1(KEYINPUT46), .C2(new_n800), .ZN(new_n801));
  AND3_X1   g615(.A1(new_n801), .A2(new_n569), .A3(new_n691), .ZN(new_n802));
  OR3_X1    g616(.A1(new_n648), .A2(KEYINPUT105), .A3(new_n673), .ZN(new_n803));
  OAI21_X1  g617(.A(KEYINPUT105), .B1(new_n648), .B2(new_n673), .ZN(new_n804));
  AND3_X1   g618(.A1(new_n654), .A2(new_n639), .A3(new_n655), .ZN(new_n805));
  XNOR2_X1  g619(.A(new_n805), .B(KEYINPUT43), .ZN(new_n806));
  NAND3_X1  g620(.A1(new_n803), .A2(new_n804), .A3(new_n806), .ZN(new_n807));
  INV_X1    g621(.A(KEYINPUT44), .ZN(new_n808));
  NAND2_X1  g622(.A1(new_n807), .A2(new_n808), .ZN(new_n809));
  NAND4_X1  g623(.A1(new_n803), .A2(KEYINPUT44), .A3(new_n804), .A4(new_n806), .ZN(new_n810));
  NAND3_X1  g624(.A1(new_n809), .A2(new_n771), .A3(new_n810), .ZN(new_n811));
  NAND2_X1  g625(.A1(new_n811), .A2(KEYINPUT106), .ZN(new_n812));
  INV_X1    g626(.A(KEYINPUT106), .ZN(new_n813));
  NAND4_X1  g627(.A1(new_n809), .A2(new_n813), .A3(new_n771), .A4(new_n810), .ZN(new_n814));
  NAND3_X1  g628(.A1(new_n802), .A2(new_n812), .A3(new_n814), .ZN(new_n815));
  XNOR2_X1  g629(.A(new_n815), .B(G137), .ZN(G39));
  NAND2_X1  g630(.A1(new_n801), .A2(new_n569), .ZN(new_n817));
  XNOR2_X1  g631(.A(KEYINPUT107), .B(KEYINPUT47), .ZN(new_n818));
  INV_X1    g632(.A(new_n818), .ZN(new_n819));
  NAND2_X1  g633(.A1(new_n817), .A2(new_n819), .ZN(new_n820));
  NAND3_X1  g634(.A1(new_n801), .A2(new_n569), .A3(new_n818), .ZN(new_n821));
  NAND2_X1  g635(.A1(new_n771), .A2(new_n711), .ZN(new_n822));
  NOR3_X1   g636(.A1(new_n822), .A2(new_n322), .A3(new_n365), .ZN(new_n823));
  NAND3_X1  g637(.A1(new_n820), .A2(new_n821), .A3(new_n823), .ZN(new_n824));
  NAND2_X1  g638(.A1(new_n824), .A2(KEYINPUT108), .ZN(new_n825));
  INV_X1    g639(.A(KEYINPUT108), .ZN(new_n826));
  NAND4_X1  g640(.A1(new_n820), .A2(new_n826), .A3(new_n821), .A4(new_n823), .ZN(new_n827));
  NAND2_X1  g641(.A1(new_n825), .A2(new_n827), .ZN(new_n828));
  XNOR2_X1  g642(.A(new_n828), .B(G140), .ZN(G42));
  OAI21_X1  g643(.A(new_n622), .B1(new_n621), .B2(new_n626), .ZN(new_n830));
  NAND2_X1  g644(.A1(new_n806), .A2(new_n560), .ZN(new_n831));
  NOR2_X1   g645(.A1(new_n831), .A2(KEYINPUT112), .ZN(new_n832));
  INV_X1    g646(.A(new_n832), .ZN(new_n833));
  NAND2_X1  g647(.A1(new_n831), .A2(KEYINPUT112), .ZN(new_n834));
  AOI211_X1 g648(.A(new_n739), .B(new_n830), .C1(new_n833), .C2(new_n834), .ZN(new_n835));
  INV_X1    g649(.A(new_n770), .ZN(new_n836));
  XOR2_X1   g650(.A(KEYINPUT117), .B(KEYINPUT48), .Z(new_n837));
  NAND3_X1  g651(.A1(new_n835), .A2(new_n836), .A3(new_n837), .ZN(new_n838));
  INV_X1    g652(.A(new_n837), .ZN(new_n839));
  NOR2_X1   g653(.A1(new_n830), .A2(new_n739), .ZN(new_n840));
  INV_X1    g654(.A(new_n834), .ZN(new_n841));
  OAI21_X1  g655(.A(new_n840), .B1(new_n841), .B2(new_n832), .ZN(new_n842));
  OAI21_X1  g656(.A(new_n839), .B1(new_n842), .B2(new_n770), .ZN(new_n843));
  AOI21_X1  g657(.A(new_n761), .B1(new_n833), .B2(new_n834), .ZN(new_n844));
  NAND2_X1  g658(.A1(new_n844), .A2(new_n743), .ZN(new_n845));
  XOR2_X1   g659(.A(new_n556), .B(KEYINPUT116), .Z(new_n846));
  INV_X1    g660(.A(new_n698), .ZN(new_n847));
  AND4_X1   g661(.A1(new_n365), .A2(new_n847), .A3(new_n560), .A4(new_n840), .ZN(new_n848));
  AOI21_X1  g662(.A(new_n846), .B1(new_n848), .B2(new_n641), .ZN(new_n849));
  NAND4_X1  g663(.A1(new_n838), .A2(new_n843), .A3(new_n845), .A4(new_n849), .ZN(new_n850));
  NAND2_X1  g664(.A1(new_n844), .A2(new_n771), .ZN(new_n851));
  XNOR2_X1  g665(.A(new_n851), .B(KEYINPUT113), .ZN(new_n852));
  AOI22_X1  g666(.A1(new_n820), .A2(new_n821), .B1(new_n649), .B2(new_n723), .ZN(new_n853));
  OR2_X1    g667(.A1(new_n852), .A2(new_n853), .ZN(new_n854));
  NOR2_X1   g668(.A1(new_n639), .A2(new_n507), .ZN(new_n855));
  NAND2_X1  g669(.A1(new_n848), .A2(new_n855), .ZN(new_n856));
  NAND3_X1  g670(.A1(new_n756), .A2(new_n734), .A3(new_n760), .ZN(new_n857));
  OAI21_X1  g671(.A(new_n856), .B1(new_n842), .B2(new_n857), .ZN(new_n858));
  NAND3_X1  g672(.A1(new_n707), .A2(new_n623), .A3(new_n740), .ZN(new_n859));
  XNOR2_X1  g673(.A(new_n859), .B(KEYINPUT114), .ZN(new_n860));
  INV_X1    g674(.A(new_n860), .ZN(new_n861));
  NAND3_X1  g675(.A1(new_n861), .A2(KEYINPUT50), .A3(new_n844), .ZN(new_n862));
  INV_X1    g676(.A(KEYINPUT50), .ZN(new_n863));
  INV_X1    g677(.A(new_n761), .ZN(new_n864));
  OAI21_X1  g678(.A(new_n864), .B1(new_n841), .B2(new_n832), .ZN(new_n865));
  OAI21_X1  g679(.A(new_n863), .B1(new_n865), .B2(new_n860), .ZN(new_n866));
  AOI21_X1  g680(.A(new_n858), .B1(new_n862), .B2(new_n866), .ZN(new_n867));
  AND2_X1   g681(.A1(new_n867), .A2(KEYINPUT51), .ZN(new_n868));
  AOI21_X1  g682(.A(new_n850), .B1(new_n854), .B2(new_n868), .ZN(new_n869));
  INV_X1    g683(.A(KEYINPUT51), .ZN(new_n870));
  INV_X1    g684(.A(KEYINPUT115), .ZN(new_n871));
  OAI22_X1  g685(.A1(new_n852), .A2(new_n853), .B1(new_n867), .B2(new_n871), .ZN(new_n872));
  AND2_X1   g686(.A1(new_n867), .A2(new_n871), .ZN(new_n873));
  OAI21_X1  g687(.A(new_n870), .B1(new_n872), .B2(new_n873), .ZN(new_n874));
  NAND2_X1  g688(.A1(new_n869), .A2(new_n874), .ZN(new_n875));
  INV_X1    g689(.A(new_n767), .ZN(new_n876));
  NOR2_X1   g690(.A1(new_n734), .A2(new_n687), .ZN(new_n877));
  NAND4_X1  g691(.A1(new_n763), .A2(new_n698), .A3(new_n776), .A4(new_n877), .ZN(new_n878));
  NAND4_X1  g692(.A1(new_n716), .A2(new_n689), .A3(new_n876), .A4(new_n878), .ZN(new_n879));
  NAND2_X1  g693(.A1(new_n879), .A2(KEYINPUT52), .ZN(new_n880));
  AND3_X1   g694(.A1(new_n322), .A2(new_n683), .A3(new_n734), .ZN(new_n881));
  AND2_X1   g695(.A1(new_n684), .A2(new_n688), .ZN(new_n882));
  AOI21_X1  g696(.A(new_n767), .B1(new_n881), .B2(new_n882), .ZN(new_n883));
  INV_X1    g697(.A(KEYINPUT52), .ZN(new_n884));
  NAND4_X1  g698(.A1(new_n883), .A2(new_n884), .A3(new_n716), .A4(new_n878), .ZN(new_n885));
  AND2_X1   g699(.A1(new_n880), .A2(new_n885), .ZN(new_n886));
  NAND2_X1  g700(.A1(new_n683), .A2(new_n568), .ZN(new_n887));
  NOR3_X1   g701(.A1(new_n887), .A2(new_n623), .A3(new_n706), .ZN(new_n888));
  OAI21_X1  g702(.A(new_n888), .B1(new_n718), .B2(new_n674), .ZN(new_n889));
  AOI21_X1  g703(.A(new_n563), .B1(new_n657), .B2(new_n640), .ZN(new_n890));
  NAND4_X1  g704(.A1(new_n627), .A2(new_n648), .A3(new_n650), .A4(new_n890), .ZN(new_n891));
  AOI21_X1  g705(.A(KEYINPUT109), .B1(new_n889), .B2(new_n891), .ZN(new_n892));
  AND4_X1   g706(.A1(KEYINPUT109), .A2(new_n628), .A3(new_n675), .A4(new_n891), .ZN(new_n893));
  NOR2_X1   g707(.A1(new_n892), .A2(new_n893), .ZN(new_n894));
  AND3_X1   g708(.A1(new_n726), .A2(new_n322), .A3(new_n365), .ZN(new_n895));
  AOI22_X1  g709(.A1(new_n895), .A2(new_n644), .B1(new_n762), .B2(new_n763), .ZN(new_n896));
  NAND3_X1  g710(.A1(new_n745), .A2(new_n896), .A3(new_n731), .ZN(new_n897));
  NOR2_X1   g711(.A1(new_n894), .A2(new_n897), .ZN(new_n898));
  AND3_X1   g712(.A1(new_n548), .A2(new_n324), .A3(new_n565), .ZN(new_n899));
  AOI21_X1  g713(.A(new_n565), .B1(new_n548), .B2(new_n324), .ZN(new_n900));
  NOR3_X1   g714(.A1(new_n899), .A2(new_n900), .A3(new_n687), .ZN(new_n901));
  INV_X1    g715(.A(KEYINPUT110), .ZN(new_n902));
  NAND4_X1  g716(.A1(new_n901), .A2(new_n654), .A3(new_n655), .A4(new_n902), .ZN(new_n903));
  NAND3_X1  g717(.A1(new_n552), .A2(new_n566), .A3(new_n710), .ZN(new_n904));
  OAI21_X1  g718(.A(KEYINPUT110), .B1(new_n507), .B2(new_n904), .ZN(new_n905));
  NAND2_X1  g719(.A1(new_n903), .A2(new_n905), .ZN(new_n906));
  NOR2_X1   g720(.A1(new_n830), .A2(new_n906), .ZN(new_n907));
  NAND3_X1  g721(.A1(new_n682), .A2(new_n683), .A3(new_n907), .ZN(new_n908));
  OR2_X1    g722(.A1(new_n766), .A2(new_n779), .ZN(new_n909));
  NAND3_X1  g723(.A1(new_n908), .A2(new_n786), .A3(new_n909), .ZN(new_n910));
  NOR2_X1   g724(.A1(new_n910), .A2(new_n783), .ZN(new_n911));
  INV_X1    g725(.A(KEYINPUT53), .ZN(new_n912));
  NAND2_X1  g726(.A1(new_n689), .A2(new_n876), .ZN(new_n913));
  AOI21_X1  g727(.A(new_n912), .B1(new_n913), .B2(KEYINPUT52), .ZN(new_n914));
  NAND4_X1  g728(.A1(new_n886), .A2(new_n898), .A3(new_n911), .A4(new_n914), .ZN(new_n915));
  INV_X1    g729(.A(KEYINPUT54), .ZN(new_n916));
  NAND3_X1  g730(.A1(new_n628), .A2(new_n675), .A3(new_n891), .ZN(new_n917));
  INV_X1    g731(.A(KEYINPUT109), .ZN(new_n918));
  NAND2_X1  g732(.A1(new_n917), .A2(new_n918), .ZN(new_n919));
  NAND3_X1  g733(.A1(new_n889), .A2(KEYINPUT109), .A3(new_n891), .ZN(new_n920));
  NAND2_X1  g734(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  AND3_X1   g735(.A1(new_n764), .A2(new_n731), .A3(new_n727), .ZN(new_n922));
  NAND4_X1  g736(.A1(new_n921), .A2(new_n911), .A3(new_n745), .A4(new_n922), .ZN(new_n923));
  NAND2_X1  g737(.A1(new_n880), .A2(new_n885), .ZN(new_n924));
  OAI21_X1  g738(.A(new_n912), .B1(new_n923), .B2(new_n924), .ZN(new_n925));
  NAND3_X1  g739(.A1(new_n915), .A2(new_n916), .A3(new_n925), .ZN(new_n926));
  NAND2_X1  g740(.A1(new_n926), .A2(KEYINPUT111), .ZN(new_n927));
  AND4_X1   g741(.A1(new_n745), .A2(new_n921), .A3(new_n911), .A4(new_n922), .ZN(new_n928));
  AOI21_X1  g742(.A(KEYINPUT53), .B1(new_n928), .B2(new_n886), .ZN(new_n929));
  AOI21_X1  g743(.A(KEYINPUT53), .B1(new_n913), .B2(KEYINPUT52), .ZN(new_n930));
  NOR3_X1   g744(.A1(new_n923), .A2(new_n924), .A3(new_n930), .ZN(new_n931));
  OAI21_X1  g745(.A(KEYINPUT54), .B1(new_n929), .B2(new_n931), .ZN(new_n932));
  INV_X1    g746(.A(KEYINPUT111), .ZN(new_n933));
  NAND4_X1  g747(.A1(new_n915), .A2(new_n925), .A3(new_n933), .A4(new_n916), .ZN(new_n934));
  NAND3_X1  g748(.A1(new_n927), .A2(new_n932), .A3(new_n934), .ZN(new_n935));
  OAI22_X1  g749(.A1(new_n875), .A2(new_n935), .B1(G952), .B2(G953), .ZN(new_n936));
  XNOR2_X1  g750(.A(new_n723), .B(KEYINPUT49), .ZN(new_n937));
  NOR2_X1   g751(.A1(new_n649), .A2(new_n623), .ZN(new_n938));
  AND3_X1   g752(.A1(new_n937), .A2(new_n754), .A3(new_n938), .ZN(new_n939));
  NAND4_X1  g753(.A1(new_n939), .A2(new_n707), .A3(new_n847), .A4(new_n805), .ZN(new_n940));
  NAND2_X1  g754(.A1(new_n936), .A2(new_n940), .ZN(G75));
  OR3_X1    g755(.A1(new_n352), .A2(KEYINPUT118), .A3(G952), .ZN(new_n942));
  OAI21_X1  g756(.A(KEYINPUT118), .B1(new_n352), .B2(G952), .ZN(new_n943));
  NAND2_X1  g757(.A1(new_n942), .A2(new_n943), .ZN(new_n944));
  XNOR2_X1  g758(.A(new_n944), .B(KEYINPUT119), .ZN(new_n945));
  INV_X1    g759(.A(new_n945), .ZN(new_n946));
  AOI21_X1  g760(.A(new_n324), .B1(new_n915), .B2(new_n925), .ZN(new_n947));
  AOI21_X1  g761(.A(KEYINPUT56), .B1(new_n947), .B2(G210), .ZN(new_n948));
  AND2_X1   g762(.A1(new_n588), .A2(new_n595), .ZN(new_n949));
  XNOR2_X1  g763(.A(new_n949), .B(new_n593), .ZN(new_n950));
  XNOR2_X1  g764(.A(new_n950), .B(KEYINPUT55), .ZN(new_n951));
  INV_X1    g765(.A(new_n951), .ZN(new_n952));
  OAI21_X1  g766(.A(new_n946), .B1(new_n948), .B2(new_n952), .ZN(new_n953));
  AOI21_X1  g767(.A(new_n953), .B1(new_n948), .B2(new_n952), .ZN(G51));
  INV_X1    g768(.A(new_n914), .ZN(new_n955));
  NOR3_X1   g769(.A1(new_n923), .A2(new_n924), .A3(new_n955), .ZN(new_n956));
  OAI21_X1  g770(.A(KEYINPUT54), .B1(new_n929), .B2(new_n956), .ZN(new_n957));
  INV_X1    g771(.A(KEYINPUT120), .ZN(new_n958));
  NAND3_X1  g772(.A1(new_n957), .A2(new_n958), .A3(new_n926), .ZN(new_n959));
  NAND2_X1  g773(.A1(new_n915), .A2(new_n925), .ZN(new_n960));
  NAND3_X1  g774(.A1(new_n960), .A2(KEYINPUT120), .A3(KEYINPUT54), .ZN(new_n961));
  XOR2_X1   g775(.A(new_n772), .B(KEYINPUT57), .Z(new_n962));
  NAND3_X1  g776(.A1(new_n959), .A2(new_n961), .A3(new_n962), .ZN(new_n963));
  NAND2_X1  g777(.A1(new_n963), .A2(new_n720), .ZN(new_n964));
  XOR2_X1   g778(.A(new_n793), .B(KEYINPUT121), .Z(new_n965));
  NAND2_X1  g779(.A1(new_n947), .A2(new_n965), .ZN(new_n966));
  AOI21_X1  g780(.A(new_n944), .B1(new_n964), .B2(new_n966), .ZN(G54));
  NAND2_X1  g781(.A1(KEYINPUT58), .A2(G475), .ZN(new_n968));
  INV_X1    g782(.A(new_n968), .ZN(new_n969));
  NAND2_X1  g783(.A1(new_n947), .A2(new_n969), .ZN(new_n970));
  OAI21_X1  g784(.A(new_n970), .B1(new_n491), .B2(new_n472), .ZN(new_n971));
  NAND3_X1  g785(.A1(new_n947), .A2(new_n484), .A3(new_n969), .ZN(new_n972));
  AOI21_X1  g786(.A(new_n944), .B1(new_n971), .B2(new_n972), .ZN(G60));
  NAND2_X1  g787(.A1(G478), .A2(G902), .ZN(new_n974));
  XNOR2_X1  g788(.A(new_n974), .B(KEYINPUT59), .ZN(new_n975));
  NAND2_X1  g789(.A1(new_n935), .A2(new_n975), .ZN(new_n976));
  NAND2_X1  g790(.A1(new_n976), .A2(new_n637), .ZN(new_n977));
  INV_X1    g791(.A(KEYINPUT122), .ZN(new_n978));
  INV_X1    g792(.A(new_n637), .ZN(new_n979));
  AND2_X1   g793(.A1(new_n979), .A2(new_n975), .ZN(new_n980));
  NAND3_X1  g794(.A1(new_n959), .A2(new_n961), .A3(new_n980), .ZN(new_n981));
  NAND4_X1  g795(.A1(new_n977), .A2(new_n978), .A3(new_n946), .A4(new_n981), .ZN(new_n982));
  NAND2_X1  g796(.A1(new_n981), .A2(new_n946), .ZN(new_n983));
  AOI21_X1  g797(.A(new_n979), .B1(new_n935), .B2(new_n975), .ZN(new_n984));
  OAI21_X1  g798(.A(KEYINPUT122), .B1(new_n983), .B2(new_n984), .ZN(new_n985));
  NAND2_X1  g799(.A1(new_n982), .A2(new_n985), .ZN(G63));
  NAND2_X1  g800(.A1(G217), .A2(G902), .ZN(new_n987));
  XNOR2_X1  g801(.A(new_n987), .B(KEYINPUT123), .ZN(new_n988));
  XNOR2_X1  g802(.A(new_n988), .B(KEYINPUT60), .ZN(new_n989));
  AND2_X1   g803(.A1(new_n960), .A2(new_n989), .ZN(new_n990));
  OR2_X1    g804(.A1(new_n990), .A2(new_n357), .ZN(new_n991));
  NAND2_X1  g805(.A1(new_n990), .A2(new_n671), .ZN(new_n992));
  NAND3_X1  g806(.A1(new_n991), .A2(new_n946), .A3(new_n992), .ZN(new_n993));
  INV_X1    g807(.A(KEYINPUT61), .ZN(new_n994));
  NAND2_X1  g808(.A1(new_n993), .A2(new_n994), .ZN(new_n995));
  NAND4_X1  g809(.A1(new_n991), .A2(KEYINPUT61), .A3(new_n946), .A4(new_n992), .ZN(new_n996));
  NAND2_X1  g810(.A1(new_n995), .A2(new_n996), .ZN(G66));
  INV_X1    g811(.A(new_n561), .ZN(new_n998));
  AOI21_X1  g812(.A(new_n352), .B1(new_n998), .B2(G224), .ZN(new_n999));
  INV_X1    g813(.A(new_n898), .ZN(new_n1000));
  AOI21_X1  g814(.A(new_n999), .B1(new_n1000), .B2(new_n352), .ZN(new_n1001));
  INV_X1    g815(.A(G898), .ZN(new_n1002));
  AOI21_X1  g816(.A(new_n949), .B1(new_n1002), .B2(G953), .ZN(new_n1003));
  XNOR2_X1  g817(.A(new_n1001), .B(new_n1003), .ZN(G69));
  INV_X1    g818(.A(G900), .ZN(new_n1005));
  OAI21_X1  g819(.A(G953), .B1(new_n400), .B2(new_n1005), .ZN(new_n1006));
  XOR2_X1   g820(.A(new_n1006), .B(KEYINPUT124), .Z(new_n1007));
  INV_X1    g821(.A(new_n1007), .ZN(new_n1008));
  INV_X1    g822(.A(KEYINPUT125), .ZN(new_n1009));
  NAND3_X1  g823(.A1(new_n708), .A2(new_n716), .A3(new_n883), .ZN(new_n1010));
  INV_X1    g824(.A(KEYINPUT62), .ZN(new_n1011));
  XNOR2_X1  g825(.A(new_n1010), .B(new_n1011), .ZN(new_n1012));
  AOI21_X1  g826(.A(new_n692), .B1(new_n640), .B2(new_n657), .ZN(new_n1013));
  NAND3_X1  g827(.A1(new_n1013), .A2(new_n718), .A3(new_n771), .ZN(new_n1014));
  AND3_X1   g828(.A1(new_n1012), .A2(new_n815), .A3(new_n1014), .ZN(new_n1015));
  AOI21_X1  g829(.A(G953), .B1(new_n828), .B2(new_n1015), .ZN(new_n1016));
  NAND2_X1  g830(.A1(new_n314), .A2(new_n282), .ZN(new_n1017));
  XNOR2_X1  g831(.A(new_n1017), .B(new_n456), .ZN(new_n1018));
  INV_X1    g832(.A(new_n1018), .ZN(new_n1019));
  OAI21_X1  g833(.A(new_n1009), .B1(new_n1016), .B2(new_n1019), .ZN(new_n1020));
  AOI21_X1  g834(.A(new_n1018), .B1(G900), .B2(G953), .ZN(new_n1021));
  INV_X1    g835(.A(new_n1021), .ZN(new_n1022));
  NAND3_X1  g836(.A1(new_n802), .A2(new_n763), .A3(new_n836), .ZN(new_n1023));
  INV_X1    g837(.A(new_n783), .ZN(new_n1024));
  AND4_X1   g838(.A1(new_n716), .A2(new_n1024), .A3(new_n786), .A4(new_n883), .ZN(new_n1025));
  NAND3_X1  g839(.A1(new_n815), .A2(new_n1023), .A3(new_n1025), .ZN(new_n1026));
  AOI21_X1  g840(.A(new_n1026), .B1(new_n827), .B2(new_n825), .ZN(new_n1027));
  AOI21_X1  g841(.A(new_n1022), .B1(new_n1027), .B2(new_n352), .ZN(new_n1028));
  OAI21_X1  g842(.A(new_n1008), .B1(new_n1020), .B2(new_n1028), .ZN(new_n1029));
  NAND2_X1  g843(.A1(new_n1027), .A2(new_n352), .ZN(new_n1030));
  NAND2_X1  g844(.A1(new_n1030), .A2(new_n1021), .ZN(new_n1031));
  NAND3_X1  g845(.A1(new_n1012), .A2(new_n815), .A3(new_n1014), .ZN(new_n1032));
  AOI21_X1  g846(.A(new_n1032), .B1(new_n827), .B2(new_n825), .ZN(new_n1033));
  OAI21_X1  g847(.A(new_n1018), .B1(new_n1033), .B2(G953), .ZN(new_n1034));
  NAND4_X1  g848(.A1(new_n1031), .A2(new_n1034), .A3(new_n1009), .A4(new_n1007), .ZN(new_n1035));
  AND2_X1   g849(.A1(new_n1029), .A2(new_n1035), .ZN(G72));
  NAND2_X1  g850(.A1(new_n315), .A2(new_n192), .ZN(new_n1037));
  XNOR2_X1  g851(.A(KEYINPUT126), .B(KEYINPUT63), .ZN(new_n1038));
  NAND2_X1  g852(.A1(G472), .A2(G902), .ZN(new_n1039));
  XNOR2_X1  g853(.A(new_n1038), .B(new_n1039), .ZN(new_n1040));
  INV_X1    g854(.A(new_n1040), .ZN(new_n1041));
  NOR2_X1   g855(.A1(new_n696), .A2(new_n1041), .ZN(new_n1042));
  OAI211_X1 g856(.A(new_n1037), .B(new_n1042), .C1(new_n929), .C2(new_n931), .ZN(new_n1043));
  AOI21_X1  g857(.A(new_n1041), .B1(new_n1033), .B2(new_n898), .ZN(new_n1044));
  INV_X1    g858(.A(new_n696), .ZN(new_n1045));
  OAI21_X1  g859(.A(new_n1043), .B1(new_n1044), .B2(new_n1045), .ZN(new_n1046));
  INV_X1    g860(.A(KEYINPUT127), .ZN(new_n1047));
  INV_X1    g861(.A(new_n1026), .ZN(new_n1048));
  NAND3_X1  g862(.A1(new_n828), .A2(new_n1048), .A3(new_n898), .ZN(new_n1049));
  AOI21_X1  g863(.A(new_n1037), .B1(new_n1049), .B2(new_n1040), .ZN(new_n1050));
  OAI21_X1  g864(.A(new_n1047), .B1(new_n1050), .B2(new_n944), .ZN(new_n1051));
  INV_X1    g865(.A(new_n944), .ZN(new_n1052));
  AOI21_X1  g866(.A(new_n1041), .B1(new_n1027), .B2(new_n898), .ZN(new_n1053));
  OAI211_X1 g867(.A(KEYINPUT127), .B(new_n1052), .C1(new_n1053), .C2(new_n1037), .ZN(new_n1054));
  AOI21_X1  g868(.A(new_n1046), .B1(new_n1051), .B2(new_n1054), .ZN(G57));
endmodule


