

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357,
         n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368,
         n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379,
         n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390,
         n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
         n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412,
         n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423,
         n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
         n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445,
         n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456,
         n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467,
         n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478,
         n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489,
         n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500,
         n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511,
         n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589,
         n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, n600,
         n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, n611,
         n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, n622,
         n623, n624, n625, n626, n627, n628, n629, n630, n631, n632, n633,
         n634, n635, n636, n637, n638, n639, n640, n641, n642, n643, n644,
         n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, n655,
         n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666,
         n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, n677,
         n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688,
         n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n699,
         n700, n701, n702, n703, n704, n705, n706, n707, n708, n709, n710,
         n711, n712, n713, n714, n715, n716, n717, n718, n719, n720, n721,
         n722, n723, n724, n725, n726, n727, n728, n729, n730, n731, n732,
         n733, n734, n735, n736, n737, n738, n739, n740, n741, n742;

  INV_X1 U370 ( .A(n650), .ZN(n347) );
  BUF_X1 U371 ( .A(n548), .Z(n349) );
  NOR2_X1 U372 ( .A1(n549), .A2(n553), .ZN(n679) );
  XNOR2_X1 U373 ( .A(n596), .B(KEYINPUT1), .ZN(n548) );
  XNOR2_X1 U374 ( .A(n513), .B(n501), .ZN(n730) );
  INV_X1 U375 ( .A(n353), .ZN(n350) );
  XNOR2_X1 U376 ( .A(n499), .B(n500), .ZN(n513) );
  XNOR2_X1 U377 ( .A(n391), .B(G143), .ZN(n539) );
  XNOR2_X1 U378 ( .A(n392), .B(KEYINPUT90), .ZN(n552) );
  NAND2_X2 U379 ( .A1(n468), .A2(G210), .ZN(n354) );
  NAND2_X1 U380 ( .A1(n348), .A2(n347), .ZN(n380) );
  INV_X1 U381 ( .A(n629), .ZN(n348) );
  XOR2_X2 U382 ( .A(KEYINPUT72), .B(KEYINPUT34), .Z(n516) );
  NOR2_X1 U383 ( .A1(n351), .A2(n350), .ZN(n396) );
  INV_X1 U384 ( .A(n389), .ZN(n351) );
  INV_X1 U385 ( .A(G953), .ZN(n736) );
  XNOR2_X2 U386 ( .A(G128), .B(KEYINPUT65), .ZN(n391) );
  XNOR2_X2 U387 ( .A(n554), .B(KEYINPUT31), .ZN(n650) );
  NAND2_X2 U388 ( .A1(n541), .A2(n589), .ZN(n542) );
  NAND2_X2 U389 ( .A1(n396), .A2(n451), .ZN(n404) );
  XNOR2_X2 U390 ( .A(n464), .B(n463), .ZN(n454) );
  INV_X1 U391 ( .A(G146), .ZN(n502) );
  INV_X1 U392 ( .A(G116), .ZN(n463) );
  NOR2_X1 U393 ( .A1(n734), .A2(n435), .ZN(n434) );
  AND2_X2 U394 ( .A1(n552), .A2(n551), .ZN(n629) );
  XNOR2_X1 U395 ( .A(n549), .B(KEYINPUT6), .ZN(n583) );
  NOR2_X1 U396 ( .A1(n697), .A2(G902), .ZN(n507) );
  XNOR2_X1 U397 ( .A(n730), .B(n446), .ZN(n697) );
  XNOR2_X1 U398 ( .A(n505), .B(n504), .ZN(n446) );
  XNOR2_X1 U399 ( .A(n503), .B(n502), .ZN(n504) );
  XNOR2_X1 U400 ( .A(G122), .B(KEYINPUT16), .ZN(n453) );
  NAND2_X1 U401 ( .A1(n433), .A2(n395), .ZN(n352) );
  NAND2_X1 U402 ( .A1(n433), .A2(n395), .ZN(n432) );
  XNOR2_X1 U403 ( .A(G902), .B(KEYINPUT15), .ZN(n458) );
  XNOR2_X1 U404 ( .A(n405), .B(n436), .ZN(n621) );
  XNOR2_X1 U405 ( .A(n505), .B(n437), .ZN(n436) );
  XNOR2_X1 U406 ( .A(n715), .B(n498), .ZN(n405) );
  XNOR2_X1 U407 ( .A(n461), .B(n438), .ZN(n437) );
  XNOR2_X1 U408 ( .A(n481), .B(n419), .ZN(n729) );
  INV_X1 U409 ( .A(KEYINPUT10), .ZN(n419) );
  NAND2_X1 U410 ( .A1(n365), .A2(n359), .ZN(n734) );
  XNOR2_X1 U411 ( .A(n366), .B(n398), .ZN(n365) );
  INV_X1 U412 ( .A(n654), .ZN(n397) );
  INV_X1 U413 ( .A(KEYINPUT47), .ZN(n413) );
  INV_X1 U414 ( .A(KEYINPUT46), .ZN(n415) );
  XNOR2_X1 U415 ( .A(n539), .B(n355), .ZN(n499) );
  NOR2_X1 U416 ( .A1(n613), .A2(n448), .ZN(n447) );
  XNOR2_X1 U417 ( .A(n371), .B(G101), .ZN(n508) );
  INV_X1 U418 ( .A(KEYINPUT67), .ZN(n371) );
  NOR2_X2 U419 ( .A1(n564), .A2(n544), .ZN(n673) );
  XNOR2_X1 U420 ( .A(n495), .B(n494), .ZN(n668) );
  XNOR2_X1 U421 ( .A(n493), .B(KEYINPUT25), .ZN(n494) );
  XOR2_X1 U422 ( .A(KEYINPUT5), .B(KEYINPUT96), .Z(n512) );
  XNOR2_X1 U423 ( .A(G146), .B(G137), .ZN(n511) );
  XNOR2_X1 U424 ( .A(G134), .B(G131), .ZN(n500) );
  XNOR2_X1 U425 ( .A(KEYINPUT91), .B(KEYINPUT80), .ZN(n484) );
  XNOR2_X1 U426 ( .A(n501), .B(KEYINPUT93), .ZN(n482) );
  XOR2_X1 U427 ( .A(KEYINPUT23), .B(G110), .Z(n480) );
  XNOR2_X1 U428 ( .A(G107), .B(G134), .ZN(n531) );
  XNOR2_X1 U429 ( .A(G116), .B(G122), .ZN(n530) );
  XNOR2_X1 U430 ( .A(n443), .B(n441), .ZN(n703) );
  XNOR2_X1 U431 ( .A(n527), .B(n442), .ZN(n441) );
  XNOR2_X1 U432 ( .A(n526), .B(n523), .ZN(n442) );
  INV_X1 U433 ( .A(n734), .ZN(n395) );
  NOR2_X1 U434 ( .A1(n592), .A2(n579), .ZN(n580) );
  INV_X1 U435 ( .A(n543), .ZN(n556) );
  XNOR2_X1 U436 ( .A(KEYINPUT28), .B(KEYINPUT106), .ZN(n594) );
  INV_X1 U437 ( .A(KEYINPUT102), .ZN(n378) );
  XNOR2_X1 U438 ( .A(n542), .B(KEYINPUT35), .ZN(n377) );
  XNOR2_X1 U439 ( .A(n462), .B(n357), .ZN(n438) );
  XNOR2_X1 U440 ( .A(n420), .B(G146), .ZN(n481) );
  INV_X1 U441 ( .A(G125), .ZN(n420) );
  NOR2_X1 U442 ( .A1(G953), .A2(G237), .ZN(n525) );
  XNOR2_X1 U443 ( .A(n597), .B(n413), .ZN(n412) );
  INV_X1 U444 ( .A(KEYINPUT48), .ZN(n398) );
  XNOR2_X1 U445 ( .A(G113), .B(G131), .ZN(n523) );
  XNOR2_X1 U446 ( .A(G143), .B(G122), .ZN(n518) );
  XOR2_X1 U447 ( .A(G140), .B(G104), .Z(n519) );
  XOR2_X1 U448 ( .A(G137), .B(G140), .Z(n501) );
  NAND2_X1 U449 ( .A1(G237), .A2(G234), .ZN(n471) );
  XOR2_X1 U450 ( .A(KEYINPUT14), .B(KEYINPUT88), .Z(n472) );
  NOR2_X1 U451 ( .A1(G902), .A2(G237), .ZN(n467) );
  XOR2_X1 U452 ( .A(n590), .B(KEYINPUT38), .Z(n658) );
  NAND2_X1 U453 ( .A1(n466), .A2(n354), .ZN(n452) );
  XNOR2_X1 U454 ( .A(n528), .B(n439), .ZN(n543) );
  XNOR2_X1 U455 ( .A(n529), .B(n440), .ZN(n439) );
  INV_X1 U456 ( .A(G475), .ZN(n440) );
  NAND2_X1 U457 ( .A1(n543), .A2(n555), .ZN(n660) );
  XNOR2_X1 U458 ( .A(n459), .B(G110), .ZN(n713) );
  NAND2_X1 U459 ( .A1(n432), .A2(n430), .ZN(n429) );
  AND2_X1 U460 ( .A1(n434), .A2(n447), .ZN(n428) );
  XNOR2_X1 U461 ( .A(n460), .B(n713), .ZN(n505) );
  XNOR2_X1 U462 ( .A(n508), .B(KEYINPUT71), .ZN(n460) );
  XNOR2_X1 U463 ( .A(KEYINPUT104), .B(KEYINPUT33), .ZN(n444) );
  NAND2_X1 U464 ( .A1(n390), .A2(n583), .ZN(n445) );
  AND2_X1 U465 ( .A1(n548), .A2(n673), .ZN(n390) );
  XNOR2_X1 U466 ( .A(n369), .B(n368), .ZN(n619) );
  XNOR2_X1 U467 ( .A(n510), .B(n457), .ZN(n368) );
  XNOR2_X1 U468 ( .A(n513), .B(n370), .ZN(n369) );
  XNOR2_X1 U469 ( .A(G128), .B(G119), .ZN(n479) );
  XNOR2_X1 U470 ( .A(n539), .B(n538), .ZN(n614) );
  XNOR2_X1 U471 ( .A(n703), .B(n702), .ZN(n704) );
  NAND2_X1 U472 ( .A1(n426), .A2(n425), .ZN(n612) );
  INV_X1 U473 ( .A(KEYINPUT40), .ZN(n367) );
  XNOR2_X1 U474 ( .A(n422), .B(n421), .ZN(n644) );
  INV_X1 U475 ( .A(KEYINPUT78), .ZN(n421) );
  NOR2_X1 U476 ( .A1(n601), .A2(n407), .ZN(n422) );
  AND2_X1 U477 ( .A1(n452), .A2(n450), .ZN(n353) );
  XOR2_X1 U478 ( .A(KEYINPUT4), .B(KEYINPUT68), .Z(n355) );
  OR2_X1 U479 ( .A1(n466), .A2(n354), .ZN(n356) );
  XNOR2_X1 U480 ( .A(KEYINPUT17), .B(KEYINPUT77), .ZN(n357) );
  AND2_X1 U481 ( .A1(n451), .A2(n452), .ZN(n358) );
  AND2_X1 U482 ( .A1(n657), .A2(n397), .ZN(n359) );
  OR2_X1 U483 ( .A1(n548), .A2(n564), .ZN(n360) );
  OR2_X1 U484 ( .A1(n652), .A2(n641), .ZN(n361) );
  XOR2_X1 U485 ( .A(n619), .B(KEYINPUT62), .Z(n362) );
  XNOR2_X1 U486 ( .A(KEYINPUT64), .B(KEYINPUT45), .ZN(n363) );
  INV_X1 U487 ( .A(n610), .ZN(n435) );
  XOR2_X1 U488 ( .A(KEYINPUT85), .B(n616), .Z(n712) );
  INV_X1 U489 ( .A(n712), .ZN(n626) );
  XOR2_X1 U490 ( .A(n627), .B(KEYINPUT81), .Z(n364) );
  NAND2_X1 U491 ( .A1(n411), .A2(n414), .ZN(n366) );
  XNOR2_X1 U492 ( .A(n418), .B(G131), .ZN(G33) );
  XNOR2_X1 U493 ( .A(n599), .B(n367), .ZN(n418) );
  XNOR2_X1 U494 ( .A(n514), .B(n509), .ZN(n370) );
  NAND2_X1 U495 ( .A1(n376), .A2(n372), .ZN(n394) );
  XNOR2_X1 U496 ( .A(n373), .B(n378), .ZN(n372) );
  NAND2_X1 U497 ( .A1(n375), .A2(n374), .ZN(n373) );
  INV_X1 U498 ( .A(n628), .ZN(n374) );
  NAND2_X1 U499 ( .A1(n380), .A2(n379), .ZN(n375) );
  NAND2_X1 U500 ( .A1(n377), .A2(KEYINPUT44), .ZN(n376) );
  INV_X1 U501 ( .A(n662), .ZN(n379) );
  INV_X1 U502 ( .A(n499), .ZN(n498) );
  BUF_X1 U503 ( .A(n621), .Z(n381) );
  BUF_X1 U504 ( .A(n433), .Z(n382) );
  NAND2_X1 U505 ( .A1(n429), .A2(n427), .ZN(n383) );
  NOR2_X1 U506 ( .A1(n563), .A2(n384), .ZN(n628) );
  OR2_X1 U507 ( .A1(n583), .A2(n360), .ZN(n384) );
  NAND2_X1 U508 ( .A1(n429), .A2(n427), .ZN(n701) );
  XNOR2_X1 U509 ( .A(n542), .B(KEYINPUT35), .ZN(n385) );
  NAND2_X1 U510 ( .A1(n381), .A2(n354), .ZN(n386) );
  BUF_X1 U511 ( .A(n383), .Z(n708) );
  BUF_X1 U512 ( .A(n424), .Z(n407) );
  NOR2_X1 U513 ( .A1(n431), .A2(n610), .ZN(n430) );
  XNOR2_X1 U514 ( .A(n416), .B(n415), .ZN(n414) );
  NAND2_X1 U515 ( .A1(n387), .A2(n578), .ZN(n592) );
  XNOR2_X1 U516 ( .A(n573), .B(KEYINPUT30), .ZN(n387) );
  NAND2_X1 U517 ( .A1(n621), .A2(n354), .ZN(n389) );
  XNOR2_X2 U518 ( .A(n388), .B(n363), .ZN(n433) );
  NAND2_X1 U519 ( .A1(n399), .A2(n401), .ZN(n388) );
  NAND2_X1 U520 ( .A1(n428), .A2(n433), .ZN(n427) );
  NOR2_X1 U521 ( .A1(n617), .A2(n712), .ZN(n618) );
  NOR2_X1 U522 ( .A1(n706), .A2(n712), .ZN(n408) );
  NAND2_X1 U523 ( .A1(n358), .A2(n386), .ZN(n608) );
  XNOR2_X2 U524 ( .A(n515), .B(G472), .ZN(n549) );
  XNOR2_X2 U525 ( .A(n507), .B(n506), .ZN(n596) );
  NAND2_X1 U526 ( .A1(n392), .A2(n679), .ZN(n554) );
  AND2_X1 U527 ( .A1(n392), .A2(n545), .ZN(n547) );
  XNOR2_X2 U528 ( .A(n478), .B(KEYINPUT0), .ZN(n392) );
  NAND2_X1 U529 ( .A1(n393), .A2(n568), .ZN(n569) );
  XNOR2_X1 U530 ( .A(n394), .B(KEYINPUT83), .ZN(n393) );
  INV_X1 U531 ( .A(n382), .ZN(n724) );
  OR2_X1 U532 ( .A1(n621), .A2(n356), .ZN(n451) );
  XNOR2_X1 U533 ( .A(n569), .B(n400), .ZN(n399) );
  INV_X1 U534 ( .A(KEYINPUT82), .ZN(n400) );
  INV_X1 U535 ( .A(n572), .ZN(n401) );
  XNOR2_X2 U536 ( .A(n402), .B(n470), .ZN(n424) );
  NOR2_X1 U537 ( .A1(n603), .A2(n402), .ZN(n586) );
  XNOR2_X2 U538 ( .A(n404), .B(KEYINPUT84), .ZN(n402) );
  XNOR2_X1 U539 ( .A(n488), .B(n487), .ZN(n489) );
  NAND2_X1 U540 ( .A1(n383), .A2(G472), .ZN(n620) );
  XNOR2_X1 U541 ( .A(n403), .B(KEYINPUT63), .ZN(G57) );
  NAND2_X1 U542 ( .A1(n406), .A2(n626), .ZN(n403) );
  NOR2_X1 U543 ( .A1(n563), .A2(n583), .ZN(n559) );
  XNOR2_X1 U544 ( .A(n620), .B(n362), .ZN(n406) );
  XNOR2_X1 U545 ( .A(n408), .B(n707), .ZN(G60) );
  XNOR2_X1 U546 ( .A(n409), .B(n364), .ZN(G51) );
  NAND2_X1 U547 ( .A1(n410), .A2(n626), .ZN(n409) );
  XNOR2_X1 U548 ( .A(n625), .B(n624), .ZN(n410) );
  NOR2_X1 U549 ( .A1(n412), .A2(n361), .ZN(n411) );
  NAND2_X1 U550 ( .A1(n418), .A2(n417), .ZN(n416) );
  INV_X1 U551 ( .A(n742), .ZN(n417) );
  NAND2_X1 U552 ( .A1(n423), .A2(n596), .ZN(n601) );
  XNOR2_X1 U553 ( .A(n595), .B(n594), .ZN(n423) );
  NOR2_X2 U554 ( .A1(n424), .A2(n477), .ZN(n478) );
  NAND2_X1 U555 ( .A1(n382), .A2(n434), .ZN(n425) );
  NAND2_X1 U556 ( .A1(n352), .A2(n435), .ZN(n426) );
  INV_X1 U557 ( .A(n447), .ZN(n431) );
  XNOR2_X1 U558 ( .A(n729), .B(n482), .ZN(n488) );
  XNOR2_X1 U559 ( .A(n524), .B(n729), .ZN(n443) );
  NAND2_X1 U560 ( .A1(n552), .A2(n687), .ZN(n517) );
  XNOR2_X2 U561 ( .A(n445), .B(n444), .ZN(n687) );
  NAND2_X1 U562 ( .A1(n612), .A2(n611), .ZN(n449) );
  INV_X1 U563 ( .A(n611), .ZN(n448) );
  NAND2_X1 U564 ( .A1(n449), .A2(n692), .ZN(n693) );
  INV_X1 U565 ( .A(n604), .ZN(n450) );
  XNOR2_X2 U566 ( .A(n514), .B(n453), .ZN(n715) );
  XNOR2_X2 U567 ( .A(n454), .B(n465), .ZN(n514) );
  XNOR2_X1 U568 ( .A(n699), .B(n698), .ZN(n700) );
  XNOR2_X2 U569 ( .A(G113), .B(KEYINPUT3), .ZN(n464) );
  XOR2_X1 U570 ( .A(n485), .B(n484), .Z(n455) );
  XOR2_X1 U571 ( .A(n696), .B(n695), .Z(n456) );
  XOR2_X1 U572 ( .A(n512), .B(n511), .Z(n457) );
  INV_X1 U573 ( .A(KEYINPUT19), .ZN(n470) );
  XNOR2_X1 U574 ( .A(n486), .B(n455), .ZN(n487) );
  XNOR2_X1 U575 ( .A(n705), .B(n704), .ZN(n706) );
  INV_X1 U576 ( .A(KEYINPUT56), .ZN(n627) );
  XNOR2_X1 U577 ( .A(n458), .B(KEYINPUT86), .ZN(n613) );
  INV_X1 U578 ( .A(n613), .ZN(n466) );
  XNOR2_X1 U579 ( .A(G107), .B(G104), .ZN(n459) );
  XNOR2_X1 U580 ( .A(n481), .B(KEYINPUT18), .ZN(n461) );
  NAND2_X1 U581 ( .A1(G224), .A2(n736), .ZN(n462) );
  XOR2_X1 U582 ( .A(KEYINPUT70), .B(G119), .Z(n465) );
  XOR2_X1 U583 ( .A(KEYINPUT74), .B(n467), .Z(n468) );
  NAND2_X1 U584 ( .A1(G214), .A2(n468), .ZN(n469) );
  XNOR2_X1 U585 ( .A(n469), .B(KEYINPUT87), .ZN(n604) );
  XOR2_X1 U586 ( .A(n472), .B(n471), .Z(n474) );
  NAND2_X1 U587 ( .A1(n474), .A2(G952), .ZN(n473) );
  XOR2_X1 U588 ( .A(KEYINPUT89), .B(n473), .Z(n686) );
  NOR2_X1 U589 ( .A1(G953), .A2(n686), .ZN(n576) );
  AND2_X1 U590 ( .A1(n474), .A2(G953), .ZN(n475) );
  NAND2_X1 U591 ( .A1(G902), .A2(n475), .ZN(n574) );
  NOR2_X1 U592 ( .A1(n574), .A2(G898), .ZN(n476) );
  NOR2_X1 U593 ( .A1(n576), .A2(n476), .ZN(n477) );
  XNOR2_X1 U594 ( .A(n480), .B(n479), .ZN(n490) );
  NAND2_X1 U595 ( .A1(G234), .A2(n736), .ZN(n483) );
  XOR2_X1 U596 ( .A(KEYINPUT8), .B(n483), .Z(n535) );
  NAND2_X1 U597 ( .A1(G221), .A2(n535), .ZN(n486) );
  XOR2_X1 U598 ( .A(KEYINPUT92), .B(KEYINPUT24), .Z(n485) );
  XNOR2_X1 U599 ( .A(n490), .B(n489), .ZN(n710) );
  NOR2_X1 U600 ( .A1(n710), .A2(G902), .ZN(n495) );
  NAND2_X1 U601 ( .A1(n613), .A2(G234), .ZN(n492) );
  XNOR2_X1 U602 ( .A(KEYINPUT94), .B(KEYINPUT20), .ZN(n491) );
  XNOR2_X1 U603 ( .A(n492), .B(n491), .ZN(n496) );
  NAND2_X1 U604 ( .A1(n496), .A2(G217), .ZN(n493) );
  INV_X1 U605 ( .A(n668), .ZN(n564) );
  NAND2_X1 U606 ( .A1(G221), .A2(n496), .ZN(n497) );
  XOR2_X1 U607 ( .A(KEYINPUT21), .B(n497), .Z(n669) );
  XNOR2_X1 U608 ( .A(KEYINPUT95), .B(n669), .ZN(n544) );
  NAND2_X1 U609 ( .A1(G227), .A2(n736), .ZN(n503) );
  XNOR2_X1 U610 ( .A(KEYINPUT69), .B(G469), .ZN(n506) );
  XOR2_X1 U611 ( .A(n508), .B(KEYINPUT75), .Z(n510) );
  NAND2_X1 U612 ( .A1(n525), .A2(G210), .ZN(n509) );
  NOR2_X1 U613 ( .A1(n619), .A2(G902), .ZN(n515) );
  XNOR2_X1 U614 ( .A(n517), .B(n516), .ZN(n541) );
  XNOR2_X1 U615 ( .A(KEYINPUT100), .B(KEYINPUT13), .ZN(n529) );
  XNOR2_X1 U616 ( .A(n519), .B(n518), .ZN(n527) );
  XOR2_X1 U617 ( .A(KEYINPUT98), .B(KEYINPUT11), .Z(n521) );
  XNOR2_X1 U618 ( .A(KEYINPUT12), .B(KEYINPUT97), .ZN(n520) );
  XNOR2_X1 U619 ( .A(n521), .B(n520), .ZN(n522) );
  XOR2_X1 U620 ( .A(n522), .B(KEYINPUT99), .Z(n524) );
  NAND2_X1 U621 ( .A1(n525), .A2(G214), .ZN(n526) );
  NOR2_X1 U622 ( .A1(G902), .A2(n703), .ZN(n528) );
  XNOR2_X1 U623 ( .A(n530), .B(KEYINPUT101), .ZN(n534) );
  XOR2_X1 U624 ( .A(KEYINPUT7), .B(KEYINPUT9), .Z(n532) );
  XNOR2_X1 U625 ( .A(n532), .B(n531), .ZN(n533) );
  XOR2_X1 U626 ( .A(n534), .B(n533), .Z(n537) );
  NAND2_X1 U627 ( .A1(G217), .A2(n535), .ZN(n536) );
  XNOR2_X1 U628 ( .A(n537), .B(n536), .ZN(n538) );
  NOR2_X1 U629 ( .A1(G902), .A2(n614), .ZN(n540) );
  XNOR2_X1 U630 ( .A(G478), .B(n540), .ZN(n555) );
  NOR2_X1 U631 ( .A1(n543), .A2(n555), .ZN(n589) );
  NOR2_X1 U632 ( .A1(n660), .A2(n544), .ZN(n545) );
  XNOR2_X1 U633 ( .A(KEYINPUT22), .B(KEYINPUT73), .ZN(n546) );
  XNOR2_X1 U634 ( .A(n547), .B(n546), .ZN(n563) );
  NAND2_X1 U635 ( .A1(n596), .A2(n673), .ZN(n577) );
  INV_X1 U636 ( .A(n577), .ZN(n550) );
  AND2_X1 U637 ( .A1(n549), .A2(n550), .ZN(n551) );
  NAND2_X1 U638 ( .A1(n673), .A2(n548), .ZN(n553) );
  NAND2_X1 U639 ( .A1(n556), .A2(n555), .ZN(n643) );
  INV_X1 U640 ( .A(n643), .ZN(n647) );
  NOR2_X1 U641 ( .A1(n556), .A2(n555), .ZN(n649) );
  NOR2_X1 U642 ( .A1(n647), .A2(n649), .ZN(n662) );
  XNOR2_X1 U643 ( .A(KEYINPUT66), .B(KEYINPUT32), .ZN(n562) );
  NAND2_X1 U644 ( .A1(n564), .A2(n349), .ZN(n558) );
  XNOR2_X1 U645 ( .A(KEYINPUT103), .B(n558), .ZN(n560) );
  NAND2_X1 U646 ( .A1(n560), .A2(n559), .ZN(n561) );
  XNOR2_X1 U647 ( .A(n562), .B(n561), .ZN(n741) );
  INV_X1 U648 ( .A(n349), .ZN(n588) );
  BUF_X1 U649 ( .A(n563), .Z(n566) );
  NAND2_X1 U650 ( .A1(n564), .A2(n549), .ZN(n565) );
  NOR2_X1 U651 ( .A1(n566), .A2(n565), .ZN(n567) );
  NAND2_X1 U652 ( .A1(n588), .A2(n567), .ZN(n635) );
  NAND2_X1 U653 ( .A1(n741), .A2(n635), .ZN(n570) );
  NAND2_X1 U654 ( .A1(KEYINPUT44), .A2(n570), .ZN(n568) );
  OR2_X1 U655 ( .A1(n570), .A2(n385), .ZN(n571) );
  NOR2_X1 U656 ( .A1(KEYINPUT44), .A2(n571), .ZN(n572) );
  NOR2_X1 U657 ( .A1(n604), .A2(n549), .ZN(n573) );
  NOR2_X1 U658 ( .A1(G900), .A2(n574), .ZN(n575) );
  NOR2_X1 U659 ( .A1(n576), .A2(n575), .ZN(n581) );
  NOR2_X1 U660 ( .A1(n581), .A2(n577), .ZN(n578) );
  INV_X1 U661 ( .A(n608), .ZN(n590) );
  INV_X1 U662 ( .A(n658), .ZN(n579) );
  XNOR2_X1 U663 ( .A(n580), .B(KEYINPUT39), .ZN(n598) );
  INV_X1 U664 ( .A(n649), .ZN(n637) );
  NOR2_X1 U665 ( .A1(n598), .A2(n637), .ZN(n654) );
  NOR2_X1 U666 ( .A1(n581), .A2(n668), .ZN(n582) );
  NAND2_X1 U667 ( .A1(n582), .A2(n669), .ZN(n593) );
  INV_X1 U668 ( .A(n583), .ZN(n584) );
  NOR2_X1 U669 ( .A1(n593), .A2(n584), .ZN(n585) );
  NAND2_X1 U670 ( .A1(n647), .A2(n585), .ZN(n603) );
  XOR2_X1 U671 ( .A(KEYINPUT36), .B(n586), .Z(n587) );
  NOR2_X1 U672 ( .A1(n588), .A2(n587), .ZN(n652) );
  NAND2_X1 U673 ( .A1(n590), .A2(n589), .ZN(n591) );
  NOR2_X1 U674 ( .A1(n592), .A2(n591), .ZN(n641) );
  NOR2_X1 U675 ( .A1(n593), .A2(n549), .ZN(n595) );
  NOR2_X1 U676 ( .A1(n644), .A2(n662), .ZN(n597) );
  NOR2_X1 U677 ( .A1(n598), .A2(n643), .ZN(n599) );
  NAND2_X1 U678 ( .A1(n658), .A2(n450), .ZN(n661) );
  NOR2_X1 U679 ( .A1(n660), .A2(n661), .ZN(n600) );
  XNOR2_X1 U680 ( .A(n600), .B(KEYINPUT41), .ZN(n688) );
  NOR2_X1 U681 ( .A1(n601), .A2(n688), .ZN(n602) );
  XNOR2_X1 U682 ( .A(n602), .B(KEYINPUT42), .ZN(n742) );
  XNOR2_X1 U683 ( .A(KEYINPUT105), .B(KEYINPUT43), .ZN(n607) );
  OR2_X1 U684 ( .A1(n349), .A2(n603), .ZN(n605) );
  NOR2_X1 U685 ( .A1(n605), .A2(n604), .ZN(n606) );
  XNOR2_X1 U686 ( .A(n607), .B(n606), .ZN(n609) );
  NAND2_X1 U687 ( .A1(n609), .A2(n608), .ZN(n657) );
  NAND2_X1 U688 ( .A1(KEYINPUT2), .A2(KEYINPUT76), .ZN(n610) );
  OR2_X1 U689 ( .A1(KEYINPUT2), .A2(KEYINPUT76), .ZN(n611) );
  NAND2_X1 U690 ( .A1(n701), .A2(G478), .ZN(n615) );
  XNOR2_X1 U691 ( .A(n615), .B(n614), .ZN(n617) );
  NOR2_X1 U692 ( .A1(G952), .A2(n736), .ZN(n616) );
  XNOR2_X1 U693 ( .A(n618), .B(KEYINPUT122), .ZN(G63) );
  NAND2_X1 U694 ( .A1(n383), .A2(G210), .ZN(n625) );
  XOR2_X1 U695 ( .A(KEYINPUT54), .B(KEYINPUT55), .Z(n623) );
  XNOR2_X1 U696 ( .A(n381), .B(KEYINPUT79), .ZN(n622) );
  XNOR2_X1 U697 ( .A(n623), .B(n622), .ZN(n624) );
  XOR2_X1 U698 ( .A(n628), .B(G101), .Z(G3) );
  NAND2_X1 U699 ( .A1(n629), .A2(n647), .ZN(n630) );
  XNOR2_X1 U700 ( .A(n630), .B(G104), .ZN(G6) );
  XOR2_X1 U701 ( .A(KEYINPUT26), .B(KEYINPUT107), .Z(n632) );
  NAND2_X1 U702 ( .A1(n629), .A2(n649), .ZN(n631) );
  XNOR2_X1 U703 ( .A(n632), .B(n631), .ZN(n634) );
  XOR2_X1 U704 ( .A(G107), .B(KEYINPUT27), .Z(n633) );
  XNOR2_X1 U705 ( .A(n634), .B(n633), .ZN(G9) );
  XNOR2_X1 U706 ( .A(G110), .B(KEYINPUT108), .ZN(n636) );
  XNOR2_X1 U707 ( .A(n636), .B(n635), .ZN(G12) );
  NOR2_X1 U708 ( .A1(n644), .A2(n637), .ZN(n639) );
  XNOR2_X1 U709 ( .A(KEYINPUT109), .B(KEYINPUT29), .ZN(n638) );
  XNOR2_X1 U710 ( .A(n639), .B(n638), .ZN(n640) );
  XOR2_X1 U711 ( .A(G128), .B(n640), .Z(G30) );
  XOR2_X1 U712 ( .A(G143), .B(n641), .Z(n642) );
  XNOR2_X1 U713 ( .A(KEYINPUT110), .B(n642), .ZN(G45) );
  NOR2_X1 U714 ( .A1(n644), .A2(n643), .ZN(n646) );
  XNOR2_X1 U715 ( .A(G146), .B(KEYINPUT111), .ZN(n645) );
  XNOR2_X1 U716 ( .A(n646), .B(n645), .ZN(G48) );
  NAND2_X1 U717 ( .A1(n650), .A2(n647), .ZN(n648) );
  XNOR2_X1 U718 ( .A(n648), .B(G113), .ZN(G15) );
  NAND2_X1 U719 ( .A1(n650), .A2(n649), .ZN(n651) );
  XNOR2_X1 U720 ( .A(n651), .B(G116), .ZN(G18) );
  XNOR2_X1 U721 ( .A(G125), .B(n652), .ZN(n653) );
  XNOR2_X1 U722 ( .A(n653), .B(KEYINPUT37), .ZN(G27) );
  XOR2_X1 U723 ( .A(G134), .B(n654), .Z(n655) );
  XNOR2_X1 U724 ( .A(KEYINPUT112), .B(n655), .ZN(G36) );
  XOR2_X1 U725 ( .A(G140), .B(KEYINPUT113), .Z(n656) );
  XNOR2_X1 U726 ( .A(n657), .B(n656), .ZN(G42) );
  NOR2_X1 U727 ( .A1(n658), .A2(n450), .ZN(n659) );
  NOR2_X1 U728 ( .A1(n660), .A2(n659), .ZN(n664) );
  NOR2_X1 U729 ( .A1(n662), .A2(n661), .ZN(n663) );
  NOR2_X1 U730 ( .A1(n664), .A2(n663), .ZN(n665) );
  XOR2_X1 U731 ( .A(KEYINPUT116), .B(n665), .Z(n666) );
  NAND2_X1 U732 ( .A1(n666), .A2(n687), .ZN(n667) );
  XNOR2_X1 U733 ( .A(n667), .B(KEYINPUT117), .ZN(n683) );
  NOR2_X1 U734 ( .A1(n669), .A2(n668), .ZN(n670) );
  XNOR2_X1 U735 ( .A(n670), .B(KEYINPUT49), .ZN(n671) );
  NAND2_X1 U736 ( .A1(n671), .A2(n549), .ZN(n672) );
  XNOR2_X1 U737 ( .A(KEYINPUT114), .B(n672), .ZN(n677) );
  NOR2_X1 U738 ( .A1(n673), .A2(n349), .ZN(n674) );
  XOR2_X1 U739 ( .A(KEYINPUT115), .B(n674), .Z(n675) );
  XNOR2_X1 U740 ( .A(n675), .B(KEYINPUT50), .ZN(n676) );
  NOR2_X1 U741 ( .A1(n677), .A2(n676), .ZN(n678) );
  NOR2_X1 U742 ( .A1(n679), .A2(n678), .ZN(n680) );
  XOR2_X1 U743 ( .A(KEYINPUT51), .B(n680), .Z(n681) );
  NOR2_X1 U744 ( .A1(n688), .A2(n681), .ZN(n682) );
  NOR2_X1 U745 ( .A1(n683), .A2(n682), .ZN(n684) );
  XNOR2_X1 U746 ( .A(n684), .B(KEYINPUT52), .ZN(n685) );
  NOR2_X1 U747 ( .A1(n686), .A2(n685), .ZN(n691) );
  INV_X1 U748 ( .A(n687), .ZN(n689) );
  NOR2_X1 U749 ( .A1(n689), .A2(n688), .ZN(n690) );
  NOR2_X1 U750 ( .A1(n691), .A2(n690), .ZN(n692) );
  NOR2_X1 U751 ( .A1(n693), .A2(G953), .ZN(n694) );
  XNOR2_X1 U752 ( .A(n694), .B(KEYINPUT53), .ZN(G75) );
  NAND2_X1 U753 ( .A1(n708), .A2(G469), .ZN(n699) );
  XOR2_X1 U754 ( .A(KEYINPUT118), .B(KEYINPUT119), .Z(n696) );
  XNOR2_X1 U755 ( .A(KEYINPUT58), .B(KEYINPUT57), .ZN(n695) );
  XNOR2_X1 U756 ( .A(n697), .B(n456), .ZN(n698) );
  NOR2_X1 U757 ( .A1(n712), .A2(n700), .ZN(G54) );
  NAND2_X1 U758 ( .A1(n701), .A2(G475), .ZN(n705) );
  XOR2_X1 U759 ( .A(KEYINPUT120), .B(KEYINPUT59), .Z(n702) );
  XOR2_X1 U760 ( .A(KEYINPUT60), .B(KEYINPUT121), .Z(n707) );
  NAND2_X1 U761 ( .A1(G217), .A2(n708), .ZN(n709) );
  XNOR2_X1 U762 ( .A(n710), .B(n709), .ZN(n711) );
  NOR2_X1 U763 ( .A1(n712), .A2(n711), .ZN(G66) );
  XNOR2_X1 U764 ( .A(n713), .B(G101), .ZN(n714) );
  XNOR2_X1 U765 ( .A(n714), .B(KEYINPUT124), .ZN(n716) );
  XNOR2_X1 U766 ( .A(n715), .B(n716), .ZN(n718) );
  NOR2_X1 U767 ( .A1(n736), .A2(G898), .ZN(n717) );
  NOR2_X1 U768 ( .A1(n718), .A2(n717), .ZN(n719) );
  XNOR2_X1 U769 ( .A(KEYINPUT125), .B(n719), .ZN(n728) );
  INV_X1 U770 ( .A(G898), .ZN(n723) );
  NAND2_X1 U771 ( .A1(G224), .A2(G953), .ZN(n720) );
  XNOR2_X1 U772 ( .A(n720), .B(KEYINPUT123), .ZN(n721) );
  XNOR2_X1 U773 ( .A(n721), .B(KEYINPUT61), .ZN(n722) );
  NOR2_X1 U774 ( .A1(n723), .A2(n722), .ZN(n726) );
  NOR2_X1 U775 ( .A1(G953), .A2(n724), .ZN(n725) );
  NOR2_X1 U776 ( .A1(n726), .A2(n725), .ZN(n727) );
  XNOR2_X1 U777 ( .A(n728), .B(n727), .ZN(G69) );
  XOR2_X1 U778 ( .A(n730), .B(n729), .Z(n735) );
  XNOR2_X1 U779 ( .A(G227), .B(n735), .ZN(n731) );
  XNOR2_X1 U780 ( .A(KEYINPUT126), .B(n731), .ZN(n732) );
  NOR2_X1 U781 ( .A1(n736), .A2(n732), .ZN(n733) );
  NAND2_X1 U782 ( .A1(n733), .A2(G900), .ZN(n739) );
  XNOR2_X1 U783 ( .A(n735), .B(n734), .ZN(n737) );
  NAND2_X1 U784 ( .A1(n737), .A2(n736), .ZN(n738) );
  NAND2_X1 U785 ( .A1(n739), .A2(n738), .ZN(n740) );
  XNOR2_X1 U786 ( .A(n740), .B(KEYINPUT127), .ZN(G72) );
  XOR2_X1 U787 ( .A(n385), .B(G122), .Z(G24) );
  XNOR2_X1 U788 ( .A(G119), .B(n741), .ZN(G21) );
  XOR2_X1 U789 ( .A(n742), .B(G137), .Z(G39) );
endmodule

