//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 1 0 0 0 1 0 0 1 0 1 1 0 0 1 1 0 0 1 1 0 1 0 0 0 0 0 1 0 0 0 1 1 0 0 0 0 1 0 1 1 1 0 0 0 0 1 0 1 1 1 1 0 0 0 0 1 1 1 0 1 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:34:51 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n527, new_n528, new_n529, new_n530, new_n531, new_n532,
    new_n533, new_n534, new_n535, new_n536, new_n537, new_n539, new_n540,
    new_n541, new_n542, new_n543, new_n544, new_n545, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n555, new_n556, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n572, new_n573, new_n574, new_n576, new_n577,
    new_n578, new_n579, new_n580, new_n581, new_n582, new_n583, new_n584,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n605, new_n606, new_n607, new_n610, new_n612,
    new_n613, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n898, new_n899, new_n900, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1179, new_n1180, new_n1181;
  BUF_X1    g000(.A(G452), .Z(G350));
  XNOR2_X1  g001(.A(KEYINPUT64), .B(G452), .ZN(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  XNOR2_X1  g014(.A(KEYINPUT65), .B(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n450));
  XNOR2_X1  g025(.A(new_n450), .B(KEYINPUT2), .ZN(new_n451));
  NOR4_X1   g026(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n452));
  NAND2_X1  g027(.A1(new_n451), .A2(new_n452), .ZN(G261));
  INV_X1    g028(.A(G261), .ZN(G325));
  INV_X1    g029(.A(new_n451), .ZN(new_n455));
  NAND2_X1  g030(.A1(new_n455), .A2(G2106), .ZN(new_n456));
  INV_X1    g031(.A(KEYINPUT66), .ZN(new_n457));
  INV_X1    g032(.A(G567), .ZN(new_n458));
  OAI22_X1  g033(.A1(new_n456), .A2(new_n457), .B1(new_n458), .B2(new_n452), .ZN(new_n459));
  AOI21_X1  g034(.A(new_n459), .B1(new_n457), .B2(new_n456), .ZN(G319));
  INV_X1    g035(.A(G2105), .ZN(new_n461));
  XNOR2_X1  g036(.A(KEYINPUT3), .B(G2104), .ZN(new_n462));
  NAND2_X1  g037(.A1(new_n462), .A2(G125), .ZN(new_n463));
  NAND2_X1  g038(.A1(G113), .A2(G2104), .ZN(new_n464));
  INV_X1    g039(.A(KEYINPUT67), .ZN(new_n465));
  XNOR2_X1  g040(.A(new_n464), .B(new_n465), .ZN(new_n466));
  AOI21_X1  g041(.A(new_n461), .B1(new_n463), .B2(new_n466), .ZN(new_n467));
  AND2_X1   g042(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n468));
  NOR2_X1   g043(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n469));
  OAI211_X1 g044(.A(G137), .B(new_n461), .C1(new_n468), .C2(new_n469), .ZN(new_n470));
  AND2_X1   g045(.A1(new_n461), .A2(G2104), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n471), .A2(G101), .ZN(new_n472));
  INV_X1    g047(.A(KEYINPUT68), .ZN(new_n473));
  NAND3_X1  g048(.A1(new_n470), .A2(new_n472), .A3(new_n473), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n470), .A2(new_n472), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n475), .A2(KEYINPUT68), .ZN(new_n476));
  AOI21_X1  g051(.A(new_n467), .B1(new_n474), .B2(new_n476), .ZN(G160));
  OAI21_X1  g052(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n478));
  INV_X1    g053(.A(G112), .ZN(new_n479));
  AOI21_X1  g054(.A(new_n478), .B1(new_n479), .B2(G2105), .ZN(new_n480));
  NOR2_X1   g055(.A1(new_n468), .A2(new_n469), .ZN(new_n481));
  NOR2_X1   g056(.A1(new_n481), .A2(new_n461), .ZN(new_n482));
  NAND2_X1  g057(.A1(new_n482), .A2(G124), .ZN(new_n483));
  XNOR2_X1  g058(.A(new_n483), .B(KEYINPUT69), .ZN(new_n484));
  NOR2_X1   g059(.A1(new_n481), .A2(G2105), .ZN(new_n485));
  AOI211_X1 g060(.A(new_n480), .B(new_n484), .C1(G136), .C2(new_n485), .ZN(G162));
  OAI21_X1  g061(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n487));
  INV_X1    g062(.A(G114), .ZN(new_n488));
  AOI21_X1  g063(.A(new_n487), .B1(new_n488), .B2(G2105), .ZN(new_n489));
  AND2_X1   g064(.A1(G126), .A2(G2105), .ZN(new_n490));
  OAI21_X1  g065(.A(new_n490), .B1(new_n468), .B2(new_n469), .ZN(new_n491));
  NAND2_X1  g066(.A1(new_n491), .A2(KEYINPUT70), .ZN(new_n492));
  INV_X1    g067(.A(KEYINPUT70), .ZN(new_n493));
  OAI211_X1 g068(.A(new_n493), .B(new_n490), .C1(new_n468), .C2(new_n469), .ZN(new_n494));
  AOI21_X1  g069(.A(new_n489), .B1(new_n492), .B2(new_n494), .ZN(new_n495));
  OAI211_X1 g070(.A(G138), .B(new_n461), .C1(new_n468), .C2(new_n469), .ZN(new_n496));
  NAND2_X1  g071(.A1(new_n496), .A2(KEYINPUT4), .ZN(new_n497));
  INV_X1    g072(.A(KEYINPUT4), .ZN(new_n498));
  NAND4_X1  g073(.A1(new_n462), .A2(new_n498), .A3(G138), .A4(new_n461), .ZN(new_n499));
  NAND2_X1  g074(.A1(new_n497), .A2(new_n499), .ZN(new_n500));
  AND3_X1   g075(.A1(new_n495), .A2(KEYINPUT71), .A3(new_n500), .ZN(new_n501));
  AOI21_X1  g076(.A(KEYINPUT71), .B1(new_n495), .B2(new_n500), .ZN(new_n502));
  NOR2_X1   g077(.A1(new_n501), .A2(new_n502), .ZN(G164));
  INV_X1    g078(.A(G62), .ZN(new_n504));
  OR2_X1    g079(.A1(KEYINPUT5), .A2(G543), .ZN(new_n505));
  NAND2_X1  g080(.A1(KEYINPUT5), .A2(G543), .ZN(new_n506));
  AOI21_X1  g081(.A(new_n504), .B1(new_n505), .B2(new_n506), .ZN(new_n507));
  NAND2_X1  g082(.A1(new_n507), .A2(KEYINPUT73), .ZN(new_n508));
  INV_X1    g083(.A(new_n508), .ZN(new_n509));
  NAND2_X1  g084(.A1(G75), .A2(G543), .ZN(new_n510));
  OAI21_X1  g085(.A(new_n510), .B1(new_n507), .B2(KEYINPUT73), .ZN(new_n511));
  OAI21_X1  g086(.A(G651), .B1(new_n509), .B2(new_n511), .ZN(new_n512));
  OR2_X1    g087(.A1(KEYINPUT6), .A2(G651), .ZN(new_n513));
  NAND2_X1  g088(.A1(KEYINPUT6), .A2(G651), .ZN(new_n514));
  AOI22_X1  g089(.A1(new_n513), .A2(new_n514), .B1(new_n505), .B2(new_n506), .ZN(new_n515));
  INV_X1    g090(.A(G543), .ZN(new_n516));
  AOI21_X1  g091(.A(new_n516), .B1(new_n513), .B2(new_n514), .ZN(new_n517));
  AOI22_X1  g092(.A1(new_n515), .A2(G88), .B1(new_n517), .B2(G50), .ZN(new_n518));
  INV_X1    g093(.A(KEYINPUT72), .ZN(new_n519));
  AND2_X1   g094(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  NOR2_X1   g095(.A1(new_n518), .A2(new_n519), .ZN(new_n521));
  OAI21_X1  g096(.A(new_n512), .B1(new_n520), .B2(new_n521), .ZN(new_n522));
  NAND2_X1  g097(.A1(new_n522), .A2(KEYINPUT74), .ZN(new_n523));
  INV_X1    g098(.A(KEYINPUT74), .ZN(new_n524));
  OAI211_X1 g099(.A(new_n524), .B(new_n512), .C1(new_n520), .C2(new_n521), .ZN(new_n525));
  NAND2_X1  g100(.A1(new_n523), .A2(new_n525), .ZN(G166));
  NAND2_X1  g101(.A1(new_n505), .A2(new_n506), .ZN(new_n527));
  INV_X1    g102(.A(new_n527), .ZN(new_n528));
  XNOR2_X1  g103(.A(KEYINPUT6), .B(G651), .ZN(new_n529));
  NAND2_X1  g104(.A1(new_n529), .A2(G89), .ZN(new_n530));
  NAND2_X1  g105(.A1(G63), .A2(G651), .ZN(new_n531));
  AOI21_X1  g106(.A(new_n528), .B1(new_n530), .B2(new_n531), .ZN(new_n532));
  NAND3_X1  g107(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n533));
  XNOR2_X1  g108(.A(new_n533), .B(KEYINPUT7), .ZN(new_n534));
  NAND2_X1  g109(.A1(new_n529), .A2(G543), .ZN(new_n535));
  XOR2_X1   g110(.A(KEYINPUT75), .B(G51), .Z(new_n536));
  OAI21_X1  g111(.A(new_n534), .B1(new_n535), .B2(new_n536), .ZN(new_n537));
  NOR2_X1   g112(.A1(new_n532), .A2(new_n537), .ZN(G168));
  AOI22_X1  g113(.A1(new_n527), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n539));
  INV_X1    g114(.A(G651), .ZN(new_n540));
  NOR2_X1   g115(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  NAND2_X1  g116(.A1(new_n527), .A2(new_n529), .ZN(new_n542));
  INV_X1    g117(.A(G90), .ZN(new_n543));
  INV_X1    g118(.A(G52), .ZN(new_n544));
  OAI22_X1  g119(.A1(new_n542), .A2(new_n543), .B1(new_n535), .B2(new_n544), .ZN(new_n545));
  NOR2_X1   g120(.A1(new_n541), .A2(new_n545), .ZN(G171));
  AOI22_X1  g121(.A1(new_n527), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n547));
  NOR2_X1   g122(.A1(new_n547), .A2(new_n540), .ZN(new_n548));
  XOR2_X1   g123(.A(KEYINPUT76), .B(G81), .Z(new_n549));
  INV_X1    g124(.A(G43), .ZN(new_n550));
  OAI22_X1  g125(.A1(new_n542), .A2(new_n549), .B1(new_n535), .B2(new_n550), .ZN(new_n551));
  NOR2_X1   g126(.A1(new_n548), .A2(new_n551), .ZN(new_n552));
  NAND2_X1  g127(.A1(new_n552), .A2(G860), .ZN(G153));
  NAND4_X1  g128(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g129(.A1(G1), .A2(G3), .ZN(new_n555));
  XNOR2_X1  g130(.A(new_n555), .B(KEYINPUT8), .ZN(new_n556));
  NAND4_X1  g131(.A1(G319), .A2(G483), .A3(G661), .A4(new_n556), .ZN(G188));
  INV_X1    g132(.A(KEYINPUT77), .ZN(new_n558));
  INV_X1    g133(.A(G91), .ZN(new_n559));
  OAI21_X1  g134(.A(new_n558), .B1(new_n542), .B2(new_n559), .ZN(new_n560));
  NAND3_X1  g135(.A1(new_n515), .A2(KEYINPUT77), .A3(G91), .ZN(new_n561));
  NAND2_X1  g136(.A1(G78), .A2(G543), .ZN(new_n562));
  INV_X1    g137(.A(G65), .ZN(new_n563));
  OAI21_X1  g138(.A(new_n562), .B1(new_n528), .B2(new_n563), .ZN(new_n564));
  AOI22_X1  g139(.A1(new_n560), .A2(new_n561), .B1(new_n564), .B2(G651), .ZN(new_n565));
  NAND2_X1  g140(.A1(new_n517), .A2(G53), .ZN(new_n566));
  XNOR2_X1  g141(.A(new_n566), .B(KEYINPUT9), .ZN(new_n567));
  NAND2_X1  g142(.A1(new_n565), .A2(new_n567), .ZN(G299));
  INV_X1    g143(.A(G171), .ZN(G301));
  INV_X1    g144(.A(G168), .ZN(G286));
  INV_X1    g145(.A(G166), .ZN(G303));
  NAND2_X1  g146(.A1(new_n515), .A2(G87), .ZN(new_n572));
  OAI21_X1  g147(.A(G651), .B1(new_n527), .B2(G74), .ZN(new_n573));
  NAND2_X1  g148(.A1(new_n517), .A2(G49), .ZN(new_n574));
  NAND3_X1  g149(.A1(new_n572), .A2(new_n573), .A3(new_n574), .ZN(G288));
  AOI22_X1  g150(.A1(new_n515), .A2(G86), .B1(new_n517), .B2(G48), .ZN(new_n576));
  INV_X1    g151(.A(G61), .ZN(new_n577));
  AOI21_X1  g152(.A(new_n577), .B1(new_n505), .B2(new_n506), .ZN(new_n578));
  NAND2_X1  g153(.A1(G73), .A2(G543), .ZN(new_n579));
  NAND2_X1  g154(.A1(new_n579), .A2(KEYINPUT78), .ZN(new_n580));
  INV_X1    g155(.A(KEYINPUT78), .ZN(new_n581));
  NAND3_X1  g156(.A1(new_n581), .A2(G73), .A3(G543), .ZN(new_n582));
  NAND2_X1  g157(.A1(new_n580), .A2(new_n582), .ZN(new_n583));
  OAI21_X1  g158(.A(G651), .B1(new_n578), .B2(new_n583), .ZN(new_n584));
  NAND2_X1  g159(.A1(new_n576), .A2(new_n584), .ZN(G305));
  NAND2_X1  g160(.A1(G72), .A2(G543), .ZN(new_n586));
  INV_X1    g161(.A(G60), .ZN(new_n587));
  OAI21_X1  g162(.A(new_n586), .B1(new_n528), .B2(new_n587), .ZN(new_n588));
  INV_X1    g163(.A(KEYINPUT79), .ZN(new_n589));
  AOI21_X1  g164(.A(new_n540), .B1(new_n588), .B2(new_n589), .ZN(new_n590));
  OAI21_X1  g165(.A(new_n590), .B1(new_n589), .B2(new_n588), .ZN(new_n591));
  AOI22_X1  g166(.A1(new_n515), .A2(G85), .B1(new_n517), .B2(G47), .ZN(new_n592));
  NAND2_X1  g167(.A1(new_n591), .A2(new_n592), .ZN(G290));
  NAND2_X1  g168(.A1(G301), .A2(G868), .ZN(new_n594));
  AND3_X1   g169(.A1(new_n527), .A2(new_n529), .A3(G92), .ZN(new_n595));
  XNOR2_X1  g170(.A(new_n595), .B(KEYINPUT10), .ZN(new_n596));
  NAND2_X1  g171(.A1(G79), .A2(G543), .ZN(new_n597));
  INV_X1    g172(.A(G66), .ZN(new_n598));
  OAI21_X1  g173(.A(new_n597), .B1(new_n528), .B2(new_n598), .ZN(new_n599));
  AOI22_X1  g174(.A1(new_n599), .A2(G651), .B1(G54), .B2(new_n517), .ZN(new_n600));
  NAND2_X1  g175(.A1(new_n596), .A2(new_n600), .ZN(new_n601));
  INV_X1    g176(.A(new_n601), .ZN(new_n602));
  OAI21_X1  g177(.A(new_n594), .B1(new_n602), .B2(G868), .ZN(G284));
  OAI21_X1  g178(.A(new_n594), .B1(new_n602), .B2(G868), .ZN(G321));
  NAND2_X1  g179(.A1(G286), .A2(G868), .ZN(new_n605));
  XNOR2_X1  g180(.A(new_n605), .B(KEYINPUT80), .ZN(new_n606));
  INV_X1    g181(.A(G299), .ZN(new_n607));
  OAI21_X1  g182(.A(new_n606), .B1(G868), .B2(new_n607), .ZN(G297));
  OAI21_X1  g183(.A(new_n606), .B1(G868), .B2(new_n607), .ZN(G280));
  XNOR2_X1  g184(.A(KEYINPUT81), .B(G559), .ZN(new_n610));
  OAI21_X1  g185(.A(new_n602), .B1(G860), .B2(new_n610), .ZN(G148));
  NAND2_X1  g186(.A1(new_n602), .A2(new_n610), .ZN(new_n612));
  NAND2_X1  g187(.A1(new_n612), .A2(G868), .ZN(new_n613));
  OAI21_X1  g188(.A(new_n613), .B1(G868), .B2(new_n552), .ZN(G323));
  XNOR2_X1  g189(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g190(.A1(new_n462), .A2(new_n471), .ZN(new_n616));
  XOR2_X1   g191(.A(KEYINPUT82), .B(KEYINPUT12), .Z(new_n617));
  XNOR2_X1  g192(.A(new_n616), .B(new_n617), .ZN(new_n618));
  XNOR2_X1  g193(.A(new_n618), .B(KEYINPUT13), .ZN(new_n619));
  INV_X1    g194(.A(G2100), .ZN(new_n620));
  OR2_X1    g195(.A1(new_n619), .A2(new_n620), .ZN(new_n621));
  NAND2_X1  g196(.A1(new_n619), .A2(new_n620), .ZN(new_n622));
  NAND2_X1  g197(.A1(new_n485), .A2(G135), .ZN(new_n623));
  NAND2_X1  g198(.A1(new_n482), .A2(G123), .ZN(new_n624));
  NOR2_X1   g199(.A1(new_n461), .A2(G111), .ZN(new_n625));
  OAI21_X1  g200(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n626));
  OAI211_X1 g201(.A(new_n623), .B(new_n624), .C1(new_n625), .C2(new_n626), .ZN(new_n627));
  XOR2_X1   g202(.A(new_n627), .B(G2096), .Z(new_n628));
  NAND3_X1  g203(.A1(new_n621), .A2(new_n622), .A3(new_n628), .ZN(G156));
  XNOR2_X1  g204(.A(KEYINPUT15), .B(G2435), .ZN(new_n630));
  XNOR2_X1  g205(.A(KEYINPUT83), .B(G2438), .ZN(new_n631));
  XNOR2_X1  g206(.A(new_n630), .B(new_n631), .ZN(new_n632));
  XNOR2_X1  g207(.A(G2427), .B(G2430), .ZN(new_n633));
  OR2_X1    g208(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  NAND2_X1  g209(.A1(new_n632), .A2(new_n633), .ZN(new_n635));
  NAND3_X1  g210(.A1(new_n634), .A2(KEYINPUT14), .A3(new_n635), .ZN(new_n636));
  XNOR2_X1  g211(.A(G2451), .B(G2454), .ZN(new_n637));
  XNOR2_X1  g212(.A(new_n637), .B(KEYINPUT16), .ZN(new_n638));
  XOR2_X1   g213(.A(G1341), .B(G1348), .Z(new_n639));
  XNOR2_X1  g214(.A(new_n638), .B(new_n639), .ZN(new_n640));
  XNOR2_X1  g215(.A(new_n636), .B(new_n640), .ZN(new_n641));
  XOR2_X1   g216(.A(G2443), .B(G2446), .Z(new_n642));
  OAI21_X1  g217(.A(G14), .B1(new_n641), .B2(new_n642), .ZN(new_n643));
  AOI21_X1  g218(.A(new_n643), .B1(new_n642), .B2(new_n641), .ZN(G401));
  XOR2_X1   g219(.A(G2072), .B(G2078), .Z(new_n645));
  XOR2_X1   g220(.A(KEYINPUT85), .B(KEYINPUT17), .Z(new_n646));
  XNOR2_X1  g221(.A(new_n645), .B(new_n646), .ZN(new_n647));
  XNOR2_X1  g222(.A(G2067), .B(G2678), .ZN(new_n648));
  INV_X1    g223(.A(new_n648), .ZN(new_n649));
  NOR2_X1   g224(.A1(new_n647), .A2(new_n649), .ZN(new_n650));
  INV_X1    g225(.A(KEYINPUT84), .ZN(new_n651));
  XOR2_X1   g226(.A(G2084), .B(G2090), .Z(new_n652));
  AOI21_X1  g227(.A(new_n652), .B1(new_n649), .B2(new_n645), .ZN(new_n653));
  AOI21_X1  g228(.A(new_n650), .B1(new_n651), .B2(new_n653), .ZN(new_n654));
  OAI21_X1  g229(.A(new_n654), .B1(new_n651), .B2(new_n653), .ZN(new_n655));
  INV_X1    g230(.A(new_n645), .ZN(new_n656));
  NAND3_X1  g231(.A1(new_n656), .A2(new_n652), .A3(new_n648), .ZN(new_n657));
  XOR2_X1   g232(.A(new_n657), .B(KEYINPUT18), .Z(new_n658));
  NAND3_X1  g233(.A1(new_n647), .A2(new_n652), .A3(new_n649), .ZN(new_n659));
  NAND3_X1  g234(.A1(new_n655), .A2(new_n658), .A3(new_n659), .ZN(new_n660));
  XOR2_X1   g235(.A(G2096), .B(G2100), .Z(new_n661));
  XNOR2_X1  g236(.A(new_n660), .B(new_n661), .ZN(G227));
  XOR2_X1   g237(.A(G1956), .B(G2474), .Z(new_n663));
  XNOR2_X1  g238(.A(new_n663), .B(KEYINPUT86), .ZN(new_n664));
  XNOR2_X1  g239(.A(G1961), .B(G1966), .ZN(new_n665));
  INV_X1    g240(.A(new_n665), .ZN(new_n666));
  NAND2_X1  g241(.A1(new_n664), .A2(new_n666), .ZN(new_n667));
  XNOR2_X1  g242(.A(G1971), .B(G1976), .ZN(new_n668));
  XNOR2_X1  g243(.A(new_n668), .B(KEYINPUT19), .ZN(new_n669));
  NOR2_X1   g244(.A1(new_n667), .A2(new_n669), .ZN(new_n670));
  XOR2_X1   g245(.A(new_n670), .B(KEYINPUT20), .Z(new_n671));
  NOR2_X1   g246(.A1(new_n664), .A2(new_n666), .ZN(new_n672));
  INV_X1    g247(.A(new_n672), .ZN(new_n673));
  NAND3_X1  g248(.A1(new_n673), .A2(new_n669), .A3(new_n667), .ZN(new_n674));
  OAI211_X1 g249(.A(new_n671), .B(new_n674), .C1(new_n669), .C2(new_n673), .ZN(new_n675));
  XNOR2_X1  g250(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n676));
  XNOR2_X1  g251(.A(new_n675), .B(new_n676), .ZN(new_n677));
  XNOR2_X1  g252(.A(G1991), .B(G1996), .ZN(new_n678));
  XNOR2_X1  g253(.A(new_n678), .B(KEYINPUT87), .ZN(new_n679));
  XNOR2_X1  g254(.A(new_n677), .B(new_n679), .ZN(new_n680));
  XNOR2_X1  g255(.A(G1981), .B(G1986), .ZN(new_n681));
  INV_X1    g256(.A(new_n681), .ZN(new_n682));
  OR2_X1    g257(.A1(new_n680), .A2(new_n682), .ZN(new_n683));
  NAND2_X1  g258(.A1(new_n680), .A2(new_n682), .ZN(new_n684));
  NAND2_X1  g259(.A1(new_n683), .A2(new_n684), .ZN(G229));
  MUX2_X1   g260(.A(G6), .B(G305), .S(G16), .Z(new_n686));
  XNOR2_X1  g261(.A(new_n686), .B(KEYINPUT32), .ZN(new_n687));
  INV_X1    g262(.A(G1981), .ZN(new_n688));
  XNOR2_X1  g263(.A(new_n687), .B(new_n688), .ZN(new_n689));
  INV_X1    g264(.A(G16), .ZN(new_n690));
  NAND2_X1  g265(.A1(new_n690), .A2(G22), .ZN(new_n691));
  OAI21_X1  g266(.A(new_n691), .B1(G166), .B2(new_n690), .ZN(new_n692));
  OR2_X1    g267(.A1(new_n692), .A2(G1971), .ZN(new_n693));
  NAND2_X1  g268(.A1(new_n692), .A2(G1971), .ZN(new_n694));
  NOR2_X1   g269(.A1(G16), .A2(G23), .ZN(new_n695));
  XNOR2_X1  g270(.A(new_n695), .B(KEYINPUT88), .ZN(new_n696));
  OAI21_X1  g271(.A(new_n696), .B1(G288), .B2(new_n690), .ZN(new_n697));
  XOR2_X1   g272(.A(new_n697), .B(KEYINPUT33), .Z(new_n698));
  XNOR2_X1  g273(.A(new_n698), .B(G1976), .ZN(new_n699));
  NAND4_X1  g274(.A1(new_n689), .A2(new_n693), .A3(new_n694), .A4(new_n699), .ZN(new_n700));
  OR2_X1    g275(.A1(new_n700), .A2(KEYINPUT34), .ZN(new_n701));
  NAND2_X1  g276(.A1(new_n700), .A2(KEYINPUT34), .ZN(new_n702));
  MUX2_X1   g277(.A(G24), .B(G290), .S(G16), .Z(new_n703));
  AND2_X1   g278(.A1(new_n703), .A2(G1986), .ZN(new_n704));
  NOR2_X1   g279(.A1(new_n703), .A2(G1986), .ZN(new_n705));
  NAND2_X1  g280(.A1(new_n485), .A2(G131), .ZN(new_n706));
  NAND2_X1  g281(.A1(new_n482), .A2(G119), .ZN(new_n707));
  NOR2_X1   g282(.A1(new_n461), .A2(G107), .ZN(new_n708));
  OAI21_X1  g283(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n709));
  OAI211_X1 g284(.A(new_n706), .B(new_n707), .C1(new_n708), .C2(new_n709), .ZN(new_n710));
  MUX2_X1   g285(.A(G25), .B(new_n710), .S(G29), .Z(new_n711));
  XOR2_X1   g286(.A(KEYINPUT35), .B(G1991), .Z(new_n712));
  INV_X1    g287(.A(new_n712), .ZN(new_n713));
  XNOR2_X1  g288(.A(new_n711), .B(new_n713), .ZN(new_n714));
  NOR3_X1   g289(.A1(new_n704), .A2(new_n705), .A3(new_n714), .ZN(new_n715));
  NAND3_X1  g290(.A1(new_n701), .A2(new_n702), .A3(new_n715), .ZN(new_n716));
  XOR2_X1   g291(.A(new_n716), .B(KEYINPUT36), .Z(new_n717));
  AOI22_X1  g292(.A1(new_n485), .A2(G141), .B1(G105), .B2(new_n471), .ZN(new_n718));
  NAND2_X1  g293(.A1(new_n482), .A2(G129), .ZN(new_n719));
  NAND3_X1  g294(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n720));
  XOR2_X1   g295(.A(new_n720), .B(KEYINPUT26), .Z(new_n721));
  NAND3_X1  g296(.A1(new_n718), .A2(new_n719), .A3(new_n721), .ZN(new_n722));
  OR2_X1    g297(.A1(new_n722), .A2(KEYINPUT92), .ZN(new_n723));
  NAND2_X1  g298(.A1(new_n722), .A2(KEYINPUT92), .ZN(new_n724));
  NAND2_X1  g299(.A1(new_n723), .A2(new_n724), .ZN(new_n725));
  INV_X1    g300(.A(new_n725), .ZN(new_n726));
  INV_X1    g301(.A(G29), .ZN(new_n727));
  NOR2_X1   g302(.A1(new_n726), .A2(new_n727), .ZN(new_n728));
  AOI21_X1  g303(.A(new_n728), .B1(new_n727), .B2(G32), .ZN(new_n729));
  XOR2_X1   g304(.A(KEYINPUT27), .B(G1996), .Z(new_n730));
  XNOR2_X1  g305(.A(new_n730), .B(KEYINPUT93), .ZN(new_n731));
  NAND2_X1  g306(.A1(new_n729), .A2(new_n731), .ZN(new_n732));
  XOR2_X1   g307(.A(new_n732), .B(KEYINPUT94), .Z(new_n733));
  NAND2_X1  g308(.A1(new_n727), .A2(G27), .ZN(new_n734));
  OAI21_X1  g309(.A(new_n734), .B1(G164), .B2(new_n727), .ZN(new_n735));
  INV_X1    g310(.A(G2078), .ZN(new_n736));
  XNOR2_X1  g311(.A(new_n735), .B(new_n736), .ZN(new_n737));
  INV_X1    g312(.A(G2084), .ZN(new_n738));
  INV_X1    g313(.A(G34), .ZN(new_n739));
  AOI21_X1  g314(.A(G29), .B1(new_n739), .B2(KEYINPUT24), .ZN(new_n740));
  OAI21_X1  g315(.A(new_n740), .B1(KEYINPUT24), .B2(new_n739), .ZN(new_n741));
  INV_X1    g316(.A(G160), .ZN(new_n742));
  OAI21_X1  g317(.A(new_n741), .B1(new_n742), .B2(new_n727), .ZN(new_n743));
  OAI22_X1  g318(.A1(new_n729), .A2(new_n731), .B1(new_n738), .B2(new_n743), .ZN(new_n744));
  NAND2_X1  g319(.A1(new_n727), .A2(G33), .ZN(new_n745));
  NAND3_X1  g320(.A1(new_n461), .A2(G103), .A3(G2104), .ZN(new_n746));
  XNOR2_X1  g321(.A(new_n746), .B(KEYINPUT25), .ZN(new_n747));
  AOI21_X1  g322(.A(new_n747), .B1(G139), .B2(new_n485), .ZN(new_n748));
  AOI22_X1  g323(.A1(new_n462), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n749));
  OR2_X1    g324(.A1(new_n749), .A2(new_n461), .ZN(new_n750));
  AND2_X1   g325(.A1(new_n748), .A2(new_n750), .ZN(new_n751));
  OAI21_X1  g326(.A(new_n745), .B1(new_n751), .B2(new_n727), .ZN(new_n752));
  XOR2_X1   g327(.A(new_n752), .B(G2072), .Z(new_n753));
  INV_X1    g328(.A(G1961), .ZN(new_n754));
  NOR2_X1   g329(.A1(G171), .A2(new_n690), .ZN(new_n755));
  AOI21_X1  g330(.A(new_n755), .B1(G5), .B2(new_n690), .ZN(new_n756));
  OAI21_X1  g331(.A(new_n753), .B1(new_n754), .B2(new_n756), .ZN(new_n757));
  NOR2_X1   g332(.A1(new_n552), .A2(new_n690), .ZN(new_n758));
  AOI21_X1  g333(.A(new_n758), .B1(new_n690), .B2(G19), .ZN(new_n759));
  INV_X1    g334(.A(new_n759), .ZN(new_n760));
  OR2_X1    g335(.A1(new_n760), .A2(G1341), .ZN(new_n761));
  XOR2_X1   g336(.A(KEYINPUT31), .B(G11), .Z(new_n762));
  NOR2_X1   g337(.A1(new_n627), .A2(new_n727), .ZN(new_n763));
  XNOR2_X1  g338(.A(KEYINPUT30), .B(G28), .ZN(new_n764));
  AOI211_X1 g339(.A(new_n762), .B(new_n763), .C1(new_n727), .C2(new_n764), .ZN(new_n765));
  NAND2_X1  g340(.A1(new_n756), .A2(new_n754), .ZN(new_n766));
  NAND2_X1  g341(.A1(new_n760), .A2(G1341), .ZN(new_n767));
  NAND4_X1  g342(.A1(new_n761), .A2(new_n765), .A3(new_n766), .A4(new_n767), .ZN(new_n768));
  NOR3_X1   g343(.A1(new_n744), .A2(new_n757), .A3(new_n768), .ZN(new_n769));
  NAND2_X1  g344(.A1(new_n743), .A2(new_n738), .ZN(new_n770));
  XOR2_X1   g345(.A(new_n770), .B(KEYINPUT95), .Z(new_n771));
  NAND4_X1  g346(.A1(new_n733), .A2(new_n737), .A3(new_n769), .A4(new_n771), .ZN(new_n772));
  NAND2_X1  g347(.A1(new_n727), .A2(G35), .ZN(new_n773));
  OAI21_X1  g348(.A(new_n773), .B1(G162), .B2(new_n727), .ZN(new_n774));
  XNOR2_X1  g349(.A(new_n774), .B(KEYINPUT29), .ZN(new_n775));
  OR2_X1    g350(.A1(new_n775), .A2(G2090), .ZN(new_n776));
  NOR2_X1   g351(.A1(new_n602), .A2(new_n690), .ZN(new_n777));
  AOI21_X1  g352(.A(new_n777), .B1(G4), .B2(new_n690), .ZN(new_n778));
  XNOR2_X1  g353(.A(KEYINPUT89), .B(G1348), .ZN(new_n779));
  AND2_X1   g354(.A1(new_n778), .A2(new_n779), .ZN(new_n780));
  NOR2_X1   g355(.A1(new_n778), .A2(new_n779), .ZN(new_n781));
  XNOR2_X1  g356(.A(KEYINPUT90), .B(KEYINPUT28), .ZN(new_n782));
  XNOR2_X1  g357(.A(new_n782), .B(KEYINPUT91), .ZN(new_n783));
  NAND2_X1  g358(.A1(new_n727), .A2(G26), .ZN(new_n784));
  XOR2_X1   g359(.A(new_n783), .B(new_n784), .Z(new_n785));
  NAND2_X1  g360(.A1(new_n485), .A2(G140), .ZN(new_n786));
  NAND2_X1  g361(.A1(new_n482), .A2(G128), .ZN(new_n787));
  OR2_X1    g362(.A1(G104), .A2(G2105), .ZN(new_n788));
  OAI211_X1 g363(.A(new_n788), .B(G2104), .C1(G116), .C2(new_n461), .ZN(new_n789));
  NAND3_X1  g364(.A1(new_n786), .A2(new_n787), .A3(new_n789), .ZN(new_n790));
  AOI21_X1  g365(.A(new_n785), .B1(G29), .B2(new_n790), .ZN(new_n791));
  INV_X1    g366(.A(G2067), .ZN(new_n792));
  XNOR2_X1  g367(.A(new_n791), .B(new_n792), .ZN(new_n793));
  NAND2_X1  g368(.A1(new_n690), .A2(G21), .ZN(new_n794));
  OAI21_X1  g369(.A(new_n794), .B1(G168), .B2(new_n690), .ZN(new_n795));
  XNOR2_X1  g370(.A(new_n795), .B(G1966), .ZN(new_n796));
  NOR4_X1   g371(.A1(new_n780), .A2(new_n781), .A3(new_n793), .A4(new_n796), .ZN(new_n797));
  NAND2_X1  g372(.A1(new_n775), .A2(G2090), .ZN(new_n798));
  NAND2_X1  g373(.A1(new_n690), .A2(G20), .ZN(new_n799));
  XOR2_X1   g374(.A(new_n799), .B(KEYINPUT96), .Z(new_n800));
  XNOR2_X1  g375(.A(new_n800), .B(KEYINPUT23), .ZN(new_n801));
  AOI21_X1  g376(.A(new_n801), .B1(G299), .B2(G16), .ZN(new_n802));
  XNOR2_X1  g377(.A(new_n802), .B(G1956), .ZN(new_n803));
  NAND4_X1  g378(.A1(new_n776), .A2(new_n797), .A3(new_n798), .A4(new_n803), .ZN(new_n804));
  OR2_X1    g379(.A1(new_n772), .A2(new_n804), .ZN(new_n805));
  NOR2_X1   g380(.A1(new_n717), .A2(new_n805), .ZN(G311));
  INV_X1    g381(.A(G311), .ZN(G150));
  AOI22_X1  g382(.A1(new_n527), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n808));
  NOR2_X1   g383(.A1(new_n808), .A2(new_n540), .ZN(new_n809));
  INV_X1    g384(.A(G93), .ZN(new_n810));
  INV_X1    g385(.A(G55), .ZN(new_n811));
  OAI22_X1  g386(.A1(new_n542), .A2(new_n810), .B1(new_n535), .B2(new_n811), .ZN(new_n812));
  OR2_X1    g387(.A1(new_n809), .A2(new_n812), .ZN(new_n813));
  NAND2_X1  g388(.A1(new_n813), .A2(G860), .ZN(new_n814));
  XNOR2_X1  g389(.A(new_n814), .B(KEYINPUT98), .ZN(new_n815));
  XNOR2_X1  g390(.A(new_n815), .B(KEYINPUT37), .ZN(new_n816));
  NAND2_X1  g391(.A1(new_n602), .A2(G559), .ZN(new_n817));
  XNOR2_X1  g392(.A(new_n817), .B(KEYINPUT38), .ZN(new_n818));
  OR2_X1    g393(.A1(new_n548), .A2(new_n551), .ZN(new_n819));
  NAND2_X1  g394(.A1(new_n819), .A2(new_n813), .ZN(new_n820));
  NOR2_X1   g395(.A1(new_n809), .A2(new_n812), .ZN(new_n821));
  NAND2_X1  g396(.A1(new_n552), .A2(new_n821), .ZN(new_n822));
  NAND2_X1  g397(.A1(new_n820), .A2(new_n822), .ZN(new_n823));
  XNOR2_X1  g398(.A(new_n818), .B(new_n823), .ZN(new_n824));
  INV_X1    g399(.A(KEYINPUT39), .ZN(new_n825));
  NAND2_X1  g400(.A1(new_n824), .A2(new_n825), .ZN(new_n826));
  XOR2_X1   g401(.A(new_n826), .B(KEYINPUT97), .Z(new_n827));
  INV_X1    g402(.A(G860), .ZN(new_n828));
  OAI21_X1  g403(.A(new_n828), .B1(new_n824), .B2(new_n825), .ZN(new_n829));
  OAI21_X1  g404(.A(new_n816), .B1(new_n827), .B2(new_n829), .ZN(G145));
  XOR2_X1   g405(.A(G162), .B(new_n627), .Z(new_n831));
  XNOR2_X1  g406(.A(G160), .B(KEYINPUT99), .ZN(new_n832));
  XOR2_X1   g407(.A(new_n831), .B(new_n832), .Z(new_n833));
  INV_X1    g408(.A(new_n790), .ZN(new_n834));
  NAND3_X1  g409(.A1(new_n723), .A2(new_n834), .A3(new_n724), .ZN(new_n835));
  INV_X1    g410(.A(new_n835), .ZN(new_n836));
  AOI21_X1  g411(.A(new_n834), .B1(new_n723), .B2(new_n724), .ZN(new_n837));
  OAI211_X1 g412(.A(new_n500), .B(new_n495), .C1(new_n836), .C2(new_n837), .ZN(new_n838));
  INV_X1    g413(.A(new_n837), .ZN(new_n839));
  NAND2_X1  g414(.A1(new_n495), .A2(new_n500), .ZN(new_n840));
  NAND3_X1  g415(.A1(new_n839), .A2(new_n840), .A3(new_n835), .ZN(new_n841));
  NAND2_X1  g416(.A1(new_n838), .A2(new_n841), .ZN(new_n842));
  INV_X1    g417(.A(new_n751), .ZN(new_n843));
  NAND2_X1  g418(.A1(new_n842), .A2(new_n843), .ZN(new_n844));
  NAND3_X1  g419(.A1(new_n838), .A2(new_n751), .A3(new_n841), .ZN(new_n845));
  NAND2_X1  g420(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  XOR2_X1   g421(.A(new_n710), .B(new_n618), .Z(new_n847));
  NAND2_X1  g422(.A1(new_n482), .A2(G130), .ZN(new_n848));
  OR2_X1    g423(.A1(G106), .A2(G2105), .ZN(new_n849));
  OAI211_X1 g424(.A(new_n849), .B(G2104), .C1(G118), .C2(new_n461), .ZN(new_n850));
  NAND2_X1  g425(.A1(new_n848), .A2(new_n850), .ZN(new_n851));
  AOI21_X1  g426(.A(new_n851), .B1(G142), .B2(new_n485), .ZN(new_n852));
  XNOR2_X1  g427(.A(new_n847), .B(new_n852), .ZN(new_n853));
  INV_X1    g428(.A(new_n853), .ZN(new_n854));
  NAND2_X1  g429(.A1(new_n846), .A2(new_n854), .ZN(new_n855));
  NAND3_X1  g430(.A1(new_n844), .A2(new_n853), .A3(new_n845), .ZN(new_n856));
  NAND3_X1  g431(.A1(new_n833), .A2(new_n855), .A3(new_n856), .ZN(new_n857));
  INV_X1    g432(.A(G37), .ZN(new_n858));
  AND2_X1   g433(.A1(new_n857), .A2(new_n858), .ZN(new_n859));
  INV_X1    g434(.A(KEYINPUT100), .ZN(new_n860));
  NAND2_X1  g435(.A1(new_n856), .A2(new_n860), .ZN(new_n861));
  NAND2_X1  g436(.A1(new_n861), .A2(new_n855), .ZN(new_n862));
  NAND3_X1  g437(.A1(new_n846), .A2(new_n860), .A3(new_n854), .ZN(new_n863));
  AOI21_X1  g438(.A(new_n833), .B1(new_n862), .B2(new_n863), .ZN(new_n864));
  NOR2_X1   g439(.A1(new_n864), .A2(KEYINPUT101), .ZN(new_n865));
  INV_X1    g440(.A(KEYINPUT101), .ZN(new_n866));
  AOI211_X1 g441(.A(new_n866), .B(new_n833), .C1(new_n862), .C2(new_n863), .ZN(new_n867));
  OAI21_X1  g442(.A(new_n859), .B1(new_n865), .B2(new_n867), .ZN(new_n868));
  XNOR2_X1  g443(.A(new_n868), .B(KEYINPUT40), .ZN(G395));
  XOR2_X1   g444(.A(new_n612), .B(new_n823), .Z(new_n870));
  NAND2_X1  g445(.A1(new_n602), .A2(new_n607), .ZN(new_n871));
  NAND2_X1  g446(.A1(new_n601), .A2(G299), .ZN(new_n872));
  NAND2_X1  g447(.A1(new_n871), .A2(new_n872), .ZN(new_n873));
  INV_X1    g448(.A(KEYINPUT41), .ZN(new_n874));
  NAND2_X1  g449(.A1(new_n873), .A2(new_n874), .ZN(new_n875));
  AND2_X1   g450(.A1(new_n871), .A2(new_n872), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n876), .A2(KEYINPUT41), .ZN(new_n877));
  NAND3_X1  g452(.A1(new_n870), .A2(new_n875), .A3(new_n877), .ZN(new_n878));
  OAI21_X1  g453(.A(new_n878), .B1(new_n870), .B2(new_n873), .ZN(new_n879));
  INV_X1    g454(.A(KEYINPUT102), .ZN(new_n880));
  NOR2_X1   g455(.A1(new_n879), .A2(new_n880), .ZN(new_n881));
  XNOR2_X1  g456(.A(G166), .B(G288), .ZN(new_n882));
  XNOR2_X1  g457(.A(G290), .B(G305), .ZN(new_n883));
  OR2_X1    g458(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  NAND2_X1  g459(.A1(new_n882), .A2(new_n883), .ZN(new_n885));
  NAND2_X1  g460(.A1(new_n884), .A2(new_n885), .ZN(new_n886));
  INV_X1    g461(.A(KEYINPUT42), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n886), .A2(new_n887), .ZN(new_n888));
  NAND3_X1  g463(.A1(new_n884), .A2(KEYINPUT42), .A3(new_n885), .ZN(new_n889));
  NAND2_X1  g464(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n879), .A2(new_n880), .ZN(new_n891));
  AOI21_X1  g466(.A(new_n881), .B1(new_n890), .B2(new_n891), .ZN(new_n892));
  AOI211_X1 g467(.A(new_n880), .B(new_n879), .C1(new_n888), .C2(new_n889), .ZN(new_n893));
  OAI21_X1  g468(.A(G868), .B1(new_n892), .B2(new_n893), .ZN(new_n894));
  NOR2_X1   g469(.A1(new_n821), .A2(G868), .ZN(new_n895));
  INV_X1    g470(.A(new_n895), .ZN(new_n896));
  NAND2_X1  g471(.A1(new_n894), .A2(new_n896), .ZN(G331));
  NOR2_X1   g472(.A1(G331), .A2(KEYINPUT103), .ZN(new_n898));
  INV_X1    g473(.A(KEYINPUT103), .ZN(new_n899));
  AOI21_X1  g474(.A(new_n899), .B1(new_n894), .B2(new_n896), .ZN(new_n900));
  NOR2_X1   g475(.A1(new_n898), .A2(new_n900), .ZN(G295));
  INV_X1    g476(.A(KEYINPUT104), .ZN(new_n902));
  NAND3_X1  g477(.A1(new_n820), .A2(G301), .A3(new_n822), .ZN(new_n903));
  INV_X1    g478(.A(new_n903), .ZN(new_n904));
  AOI21_X1  g479(.A(G301), .B1(new_n820), .B2(new_n822), .ZN(new_n905));
  OAI21_X1  g480(.A(G286), .B1(new_n904), .B2(new_n905), .ZN(new_n906));
  INV_X1    g481(.A(new_n905), .ZN(new_n907));
  NAND3_X1  g482(.A1(new_n907), .A2(G168), .A3(new_n903), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n906), .A2(new_n908), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n909), .A2(new_n876), .ZN(new_n910));
  NAND4_X1  g485(.A1(new_n877), .A2(new_n906), .A3(new_n875), .A4(new_n908), .ZN(new_n911));
  AOI21_X1  g486(.A(new_n902), .B1(new_n910), .B2(new_n911), .ZN(new_n912));
  AND2_X1   g487(.A1(new_n911), .A2(new_n902), .ZN(new_n913));
  OAI21_X1  g488(.A(new_n886), .B1(new_n912), .B2(new_n913), .ZN(new_n914));
  INV_X1    g489(.A(KEYINPUT105), .ZN(new_n915));
  NAND3_X1  g490(.A1(new_n914), .A2(new_n915), .A3(new_n858), .ZN(new_n916));
  OR3_X1    g491(.A1(new_n886), .A2(new_n912), .A3(new_n913), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n916), .A2(new_n917), .ZN(new_n918));
  AOI21_X1  g493(.A(new_n915), .B1(new_n914), .B2(new_n858), .ZN(new_n919));
  OAI21_X1  g494(.A(KEYINPUT43), .B1(new_n918), .B2(new_n919), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n910), .A2(new_n911), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n886), .A2(new_n921), .ZN(new_n922));
  XNOR2_X1  g497(.A(new_n922), .B(KEYINPUT106), .ZN(new_n923));
  INV_X1    g498(.A(KEYINPUT43), .ZN(new_n924));
  NAND4_X1  g499(.A1(new_n923), .A2(new_n924), .A3(new_n858), .A4(new_n917), .ZN(new_n925));
  NAND2_X1  g500(.A1(new_n920), .A2(new_n925), .ZN(new_n926));
  INV_X1    g501(.A(KEYINPUT44), .ZN(new_n927));
  NAND2_X1  g502(.A1(new_n926), .A2(new_n927), .ZN(new_n928));
  OAI21_X1  g503(.A(new_n924), .B1(new_n918), .B2(new_n919), .ZN(new_n929));
  NAND4_X1  g504(.A1(new_n923), .A2(KEYINPUT43), .A3(new_n858), .A4(new_n917), .ZN(new_n930));
  AND2_X1   g505(.A1(new_n929), .A2(new_n930), .ZN(new_n931));
  OAI21_X1  g506(.A(new_n928), .B1(new_n927), .B2(new_n931), .ZN(G397));
  INV_X1    g507(.A(KEYINPUT117), .ZN(new_n933));
  AOI21_X1  g508(.A(G1384), .B1(new_n495), .B2(new_n500), .ZN(new_n934));
  INV_X1    g509(.A(KEYINPUT50), .ZN(new_n935));
  NAND2_X1  g510(.A1(new_n934), .A2(new_n935), .ZN(new_n936));
  INV_X1    g511(.A(G125), .ZN(new_n937));
  NOR2_X1   g512(.A1(new_n481), .A2(new_n937), .ZN(new_n938));
  XNOR2_X1  g513(.A(new_n464), .B(KEYINPUT67), .ZN(new_n939));
  OAI21_X1  g514(.A(G2105), .B1(new_n938), .B2(new_n939), .ZN(new_n940));
  AND3_X1   g515(.A1(new_n470), .A2(new_n472), .A3(new_n473), .ZN(new_n941));
  AOI21_X1  g516(.A(new_n473), .B1(new_n470), .B2(new_n472), .ZN(new_n942));
  OAI211_X1 g517(.A(new_n940), .B(G40), .C1(new_n941), .C2(new_n942), .ZN(new_n943));
  NOR2_X1   g518(.A1(new_n943), .A2(G2090), .ZN(new_n944));
  INV_X1    g519(.A(G1384), .ZN(new_n945));
  OAI21_X1  g520(.A(new_n945), .B1(new_n501), .B2(new_n502), .ZN(new_n946));
  AND3_X1   g521(.A1(new_n946), .A2(KEYINPUT107), .A3(KEYINPUT50), .ZN(new_n947));
  AOI21_X1  g522(.A(KEYINPUT107), .B1(new_n946), .B2(KEYINPUT50), .ZN(new_n948));
  OAI211_X1 g523(.A(new_n936), .B(new_n944), .C1(new_n947), .C2(new_n948), .ZN(new_n949));
  NAND2_X1  g524(.A1(new_n949), .A2(KEYINPUT108), .ZN(new_n950));
  INV_X1    g525(.A(KEYINPUT107), .ZN(new_n951));
  INV_X1    g526(.A(KEYINPUT71), .ZN(new_n952));
  NAND2_X1  g527(.A1(new_n840), .A2(new_n952), .ZN(new_n953));
  NAND3_X1  g528(.A1(new_n495), .A2(KEYINPUT71), .A3(new_n500), .ZN(new_n954));
  AOI21_X1  g529(.A(G1384), .B1(new_n953), .B2(new_n954), .ZN(new_n955));
  OAI21_X1  g530(.A(new_n951), .B1(new_n955), .B2(new_n935), .ZN(new_n956));
  NAND3_X1  g531(.A1(new_n946), .A2(KEYINPUT107), .A3(KEYINPUT50), .ZN(new_n957));
  NAND2_X1  g532(.A1(new_n956), .A2(new_n957), .ZN(new_n958));
  INV_X1    g533(.A(KEYINPUT108), .ZN(new_n959));
  NAND4_X1  g534(.A1(new_n958), .A2(new_n959), .A3(new_n936), .A4(new_n944), .ZN(new_n960));
  NAND2_X1  g535(.A1(new_n934), .A2(KEYINPUT45), .ZN(new_n961));
  INV_X1    g536(.A(new_n943), .ZN(new_n962));
  NAND2_X1  g537(.A1(new_n961), .A2(new_n962), .ZN(new_n963));
  INV_X1    g538(.A(KEYINPUT45), .ZN(new_n964));
  AOI21_X1  g539(.A(new_n963), .B1(new_n964), .B2(new_n946), .ZN(new_n965));
  NOR2_X1   g540(.A1(new_n965), .A2(G1971), .ZN(new_n966));
  INV_X1    g541(.A(new_n966), .ZN(new_n967));
  NAND3_X1  g542(.A1(new_n950), .A2(new_n960), .A3(new_n967), .ZN(new_n968));
  NAND2_X1  g543(.A1(new_n968), .A2(G8), .ZN(new_n969));
  NAND3_X1  g544(.A1(new_n523), .A2(G8), .A3(new_n525), .ZN(new_n970));
  XNOR2_X1  g545(.A(new_n970), .B(KEYINPUT55), .ZN(new_n971));
  NAND2_X1  g546(.A1(new_n969), .A2(new_n971), .ZN(new_n972));
  INV_X1    g547(.A(G8), .ZN(new_n973));
  AOI21_X1  g548(.A(new_n966), .B1(new_n949), .B2(KEYINPUT108), .ZN(new_n974));
  AOI211_X1 g549(.A(new_n973), .B(new_n971), .C1(new_n974), .C2(new_n960), .ZN(new_n975));
  OAI211_X1 g550(.A(G40), .B(G160), .C1(new_n934), .C2(KEYINPUT45), .ZN(new_n976));
  AOI21_X1  g551(.A(new_n976), .B1(new_n955), .B2(KEYINPUT45), .ZN(new_n977));
  OAI21_X1  g552(.A(KEYINPUT116), .B1(new_n977), .B2(G1966), .ZN(new_n978));
  NAND2_X1  g553(.A1(new_n840), .A2(new_n945), .ZN(new_n979));
  AOI21_X1  g554(.A(new_n943), .B1(new_n979), .B2(new_n964), .ZN(new_n980));
  OAI21_X1  g555(.A(new_n980), .B1(new_n946), .B2(new_n964), .ZN(new_n981));
  INV_X1    g556(.A(KEYINPUT116), .ZN(new_n982));
  INV_X1    g557(.A(G1966), .ZN(new_n983));
  NAND3_X1  g558(.A1(new_n981), .A2(new_n982), .A3(new_n983), .ZN(new_n984));
  NAND2_X1  g559(.A1(new_n978), .A2(new_n984), .ZN(new_n985));
  NAND4_X1  g560(.A1(new_n958), .A2(new_n738), .A3(new_n962), .A4(new_n936), .ZN(new_n986));
  AOI21_X1  g561(.A(new_n973), .B1(new_n985), .B2(new_n986), .ZN(new_n987));
  OAI21_X1  g562(.A(G8), .B1(new_n979), .B2(new_n943), .ZN(new_n988));
  NAND3_X1  g563(.A1(new_n527), .A2(new_n529), .A3(G86), .ZN(new_n989));
  NAND2_X1  g564(.A1(new_n517), .A2(G48), .ZN(new_n990));
  NAND4_X1  g565(.A1(new_n584), .A2(new_n688), .A3(new_n989), .A4(new_n990), .ZN(new_n991));
  NAND2_X1  g566(.A1(new_n991), .A2(KEYINPUT111), .ZN(new_n992));
  INV_X1    g567(.A(KEYINPUT111), .ZN(new_n993));
  NAND4_X1  g568(.A1(new_n576), .A2(new_n993), .A3(new_n688), .A4(new_n584), .ZN(new_n994));
  NAND2_X1  g569(.A1(new_n992), .A2(new_n994), .ZN(new_n995));
  NAND2_X1  g570(.A1(G305), .A2(G1981), .ZN(new_n996));
  NAND3_X1  g571(.A1(new_n995), .A2(KEYINPUT49), .A3(new_n996), .ZN(new_n997));
  INV_X1    g572(.A(KEYINPUT113), .ZN(new_n998));
  AOI21_X1  g573(.A(new_n988), .B1(new_n997), .B2(new_n998), .ZN(new_n999));
  AOI22_X1  g574(.A1(new_n992), .A2(new_n994), .B1(G305), .B2(G1981), .ZN(new_n1000));
  NAND3_X1  g575(.A1(new_n1000), .A2(KEYINPUT113), .A3(KEYINPUT49), .ZN(new_n1001));
  INV_X1    g576(.A(KEYINPUT112), .ZN(new_n1002));
  AND2_X1   g577(.A1(new_n1000), .A2(new_n1002), .ZN(new_n1003));
  INV_X1    g578(.A(KEYINPUT49), .ZN(new_n1004));
  OAI21_X1  g579(.A(new_n1004), .B1(new_n1000), .B2(new_n1002), .ZN(new_n1005));
  OAI211_X1 g580(.A(new_n999), .B(new_n1001), .C1(new_n1003), .C2(new_n1005), .ZN(new_n1006));
  AND3_X1   g581(.A1(new_n572), .A2(new_n573), .A3(new_n574), .ZN(new_n1007));
  NAND2_X1  g582(.A1(new_n1007), .A2(G1976), .ZN(new_n1008));
  OAI211_X1 g583(.A(new_n1008), .B(G8), .C1(new_n979), .C2(new_n943), .ZN(new_n1009));
  INV_X1    g584(.A(KEYINPUT110), .ZN(new_n1010));
  INV_X1    g585(.A(KEYINPUT52), .ZN(new_n1011));
  OAI21_X1  g586(.A(new_n1011), .B1(new_n1007), .B2(G1976), .ZN(new_n1012));
  OR3_X1    g587(.A1(new_n1009), .A2(new_n1010), .A3(new_n1012), .ZN(new_n1013));
  OAI21_X1  g588(.A(new_n1010), .B1(new_n1009), .B2(new_n1012), .ZN(new_n1014));
  NAND2_X1  g589(.A1(new_n1013), .A2(new_n1014), .ZN(new_n1015));
  NAND2_X1  g590(.A1(new_n1009), .A2(KEYINPUT52), .ZN(new_n1016));
  INV_X1    g591(.A(KEYINPUT109), .ZN(new_n1017));
  NAND2_X1  g592(.A1(new_n1016), .A2(new_n1017), .ZN(new_n1018));
  NAND3_X1  g593(.A1(new_n1009), .A2(KEYINPUT109), .A3(KEYINPUT52), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n1018), .A2(new_n1019), .ZN(new_n1020));
  AND3_X1   g595(.A1(new_n1006), .A2(new_n1015), .A3(new_n1020), .ZN(new_n1021));
  NAND4_X1  g596(.A1(new_n987), .A2(new_n1021), .A3(KEYINPUT63), .A4(G168), .ZN(new_n1022));
  NOR2_X1   g597(.A1(new_n975), .A2(new_n1022), .ZN(new_n1023));
  INV_X1    g598(.A(new_n971), .ZN(new_n1024));
  NAND3_X1  g599(.A1(new_n968), .A2(G8), .A3(new_n1024), .ZN(new_n1025));
  NOR2_X1   g600(.A1(KEYINPUT50), .A2(G1384), .ZN(new_n1026));
  OAI21_X1  g601(.A(new_n1026), .B1(new_n501), .B2(new_n502), .ZN(new_n1027));
  INV_X1    g602(.A(KEYINPUT114), .ZN(new_n1028));
  NAND2_X1  g603(.A1(new_n1027), .A2(new_n1028), .ZN(new_n1029));
  OAI211_X1 g604(.A(KEYINPUT114), .B(new_n1026), .C1(new_n501), .C2(new_n502), .ZN(new_n1030));
  OAI211_X1 g605(.A(G40), .B(G160), .C1(new_n934), .C2(new_n935), .ZN(new_n1031));
  INV_X1    g606(.A(new_n1031), .ZN(new_n1032));
  NAND3_X1  g607(.A1(new_n1029), .A2(new_n1030), .A3(new_n1032), .ZN(new_n1033));
  AOI21_X1  g608(.A(G2090), .B1(new_n1033), .B2(KEYINPUT115), .ZN(new_n1034));
  AOI21_X1  g609(.A(new_n1031), .B1(new_n1028), .B2(new_n1027), .ZN(new_n1035));
  INV_X1    g610(.A(KEYINPUT115), .ZN(new_n1036));
  NAND3_X1  g611(.A1(new_n1035), .A2(new_n1036), .A3(new_n1030), .ZN(new_n1037));
  AOI21_X1  g612(.A(new_n966), .B1(new_n1034), .B2(new_n1037), .ZN(new_n1038));
  OAI21_X1  g613(.A(new_n971), .B1(new_n1038), .B2(new_n973), .ZN(new_n1039));
  AOI211_X1 g614(.A(new_n973), .B(G286), .C1(new_n985), .C2(new_n986), .ZN(new_n1040));
  NAND4_X1  g615(.A1(new_n1025), .A2(new_n1039), .A3(new_n1040), .A4(new_n1021), .ZN(new_n1041));
  INV_X1    g616(.A(KEYINPUT63), .ZN(new_n1042));
  AOI22_X1  g617(.A1(new_n972), .A2(new_n1023), .B1(new_n1041), .B2(new_n1042), .ZN(new_n1043));
  NAND2_X1  g618(.A1(new_n975), .A2(new_n1021), .ZN(new_n1044));
  NOR2_X1   g619(.A1(G288), .A2(G1976), .ZN(new_n1045));
  AND2_X1   g620(.A1(new_n1006), .A2(new_n1045), .ZN(new_n1046));
  INV_X1    g621(.A(new_n995), .ZN(new_n1047));
  OAI221_X1 g622(.A(G8), .B1(new_n943), .B2(new_n979), .C1(new_n1046), .C2(new_n1047), .ZN(new_n1048));
  NAND2_X1  g623(.A1(new_n1044), .A2(new_n1048), .ZN(new_n1049));
  OAI21_X1  g624(.A(new_n933), .B1(new_n1043), .B2(new_n1049), .ZN(new_n1050));
  NAND2_X1  g625(.A1(new_n1041), .A2(new_n1042), .ZN(new_n1051));
  AND2_X1   g626(.A1(new_n1021), .A2(KEYINPUT63), .ZN(new_n1052));
  NAND4_X1  g627(.A1(new_n972), .A2(new_n1025), .A3(new_n1040), .A4(new_n1052), .ZN(new_n1053));
  NAND2_X1  g628(.A1(new_n1051), .A2(new_n1053), .ZN(new_n1054));
  INV_X1    g629(.A(new_n1049), .ZN(new_n1055));
  NAND3_X1  g630(.A1(new_n1054), .A2(KEYINPUT117), .A3(new_n1055), .ZN(new_n1056));
  XOR2_X1   g631(.A(G299), .B(KEYINPUT57), .Z(new_n1057));
  INV_X1    g632(.A(new_n1057), .ZN(new_n1058));
  AOI21_X1  g633(.A(G1956), .B1(new_n1035), .B2(new_n1030), .ZN(new_n1059));
  AOI21_X1  g634(.A(new_n943), .B1(KEYINPUT45), .B2(new_n934), .ZN(new_n1060));
  XNOR2_X1  g635(.A(KEYINPUT56), .B(G2072), .ZN(new_n1061));
  OAI211_X1 g636(.A(new_n1060), .B(new_n1061), .C1(new_n955), .C2(KEYINPUT45), .ZN(new_n1062));
  INV_X1    g637(.A(new_n1062), .ZN(new_n1063));
  OAI21_X1  g638(.A(new_n1058), .B1(new_n1059), .B2(new_n1063), .ZN(new_n1064));
  INV_X1    g639(.A(G1956), .ZN(new_n1065));
  NAND2_X1  g640(.A1(new_n1033), .A2(new_n1065), .ZN(new_n1066));
  NAND3_X1  g641(.A1(new_n1066), .A2(new_n1057), .A3(new_n1062), .ZN(new_n1067));
  AND3_X1   g642(.A1(new_n1064), .A2(new_n1067), .A3(KEYINPUT61), .ZN(new_n1068));
  AOI21_X1  g643(.A(KEYINPUT61), .B1(new_n1064), .B2(new_n1067), .ZN(new_n1069));
  NOR2_X1   g644(.A1(new_n1068), .A2(new_n1069), .ZN(new_n1070));
  INV_X1    g645(.A(KEYINPUT60), .ZN(new_n1071));
  AOI22_X1  g646(.A1(new_n956), .A2(new_n957), .B1(new_n935), .B2(new_n934), .ZN(new_n1072));
  AOI21_X1  g647(.A(G1348), .B1(new_n1072), .B2(new_n962), .ZN(new_n1073));
  INV_X1    g648(.A(KEYINPUT118), .ZN(new_n1074));
  NAND3_X1  g649(.A1(new_n962), .A2(new_n1074), .A3(new_n934), .ZN(new_n1075));
  OAI21_X1  g650(.A(KEYINPUT118), .B1(new_n979), .B2(new_n943), .ZN(new_n1076));
  AOI21_X1  g651(.A(G2067), .B1(new_n1075), .B2(new_n1076), .ZN(new_n1077));
  INV_X1    g652(.A(KEYINPUT119), .ZN(new_n1078));
  XNOR2_X1  g653(.A(new_n1077), .B(new_n1078), .ZN(new_n1079));
  OAI21_X1  g654(.A(new_n1071), .B1(new_n1073), .B2(new_n1079), .ZN(new_n1080));
  OAI211_X1 g655(.A(new_n962), .B(new_n936), .C1(new_n947), .C2(new_n948), .ZN(new_n1081));
  INV_X1    g656(.A(G1348), .ZN(new_n1082));
  NAND2_X1  g657(.A1(new_n1081), .A2(new_n1082), .ZN(new_n1083));
  XNOR2_X1  g658(.A(new_n1077), .B(KEYINPUT119), .ZN(new_n1084));
  INV_X1    g659(.A(KEYINPUT123), .ZN(new_n1085));
  AOI21_X1  g660(.A(new_n1071), .B1(new_n602), .B2(new_n1085), .ZN(new_n1086));
  NAND3_X1  g661(.A1(new_n1083), .A2(new_n1084), .A3(new_n1086), .ZN(new_n1087));
  NOR2_X1   g662(.A1(new_n602), .A2(new_n1085), .ZN(new_n1088));
  INV_X1    g663(.A(new_n1088), .ZN(new_n1089));
  NAND3_X1  g664(.A1(new_n1080), .A2(new_n1087), .A3(new_n1089), .ZN(new_n1090));
  NAND4_X1  g665(.A1(new_n1083), .A2(new_n1084), .A3(new_n1086), .A4(new_n1088), .ZN(new_n1091));
  INV_X1    g666(.A(G1996), .ZN(new_n1092));
  OAI211_X1 g667(.A(new_n1092), .B(new_n1060), .C1(new_n955), .C2(KEYINPUT45), .ZN(new_n1093));
  XOR2_X1   g668(.A(KEYINPUT58), .B(G1341), .Z(new_n1094));
  NAND3_X1  g669(.A1(new_n1075), .A2(new_n1076), .A3(new_n1094), .ZN(new_n1095));
  AOI21_X1  g670(.A(new_n819), .B1(new_n1093), .B2(new_n1095), .ZN(new_n1096));
  AND4_X1   g671(.A1(KEYINPUT121), .A2(new_n1096), .A3(KEYINPUT122), .A4(KEYINPUT59), .ZN(new_n1097));
  NOR2_X1   g672(.A1(new_n1096), .A2(KEYINPUT121), .ZN(new_n1098));
  AOI21_X1  g673(.A(KEYINPUT59), .B1(new_n1096), .B2(KEYINPUT122), .ZN(new_n1099));
  NOR3_X1   g674(.A1(new_n1097), .A2(new_n1098), .A3(new_n1099), .ZN(new_n1100));
  NAND4_X1  g675(.A1(new_n1070), .A2(new_n1090), .A3(new_n1091), .A4(new_n1100), .ZN(new_n1101));
  AOI21_X1  g676(.A(new_n601), .B1(new_n1083), .B2(new_n1084), .ZN(new_n1102));
  INV_X1    g677(.A(KEYINPUT120), .ZN(new_n1103));
  OAI21_X1  g678(.A(new_n1064), .B1(new_n1102), .B2(new_n1103), .ZN(new_n1104));
  AOI211_X1 g679(.A(KEYINPUT120), .B(new_n601), .C1(new_n1083), .C2(new_n1084), .ZN(new_n1105));
  OAI21_X1  g680(.A(new_n1067), .B1(new_n1104), .B2(new_n1105), .ZN(new_n1106));
  NAND2_X1  g681(.A1(new_n1101), .A2(new_n1106), .ZN(new_n1107));
  AOI21_X1  g682(.A(KEYINPUT53), .B1(new_n965), .B2(new_n736), .ZN(new_n1108));
  AOI21_X1  g683(.A(new_n1108), .B1(new_n1081), .B2(new_n754), .ZN(new_n1109));
  AND2_X1   g684(.A1(new_n736), .A2(KEYINPUT53), .ZN(new_n1110));
  NAND3_X1  g685(.A1(new_n980), .A2(new_n961), .A3(new_n1110), .ZN(new_n1111));
  NAND3_X1  g686(.A1(new_n1109), .A2(G301), .A3(new_n1111), .ZN(new_n1112));
  OR2_X1    g687(.A1(new_n1112), .A2(KEYINPUT126), .ZN(new_n1113));
  INV_X1    g688(.A(KEYINPUT54), .ZN(new_n1114));
  NAND2_X1  g689(.A1(new_n977), .A2(new_n1110), .ZN(new_n1115));
  AOI21_X1  g690(.A(G301), .B1(new_n1109), .B2(new_n1115), .ZN(new_n1116));
  NAND2_X1  g691(.A1(new_n1112), .A2(KEYINPUT126), .ZN(new_n1117));
  OAI211_X1 g692(.A(new_n1113), .B(new_n1114), .C1(new_n1116), .C2(new_n1117), .ZN(new_n1118));
  AND3_X1   g693(.A1(new_n1109), .A2(G301), .A3(new_n1115), .ZN(new_n1119));
  AOI21_X1  g694(.A(G301), .B1(new_n1109), .B2(new_n1111), .ZN(new_n1120));
  NOR3_X1   g695(.A1(new_n1119), .A2(new_n1120), .A3(new_n1114), .ZN(new_n1121));
  NAND3_X1  g696(.A1(new_n1025), .A2(new_n1039), .A3(new_n1021), .ZN(new_n1122));
  NOR2_X1   g697(.A1(new_n1121), .A2(new_n1122), .ZN(new_n1123));
  NAND2_X1  g698(.A1(G286), .A2(G8), .ZN(new_n1124));
  XOR2_X1   g699(.A(new_n1124), .B(KEYINPUT124), .Z(new_n1125));
  INV_X1    g700(.A(new_n1125), .ZN(new_n1126));
  AND3_X1   g701(.A1(new_n981), .A2(new_n982), .A3(new_n983), .ZN(new_n1127));
  AOI21_X1  g702(.A(new_n982), .B1(new_n981), .B2(new_n983), .ZN(new_n1128));
  OAI22_X1  g703(.A1(new_n1081), .A2(G2084), .B1(new_n1127), .B2(new_n1128), .ZN(new_n1129));
  AOI221_X4 g704(.A(new_n1126), .B1(KEYINPUT125), .B2(KEYINPUT51), .C1(new_n1129), .C2(G8), .ZN(new_n1130));
  OAI21_X1  g705(.A(KEYINPUT51), .B1(new_n987), .B2(KEYINPUT125), .ZN(new_n1131));
  INV_X1    g706(.A(new_n1131), .ZN(new_n1132));
  AOI21_X1  g707(.A(new_n1125), .B1(new_n985), .B2(new_n986), .ZN(new_n1133));
  NAND2_X1  g708(.A1(new_n1129), .A2(G8), .ZN(new_n1134));
  AOI21_X1  g709(.A(new_n1133), .B1(new_n1134), .B2(new_n1125), .ZN(new_n1135));
  AOI21_X1  g710(.A(new_n1130), .B1(new_n1132), .B2(new_n1135), .ZN(new_n1136));
  NAND4_X1  g711(.A1(new_n1107), .A2(new_n1118), .A3(new_n1123), .A4(new_n1136), .ZN(new_n1137));
  INV_X1    g712(.A(KEYINPUT125), .ZN(new_n1138));
  INV_X1    g713(.A(KEYINPUT51), .ZN(new_n1139));
  OAI211_X1 g714(.A(new_n1134), .B(new_n1125), .C1(new_n1138), .C2(new_n1139), .ZN(new_n1140));
  NAND2_X1  g715(.A1(new_n1129), .A2(new_n1126), .ZN(new_n1141));
  OAI21_X1  g716(.A(new_n1141), .B1(new_n987), .B2(new_n1126), .ZN(new_n1142));
  OAI21_X1  g717(.A(new_n1140), .B1(new_n1142), .B2(new_n1131), .ZN(new_n1143));
  INV_X1    g718(.A(KEYINPUT62), .ZN(new_n1144));
  NAND2_X1  g719(.A1(new_n1143), .A2(new_n1144), .ZN(new_n1145));
  INV_X1    g720(.A(new_n1122), .ZN(new_n1146));
  OAI211_X1 g721(.A(new_n1140), .B(KEYINPUT62), .C1(new_n1142), .C2(new_n1131), .ZN(new_n1147));
  NAND4_X1  g722(.A1(new_n1145), .A2(new_n1146), .A3(new_n1116), .A4(new_n1147), .ZN(new_n1148));
  NAND4_X1  g723(.A1(new_n1050), .A2(new_n1056), .A3(new_n1137), .A4(new_n1148), .ZN(new_n1149));
  NOR2_X1   g724(.A1(new_n934), .A2(KEYINPUT45), .ZN(new_n1150));
  NAND2_X1  g725(.A1(new_n1150), .A2(new_n962), .ZN(new_n1151));
  INV_X1    g726(.A(new_n1151), .ZN(new_n1152));
  XNOR2_X1  g727(.A(new_n790), .B(new_n792), .ZN(new_n1153));
  OAI21_X1  g728(.A(new_n1153), .B1(new_n726), .B2(new_n1092), .ZN(new_n1154));
  AOI21_X1  g729(.A(new_n1154), .B1(new_n1092), .B2(new_n726), .ZN(new_n1155));
  XNOR2_X1  g730(.A(new_n710), .B(new_n712), .ZN(new_n1156));
  NAND2_X1  g731(.A1(new_n1155), .A2(new_n1156), .ZN(new_n1157));
  XNOR2_X1  g732(.A(G290), .B(G1986), .ZN(new_n1158));
  OAI21_X1  g733(.A(new_n1152), .B1(new_n1157), .B2(new_n1158), .ZN(new_n1159));
  NAND2_X1  g734(.A1(new_n1149), .A2(new_n1159), .ZN(new_n1160));
  NAND2_X1  g735(.A1(new_n1152), .A2(new_n1092), .ZN(new_n1161));
  XNOR2_X1  g736(.A(new_n1161), .B(KEYINPUT46), .ZN(new_n1162));
  AND2_X1   g737(.A1(new_n726), .A2(new_n1153), .ZN(new_n1163));
  OAI21_X1  g738(.A(new_n1162), .B1(new_n1151), .B2(new_n1163), .ZN(new_n1164));
  XOR2_X1   g739(.A(new_n1164), .B(KEYINPUT127), .Z(new_n1165));
  OR2_X1    g740(.A1(new_n1165), .A2(KEYINPUT47), .ZN(new_n1166));
  NAND2_X1  g741(.A1(new_n1165), .A2(KEYINPUT47), .ZN(new_n1167));
  NOR2_X1   g742(.A1(new_n710), .A2(new_n713), .ZN(new_n1168));
  NAND2_X1  g743(.A1(new_n1155), .A2(new_n1168), .ZN(new_n1169));
  NAND2_X1  g744(.A1(new_n834), .A2(new_n792), .ZN(new_n1170));
  AOI21_X1  g745(.A(new_n1151), .B1(new_n1169), .B2(new_n1170), .ZN(new_n1171));
  NAND2_X1  g746(.A1(new_n1157), .A2(new_n1152), .ZN(new_n1172));
  NOR3_X1   g747(.A1(new_n1151), .A2(G290), .A3(G1986), .ZN(new_n1173));
  XOR2_X1   g748(.A(new_n1173), .B(KEYINPUT48), .Z(new_n1174));
  AOI21_X1  g749(.A(new_n1171), .B1(new_n1172), .B2(new_n1174), .ZN(new_n1175));
  AND3_X1   g750(.A1(new_n1166), .A2(new_n1167), .A3(new_n1175), .ZN(new_n1176));
  NAND2_X1  g751(.A1(new_n1160), .A2(new_n1176), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g752(.A(G319), .ZN(new_n1179));
  OR2_X1    g753(.A1(G227), .A2(new_n1179), .ZN(new_n1180));
  NOR3_X1   g754(.A1(G229), .A2(G401), .A3(new_n1180), .ZN(new_n1181));
  NAND3_X1  g755(.A1(new_n1181), .A2(new_n868), .A3(new_n926), .ZN(G225));
  INV_X1    g756(.A(G225), .ZN(G308));
endmodule


