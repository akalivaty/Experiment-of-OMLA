//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 1 0 1 1 1 0 0 0 0 1 0 1 0 1 0 0 1 0 0 0 0 0 1 1 1 0 1 1 0 0 1 0 0 0 1 0 1 1 0 0 0 1 1 1 0 1 1 0 1 1 0 0 1 1 0 0 1 0 1 0 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:39:01 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n205, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n690, new_n691, new_n692, new_n693, new_n694, new_n695, new_n696,
    new_n697, new_n698, new_n699, new_n700, new_n701, new_n702, new_n703,
    new_n704, new_n705, new_n706, new_n707, new_n708, new_n709, new_n710,
    new_n711, new_n712, new_n713, new_n714, new_n715, new_n716, new_n717,
    new_n718, new_n719, new_n720, new_n721, new_n722, new_n723, new_n724,
    new_n725, new_n726, new_n727, new_n728, new_n729, new_n730, new_n731,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n772, new_n773, new_n774, new_n775,
    new_n776, new_n777, new_n778, new_n779, new_n780, new_n781, new_n782,
    new_n783, new_n784, new_n785, new_n786, new_n787, new_n788, new_n789,
    new_n790, new_n791, new_n792, new_n793, new_n794, new_n795, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1087,
    new_n1088, new_n1089, new_n1090, new_n1091, new_n1092, new_n1093,
    new_n1094, new_n1095, new_n1096, new_n1097, new_n1098, new_n1099,
    new_n1100, new_n1101, new_n1102, new_n1103, new_n1104, new_n1105,
    new_n1106, new_n1107, new_n1108, new_n1109, new_n1110, new_n1111,
    new_n1112, new_n1113, new_n1114, new_n1115, new_n1116, new_n1118,
    new_n1119, new_n1120, new_n1121, new_n1122, new_n1123, new_n1124,
    new_n1125, new_n1126, new_n1127, new_n1128, new_n1129, new_n1130,
    new_n1131, new_n1132, new_n1133, new_n1134, new_n1135, new_n1136,
    new_n1137, new_n1138, new_n1139, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1186, new_n1187, new_n1188, new_n1189, new_n1190, new_n1191,
    new_n1192, new_n1193, new_n1194, new_n1195, new_n1196, new_n1197,
    new_n1198, new_n1199, new_n1200, new_n1201, new_n1202, new_n1203,
    new_n1204, new_n1205, new_n1206, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1251, new_n1252,
    new_n1253, new_n1254, new_n1255, new_n1256, new_n1257, new_n1258,
    new_n1259, new_n1260, new_n1261, new_n1262, new_n1263, new_n1264,
    new_n1265, new_n1266, new_n1267, new_n1268, new_n1269, new_n1270,
    new_n1271, new_n1272, new_n1273, new_n1274, new_n1276, new_n1277,
    new_n1278, new_n1279, new_n1280, new_n1281, new_n1282, new_n1283,
    new_n1284, new_n1285, new_n1286, new_n1287, new_n1288, new_n1289,
    new_n1290, new_n1291, new_n1292, new_n1293, new_n1294, new_n1295,
    new_n1296, new_n1297, new_n1298, new_n1299, new_n1300, new_n1301,
    new_n1303, new_n1304, new_n1305, new_n1306, new_n1307, new_n1308,
    new_n1309, new_n1310, new_n1311, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1346,
    new_n1347, new_n1348, new_n1349, new_n1350, new_n1351, new_n1352,
    new_n1353, new_n1354, new_n1355, new_n1356, new_n1357, new_n1358,
    new_n1359, new_n1360, new_n1361, new_n1362, new_n1363, new_n1364,
    new_n1365, new_n1366, new_n1367, new_n1368, new_n1369, new_n1370,
    new_n1371, new_n1372, new_n1373, new_n1374, new_n1375, new_n1376,
    new_n1377, new_n1378, new_n1379, new_n1380, new_n1381, new_n1382,
    new_n1383, new_n1384, new_n1385, new_n1386, new_n1388, new_n1389,
    new_n1390, new_n1391, new_n1392, new_n1393, new_n1394;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(new_n205));
  XNOR2_X1  g0005(.A(new_n205), .B(KEYINPUT64), .ZN(G355));
  NAND2_X1  g0006(.A1(G1), .A2(G20), .ZN(new_n207));
  NOR2_X1   g0007(.A1(new_n207), .A2(G13), .ZN(new_n208));
  OAI211_X1 g0008(.A(new_n208), .B(G250), .C1(G257), .C2(G264), .ZN(new_n209));
  INV_X1    g0009(.A(KEYINPUT0), .ZN(new_n210));
  INV_X1    g0010(.A(new_n201), .ZN(new_n211));
  NAND2_X1  g0011(.A1(new_n211), .A2(G50), .ZN(new_n212));
  INV_X1    g0012(.A(new_n212), .ZN(new_n213));
  NAND2_X1  g0013(.A1(G1), .A2(G13), .ZN(new_n214));
  INV_X1    g0014(.A(G20), .ZN(new_n215));
  NOR2_X1   g0015(.A1(new_n214), .A2(new_n215), .ZN(new_n216));
  AOI22_X1  g0016(.A1(new_n209), .A2(new_n210), .B1(new_n213), .B2(new_n216), .ZN(new_n217));
  AOI22_X1  g0017(.A1(G87), .A2(G250), .B1(G107), .B2(G264), .ZN(new_n218));
  INV_X1    g0018(.A(G58), .ZN(new_n219));
  INV_X1    g0019(.A(G232), .ZN(new_n220));
  INV_X1    g0020(.A(G97), .ZN(new_n221));
  INV_X1    g0021(.A(G257), .ZN(new_n222));
  OAI221_X1 g0022(.A(new_n218), .B1(new_n219), .B2(new_n220), .C1(new_n221), .C2(new_n222), .ZN(new_n223));
  NAND2_X1  g0023(.A1(new_n223), .A2(KEYINPUT66), .ZN(new_n224));
  XNOR2_X1  g0024(.A(KEYINPUT65), .B(G77), .ZN(new_n225));
  NAND2_X1  g0025(.A1(new_n225), .A2(G244), .ZN(new_n226));
  NAND2_X1  g0026(.A1(G68), .A2(G238), .ZN(new_n227));
  AOI22_X1  g0027(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n228));
  NAND4_X1  g0028(.A1(new_n224), .A2(new_n226), .A3(new_n227), .A4(new_n228), .ZN(new_n229));
  NOR2_X1   g0029(.A1(new_n223), .A2(KEYINPUT66), .ZN(new_n230));
  OAI21_X1  g0030(.A(new_n207), .B1(new_n229), .B2(new_n230), .ZN(new_n231));
  OAI221_X1 g0031(.A(new_n217), .B1(new_n210), .B2(new_n209), .C1(new_n231), .C2(KEYINPUT1), .ZN(new_n232));
  AOI21_X1  g0032(.A(new_n232), .B1(KEYINPUT1), .B2(new_n231), .ZN(G361));
  XNOR2_X1  g0033(.A(G238), .B(G244), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n234), .B(KEYINPUT2), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n235), .B(G226), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n236), .B(new_n220), .ZN(new_n237));
  XOR2_X1   g0037(.A(new_n237), .B(KEYINPUT67), .Z(new_n238));
  XNOR2_X1  g0038(.A(G250), .B(G257), .ZN(new_n239));
  XNOR2_X1  g0039(.A(G264), .B(G270), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n238), .B(new_n241), .ZN(G358));
  XOR2_X1   g0042(.A(G68), .B(G77), .Z(new_n243));
  XNOR2_X1  g0043(.A(G50), .B(G58), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XOR2_X1   g0045(.A(G87), .B(G97), .Z(new_n246));
  XNOR2_X1  g0046(.A(G107), .B(G116), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n246), .B(new_n247), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n245), .B(new_n248), .ZN(G351));
  INV_X1    g0049(.A(KEYINPUT77), .ZN(new_n250));
  INV_X1    g0050(.A(G41), .ZN(new_n251));
  INV_X1    g0051(.A(G45), .ZN(new_n252));
  NAND2_X1  g0052(.A1(new_n251), .A2(new_n252), .ZN(new_n253));
  INV_X1    g0053(.A(new_n253), .ZN(new_n254));
  INV_X1    g0054(.A(G274), .ZN(new_n255));
  OR3_X1    g0055(.A1(new_n254), .A2(G1), .A3(new_n255), .ZN(new_n256));
  OR2_X1    g0056(.A1(KEYINPUT68), .A2(G1), .ZN(new_n257));
  NAND2_X1  g0057(.A1(KEYINPUT68), .A2(G1), .ZN(new_n258));
  NAND3_X1  g0058(.A1(new_n257), .A2(new_n253), .A3(new_n258), .ZN(new_n259));
  AND2_X1   g0059(.A1(G1), .A2(G13), .ZN(new_n260));
  NAND2_X1  g0060(.A1(G33), .A2(G41), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n260), .A2(new_n261), .ZN(new_n262));
  NAND2_X1  g0062(.A1(new_n259), .A2(new_n262), .ZN(new_n263));
  INV_X1    g0063(.A(G238), .ZN(new_n264));
  OAI21_X1  g0064(.A(new_n256), .B1(new_n263), .B2(new_n264), .ZN(new_n265));
  INV_X1    g0065(.A(new_n265), .ZN(new_n266));
  INV_X1    g0066(.A(KEYINPUT3), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n267), .A2(G33), .ZN(new_n268));
  INV_X1    g0068(.A(G33), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n269), .A2(KEYINPUT3), .ZN(new_n270));
  INV_X1    g0070(.A(G1698), .ZN(new_n271));
  NAND4_X1  g0071(.A1(new_n268), .A2(new_n270), .A3(G226), .A4(new_n271), .ZN(new_n272));
  INV_X1    g0072(.A(KEYINPUT73), .ZN(new_n273));
  NAND2_X1  g0073(.A1(new_n272), .A2(new_n273), .ZN(new_n274));
  XNOR2_X1  g0074(.A(KEYINPUT3), .B(G33), .ZN(new_n275));
  NAND4_X1  g0075(.A1(new_n275), .A2(KEYINPUT73), .A3(G226), .A4(new_n271), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n274), .A2(new_n276), .ZN(new_n277));
  NAND4_X1  g0077(.A1(new_n268), .A2(new_n270), .A3(G232), .A4(G1698), .ZN(new_n278));
  NAND2_X1  g0078(.A1(G33), .A2(G97), .ZN(new_n279));
  NAND2_X1  g0079(.A1(new_n278), .A2(new_n279), .ZN(new_n280));
  INV_X1    g0080(.A(new_n280), .ZN(new_n281));
  NAND2_X1  g0081(.A1(new_n277), .A2(new_n281), .ZN(new_n282));
  INV_X1    g0082(.A(new_n262), .ZN(new_n283));
  AOI21_X1  g0083(.A(KEYINPUT74), .B1(new_n282), .B2(new_n283), .ZN(new_n284));
  AOI21_X1  g0084(.A(new_n280), .B1(new_n274), .B2(new_n276), .ZN(new_n285));
  INV_X1    g0085(.A(KEYINPUT74), .ZN(new_n286));
  NOR3_X1   g0086(.A1(new_n285), .A2(new_n286), .A3(new_n262), .ZN(new_n287));
  OAI21_X1  g0087(.A(new_n266), .B1(new_n284), .B2(new_n287), .ZN(new_n288));
  INV_X1    g0088(.A(KEYINPUT75), .ZN(new_n289));
  NAND3_X1  g0089(.A1(new_n288), .A2(new_n289), .A3(KEYINPUT13), .ZN(new_n290));
  OAI21_X1  g0090(.A(new_n286), .B1(new_n285), .B2(new_n262), .ZN(new_n291));
  NAND3_X1  g0091(.A1(new_n282), .A2(KEYINPUT74), .A3(new_n283), .ZN(new_n292));
  AOI21_X1  g0092(.A(new_n265), .B1(new_n291), .B2(new_n292), .ZN(new_n293));
  INV_X1    g0093(.A(KEYINPUT13), .ZN(new_n294));
  OAI21_X1  g0094(.A(KEYINPUT75), .B1(new_n293), .B2(new_n294), .ZN(new_n295));
  AOI22_X1  g0095(.A1(new_n290), .A2(new_n295), .B1(new_n294), .B2(new_n293), .ZN(new_n296));
  INV_X1    g0096(.A(G169), .ZN(new_n297));
  AOI21_X1  g0097(.A(new_n297), .B1(KEYINPUT76), .B2(KEYINPUT14), .ZN(new_n298));
  INV_X1    g0098(.A(new_n298), .ZN(new_n299));
  OAI22_X1  g0099(.A1(new_n296), .A2(new_n299), .B1(KEYINPUT76), .B2(KEYINPUT14), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n293), .A2(new_n294), .ZN(new_n301));
  AOI21_X1  g0101(.A(new_n289), .B1(new_n288), .B2(KEYINPUT13), .ZN(new_n302));
  NOR3_X1   g0102(.A1(new_n293), .A2(KEYINPUT75), .A3(new_n294), .ZN(new_n303));
  OAI21_X1  g0103(.A(new_n301), .B1(new_n302), .B2(new_n303), .ZN(new_n304));
  NOR2_X1   g0104(.A1(KEYINPUT76), .A2(KEYINPUT14), .ZN(new_n305));
  NAND3_X1  g0105(.A1(new_n304), .A2(new_n298), .A3(new_n305), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n288), .A2(KEYINPUT13), .ZN(new_n307));
  NAND3_X1  g0107(.A1(new_n307), .A2(G179), .A3(new_n301), .ZN(new_n308));
  NAND3_X1  g0108(.A1(new_n300), .A2(new_n306), .A3(new_n308), .ZN(new_n309));
  NAND3_X1  g0109(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n310), .A2(new_n214), .ZN(new_n311));
  INV_X1    g0111(.A(new_n311), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n257), .A2(new_n258), .ZN(new_n313));
  OAI21_X1  g0113(.A(new_n312), .B1(new_n313), .B2(new_n215), .ZN(new_n314));
  INV_X1    g0114(.A(new_n314), .ZN(new_n315));
  NOR2_X1   g0115(.A1(G20), .A2(G33), .ZN(new_n316));
  INV_X1    g0116(.A(new_n316), .ZN(new_n317));
  OAI22_X1  g0117(.A1(new_n317), .A2(new_n202), .B1(new_n215), .B2(G68), .ZN(new_n318));
  INV_X1    g0118(.A(G77), .ZN(new_n319));
  NOR3_X1   g0119(.A1(new_n269), .A2(new_n319), .A3(G20), .ZN(new_n320));
  OAI21_X1  g0120(.A(new_n311), .B1(new_n318), .B2(new_n320), .ZN(new_n321));
  INV_X1    g0121(.A(KEYINPUT11), .ZN(new_n322));
  AOI22_X1  g0122(.A1(G68), .A2(new_n315), .B1(new_n321), .B2(new_n322), .ZN(new_n323));
  OAI21_X1  g0123(.A(new_n323), .B1(new_n322), .B2(new_n321), .ZN(new_n324));
  NAND4_X1  g0124(.A1(new_n257), .A2(G13), .A3(G20), .A4(new_n258), .ZN(new_n325));
  NOR2_X1   g0125(.A1(new_n325), .A2(G68), .ZN(new_n326));
  XNOR2_X1  g0126(.A(new_n326), .B(KEYINPUT12), .ZN(new_n327));
  NOR2_X1   g0127(.A1(new_n324), .A2(new_n327), .ZN(new_n328));
  INV_X1    g0128(.A(new_n328), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n309), .A2(new_n329), .ZN(new_n330));
  NAND3_X1  g0130(.A1(new_n307), .A2(G190), .A3(new_n301), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n331), .A2(new_n328), .ZN(new_n332));
  AOI21_X1  g0132(.A(new_n332), .B1(G200), .B2(new_n304), .ZN(new_n333));
  INV_X1    g0133(.A(new_n333), .ZN(new_n334));
  AOI21_X1  g0134(.A(new_n250), .B1(new_n330), .B2(new_n334), .ZN(new_n335));
  AOI211_X1 g0135(.A(KEYINPUT77), .B(new_n333), .C1(new_n309), .C2(new_n329), .ZN(new_n336));
  XNOR2_X1  g0136(.A(KEYINPUT70), .B(G58), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n337), .A2(G68), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n338), .A2(new_n211), .ZN(new_n339));
  AOI22_X1  g0139(.A1(new_n339), .A2(G20), .B1(G159), .B2(new_n316), .ZN(new_n340));
  OAI21_X1  g0140(.A(KEYINPUT79), .B1(new_n269), .B2(KEYINPUT3), .ZN(new_n341));
  INV_X1    g0141(.A(KEYINPUT79), .ZN(new_n342));
  NAND3_X1  g0142(.A1(new_n342), .A2(new_n267), .A3(G33), .ZN(new_n343));
  NAND2_X1  g0143(.A1(new_n341), .A2(new_n343), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n269), .A2(KEYINPUT78), .ZN(new_n345));
  INV_X1    g0145(.A(KEYINPUT78), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n346), .A2(G33), .ZN(new_n347));
  NAND3_X1  g0147(.A1(new_n345), .A2(new_n347), .A3(KEYINPUT3), .ZN(new_n348));
  AOI21_X1  g0148(.A(G20), .B1(new_n344), .B2(new_n348), .ZN(new_n349));
  INV_X1    g0149(.A(KEYINPUT7), .ZN(new_n350));
  OAI21_X1  g0150(.A(G68), .B1(new_n349), .B2(new_n350), .ZN(new_n351));
  XNOR2_X1  g0151(.A(KEYINPUT78), .B(G33), .ZN(new_n352));
  AOI22_X1  g0152(.A1(new_n352), .A2(KEYINPUT3), .B1(new_n341), .B2(new_n343), .ZN(new_n353));
  NOR3_X1   g0153(.A1(new_n353), .A2(KEYINPUT7), .A3(G20), .ZN(new_n354));
  OAI211_X1 g0154(.A(new_n340), .B(KEYINPUT16), .C1(new_n351), .C2(new_n354), .ZN(new_n355));
  INV_X1    g0155(.A(KEYINPUT16), .ZN(new_n356));
  INV_X1    g0156(.A(G68), .ZN(new_n357));
  NOR2_X1   g0157(.A1(new_n350), .A2(G20), .ZN(new_n358));
  AOI21_X1  g0158(.A(KEYINPUT3), .B1(new_n345), .B2(new_n347), .ZN(new_n359));
  INV_X1    g0159(.A(new_n270), .ZN(new_n360));
  OAI21_X1  g0160(.A(new_n358), .B1(new_n359), .B2(new_n360), .ZN(new_n361));
  OAI21_X1  g0161(.A(new_n350), .B1(new_n275), .B2(G20), .ZN(new_n362));
  AOI21_X1  g0162(.A(new_n357), .B1(new_n361), .B2(new_n362), .ZN(new_n363));
  AOI21_X1  g0163(.A(new_n201), .B1(new_n337), .B2(G68), .ZN(new_n364));
  INV_X1    g0164(.A(G159), .ZN(new_n365));
  OAI22_X1  g0165(.A1(new_n364), .A2(new_n215), .B1(new_n365), .B2(new_n317), .ZN(new_n366));
  OAI21_X1  g0166(.A(new_n356), .B1(new_n363), .B2(new_n366), .ZN(new_n367));
  NAND3_X1  g0167(.A1(new_n355), .A2(new_n367), .A3(new_n311), .ZN(new_n368));
  INV_X1    g0168(.A(G200), .ZN(new_n369));
  NAND3_X1  g0169(.A1(new_n259), .A2(G232), .A3(new_n262), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n370), .A2(KEYINPUT81), .ZN(new_n371));
  INV_X1    g0171(.A(KEYINPUT81), .ZN(new_n372));
  NAND4_X1  g0172(.A1(new_n259), .A2(new_n372), .A3(G232), .A4(new_n262), .ZN(new_n373));
  NAND3_X1  g0173(.A1(new_n371), .A2(new_n256), .A3(new_n373), .ZN(new_n374));
  NAND2_X1  g0174(.A1(G226), .A2(G1698), .ZN(new_n375));
  INV_X1    g0175(.A(G223), .ZN(new_n376));
  OAI21_X1  g0176(.A(new_n375), .B1(new_n376), .B2(G1698), .ZN(new_n377));
  NAND3_X1  g0177(.A1(new_n344), .A2(new_n348), .A3(new_n377), .ZN(new_n378));
  NAND2_X1  g0178(.A1(G33), .A2(G87), .ZN(new_n379));
  AOI21_X1  g0179(.A(new_n262), .B1(new_n378), .B2(new_n379), .ZN(new_n380));
  OAI21_X1  g0180(.A(new_n369), .B1(new_n374), .B2(new_n380), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n378), .A2(new_n379), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n382), .A2(new_n283), .ZN(new_n383));
  AND2_X1   g0183(.A1(new_n256), .A2(new_n373), .ZN(new_n384));
  INV_X1    g0184(.A(G190), .ZN(new_n385));
  NAND4_X1  g0185(.A1(new_n383), .A2(new_n384), .A3(new_n385), .A4(new_n371), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n381), .A2(new_n386), .ZN(new_n387));
  NOR2_X1   g0187(.A1(KEYINPUT8), .A2(G58), .ZN(new_n388));
  AOI21_X1  g0188(.A(new_n388), .B1(new_n337), .B2(KEYINPUT8), .ZN(new_n389));
  INV_X1    g0189(.A(new_n325), .ZN(new_n390));
  OR2_X1    g0190(.A1(new_n389), .A2(new_n390), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n314), .A2(new_n389), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n391), .A2(new_n392), .ZN(new_n393));
  NAND3_X1  g0193(.A1(new_n368), .A2(new_n387), .A3(new_n393), .ZN(new_n394));
  INV_X1    g0194(.A(KEYINPUT82), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n394), .A2(new_n395), .ZN(new_n396));
  NAND4_X1  g0196(.A1(new_n368), .A2(new_n387), .A3(KEYINPUT82), .A4(new_n393), .ZN(new_n397));
  NAND3_X1  g0197(.A1(new_n396), .A2(KEYINPUT17), .A3(new_n397), .ZN(new_n398));
  OR2_X1    g0198(.A1(new_n394), .A2(KEYINPUT17), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n398), .A2(new_n399), .ZN(new_n400));
  INV_X1    g0200(.A(KEYINPUT80), .ZN(new_n401));
  AND3_X1   g0201(.A1(new_n368), .A2(new_n401), .A3(new_n393), .ZN(new_n402));
  AOI21_X1  g0202(.A(new_n401), .B1(new_n368), .B2(new_n393), .ZN(new_n403));
  NOR2_X1   g0203(.A1(new_n402), .A2(new_n403), .ZN(new_n404));
  NOR2_X1   g0204(.A1(new_n374), .A2(new_n380), .ZN(new_n405));
  NOR2_X1   g0205(.A1(new_n405), .A2(G169), .ZN(new_n406));
  INV_X1    g0206(.A(G179), .ZN(new_n407));
  AOI21_X1  g0207(.A(new_n406), .B1(new_n407), .B2(new_n405), .ZN(new_n408));
  AOI21_X1  g0208(.A(KEYINPUT18), .B1(new_n404), .B2(new_n408), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n368), .A2(new_n393), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n410), .A2(KEYINPUT80), .ZN(new_n411));
  NAND3_X1  g0211(.A1(new_n368), .A2(new_n401), .A3(new_n393), .ZN(new_n412));
  AND4_X1   g0212(.A1(KEYINPUT18), .A2(new_n411), .A3(new_n412), .A4(new_n408), .ZN(new_n413));
  INV_X1    g0213(.A(KEYINPUT72), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n275), .A2(G1698), .ZN(new_n415));
  INV_X1    g0215(.A(new_n225), .ZN(new_n416));
  OAI22_X1  g0216(.A1(new_n415), .A2(new_n376), .B1(new_n416), .B2(new_n275), .ZN(new_n417));
  INV_X1    g0217(.A(new_n417), .ZN(new_n418));
  NAND3_X1  g0218(.A1(new_n275), .A2(G222), .A3(new_n271), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n419), .A2(KEYINPUT69), .ZN(new_n420));
  INV_X1    g0220(.A(KEYINPUT69), .ZN(new_n421));
  NAND4_X1  g0221(.A1(new_n275), .A2(new_n421), .A3(G222), .A4(new_n271), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n420), .A2(new_n422), .ZN(new_n423));
  AOI21_X1  g0223(.A(new_n262), .B1(new_n418), .B2(new_n423), .ZN(new_n424));
  INV_X1    g0224(.A(G226), .ZN(new_n425));
  OAI21_X1  g0225(.A(new_n256), .B1(new_n263), .B2(new_n425), .ZN(new_n426));
  OAI21_X1  g0226(.A(G200), .B1(new_n424), .B2(new_n426), .ZN(new_n427));
  INV_X1    g0227(.A(new_n426), .ZN(new_n428));
  AOI21_X1  g0228(.A(new_n417), .B1(new_n422), .B2(new_n420), .ZN(new_n429));
  OAI211_X1 g0229(.A(G190), .B(new_n428), .C1(new_n429), .C2(new_n262), .ZN(new_n430));
  INV_X1    g0230(.A(KEYINPUT9), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n314), .A2(G50), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n325), .A2(new_n202), .ZN(new_n433));
  AND2_X1   g0233(.A1(new_n432), .A2(new_n433), .ZN(new_n434));
  NOR2_X1   g0234(.A1(new_n269), .A2(G20), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n389), .A2(new_n435), .ZN(new_n436));
  AOI22_X1  g0236(.A1(new_n203), .A2(G20), .B1(G150), .B2(new_n316), .ZN(new_n437));
  AOI21_X1  g0237(.A(new_n312), .B1(new_n436), .B2(new_n437), .ZN(new_n438));
  OAI21_X1  g0238(.A(new_n431), .B1(new_n434), .B2(new_n438), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n432), .A2(new_n433), .ZN(new_n440));
  INV_X1    g0240(.A(new_n437), .ZN(new_n441));
  AOI21_X1  g0241(.A(new_n441), .B1(new_n389), .B2(new_n435), .ZN(new_n442));
  OAI211_X1 g0242(.A(KEYINPUT9), .B(new_n440), .C1(new_n442), .C2(new_n312), .ZN(new_n443));
  NAND4_X1  g0243(.A1(new_n427), .A2(new_n430), .A3(new_n439), .A4(new_n443), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n444), .A2(KEYINPUT10), .ZN(new_n445));
  AND2_X1   g0245(.A1(new_n439), .A2(new_n443), .ZN(new_n446));
  INV_X1    g0246(.A(KEYINPUT10), .ZN(new_n447));
  NAND4_X1  g0247(.A1(new_n446), .A2(new_n447), .A3(new_n430), .A4(new_n427), .ZN(new_n448));
  NAND2_X1  g0248(.A1(new_n445), .A2(new_n448), .ZN(new_n449));
  NOR2_X1   g0249(.A1(new_n434), .A2(new_n438), .ZN(new_n450));
  OAI21_X1  g0250(.A(G169), .B1(new_n424), .B2(new_n426), .ZN(new_n451));
  OAI211_X1 g0251(.A(G179), .B(new_n428), .C1(new_n429), .C2(new_n262), .ZN(new_n452));
  AOI21_X1  g0252(.A(new_n450), .B1(new_n451), .B2(new_n452), .ZN(new_n453));
  INV_X1    g0253(.A(new_n453), .ZN(new_n454));
  INV_X1    g0254(.A(new_n256), .ZN(new_n455));
  INV_X1    g0255(.A(new_n263), .ZN(new_n456));
  AOI21_X1  g0256(.A(new_n455), .B1(new_n456), .B2(G244), .ZN(new_n457));
  NAND3_X1  g0257(.A1(new_n275), .A2(G232), .A3(new_n271), .ZN(new_n458));
  INV_X1    g0258(.A(G107), .ZN(new_n459));
  OAI221_X1 g0259(.A(new_n458), .B1(new_n459), .B2(new_n275), .C1(new_n415), .C2(new_n264), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n460), .A2(new_n283), .ZN(new_n461));
  NAND2_X1  g0261(.A1(new_n457), .A2(new_n461), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n462), .A2(G200), .ZN(new_n463));
  XOR2_X1   g0263(.A(KEYINPUT8), .B(G58), .Z(new_n464));
  AOI22_X1  g0264(.A1(new_n464), .A2(new_n316), .B1(new_n225), .B2(G20), .ZN(new_n465));
  XNOR2_X1  g0265(.A(KEYINPUT15), .B(G87), .ZN(new_n466));
  INV_X1    g0266(.A(new_n466), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n467), .A2(new_n435), .ZN(new_n468));
  AOI21_X1  g0268(.A(new_n312), .B1(new_n465), .B2(new_n468), .ZN(new_n469));
  OAI22_X1  g0269(.A1(new_n314), .A2(new_n319), .B1(new_n225), .B2(new_n325), .ZN(new_n470));
  NOR2_X1   g0270(.A1(new_n469), .A2(new_n470), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n471), .A2(KEYINPUT71), .ZN(new_n472));
  NAND3_X1  g0272(.A1(new_n457), .A2(new_n461), .A3(G190), .ZN(new_n473));
  INV_X1    g0273(.A(KEYINPUT71), .ZN(new_n474));
  OAI21_X1  g0274(.A(new_n474), .B1(new_n469), .B2(new_n470), .ZN(new_n475));
  NAND4_X1  g0275(.A1(new_n463), .A2(new_n472), .A3(new_n473), .A4(new_n475), .ZN(new_n476));
  AND3_X1   g0276(.A1(new_n457), .A2(new_n461), .A3(G179), .ZN(new_n477));
  AOI21_X1  g0277(.A(new_n297), .B1(new_n457), .B2(new_n461), .ZN(new_n478));
  OAI22_X1  g0278(.A1(new_n477), .A2(new_n478), .B1(new_n469), .B2(new_n470), .ZN(new_n479));
  AND2_X1   g0279(.A1(new_n476), .A2(new_n479), .ZN(new_n480));
  AND4_X1   g0280(.A1(new_n414), .A2(new_n449), .A3(new_n454), .A4(new_n480), .ZN(new_n481));
  AOI21_X1  g0281(.A(new_n453), .B1(new_n445), .B2(new_n448), .ZN(new_n482));
  AOI21_X1  g0282(.A(new_n414), .B1(new_n482), .B2(new_n480), .ZN(new_n483));
  OAI221_X1 g0283(.A(new_n400), .B1(new_n409), .B2(new_n413), .C1(new_n481), .C2(new_n483), .ZN(new_n484));
  NOR3_X1   g0284(.A1(new_n335), .A2(new_n336), .A3(new_n484), .ZN(new_n485));
  NAND2_X1  g0285(.A1(G257), .A2(G1698), .ZN(new_n486));
  INV_X1    g0286(.A(G250), .ZN(new_n487));
  OAI21_X1  g0287(.A(new_n486), .B1(new_n487), .B2(G1698), .ZN(new_n488));
  NAND3_X1  g0288(.A1(new_n344), .A2(new_n348), .A3(new_n488), .ZN(new_n489));
  XOR2_X1   g0289(.A(KEYINPUT91), .B(G294), .Z(new_n490));
  NAND2_X1  g0290(.A1(new_n345), .A2(new_n347), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  AOI21_X1  g0292(.A(new_n262), .B1(new_n489), .B2(new_n492), .ZN(new_n493));
  NAND3_X1  g0293(.A1(new_n257), .A2(G45), .A3(new_n258), .ZN(new_n494));
  AND2_X1   g0294(.A1(KEYINPUT5), .A2(G41), .ZN(new_n495));
  NOR2_X1   g0295(.A1(KEYINPUT5), .A2(G41), .ZN(new_n496));
  NOR2_X1   g0296(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  OAI211_X1 g0297(.A(G264), .B(new_n262), .C1(new_n494), .C2(new_n497), .ZN(new_n498));
  INV_X1    g0298(.A(new_n498), .ZN(new_n499));
  XOR2_X1   g0299(.A(KEYINPUT68), .B(G1), .Z(new_n500));
  AOI21_X1  g0300(.A(new_n255), .B1(new_n260), .B2(new_n261), .ZN(new_n501));
  XNOR2_X1  g0301(.A(KEYINPUT5), .B(G41), .ZN(new_n502));
  NAND4_X1  g0302(.A1(new_n500), .A2(new_n501), .A3(G45), .A4(new_n502), .ZN(new_n503));
  INV_X1    g0303(.A(new_n503), .ZN(new_n504));
  NOR3_X1   g0304(.A1(new_n493), .A2(new_n499), .A3(new_n504), .ZN(new_n505));
  INV_X1    g0305(.A(new_n505), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n506), .A2(G169), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n505), .A2(G179), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  INV_X1    g0309(.A(KEYINPUT24), .ZN(new_n510));
  INV_X1    g0310(.A(KEYINPUT90), .ZN(new_n511));
  INV_X1    g0311(.A(G87), .ZN(new_n512));
  NOR2_X1   g0312(.A1(new_n512), .A2(G20), .ZN(new_n513));
  NAND3_X1  g0313(.A1(new_n513), .A2(new_n268), .A3(new_n270), .ZN(new_n514));
  INV_X1    g0314(.A(KEYINPUT22), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  NOR2_X1   g0316(.A1(new_n346), .A2(G33), .ZN(new_n517));
  NOR2_X1   g0317(.A1(new_n269), .A2(KEYINPUT78), .ZN(new_n518));
  OAI211_X1 g0318(.A(new_n215), .B(G116), .C1(new_n517), .C2(new_n518), .ZN(new_n519));
  OAI21_X1  g0319(.A(KEYINPUT23), .B1(new_n215), .B2(G107), .ZN(new_n520));
  INV_X1    g0320(.A(KEYINPUT23), .ZN(new_n521));
  NAND3_X1  g0321(.A1(new_n521), .A2(new_n459), .A3(G20), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n520), .A2(new_n522), .ZN(new_n523));
  INV_X1    g0323(.A(new_n523), .ZN(new_n524));
  AND3_X1   g0324(.A1(new_n516), .A2(new_n519), .A3(new_n524), .ZN(new_n525));
  NOR2_X1   g0325(.A1(new_n515), .A2(new_n512), .ZN(new_n526));
  NAND4_X1  g0326(.A1(new_n344), .A2(new_n348), .A3(new_n215), .A4(new_n526), .ZN(new_n527));
  AOI21_X1  g0327(.A(new_n511), .B1(new_n525), .B2(new_n527), .ZN(new_n528));
  INV_X1    g0328(.A(G116), .ZN(new_n529));
  AOI21_X1  g0329(.A(new_n529), .B1(new_n345), .B2(new_n347), .ZN(new_n530));
  AOI21_X1  g0330(.A(new_n523), .B1(new_n530), .B2(new_n215), .ZN(new_n531));
  AND4_X1   g0331(.A1(new_n511), .A2(new_n531), .A3(new_n527), .A4(new_n516), .ZN(new_n532));
  OAI21_X1  g0332(.A(new_n510), .B1(new_n528), .B2(new_n532), .ZN(new_n533));
  NAND3_X1  g0333(.A1(new_n525), .A2(new_n511), .A3(new_n527), .ZN(new_n534));
  NAND3_X1  g0334(.A1(new_n531), .A2(new_n527), .A3(new_n516), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n535), .A2(KEYINPUT90), .ZN(new_n536));
  NAND3_X1  g0336(.A1(new_n534), .A2(new_n536), .A3(KEYINPUT24), .ZN(new_n537));
  NAND3_X1  g0337(.A1(new_n533), .A2(new_n311), .A3(new_n537), .ZN(new_n538));
  INV_X1    g0338(.A(new_n538), .ZN(new_n539));
  NAND3_X1  g0339(.A1(new_n257), .A2(G33), .A3(new_n258), .ZN(new_n540));
  NAND3_X1  g0340(.A1(new_n325), .A2(new_n312), .A3(new_n540), .ZN(new_n541));
  INV_X1    g0341(.A(new_n541), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n542), .A2(G107), .ZN(new_n543));
  OR3_X1    g0343(.A1(new_n325), .A2(KEYINPUT25), .A3(G107), .ZN(new_n544));
  OAI21_X1  g0344(.A(KEYINPUT25), .B1(new_n325), .B2(G107), .ZN(new_n545));
  NAND3_X1  g0345(.A1(new_n543), .A2(new_n544), .A3(new_n545), .ZN(new_n546));
  OAI21_X1  g0346(.A(new_n509), .B1(new_n539), .B2(new_n546), .ZN(new_n547));
  INV_X1    g0347(.A(new_n546), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n505), .A2(new_n385), .ZN(new_n549));
  OAI21_X1  g0349(.A(new_n549), .B1(G200), .B2(new_n505), .ZN(new_n550));
  NAND3_X1  g0350(.A1(new_n538), .A2(new_n548), .A3(new_n550), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n547), .A2(new_n551), .ZN(new_n552));
  NAND2_X1  g0352(.A1(G264), .A2(G1698), .ZN(new_n553));
  OAI21_X1  g0353(.A(new_n553), .B1(new_n222), .B2(G1698), .ZN(new_n554));
  NAND3_X1  g0354(.A1(new_n344), .A2(new_n348), .A3(new_n554), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n268), .A2(new_n270), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n556), .A2(G303), .ZN(new_n557));
  AOI21_X1  g0357(.A(new_n262), .B1(new_n555), .B2(new_n557), .ZN(new_n558));
  OAI211_X1 g0358(.A(G270), .B(new_n262), .C1(new_n494), .C2(new_n497), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n559), .A2(new_n503), .ZN(new_n560));
  OAI21_X1  g0360(.A(G169), .B1(new_n558), .B2(new_n560), .ZN(new_n561));
  NAND2_X1  g0361(.A1(G33), .A2(G283), .ZN(new_n562));
  OAI21_X1  g0362(.A(new_n562), .B1(new_n221), .B2(G33), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n563), .A2(new_n215), .ZN(new_n564));
  NOR2_X1   g0364(.A1(new_n215), .A2(new_n529), .ZN(new_n565));
  INV_X1    g0365(.A(new_n565), .ZN(new_n566));
  AOI21_X1  g0366(.A(new_n312), .B1(new_n564), .B2(new_n566), .ZN(new_n567));
  NAND3_X1  g0367(.A1(new_n567), .A2(KEYINPUT88), .A3(KEYINPUT20), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n269), .A2(G97), .ZN(new_n569));
  AOI21_X1  g0369(.A(G20), .B1(new_n569), .B2(new_n562), .ZN(new_n570));
  OAI211_X1 g0370(.A(KEYINPUT20), .B(new_n311), .C1(new_n570), .C2(new_n565), .ZN(new_n571));
  INV_X1    g0371(.A(KEYINPUT88), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n571), .A2(new_n572), .ZN(new_n573));
  INV_X1    g0373(.A(KEYINPUT20), .ZN(new_n574));
  AOI21_X1  g0374(.A(new_n565), .B1(new_n563), .B2(new_n215), .ZN(new_n575));
  OAI21_X1  g0375(.A(new_n574), .B1(new_n575), .B2(new_n312), .ZN(new_n576));
  NAND3_X1  g0376(.A1(new_n568), .A2(new_n573), .A3(new_n576), .ZN(new_n577));
  NOR2_X1   g0377(.A1(new_n325), .A2(G116), .ZN(new_n578));
  AOI21_X1  g0378(.A(new_n578), .B1(new_n542), .B2(G116), .ZN(new_n579));
  AOI21_X1  g0379(.A(new_n561), .B1(new_n577), .B2(new_n579), .ZN(new_n580));
  OAI21_X1  g0380(.A(KEYINPUT89), .B1(new_n580), .B2(KEYINPUT21), .ZN(new_n581));
  INV_X1    g0381(.A(new_n561), .ZN(new_n582));
  OAI21_X1  g0382(.A(new_n576), .B1(new_n572), .B2(new_n571), .ZN(new_n583));
  AOI21_X1  g0383(.A(KEYINPUT88), .B1(new_n567), .B2(KEYINPUT20), .ZN(new_n584));
  OAI21_X1  g0384(.A(new_n579), .B1(new_n583), .B2(new_n584), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n582), .A2(new_n585), .ZN(new_n586));
  INV_X1    g0386(.A(KEYINPUT89), .ZN(new_n587));
  INV_X1    g0387(.A(KEYINPUT21), .ZN(new_n588));
  NAND3_X1  g0388(.A1(new_n586), .A2(new_n587), .A3(new_n588), .ZN(new_n589));
  NOR2_X1   g0389(.A1(new_n558), .A2(new_n560), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n590), .A2(G179), .ZN(new_n591));
  OAI21_X1  g0391(.A(new_n591), .B1(new_n588), .B2(new_n561), .ZN(new_n592));
  AOI22_X1  g0392(.A1(new_n581), .A2(new_n589), .B1(new_n585), .B2(new_n592), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n590), .A2(new_n385), .ZN(new_n594));
  OAI21_X1  g0394(.A(new_n594), .B1(G200), .B2(new_n590), .ZN(new_n595));
  INV_X1    g0395(.A(new_n585), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n595), .A2(new_n596), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n593), .A2(new_n597), .ZN(new_n598));
  INV_X1    g0398(.A(KEYINPUT84), .ZN(new_n599));
  INV_X1    g0399(.A(new_n358), .ZN(new_n600));
  OAI21_X1  g0400(.A(new_n267), .B1(new_n517), .B2(new_n518), .ZN(new_n601));
  AOI21_X1  g0401(.A(new_n600), .B1(new_n601), .B2(new_n270), .ZN(new_n602));
  AOI21_X1  g0402(.A(KEYINPUT7), .B1(new_n556), .B2(new_n215), .ZN(new_n603));
  OAI21_X1  g0403(.A(G107), .B1(new_n602), .B2(new_n603), .ZN(new_n604));
  XNOR2_X1  g0404(.A(G97), .B(G107), .ZN(new_n605));
  INV_X1    g0405(.A(KEYINPUT6), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n605), .A2(new_n606), .ZN(new_n607));
  INV_X1    g0407(.A(KEYINPUT83), .ZN(new_n608));
  NAND2_X1  g0408(.A1(KEYINPUT6), .A2(G97), .ZN(new_n609));
  OAI21_X1  g0409(.A(new_n608), .B1(new_n609), .B2(G107), .ZN(new_n610));
  NAND4_X1  g0410(.A1(new_n459), .A2(KEYINPUT83), .A3(KEYINPUT6), .A4(G97), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n607), .A2(new_n612), .ZN(new_n613));
  AOI22_X1  g0413(.A1(new_n613), .A2(G20), .B1(G77), .B2(new_n316), .ZN(new_n614));
  AOI21_X1  g0414(.A(new_n312), .B1(new_n604), .B2(new_n614), .ZN(new_n615));
  NOR2_X1   g0415(.A1(new_n325), .A2(G97), .ZN(new_n616));
  AOI21_X1  g0416(.A(new_n616), .B1(new_n542), .B2(G97), .ZN(new_n617));
  INV_X1    g0417(.A(new_n617), .ZN(new_n618));
  OAI21_X1  g0418(.A(new_n599), .B1(new_n615), .B2(new_n618), .ZN(new_n619));
  AOI21_X1  g0419(.A(new_n459), .B1(new_n361), .B2(new_n362), .ZN(new_n620));
  AOI22_X1  g0420(.A1(new_n606), .A2(new_n605), .B1(new_n610), .B2(new_n611), .ZN(new_n621));
  OAI22_X1  g0421(.A1(new_n621), .A2(new_n215), .B1(new_n319), .B2(new_n317), .ZN(new_n622));
  OAI21_X1  g0422(.A(new_n311), .B1(new_n620), .B2(new_n622), .ZN(new_n623));
  NAND3_X1  g0423(.A1(new_n623), .A2(KEYINPUT84), .A3(new_n617), .ZN(new_n624));
  NAND4_X1  g0424(.A1(new_n344), .A2(new_n348), .A3(G244), .A4(new_n271), .ZN(new_n625));
  INV_X1    g0425(.A(KEYINPUT4), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  AND2_X1   g0427(.A1(KEYINPUT4), .A2(G244), .ZN(new_n628));
  NAND4_X1  g0428(.A1(new_n268), .A2(new_n270), .A3(new_n628), .A4(new_n271), .ZN(new_n629));
  INV_X1    g0429(.A(KEYINPUT85), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  NAND4_X1  g0431(.A1(new_n275), .A2(KEYINPUT85), .A3(new_n271), .A4(new_n628), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n631), .A2(new_n632), .ZN(new_n633));
  NAND4_X1  g0433(.A1(new_n268), .A2(new_n270), .A3(G250), .A4(G1698), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n634), .A2(new_n562), .ZN(new_n635));
  INV_X1    g0435(.A(new_n635), .ZN(new_n636));
  NAND3_X1  g0436(.A1(new_n627), .A2(new_n633), .A3(new_n636), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n637), .A2(new_n283), .ZN(new_n638));
  NAND3_X1  g0438(.A1(new_n500), .A2(G45), .A3(new_n502), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n639), .A2(new_n262), .ZN(new_n640));
  OAI21_X1  g0440(.A(new_n503), .B1(new_n640), .B2(new_n222), .ZN(new_n641));
  INV_X1    g0441(.A(new_n641), .ZN(new_n642));
  AOI21_X1  g0442(.A(G200), .B1(new_n638), .B2(new_n642), .ZN(new_n643));
  AOI21_X1  g0443(.A(new_n635), .B1(new_n631), .B2(new_n632), .ZN(new_n644));
  AOI21_X1  g0444(.A(new_n262), .B1(new_n644), .B2(new_n627), .ZN(new_n645));
  NOR3_X1   g0445(.A1(new_n645), .A2(G190), .A3(new_n641), .ZN(new_n646));
  OAI211_X1 g0446(.A(new_n619), .B(new_n624), .C1(new_n643), .C2(new_n646), .ZN(new_n647));
  NAND3_X1  g0447(.A1(new_n638), .A2(new_n407), .A3(new_n642), .ZN(new_n648));
  OAI21_X1  g0448(.A(new_n297), .B1(new_n645), .B2(new_n641), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n623), .A2(new_n617), .ZN(new_n650));
  NAND3_X1  g0450(.A1(new_n648), .A2(new_n649), .A3(new_n650), .ZN(new_n651));
  NOR2_X1   g0451(.A1(new_n467), .A2(new_n325), .ZN(new_n652));
  NAND4_X1  g0452(.A1(new_n344), .A2(new_n348), .A3(new_n215), .A4(G68), .ZN(new_n653));
  NOR2_X1   g0453(.A1(G87), .A2(G97), .ZN(new_n654));
  AOI22_X1  g0454(.A1(new_n654), .A2(new_n459), .B1(new_n279), .B2(new_n215), .ZN(new_n655));
  INV_X1    g0455(.A(KEYINPUT19), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n656), .A2(new_n215), .ZN(new_n657));
  OAI22_X1  g0457(.A1(new_n655), .A2(new_n656), .B1(new_n279), .B2(new_n657), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n653), .A2(new_n658), .ZN(new_n659));
  AOI21_X1  g0459(.A(new_n652), .B1(new_n659), .B2(new_n311), .ZN(new_n660));
  OAI21_X1  g0460(.A(new_n660), .B1(new_n466), .B2(new_n541), .ZN(new_n661));
  NAND4_X1  g0461(.A1(new_n344), .A2(new_n348), .A3(G244), .A4(G1698), .ZN(new_n662));
  NOR2_X1   g0462(.A1(new_n264), .A2(G1698), .ZN(new_n663));
  NAND3_X1  g0463(.A1(new_n344), .A2(new_n348), .A3(new_n663), .ZN(new_n664));
  INV_X1    g0464(.A(new_n530), .ZN(new_n665));
  NAND3_X1  g0465(.A1(new_n662), .A2(new_n664), .A3(new_n665), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n666), .A2(new_n283), .ZN(new_n667));
  INV_X1    g0467(.A(KEYINPUT86), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n262), .A2(G274), .ZN(new_n669));
  OAI21_X1  g0469(.A(new_n668), .B1(new_n669), .B2(new_n494), .ZN(new_n670));
  NAND4_X1  g0470(.A1(new_n500), .A2(new_n501), .A3(KEYINPUT86), .A4(G45), .ZN(new_n671));
  NOR2_X1   g0471(.A1(new_n283), .A2(new_n487), .ZN(new_n672));
  AOI22_X1  g0472(.A1(new_n670), .A2(new_n671), .B1(new_n672), .B2(new_n494), .ZN(new_n673));
  NAND3_X1  g0473(.A1(new_n667), .A2(new_n673), .A3(new_n407), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n667), .A2(new_n673), .ZN(new_n675));
  INV_X1    g0475(.A(new_n675), .ZN(new_n676));
  OAI211_X1 g0476(.A(new_n661), .B(new_n674), .C1(new_n676), .C2(G169), .ZN(new_n677));
  NAND3_X1  g0477(.A1(new_n667), .A2(new_n673), .A3(G190), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n678), .A2(KEYINPUT87), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n675), .A2(G200), .ZN(new_n680));
  INV_X1    g0480(.A(KEYINPUT87), .ZN(new_n681));
  NAND4_X1  g0481(.A1(new_n667), .A2(new_n673), .A3(new_n681), .A4(G190), .ZN(new_n682));
  AOI21_X1  g0482(.A(new_n312), .B1(new_n653), .B2(new_n658), .ZN(new_n683));
  NOR2_X1   g0483(.A1(new_n541), .A2(new_n512), .ZN(new_n684));
  NOR3_X1   g0484(.A1(new_n683), .A2(new_n652), .A3(new_n684), .ZN(new_n685));
  NAND4_X1  g0485(.A1(new_n679), .A2(new_n680), .A3(new_n682), .A4(new_n685), .ZN(new_n686));
  NAND4_X1  g0486(.A1(new_n647), .A2(new_n651), .A3(new_n677), .A4(new_n686), .ZN(new_n687));
  NOR3_X1   g0487(.A1(new_n552), .A2(new_n598), .A3(new_n687), .ZN(new_n688));
  AND2_X1   g0488(.A1(new_n485), .A2(new_n688), .ZN(G372));
  AND2_X1   g0489(.A1(new_n647), .A2(new_n651), .ZN(new_n690));
  INV_X1    g0490(.A(KEYINPUT93), .ZN(new_n691));
  INV_X1    g0491(.A(new_n684), .ZN(new_n692));
  AOI21_X1  g0492(.A(KEYINPUT92), .B1(new_n660), .B2(new_n692), .ZN(new_n693));
  INV_X1    g0493(.A(KEYINPUT92), .ZN(new_n694));
  NOR4_X1   g0494(.A1(new_n683), .A2(new_n684), .A3(new_n694), .A4(new_n652), .ZN(new_n695));
  OAI211_X1 g0495(.A(new_n680), .B(new_n678), .C1(new_n693), .C2(new_n695), .ZN(new_n696));
  AND2_X1   g0496(.A1(new_n696), .A2(new_n677), .ZN(new_n697));
  NAND4_X1  g0497(.A1(new_n690), .A2(new_n691), .A3(new_n551), .A4(new_n697), .ZN(new_n698));
  NAND3_X1  g0498(.A1(new_n551), .A2(new_n647), .A3(new_n651), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n696), .A2(new_n677), .ZN(new_n700));
  OAI21_X1  g0500(.A(KEYINPUT93), .B1(new_n699), .B2(new_n700), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n592), .A2(new_n585), .ZN(new_n702));
  AOI21_X1  g0502(.A(new_n587), .B1(new_n586), .B2(new_n588), .ZN(new_n703));
  AOI211_X1 g0503(.A(KEYINPUT89), .B(KEYINPUT21), .C1(new_n582), .C2(new_n585), .ZN(new_n704));
  OAI21_X1  g0504(.A(new_n702), .B1(new_n703), .B2(new_n704), .ZN(new_n705));
  AOI22_X1  g0505(.A1(new_n538), .A2(new_n548), .B1(new_n508), .B2(new_n507), .ZN(new_n706));
  OAI21_X1  g0506(.A(KEYINPUT94), .B1(new_n705), .B2(new_n706), .ZN(new_n707));
  INV_X1    g0507(.A(KEYINPUT94), .ZN(new_n708));
  NAND3_X1  g0508(.A1(new_n547), .A2(new_n593), .A3(new_n708), .ZN(new_n709));
  NAND4_X1  g0509(.A1(new_n698), .A2(new_n701), .A3(new_n707), .A4(new_n709), .ZN(new_n710));
  NAND2_X1  g0510(.A1(new_n648), .A2(new_n649), .ZN(new_n711));
  AOI21_X1  g0511(.A(new_n711), .B1(new_n619), .B2(new_n624), .ZN(new_n712));
  INV_X1    g0512(.A(KEYINPUT26), .ZN(new_n713));
  NAND3_X1  g0513(.A1(new_n697), .A2(new_n712), .A3(new_n713), .ZN(new_n714));
  AND3_X1   g0514(.A1(new_n648), .A2(new_n650), .A3(new_n649), .ZN(new_n715));
  NAND3_X1  g0515(.A1(new_n715), .A2(new_n677), .A3(new_n686), .ZN(new_n716));
  NAND2_X1  g0516(.A1(new_n716), .A2(KEYINPUT26), .ZN(new_n717));
  NAND3_X1  g0517(.A1(new_n714), .A2(new_n717), .A3(new_n677), .ZN(new_n718));
  INV_X1    g0518(.A(KEYINPUT95), .ZN(new_n719));
  NAND2_X1  g0519(.A1(new_n718), .A2(new_n719), .ZN(new_n720));
  NAND4_X1  g0520(.A1(new_n714), .A2(new_n717), .A3(KEYINPUT95), .A4(new_n677), .ZN(new_n721));
  NAND3_X1  g0521(.A1(new_n710), .A2(new_n720), .A3(new_n721), .ZN(new_n722));
  NAND2_X1  g0522(.A1(new_n485), .A2(new_n722), .ZN(new_n723));
  NAND2_X1  g0523(.A1(new_n408), .A2(new_n410), .ZN(new_n724));
  INV_X1    g0524(.A(KEYINPUT18), .ZN(new_n725));
  XNOR2_X1  g0525(.A(new_n724), .B(new_n725), .ZN(new_n726));
  INV_X1    g0526(.A(new_n479), .ZN(new_n727));
  AOI22_X1  g0527(.A1(new_n309), .A2(new_n329), .B1(new_n334), .B2(new_n727), .ZN(new_n728));
  INV_X1    g0528(.A(new_n400), .ZN(new_n729));
  OAI21_X1  g0529(.A(new_n726), .B1(new_n728), .B2(new_n729), .ZN(new_n730));
  AOI21_X1  g0530(.A(new_n453), .B1(new_n730), .B2(new_n449), .ZN(new_n731));
  NAND2_X1  g0531(.A1(new_n723), .A2(new_n731), .ZN(G369));
  AND2_X1   g0532(.A1(new_n215), .A2(G13), .ZN(new_n733));
  NAND2_X1  g0533(.A1(new_n500), .A2(new_n733), .ZN(new_n734));
  OR2_X1    g0534(.A1(new_n734), .A2(KEYINPUT27), .ZN(new_n735));
  NAND2_X1  g0535(.A1(new_n734), .A2(KEYINPUT27), .ZN(new_n736));
  AND3_X1   g0536(.A1(new_n735), .A2(G213), .A3(new_n736), .ZN(new_n737));
  NAND2_X1  g0537(.A1(new_n737), .A2(G343), .ZN(new_n738));
  NOR2_X1   g0538(.A1(new_n596), .A2(new_n738), .ZN(new_n739));
  NAND2_X1  g0539(.A1(new_n705), .A2(new_n739), .ZN(new_n740));
  OAI21_X1  g0540(.A(new_n740), .B1(new_n598), .B2(new_n739), .ZN(new_n741));
  XNOR2_X1  g0541(.A(new_n741), .B(KEYINPUT96), .ZN(new_n742));
  NAND2_X1  g0542(.A1(new_n742), .A2(G330), .ZN(new_n743));
  INV_X1    g0543(.A(new_n743), .ZN(new_n744));
  INV_X1    g0544(.A(new_n738), .ZN(new_n745));
  OAI21_X1  g0545(.A(new_n745), .B1(new_n539), .B2(new_n546), .ZN(new_n746));
  AOI21_X1  g0546(.A(new_n706), .B1(new_n746), .B2(new_n551), .ZN(new_n747));
  NAND2_X1  g0547(.A1(new_n706), .A2(new_n738), .ZN(new_n748));
  INV_X1    g0548(.A(new_n748), .ZN(new_n749));
  NOR2_X1   g0549(.A1(new_n747), .A2(new_n749), .ZN(new_n750));
  NAND2_X1  g0550(.A1(new_n744), .A2(new_n750), .ZN(new_n751));
  NOR2_X1   g0551(.A1(new_n593), .A2(new_n745), .ZN(new_n752));
  AND2_X1   g0552(.A1(new_n750), .A2(new_n752), .ZN(new_n753));
  NOR2_X1   g0553(.A1(new_n753), .A2(new_n749), .ZN(new_n754));
  NAND2_X1  g0554(.A1(new_n751), .A2(new_n754), .ZN(G399));
  INV_X1    g0555(.A(new_n208), .ZN(new_n756));
  NOR2_X1   g0556(.A1(new_n756), .A2(G41), .ZN(new_n757));
  INV_X1    g0557(.A(new_n757), .ZN(new_n758));
  NAND2_X1  g0558(.A1(new_n758), .A2(G1), .ZN(new_n759));
  NAND3_X1  g0559(.A1(new_n654), .A2(new_n459), .A3(new_n529), .ZN(new_n760));
  OAI22_X1  g0560(.A1(new_n759), .A2(new_n760), .B1(new_n212), .B2(new_n758), .ZN(new_n761));
  XNOR2_X1  g0561(.A(new_n761), .B(KEYINPUT28), .ZN(new_n762));
  AOI211_X1 g0562(.A(new_n700), .B(new_n699), .C1(new_n593), .C2(new_n547), .ZN(new_n763));
  NAND2_X1  g0563(.A1(new_n619), .A2(new_n624), .ZN(new_n764));
  NAND3_X1  g0564(.A1(new_n764), .A2(new_n648), .A3(new_n649), .ZN(new_n765));
  OAI21_X1  g0565(.A(KEYINPUT26), .B1(new_n765), .B2(new_n700), .ZN(new_n766));
  OAI211_X1 g0566(.A(new_n766), .B(new_n677), .C1(KEYINPUT26), .C2(new_n716), .ZN(new_n767));
  OAI21_X1  g0567(.A(new_n738), .B1(new_n763), .B2(new_n767), .ZN(new_n768));
  NAND2_X1  g0568(.A1(new_n768), .A2(KEYINPUT29), .ZN(new_n769));
  NAND2_X1  g0569(.A1(new_n722), .A2(new_n738), .ZN(new_n770));
  OAI21_X1  g0570(.A(new_n769), .B1(new_n770), .B2(KEYINPUT29), .ZN(new_n771));
  INV_X1    g0571(.A(G330), .ZN(new_n772));
  NOR2_X1   g0572(.A1(new_n493), .A2(new_n499), .ZN(new_n773));
  INV_X1    g0573(.A(new_n773), .ZN(new_n774));
  NOR3_X1   g0574(.A1(new_n591), .A2(new_n675), .A3(new_n774), .ZN(new_n775));
  NOR2_X1   g0575(.A1(new_n645), .A2(new_n641), .ZN(new_n776));
  NOR2_X1   g0576(.A1(KEYINPUT97), .A2(KEYINPUT30), .ZN(new_n777));
  AND3_X1   g0577(.A1(new_n775), .A2(new_n776), .A3(new_n777), .ZN(new_n778));
  INV_X1    g0578(.A(KEYINPUT97), .ZN(new_n779));
  INV_X1    g0579(.A(KEYINPUT30), .ZN(new_n780));
  AOI22_X1  g0580(.A1(new_n775), .A2(new_n776), .B1(new_n779), .B2(new_n780), .ZN(new_n781));
  NOR2_X1   g0581(.A1(new_n590), .A2(G179), .ZN(new_n782));
  NAND3_X1  g0582(.A1(new_n782), .A2(new_n506), .A3(new_n675), .ZN(new_n783));
  OAI22_X1  g0583(.A1(new_n778), .A2(new_n781), .B1(new_n776), .B2(new_n783), .ZN(new_n784));
  OAI21_X1  g0584(.A(new_n745), .B1(new_n784), .B2(KEYINPUT31), .ZN(new_n785));
  INV_X1    g0585(.A(KEYINPUT31), .ZN(new_n786));
  OAI21_X1  g0586(.A(new_n785), .B1(new_n688), .B2(new_n786), .ZN(new_n787));
  NOR2_X1   g0587(.A1(new_n738), .A2(new_n786), .ZN(new_n788));
  NAND2_X1  g0588(.A1(new_n784), .A2(new_n788), .ZN(new_n789));
  INV_X1    g0589(.A(KEYINPUT98), .ZN(new_n790));
  NAND2_X1  g0590(.A1(new_n789), .A2(new_n790), .ZN(new_n791));
  NAND3_X1  g0591(.A1(new_n784), .A2(KEYINPUT98), .A3(new_n788), .ZN(new_n792));
  NAND2_X1  g0592(.A1(new_n791), .A2(new_n792), .ZN(new_n793));
  AOI21_X1  g0593(.A(new_n772), .B1(new_n787), .B2(new_n793), .ZN(new_n794));
  NOR2_X1   g0594(.A1(new_n771), .A2(new_n794), .ZN(new_n795));
  OAI21_X1  g0595(.A(new_n762), .B1(new_n795), .B2(G1), .ZN(G364));
  NAND2_X1  g0596(.A1(new_n733), .A2(G45), .ZN(new_n797));
  NAND3_X1  g0597(.A1(new_n758), .A2(G1), .A3(new_n797), .ZN(new_n798));
  INV_X1    g0598(.A(new_n798), .ZN(new_n799));
  NOR2_X1   g0599(.A1(new_n744), .A2(new_n799), .ZN(new_n800));
  OAI21_X1  g0600(.A(new_n800), .B1(G330), .B2(new_n742), .ZN(new_n801));
  NOR2_X1   g0601(.A1(new_n756), .A2(new_n556), .ZN(new_n802));
  AOI22_X1  g0602(.A1(new_n802), .A2(G355), .B1(new_n529), .B2(new_n756), .ZN(new_n803));
  NOR2_X1   g0603(.A1(new_n353), .A2(new_n756), .ZN(new_n804));
  INV_X1    g0604(.A(new_n804), .ZN(new_n805));
  AOI21_X1  g0605(.A(new_n805), .B1(new_n252), .B2(new_n213), .ZN(new_n806));
  NAND2_X1  g0606(.A1(new_n806), .A2(KEYINPUT99), .ZN(new_n807));
  OAI21_X1  g0607(.A(new_n807), .B1(new_n252), .B2(new_n245), .ZN(new_n808));
  NOR2_X1   g0608(.A1(new_n806), .A2(KEYINPUT99), .ZN(new_n809));
  OAI21_X1  g0609(.A(new_n803), .B1(new_n808), .B2(new_n809), .ZN(new_n810));
  NOR2_X1   g0610(.A1(G13), .A2(G33), .ZN(new_n811));
  INV_X1    g0611(.A(new_n811), .ZN(new_n812));
  NOR2_X1   g0612(.A1(new_n812), .A2(G20), .ZN(new_n813));
  AOI21_X1  g0613(.A(new_n214), .B1(G20), .B2(new_n297), .ZN(new_n814));
  NOR2_X1   g0614(.A1(new_n813), .A2(new_n814), .ZN(new_n815));
  AND2_X1   g0615(.A1(new_n810), .A2(new_n815), .ZN(new_n816));
  NAND2_X1  g0616(.A1(new_n385), .A2(G20), .ZN(new_n817));
  INV_X1    g0617(.A(KEYINPUT101), .ZN(new_n818));
  XNOR2_X1  g0618(.A(new_n817), .B(new_n818), .ZN(new_n819));
  NOR3_X1   g0619(.A1(new_n819), .A2(G179), .A3(new_n369), .ZN(new_n820));
  INV_X1    g0620(.A(new_n820), .ZN(new_n821));
  INV_X1    g0621(.A(G283), .ZN(new_n822));
  INV_X1    g0622(.A(G326), .ZN(new_n823));
  NAND2_X1  g0623(.A1(G20), .A2(G179), .ZN(new_n824));
  XOR2_X1   g0624(.A(new_n824), .B(KEYINPUT100), .Z(new_n825));
  NOR2_X1   g0625(.A1(new_n385), .A2(new_n369), .ZN(new_n826));
  NAND2_X1  g0626(.A1(new_n825), .A2(new_n826), .ZN(new_n827));
  OAI22_X1  g0627(.A1(new_n821), .A2(new_n822), .B1(new_n823), .B2(new_n827), .ZN(new_n828));
  NOR3_X1   g0628(.A1(new_n385), .A2(G179), .A3(G200), .ZN(new_n829));
  NOR2_X1   g0629(.A1(new_n829), .A2(new_n215), .ZN(new_n830));
  INV_X1    g0630(.A(new_n830), .ZN(new_n831));
  AND2_X1   g0631(.A1(new_n831), .A2(new_n490), .ZN(new_n832));
  NOR4_X1   g0632(.A1(new_n215), .A2(new_n385), .A3(new_n369), .A4(G179), .ZN(new_n833));
  INV_X1    g0633(.A(new_n833), .ZN(new_n834));
  INV_X1    g0634(.A(G303), .ZN(new_n835));
  OAI21_X1  g0635(.A(new_n556), .B1(new_n834), .B2(new_n835), .ZN(new_n836));
  NOR3_X1   g0636(.A1(new_n819), .A2(G179), .A3(G200), .ZN(new_n837));
  AOI211_X1 g0637(.A(new_n832), .B(new_n836), .C1(G329), .C2(new_n837), .ZN(new_n838));
  INV_X1    g0638(.A(G311), .ZN(new_n839));
  NAND3_X1  g0639(.A1(new_n825), .A2(new_n385), .A3(new_n369), .ZN(new_n840));
  NAND2_X1  g0640(.A1(new_n825), .A2(new_n385), .ZN(new_n841));
  NOR2_X1   g0641(.A1(new_n841), .A2(new_n369), .ZN(new_n842));
  INV_X1    g0642(.A(new_n842), .ZN(new_n843));
  XOR2_X1   g0643(.A(KEYINPUT33), .B(G317), .Z(new_n844));
  OAI221_X1 g0644(.A(new_n838), .B1(new_n839), .B2(new_n840), .C1(new_n843), .C2(new_n844), .ZN(new_n845));
  NOR2_X1   g0645(.A1(new_n385), .A2(G200), .ZN(new_n846));
  AND2_X1   g0646(.A1(new_n825), .A2(new_n846), .ZN(new_n847));
  AOI211_X1 g0647(.A(new_n828), .B(new_n845), .C1(G322), .C2(new_n847), .ZN(new_n848));
  OR2_X1    g0648(.A1(new_n848), .A2(KEYINPUT103), .ZN(new_n849));
  NAND2_X1  g0649(.A1(new_n848), .A2(KEYINPUT103), .ZN(new_n850));
  INV_X1    g0650(.A(new_n837), .ZN(new_n851));
  XOR2_X1   g0651(.A(KEYINPUT102), .B(G159), .Z(new_n852));
  NOR2_X1   g0652(.A1(new_n851), .A2(new_n852), .ZN(new_n853));
  XNOR2_X1  g0653(.A(new_n853), .B(KEYINPUT32), .ZN(new_n854));
  INV_X1    g0654(.A(new_n847), .ZN(new_n855));
  INV_X1    g0655(.A(new_n337), .ZN(new_n856));
  OAI22_X1  g0656(.A1(new_n855), .A2(new_n856), .B1(new_n202), .B2(new_n827), .ZN(new_n857));
  NOR2_X1   g0657(.A1(new_n821), .A2(new_n459), .ZN(new_n858));
  OAI221_X1 g0658(.A(new_n275), .B1(new_n221), .B2(new_n830), .C1(new_n834), .C2(new_n512), .ZN(new_n859));
  NOR3_X1   g0659(.A1(new_n857), .A2(new_n858), .A3(new_n859), .ZN(new_n860));
  INV_X1    g0660(.A(new_n840), .ZN(new_n861));
  AOI22_X1  g0661(.A1(G68), .A2(new_n842), .B1(new_n861), .B2(new_n225), .ZN(new_n862));
  NAND3_X1  g0662(.A1(new_n854), .A2(new_n860), .A3(new_n862), .ZN(new_n863));
  NAND3_X1  g0663(.A1(new_n849), .A2(new_n850), .A3(new_n863), .ZN(new_n864));
  AOI211_X1 g0664(.A(new_n816), .B(new_n798), .C1(new_n864), .C2(new_n814), .ZN(new_n865));
  INV_X1    g0665(.A(new_n813), .ZN(new_n866));
  OAI21_X1  g0666(.A(new_n865), .B1(new_n742), .B2(new_n866), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n801), .A2(new_n867), .ZN(G396));
  OAI21_X1  g0668(.A(new_n476), .B1(new_n471), .B2(new_n738), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n869), .A2(new_n479), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n727), .A2(new_n738), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n870), .A2(new_n871), .ZN(new_n872));
  INV_X1    g0672(.A(new_n872), .ZN(new_n873));
  XNOR2_X1  g0673(.A(new_n770), .B(new_n873), .ZN(new_n874));
  AOI21_X1  g0674(.A(new_n799), .B1(new_n874), .B2(new_n794), .ZN(new_n875));
  OAI21_X1  g0675(.A(new_n875), .B1(new_n794), .B2(new_n874), .ZN(new_n876));
  INV_X1    g0676(.A(new_n827), .ZN(new_n877));
  AOI22_X1  g0677(.A1(G137), .A2(new_n877), .B1(new_n847), .B2(G143), .ZN(new_n878));
  INV_X1    g0678(.A(G150), .ZN(new_n879));
  OAI221_X1 g0679(.A(new_n878), .B1(new_n840), .B2(new_n852), .C1(new_n879), .C2(new_n843), .ZN(new_n880));
  XOR2_X1   g0680(.A(new_n880), .B(KEYINPUT34), .Z(new_n881));
  OAI221_X1 g0681(.A(new_n353), .B1(new_n856), .B2(new_n830), .C1(new_n834), .C2(new_n202), .ZN(new_n882));
  NOR2_X1   g0682(.A1(new_n821), .A2(new_n357), .ZN(new_n883));
  INV_X1    g0683(.A(new_n883), .ZN(new_n884));
  INV_X1    g0684(.A(G132), .ZN(new_n885));
  OAI21_X1  g0685(.A(new_n884), .B1(new_n885), .B2(new_n851), .ZN(new_n886));
  NOR3_X1   g0686(.A1(new_n881), .A2(new_n882), .A3(new_n886), .ZN(new_n887));
  OAI221_X1 g0687(.A(new_n556), .B1(new_n221), .B2(new_n830), .C1(new_n834), .C2(new_n459), .ZN(new_n888));
  AOI21_X1  g0688(.A(new_n888), .B1(new_n877), .B2(G303), .ZN(new_n889));
  OAI221_X1 g0689(.A(new_n889), .B1(new_n529), .B2(new_n840), .C1(new_n822), .C2(new_n843), .ZN(new_n890));
  NOR2_X1   g0690(.A1(new_n821), .A2(new_n512), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n847), .A2(G294), .ZN(new_n892));
  OAI21_X1  g0692(.A(new_n892), .B1(new_n851), .B2(new_n839), .ZN(new_n893));
  NOR3_X1   g0693(.A1(new_n890), .A2(new_n891), .A3(new_n893), .ZN(new_n894));
  OAI21_X1  g0694(.A(new_n814), .B1(new_n887), .B2(new_n894), .ZN(new_n895));
  NOR2_X1   g0695(.A1(new_n814), .A2(new_n811), .ZN(new_n896));
  AOI21_X1  g0696(.A(new_n798), .B1(new_n319), .B2(new_n896), .ZN(new_n897));
  OAI211_X1 g0697(.A(new_n895), .B(new_n897), .C1(new_n812), .C2(new_n873), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n876), .A2(new_n898), .ZN(G384));
  OAI211_X1 g0699(.A(G116), .B(new_n216), .C1(new_n613), .C2(KEYINPUT35), .ZN(new_n900));
  AOI21_X1  g0700(.A(new_n900), .B1(KEYINPUT35), .B2(new_n613), .ZN(new_n901));
  XNOR2_X1  g0701(.A(new_n901), .B(KEYINPUT36), .ZN(new_n902));
  NAND3_X1  g0702(.A1(new_n213), .A2(new_n338), .A3(new_n225), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n202), .A2(G68), .ZN(new_n904));
  AOI211_X1 g0704(.A(G13), .B(new_n500), .C1(new_n903), .C2(new_n904), .ZN(new_n905));
  NOR2_X1   g0705(.A1(new_n902), .A2(new_n905), .ZN(new_n906));
  AND3_X1   g0706(.A1(new_n398), .A2(KEYINPUT106), .A3(new_n399), .ZN(new_n907));
  AOI21_X1  g0707(.A(KEYINPUT106), .B1(new_n398), .B2(new_n399), .ZN(new_n908));
  OAI21_X1  g0708(.A(new_n726), .B1(new_n907), .B2(new_n908), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n404), .A2(new_n737), .ZN(new_n910));
  INV_X1    g0710(.A(new_n910), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n411), .A2(new_n412), .ZN(new_n912));
  INV_X1    g0712(.A(new_n408), .ZN(new_n913));
  OAI21_X1  g0713(.A(KEYINPUT105), .B1(new_n912), .B2(new_n913), .ZN(new_n914));
  INV_X1    g0714(.A(KEYINPUT37), .ZN(new_n915));
  AND3_X1   g0715(.A1(new_n396), .A2(new_n915), .A3(new_n397), .ZN(new_n916));
  INV_X1    g0716(.A(KEYINPUT105), .ZN(new_n917));
  NAND4_X1  g0717(.A1(new_n411), .A2(new_n917), .A3(new_n408), .A4(new_n412), .ZN(new_n918));
  NAND4_X1  g0718(.A1(new_n914), .A2(new_n916), .A3(new_n918), .A4(new_n910), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n724), .A2(new_n394), .ZN(new_n920));
  OAI21_X1  g0720(.A(KEYINPUT37), .B1(new_n911), .B2(new_n920), .ZN(new_n921));
  AOI22_X1  g0721(.A1(new_n909), .A2(new_n911), .B1(new_n919), .B2(new_n921), .ZN(new_n922));
  NOR2_X1   g0722(.A1(new_n922), .A2(KEYINPUT38), .ZN(new_n923));
  OAI21_X1  g0723(.A(new_n400), .B1(new_n409), .B2(new_n413), .ZN(new_n924));
  OAI21_X1  g0724(.A(new_n340), .B1(new_n351), .B2(new_n354), .ZN(new_n925));
  AND2_X1   g0725(.A1(new_n925), .A2(new_n356), .ZN(new_n926));
  NAND2_X1  g0726(.A1(new_n355), .A2(new_n311), .ZN(new_n927));
  OAI21_X1  g0727(.A(new_n393), .B1(new_n926), .B2(new_n927), .ZN(new_n928));
  AND2_X1   g0728(.A1(new_n928), .A2(new_n737), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n924), .A2(new_n929), .ZN(new_n930));
  OAI21_X1  g0730(.A(new_n928), .B1(new_n408), .B2(new_n737), .ZN(new_n931));
  NAND3_X1  g0731(.A1(new_n931), .A2(new_n396), .A3(new_n397), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n932), .A2(KEYINPUT37), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n919), .A2(new_n933), .ZN(new_n934));
  AND3_X1   g0734(.A1(new_n930), .A2(new_n934), .A3(KEYINPUT38), .ZN(new_n935));
  OAI21_X1  g0735(.A(KEYINPUT40), .B1(new_n923), .B2(new_n935), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n329), .A2(new_n745), .ZN(new_n937));
  NAND3_X1  g0737(.A1(new_n330), .A2(new_n334), .A3(new_n937), .ZN(new_n938));
  OAI211_X1 g0738(.A(new_n329), .B(new_n745), .C1(new_n309), .C2(new_n333), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n938), .A2(new_n939), .ZN(new_n940));
  AOI21_X1  g0740(.A(new_n872), .B1(new_n787), .B2(new_n789), .ZN(new_n941));
  NAND2_X1  g0741(.A1(new_n940), .A2(new_n941), .ZN(new_n942));
  INV_X1    g0742(.A(KEYINPUT108), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n942), .A2(new_n943), .ZN(new_n944));
  NAND3_X1  g0744(.A1(new_n940), .A2(new_n941), .A3(KEYINPUT108), .ZN(new_n945));
  AOI21_X1  g0745(.A(new_n936), .B1(new_n944), .B2(new_n945), .ZN(new_n946));
  XNOR2_X1  g0746(.A(KEYINPUT107), .B(KEYINPUT40), .ZN(new_n947));
  INV_X1    g0747(.A(new_n942), .ZN(new_n948));
  AOI21_X1  g0748(.A(KEYINPUT38), .B1(new_n930), .B2(new_n934), .ZN(new_n949));
  NOR2_X1   g0749(.A1(new_n935), .A2(new_n949), .ZN(new_n950));
  INV_X1    g0750(.A(new_n950), .ZN(new_n951));
  AOI21_X1  g0751(.A(new_n947), .B1(new_n948), .B2(new_n951), .ZN(new_n952));
  NOR2_X1   g0752(.A1(new_n946), .A2(new_n952), .ZN(new_n953));
  NAND2_X1  g0753(.A1(new_n787), .A2(new_n789), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n485), .A2(new_n954), .ZN(new_n955));
  XOR2_X1   g0755(.A(new_n953), .B(new_n955), .Z(new_n956));
  NOR2_X1   g0756(.A1(new_n956), .A2(new_n772), .ZN(new_n957));
  NAND3_X1  g0757(.A1(new_n722), .A2(new_n738), .A3(new_n873), .ZN(new_n958));
  NAND2_X1  g0758(.A1(new_n958), .A2(new_n871), .ZN(new_n959));
  NAND2_X1  g0759(.A1(new_n959), .A2(new_n940), .ZN(new_n960));
  NAND2_X1  g0760(.A1(new_n960), .A2(KEYINPUT104), .ZN(new_n961));
  AOI22_X1  g0761(.A1(new_n958), .A2(new_n871), .B1(new_n938), .B2(new_n939), .ZN(new_n962));
  INV_X1    g0762(.A(KEYINPUT104), .ZN(new_n963));
  NAND2_X1  g0763(.A1(new_n962), .A2(new_n963), .ZN(new_n964));
  AOI21_X1  g0764(.A(new_n950), .B1(new_n961), .B2(new_n964), .ZN(new_n965));
  OAI21_X1  g0765(.A(KEYINPUT39), .B1(new_n935), .B2(new_n949), .ZN(new_n966));
  INV_X1    g0766(.A(KEYINPUT39), .ZN(new_n967));
  NAND3_X1  g0767(.A1(new_n930), .A2(new_n934), .A3(KEYINPUT38), .ZN(new_n968));
  OAI211_X1 g0768(.A(new_n967), .B(new_n968), .C1(new_n922), .C2(KEYINPUT38), .ZN(new_n969));
  NAND2_X1  g0769(.A1(new_n966), .A2(new_n969), .ZN(new_n970));
  NOR2_X1   g0770(.A1(new_n330), .A2(new_n745), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n970), .A2(new_n971), .ZN(new_n972));
  INV_X1    g0772(.A(new_n726), .ZN(new_n973));
  INV_X1    g0773(.A(new_n737), .ZN(new_n974));
  NAND2_X1  g0774(.A1(new_n973), .A2(new_n974), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n972), .A2(new_n975), .ZN(new_n976));
  NOR2_X1   g0776(.A1(new_n965), .A2(new_n976), .ZN(new_n977));
  NAND2_X1  g0777(.A1(new_n485), .A2(new_n771), .ZN(new_n978));
  NAND2_X1  g0778(.A1(new_n978), .A2(new_n731), .ZN(new_n979));
  XNOR2_X1  g0779(.A(new_n977), .B(new_n979), .ZN(new_n980));
  OAI22_X1  g0780(.A1(new_n957), .A2(new_n980), .B1(new_n500), .B2(new_n733), .ZN(new_n981));
  AND2_X1   g0781(.A1(new_n957), .A2(new_n980), .ZN(new_n982));
  OAI21_X1  g0782(.A(new_n906), .B1(new_n981), .B2(new_n982), .ZN(G367));
  NAND2_X1  g0783(.A1(new_n764), .A2(new_n745), .ZN(new_n984));
  NAND2_X1  g0784(.A1(new_n690), .A2(new_n984), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n712), .A2(new_n745), .ZN(new_n986));
  NAND2_X1  g0786(.A1(new_n985), .A2(new_n986), .ZN(new_n987));
  NAND2_X1  g0787(.A1(new_n753), .A2(new_n987), .ZN(new_n988));
  XOR2_X1   g0788(.A(new_n988), .B(KEYINPUT42), .Z(new_n989));
  INV_X1    g0789(.A(new_n987), .ZN(new_n990));
  OAI21_X1  g0790(.A(new_n651), .B1(new_n990), .B2(new_n547), .ZN(new_n991));
  NAND2_X1  g0791(.A1(new_n991), .A2(new_n738), .ZN(new_n992));
  NAND2_X1  g0792(.A1(new_n989), .A2(new_n992), .ZN(new_n993));
  INV_X1    g0793(.A(KEYINPUT109), .ZN(new_n994));
  NAND2_X1  g0794(.A1(new_n993), .A2(new_n994), .ZN(new_n995));
  NAND3_X1  g0795(.A1(new_n989), .A2(KEYINPUT109), .A3(new_n992), .ZN(new_n996));
  NOR2_X1   g0796(.A1(new_n693), .A2(new_n695), .ZN(new_n997));
  NAND2_X1  g0797(.A1(new_n997), .A2(new_n745), .ZN(new_n998));
  NAND2_X1  g0798(.A1(new_n700), .A2(new_n998), .ZN(new_n999));
  NAND3_X1  g0799(.A1(new_n677), .A2(new_n997), .A3(new_n745), .ZN(new_n1000));
  NAND2_X1  g0800(.A1(new_n999), .A2(new_n1000), .ZN(new_n1001));
  XNOR2_X1  g0801(.A(new_n1001), .B(KEYINPUT43), .ZN(new_n1002));
  NAND3_X1  g0802(.A1(new_n995), .A2(new_n996), .A3(new_n1002), .ZN(new_n1003));
  INV_X1    g0803(.A(new_n1003), .ZN(new_n1004));
  INV_X1    g0804(.A(new_n1001), .ZN(new_n1005));
  NOR2_X1   g0805(.A1(new_n1005), .A2(KEYINPUT43), .ZN(new_n1006));
  INV_X1    g0806(.A(new_n1006), .ZN(new_n1007));
  AOI21_X1  g0807(.A(new_n1007), .B1(new_n995), .B2(new_n996), .ZN(new_n1008));
  OAI22_X1  g0808(.A1(new_n1004), .A2(new_n1008), .B1(new_n751), .B2(new_n990), .ZN(new_n1009));
  INV_X1    g0809(.A(new_n1008), .ZN(new_n1010));
  NOR2_X1   g0810(.A1(new_n751), .A2(new_n990), .ZN(new_n1011));
  NAND3_X1  g0811(.A1(new_n1010), .A2(new_n1003), .A3(new_n1011), .ZN(new_n1012));
  NAND2_X1  g0812(.A1(new_n1009), .A2(new_n1012), .ZN(new_n1013));
  INV_X1    g0813(.A(new_n1013), .ZN(new_n1014));
  XOR2_X1   g0814(.A(new_n757), .B(KEYINPUT41), .Z(new_n1015));
  INV_X1    g0815(.A(new_n754), .ZN(new_n1016));
  OAI21_X1  g0816(.A(KEYINPUT110), .B1(new_n1016), .B2(new_n990), .ZN(new_n1017));
  INV_X1    g0817(.A(KEYINPUT110), .ZN(new_n1018));
  NAND3_X1  g0818(.A1(new_n754), .A2(new_n1018), .A3(new_n987), .ZN(new_n1019));
  NAND2_X1  g0819(.A1(new_n1017), .A2(new_n1019), .ZN(new_n1020));
  INV_X1    g0820(.A(KEYINPUT45), .ZN(new_n1021));
  NAND2_X1  g0821(.A1(new_n1020), .A2(new_n1021), .ZN(new_n1022));
  NOR2_X1   g0822(.A1(new_n754), .A2(new_n987), .ZN(new_n1023));
  XNOR2_X1  g0823(.A(new_n1023), .B(KEYINPUT44), .ZN(new_n1024));
  NAND3_X1  g0824(.A1(new_n1017), .A2(KEYINPUT45), .A3(new_n1019), .ZN(new_n1025));
  INV_X1    g0825(.A(KEYINPUT112), .ZN(new_n1026));
  NAND3_X1  g0826(.A1(new_n744), .A2(new_n1026), .A3(new_n750), .ZN(new_n1027));
  NAND4_X1  g0827(.A1(new_n1022), .A2(new_n1024), .A3(new_n1025), .A4(new_n1027), .ZN(new_n1028));
  NAND2_X1  g0828(.A1(new_n751), .A2(KEYINPUT112), .ZN(new_n1029));
  INV_X1    g0829(.A(new_n1029), .ZN(new_n1030));
  NAND2_X1  g0830(.A1(new_n1028), .A2(new_n1030), .ZN(new_n1031));
  AND2_X1   g0831(.A1(new_n1025), .A2(new_n1027), .ZN(new_n1032));
  NAND4_X1  g0832(.A1(new_n1032), .A2(new_n1022), .A3(new_n1024), .A4(new_n1029), .ZN(new_n1033));
  NAND2_X1  g0833(.A1(new_n1031), .A2(new_n1033), .ZN(new_n1034));
  XNOR2_X1  g0834(.A(new_n750), .B(new_n752), .ZN(new_n1035));
  INV_X1    g0835(.A(KEYINPUT111), .ZN(new_n1036));
  AOI21_X1  g0836(.A(new_n1035), .B1(new_n743), .B2(new_n1036), .ZN(new_n1037));
  NOR2_X1   g0837(.A1(new_n743), .A2(new_n1036), .ZN(new_n1038));
  XNOR2_X1  g0838(.A(new_n1037), .B(new_n1038), .ZN(new_n1039));
  INV_X1    g0839(.A(new_n795), .ZN(new_n1040));
  NOR2_X1   g0840(.A1(new_n1039), .A2(new_n1040), .ZN(new_n1041));
  NAND2_X1  g0841(.A1(new_n1034), .A2(new_n1041), .ZN(new_n1042));
  AOI21_X1  g0842(.A(new_n1015), .B1(new_n1042), .B2(new_n795), .ZN(new_n1043));
  NAND2_X1  g0843(.A1(new_n797), .A2(G1), .ZN(new_n1044));
  OAI21_X1  g0844(.A(new_n1014), .B1(new_n1043), .B2(new_n1044), .ZN(new_n1045));
  INV_X1    g0845(.A(new_n815), .ZN(new_n1046));
  AOI21_X1  g0846(.A(new_n1046), .B1(new_n756), .B2(new_n467), .ZN(new_n1047));
  NAND2_X1  g0847(.A1(new_n804), .A2(new_n241), .ZN(new_n1048));
  AOI21_X1  g0848(.A(new_n798), .B1(new_n1047), .B2(new_n1048), .ZN(new_n1049));
  AOI22_X1  g0849(.A1(G143), .A2(new_n877), .B1(new_n820), .B2(new_n225), .ZN(new_n1050));
  INV_X1    g0850(.A(G137), .ZN(new_n1051));
  OAI21_X1  g0851(.A(new_n1050), .B1(new_n1051), .B2(new_n851), .ZN(new_n1052));
  AOI21_X1  g0852(.A(new_n556), .B1(new_n833), .B2(new_n337), .ZN(new_n1053));
  OAI221_X1 g0853(.A(new_n1053), .B1(new_n357), .B2(new_n830), .C1(new_n855), .C2(new_n879), .ZN(new_n1054));
  NOR2_X1   g0854(.A1(new_n843), .A2(new_n852), .ZN(new_n1055));
  NOR2_X1   g0855(.A1(new_n840), .A2(new_n202), .ZN(new_n1056));
  NOR4_X1   g0856(.A1(new_n1052), .A2(new_n1054), .A3(new_n1055), .A4(new_n1056), .ZN(new_n1057));
  XNOR2_X1  g0857(.A(new_n1057), .B(KEYINPUT113), .ZN(new_n1058));
  AOI22_X1  g0858(.A1(new_n837), .A2(G317), .B1(new_n847), .B2(G303), .ZN(new_n1059));
  NAND2_X1  g0859(.A1(new_n820), .A2(G97), .ZN(new_n1060));
  OAI211_X1 g0860(.A(new_n1059), .B(new_n1060), .C1(new_n839), .C2(new_n827), .ZN(new_n1061));
  NOR2_X1   g0861(.A1(new_n840), .A2(new_n822), .ZN(new_n1062));
  NOR2_X1   g0862(.A1(new_n834), .A2(new_n529), .ZN(new_n1063));
  OR2_X1    g0863(.A1(new_n1063), .A2(KEYINPUT46), .ZN(new_n1064));
  AOI22_X1  g0864(.A1(new_n1063), .A2(KEYINPUT46), .B1(G107), .B2(new_n831), .ZN(new_n1065));
  INV_X1    g0865(.A(new_n353), .ZN(new_n1066));
  NAND3_X1  g0866(.A1(new_n1064), .A2(new_n1065), .A3(new_n1066), .ZN(new_n1067));
  AND2_X1   g0867(.A1(new_n842), .A2(new_n490), .ZN(new_n1068));
  OR4_X1    g0868(.A1(new_n1061), .A2(new_n1062), .A3(new_n1067), .A4(new_n1068), .ZN(new_n1069));
  NAND3_X1  g0869(.A1(new_n1058), .A2(KEYINPUT47), .A3(new_n1069), .ZN(new_n1070));
  NAND2_X1  g0870(.A1(new_n1070), .A2(new_n814), .ZN(new_n1071));
  AOI21_X1  g0871(.A(KEYINPUT47), .B1(new_n1058), .B2(new_n1069), .ZN(new_n1072));
  OAI221_X1 g0872(.A(new_n1049), .B1(new_n866), .B2(new_n1005), .C1(new_n1071), .C2(new_n1072), .ZN(new_n1073));
  NAND2_X1  g0873(.A1(new_n1045), .A2(new_n1073), .ZN(G387));
  NAND2_X1  g0874(.A1(new_n802), .A2(new_n760), .ZN(new_n1075));
  OAI21_X1  g0875(.A(new_n1075), .B1(G107), .B2(new_n208), .ZN(new_n1076));
  NAND2_X1  g0876(.A1(new_n237), .A2(G45), .ZN(new_n1077));
  NAND2_X1  g0877(.A1(new_n464), .A2(new_n202), .ZN(new_n1078));
  XOR2_X1   g0878(.A(new_n1078), .B(KEYINPUT50), .Z(new_n1079));
  AOI211_X1 g0879(.A(G45), .B(new_n760), .C1(G68), .C2(G77), .ZN(new_n1080));
  AOI21_X1  g0880(.A(new_n805), .B1(new_n1079), .B2(new_n1080), .ZN(new_n1081));
  AOI21_X1  g0881(.A(new_n1076), .B1(new_n1077), .B2(new_n1081), .ZN(new_n1082));
  OAI21_X1  g0882(.A(new_n799), .B1(new_n1082), .B2(new_n1046), .ZN(new_n1083));
  AOI21_X1  g0883(.A(new_n353), .B1(new_n820), .B2(G116), .ZN(new_n1084));
  AOI22_X1  g0884(.A1(G322), .A2(new_n877), .B1(new_n847), .B2(G317), .ZN(new_n1085));
  OAI21_X1  g0885(.A(new_n1085), .B1(new_n835), .B2(new_n840), .ZN(new_n1086));
  AOI21_X1  g0886(.A(new_n1086), .B1(G311), .B2(new_n842), .ZN(new_n1087));
  OR2_X1    g0887(.A1(new_n1087), .A2(KEYINPUT48), .ZN(new_n1088));
  NAND2_X1  g0888(.A1(new_n1087), .A2(KEYINPUT48), .ZN(new_n1089));
  AOI22_X1  g0889(.A1(new_n831), .A2(G283), .B1(new_n490), .B2(new_n833), .ZN(new_n1090));
  NAND3_X1  g0890(.A1(new_n1088), .A2(new_n1089), .A3(new_n1090), .ZN(new_n1091));
  INV_X1    g0891(.A(KEYINPUT49), .ZN(new_n1092));
  OAI221_X1 g0892(.A(new_n1084), .B1(new_n823), .B2(new_n851), .C1(new_n1091), .C2(new_n1092), .ZN(new_n1093));
  AND2_X1   g0893(.A1(new_n1091), .A2(new_n1092), .ZN(new_n1094));
  AOI22_X1  g0894(.A1(new_n837), .A2(G150), .B1(new_n847), .B2(G50), .ZN(new_n1095));
  OAI211_X1 g0895(.A(new_n1095), .B(new_n1060), .C1(new_n365), .C2(new_n827), .ZN(new_n1096));
  NAND2_X1  g0896(.A1(new_n831), .A2(new_n467), .ZN(new_n1097));
  OAI211_X1 g0897(.A(new_n1097), .B(new_n353), .C1(new_n416), .C2(new_n834), .ZN(new_n1098));
  AOI21_X1  g0898(.A(new_n1098), .B1(new_n842), .B2(new_n389), .ZN(new_n1099));
  OAI21_X1  g0899(.A(new_n1099), .B1(new_n357), .B2(new_n840), .ZN(new_n1100));
  OAI22_X1  g0900(.A1(new_n1093), .A2(new_n1094), .B1(new_n1096), .B2(new_n1100), .ZN(new_n1101));
  AOI21_X1  g0901(.A(new_n1083), .B1(new_n1101), .B2(new_n814), .ZN(new_n1102));
  OAI21_X1  g0902(.A(new_n1102), .B1(new_n750), .B2(new_n866), .ZN(new_n1103));
  XNOR2_X1  g0903(.A(new_n1103), .B(KEYINPUT114), .ZN(new_n1104));
  INV_X1    g0904(.A(new_n1044), .ZN(new_n1105));
  OAI21_X1  g0905(.A(new_n1104), .B1(new_n1039), .B2(new_n1105), .ZN(new_n1106));
  INV_X1    g0906(.A(new_n1106), .ZN(new_n1107));
  INV_X1    g0907(.A(new_n1041), .ZN(new_n1108));
  XNOR2_X1  g0908(.A(new_n757), .B(KEYINPUT115), .ZN(new_n1109));
  NAND3_X1  g0909(.A1(new_n1108), .A2(KEYINPUT116), .A3(new_n1109), .ZN(new_n1110));
  NAND2_X1  g0910(.A1(new_n1039), .A2(new_n1040), .ZN(new_n1111));
  NAND2_X1  g0911(.A1(new_n1110), .A2(new_n1111), .ZN(new_n1112));
  INV_X1    g0912(.A(KEYINPUT116), .ZN(new_n1113));
  INV_X1    g0913(.A(new_n1109), .ZN(new_n1114));
  OAI21_X1  g0914(.A(new_n1113), .B1(new_n1041), .B2(new_n1114), .ZN(new_n1115));
  INV_X1    g0915(.A(new_n1115), .ZN(new_n1116));
  OAI21_X1  g0916(.A(new_n1107), .B1(new_n1112), .B2(new_n1116), .ZN(G393));
  NAND3_X1  g0917(.A1(new_n1031), .A2(new_n1108), .A3(new_n1033), .ZN(new_n1118));
  NAND3_X1  g0918(.A1(new_n1042), .A2(new_n1109), .A3(new_n1118), .ZN(new_n1119));
  NAND2_X1  g0919(.A1(new_n990), .A2(new_n813), .ZN(new_n1120));
  OAI221_X1 g0920(.A(new_n815), .B1(new_n221), .B2(new_n208), .C1(new_n805), .C2(new_n248), .ZN(new_n1121));
  NAND2_X1  g0921(.A1(new_n1121), .A2(new_n799), .ZN(new_n1122));
  AOI22_X1  g0922(.A1(G317), .A2(new_n877), .B1(new_n847), .B2(G311), .ZN(new_n1123));
  XOR2_X1   g0923(.A(new_n1123), .B(KEYINPUT52), .Z(new_n1124));
  OAI221_X1 g0924(.A(new_n556), .B1(new_n529), .B2(new_n830), .C1(new_n834), .C2(new_n822), .ZN(new_n1125));
  AOI211_X1 g0925(.A(new_n1125), .B(new_n858), .C1(G322), .C2(new_n837), .ZN(new_n1126));
  AOI22_X1  g0926(.A1(G303), .A2(new_n842), .B1(new_n861), .B2(G294), .ZN(new_n1127));
  NAND3_X1  g0927(.A1(new_n1124), .A2(new_n1126), .A3(new_n1127), .ZN(new_n1128));
  NAND2_X1  g0928(.A1(new_n861), .A2(new_n464), .ZN(new_n1129));
  OAI221_X1 g0929(.A(new_n1129), .B1(new_n319), .B2(new_n830), .C1(new_n843), .C2(new_n202), .ZN(new_n1130));
  XOR2_X1   g0930(.A(new_n1130), .B(KEYINPUT117), .Z(new_n1131));
  AOI211_X1 g0931(.A(new_n1066), .B(new_n891), .C1(G68), .C2(new_n833), .ZN(new_n1132));
  OAI22_X1  g0932(.A1(new_n855), .A2(new_n365), .B1(new_n879), .B2(new_n827), .ZN(new_n1133));
  XNOR2_X1  g0933(.A(new_n1133), .B(KEYINPUT51), .ZN(new_n1134));
  NAND2_X1  g0934(.A1(new_n837), .A2(G143), .ZN(new_n1135));
  NAND3_X1  g0935(.A1(new_n1132), .A2(new_n1134), .A3(new_n1135), .ZN(new_n1136));
  OAI21_X1  g0936(.A(new_n1128), .B1(new_n1131), .B2(new_n1136), .ZN(new_n1137));
  AOI21_X1  g0937(.A(new_n1122), .B1(new_n1137), .B2(new_n814), .ZN(new_n1138));
  AOI22_X1  g0938(.A1(new_n1034), .A2(new_n1044), .B1(new_n1120), .B2(new_n1138), .ZN(new_n1139));
  NAND2_X1  g0939(.A1(new_n1119), .A2(new_n1139), .ZN(G390));
  INV_X1    g0940(.A(new_n870), .ZN(new_n1141));
  OAI21_X1  g0941(.A(new_n871), .B1(new_n768), .B2(new_n1141), .ZN(new_n1142));
  INV_X1    g0942(.A(KEYINPUT118), .ZN(new_n1143));
  AND3_X1   g0943(.A1(new_n938), .A2(new_n1143), .A3(new_n939), .ZN(new_n1144));
  AOI21_X1  g0944(.A(new_n1143), .B1(new_n938), .B2(new_n939), .ZN(new_n1145));
  OAI21_X1  g0945(.A(new_n1142), .B1(new_n1144), .B2(new_n1145), .ZN(new_n1146));
  INV_X1    g0946(.A(KEYINPUT38), .ZN(new_n1147));
  AND2_X1   g0947(.A1(new_n909), .A2(new_n911), .ZN(new_n1148));
  AND2_X1   g0948(.A1(new_n921), .A2(new_n919), .ZN(new_n1149));
  OAI21_X1  g0949(.A(new_n1147), .B1(new_n1148), .B2(new_n1149), .ZN(new_n1150));
  AOI21_X1  g0950(.A(new_n971), .B1(new_n1150), .B2(new_n968), .ZN(new_n1151));
  NAND2_X1  g0951(.A1(new_n1146), .A2(new_n1151), .ZN(new_n1152));
  OAI211_X1 g0952(.A(new_n966), .B(new_n969), .C1(new_n962), .C2(new_n971), .ZN(new_n1153));
  AOI211_X1 g0953(.A(new_n772), .B(new_n872), .C1(new_n787), .C2(new_n793), .ZN(new_n1154));
  NAND2_X1  g0954(.A1(new_n1154), .A2(new_n940), .ZN(new_n1155));
  NAND3_X1  g0955(.A1(new_n1152), .A2(new_n1153), .A3(new_n1155), .ZN(new_n1156));
  INV_X1    g0956(.A(new_n971), .ZN(new_n1157));
  NAND2_X1  g0957(.A1(new_n960), .A2(new_n1157), .ZN(new_n1158));
  AND2_X1   g0958(.A1(new_n966), .A2(new_n969), .ZN(new_n1159));
  AOI22_X1  g0959(.A1(new_n1158), .A2(new_n1159), .B1(new_n1146), .B2(new_n1151), .ZN(new_n1160));
  NAND3_X1  g0960(.A1(new_n940), .A2(new_n941), .A3(G330), .ZN(new_n1161));
  OAI21_X1  g0961(.A(new_n1156), .B1(new_n1160), .B2(new_n1161), .ZN(new_n1162));
  INV_X1    g0962(.A(new_n1162), .ZN(new_n1163));
  OAI21_X1  g0963(.A(new_n1161), .B1(new_n1154), .B2(new_n940), .ZN(new_n1164));
  NAND2_X1  g0964(.A1(new_n1164), .A2(new_n959), .ZN(new_n1165));
  NAND2_X1  g0965(.A1(new_n940), .A2(KEYINPUT118), .ZN(new_n1166));
  NAND2_X1  g0966(.A1(new_n941), .A2(G330), .ZN(new_n1167));
  NAND3_X1  g0967(.A1(new_n938), .A2(new_n1143), .A3(new_n939), .ZN(new_n1168));
  NAND3_X1  g0968(.A1(new_n1166), .A2(new_n1167), .A3(new_n1168), .ZN(new_n1169));
  AOI21_X1  g0969(.A(new_n1142), .B1(new_n1154), .B2(new_n940), .ZN(new_n1170));
  NAND2_X1  g0970(.A1(new_n1169), .A2(new_n1170), .ZN(new_n1171));
  NAND2_X1  g0971(.A1(new_n1165), .A2(new_n1171), .ZN(new_n1172));
  NAND2_X1  g0972(.A1(new_n330), .A2(new_n334), .ZN(new_n1173));
  AOI21_X1  g0973(.A(new_n484), .B1(new_n1173), .B2(KEYINPUT77), .ZN(new_n1174));
  INV_X1    g0974(.A(new_n336), .ZN(new_n1175));
  NAND4_X1  g0975(.A1(new_n1174), .A2(G330), .A3(new_n1175), .A4(new_n954), .ZN(new_n1176));
  NAND3_X1  g0976(.A1(new_n978), .A2(new_n731), .A3(new_n1176), .ZN(new_n1177));
  NAND2_X1  g0977(.A1(new_n1177), .A2(KEYINPUT119), .ZN(new_n1178));
  INV_X1    g0978(.A(KEYINPUT119), .ZN(new_n1179));
  NAND4_X1  g0979(.A1(new_n978), .A2(new_n1176), .A3(new_n1179), .A4(new_n731), .ZN(new_n1180));
  NAND3_X1  g0980(.A1(new_n1172), .A2(new_n1178), .A3(new_n1180), .ZN(new_n1181));
  INV_X1    g0981(.A(new_n1181), .ZN(new_n1182));
  AOI21_X1  g0982(.A(new_n1114), .B1(new_n1163), .B2(new_n1182), .ZN(new_n1183));
  OAI21_X1  g0983(.A(new_n1183), .B1(new_n1163), .B2(new_n1182), .ZN(new_n1184));
  NAND2_X1  g0984(.A1(new_n1159), .A2(new_n811), .ZN(new_n1185));
  INV_X1    g0985(.A(new_n896), .ZN(new_n1186));
  OAI21_X1  g0986(.A(new_n799), .B1(new_n389), .B2(new_n1186), .ZN(new_n1187));
  OAI21_X1  g0987(.A(new_n556), .B1(new_n834), .B2(new_n512), .ZN(new_n1188));
  AOI211_X1 g0988(.A(new_n1188), .B(new_n883), .C1(G77), .C2(new_n831), .ZN(new_n1189));
  OAI221_X1 g0989(.A(new_n1189), .B1(new_n221), .B2(new_n840), .C1(new_n459), .C2(new_n843), .ZN(new_n1190));
  AOI22_X1  g0990(.A1(new_n837), .A2(G294), .B1(new_n847), .B2(G116), .ZN(new_n1191));
  OAI21_X1  g0991(.A(new_n1191), .B1(new_n822), .B2(new_n827), .ZN(new_n1192));
  AOI22_X1  g0992(.A1(G50), .A2(new_n820), .B1(new_n837), .B2(G125), .ZN(new_n1193));
  NAND2_X1  g0993(.A1(new_n833), .A2(G150), .ZN(new_n1194));
  XOR2_X1   g0994(.A(new_n1194), .B(KEYINPUT53), .Z(new_n1195));
  OAI211_X1 g0995(.A(new_n1193), .B(new_n1195), .C1(new_n885), .C2(new_n855), .ZN(new_n1196));
  NAND2_X1  g0996(.A1(new_n842), .A2(G137), .ZN(new_n1197));
  XNOR2_X1  g0997(.A(KEYINPUT54), .B(G143), .ZN(new_n1198));
  XNOR2_X1  g0998(.A(new_n1198), .B(KEYINPUT120), .ZN(new_n1199));
  NAND2_X1  g0999(.A1(new_n861), .A2(new_n1199), .ZN(new_n1200));
  NAND2_X1  g1000(.A1(new_n877), .A2(G128), .ZN(new_n1201));
  AOI21_X1  g1001(.A(new_n556), .B1(new_n831), .B2(G159), .ZN(new_n1202));
  NAND4_X1  g1002(.A1(new_n1197), .A2(new_n1200), .A3(new_n1201), .A4(new_n1202), .ZN(new_n1203));
  OAI22_X1  g1003(.A1(new_n1190), .A2(new_n1192), .B1(new_n1196), .B2(new_n1203), .ZN(new_n1204));
  AOI21_X1  g1004(.A(new_n1187), .B1(new_n1204), .B2(new_n814), .ZN(new_n1205));
  AOI22_X1  g1005(.A1(new_n1163), .A2(new_n1044), .B1(new_n1185), .B2(new_n1205), .ZN(new_n1206));
  NAND2_X1  g1006(.A1(new_n1184), .A2(new_n1206), .ZN(G378));
  AOI221_X4 g1007(.A(KEYINPUT104), .B1(new_n938), .B2(new_n939), .C1(new_n958), .C2(new_n871), .ZN(new_n1208));
  AOI21_X1  g1008(.A(new_n963), .B1(new_n959), .B2(new_n940), .ZN(new_n1209));
  OAI21_X1  g1009(.A(new_n951), .B1(new_n1208), .B2(new_n1209), .ZN(new_n1210));
  AOI22_X1  g1010(.A1(new_n970), .A2(new_n971), .B1(new_n973), .B2(new_n974), .ZN(new_n1211));
  NOR2_X1   g1011(.A1(new_n974), .A2(new_n450), .ZN(new_n1212));
  XNOR2_X1  g1012(.A(new_n482), .B(new_n1212), .ZN(new_n1213));
  XOR2_X1   g1013(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1214));
  XNOR2_X1  g1014(.A(new_n1213), .B(new_n1214), .ZN(new_n1215));
  AND3_X1   g1015(.A1(new_n1210), .A2(new_n1211), .A3(new_n1215), .ZN(new_n1216));
  AOI21_X1  g1016(.A(new_n1215), .B1(new_n1210), .B2(new_n1211), .ZN(new_n1217));
  NOR3_X1   g1017(.A1(new_n946), .A2(new_n952), .A3(new_n772), .ZN(new_n1218));
  NOR3_X1   g1018(.A1(new_n1216), .A2(new_n1217), .A3(new_n1218), .ZN(new_n1219));
  NAND2_X1  g1019(.A1(new_n944), .A2(new_n945), .ZN(new_n1220));
  NAND2_X1  g1020(.A1(new_n1150), .A2(new_n968), .ZN(new_n1221));
  NAND3_X1  g1021(.A1(new_n1220), .A2(KEYINPUT40), .A3(new_n1221), .ZN(new_n1222));
  INV_X1    g1022(.A(new_n952), .ZN(new_n1223));
  NAND3_X1  g1023(.A1(new_n1222), .A2(G330), .A3(new_n1223), .ZN(new_n1224));
  INV_X1    g1024(.A(new_n1215), .ZN(new_n1225));
  OAI21_X1  g1025(.A(new_n1225), .B1(new_n965), .B2(new_n976), .ZN(new_n1226));
  NAND3_X1  g1026(.A1(new_n1210), .A2(new_n1211), .A3(new_n1215), .ZN(new_n1227));
  AOI21_X1  g1027(.A(new_n1224), .B1(new_n1226), .B2(new_n1227), .ZN(new_n1228));
  OAI21_X1  g1028(.A(KEYINPUT121), .B1(new_n1219), .B2(new_n1228), .ZN(new_n1229));
  OAI21_X1  g1029(.A(new_n1218), .B1(new_n1216), .B2(new_n1217), .ZN(new_n1230));
  INV_X1    g1030(.A(KEYINPUT121), .ZN(new_n1231));
  NAND3_X1  g1031(.A1(new_n1226), .A2(new_n1224), .A3(new_n1227), .ZN(new_n1232));
  NAND3_X1  g1032(.A1(new_n1230), .A2(new_n1231), .A3(new_n1232), .ZN(new_n1233));
  AND2_X1   g1033(.A1(new_n1178), .A2(new_n1180), .ZN(new_n1234));
  AND2_X1   g1034(.A1(new_n1165), .A2(new_n1171), .ZN(new_n1235));
  OAI21_X1  g1035(.A(new_n1234), .B1(new_n1162), .B2(new_n1235), .ZN(new_n1236));
  NAND3_X1  g1036(.A1(new_n1229), .A2(new_n1233), .A3(new_n1236), .ZN(new_n1237));
  INV_X1    g1037(.A(KEYINPUT57), .ZN(new_n1238));
  NAND2_X1  g1038(.A1(new_n1237), .A2(new_n1238), .ZN(new_n1239));
  NOR2_X1   g1039(.A1(new_n1219), .A2(new_n1228), .ZN(new_n1240));
  NAND2_X1  g1040(.A1(new_n1236), .A2(KEYINPUT57), .ZN(new_n1241));
  OAI21_X1  g1041(.A(new_n1109), .B1(new_n1240), .B2(new_n1241), .ZN(new_n1242));
  INV_X1    g1042(.A(new_n1242), .ZN(new_n1243));
  NAND2_X1  g1043(.A1(new_n1239), .A2(new_n1243), .ZN(new_n1244));
  NAND3_X1  g1044(.A1(new_n1229), .A2(new_n1233), .A3(new_n1044), .ZN(new_n1245));
  NAND2_X1  g1045(.A1(new_n1215), .A2(new_n811), .ZN(new_n1246));
  OAI21_X1  g1046(.A(new_n799), .B1(G50), .B2(new_n1186), .ZN(new_n1247));
  NAND2_X1  g1047(.A1(new_n877), .A2(G116), .ZN(new_n1248));
  NAND2_X1  g1048(.A1(new_n820), .A2(new_n337), .ZN(new_n1249));
  AND2_X1   g1049(.A1(new_n1248), .A2(new_n1249), .ZN(new_n1250));
  OAI221_X1 g1050(.A(new_n1250), .B1(new_n459), .B2(new_n855), .C1(new_n822), .C2(new_n851), .ZN(new_n1251));
  OAI22_X1  g1051(.A1(new_n834), .A2(new_n416), .B1(new_n357), .B2(new_n830), .ZN(new_n1252));
  NOR2_X1   g1052(.A1(new_n353), .A2(G41), .ZN(new_n1253));
  INV_X1    g1053(.A(new_n1253), .ZN(new_n1254));
  AOI211_X1 g1054(.A(new_n1252), .B(new_n1254), .C1(new_n467), .C2(new_n861), .ZN(new_n1255));
  OAI21_X1  g1055(.A(new_n1255), .B1(new_n221), .B2(new_n843), .ZN(new_n1256));
  NOR2_X1   g1056(.A1(new_n1251), .A2(new_n1256), .ZN(new_n1257));
  OR2_X1    g1057(.A1(new_n1257), .A2(KEYINPUT58), .ZN(new_n1258));
  AOI22_X1  g1058(.A1(G132), .A2(new_n842), .B1(new_n861), .B2(G137), .ZN(new_n1259));
  AOI22_X1  g1059(.A1(new_n847), .A2(G128), .B1(G150), .B2(new_n831), .ZN(new_n1260));
  AOI22_X1  g1060(.A1(new_n877), .A2(G125), .B1(new_n833), .B2(new_n1199), .ZN(new_n1261));
  NAND3_X1  g1061(.A1(new_n1259), .A2(new_n1260), .A3(new_n1261), .ZN(new_n1262));
  OR2_X1    g1062(.A1(new_n1262), .A2(KEYINPUT59), .ZN(new_n1263));
  NAND2_X1  g1063(.A1(new_n1262), .A2(KEYINPUT59), .ZN(new_n1264));
  OAI211_X1 g1064(.A(new_n269), .B(new_n251), .C1(new_n821), .C2(new_n852), .ZN(new_n1265));
  AOI21_X1  g1065(.A(new_n1265), .B1(G124), .B2(new_n837), .ZN(new_n1266));
  NAND3_X1  g1066(.A1(new_n1263), .A2(new_n1264), .A3(new_n1266), .ZN(new_n1267));
  NAND2_X1  g1067(.A1(new_n1257), .A2(KEYINPUT58), .ZN(new_n1268));
  OAI211_X1 g1068(.A(new_n1254), .B(new_n202), .C1(G33), .C2(G41), .ZN(new_n1269));
  NAND4_X1  g1069(.A1(new_n1258), .A2(new_n1267), .A3(new_n1268), .A4(new_n1269), .ZN(new_n1270));
  AOI21_X1  g1070(.A(new_n1247), .B1(new_n1270), .B2(new_n814), .ZN(new_n1271));
  NAND2_X1  g1071(.A1(new_n1246), .A2(new_n1271), .ZN(new_n1272));
  NAND2_X1  g1072(.A1(new_n1245), .A2(new_n1272), .ZN(new_n1273));
  INV_X1    g1073(.A(new_n1273), .ZN(new_n1274));
  NAND2_X1  g1074(.A1(new_n1244), .A2(new_n1274), .ZN(G375));
  NAND2_X1  g1075(.A1(new_n1178), .A2(new_n1180), .ZN(new_n1276));
  NAND2_X1  g1076(.A1(new_n1276), .A2(new_n1235), .ZN(new_n1277));
  XOR2_X1   g1077(.A(new_n1015), .B(KEYINPUT122), .Z(new_n1278));
  NAND3_X1  g1078(.A1(new_n1277), .A2(new_n1181), .A3(new_n1278), .ZN(new_n1279));
  NOR2_X1   g1079(.A1(new_n1235), .A2(new_n1105), .ZN(new_n1280));
  AOI22_X1  g1080(.A1(G294), .A2(new_n877), .B1(new_n847), .B2(G283), .ZN(new_n1281));
  OAI21_X1  g1081(.A(new_n1281), .B1(new_n319), .B2(new_n821), .ZN(new_n1282));
  OAI211_X1 g1082(.A(new_n1097), .B(new_n556), .C1(new_n221), .C2(new_n834), .ZN(new_n1283));
  AOI21_X1  g1083(.A(new_n1283), .B1(G303), .B2(new_n837), .ZN(new_n1284));
  OAI21_X1  g1084(.A(new_n1284), .B1(new_n459), .B2(new_n840), .ZN(new_n1285));
  AOI211_X1 g1085(.A(new_n1282), .B(new_n1285), .C1(G116), .C2(new_n842), .ZN(new_n1286));
  OAI221_X1 g1086(.A(new_n353), .B1(new_n202), .B2(new_n830), .C1(new_n834), .C2(new_n365), .ZN(new_n1287));
  INV_X1    g1087(.A(G128), .ZN(new_n1288));
  OAI21_X1  g1088(.A(new_n1249), .B1(new_n851), .B2(new_n1288), .ZN(new_n1289));
  AOI211_X1 g1089(.A(new_n1287), .B(new_n1289), .C1(G150), .C2(new_n861), .ZN(new_n1290));
  XNOR2_X1  g1090(.A(new_n1290), .B(KEYINPUT124), .ZN(new_n1291));
  OAI22_X1  g1091(.A1(new_n855), .A2(new_n1051), .B1(new_n885), .B2(new_n827), .ZN(new_n1292));
  AOI21_X1  g1092(.A(new_n1292), .B1(new_n842), .B2(new_n1199), .ZN(new_n1293));
  AOI21_X1  g1093(.A(new_n1286), .B1(new_n1291), .B2(new_n1293), .ZN(new_n1294));
  INV_X1    g1094(.A(new_n814), .ZN(new_n1295));
  OAI221_X1 g1095(.A(new_n799), .B1(G68), .B2(new_n1186), .C1(new_n1294), .C2(new_n1295), .ZN(new_n1296));
  NOR3_X1   g1096(.A1(new_n1144), .A2(new_n1145), .A3(new_n812), .ZN(new_n1297));
  OR2_X1    g1097(.A1(new_n1297), .A2(KEYINPUT123), .ZN(new_n1298));
  NAND2_X1  g1098(.A1(new_n1297), .A2(KEYINPUT123), .ZN(new_n1299));
  AOI21_X1  g1099(.A(new_n1296), .B1(new_n1298), .B2(new_n1299), .ZN(new_n1300));
  NOR2_X1   g1100(.A1(new_n1280), .A2(new_n1300), .ZN(new_n1301));
  NAND2_X1  g1101(.A1(new_n1279), .A2(new_n1301), .ZN(G381));
  AOI21_X1  g1102(.A(new_n1273), .B1(new_n1239), .B2(new_n1243), .ZN(new_n1303));
  INV_X1    g1103(.A(G378), .ZN(new_n1304));
  NAND2_X1  g1104(.A1(new_n1303), .A2(new_n1304), .ZN(new_n1305));
  INV_X1    g1105(.A(G390), .ZN(new_n1306));
  INV_X1    g1106(.A(G384), .ZN(new_n1307));
  NOR2_X1   g1107(.A1(new_n1041), .A2(new_n1114), .ZN(new_n1308));
  AOI22_X1  g1108(.A1(new_n1308), .A2(KEYINPUT116), .B1(new_n1040), .B2(new_n1039), .ZN(new_n1309));
  AOI211_X1 g1109(.A(G396), .B(new_n1106), .C1(new_n1309), .C2(new_n1115), .ZN(new_n1310));
  NAND3_X1  g1110(.A1(new_n1306), .A2(new_n1307), .A3(new_n1310), .ZN(new_n1311));
  OR4_X1    g1111(.A1(G387), .A2(new_n1305), .A3(G381), .A4(new_n1311), .ZN(G407));
  OAI211_X1 g1112(.A(G407), .B(G213), .C1(G343), .C2(new_n1305), .ZN(G409));
  INV_X1    g1113(.A(G343), .ZN(new_n1314));
  NAND2_X1  g1114(.A1(new_n1314), .A2(G213), .ZN(new_n1315));
  INV_X1    g1115(.A(KEYINPUT125), .ZN(new_n1316));
  NAND2_X1  g1116(.A1(new_n1181), .A2(new_n1109), .ZN(new_n1317));
  NAND2_X1  g1117(.A1(new_n1277), .A2(KEYINPUT60), .ZN(new_n1318));
  INV_X1    g1118(.A(KEYINPUT60), .ZN(new_n1319));
  NAND3_X1  g1119(.A1(new_n1276), .A2(new_n1235), .A3(new_n1319), .ZN(new_n1320));
  AOI21_X1  g1120(.A(new_n1317), .B1(new_n1318), .B2(new_n1320), .ZN(new_n1321));
  INV_X1    g1121(.A(new_n1301), .ZN(new_n1322));
  OAI211_X1 g1122(.A(new_n1316), .B(new_n1307), .C1(new_n1321), .C2(new_n1322), .ZN(new_n1323));
  AND2_X1   g1123(.A1(new_n1181), .A2(new_n1109), .ZN(new_n1324));
  INV_X1    g1124(.A(new_n1320), .ZN(new_n1325));
  AOI21_X1  g1125(.A(new_n1319), .B1(new_n1276), .B2(new_n1235), .ZN(new_n1326));
  OAI21_X1  g1126(.A(new_n1324), .B1(new_n1325), .B2(new_n1326), .ZN(new_n1327));
  NAND3_X1  g1127(.A1(new_n1327), .A2(G384), .A3(new_n1301), .ZN(new_n1328));
  NAND2_X1  g1128(.A1(new_n1323), .A2(new_n1328), .ZN(new_n1329));
  NAND2_X1  g1129(.A1(new_n1327), .A2(new_n1301), .ZN(new_n1330));
  AOI21_X1  g1130(.A(new_n1316), .B1(new_n1330), .B2(new_n1307), .ZN(new_n1331));
  NOR2_X1   g1131(.A1(new_n1329), .A2(new_n1331), .ZN(new_n1332));
  AOI21_X1  g1132(.A(new_n1242), .B1(new_n1238), .B2(new_n1237), .ZN(new_n1333));
  NOR3_X1   g1133(.A1(new_n1333), .A2(new_n1304), .A3(new_n1273), .ZN(new_n1334));
  INV_X1    g1134(.A(new_n1240), .ZN(new_n1335));
  AOI22_X1  g1135(.A1(new_n1335), .A2(new_n1044), .B1(new_n1246), .B2(new_n1271), .ZN(new_n1336));
  NAND4_X1  g1136(.A1(new_n1229), .A2(new_n1233), .A3(new_n1236), .A4(new_n1278), .ZN(new_n1337));
  AOI21_X1  g1137(.A(G378), .B1(new_n1336), .B2(new_n1337), .ZN(new_n1338));
  OAI211_X1 g1138(.A(new_n1315), .B(new_n1332), .C1(new_n1334), .C2(new_n1338), .ZN(new_n1339));
  NAND2_X1  g1139(.A1(new_n1339), .A2(KEYINPUT62), .ZN(new_n1340));
  INV_X1    g1140(.A(KEYINPUT61), .ZN(new_n1341));
  NAND3_X1  g1141(.A1(new_n1244), .A2(G378), .A3(new_n1274), .ZN(new_n1342));
  INV_X1    g1142(.A(new_n1338), .ZN(new_n1343));
  NAND2_X1  g1143(.A1(new_n1342), .A2(new_n1343), .ZN(new_n1344));
  INV_X1    g1144(.A(KEYINPUT62), .ZN(new_n1345));
  NAND4_X1  g1145(.A1(new_n1344), .A2(new_n1345), .A3(new_n1315), .A4(new_n1332), .ZN(new_n1346));
  INV_X1    g1146(.A(new_n1315), .ZN(new_n1347));
  NAND2_X1  g1147(.A1(new_n1347), .A2(G2897), .ZN(new_n1348));
  XOR2_X1   g1148(.A(new_n1348), .B(KEYINPUT126), .Z(new_n1349));
  OAI21_X1  g1149(.A(new_n1349), .B1(new_n1329), .B2(new_n1331), .ZN(new_n1350));
  OAI21_X1  g1150(.A(new_n1307), .B1(new_n1321), .B2(new_n1322), .ZN(new_n1351));
  NAND2_X1  g1151(.A1(new_n1351), .A2(KEYINPUT125), .ZN(new_n1352));
  INV_X1    g1152(.A(new_n1349), .ZN(new_n1353));
  NAND4_X1  g1153(.A1(new_n1352), .A2(new_n1323), .A3(new_n1328), .A4(new_n1353), .ZN(new_n1354));
  AND2_X1   g1154(.A1(new_n1350), .A2(new_n1354), .ZN(new_n1355));
  AOI21_X1  g1155(.A(new_n1338), .B1(new_n1303), .B2(G378), .ZN(new_n1356));
  OAI21_X1  g1156(.A(new_n1355), .B1(new_n1356), .B2(new_n1347), .ZN(new_n1357));
  NAND4_X1  g1157(.A1(new_n1340), .A2(new_n1341), .A3(new_n1346), .A4(new_n1357), .ZN(new_n1358));
  INV_X1    g1158(.A(new_n1015), .ZN(new_n1359));
  AOI21_X1  g1159(.A(new_n1108), .B1(new_n1031), .B2(new_n1033), .ZN(new_n1360));
  OAI21_X1  g1160(.A(new_n1359), .B1(new_n1360), .B2(new_n1040), .ZN(new_n1361));
  AOI21_X1  g1161(.A(new_n1013), .B1(new_n1361), .B2(new_n1105), .ZN(new_n1362));
  INV_X1    g1162(.A(new_n1073), .ZN(new_n1363));
  OAI21_X1  g1163(.A(new_n1306), .B1(new_n1362), .B2(new_n1363), .ZN(new_n1364));
  NAND3_X1  g1164(.A1(new_n1045), .A2(new_n1073), .A3(G390), .ZN(new_n1365));
  INV_X1    g1165(.A(KEYINPUT127), .ZN(new_n1366));
  NAND2_X1  g1166(.A1(G393), .A2(G396), .ZN(new_n1367));
  NAND2_X1  g1167(.A1(new_n1309), .A2(new_n1115), .ZN(new_n1368));
  INV_X1    g1168(.A(G396), .ZN(new_n1369));
  NAND3_X1  g1169(.A1(new_n1368), .A2(new_n1369), .A3(new_n1107), .ZN(new_n1370));
  AOI21_X1  g1170(.A(new_n1366), .B1(new_n1367), .B2(new_n1370), .ZN(new_n1371));
  NAND3_X1  g1171(.A1(new_n1364), .A2(new_n1365), .A3(new_n1371), .ZN(new_n1372));
  AOI21_X1  g1172(.A(new_n1369), .B1(new_n1368), .B2(new_n1107), .ZN(new_n1373));
  OAI21_X1  g1173(.A(KEYINPUT127), .B1(new_n1373), .B2(new_n1310), .ZN(new_n1374));
  NAND3_X1  g1174(.A1(new_n1374), .A2(G387), .A3(new_n1306), .ZN(new_n1375));
  NOR2_X1   g1175(.A1(new_n1373), .A2(new_n1310), .ZN(new_n1376));
  NAND4_X1  g1176(.A1(new_n1376), .A2(new_n1045), .A3(new_n1073), .A4(G390), .ZN(new_n1377));
  AND3_X1   g1177(.A1(new_n1372), .A2(new_n1375), .A3(new_n1377), .ZN(new_n1378));
  NAND2_X1  g1178(.A1(new_n1358), .A2(new_n1378), .ZN(new_n1379));
  NAND4_X1  g1179(.A1(new_n1344), .A2(KEYINPUT63), .A3(new_n1315), .A4(new_n1332), .ZN(new_n1380));
  NOR2_X1   g1180(.A1(new_n1378), .A2(KEYINPUT61), .ZN(new_n1381));
  INV_X1    g1181(.A(KEYINPUT63), .ZN(new_n1382));
  NAND2_X1  g1182(.A1(new_n1344), .A2(new_n1315), .ZN(new_n1383));
  AOI21_X1  g1183(.A(new_n1382), .B1(new_n1383), .B2(new_n1355), .ZN(new_n1384));
  INV_X1    g1184(.A(new_n1339), .ZN(new_n1385));
  OAI211_X1 g1185(.A(new_n1380), .B(new_n1381), .C1(new_n1384), .C2(new_n1385), .ZN(new_n1386));
  NAND2_X1  g1186(.A1(new_n1379), .A2(new_n1386), .ZN(G405));
  NAND2_X1  g1187(.A1(G375), .A2(G378), .ZN(new_n1388));
  NAND3_X1  g1188(.A1(new_n1378), .A2(new_n1305), .A3(new_n1388), .ZN(new_n1389));
  NAND2_X1  g1189(.A1(new_n1388), .A2(new_n1305), .ZN(new_n1390));
  NAND3_X1  g1190(.A1(new_n1372), .A2(new_n1375), .A3(new_n1377), .ZN(new_n1391));
  NAND2_X1  g1191(.A1(new_n1390), .A2(new_n1391), .ZN(new_n1392));
  AND3_X1   g1192(.A1(new_n1389), .A2(new_n1392), .A3(new_n1332), .ZN(new_n1393));
  AOI21_X1  g1193(.A(new_n1332), .B1(new_n1389), .B2(new_n1392), .ZN(new_n1394));
  NOR2_X1   g1194(.A1(new_n1393), .A2(new_n1394), .ZN(G402));
endmodule


