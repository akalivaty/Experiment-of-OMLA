//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 1 0 0 0 1 0 0 0 0 1 1 1 1 1 1 1 0 0 1 1 1 0 1 0 0 1 0 1 0 0 1 1 0 1 0 0 1 0 0 1 0 0 0 0 1 1 0 1 1 0 0 0 1 1 0 1 1 1 0 0 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:24:26 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n619, new_n620, new_n621, new_n622,
    new_n623, new_n624, new_n625, new_n627, new_n628, new_n629, new_n630,
    new_n631, new_n632, new_n633, new_n635, new_n636, new_n637, new_n638,
    new_n639, new_n640, new_n641, new_n642, new_n643, new_n644, new_n645,
    new_n646, new_n647, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n702, new_n704, new_n705, new_n706,
    new_n707, new_n709, new_n710, new_n711, new_n712, new_n713, new_n714,
    new_n715, new_n716, new_n717, new_n718, new_n719, new_n720, new_n721,
    new_n722, new_n723, new_n725, new_n726, new_n727, new_n728, new_n729,
    new_n730, new_n731, new_n732, new_n733, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n753, new_n754, new_n755, new_n756, new_n757, new_n758, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n786, new_n787, new_n788, new_n789,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n919,
    new_n920, new_n921, new_n923, new_n924, new_n925, new_n926, new_n927,
    new_n928, new_n930, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n939, new_n941, new_n942, new_n943,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n972, new_n973,
    new_n974, new_n975, new_n976, new_n977, new_n978, new_n979, new_n980,
    new_n981, new_n982, new_n983, new_n984, new_n985, new_n986, new_n987;
  INV_X1    g000(.A(KEYINPUT67), .ZN(new_n187));
  INV_X1    g001(.A(G134), .ZN(new_n188));
  OAI21_X1  g002(.A(KEYINPUT11), .B1(new_n188), .B2(G137), .ZN(new_n189));
  INV_X1    g003(.A(KEYINPUT11), .ZN(new_n190));
  INV_X1    g004(.A(G137), .ZN(new_n191));
  NAND3_X1  g005(.A1(new_n190), .A2(new_n191), .A3(G134), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n189), .A2(new_n192), .ZN(new_n193));
  INV_X1    g007(.A(G131), .ZN(new_n194));
  INV_X1    g008(.A(KEYINPUT64), .ZN(new_n195));
  OAI21_X1  g009(.A(new_n195), .B1(new_n191), .B2(G134), .ZN(new_n196));
  NAND3_X1  g010(.A1(new_n188), .A2(KEYINPUT64), .A3(G137), .ZN(new_n197));
  NAND4_X1  g011(.A1(new_n193), .A2(new_n194), .A3(new_n196), .A4(new_n197), .ZN(new_n198));
  INV_X1    g012(.A(KEYINPUT65), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n198), .A2(new_n199), .ZN(new_n200));
  AND2_X1   g014(.A1(new_n196), .A2(new_n197), .ZN(new_n201));
  NAND4_X1  g015(.A1(new_n201), .A2(KEYINPUT65), .A3(new_n194), .A4(new_n193), .ZN(new_n202));
  AND2_X1   g016(.A1(new_n200), .A2(new_n202), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n191), .A2(G134), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n188), .A2(G137), .ZN(new_n205));
  AOI21_X1  g019(.A(new_n194), .B1(new_n204), .B2(new_n205), .ZN(new_n206));
  OAI21_X1  g020(.A(new_n187), .B1(new_n203), .B2(new_n206), .ZN(new_n207));
  AOI21_X1  g021(.A(new_n206), .B1(new_n200), .B2(new_n202), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n208), .A2(KEYINPUT67), .ZN(new_n209));
  INV_X1    g023(.A(G146), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n210), .A2(G143), .ZN(new_n211));
  INV_X1    g025(.A(G143), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n212), .A2(G146), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n211), .A2(new_n213), .ZN(new_n214));
  INV_X1    g028(.A(KEYINPUT1), .ZN(new_n215));
  AOI21_X1  g029(.A(new_n215), .B1(G143), .B2(new_n210), .ZN(new_n216));
  INV_X1    g030(.A(G128), .ZN(new_n217));
  OAI21_X1  g031(.A(new_n214), .B1(new_n216), .B2(new_n217), .ZN(new_n218));
  XNOR2_X1  g032(.A(G143), .B(G146), .ZN(new_n219));
  NOR2_X1   g033(.A1(new_n217), .A2(KEYINPUT1), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n219), .A2(new_n220), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n218), .A2(new_n221), .ZN(new_n222));
  NAND3_X1  g036(.A1(new_n207), .A2(new_n209), .A3(new_n222), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n200), .A2(new_n202), .ZN(new_n224));
  AOI21_X1  g038(.A(new_n194), .B1(new_n201), .B2(new_n193), .ZN(new_n225));
  INV_X1    g039(.A(new_n225), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n224), .A2(new_n226), .ZN(new_n227));
  INV_X1    g041(.A(KEYINPUT66), .ZN(new_n228));
  INV_X1    g042(.A(KEYINPUT0), .ZN(new_n229));
  OAI211_X1 g043(.A(new_n211), .B(new_n213), .C1(new_n229), .C2(new_n217), .ZN(new_n230));
  XOR2_X1   g044(.A(KEYINPUT0), .B(G128), .Z(new_n231));
  OAI21_X1  g045(.A(new_n230), .B1(new_n231), .B2(new_n219), .ZN(new_n232));
  NAND3_X1  g046(.A1(new_n227), .A2(new_n228), .A3(new_n232), .ZN(new_n233));
  AOI21_X1  g047(.A(new_n225), .B1(new_n200), .B2(new_n202), .ZN(new_n234));
  INV_X1    g048(.A(new_n232), .ZN(new_n235));
  OAI21_X1  g049(.A(KEYINPUT66), .B1(new_n234), .B2(new_n235), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n233), .A2(new_n236), .ZN(new_n237));
  INV_X1    g051(.A(KEYINPUT30), .ZN(new_n238));
  NAND3_X1  g052(.A1(new_n223), .A2(new_n237), .A3(new_n238), .ZN(new_n239));
  INV_X1    g053(.A(KEYINPUT68), .ZN(new_n240));
  XNOR2_X1  g054(.A(new_n232), .B(new_n240), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n227), .A2(new_n241), .ZN(new_n242));
  OAI21_X1  g056(.A(new_n222), .B1(new_n208), .B2(KEYINPUT69), .ZN(new_n243));
  INV_X1    g057(.A(KEYINPUT69), .ZN(new_n244));
  AOI211_X1 g058(.A(new_n244), .B(new_n206), .C1(new_n200), .C2(new_n202), .ZN(new_n245));
  OAI21_X1  g059(.A(new_n242), .B1(new_n243), .B2(new_n245), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n246), .A2(KEYINPUT30), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n239), .A2(new_n247), .ZN(new_n248));
  XOR2_X1   g062(.A(G116), .B(G119), .Z(new_n249));
  XNOR2_X1  g063(.A(KEYINPUT2), .B(G113), .ZN(new_n250));
  XNOR2_X1  g064(.A(new_n249), .B(new_n250), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n248), .A2(new_n251), .ZN(new_n252));
  INV_X1    g066(.A(new_n251), .ZN(new_n253));
  OAI211_X1 g067(.A(new_n253), .B(new_n242), .C1(new_n243), .C2(new_n245), .ZN(new_n254));
  NOR2_X1   g068(.A1(G237), .A2(G953), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n255), .A2(G210), .ZN(new_n256));
  XOR2_X1   g070(.A(new_n256), .B(KEYINPUT27), .Z(new_n257));
  XNOR2_X1  g071(.A(KEYINPUT26), .B(G101), .ZN(new_n258));
  XOR2_X1   g072(.A(new_n257), .B(new_n258), .Z(new_n259));
  NAND3_X1  g073(.A1(new_n252), .A2(new_n254), .A3(new_n259), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n260), .A2(KEYINPUT31), .ZN(new_n261));
  INV_X1    g075(.A(new_n259), .ZN(new_n262));
  INV_X1    g076(.A(KEYINPUT28), .ZN(new_n263));
  AOI21_X1  g077(.A(KEYINPUT70), .B1(new_n254), .B2(new_n263), .ZN(new_n264));
  INV_X1    g078(.A(new_n264), .ZN(new_n265));
  NAND3_X1  g079(.A1(new_n254), .A2(KEYINPUT70), .A3(new_n263), .ZN(new_n266));
  NAND2_X1  g080(.A1(new_n265), .A2(new_n266), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n223), .A2(new_n237), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n268), .A2(new_n251), .ZN(new_n269));
  AOI21_X1  g083(.A(new_n263), .B1(new_n269), .B2(new_n254), .ZN(new_n270));
  OAI21_X1  g084(.A(new_n262), .B1(new_n267), .B2(new_n270), .ZN(new_n271));
  INV_X1    g085(.A(new_n254), .ZN(new_n272));
  AOI21_X1  g086(.A(new_n272), .B1(new_n248), .B2(new_n251), .ZN(new_n273));
  INV_X1    g087(.A(KEYINPUT31), .ZN(new_n274));
  NAND3_X1  g088(.A1(new_n273), .A2(new_n274), .A3(new_n259), .ZN(new_n275));
  NAND3_X1  g089(.A1(new_n261), .A2(new_n271), .A3(new_n275), .ZN(new_n276));
  NOR2_X1   g090(.A1(G472), .A2(G902), .ZN(new_n277));
  INV_X1    g091(.A(new_n277), .ZN(new_n278));
  INV_X1    g092(.A(KEYINPUT32), .ZN(new_n279));
  NOR2_X1   g093(.A1(new_n278), .A2(new_n279), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n276), .A2(new_n280), .ZN(new_n281));
  AND3_X1   g095(.A1(new_n254), .A2(KEYINPUT70), .A3(new_n263), .ZN(new_n282));
  NOR2_X1   g096(.A1(new_n282), .A2(new_n264), .ZN(new_n283));
  AOI21_X1  g097(.A(new_n253), .B1(new_n223), .B2(new_n237), .ZN(new_n284));
  OAI21_X1  g098(.A(KEYINPUT28), .B1(new_n284), .B2(new_n272), .ZN(new_n285));
  NAND3_X1  g099(.A1(new_n283), .A2(new_n285), .A3(new_n259), .ZN(new_n286));
  INV_X1    g100(.A(KEYINPUT29), .ZN(new_n287));
  AOI21_X1  g101(.A(new_n253), .B1(new_n239), .B2(new_n247), .ZN(new_n288));
  OAI21_X1  g102(.A(new_n262), .B1(new_n288), .B2(new_n272), .ZN(new_n289));
  NAND3_X1  g103(.A1(new_n286), .A2(new_n287), .A3(new_n289), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n246), .A2(new_n251), .ZN(new_n291));
  AOI21_X1  g105(.A(new_n263), .B1(new_n291), .B2(new_n254), .ZN(new_n292));
  NOR3_X1   g106(.A1(new_n292), .A2(new_n282), .A3(new_n264), .ZN(new_n293));
  NOR2_X1   g107(.A1(new_n262), .A2(new_n287), .ZN(new_n294));
  AOI21_X1  g108(.A(G902), .B1(new_n293), .B2(new_n294), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n290), .A2(new_n295), .ZN(new_n296));
  NAND2_X1  g110(.A1(new_n296), .A2(G472), .ZN(new_n297));
  AOI21_X1  g111(.A(new_n274), .B1(new_n273), .B2(new_n259), .ZN(new_n298));
  NOR4_X1   g112(.A1(new_n288), .A2(KEYINPUT31), .A3(new_n272), .A4(new_n262), .ZN(new_n299));
  NOR2_X1   g113(.A1(new_n298), .A2(new_n299), .ZN(new_n300));
  AOI21_X1  g114(.A(new_n278), .B1(new_n300), .B2(new_n271), .ZN(new_n301));
  OAI211_X1 g115(.A(new_n281), .B(new_n297), .C1(new_n301), .C2(KEYINPUT32), .ZN(new_n302));
  INV_X1    g116(.A(KEYINPUT23), .ZN(new_n303));
  INV_X1    g117(.A(G119), .ZN(new_n304));
  OAI21_X1  g118(.A(new_n303), .B1(new_n304), .B2(G128), .ZN(new_n305));
  NAND3_X1  g119(.A1(new_n217), .A2(KEYINPUT23), .A3(G119), .ZN(new_n306));
  OAI211_X1 g120(.A(new_n305), .B(new_n306), .C1(G119), .C2(new_n217), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n307), .A2(G110), .ZN(new_n308));
  XOR2_X1   g122(.A(KEYINPUT24), .B(G110), .Z(new_n309));
  XNOR2_X1  g123(.A(G119), .B(G128), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n309), .A2(new_n310), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n308), .A2(new_n311), .ZN(new_n312));
  INV_X1    g126(.A(G140), .ZN(new_n313));
  NAND2_X1  g127(.A1(new_n313), .A2(G125), .ZN(new_n314));
  NOR2_X1   g128(.A1(new_n314), .A2(KEYINPUT16), .ZN(new_n315));
  INV_X1    g129(.A(KEYINPUT72), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n315), .A2(new_n316), .ZN(new_n317));
  XNOR2_X1  g131(.A(G125), .B(G140), .ZN(new_n318));
  AOI21_X1  g132(.A(KEYINPUT72), .B1(new_n318), .B2(KEYINPUT16), .ZN(new_n319));
  OAI21_X1  g133(.A(new_n317), .B1(new_n319), .B2(new_n315), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n320), .A2(new_n210), .ZN(new_n321));
  OAI211_X1 g135(.A(G146), .B(new_n317), .C1(new_n319), .C2(new_n315), .ZN(new_n322));
  AOI21_X1  g136(.A(new_n312), .B1(new_n321), .B2(new_n322), .ZN(new_n323));
  XOR2_X1   g137(.A(KEYINPUT73), .B(G110), .Z(new_n324));
  OAI22_X1  g138(.A1(new_n307), .A2(new_n324), .B1(new_n310), .B2(new_n309), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n318), .A2(new_n210), .ZN(new_n326));
  AND3_X1   g140(.A1(new_n322), .A2(new_n325), .A3(new_n326), .ZN(new_n327));
  XNOR2_X1  g141(.A(KEYINPUT22), .B(G137), .ZN(new_n328));
  INV_X1    g142(.A(G953), .ZN(new_n329));
  AND3_X1   g143(.A1(new_n329), .A2(G221), .A3(G234), .ZN(new_n330));
  XNOR2_X1  g144(.A(new_n328), .B(new_n330), .ZN(new_n331));
  OR3_X1    g145(.A1(new_n323), .A2(new_n327), .A3(new_n331), .ZN(new_n332));
  INV_X1    g146(.A(G902), .ZN(new_n333));
  OAI21_X1  g147(.A(new_n331), .B1(new_n323), .B2(new_n327), .ZN(new_n334));
  NAND3_X1  g148(.A1(new_n332), .A2(new_n333), .A3(new_n334), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n335), .A2(KEYINPUT74), .ZN(new_n336));
  INV_X1    g150(.A(KEYINPUT75), .ZN(new_n337));
  INV_X1    g151(.A(KEYINPUT25), .ZN(new_n338));
  INV_X1    g152(.A(KEYINPUT74), .ZN(new_n339));
  NAND4_X1  g153(.A1(new_n332), .A2(new_n339), .A3(new_n333), .A4(new_n334), .ZN(new_n340));
  NAND4_X1  g154(.A1(new_n336), .A2(new_n337), .A3(new_n338), .A4(new_n340), .ZN(new_n341));
  XNOR2_X1  g155(.A(KEYINPUT71), .B(G217), .ZN(new_n342));
  AOI21_X1  g156(.A(new_n342), .B1(G234), .B2(new_n333), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n341), .A2(new_n343), .ZN(new_n344));
  INV_X1    g158(.A(new_n344), .ZN(new_n345));
  OAI21_X1  g159(.A(KEYINPUT75), .B1(new_n335), .B2(new_n338), .ZN(new_n346));
  AOI21_X1  g160(.A(KEYINPUT25), .B1(new_n335), .B2(KEYINPUT74), .ZN(new_n347));
  AOI21_X1  g161(.A(new_n346), .B1(new_n340), .B2(new_n347), .ZN(new_n348));
  INV_X1    g162(.A(new_n348), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n345), .A2(new_n349), .ZN(new_n350));
  NOR2_X1   g164(.A1(new_n343), .A2(G902), .ZN(new_n351));
  NAND3_X1  g165(.A1(new_n332), .A2(new_n334), .A3(new_n351), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n350), .A2(new_n352), .ZN(new_n353));
  INV_X1    g167(.A(new_n353), .ZN(new_n354));
  INV_X1    g168(.A(G237), .ZN(new_n355));
  NAND3_X1  g169(.A1(new_n355), .A2(new_n329), .A3(G214), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n356), .A2(new_n212), .ZN(new_n357));
  NAND3_X1  g171(.A1(new_n255), .A2(G143), .A3(G214), .ZN(new_n358));
  NAND2_X1  g172(.A1(new_n357), .A2(new_n358), .ZN(new_n359));
  AOI21_X1  g173(.A(KEYINPUT88), .B1(new_n359), .B2(G131), .ZN(new_n360));
  INV_X1    g174(.A(KEYINPUT88), .ZN(new_n361));
  AOI211_X1 g175(.A(new_n361), .B(new_n194), .C1(new_n357), .C2(new_n358), .ZN(new_n362));
  OAI21_X1  g176(.A(KEYINPUT17), .B1(new_n360), .B2(new_n362), .ZN(new_n363));
  AND4_X1   g177(.A1(G143), .A2(new_n355), .A3(new_n329), .A4(G214), .ZN(new_n364));
  AOI21_X1  g178(.A(G143), .B1(new_n255), .B2(G214), .ZN(new_n365));
  OAI21_X1  g179(.A(G131), .B1(new_n364), .B2(new_n365), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n366), .A2(new_n361), .ZN(new_n367));
  INV_X1    g181(.A(KEYINPUT17), .ZN(new_n368));
  OAI211_X1 g182(.A(KEYINPUT88), .B(G131), .C1(new_n364), .C2(new_n365), .ZN(new_n369));
  NAND3_X1  g183(.A1(new_n357), .A2(new_n194), .A3(new_n358), .ZN(new_n370));
  NAND4_X1  g184(.A1(new_n367), .A2(new_n368), .A3(new_n369), .A4(new_n370), .ZN(new_n371));
  NAND4_X1  g185(.A1(new_n363), .A2(new_n371), .A3(new_n321), .A4(new_n322), .ZN(new_n372));
  XNOR2_X1  g186(.A(G113), .B(G122), .ZN(new_n373));
  INV_X1    g187(.A(G104), .ZN(new_n374));
  XNOR2_X1  g188(.A(new_n373), .B(new_n374), .ZN(new_n375));
  INV_X1    g189(.A(KEYINPUT86), .ZN(new_n376));
  INV_X1    g190(.A(G125), .ZN(new_n377));
  NOR2_X1   g191(.A1(new_n377), .A2(G140), .ZN(new_n378));
  NOR2_X1   g192(.A1(new_n313), .A2(G125), .ZN(new_n379));
  OAI21_X1  g193(.A(new_n376), .B1(new_n378), .B2(new_n379), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n377), .A2(G140), .ZN(new_n381));
  NAND3_X1  g195(.A1(new_n314), .A2(new_n381), .A3(KEYINPUT86), .ZN(new_n382));
  NAND3_X1  g196(.A1(new_n380), .A2(G146), .A3(new_n382), .ZN(new_n383));
  NAND2_X1  g197(.A1(new_n383), .A2(new_n326), .ZN(new_n384));
  NOR2_X1   g198(.A1(new_n364), .A2(new_n365), .ZN(new_n385));
  INV_X1    g199(.A(KEYINPUT87), .ZN(new_n386));
  AOI22_X1  g200(.A1(new_n385), .A2(new_n386), .B1(KEYINPUT18), .B2(G131), .ZN(new_n387));
  NAND2_X1  g201(.A1(KEYINPUT18), .A2(G131), .ZN(new_n388));
  NOR3_X1   g202(.A1(new_n359), .A2(KEYINPUT87), .A3(new_n388), .ZN(new_n389));
  OAI21_X1  g203(.A(new_n384), .B1(new_n387), .B2(new_n389), .ZN(new_n390));
  NAND3_X1  g204(.A1(new_n372), .A2(new_n375), .A3(new_n390), .ZN(new_n391));
  INV_X1    g205(.A(new_n391), .ZN(new_n392));
  AOI21_X1  g206(.A(new_n375), .B1(new_n372), .B2(new_n390), .ZN(new_n393));
  OAI21_X1  g207(.A(new_n333), .B1(new_n392), .B2(new_n393), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n394), .A2(G475), .ZN(new_n395));
  NOR2_X1   g209(.A1(G475), .A2(G902), .ZN(new_n396));
  INV_X1    g210(.A(new_n396), .ZN(new_n397));
  AND3_X1   g211(.A1(new_n367), .A2(new_n369), .A3(new_n370), .ZN(new_n398));
  NAND3_X1  g212(.A1(new_n380), .A2(KEYINPUT19), .A3(new_n382), .ZN(new_n399));
  INV_X1    g213(.A(KEYINPUT19), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n318), .A2(new_n400), .ZN(new_n401));
  NAND3_X1  g215(.A1(new_n399), .A2(new_n210), .A3(new_n401), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n402), .A2(new_n322), .ZN(new_n403));
  OAI21_X1  g217(.A(new_n390), .B1(new_n398), .B2(new_n403), .ZN(new_n404));
  INV_X1    g218(.A(new_n375), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n404), .A2(new_n405), .ZN(new_n406));
  AOI21_X1  g220(.A(new_n397), .B1(new_n391), .B2(new_n406), .ZN(new_n407));
  NAND2_X1  g221(.A1(new_n391), .A2(new_n406), .ZN(new_n408));
  NAND2_X1  g222(.A1(new_n408), .A2(KEYINPUT89), .ZN(new_n409));
  INV_X1    g223(.A(KEYINPUT20), .ZN(new_n410));
  AOI21_X1  g224(.A(new_n407), .B1(new_n409), .B2(new_n410), .ZN(new_n411));
  INV_X1    g225(.A(KEYINPUT89), .ZN(new_n412));
  AND4_X1   g226(.A1(new_n412), .A2(new_n408), .A3(new_n410), .A4(new_n396), .ZN(new_n413));
  OAI21_X1  g227(.A(new_n395), .B1(new_n411), .B2(new_n413), .ZN(new_n414));
  INV_X1    g228(.A(KEYINPUT90), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n414), .A2(new_n415), .ZN(new_n416));
  NAND2_X1  g230(.A1(new_n408), .A2(new_n396), .ZN(new_n417));
  AOI21_X1  g231(.A(new_n412), .B1(new_n391), .B2(new_n406), .ZN(new_n418));
  OAI21_X1  g232(.A(new_n417), .B1(KEYINPUT20), .B2(new_n418), .ZN(new_n419));
  NAND3_X1  g233(.A1(new_n409), .A2(new_n410), .A3(new_n407), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n419), .A2(new_n420), .ZN(new_n421));
  NAND3_X1  g235(.A1(new_n421), .A2(KEYINPUT90), .A3(new_n395), .ZN(new_n422));
  INV_X1    g236(.A(G107), .ZN(new_n423));
  INV_X1    g237(.A(G122), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n424), .A2(G116), .ZN(new_n425));
  AOI21_X1  g239(.A(new_n423), .B1(new_n425), .B2(KEYINPUT14), .ZN(new_n426));
  XNOR2_X1  g240(.A(G116), .B(G122), .ZN(new_n427));
  XNOR2_X1  g241(.A(new_n426), .B(new_n427), .ZN(new_n428));
  XNOR2_X1  g242(.A(G128), .B(G143), .ZN(new_n429));
  XNOR2_X1  g243(.A(new_n429), .B(KEYINPUT92), .ZN(new_n430));
  AND2_X1   g244(.A1(new_n430), .A2(G134), .ZN(new_n431));
  NOR2_X1   g245(.A1(new_n430), .A2(G134), .ZN(new_n432));
  OAI21_X1  g246(.A(new_n428), .B1(new_n431), .B2(new_n432), .ZN(new_n433));
  XOR2_X1   g247(.A(KEYINPUT91), .B(KEYINPUT13), .Z(new_n434));
  NAND3_X1  g248(.A1(new_n434), .A2(G128), .A3(new_n212), .ZN(new_n435));
  INV_X1    g249(.A(new_n429), .ZN(new_n436));
  OAI211_X1 g250(.A(new_n435), .B(G134), .C1(new_n436), .C2(new_n434), .ZN(new_n437));
  XNOR2_X1  g251(.A(new_n427), .B(new_n423), .ZN(new_n438));
  OAI211_X1 g252(.A(new_n437), .B(new_n438), .C1(G134), .C2(new_n430), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n433), .A2(new_n439), .ZN(new_n440));
  XNOR2_X1  g254(.A(KEYINPUT9), .B(G234), .ZN(new_n441));
  NOR3_X1   g255(.A1(new_n342), .A2(new_n441), .A3(G953), .ZN(new_n442));
  INV_X1    g256(.A(new_n442), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n440), .A2(new_n443), .ZN(new_n444));
  NAND3_X1  g258(.A1(new_n433), .A2(new_n439), .A3(new_n442), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n444), .A2(new_n445), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n446), .A2(new_n333), .ZN(new_n447));
  INV_X1    g261(.A(G478), .ZN(new_n448));
  NOR2_X1   g262(.A1(new_n448), .A2(KEYINPUT15), .ZN(new_n449));
  AND2_X1   g263(.A1(new_n447), .A2(new_n449), .ZN(new_n450));
  NOR2_X1   g264(.A1(new_n447), .A2(new_n449), .ZN(new_n451));
  NOR2_X1   g265(.A1(new_n450), .A2(new_n451), .ZN(new_n452));
  NAND3_X1  g266(.A1(new_n416), .A2(new_n422), .A3(new_n452), .ZN(new_n453));
  INV_X1    g267(.A(new_n453), .ZN(new_n454));
  INV_X1    g268(.A(G469), .ZN(new_n455));
  XNOR2_X1  g269(.A(G110), .B(G140), .ZN(new_n456));
  XNOR2_X1  g270(.A(new_n456), .B(KEYINPUT76), .ZN(new_n457));
  INV_X1    g271(.A(G227), .ZN(new_n458));
  NOR2_X1   g272(.A1(new_n458), .A2(G953), .ZN(new_n459));
  XOR2_X1   g273(.A(new_n457), .B(new_n459), .Z(new_n460));
  NAND2_X1  g274(.A1(new_n423), .A2(G104), .ZN(new_n461));
  AND2_X1   g275(.A1(KEYINPUT77), .A2(KEYINPUT3), .ZN(new_n462));
  NOR2_X1   g276(.A1(KEYINPUT77), .A2(KEYINPUT3), .ZN(new_n463));
  OAI21_X1  g277(.A(new_n461), .B1(new_n462), .B2(new_n463), .ZN(new_n464));
  INV_X1    g278(.A(G101), .ZN(new_n465));
  NAND2_X1  g279(.A1(new_n374), .A2(G107), .ZN(new_n466));
  NAND2_X1  g280(.A1(KEYINPUT77), .A2(KEYINPUT3), .ZN(new_n467));
  NAND3_X1  g281(.A1(new_n467), .A2(G104), .A3(new_n423), .ZN(new_n468));
  NAND4_X1  g282(.A1(new_n464), .A2(new_n465), .A3(new_n466), .A4(new_n468), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n466), .A2(new_n461), .ZN(new_n470));
  NAND2_X1  g284(.A1(new_n470), .A2(G101), .ZN(new_n471));
  AND2_X1   g285(.A1(new_n469), .A2(new_n471), .ZN(new_n472));
  NOR2_X1   g286(.A1(new_n216), .A2(KEYINPUT80), .ZN(new_n473));
  INV_X1    g287(.A(new_n473), .ZN(new_n474));
  AOI21_X1  g288(.A(new_n217), .B1(new_n216), .B2(KEYINPUT80), .ZN(new_n475));
  AOI21_X1  g289(.A(new_n219), .B1(new_n474), .B2(new_n475), .ZN(new_n476));
  INV_X1    g290(.A(KEYINPUT79), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n221), .A2(new_n477), .ZN(new_n478));
  NAND3_X1  g292(.A1(new_n219), .A2(KEYINPUT79), .A3(new_n220), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n478), .A2(new_n479), .ZN(new_n480));
  OAI21_X1  g294(.A(new_n472), .B1(new_n476), .B2(new_n480), .ZN(new_n481));
  OAI21_X1  g295(.A(new_n481), .B1(new_n222), .B2(new_n472), .ZN(new_n482));
  INV_X1    g296(.A(KEYINPUT12), .ZN(new_n483));
  NAND4_X1  g297(.A1(new_n482), .A2(KEYINPUT81), .A3(new_n483), .A4(new_n227), .ZN(new_n484));
  OR2_X1    g298(.A1(new_n483), .A2(KEYINPUT81), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n483), .A2(KEYINPUT81), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n469), .A2(new_n471), .ZN(new_n487));
  AND3_X1   g301(.A1(new_n219), .A2(KEYINPUT79), .A3(new_n220), .ZN(new_n488));
  AOI21_X1  g302(.A(KEYINPUT79), .B1(new_n219), .B2(new_n220), .ZN(new_n489));
  NOR2_X1   g303(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  NAND2_X1  g304(.A1(new_n211), .A2(KEYINPUT1), .ZN(new_n491));
  INV_X1    g305(.A(KEYINPUT80), .ZN(new_n492));
  OAI21_X1  g306(.A(G128), .B1(new_n491), .B2(new_n492), .ZN(new_n493));
  OAI21_X1  g307(.A(new_n214), .B1(new_n493), .B2(new_n473), .ZN(new_n494));
  AOI21_X1  g308(.A(new_n487), .B1(new_n490), .B2(new_n494), .ZN(new_n495));
  AOI21_X1  g309(.A(new_n222), .B1(new_n471), .B2(new_n469), .ZN(new_n496));
  NOR2_X1   g310(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  OAI211_X1 g311(.A(new_n485), .B(new_n486), .C1(new_n497), .C2(new_n234), .ZN(new_n498));
  INV_X1    g312(.A(KEYINPUT78), .ZN(new_n499));
  OR2_X1    g313(.A1(KEYINPUT77), .A2(KEYINPUT3), .ZN(new_n500));
  AOI22_X1  g314(.A1(new_n500), .A2(new_n467), .B1(G104), .B2(new_n423), .ZN(new_n501));
  NAND2_X1  g315(.A1(new_n468), .A2(new_n466), .ZN(new_n502));
  OAI21_X1  g316(.A(new_n499), .B1(new_n501), .B2(new_n502), .ZN(new_n503));
  NAND4_X1  g317(.A1(new_n464), .A2(KEYINPUT78), .A3(new_n466), .A4(new_n468), .ZN(new_n504));
  NAND3_X1  g318(.A1(new_n503), .A2(G101), .A3(new_n504), .ZN(new_n505));
  AND2_X1   g319(.A1(new_n469), .A2(KEYINPUT4), .ZN(new_n506));
  NAND2_X1  g320(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  INV_X1    g321(.A(KEYINPUT4), .ZN(new_n508));
  NAND4_X1  g322(.A1(new_n503), .A2(new_n508), .A3(G101), .A4(new_n504), .ZN(new_n509));
  NAND3_X1  g323(.A1(new_n241), .A2(new_n507), .A3(new_n509), .ZN(new_n510));
  INV_X1    g324(.A(KEYINPUT10), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n481), .A2(new_n511), .ZN(new_n512));
  AOI21_X1  g326(.A(new_n511), .B1(new_n218), .B2(new_n221), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n472), .A2(new_n513), .ZN(new_n514));
  NAND4_X1  g328(.A1(new_n510), .A2(new_n234), .A3(new_n512), .A4(new_n514), .ZN(new_n515));
  AND4_X1   g329(.A1(new_n460), .A2(new_n484), .A3(new_n498), .A4(new_n515), .ZN(new_n516));
  AND3_X1   g330(.A1(new_n241), .A2(new_n507), .A3(new_n509), .ZN(new_n517));
  OAI21_X1  g331(.A(new_n514), .B1(new_n495), .B2(KEYINPUT10), .ZN(new_n518));
  OAI21_X1  g332(.A(new_n227), .B1(new_n517), .B2(new_n518), .ZN(new_n519));
  AOI21_X1  g333(.A(new_n460), .B1(new_n519), .B2(new_n515), .ZN(new_n520));
  OAI211_X1 g334(.A(new_n455), .B(new_n333), .C1(new_n516), .C2(new_n520), .ZN(new_n521));
  NAND3_X1  g335(.A1(new_n484), .A2(new_n498), .A3(new_n515), .ZN(new_n522));
  INV_X1    g336(.A(new_n460), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  NAND3_X1  g338(.A1(new_n519), .A2(new_n460), .A3(new_n515), .ZN(new_n525));
  NAND3_X1  g339(.A1(new_n524), .A2(G469), .A3(new_n525), .ZN(new_n526));
  NOR2_X1   g340(.A1(new_n455), .A2(new_n333), .ZN(new_n527));
  INV_X1    g341(.A(new_n527), .ZN(new_n528));
  NAND3_X1  g342(.A1(new_n521), .A2(new_n526), .A3(new_n528), .ZN(new_n529));
  OAI21_X1  g343(.A(G221), .B1(new_n441), .B2(G902), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  NAND2_X1  g345(.A1(G234), .A2(G237), .ZN(new_n532));
  NAND3_X1  g346(.A1(new_n532), .A2(G952), .A3(new_n329), .ZN(new_n533));
  XNOR2_X1  g347(.A(new_n533), .B(KEYINPUT93), .ZN(new_n534));
  NAND2_X1  g348(.A1(new_n532), .A2(G902), .ZN(new_n535));
  INV_X1    g349(.A(G898), .ZN(new_n536));
  AOI21_X1  g350(.A(new_n329), .B1(KEYINPUT21), .B2(new_n536), .ZN(new_n537));
  OAI21_X1  g351(.A(new_n537), .B1(KEYINPUT21), .B2(new_n536), .ZN(new_n538));
  OAI21_X1  g352(.A(new_n534), .B1(new_n535), .B2(new_n538), .ZN(new_n539));
  XOR2_X1   g353(.A(new_n539), .B(KEYINPUT94), .Z(new_n540));
  OAI21_X1  g354(.A(G214), .B1(G237), .B2(G902), .ZN(new_n541));
  INV_X1    g355(.A(KEYINPUT5), .ZN(new_n542));
  NOR2_X1   g356(.A1(new_n249), .A2(new_n542), .ZN(new_n543));
  NAND3_X1  g357(.A1(new_n542), .A2(new_n304), .A3(G116), .ZN(new_n544));
  NAND2_X1  g358(.A1(new_n544), .A2(G113), .ZN(new_n545));
  OAI22_X1  g359(.A1(new_n543), .A2(new_n545), .B1(new_n249), .B2(new_n250), .ZN(new_n546));
  OR2_X1    g360(.A1(new_n546), .A2(new_n487), .ZN(new_n547));
  AND2_X1   g361(.A1(new_n505), .A2(new_n506), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n509), .A2(new_n251), .ZN(new_n549));
  OAI21_X1  g363(.A(new_n547), .B1(new_n548), .B2(new_n549), .ZN(new_n550));
  XNOR2_X1  g364(.A(G110), .B(G122), .ZN(new_n551));
  INV_X1    g365(.A(new_n551), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n550), .A2(new_n552), .ZN(new_n553));
  OAI211_X1 g367(.A(new_n547), .B(new_n551), .C1(new_n548), .C2(new_n549), .ZN(new_n554));
  NAND3_X1  g368(.A1(new_n553), .A2(KEYINPUT6), .A3(new_n554), .ZN(new_n555));
  XNOR2_X1  g369(.A(KEYINPUT83), .B(G224), .ZN(new_n556));
  NOR2_X1   g370(.A1(new_n556), .A2(G953), .ZN(new_n557));
  INV_X1    g371(.A(KEYINPUT84), .ZN(new_n558));
  XNOR2_X1  g372(.A(new_n557), .B(new_n558), .ZN(new_n559));
  XNOR2_X1  g373(.A(new_n559), .B(KEYINPUT85), .ZN(new_n560));
  OAI211_X1 g374(.A(new_n230), .B(G125), .C1(new_n231), .C2(new_n219), .ZN(new_n561));
  OAI21_X1  g375(.A(new_n561), .B1(new_n222), .B2(G125), .ZN(new_n562));
  INV_X1    g376(.A(KEYINPUT82), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n561), .A2(KEYINPUT82), .ZN(new_n565));
  NAND3_X1  g379(.A1(new_n560), .A2(new_n564), .A3(new_n565), .ZN(new_n566));
  XNOR2_X1  g380(.A(new_n557), .B(KEYINPUT84), .ZN(new_n567));
  XNOR2_X1  g381(.A(new_n567), .B(KEYINPUT85), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n564), .A2(new_n565), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n568), .A2(new_n569), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n566), .A2(new_n570), .ZN(new_n571));
  INV_X1    g385(.A(KEYINPUT6), .ZN(new_n572));
  NAND3_X1  g386(.A1(new_n550), .A2(new_n572), .A3(new_n552), .ZN(new_n573));
  NAND3_X1  g387(.A1(new_n555), .A2(new_n571), .A3(new_n573), .ZN(new_n574));
  INV_X1    g388(.A(KEYINPUT7), .ZN(new_n575));
  NOR2_X1   g389(.A1(new_n567), .A2(new_n575), .ZN(new_n576));
  AND3_X1   g390(.A1(new_n576), .A2(new_n564), .A3(new_n565), .ZN(new_n577));
  XOR2_X1   g391(.A(new_n551), .B(KEYINPUT8), .Z(new_n578));
  NAND2_X1  g392(.A1(new_n546), .A2(new_n487), .ZN(new_n579));
  AOI21_X1  g393(.A(new_n578), .B1(new_n547), .B2(new_n579), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n559), .A2(KEYINPUT7), .ZN(new_n581));
  AND2_X1   g395(.A1(new_n581), .A2(new_n562), .ZN(new_n582));
  NOR3_X1   g396(.A1(new_n577), .A2(new_n580), .A3(new_n582), .ZN(new_n583));
  AOI21_X1  g397(.A(G902), .B1(new_n583), .B2(new_n554), .ZN(new_n584));
  OAI21_X1  g398(.A(G210), .B1(G237), .B2(G902), .ZN(new_n585));
  AND3_X1   g399(.A1(new_n574), .A2(new_n584), .A3(new_n585), .ZN(new_n586));
  AOI21_X1  g400(.A(new_n585), .B1(new_n574), .B2(new_n584), .ZN(new_n587));
  OAI211_X1 g401(.A(new_n540), .B(new_n541), .C1(new_n586), .C2(new_n587), .ZN(new_n588));
  NOR2_X1   g402(.A1(new_n531), .A2(new_n588), .ZN(new_n589));
  NAND3_X1  g403(.A1(new_n454), .A2(new_n589), .A3(KEYINPUT95), .ZN(new_n590));
  INV_X1    g404(.A(KEYINPUT95), .ZN(new_n591));
  INV_X1    g405(.A(new_n541), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n574), .A2(new_n584), .ZN(new_n593));
  INV_X1    g407(.A(new_n585), .ZN(new_n594));
  NAND2_X1  g408(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  NAND3_X1  g409(.A1(new_n574), .A2(new_n584), .A3(new_n585), .ZN(new_n596));
  AOI21_X1  g410(.A(new_n592), .B1(new_n595), .B2(new_n596), .ZN(new_n597));
  NAND4_X1  g411(.A1(new_n597), .A2(new_n540), .A3(new_n530), .A4(new_n529), .ZN(new_n598));
  OAI21_X1  g412(.A(new_n591), .B1(new_n598), .B2(new_n453), .ZN(new_n599));
  NAND4_X1  g413(.A1(new_n302), .A2(new_n354), .A3(new_n590), .A4(new_n599), .ZN(new_n600));
  XNOR2_X1  g414(.A(new_n600), .B(G101), .ZN(G3));
  NAND2_X1  g415(.A1(new_n276), .A2(new_n333), .ZN(new_n602));
  AOI22_X1  g416(.A1(new_n602), .A2(G472), .B1(new_n277), .B2(new_n276), .ZN(new_n603));
  NOR2_X1   g417(.A1(new_n353), .A2(new_n531), .ZN(new_n604));
  AND2_X1   g418(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  AOI22_X1  g419(.A1(new_n444), .A2(new_n445), .B1(KEYINPUT96), .B2(KEYINPUT33), .ZN(new_n606));
  INV_X1    g420(.A(new_n446), .ZN(new_n607));
  XNOR2_X1  g421(.A(KEYINPUT96), .B(KEYINPUT33), .ZN(new_n608));
  AOI21_X1  g422(.A(new_n606), .B1(new_n607), .B2(new_n608), .ZN(new_n609));
  NOR2_X1   g423(.A1(new_n448), .A2(G902), .ZN(new_n610));
  AOI22_X1  g424(.A1(new_n609), .A2(new_n610), .B1(new_n448), .B2(new_n447), .ZN(new_n611));
  AOI21_X1  g425(.A(new_n611), .B1(new_n416), .B2(new_n422), .ZN(new_n612));
  INV_X1    g426(.A(new_n612), .ZN(new_n613));
  NOR2_X1   g427(.A1(new_n613), .A2(new_n588), .ZN(new_n614));
  NAND2_X1  g428(.A1(new_n605), .A2(new_n614), .ZN(new_n615));
  XNOR2_X1  g429(.A(new_n615), .B(KEYINPUT97), .ZN(new_n616));
  XOR2_X1   g430(.A(KEYINPUT34), .B(G104), .Z(new_n617));
  XNOR2_X1  g431(.A(new_n616), .B(new_n617), .ZN(G6));
  INV_X1    g432(.A(new_n452), .ZN(new_n619));
  XNOR2_X1  g433(.A(new_n407), .B(new_n410), .ZN(new_n620));
  AND2_X1   g434(.A1(new_n620), .A2(new_n395), .ZN(new_n621));
  XOR2_X1   g435(.A(new_n540), .B(KEYINPUT98), .Z(new_n622));
  AND4_X1   g436(.A1(new_n619), .A2(new_n597), .A3(new_n621), .A4(new_n622), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n605), .A2(new_n623), .ZN(new_n624));
  XOR2_X1   g438(.A(KEYINPUT35), .B(G107), .Z(new_n625));
  XNOR2_X1  g439(.A(new_n624), .B(new_n625), .ZN(G9));
  NOR2_X1   g440(.A1(new_n323), .A2(new_n327), .ZN(new_n627));
  NOR2_X1   g441(.A1(new_n331), .A2(KEYINPUT36), .ZN(new_n628));
  XOR2_X1   g442(.A(new_n627), .B(new_n628), .Z(new_n629));
  NAND2_X1  g443(.A1(new_n629), .A2(new_n351), .ZN(new_n630));
  OAI21_X1  g444(.A(new_n630), .B1(new_n344), .B2(new_n348), .ZN(new_n631));
  NAND4_X1  g445(.A1(new_n603), .A2(new_n599), .A3(new_n590), .A4(new_n631), .ZN(new_n632));
  XOR2_X1   g446(.A(KEYINPUT37), .B(G110), .Z(new_n633));
  XNOR2_X1  g447(.A(new_n632), .B(new_n633), .ZN(G12));
  INV_X1    g448(.A(new_n631), .ZN(new_n635));
  OAI21_X1  g449(.A(new_n541), .B1(new_n586), .B2(new_n587), .ZN(new_n636));
  NOR3_X1   g450(.A1(new_n635), .A2(new_n636), .A3(new_n531), .ZN(new_n637));
  NAND2_X1  g451(.A1(new_n297), .A2(new_n281), .ZN(new_n638));
  AOI21_X1  g452(.A(KEYINPUT32), .B1(new_n276), .B2(new_n277), .ZN(new_n639));
  OAI21_X1  g453(.A(new_n637), .B1(new_n638), .B2(new_n639), .ZN(new_n640));
  NOR3_X1   g454(.A1(new_n535), .A2(G900), .A3(new_n329), .ZN(new_n641));
  XOR2_X1   g455(.A(new_n641), .B(KEYINPUT99), .Z(new_n642));
  NAND2_X1  g456(.A1(new_n642), .A2(new_n534), .ZN(new_n643));
  XNOR2_X1  g457(.A(new_n643), .B(KEYINPUT100), .ZN(new_n644));
  INV_X1    g458(.A(new_n644), .ZN(new_n645));
  NAND3_X1  g459(.A1(new_n619), .A2(new_n621), .A3(new_n645), .ZN(new_n646));
  NOR2_X1   g460(.A1(new_n640), .A2(new_n646), .ZN(new_n647));
  XNOR2_X1  g461(.A(new_n647), .B(new_n217), .ZN(G30));
  XOR2_X1   g462(.A(new_n644), .B(KEYINPUT39), .Z(new_n649));
  INV_X1    g463(.A(new_n649), .ZN(new_n650));
  NOR2_X1   g464(.A1(new_n531), .A2(new_n650), .ZN(new_n651));
  XNOR2_X1  g465(.A(new_n651), .B(KEYINPUT40), .ZN(new_n652));
  OR2_X1    g466(.A1(new_n652), .A2(KEYINPUT101), .ZN(new_n653));
  NAND2_X1  g467(.A1(new_n652), .A2(KEYINPUT101), .ZN(new_n654));
  AOI21_X1  g468(.A(new_n259), .B1(new_n283), .B2(new_n285), .ZN(new_n655));
  NOR3_X1   g469(.A1(new_n298), .A2(new_n299), .A3(new_n655), .ZN(new_n656));
  OAI21_X1  g470(.A(new_n279), .B1(new_n656), .B2(new_n278), .ZN(new_n657));
  NOR2_X1   g471(.A1(new_n273), .A2(new_n262), .ZN(new_n658));
  NAND3_X1  g472(.A1(new_n291), .A2(new_n254), .A3(new_n262), .ZN(new_n659));
  NAND2_X1  g473(.A1(new_n659), .A2(new_n333), .ZN(new_n660));
  OAI21_X1  g474(.A(G472), .B1(new_n658), .B2(new_n660), .ZN(new_n661));
  NAND3_X1  g475(.A1(new_n657), .A2(new_n281), .A3(new_n661), .ZN(new_n662));
  NOR2_X1   g476(.A1(new_n586), .A2(new_n587), .ZN(new_n663));
  XOR2_X1   g477(.A(new_n663), .B(KEYINPUT38), .Z(new_n664));
  AOI21_X1  g478(.A(new_n452), .B1(new_n416), .B2(new_n422), .ZN(new_n665));
  AND4_X1   g479(.A1(new_n541), .A2(new_n664), .A3(new_n635), .A4(new_n665), .ZN(new_n666));
  NAND4_X1  g480(.A1(new_n653), .A2(new_n654), .A3(new_n662), .A4(new_n666), .ZN(new_n667));
  XNOR2_X1  g481(.A(new_n667), .B(G143), .ZN(G45));
  INV_X1    g482(.A(KEYINPUT103), .ZN(new_n669));
  INV_X1    g483(.A(new_n611), .ZN(new_n670));
  NOR2_X1   g484(.A1(new_n414), .A2(new_n415), .ZN(new_n671));
  AOI21_X1  g485(.A(KEYINPUT90), .B1(new_n421), .B2(new_n395), .ZN(new_n672));
  OAI211_X1 g486(.A(new_n670), .B(new_n645), .C1(new_n671), .C2(new_n672), .ZN(new_n673));
  NAND2_X1  g487(.A1(new_n673), .A2(KEYINPUT102), .ZN(new_n674));
  INV_X1    g488(.A(KEYINPUT102), .ZN(new_n675));
  NAND3_X1  g489(.A1(new_n612), .A2(new_n675), .A3(new_n645), .ZN(new_n676));
  NAND2_X1  g490(.A1(new_n674), .A2(new_n676), .ZN(new_n677));
  OAI21_X1  g491(.A(new_n669), .B1(new_n640), .B2(new_n677), .ZN(new_n678));
  NOR2_X1   g492(.A1(new_n673), .A2(KEYINPUT102), .ZN(new_n679));
  AOI21_X1  g493(.A(new_n675), .B1(new_n612), .B2(new_n645), .ZN(new_n680));
  NOR2_X1   g494(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  AND2_X1   g495(.A1(new_n529), .A2(new_n530), .ZN(new_n682));
  NAND3_X1  g496(.A1(new_n682), .A2(new_n597), .A3(new_n631), .ZN(new_n683));
  AOI22_X1  g497(.A1(G472), .A2(new_n296), .B1(new_n276), .B2(new_n280), .ZN(new_n684));
  AOI21_X1  g498(.A(new_n683), .B1(new_n684), .B2(new_n657), .ZN(new_n685));
  NAND3_X1  g499(.A1(new_n681), .A2(new_n685), .A3(KEYINPUT103), .ZN(new_n686));
  NAND2_X1  g500(.A1(new_n678), .A2(new_n686), .ZN(new_n687));
  XNOR2_X1  g501(.A(new_n687), .B(G146), .ZN(G48));
  AOI21_X1  g502(.A(new_n353), .B1(new_n684), .B2(new_n657), .ZN(new_n689));
  NAND2_X1  g503(.A1(new_n519), .A2(new_n515), .ZN(new_n690));
  NAND2_X1  g504(.A1(new_n690), .A2(new_n523), .ZN(new_n691));
  NAND4_X1  g505(.A1(new_n484), .A2(new_n498), .A3(new_n515), .A4(new_n460), .ZN(new_n692));
  NAND2_X1  g506(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  AOI21_X1  g507(.A(new_n455), .B1(new_n693), .B2(new_n333), .ZN(new_n694));
  INV_X1    g508(.A(new_n521), .ZN(new_n695));
  OR2_X1    g509(.A1(new_n694), .A2(new_n695), .ZN(new_n696));
  INV_X1    g510(.A(new_n530), .ZN(new_n697));
  NOR2_X1   g511(.A1(new_n696), .A2(new_n697), .ZN(new_n698));
  NAND3_X1  g512(.A1(new_n689), .A2(new_n614), .A3(new_n698), .ZN(new_n699));
  XNOR2_X1  g513(.A(KEYINPUT41), .B(G113), .ZN(new_n700));
  XNOR2_X1  g514(.A(new_n699), .B(new_n700), .ZN(G15));
  NAND4_X1  g515(.A1(new_n302), .A2(new_n354), .A3(new_n623), .A4(new_n698), .ZN(new_n702));
  XNOR2_X1  g516(.A(new_n702), .B(G116), .ZN(G18));
  NOR2_X1   g517(.A1(new_n694), .A2(new_n695), .ZN(new_n704));
  NAND4_X1  g518(.A1(new_n631), .A2(new_n704), .A3(new_n597), .A4(new_n530), .ZN(new_n705));
  INV_X1    g519(.A(new_n705), .ZN(new_n706));
  NAND4_X1  g520(.A1(new_n302), .A2(new_n454), .A3(new_n540), .A4(new_n706), .ZN(new_n707));
  XNOR2_X1  g521(.A(new_n707), .B(G119), .ZN(G21));
  OAI21_X1  g522(.A(new_n262), .B1(new_n267), .B2(new_n292), .ZN(new_n709));
  AOI21_X1  g523(.A(new_n278), .B1(new_n300), .B2(new_n709), .ZN(new_n710));
  INV_X1    g524(.A(new_n710), .ZN(new_n711));
  AOI21_X1  g525(.A(KEYINPUT104), .B1(new_n602), .B2(G472), .ZN(new_n712));
  INV_X1    g526(.A(KEYINPUT104), .ZN(new_n713));
  INV_X1    g527(.A(G472), .ZN(new_n714));
  AOI211_X1 g528(.A(new_n713), .B(new_n714), .C1(new_n276), .C2(new_n333), .ZN(new_n715));
  OAI211_X1 g529(.A(new_n354), .B(new_n711), .C1(new_n712), .C2(new_n715), .ZN(new_n716));
  NAND2_X1  g530(.A1(new_n597), .A2(new_n622), .ZN(new_n717));
  INV_X1    g531(.A(new_n717), .ZN(new_n718));
  NOR2_X1   g532(.A1(new_n665), .A2(KEYINPUT105), .ZN(new_n719));
  INV_X1    g533(.A(KEYINPUT105), .ZN(new_n720));
  AOI211_X1 g534(.A(new_n720), .B(new_n452), .C1(new_n416), .C2(new_n422), .ZN(new_n721));
  OAI211_X1 g535(.A(new_n698), .B(new_n718), .C1(new_n719), .C2(new_n721), .ZN(new_n722));
  NOR2_X1   g536(.A1(new_n716), .A2(new_n722), .ZN(new_n723));
  XNOR2_X1  g537(.A(new_n723), .B(new_n424), .ZN(G24));
  AND3_X1   g538(.A1(new_n674), .A2(KEYINPUT106), .A3(new_n676), .ZN(new_n725));
  AOI21_X1  g539(.A(KEYINPUT106), .B1(new_n674), .B2(new_n676), .ZN(new_n726));
  NOR2_X1   g540(.A1(new_n725), .A2(new_n726), .ZN(new_n727));
  AOI21_X1  g541(.A(G902), .B1(new_n300), .B2(new_n271), .ZN(new_n728));
  OAI21_X1  g542(.A(new_n713), .B1(new_n728), .B2(new_n714), .ZN(new_n729));
  NAND3_X1  g543(.A1(new_n602), .A2(KEYINPUT104), .A3(G472), .ZN(new_n730));
  AOI211_X1 g544(.A(new_n705), .B(new_n710), .C1(new_n729), .C2(new_n730), .ZN(new_n731));
  NAND2_X1  g545(.A1(new_n727), .A2(new_n731), .ZN(new_n732));
  XOR2_X1   g546(.A(KEYINPUT107), .B(G125), .Z(new_n733));
  XNOR2_X1  g547(.A(new_n732), .B(new_n733), .ZN(G27));
  NAND2_X1  g548(.A1(new_n663), .A2(new_n541), .ZN(new_n735));
  NOR2_X1   g549(.A1(new_n735), .A2(new_n531), .ZN(new_n736));
  INV_X1    g550(.A(KEYINPUT108), .ZN(new_n737));
  NOR2_X1   g551(.A1(new_n737), .A2(KEYINPUT42), .ZN(new_n738));
  INV_X1    g552(.A(new_n738), .ZN(new_n739));
  NAND4_X1  g553(.A1(new_n302), .A2(new_n354), .A3(new_n736), .A4(new_n739), .ZN(new_n740));
  INV_X1    g554(.A(new_n740), .ZN(new_n741));
  NAND2_X1  g555(.A1(new_n737), .A2(KEYINPUT42), .ZN(new_n742));
  NAND3_X1  g556(.A1(new_n741), .A2(new_n727), .A3(new_n742), .ZN(new_n743));
  INV_X1    g557(.A(new_n742), .ZN(new_n744));
  INV_X1    g558(.A(KEYINPUT106), .ZN(new_n745));
  OAI21_X1  g559(.A(new_n745), .B1(new_n679), .B2(new_n680), .ZN(new_n746));
  NAND3_X1  g560(.A1(new_n674), .A2(KEYINPUT106), .A3(new_n676), .ZN(new_n747));
  NAND2_X1  g561(.A1(new_n746), .A2(new_n747), .ZN(new_n748));
  OAI21_X1  g562(.A(new_n744), .B1(new_n748), .B2(new_n740), .ZN(new_n749));
  NAND2_X1  g563(.A1(new_n743), .A2(new_n749), .ZN(new_n750));
  XNOR2_X1  g564(.A(KEYINPUT109), .B(G131), .ZN(new_n751));
  XNOR2_X1  g565(.A(new_n750), .B(new_n751), .ZN(G33));
  OAI211_X1 g566(.A(new_n354), .B(new_n736), .C1(new_n638), .C2(new_n639), .ZN(new_n753));
  OAI21_X1  g567(.A(KEYINPUT110), .B1(new_n753), .B2(new_n646), .ZN(new_n754));
  INV_X1    g568(.A(KEYINPUT110), .ZN(new_n755));
  INV_X1    g569(.A(new_n646), .ZN(new_n756));
  NAND4_X1  g570(.A1(new_n689), .A2(new_n755), .A3(new_n756), .A4(new_n736), .ZN(new_n757));
  NAND2_X1  g571(.A1(new_n754), .A2(new_n757), .ZN(new_n758));
  XNOR2_X1  g572(.A(new_n758), .B(G134), .ZN(G36));
  NOR2_X1   g573(.A1(new_n671), .A2(new_n672), .ZN(new_n760));
  NAND2_X1  g574(.A1(new_n760), .A2(new_n670), .ZN(new_n761));
  OR2_X1    g575(.A1(new_n761), .A2(KEYINPUT43), .ZN(new_n762));
  NAND2_X1  g576(.A1(new_n761), .A2(KEYINPUT43), .ZN(new_n763));
  NAND2_X1  g577(.A1(new_n762), .A2(new_n763), .ZN(new_n764));
  OR2_X1    g578(.A1(new_n764), .A2(KEYINPUT111), .ZN(new_n765));
  NAND2_X1  g579(.A1(new_n764), .A2(KEYINPUT111), .ZN(new_n766));
  NOR2_X1   g580(.A1(new_n603), .A2(new_n635), .ZN(new_n767));
  NAND3_X1  g581(.A1(new_n765), .A2(new_n766), .A3(new_n767), .ZN(new_n768));
  INV_X1    g582(.A(KEYINPUT44), .ZN(new_n769));
  NAND2_X1  g583(.A1(new_n768), .A2(new_n769), .ZN(new_n770));
  NAND4_X1  g584(.A1(new_n765), .A2(KEYINPUT44), .A3(new_n766), .A4(new_n767), .ZN(new_n771));
  NAND2_X1  g585(.A1(new_n524), .A2(new_n525), .ZN(new_n772));
  INV_X1    g586(.A(KEYINPUT45), .ZN(new_n773));
  NOR2_X1   g587(.A1(new_n772), .A2(new_n773), .ZN(new_n774));
  AOI21_X1  g588(.A(KEYINPUT45), .B1(new_n524), .B2(new_n525), .ZN(new_n775));
  NOR3_X1   g589(.A1(new_n774), .A2(new_n455), .A3(new_n775), .ZN(new_n776));
  NOR2_X1   g590(.A1(new_n776), .A2(new_n527), .ZN(new_n777));
  AND2_X1   g591(.A1(new_n777), .A2(KEYINPUT46), .ZN(new_n778));
  OAI21_X1  g592(.A(new_n521), .B1(new_n777), .B2(KEYINPUT46), .ZN(new_n779));
  OAI21_X1  g593(.A(new_n530), .B1(new_n778), .B2(new_n779), .ZN(new_n780));
  OR2_X1    g594(.A1(new_n780), .A2(new_n650), .ZN(new_n781));
  XOR2_X1   g595(.A(new_n735), .B(KEYINPUT112), .Z(new_n782));
  NOR2_X1   g596(.A1(new_n781), .A2(new_n782), .ZN(new_n783));
  NAND3_X1  g597(.A1(new_n770), .A2(new_n771), .A3(new_n783), .ZN(new_n784));
  XNOR2_X1  g598(.A(new_n784), .B(G137), .ZN(G39));
  XNOR2_X1  g599(.A(new_n780), .B(KEYINPUT47), .ZN(new_n786));
  INV_X1    g600(.A(new_n786), .ZN(new_n787));
  NOR4_X1   g601(.A1(new_n677), .A2(new_n302), .A3(new_n354), .A4(new_n735), .ZN(new_n788));
  NAND2_X1  g602(.A1(new_n787), .A2(new_n788), .ZN(new_n789));
  XNOR2_X1  g603(.A(new_n789), .B(G140), .ZN(G42));
  INV_X1    g604(.A(KEYINPUT115), .ZN(new_n791));
  NOR3_X1   g605(.A1(new_n631), .A2(new_n531), .A3(new_n644), .ZN(new_n792));
  NAND2_X1  g606(.A1(new_n281), .A2(new_n661), .ZN(new_n793));
  OAI21_X1  g607(.A(new_n792), .B1(new_n793), .B2(new_n639), .ZN(new_n794));
  OAI21_X1  g608(.A(new_n597), .B1(new_n719), .B2(new_n721), .ZN(new_n795));
  NOR2_X1   g609(.A1(new_n794), .A2(new_n795), .ZN(new_n796));
  AOI21_X1  g610(.A(new_n796), .B1(new_n727), .B2(new_n731), .ZN(new_n797));
  AOI21_X1  g611(.A(new_n647), .B1(new_n678), .B2(new_n686), .ZN(new_n798));
  AND3_X1   g612(.A1(new_n797), .A2(new_n798), .A3(KEYINPUT52), .ZN(new_n799));
  AOI21_X1  g613(.A(KEYINPUT52), .B1(new_n797), .B2(new_n798), .ZN(new_n800));
  NOR2_X1   g614(.A1(new_n799), .A2(new_n800), .ZN(new_n801));
  AND3_X1   g615(.A1(new_n743), .A2(new_n758), .A3(new_n749), .ZN(new_n802));
  NOR2_X1   g616(.A1(new_n638), .A2(new_n639), .ZN(new_n803));
  NAND3_X1  g617(.A1(new_n621), .A2(new_n452), .A3(new_n645), .ZN(new_n804));
  NOR2_X1   g618(.A1(new_n735), .A2(new_n804), .ZN(new_n805));
  NAND3_X1  g619(.A1(new_n805), .A2(new_n682), .A3(new_n631), .ZN(new_n806));
  OR2_X1    g620(.A1(new_n803), .A2(new_n806), .ZN(new_n807));
  NAND3_X1  g621(.A1(new_n746), .A2(new_n747), .A3(new_n736), .ZN(new_n808));
  OAI211_X1 g622(.A(new_n631), .B(new_n711), .C1(new_n712), .C2(new_n715), .ZN(new_n809));
  OAI21_X1  g623(.A(new_n807), .B1(new_n808), .B2(new_n809), .ZN(new_n810));
  INV_X1    g624(.A(KEYINPUT113), .ZN(new_n811));
  NAND2_X1  g625(.A1(new_n416), .A2(new_n422), .ZN(new_n812));
  OAI21_X1  g626(.A(new_n811), .B1(new_n812), .B2(new_n452), .ZN(new_n813));
  NAND4_X1  g627(.A1(new_n416), .A2(new_n619), .A3(KEYINPUT113), .A4(new_n422), .ZN(new_n814));
  NAND3_X1  g628(.A1(new_n813), .A2(new_n613), .A3(new_n814), .ZN(new_n815));
  NAND4_X1  g629(.A1(new_n815), .A2(new_n603), .A3(new_n604), .A4(new_n718), .ZN(new_n816));
  NAND4_X1  g630(.A1(new_n699), .A2(new_n632), .A3(new_n702), .A4(new_n816), .ZN(new_n817));
  OAI211_X1 g631(.A(new_n600), .B(new_n707), .C1(new_n716), .C2(new_n722), .ZN(new_n818));
  NOR3_X1   g632(.A1(new_n810), .A2(new_n817), .A3(new_n818), .ZN(new_n819));
  NAND3_X1  g633(.A1(new_n802), .A2(new_n819), .A3(KEYINPUT53), .ZN(new_n820));
  OAI21_X1  g634(.A(new_n791), .B1(new_n801), .B2(new_n820), .ZN(new_n821));
  NOR2_X1   g635(.A1(new_n817), .A2(new_n818), .ZN(new_n822));
  INV_X1    g636(.A(new_n810), .ZN(new_n823));
  NAND2_X1  g637(.A1(new_n822), .A2(new_n823), .ZN(new_n824));
  NAND3_X1  g638(.A1(new_n743), .A2(new_n758), .A3(new_n749), .ZN(new_n825));
  NOR2_X1   g639(.A1(new_n824), .A2(new_n825), .ZN(new_n826));
  INV_X1    g640(.A(KEYINPUT52), .ZN(new_n827));
  INV_X1    g641(.A(new_n647), .ZN(new_n828));
  NAND2_X1  g642(.A1(new_n687), .A2(new_n828), .ZN(new_n829));
  OAI211_X1 g643(.A(new_n706), .B(new_n711), .C1(new_n712), .C2(new_n715), .ZN(new_n830));
  OAI22_X1  g644(.A1(new_n748), .A2(new_n830), .B1(new_n795), .B2(new_n794), .ZN(new_n831));
  OAI21_X1  g645(.A(new_n827), .B1(new_n829), .B2(new_n831), .ZN(new_n832));
  NAND3_X1  g646(.A1(new_n797), .A2(new_n798), .A3(KEYINPUT52), .ZN(new_n833));
  NAND2_X1  g647(.A1(new_n832), .A2(new_n833), .ZN(new_n834));
  NAND4_X1  g648(.A1(new_n826), .A2(new_n834), .A3(KEYINPUT115), .A4(KEYINPUT53), .ZN(new_n835));
  NAND2_X1  g649(.A1(new_n821), .A2(new_n835), .ZN(new_n836));
  INV_X1    g650(.A(KEYINPUT114), .ZN(new_n837));
  OAI21_X1  g651(.A(new_n837), .B1(new_n799), .B2(new_n800), .ZN(new_n838));
  NAND3_X1  g652(.A1(new_n832), .A2(KEYINPUT114), .A3(new_n833), .ZN(new_n839));
  NAND3_X1  g653(.A1(new_n838), .A2(new_n839), .A3(new_n826), .ZN(new_n840));
  INV_X1    g654(.A(KEYINPUT53), .ZN(new_n841));
  NAND2_X1  g655(.A1(new_n840), .A2(new_n841), .ZN(new_n842));
  XNOR2_X1  g656(.A(KEYINPUT116), .B(KEYINPUT54), .ZN(new_n843));
  NAND3_X1  g657(.A1(new_n836), .A2(new_n842), .A3(new_n843), .ZN(new_n844));
  NAND2_X1  g658(.A1(new_n840), .A2(KEYINPUT53), .ZN(new_n845));
  NAND3_X1  g659(.A1(new_n826), .A2(new_n834), .A3(new_n841), .ZN(new_n846));
  NAND3_X1  g660(.A1(new_n845), .A2(KEYINPUT54), .A3(new_n846), .ZN(new_n847));
  INV_X1    g661(.A(new_n534), .ZN(new_n848));
  AND3_X1   g662(.A1(new_n762), .A2(new_n848), .A3(new_n763), .ZN(new_n849));
  NOR3_X1   g663(.A1(new_n696), .A2(new_n735), .A3(new_n697), .ZN(new_n850));
  NAND2_X1  g664(.A1(new_n849), .A2(new_n850), .ZN(new_n851));
  NAND3_X1  g665(.A1(new_n850), .A2(new_n354), .A3(new_n848), .ZN(new_n852));
  OR2_X1    g666(.A1(new_n852), .A2(new_n662), .ZN(new_n853));
  NAND2_X1  g667(.A1(new_n760), .A2(new_n611), .ZN(new_n854));
  OAI22_X1  g668(.A1(new_n851), .A2(new_n809), .B1(new_n853), .B2(new_n854), .ZN(new_n855));
  OAI21_X1  g669(.A(new_n786), .B1(new_n530), .B2(new_n696), .ZN(new_n856));
  NOR4_X1   g670(.A1(new_n716), .A2(new_n764), .A3(new_n534), .A4(new_n782), .ZN(new_n857));
  AOI21_X1  g671(.A(new_n855), .B1(new_n856), .B2(new_n857), .ZN(new_n858));
  INV_X1    g672(.A(KEYINPUT50), .ZN(new_n859));
  INV_X1    g673(.A(new_n716), .ZN(new_n860));
  NAND3_X1  g674(.A1(new_n849), .A2(new_n860), .A3(new_n698), .ZN(new_n861));
  NOR2_X1   g675(.A1(new_n664), .A2(new_n541), .ZN(new_n862));
  INV_X1    g676(.A(new_n862), .ZN(new_n863));
  OAI21_X1  g677(.A(new_n859), .B1(new_n861), .B2(new_n863), .ZN(new_n864));
  NOR3_X1   g678(.A1(new_n716), .A2(new_n764), .A3(new_n534), .ZN(new_n865));
  NAND4_X1  g679(.A1(new_n865), .A2(KEYINPUT50), .A3(new_n698), .A4(new_n862), .ZN(new_n866));
  NAND2_X1  g680(.A1(new_n864), .A2(new_n866), .ZN(new_n867));
  AND3_X1   g681(.A1(new_n858), .A2(new_n867), .A3(KEYINPUT51), .ZN(new_n868));
  OAI211_X1 g682(.A(G952), .B(new_n329), .C1(new_n853), .C2(new_n613), .ZN(new_n869));
  INV_X1    g683(.A(new_n689), .ZN(new_n870));
  OR3_X1    g684(.A1(new_n851), .A2(KEYINPUT48), .A3(new_n870), .ZN(new_n871));
  OAI21_X1  g685(.A(KEYINPUT48), .B1(new_n851), .B2(new_n870), .ZN(new_n872));
  AOI21_X1  g686(.A(new_n869), .B1(new_n871), .B2(new_n872), .ZN(new_n873));
  OAI21_X1  g687(.A(new_n873), .B1(new_n636), .B2(new_n861), .ZN(new_n874));
  AOI21_X1  g688(.A(KEYINPUT51), .B1(new_n858), .B2(new_n867), .ZN(new_n875));
  NOR3_X1   g689(.A1(new_n868), .A2(new_n874), .A3(new_n875), .ZN(new_n876));
  NAND3_X1  g690(.A1(new_n844), .A2(new_n847), .A3(new_n876), .ZN(new_n877));
  NAND2_X1  g691(.A1(new_n877), .A2(KEYINPUT117), .ZN(new_n878));
  INV_X1    g692(.A(KEYINPUT117), .ZN(new_n879));
  NAND4_X1  g693(.A1(new_n844), .A2(new_n847), .A3(new_n876), .A4(new_n879), .ZN(new_n880));
  INV_X1    g694(.A(G952), .ZN(new_n881));
  NAND2_X1  g695(.A1(new_n881), .A2(new_n329), .ZN(new_n882));
  XNOR2_X1  g696(.A(new_n882), .B(KEYINPUT118), .ZN(new_n883));
  NAND3_X1  g697(.A1(new_n878), .A2(new_n880), .A3(new_n883), .ZN(new_n884));
  OR2_X1    g698(.A1(new_n696), .A2(KEYINPUT49), .ZN(new_n885));
  NAND2_X1  g699(.A1(new_n696), .A2(KEYINPUT49), .ZN(new_n886));
  NOR2_X1   g700(.A1(new_n697), .A2(new_n592), .ZN(new_n887));
  NAND4_X1  g701(.A1(new_n885), .A2(new_n354), .A3(new_n886), .A4(new_n887), .ZN(new_n888));
  OR4_X1    g702(.A1(new_n662), .A2(new_n888), .A3(new_n664), .A4(new_n761), .ZN(new_n889));
  NAND2_X1  g703(.A1(new_n884), .A2(new_n889), .ZN(new_n890));
  NAND2_X1  g704(.A1(new_n890), .A2(KEYINPUT119), .ZN(new_n891));
  INV_X1    g705(.A(KEYINPUT119), .ZN(new_n892));
  NAND3_X1  g706(.A1(new_n884), .A2(new_n892), .A3(new_n889), .ZN(new_n893));
  NAND2_X1  g707(.A1(new_n891), .A2(new_n893), .ZN(G75));
  AOI21_X1  g708(.A(new_n333), .B1(new_n836), .B2(new_n842), .ZN(new_n895));
  AND2_X1   g709(.A1(new_n895), .A2(G210), .ZN(new_n896));
  OR2_X1    g710(.A1(new_n896), .A2(KEYINPUT56), .ZN(new_n897));
  NAND2_X1  g711(.A1(new_n555), .A2(new_n573), .ZN(new_n898));
  XNOR2_X1  g712(.A(new_n898), .B(new_n571), .ZN(new_n899));
  XOR2_X1   g713(.A(new_n899), .B(KEYINPUT55), .Z(new_n900));
  AND2_X1   g714(.A1(new_n897), .A2(new_n900), .ZN(new_n901));
  NAND2_X1  g715(.A1(new_n881), .A2(G953), .ZN(new_n902));
  XOR2_X1   g716(.A(new_n902), .B(KEYINPUT120), .Z(new_n903));
  OAI21_X1  g717(.A(new_n903), .B1(new_n897), .B2(new_n900), .ZN(new_n904));
  NOR2_X1   g718(.A1(new_n901), .A2(new_n904), .ZN(G51));
  INV_X1    g719(.A(new_n903), .ZN(new_n906));
  NAND2_X1  g720(.A1(new_n836), .A2(new_n842), .ZN(new_n907));
  INV_X1    g721(.A(new_n843), .ZN(new_n908));
  NAND2_X1  g722(.A1(new_n907), .A2(new_n908), .ZN(new_n909));
  NAND2_X1  g723(.A1(new_n909), .A2(new_n844), .ZN(new_n910));
  XNOR2_X1  g724(.A(new_n527), .B(KEYINPUT57), .ZN(new_n911));
  AOI22_X1  g725(.A1(new_n910), .A2(new_n911), .B1(new_n691), .B2(new_n692), .ZN(new_n912));
  AOI22_X1  g726(.A1(new_n912), .A2(KEYINPUT121), .B1(new_n776), .B2(new_n895), .ZN(new_n913));
  NAND2_X1  g727(.A1(new_n910), .A2(new_n911), .ZN(new_n914));
  NAND2_X1  g728(.A1(new_n914), .A2(new_n693), .ZN(new_n915));
  INV_X1    g729(.A(KEYINPUT121), .ZN(new_n916));
  NAND2_X1  g730(.A1(new_n915), .A2(new_n916), .ZN(new_n917));
  AOI21_X1  g731(.A(new_n906), .B1(new_n913), .B2(new_n917), .ZN(G54));
  NAND3_X1  g732(.A1(new_n895), .A2(KEYINPUT58), .A3(G475), .ZN(new_n919));
  OR2_X1    g733(.A1(new_n919), .A2(new_n408), .ZN(new_n920));
  NAND2_X1  g734(.A1(new_n919), .A2(new_n408), .ZN(new_n921));
  AOI21_X1  g735(.A(new_n906), .B1(new_n920), .B2(new_n921), .ZN(G60));
  XOR2_X1   g736(.A(KEYINPUT122), .B(KEYINPUT59), .Z(new_n923));
  NOR2_X1   g737(.A1(new_n448), .A2(new_n333), .ZN(new_n924));
  XNOR2_X1  g738(.A(new_n923), .B(new_n924), .ZN(new_n925));
  AND3_X1   g739(.A1(new_n910), .A2(new_n609), .A3(new_n925), .ZN(new_n926));
  NAND2_X1  g740(.A1(new_n844), .A2(new_n847), .ZN(new_n927));
  AOI21_X1  g741(.A(new_n609), .B1(new_n927), .B2(new_n925), .ZN(new_n928));
  NOR3_X1   g742(.A1(new_n926), .A2(new_n928), .A3(new_n906), .ZN(G63));
  INV_X1    g743(.A(KEYINPUT61), .ZN(new_n930));
  NOR2_X1   g744(.A1(new_n930), .A2(KEYINPUT123), .ZN(new_n931));
  NAND2_X1  g745(.A1(G217), .A2(G902), .ZN(new_n932));
  XOR2_X1   g746(.A(new_n932), .B(KEYINPUT60), .Z(new_n933));
  NAND2_X1  g747(.A1(new_n907), .A2(new_n933), .ZN(new_n934));
  NAND2_X1  g748(.A1(new_n332), .A2(new_n334), .ZN(new_n935));
  AOI21_X1  g749(.A(new_n906), .B1(new_n934), .B2(new_n935), .ZN(new_n936));
  NAND3_X1  g750(.A1(new_n907), .A2(new_n629), .A3(new_n933), .ZN(new_n937));
  AOI21_X1  g751(.A(new_n931), .B1(new_n936), .B2(new_n937), .ZN(new_n938));
  AND2_X1   g752(.A1(new_n930), .A2(KEYINPUT123), .ZN(new_n939));
  XNOR2_X1  g753(.A(new_n938), .B(new_n939), .ZN(G66));
  NAND2_X1  g754(.A1(new_n556), .A2(G953), .ZN(new_n941));
  OAI211_X1 g755(.A(new_n538), .B(new_n941), .C1(new_n822), .C2(G953), .ZN(new_n942));
  OAI21_X1  g756(.A(new_n898), .B1(G898), .B2(new_n329), .ZN(new_n943));
  XNOR2_X1  g757(.A(new_n942), .B(new_n943), .ZN(G69));
  NAND2_X1  g758(.A1(new_n399), .A2(new_n401), .ZN(new_n945));
  XNOR2_X1  g759(.A(new_n248), .B(new_n945), .ZN(new_n946));
  AND2_X1   g760(.A1(new_n946), .A2(new_n329), .ZN(new_n947));
  INV_X1    g761(.A(new_n947), .ZN(new_n948));
  NAND4_X1  g762(.A1(new_n689), .A2(new_n649), .A3(new_n736), .A4(new_n815), .ZN(new_n949));
  XOR2_X1   g763(.A(new_n949), .B(KEYINPUT124), .Z(new_n950));
  NAND2_X1  g764(.A1(new_n784), .A2(new_n950), .ZN(new_n951));
  NAND2_X1  g765(.A1(new_n951), .A2(KEYINPUT125), .ZN(new_n952));
  INV_X1    g766(.A(KEYINPUT125), .ZN(new_n953));
  NAND3_X1  g767(.A1(new_n784), .A2(new_n953), .A3(new_n950), .ZN(new_n954));
  AOI22_X1  g768(.A1(new_n952), .A2(new_n954), .B1(new_n787), .B2(new_n788), .ZN(new_n955));
  AND2_X1   g769(.A1(new_n798), .A2(new_n732), .ZN(new_n956));
  NAND2_X1  g770(.A1(new_n956), .A2(new_n667), .ZN(new_n957));
  XOR2_X1   g771(.A(new_n957), .B(KEYINPUT62), .Z(new_n958));
  AOI21_X1  g772(.A(new_n948), .B1(new_n955), .B2(new_n958), .ZN(new_n959));
  NOR2_X1   g773(.A1(new_n329), .A2(G900), .ZN(new_n960));
  NOR3_X1   g774(.A1(new_n781), .A2(new_n870), .A3(new_n795), .ZN(new_n961));
  AOI21_X1  g775(.A(new_n961), .B1(new_n787), .B2(new_n788), .ZN(new_n962));
  NAND4_X1  g776(.A1(new_n784), .A2(new_n962), .A3(new_n802), .A4(new_n956), .ZN(new_n963));
  AOI211_X1 g777(.A(new_n960), .B(new_n946), .C1(new_n963), .C2(new_n329), .ZN(new_n964));
  OR3_X1    g778(.A1(new_n959), .A2(KEYINPUT126), .A3(new_n964), .ZN(new_n965));
  OAI21_X1  g779(.A(KEYINPUT126), .B1(new_n959), .B2(new_n964), .ZN(new_n966));
  INV_X1    g780(.A(G900), .ZN(new_n967));
  OAI21_X1  g781(.A(G953), .B1(new_n458), .B2(new_n967), .ZN(new_n968));
  AND3_X1   g782(.A1(new_n965), .A2(new_n966), .A3(new_n968), .ZN(new_n969));
  AOI21_X1  g783(.A(new_n968), .B1(new_n965), .B2(new_n966), .ZN(new_n970));
  NOR2_X1   g784(.A1(new_n969), .A2(new_n970), .ZN(G72));
  NAND3_X1  g785(.A1(new_n955), .A2(new_n822), .A3(new_n958), .ZN(new_n972));
  NAND2_X1  g786(.A1(G472), .A2(G902), .ZN(new_n973));
  XOR2_X1   g787(.A(new_n973), .B(KEYINPUT63), .Z(new_n974));
  NAND2_X1  g788(.A1(new_n972), .A2(new_n974), .ZN(new_n975));
  NAND2_X1  g789(.A1(new_n975), .A2(new_n658), .ZN(new_n976));
  OAI21_X1  g790(.A(new_n974), .B1(new_n273), .B2(new_n262), .ZN(new_n977));
  NOR3_X1   g791(.A1(new_n288), .A2(new_n272), .A3(new_n259), .ZN(new_n978));
  NOR2_X1   g792(.A1(new_n977), .A2(new_n978), .ZN(new_n979));
  NAND3_X1  g793(.A1(new_n845), .A2(new_n846), .A3(new_n979), .ZN(new_n980));
  INV_X1    g794(.A(new_n822), .ZN(new_n981));
  OAI21_X1  g795(.A(new_n974), .B1(new_n963), .B2(new_n981), .ZN(new_n982));
  AOI21_X1  g796(.A(new_n906), .B1(new_n982), .B2(new_n978), .ZN(new_n983));
  NAND3_X1  g797(.A1(new_n976), .A2(new_n980), .A3(new_n983), .ZN(new_n984));
  NAND2_X1  g798(.A1(new_n984), .A2(KEYINPUT127), .ZN(new_n985));
  INV_X1    g799(.A(KEYINPUT127), .ZN(new_n986));
  NAND4_X1  g800(.A1(new_n976), .A2(new_n986), .A3(new_n980), .A4(new_n983), .ZN(new_n987));
  NAND2_X1  g801(.A1(new_n985), .A2(new_n987), .ZN(G57));
endmodule


