

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n511, n512, n513, n514,
         n515, n516, n517, n518, n519, n520, n521, n522, n523, n524, n525,
         n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536,
         n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547,
         n548, n549, n550, n551, n552, n553, n555, n556, n557, n558, n559,
         n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570,
         n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581,
         n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592,
         n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603,
         n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614,
         n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625,
         n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636,
         n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647,
         n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658,
         n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669,
         n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680,
         n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691,
         n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702,
         n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713,
         n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724,
         n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735,
         n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746,
         n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757,
         n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768,
         n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, n779,
         n780, n781, n782, n783, n784, n785, n786, n787, n788, n789, n790,
         n791, n792, n793, n794, n795, n796, n797, n798, n799, n800, n801,
         n802, n803, n804, n805, n806, n807, n808, n809, n810, n811, n812,
         n813, n814, n815, n816, n817, n818, n819, n820, n821, n822, n823,
         n824, n825, n826, n827, n828, n829, n830, n831, n832, n833, n834,
         n835, n836, n837, n838, n839, n840, n841, n842, n843, n844, n845,
         n846, n847, n848, n849, n850, n851, n852, n853, n854, n855, n856,
         n857, n858, n859, n860, n861, n862, n863, n864, n865, n866, n867,
         n868, n869, n870, n871, n872, n873, n874, n875, n876, n877, n878,
         n879, n880, n881, n882, n883, n884, n885, n886, n887, n888, n889,
         n890, n891, n892, n893, n894, n895, n896, n897, n898, n899, n900,
         n901, n902, n903, n904, n905, n906, n907, n908, n909, n910, n911,
         n912, n913, n914, n915, n916, n917, n918, n919, n920, n921, n922,
         n923, n924, n925, n926, n927, n928, n929, n930, n931, n932, n933,
         n934, n935, n936, n937, n938, n939, n940, n941, n942, n943, n944,
         n945, n946, n947, n948, n949, n950, n951, n952, n953, n954, n955,
         n956, n957, n958, n959, n960, n961, n962, n963, n964, n965, n966,
         n967, n968, n969, n970, n971, n972, n973, n974, n975, n976, n977,
         n978, n979, n980, n981, n982, n983, n984, n985, n986, n987, n988,
         n989, n990, n991, n992, n993, n994, n995, n996, n997, n998, n999,
         n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009,
         n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019,
         n1020, n1021, n1022, n1023;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NOR2_X1 U545 ( .A1(G164), .A2(G1384), .ZN(n801) );
  NOR2_X1 U546 ( .A1(G651), .A2(n532), .ZN(n666) );
  INV_X2 U547 ( .A(n704), .ZN(n711) );
  XNOR2_X1 U548 ( .A(n626), .B(KEYINPUT15), .ZN(n996) );
  OR2_X1 U549 ( .A1(n717), .A2(n716), .ZN(n718) );
  NOR2_X1 U550 ( .A1(n715), .A2(n714), .ZN(n716) );
  OR2_X1 U551 ( .A1(n754), .A2(n731), .ZN(n732) );
  BUF_X1 U552 ( .A(n573), .Z(n574) );
  NOR2_X1 U553 ( .A1(G2105), .A2(n543), .ZN(n555) );
  NOR2_X2 U554 ( .A1(G2104), .A2(n548), .ZN(n893) );
  XNOR2_X1 U555 ( .A(KEYINPUT65), .B(KEYINPUT17), .ZN(n542) );
  XNOR2_X2 U556 ( .A(n759), .B(KEYINPUT95), .ZN(n773) );
  AND2_X1 U557 ( .A1(n704), .A2(G1341), .ZN(n706) );
  OR2_X1 U558 ( .A1(n706), .A2(n705), .ZN(n707) );
  INV_X1 U559 ( .A(KEYINPUT29), .ZN(n722) );
  NOR2_X1 U560 ( .A1(n735), .A2(n734), .ZN(n736) );
  INV_X1 U561 ( .A(KEYINPUT84), .ZN(n696) );
  NAND2_X1 U562 ( .A1(n618), .A2(n617), .ZN(n705) );
  INV_X1 U563 ( .A(KEYINPUT1), .ZN(n529) );
  XNOR2_X2 U564 ( .A(n530), .B(n529), .ZN(n607) );
  XNOR2_X1 U565 ( .A(KEYINPUT28), .B(n720), .ZN(n511) );
  OR2_X1 U566 ( .A1(n727), .A2(G301), .ZN(n512) );
  OR2_X1 U567 ( .A1(G299), .A2(n719), .ZN(n513) );
  XNOR2_X1 U568 ( .A(KEYINPUT96), .B(n1010), .ZN(n514) );
  XOR2_X1 U569 ( .A(n722), .B(KEYINPUT91), .Z(n515) );
  AND2_X1 U570 ( .A1(n812), .A2(n823), .ZN(n516) );
  OR2_X1 U571 ( .A1(n741), .A2(n766), .ZN(n517) );
  NOR2_X1 U572 ( .A1(n741), .A2(n762), .ZN(n518) );
  XOR2_X1 U573 ( .A(KEYINPUT31), .B(KEYINPUT92), .Z(n519) );
  AND2_X1 U574 ( .A1(n763), .A2(n518), .ZN(n520) );
  NOR2_X1 U575 ( .A1(n708), .A2(n707), .ZN(n710) );
  INV_X1 U576 ( .A(G8), .ZN(n730) );
  OR2_X1 U577 ( .A1(n751), .A2(n730), .ZN(n731) );
  INV_X1 U578 ( .A(KEYINPUT93), .ZN(n739) );
  BUF_X1 U579 ( .A(n704), .Z(n742) );
  INV_X1 U580 ( .A(n1005), .ZN(n762) );
  INV_X1 U581 ( .A(KEYINPUT85), .ZN(n728) );
  XNOR2_X1 U582 ( .A(n729), .B(n728), .ZN(n741) );
  NAND2_X1 U583 ( .A1(n993), .A2(n517), .ZN(n767) );
  NAND2_X1 U584 ( .A1(n607), .A2(G56), .ZN(n608) );
  INV_X1 U585 ( .A(KEYINPUT23), .ZN(n544) );
  NOR2_X1 U586 ( .A1(n623), .A2(n622), .ZN(n624) );
  INV_X1 U587 ( .A(KEYINPUT66), .ZN(n523) );
  INV_X1 U588 ( .A(G2105), .ZN(n548) );
  XNOR2_X1 U589 ( .A(n524), .B(n523), .ZN(n532) );
  NOR2_X2 U590 ( .A1(G651), .A2(G543), .ZN(n660) );
  BUF_X1 U591 ( .A(n555), .Z(n897) );
  NOR2_X1 U592 ( .A1(n553), .A2(n552), .ZN(n695) );
  BUF_X1 U593 ( .A(n705), .Z(n1001) );
  NAND2_X1 U594 ( .A1(G89), .A2(n660), .ZN(n521) );
  XOR2_X1 U595 ( .A(KEYINPUT4), .B(n521), .Z(n522) );
  XNOR2_X1 U596 ( .A(n522), .B(KEYINPUT73), .ZN(n526) );
  XNOR2_X1 U597 ( .A(G543), .B(KEYINPUT0), .ZN(n524) );
  INV_X1 U598 ( .A(G651), .ZN(n528) );
  NOR2_X1 U599 ( .A1(n532), .A2(n528), .ZN(n610) );
  BUF_X1 U600 ( .A(n610), .Z(n661) );
  NAND2_X1 U601 ( .A1(G76), .A2(n661), .ZN(n525) );
  NAND2_X1 U602 ( .A1(n526), .A2(n525), .ZN(n527) );
  XNOR2_X1 U603 ( .A(n527), .B(KEYINPUT5), .ZN(n538) );
  XNOR2_X1 U604 ( .A(KEYINPUT75), .B(KEYINPUT6), .ZN(n536) );
  NOR2_X1 U605 ( .A1(n528), .A2(G543), .ZN(n530) );
  NAND2_X1 U606 ( .A1(n607), .A2(G63), .ZN(n531) );
  XNOR2_X1 U607 ( .A(n531), .B(KEYINPUT74), .ZN(n534) );
  NAND2_X1 U608 ( .A1(G51), .A2(n666), .ZN(n533) );
  NAND2_X1 U609 ( .A1(n534), .A2(n533), .ZN(n535) );
  XNOR2_X1 U610 ( .A(n536), .B(n535), .ZN(n537) );
  NAND2_X1 U611 ( .A1(n538), .A2(n537), .ZN(n540) );
  XNOR2_X1 U612 ( .A(KEYINPUT76), .B(KEYINPUT7), .ZN(n539) );
  XNOR2_X1 U613 ( .A(n540), .B(n539), .ZN(G168) );
  XOR2_X1 U614 ( .A(KEYINPUT8), .B(G168), .Z(G286) );
  NOR2_X1 U615 ( .A1(G2105), .A2(G2104), .ZN(n541) );
  XNOR2_X1 U616 ( .A(n542), .B(n541), .ZN(n573) );
  NAND2_X1 U617 ( .A1(n573), .A2(G137), .ZN(n547) );
  INV_X1 U618 ( .A(G2104), .ZN(n543) );
  NAND2_X1 U619 ( .A1(n555), .A2(G101), .ZN(n545) );
  XNOR2_X1 U620 ( .A(n545), .B(n544), .ZN(n546) );
  NAND2_X1 U621 ( .A1(n547), .A2(n546), .ZN(n553) );
  NAND2_X1 U622 ( .A1(n893), .A2(G125), .ZN(n551) );
  NAND2_X1 U623 ( .A1(G2104), .A2(G2105), .ZN(n549) );
  XOR2_X1 U624 ( .A(KEYINPUT64), .B(n549), .Z(n577) );
  NAND2_X1 U625 ( .A1(G113), .A2(n577), .ZN(n550) );
  NAND2_X1 U626 ( .A1(n551), .A2(n550), .ZN(n552) );
  BUF_X1 U627 ( .A(n695), .Z(G160) );
  NAND2_X1 U628 ( .A1(G102), .A2(n897), .ZN(n557) );
  NAND2_X1 U629 ( .A1(G138), .A2(n573), .ZN(n556) );
  NAND2_X1 U630 ( .A1(n557), .A2(n556), .ZN(n561) );
  NAND2_X1 U631 ( .A1(n893), .A2(G126), .ZN(n559) );
  NAND2_X1 U632 ( .A1(G114), .A2(n577), .ZN(n558) );
  NAND2_X1 U633 ( .A1(n559), .A2(n558), .ZN(n560) );
  NOR2_X1 U634 ( .A1(n561), .A2(n560), .ZN(G164) );
  XOR2_X1 U635 ( .A(G2446), .B(G2430), .Z(n563) );
  XNOR2_X1 U636 ( .A(G2451), .B(G2454), .ZN(n562) );
  XNOR2_X1 U637 ( .A(n563), .B(n562), .ZN(n564) );
  XOR2_X1 U638 ( .A(n564), .B(G2427), .Z(n566) );
  XNOR2_X1 U639 ( .A(G1348), .B(G1341), .ZN(n565) );
  XNOR2_X1 U640 ( .A(n566), .B(n565), .ZN(n570) );
  XOR2_X1 U641 ( .A(G2443), .B(KEYINPUT102), .Z(n568) );
  XNOR2_X1 U642 ( .A(G2438), .B(G2435), .ZN(n567) );
  XNOR2_X1 U643 ( .A(n568), .B(n567), .ZN(n569) );
  XOR2_X1 U644 ( .A(n570), .B(n569), .Z(n571) );
  AND2_X1 U645 ( .A1(G14), .A2(n571), .ZN(G401) );
  AND2_X1 U646 ( .A1(G452), .A2(G94), .ZN(G173) );
  NAND2_X1 U647 ( .A1(G123), .A2(n893), .ZN(n572) );
  XNOR2_X1 U648 ( .A(n572), .B(KEYINPUT18), .ZN(n582) );
  NAND2_X1 U649 ( .A1(G99), .A2(n897), .ZN(n576) );
  NAND2_X1 U650 ( .A1(G135), .A2(n574), .ZN(n575) );
  NAND2_X1 U651 ( .A1(n576), .A2(n575), .ZN(n580) );
  BUF_X1 U652 ( .A(n577), .Z(n894) );
  NAND2_X1 U653 ( .A1(G111), .A2(n894), .ZN(n578) );
  XNOR2_X1 U654 ( .A(KEYINPUT77), .B(n578), .ZN(n579) );
  NOR2_X1 U655 ( .A1(n580), .A2(n579), .ZN(n581) );
  NAND2_X1 U656 ( .A1(n582), .A2(n581), .ZN(n919) );
  XNOR2_X1 U657 ( .A(G2096), .B(n919), .ZN(n583) );
  OR2_X1 U658 ( .A1(G2100), .A2(n583), .ZN(G156) );
  INV_X1 U659 ( .A(G57), .ZN(G237) );
  INV_X1 U660 ( .A(G132), .ZN(G219) );
  INV_X1 U661 ( .A(G82), .ZN(G220) );
  NAND2_X1 U662 ( .A1(G88), .A2(n660), .ZN(n585) );
  NAND2_X1 U663 ( .A1(G75), .A2(n661), .ZN(n584) );
  NAND2_X1 U664 ( .A1(n585), .A2(n584), .ZN(n589) );
  NAND2_X1 U665 ( .A1(G62), .A2(n607), .ZN(n587) );
  NAND2_X1 U666 ( .A1(G50), .A2(n666), .ZN(n586) );
  NAND2_X1 U667 ( .A1(n587), .A2(n586), .ZN(n588) );
  NOR2_X1 U668 ( .A1(n589), .A2(n588), .ZN(G166) );
  NAND2_X1 U669 ( .A1(G91), .A2(n660), .ZN(n591) );
  NAND2_X1 U670 ( .A1(G78), .A2(n661), .ZN(n590) );
  NAND2_X1 U671 ( .A1(n591), .A2(n590), .ZN(n594) );
  NAND2_X1 U672 ( .A1(G65), .A2(n607), .ZN(n592) );
  XNOR2_X1 U673 ( .A(KEYINPUT67), .B(n592), .ZN(n593) );
  NOR2_X1 U674 ( .A1(n594), .A2(n593), .ZN(n596) );
  NAND2_X1 U675 ( .A1(n666), .A2(G53), .ZN(n595) );
  NAND2_X1 U676 ( .A1(n596), .A2(n595), .ZN(G299) );
  NAND2_X1 U677 ( .A1(G90), .A2(n660), .ZN(n598) );
  NAND2_X1 U678 ( .A1(G77), .A2(n661), .ZN(n597) );
  NAND2_X1 U679 ( .A1(n598), .A2(n597), .ZN(n599) );
  XNOR2_X1 U680 ( .A(KEYINPUT9), .B(n599), .ZN(n603) );
  NAND2_X1 U681 ( .A1(G64), .A2(n607), .ZN(n601) );
  NAND2_X1 U682 ( .A1(G52), .A2(n666), .ZN(n600) );
  AND2_X1 U683 ( .A1(n601), .A2(n600), .ZN(n602) );
  NAND2_X1 U684 ( .A1(n603), .A2(n602), .ZN(G301) );
  NAND2_X1 U685 ( .A1(G7), .A2(G661), .ZN(n604) );
  XNOR2_X1 U686 ( .A(n604), .B(KEYINPUT10), .ZN(G223) );
  XOR2_X1 U687 ( .A(KEYINPUT68), .B(KEYINPUT11), .Z(n606) );
  INV_X1 U688 ( .A(G223), .ZN(n832) );
  NAND2_X1 U689 ( .A1(G567), .A2(n832), .ZN(n605) );
  XNOR2_X1 U690 ( .A(n606), .B(n605), .ZN(G234) );
  XNOR2_X1 U691 ( .A(KEYINPUT14), .B(n608), .ZN(n615) );
  NAND2_X1 U692 ( .A1(n660), .A2(G81), .ZN(n609) );
  XNOR2_X1 U693 ( .A(n609), .B(KEYINPUT12), .ZN(n612) );
  NAND2_X1 U694 ( .A1(G68), .A2(n610), .ZN(n611) );
  NAND2_X1 U695 ( .A1(n612), .A2(n611), .ZN(n613) );
  XNOR2_X1 U696 ( .A(n613), .B(KEYINPUT13), .ZN(n614) );
  NAND2_X1 U697 ( .A1(n615), .A2(n614), .ZN(n616) );
  XNOR2_X1 U698 ( .A(n616), .B(KEYINPUT69), .ZN(n618) );
  NAND2_X1 U699 ( .A1(n666), .A2(G43), .ZN(n617) );
  INV_X1 U700 ( .A(G860), .ZN(n633) );
  OR2_X1 U701 ( .A1(n1001), .A2(n633), .ZN(G153) );
  NAND2_X1 U702 ( .A1(G54), .A2(n666), .ZN(n625) );
  NAND2_X1 U703 ( .A1(G66), .A2(n607), .ZN(n620) );
  NAND2_X1 U704 ( .A1(G79), .A2(n661), .ZN(n619) );
  NAND2_X1 U705 ( .A1(n620), .A2(n619), .ZN(n623) );
  NAND2_X1 U706 ( .A1(n660), .A2(G92), .ZN(n621) );
  XOR2_X1 U707 ( .A(KEYINPUT70), .B(n621), .Z(n622) );
  NAND2_X1 U708 ( .A1(n625), .A2(n624), .ZN(n626) );
  NOR2_X1 U709 ( .A1(n996), .A2(G868), .ZN(n627) );
  XNOR2_X1 U710 ( .A(n627), .B(KEYINPUT71), .ZN(n629) );
  NAND2_X1 U711 ( .A1(G868), .A2(G301), .ZN(n628) );
  NAND2_X1 U712 ( .A1(n629), .A2(n628), .ZN(n630) );
  XNOR2_X1 U713 ( .A(KEYINPUT72), .B(n630), .ZN(G284) );
  NAND2_X1 U714 ( .A1(G868), .A2(G286), .ZN(n632) );
  INV_X1 U715 ( .A(G868), .ZN(n678) );
  NAND2_X1 U716 ( .A1(G299), .A2(n678), .ZN(n631) );
  NAND2_X1 U717 ( .A1(n632), .A2(n631), .ZN(G297) );
  NAND2_X1 U718 ( .A1(n633), .A2(G559), .ZN(n634) );
  NAND2_X1 U719 ( .A1(n634), .A2(n996), .ZN(n635) );
  XNOR2_X1 U720 ( .A(n635), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U721 ( .A1(G868), .A2(n1001), .ZN(n638) );
  NAND2_X1 U722 ( .A1(G868), .A2(n996), .ZN(n636) );
  NOR2_X1 U723 ( .A1(G559), .A2(n636), .ZN(n637) );
  NOR2_X1 U724 ( .A1(n638), .A2(n637), .ZN(G282) );
  NAND2_X1 U725 ( .A1(n996), .A2(G559), .ZN(n676) );
  XNOR2_X1 U726 ( .A(n1001), .B(n676), .ZN(n639) );
  NOR2_X1 U727 ( .A1(n639), .A2(G860), .ZN(n647) );
  NAND2_X1 U728 ( .A1(G93), .A2(n660), .ZN(n640) );
  XNOR2_X1 U729 ( .A(n640), .B(KEYINPUT78), .ZN(n642) );
  NAND2_X1 U730 ( .A1(n607), .A2(G67), .ZN(n641) );
  NAND2_X1 U731 ( .A1(n642), .A2(n641), .ZN(n646) );
  NAND2_X1 U732 ( .A1(G80), .A2(n661), .ZN(n644) );
  NAND2_X1 U733 ( .A1(G55), .A2(n666), .ZN(n643) );
  NAND2_X1 U734 ( .A1(n644), .A2(n643), .ZN(n645) );
  OR2_X1 U735 ( .A1(n646), .A2(n645), .ZN(n679) );
  XOR2_X1 U736 ( .A(n647), .B(n679), .Z(G145) );
  NAND2_X1 U737 ( .A1(G49), .A2(n666), .ZN(n649) );
  NAND2_X1 U738 ( .A1(G74), .A2(G651), .ZN(n648) );
  NAND2_X1 U739 ( .A1(n649), .A2(n648), .ZN(n650) );
  NOR2_X1 U740 ( .A1(n607), .A2(n650), .ZN(n652) );
  NAND2_X1 U741 ( .A1(G87), .A2(n532), .ZN(n651) );
  NAND2_X1 U742 ( .A1(n652), .A2(n651), .ZN(G288) );
  NAND2_X1 U743 ( .A1(G61), .A2(n607), .ZN(n654) );
  NAND2_X1 U744 ( .A1(G86), .A2(n660), .ZN(n653) );
  NAND2_X1 U745 ( .A1(n654), .A2(n653), .ZN(n657) );
  NAND2_X1 U746 ( .A1(n661), .A2(G73), .ZN(n655) );
  XOR2_X1 U747 ( .A(KEYINPUT2), .B(n655), .Z(n656) );
  NOR2_X1 U748 ( .A1(n657), .A2(n656), .ZN(n659) );
  NAND2_X1 U749 ( .A1(n666), .A2(G48), .ZN(n658) );
  NAND2_X1 U750 ( .A1(n659), .A2(n658), .ZN(G305) );
  AND2_X1 U751 ( .A1(n607), .A2(G60), .ZN(n665) );
  NAND2_X1 U752 ( .A1(G85), .A2(n660), .ZN(n663) );
  NAND2_X1 U753 ( .A1(G72), .A2(n661), .ZN(n662) );
  NAND2_X1 U754 ( .A1(n663), .A2(n662), .ZN(n664) );
  NOR2_X1 U755 ( .A1(n665), .A2(n664), .ZN(n668) );
  NAND2_X1 U756 ( .A1(n666), .A2(G47), .ZN(n667) );
  NAND2_X1 U757 ( .A1(n668), .A2(n667), .ZN(G290) );
  XNOR2_X1 U758 ( .A(G166), .B(G299), .ZN(n675) );
  XOR2_X1 U759 ( .A(KEYINPUT79), .B(KEYINPUT19), .Z(n669) );
  XNOR2_X1 U760 ( .A(G288), .B(n669), .ZN(n670) );
  XNOR2_X1 U761 ( .A(n670), .B(n1001), .ZN(n671) );
  XNOR2_X1 U762 ( .A(n671), .B(G305), .ZN(n672) );
  XOR2_X1 U763 ( .A(n679), .B(n672), .Z(n673) );
  XNOR2_X1 U764 ( .A(n673), .B(G290), .ZN(n674) );
  XNOR2_X1 U765 ( .A(n675), .B(n674), .ZN(n840) );
  XOR2_X1 U766 ( .A(n840), .B(n676), .Z(n677) );
  NAND2_X1 U767 ( .A1(G868), .A2(n677), .ZN(n681) );
  NAND2_X1 U768 ( .A1(n679), .A2(n678), .ZN(n680) );
  NAND2_X1 U769 ( .A1(n681), .A2(n680), .ZN(G295) );
  NAND2_X1 U770 ( .A1(G2084), .A2(G2078), .ZN(n682) );
  XOR2_X1 U771 ( .A(KEYINPUT20), .B(n682), .Z(n683) );
  NAND2_X1 U772 ( .A1(G2090), .A2(n683), .ZN(n684) );
  XNOR2_X1 U773 ( .A(KEYINPUT21), .B(n684), .ZN(n685) );
  NAND2_X1 U774 ( .A1(n685), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U775 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U776 ( .A1(G220), .A2(G219), .ZN(n686) );
  XOR2_X1 U777 ( .A(KEYINPUT22), .B(n686), .Z(n687) );
  NOR2_X1 U778 ( .A1(G218), .A2(n687), .ZN(n688) );
  NAND2_X1 U779 ( .A1(G96), .A2(n688), .ZN(n838) );
  NAND2_X1 U780 ( .A1(n838), .A2(G2106), .ZN(n692) );
  NAND2_X1 U781 ( .A1(G69), .A2(G120), .ZN(n689) );
  NOR2_X1 U782 ( .A1(G237), .A2(n689), .ZN(n690) );
  NAND2_X1 U783 ( .A1(G108), .A2(n690), .ZN(n837) );
  NAND2_X1 U784 ( .A1(n837), .A2(G567), .ZN(n691) );
  NAND2_X1 U785 ( .A1(n692), .A2(n691), .ZN(n915) );
  NAND2_X1 U786 ( .A1(G661), .A2(G483), .ZN(n693) );
  XNOR2_X1 U787 ( .A(KEYINPUT80), .B(n693), .ZN(n694) );
  NOR2_X1 U788 ( .A1(n915), .A2(n694), .ZN(n836) );
  NAND2_X1 U789 ( .A1(n836), .A2(G36), .ZN(G176) );
  INV_X1 U790 ( .A(G166), .ZN(G303) );
  NAND2_X1 U791 ( .A1(n695), .A2(G40), .ZN(n800) );
  XNOR2_X1 U792 ( .A(n800), .B(n696), .ZN(n697) );
  NAND2_X1 U793 ( .A1(n697), .A2(n801), .ZN(n704) );
  AND2_X1 U794 ( .A1(n711), .A2(G2072), .ZN(n698) );
  XNOR2_X1 U795 ( .A(n698), .B(KEYINPUT27), .ZN(n701) );
  XNOR2_X1 U796 ( .A(KEYINPUT88), .B(G1956), .ZN(n973) );
  NAND2_X1 U797 ( .A1(n704), .A2(n973), .ZN(n699) );
  XOR2_X1 U798 ( .A(KEYINPUT89), .B(n699), .Z(n700) );
  NAND2_X1 U799 ( .A1(n701), .A2(n700), .ZN(n719) );
  NAND2_X1 U800 ( .A1(n711), .A2(G1996), .ZN(n703) );
  INV_X1 U801 ( .A(KEYINPUT26), .ZN(n702) );
  XNOR2_X1 U802 ( .A(n703), .B(n702), .ZN(n708) );
  NAND2_X1 U803 ( .A1(n996), .A2(n710), .ZN(n709) );
  NAND2_X1 U804 ( .A1(n513), .A2(n709), .ZN(n717) );
  NOR2_X1 U805 ( .A1(n710), .A2(n996), .ZN(n715) );
  NAND2_X1 U806 ( .A1(G1348), .A2(n742), .ZN(n713) );
  NAND2_X1 U807 ( .A1(G2067), .A2(n711), .ZN(n712) );
  NAND2_X1 U808 ( .A1(n713), .A2(n712), .ZN(n714) );
  XNOR2_X1 U809 ( .A(n718), .B(KEYINPUT90), .ZN(n721) );
  NAND2_X1 U810 ( .A1(G299), .A2(n719), .ZN(n720) );
  NAND2_X1 U811 ( .A1(n721), .A2(n511), .ZN(n723) );
  XNOR2_X1 U812 ( .A(n723), .B(n515), .ZN(n726) );
  XOR2_X1 U813 ( .A(KEYINPUT87), .B(G1961), .Z(n977) );
  NOR2_X1 U814 ( .A1(n711), .A2(n977), .ZN(n725) );
  XOR2_X1 U815 ( .A(G2078), .B(KEYINPUT25), .Z(n950) );
  NOR2_X1 U816 ( .A1(n950), .A2(n742), .ZN(n724) );
  NOR2_X1 U817 ( .A1(n725), .A2(n724), .ZN(n727) );
  NAND2_X1 U818 ( .A1(n726), .A2(n512), .ZN(n738) );
  AND2_X1 U819 ( .A1(G301), .A2(n727), .ZN(n735) );
  NAND2_X1 U820 ( .A1(n704), .A2(G8), .ZN(n729) );
  NOR2_X1 U821 ( .A1(G1966), .A2(n741), .ZN(n754) );
  NOR2_X1 U822 ( .A1(G2084), .A2(n742), .ZN(n751) );
  XNOR2_X1 U823 ( .A(n732), .B(KEYINPUT30), .ZN(n733) );
  NOR2_X1 U824 ( .A1(n733), .A2(G168), .ZN(n734) );
  XNOR2_X1 U825 ( .A(n736), .B(n519), .ZN(n737) );
  NAND2_X1 U826 ( .A1(n738), .A2(n737), .ZN(n752) );
  NAND2_X1 U827 ( .A1(n752), .A2(G286), .ZN(n740) );
  XNOR2_X1 U828 ( .A(n740), .B(n739), .ZN(n747) );
  NOR2_X1 U829 ( .A1(G1971), .A2(n741), .ZN(n744) );
  NOR2_X1 U830 ( .A1(G2090), .A2(n742), .ZN(n743) );
  NOR2_X1 U831 ( .A1(n744), .A2(n743), .ZN(n745) );
  NAND2_X1 U832 ( .A1(G303), .A2(n745), .ZN(n746) );
  NAND2_X1 U833 ( .A1(n747), .A2(n746), .ZN(n748) );
  NAND2_X1 U834 ( .A1(n748), .A2(G8), .ZN(n750) );
  XNOR2_X1 U835 ( .A(KEYINPUT94), .B(KEYINPUT32), .ZN(n749) );
  XNOR2_X1 U836 ( .A(n750), .B(n749), .ZN(n758) );
  NAND2_X1 U837 ( .A1(n751), .A2(G8), .ZN(n756) );
  INV_X1 U838 ( .A(n752), .ZN(n753) );
  NOR2_X1 U839 ( .A1(n754), .A2(n753), .ZN(n755) );
  NAND2_X1 U840 ( .A1(n756), .A2(n755), .ZN(n757) );
  NAND2_X1 U841 ( .A1(n758), .A2(n757), .ZN(n759) );
  INV_X1 U842 ( .A(n773), .ZN(n761) );
  NOR2_X1 U843 ( .A1(G1976), .A2(G288), .ZN(n765) );
  NOR2_X1 U844 ( .A1(G1971), .A2(G303), .ZN(n760) );
  NOR2_X1 U845 ( .A1(n765), .A2(n760), .ZN(n1010) );
  NAND2_X1 U846 ( .A1(n761), .A2(n514), .ZN(n763) );
  NAND2_X1 U847 ( .A1(G1976), .A2(G288), .ZN(n1005) );
  NOR2_X1 U848 ( .A1(KEYINPUT33), .A2(n520), .ZN(n768) );
  XNOR2_X1 U849 ( .A(G1981), .B(KEYINPUT97), .ZN(n764) );
  XNOR2_X1 U850 ( .A(n764), .B(G305), .ZN(n993) );
  NAND2_X1 U851 ( .A1(n765), .A2(KEYINPUT33), .ZN(n766) );
  OR2_X1 U852 ( .A1(n768), .A2(n767), .ZN(n769) );
  XNOR2_X1 U853 ( .A(n769), .B(KEYINPUT98), .ZN(n781) );
  NOR2_X1 U854 ( .A1(G1981), .A2(G305), .ZN(n770) );
  XNOR2_X1 U855 ( .A(n770), .B(KEYINPUT24), .ZN(n771) );
  XNOR2_X1 U856 ( .A(n771), .B(KEYINPUT86), .ZN(n772) );
  INV_X1 U857 ( .A(n741), .ZN(n776) );
  AND2_X1 U858 ( .A1(n772), .A2(n776), .ZN(n779) );
  NAND2_X1 U859 ( .A1(G8), .A2(G166), .ZN(n774) );
  NOR2_X1 U860 ( .A1(G2090), .A2(n774), .ZN(n775) );
  NOR2_X1 U861 ( .A1(n773), .A2(n775), .ZN(n777) );
  NOR2_X1 U862 ( .A1(n777), .A2(n776), .ZN(n778) );
  NOR2_X1 U863 ( .A1(n779), .A2(n778), .ZN(n780) );
  NAND2_X1 U864 ( .A1(n781), .A2(n780), .ZN(n813) );
  NAND2_X1 U865 ( .A1(G95), .A2(n897), .ZN(n783) );
  NAND2_X1 U866 ( .A1(G131), .A2(n574), .ZN(n782) );
  NAND2_X1 U867 ( .A1(n783), .A2(n782), .ZN(n784) );
  XNOR2_X1 U868 ( .A(KEYINPUT81), .B(n784), .ZN(n788) );
  NAND2_X1 U869 ( .A1(n894), .A2(G107), .ZN(n786) );
  NAND2_X1 U870 ( .A1(n893), .A2(G119), .ZN(n785) );
  AND2_X1 U871 ( .A1(n786), .A2(n785), .ZN(n787) );
  NAND2_X1 U872 ( .A1(n788), .A2(n787), .ZN(n892) );
  NAND2_X1 U873 ( .A1(G1991), .A2(n892), .ZN(n798) );
  NAND2_X1 U874 ( .A1(n894), .A2(G117), .ZN(n789) );
  XNOR2_X1 U875 ( .A(n789), .B(KEYINPUT82), .ZN(n796) );
  NAND2_X1 U876 ( .A1(G141), .A2(n574), .ZN(n791) );
  NAND2_X1 U877 ( .A1(G129), .A2(n893), .ZN(n790) );
  NAND2_X1 U878 ( .A1(n791), .A2(n790), .ZN(n794) );
  NAND2_X1 U879 ( .A1(n897), .A2(G105), .ZN(n792) );
  XOR2_X1 U880 ( .A(KEYINPUT38), .B(n792), .Z(n793) );
  NOR2_X1 U881 ( .A1(n794), .A2(n793), .ZN(n795) );
  NAND2_X1 U882 ( .A1(n796), .A2(n795), .ZN(n905) );
  NAND2_X1 U883 ( .A1(G1996), .A2(n905), .ZN(n797) );
  NAND2_X1 U884 ( .A1(n798), .A2(n797), .ZN(n799) );
  XNOR2_X1 U885 ( .A(KEYINPUT83), .B(n799), .ZN(n816) );
  XOR2_X1 U886 ( .A(G1986), .B(G290), .Z(n1007) );
  NAND2_X1 U887 ( .A1(n816), .A2(n1007), .ZN(n802) );
  NOR2_X1 U888 ( .A1(n801), .A2(n800), .ZN(n828) );
  NAND2_X1 U889 ( .A1(n802), .A2(n828), .ZN(n812) );
  XNOR2_X1 U890 ( .A(KEYINPUT37), .B(G2067), .ZN(n825) );
  NAND2_X1 U891 ( .A1(G104), .A2(n897), .ZN(n804) );
  NAND2_X1 U892 ( .A1(G140), .A2(n574), .ZN(n803) );
  NAND2_X1 U893 ( .A1(n804), .A2(n803), .ZN(n805) );
  XNOR2_X1 U894 ( .A(KEYINPUT34), .B(n805), .ZN(n810) );
  NAND2_X1 U895 ( .A1(n893), .A2(G128), .ZN(n807) );
  NAND2_X1 U896 ( .A1(G116), .A2(n894), .ZN(n806) );
  NAND2_X1 U897 ( .A1(n807), .A2(n806), .ZN(n808) );
  XOR2_X1 U898 ( .A(KEYINPUT35), .B(n808), .Z(n809) );
  NOR2_X1 U899 ( .A1(n810), .A2(n809), .ZN(n811) );
  XNOR2_X1 U900 ( .A(KEYINPUT36), .B(n811), .ZN(n887) );
  NOR2_X1 U901 ( .A1(n825), .A2(n887), .ZN(n929) );
  NAND2_X1 U902 ( .A1(n828), .A2(n929), .ZN(n823) );
  NAND2_X1 U903 ( .A1(n813), .A2(n516), .ZN(n815) );
  INV_X1 U904 ( .A(KEYINPUT99), .ZN(n814) );
  XNOR2_X1 U905 ( .A(n815), .B(n814), .ZN(n830) );
  NOR2_X1 U906 ( .A1(G1996), .A2(n905), .ZN(n917) );
  INV_X1 U907 ( .A(n816), .ZN(n925) );
  NOR2_X1 U908 ( .A1(G1991), .A2(n892), .ZN(n922) );
  NOR2_X1 U909 ( .A1(G1986), .A2(G290), .ZN(n817) );
  NOR2_X1 U910 ( .A1(n922), .A2(n817), .ZN(n818) );
  XNOR2_X1 U911 ( .A(n818), .B(KEYINPUT100), .ZN(n819) );
  NOR2_X1 U912 ( .A1(n925), .A2(n819), .ZN(n820) );
  XOR2_X1 U913 ( .A(KEYINPUT101), .B(n820), .Z(n821) );
  NOR2_X1 U914 ( .A1(n917), .A2(n821), .ZN(n822) );
  XNOR2_X1 U915 ( .A(n822), .B(KEYINPUT39), .ZN(n824) );
  NAND2_X1 U916 ( .A1(n824), .A2(n823), .ZN(n826) );
  NAND2_X1 U917 ( .A1(n825), .A2(n887), .ZN(n938) );
  NAND2_X1 U918 ( .A1(n826), .A2(n938), .ZN(n827) );
  NAND2_X1 U919 ( .A1(n828), .A2(n827), .ZN(n829) );
  NAND2_X1 U920 ( .A1(n830), .A2(n829), .ZN(n831) );
  XNOR2_X1 U921 ( .A(n831), .B(KEYINPUT40), .ZN(G329) );
  INV_X1 U922 ( .A(G301), .ZN(G171) );
  NAND2_X1 U923 ( .A1(n832), .A2(G2106), .ZN(n833) );
  XOR2_X1 U924 ( .A(KEYINPUT103), .B(n833), .Z(G217) );
  AND2_X1 U925 ( .A1(G15), .A2(G2), .ZN(n834) );
  NAND2_X1 U926 ( .A1(G661), .A2(n834), .ZN(G259) );
  NAND2_X1 U927 ( .A1(G3), .A2(G1), .ZN(n835) );
  NAND2_X1 U928 ( .A1(n836), .A2(n835), .ZN(G188) );
  NOR2_X1 U930 ( .A1(n838), .A2(n837), .ZN(n839) );
  XNOR2_X1 U931 ( .A(n839), .B(KEYINPUT104), .ZN(G325) );
  XNOR2_X1 U932 ( .A(KEYINPUT105), .B(G325), .ZN(G261) );
  INV_X1 U933 ( .A(G120), .ZN(G236) );
  INV_X1 U934 ( .A(G96), .ZN(G221) );
  INV_X1 U935 ( .A(G69), .ZN(G235) );
  XNOR2_X1 U936 ( .A(n996), .B(n840), .ZN(n842) );
  XNOR2_X1 U937 ( .A(G286), .B(G171), .ZN(n841) );
  XNOR2_X1 U938 ( .A(n842), .B(n841), .ZN(n843) );
  NOR2_X1 U939 ( .A1(G37), .A2(n843), .ZN(G397) );
  XOR2_X1 U940 ( .A(G1976), .B(G1986), .Z(n845) );
  XNOR2_X1 U941 ( .A(G1996), .B(G1991), .ZN(n844) );
  XNOR2_X1 U942 ( .A(n845), .B(n844), .ZN(n855) );
  XOR2_X1 U943 ( .A(KEYINPUT111), .B(KEYINPUT110), .Z(n847) );
  XNOR2_X1 U944 ( .A(G1956), .B(KEYINPUT109), .ZN(n846) );
  XNOR2_X1 U945 ( .A(n847), .B(n846), .ZN(n851) );
  XOR2_X1 U946 ( .A(G1981), .B(G1961), .Z(n849) );
  XNOR2_X1 U947 ( .A(G1971), .B(G1966), .ZN(n848) );
  XNOR2_X1 U948 ( .A(n849), .B(n848), .ZN(n850) );
  XOR2_X1 U949 ( .A(n851), .B(n850), .Z(n853) );
  XNOR2_X1 U950 ( .A(G2474), .B(KEYINPUT41), .ZN(n852) );
  XNOR2_X1 U951 ( .A(n853), .B(n852), .ZN(n854) );
  XOR2_X1 U952 ( .A(n855), .B(n854), .Z(G229) );
  XOR2_X1 U953 ( .A(KEYINPUT106), .B(KEYINPUT42), .Z(n857) );
  XNOR2_X1 U954 ( .A(KEYINPUT108), .B(G2096), .ZN(n856) );
  XNOR2_X1 U955 ( .A(n857), .B(n856), .ZN(n858) );
  XOR2_X1 U956 ( .A(n858), .B(G2678), .Z(n860) );
  XNOR2_X1 U957 ( .A(G2067), .B(G2084), .ZN(n859) );
  XNOR2_X1 U958 ( .A(n860), .B(n859), .ZN(n864) );
  XOR2_X1 U959 ( .A(G2100), .B(G2072), .Z(n862) );
  XNOR2_X1 U960 ( .A(G2090), .B(G2078), .ZN(n861) );
  XNOR2_X1 U961 ( .A(n862), .B(n861), .ZN(n863) );
  XOR2_X1 U962 ( .A(n864), .B(n863), .Z(n866) );
  XNOR2_X1 U963 ( .A(KEYINPUT107), .B(KEYINPUT43), .ZN(n865) );
  XNOR2_X1 U964 ( .A(n866), .B(n865), .ZN(G227) );
  NAND2_X1 U965 ( .A1(G124), .A2(n893), .ZN(n867) );
  XNOR2_X1 U966 ( .A(n867), .B(KEYINPUT44), .ZN(n869) );
  NAND2_X1 U967 ( .A1(n897), .A2(G100), .ZN(n868) );
  NAND2_X1 U968 ( .A1(n869), .A2(n868), .ZN(n873) );
  NAND2_X1 U969 ( .A1(G136), .A2(n574), .ZN(n871) );
  NAND2_X1 U970 ( .A1(G112), .A2(n894), .ZN(n870) );
  NAND2_X1 U971 ( .A1(n871), .A2(n870), .ZN(n872) );
  NOR2_X1 U972 ( .A1(n873), .A2(n872), .ZN(G162) );
  XNOR2_X1 U973 ( .A(KEYINPUT113), .B(KEYINPUT114), .ZN(n878) );
  NAND2_X1 U974 ( .A1(n893), .A2(G127), .ZN(n875) );
  NAND2_X1 U975 ( .A1(G115), .A2(n894), .ZN(n874) );
  NAND2_X1 U976 ( .A1(n875), .A2(n874), .ZN(n876) );
  XNOR2_X1 U977 ( .A(n876), .B(KEYINPUT47), .ZN(n877) );
  XNOR2_X1 U978 ( .A(n878), .B(n877), .ZN(n883) );
  NAND2_X1 U979 ( .A1(G103), .A2(n897), .ZN(n880) );
  NAND2_X1 U980 ( .A1(G139), .A2(n574), .ZN(n879) );
  NAND2_X1 U981 ( .A1(n880), .A2(n879), .ZN(n881) );
  XNOR2_X1 U982 ( .A(KEYINPUT112), .B(n881), .ZN(n882) );
  NOR2_X1 U983 ( .A1(n883), .A2(n882), .ZN(n931) );
  XOR2_X1 U984 ( .A(KEYINPUT48), .B(KEYINPUT115), .Z(n885) );
  XNOR2_X1 U985 ( .A(G162), .B(KEYINPUT46), .ZN(n884) );
  XNOR2_X1 U986 ( .A(n885), .B(n884), .ZN(n886) );
  XNOR2_X1 U987 ( .A(n887), .B(n886), .ZN(n889) );
  XNOR2_X1 U988 ( .A(G160), .B(G164), .ZN(n888) );
  XNOR2_X1 U989 ( .A(n889), .B(n888), .ZN(n890) );
  XOR2_X1 U990 ( .A(n931), .B(n890), .Z(n891) );
  XNOR2_X1 U991 ( .A(n892), .B(n891), .ZN(n907) );
  NAND2_X1 U992 ( .A1(n893), .A2(G130), .ZN(n896) );
  NAND2_X1 U993 ( .A1(G118), .A2(n894), .ZN(n895) );
  NAND2_X1 U994 ( .A1(n896), .A2(n895), .ZN(n902) );
  NAND2_X1 U995 ( .A1(G106), .A2(n897), .ZN(n899) );
  NAND2_X1 U996 ( .A1(G142), .A2(n574), .ZN(n898) );
  NAND2_X1 U997 ( .A1(n899), .A2(n898), .ZN(n900) );
  XOR2_X1 U998 ( .A(n900), .B(KEYINPUT45), .Z(n901) );
  NOR2_X1 U999 ( .A1(n902), .A2(n901), .ZN(n903) );
  XNOR2_X1 U1000 ( .A(n903), .B(n919), .ZN(n904) );
  XNOR2_X1 U1001 ( .A(n905), .B(n904), .ZN(n906) );
  XNOR2_X1 U1002 ( .A(n907), .B(n906), .ZN(n908) );
  NOR2_X1 U1003 ( .A1(G37), .A2(n908), .ZN(G395) );
  NOR2_X1 U1004 ( .A1(G401), .A2(n915), .ZN(n912) );
  NOR2_X1 U1005 ( .A1(G229), .A2(G227), .ZN(n909) );
  XNOR2_X1 U1006 ( .A(KEYINPUT49), .B(n909), .ZN(n910) );
  NOR2_X1 U1007 ( .A1(G397), .A2(n910), .ZN(n911) );
  NAND2_X1 U1008 ( .A1(n912), .A2(n911), .ZN(n913) );
  NOR2_X1 U1009 ( .A1(n913), .A2(G395), .ZN(n914) );
  XNOR2_X1 U1010 ( .A(n914), .B(KEYINPUT116), .ZN(G308) );
  INV_X1 U1011 ( .A(G308), .ZN(G225) );
  INV_X1 U1012 ( .A(n915), .ZN(G319) );
  INV_X1 U1013 ( .A(G108), .ZN(G238) );
  XOR2_X1 U1014 ( .A(G2090), .B(G162), .Z(n916) );
  NOR2_X1 U1015 ( .A1(n917), .A2(n916), .ZN(n918) );
  XOR2_X1 U1016 ( .A(KEYINPUT51), .B(n918), .Z(n927) );
  XNOR2_X1 U1017 ( .A(G160), .B(G2084), .ZN(n920) );
  NAND2_X1 U1018 ( .A1(n920), .A2(n919), .ZN(n921) );
  NOR2_X1 U1019 ( .A1(n922), .A2(n921), .ZN(n923) );
  XNOR2_X1 U1020 ( .A(KEYINPUT117), .B(n923), .ZN(n924) );
  NOR2_X1 U1021 ( .A1(n925), .A2(n924), .ZN(n926) );
  NAND2_X1 U1022 ( .A1(n927), .A2(n926), .ZN(n928) );
  NOR2_X1 U1023 ( .A1(n929), .A2(n928), .ZN(n930) );
  XOR2_X1 U1024 ( .A(KEYINPUT118), .B(n930), .Z(n936) );
  XOR2_X1 U1025 ( .A(G2072), .B(n931), .Z(n933) );
  XOR2_X1 U1026 ( .A(G164), .B(G2078), .Z(n932) );
  NOR2_X1 U1027 ( .A1(n933), .A2(n932), .ZN(n934) );
  XOR2_X1 U1028 ( .A(KEYINPUT50), .B(n934), .Z(n935) );
  NOR2_X1 U1029 ( .A1(n936), .A2(n935), .ZN(n937) );
  NAND2_X1 U1030 ( .A1(n938), .A2(n937), .ZN(n939) );
  XNOR2_X1 U1031 ( .A(n939), .B(KEYINPUT119), .ZN(n940) );
  XNOR2_X1 U1032 ( .A(KEYINPUT52), .B(n940), .ZN(n942) );
  INV_X1 U1033 ( .A(KEYINPUT55), .ZN(n941) );
  NAND2_X1 U1034 ( .A1(n942), .A2(n941), .ZN(n943) );
  NAND2_X1 U1035 ( .A1(n943), .A2(G29), .ZN(n1022) );
  XOR2_X1 U1036 ( .A(G2090), .B(G35), .Z(n946) );
  XOR2_X1 U1037 ( .A(KEYINPUT54), .B(G34), .Z(n944) );
  XNOR2_X1 U1038 ( .A(n944), .B(G2084), .ZN(n945) );
  NAND2_X1 U1039 ( .A1(n946), .A2(n945), .ZN(n960) );
  XOR2_X1 U1040 ( .A(G1991), .B(G25), .Z(n947) );
  NAND2_X1 U1041 ( .A1(n947), .A2(G28), .ZN(n956) );
  XNOR2_X1 U1042 ( .A(G1996), .B(G32), .ZN(n949) );
  XNOR2_X1 U1043 ( .A(G33), .B(G2072), .ZN(n948) );
  NOR2_X1 U1044 ( .A1(n949), .A2(n948), .ZN(n954) );
  XNOR2_X1 U1045 ( .A(G2067), .B(G26), .ZN(n952) );
  XNOR2_X1 U1046 ( .A(G27), .B(n950), .ZN(n951) );
  NOR2_X1 U1047 ( .A1(n952), .A2(n951), .ZN(n953) );
  NAND2_X1 U1048 ( .A1(n954), .A2(n953), .ZN(n955) );
  NOR2_X1 U1049 ( .A1(n956), .A2(n955), .ZN(n957) );
  XNOR2_X1 U1050 ( .A(KEYINPUT53), .B(n957), .ZN(n958) );
  XNOR2_X1 U1051 ( .A(KEYINPUT120), .B(n958), .ZN(n959) );
  NOR2_X1 U1052 ( .A1(n960), .A2(n959), .ZN(n961) );
  XOR2_X1 U1053 ( .A(KEYINPUT55), .B(n961), .Z(n962) );
  NOR2_X1 U1054 ( .A1(G29), .A2(n962), .ZN(n963) );
  XNOR2_X1 U1055 ( .A(KEYINPUT121), .B(n963), .ZN(n964) );
  NAND2_X1 U1056 ( .A1(n964), .A2(G11), .ZN(n1020) );
  XNOR2_X1 U1057 ( .A(KEYINPUT123), .B(G16), .ZN(n992) );
  XNOR2_X1 U1058 ( .A(G1341), .B(G19), .ZN(n965) );
  XNOR2_X1 U1059 ( .A(n965), .B(KEYINPUT124), .ZN(n967) );
  XNOR2_X1 U1060 ( .A(G6), .B(G1981), .ZN(n966) );
  NOR2_X1 U1061 ( .A1(n967), .A2(n966), .ZN(n968) );
  XOR2_X1 U1062 ( .A(KEYINPUT125), .B(n968), .Z(n972) );
  XNOR2_X1 U1063 ( .A(KEYINPUT59), .B(G4), .ZN(n969) );
  XNOR2_X1 U1064 ( .A(n969), .B(KEYINPUT126), .ZN(n970) );
  XNOR2_X1 U1065 ( .A(G1348), .B(n970), .ZN(n971) );
  NAND2_X1 U1066 ( .A1(n972), .A2(n971), .ZN(n975) );
  XNOR2_X1 U1067 ( .A(G20), .B(n973), .ZN(n974) );
  NOR2_X1 U1068 ( .A1(n975), .A2(n974), .ZN(n976) );
  XNOR2_X1 U1069 ( .A(KEYINPUT60), .B(n976), .ZN(n981) );
  XNOR2_X1 U1070 ( .A(G1966), .B(G21), .ZN(n979) );
  XNOR2_X1 U1071 ( .A(n977), .B(G5), .ZN(n978) );
  NOR2_X1 U1072 ( .A1(n979), .A2(n978), .ZN(n980) );
  NAND2_X1 U1073 ( .A1(n981), .A2(n980), .ZN(n989) );
  XNOR2_X1 U1074 ( .A(G1986), .B(G24), .ZN(n983) );
  XNOR2_X1 U1075 ( .A(G22), .B(G1971), .ZN(n982) );
  NOR2_X1 U1076 ( .A1(n983), .A2(n982), .ZN(n986) );
  XNOR2_X1 U1077 ( .A(G1976), .B(KEYINPUT127), .ZN(n984) );
  XNOR2_X1 U1078 ( .A(n984), .B(G23), .ZN(n985) );
  NAND2_X1 U1079 ( .A1(n986), .A2(n985), .ZN(n987) );
  XNOR2_X1 U1080 ( .A(KEYINPUT58), .B(n987), .ZN(n988) );
  NOR2_X1 U1081 ( .A1(n989), .A2(n988), .ZN(n990) );
  XNOR2_X1 U1082 ( .A(KEYINPUT61), .B(n990), .ZN(n991) );
  NAND2_X1 U1083 ( .A1(n992), .A2(n991), .ZN(n1018) );
  XNOR2_X1 U1084 ( .A(KEYINPUT56), .B(G16), .ZN(n1016) );
  XNOR2_X1 U1085 ( .A(G168), .B(G1966), .ZN(n994) );
  NAND2_X1 U1086 ( .A1(n994), .A2(n993), .ZN(n995) );
  XNOR2_X1 U1087 ( .A(n995), .B(KEYINPUT57), .ZN(n1000) );
  XOR2_X1 U1088 ( .A(G1348), .B(n996), .Z(n998) );
  XOR2_X1 U1089 ( .A(G171), .B(G1961), .Z(n997) );
  NOR2_X1 U1090 ( .A1(n998), .A2(n997), .ZN(n999) );
  NAND2_X1 U1091 ( .A1(n1000), .A2(n999), .ZN(n1003) );
  XNOR2_X1 U1092 ( .A(G1341), .B(n1001), .ZN(n1002) );
  NOR2_X1 U1093 ( .A1(n1003), .A2(n1002), .ZN(n1014) );
  NAND2_X1 U1094 ( .A1(G1971), .A2(G303), .ZN(n1004) );
  NAND2_X1 U1095 ( .A1(n1005), .A2(n1004), .ZN(n1009) );
  XOR2_X1 U1096 ( .A(G1956), .B(G299), .Z(n1006) );
  NAND2_X1 U1097 ( .A1(n1007), .A2(n1006), .ZN(n1008) );
  NOR2_X1 U1098 ( .A1(n1009), .A2(n1008), .ZN(n1011) );
  NAND2_X1 U1099 ( .A1(n1011), .A2(n1010), .ZN(n1012) );
  XOR2_X1 U1100 ( .A(KEYINPUT122), .B(n1012), .Z(n1013) );
  NAND2_X1 U1101 ( .A1(n1014), .A2(n1013), .ZN(n1015) );
  NAND2_X1 U1102 ( .A1(n1016), .A2(n1015), .ZN(n1017) );
  NAND2_X1 U1103 ( .A1(n1018), .A2(n1017), .ZN(n1019) );
  NOR2_X1 U1104 ( .A1(n1020), .A2(n1019), .ZN(n1021) );
  NAND2_X1 U1105 ( .A1(n1022), .A2(n1021), .ZN(n1023) );
  XOR2_X1 U1106 ( .A(KEYINPUT62), .B(n1023), .Z(G311) );
  INV_X1 U1107 ( .A(G311), .ZN(G150) );
endmodule

