//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 1 0 0 0 0 1 0 0 0 0 1 0 1 0 0 0 1 1 0 1 0 0 1 0 1 0 0 0 1 0 0 0 1 0 1 0 0 1 0 1 0 0 1 1 1 0 0 0 1 1 1 0 1 1 1 0 0 0 1 0 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:21:34 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n677, new_n678,
    new_n679, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n726, new_n727, new_n728, new_n729, new_n730, new_n731,
    new_n732, new_n733, new_n734, new_n735, new_n736, new_n737, new_n738,
    new_n739, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n759, new_n760, new_n761,
    new_n763, new_n764, new_n765, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n780, new_n781, new_n782, new_n783, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n807, new_n808,
    new_n809, new_n810, new_n811, new_n812, new_n813, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n969, new_n970, new_n971, new_n972, new_n973,
    new_n974, new_n975, new_n976, new_n977, new_n978, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1014, new_n1015, new_n1016,
    new_n1017, new_n1018, new_n1019, new_n1020, new_n1021, new_n1022,
    new_n1024, new_n1025, new_n1026, new_n1028, new_n1029, new_n1030,
    new_n1031, new_n1032, new_n1033, new_n1034, new_n1035, new_n1036,
    new_n1037, new_n1038, new_n1039, new_n1040, new_n1041, new_n1042,
    new_n1043, new_n1044, new_n1045, new_n1046, new_n1047, new_n1048,
    new_n1049, new_n1050, new_n1052, new_n1053, new_n1054, new_n1055,
    new_n1056, new_n1057, new_n1058, new_n1059, new_n1060, new_n1061,
    new_n1062, new_n1063, new_n1064;
  XOR2_X1   g000(.A(G119), .B(G128), .Z(new_n187));
  XNOR2_X1  g001(.A(KEYINPUT24), .B(G110), .ZN(new_n188));
  NOR2_X1   g002(.A1(new_n187), .A2(new_n188), .ZN(new_n189));
  INV_X1    g003(.A(G128), .ZN(new_n190));
  AOI21_X1  g004(.A(KEYINPUT72), .B1(new_n190), .B2(G119), .ZN(new_n191));
  INV_X1    g005(.A(KEYINPUT23), .ZN(new_n192));
  OR2_X1    g006(.A1(new_n191), .A2(new_n192), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n191), .A2(new_n192), .ZN(new_n194));
  OAI211_X1 g008(.A(new_n193), .B(new_n194), .C1(G119), .C2(new_n190), .ZN(new_n195));
  AOI21_X1  g009(.A(new_n189), .B1(new_n195), .B2(G110), .ZN(new_n196));
  INV_X1    g010(.A(new_n196), .ZN(new_n197));
  XNOR2_X1  g011(.A(KEYINPUT73), .B(G125), .ZN(new_n198));
  NOR3_X1   g012(.A1(new_n198), .A2(KEYINPUT16), .A3(G140), .ZN(new_n199));
  INV_X1    g013(.A(new_n199), .ZN(new_n200));
  INV_X1    g014(.A(G140), .ZN(new_n201));
  INV_X1    g015(.A(G125), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n202), .A2(KEYINPUT73), .ZN(new_n203));
  INV_X1    g017(.A(KEYINPUT73), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n204), .A2(G125), .ZN(new_n205));
  AOI21_X1  g019(.A(new_n201), .B1(new_n203), .B2(new_n205), .ZN(new_n206));
  NOR2_X1   g020(.A1(G125), .A2(G140), .ZN(new_n207));
  OAI211_X1 g021(.A(KEYINPUT74), .B(KEYINPUT16), .C1(new_n206), .C2(new_n207), .ZN(new_n208));
  INV_X1    g022(.A(new_n208), .ZN(new_n209));
  INV_X1    g023(.A(new_n207), .ZN(new_n210));
  OAI21_X1  g024(.A(new_n210), .B1(new_n198), .B2(new_n201), .ZN(new_n211));
  AOI21_X1  g025(.A(KEYINPUT74), .B1(new_n211), .B2(KEYINPUT16), .ZN(new_n212));
  OAI21_X1  g026(.A(new_n200), .B1(new_n209), .B2(new_n212), .ZN(new_n213));
  INV_X1    g027(.A(G146), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n213), .A2(new_n214), .ZN(new_n215));
  INV_X1    g029(.A(KEYINPUT74), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n203), .A2(new_n205), .ZN(new_n217));
  AOI21_X1  g031(.A(new_n207), .B1(new_n217), .B2(G140), .ZN(new_n218));
  INV_X1    g032(.A(KEYINPUT16), .ZN(new_n219));
  OAI21_X1  g033(.A(new_n216), .B1(new_n218), .B2(new_n219), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n220), .A2(new_n208), .ZN(new_n221));
  NAND3_X1  g035(.A1(new_n221), .A2(G146), .A3(new_n200), .ZN(new_n222));
  AOI21_X1  g036(.A(new_n197), .B1(new_n215), .B2(new_n222), .ZN(new_n223));
  AOI211_X1 g037(.A(new_n214), .B(new_n199), .C1(new_n220), .C2(new_n208), .ZN(new_n224));
  NAND2_X1  g038(.A1(new_n187), .A2(new_n188), .ZN(new_n225));
  OAI21_X1  g039(.A(new_n225), .B1(new_n195), .B2(G110), .ZN(new_n226));
  INV_X1    g040(.A(KEYINPUT75), .ZN(new_n227));
  NOR2_X1   g041(.A1(new_n202), .A2(new_n201), .ZN(new_n228));
  OAI21_X1  g042(.A(new_n227), .B1(new_n228), .B2(new_n207), .ZN(new_n229));
  NAND2_X1  g043(.A1(G125), .A2(G140), .ZN(new_n230));
  NAND3_X1  g044(.A1(new_n210), .A2(KEYINPUT75), .A3(new_n230), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n229), .A2(new_n231), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n232), .A2(new_n214), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n226), .A2(new_n233), .ZN(new_n234));
  NOR2_X1   g048(.A1(new_n224), .A2(new_n234), .ZN(new_n235));
  OAI21_X1  g049(.A(KEYINPUT76), .B1(new_n223), .B2(new_n235), .ZN(new_n236));
  INV_X1    g050(.A(G953), .ZN(new_n237));
  NAND3_X1  g051(.A1(new_n237), .A2(G221), .A3(G234), .ZN(new_n238));
  XNOR2_X1  g052(.A(new_n238), .B(KEYINPUT22), .ZN(new_n239));
  XNOR2_X1  g053(.A(new_n239), .B(G137), .ZN(new_n240));
  INV_X1    g054(.A(new_n240), .ZN(new_n241));
  AOI21_X1  g055(.A(G146), .B1(new_n221), .B2(new_n200), .ZN(new_n242));
  OAI21_X1  g056(.A(new_n196), .B1(new_n242), .B2(new_n224), .ZN(new_n243));
  INV_X1    g057(.A(KEYINPUT76), .ZN(new_n244));
  NAND3_X1  g058(.A1(new_n222), .A2(new_n233), .A3(new_n226), .ZN(new_n245));
  NAND3_X1  g059(.A1(new_n243), .A2(new_n244), .A3(new_n245), .ZN(new_n246));
  NAND3_X1  g060(.A1(new_n236), .A2(new_n241), .A3(new_n246), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n243), .A2(new_n245), .ZN(new_n248));
  NAND3_X1  g062(.A1(new_n248), .A2(KEYINPUT76), .A3(new_n240), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n247), .A2(new_n249), .ZN(new_n250));
  INV_X1    g064(.A(G902), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n250), .A2(new_n251), .ZN(new_n252));
  INV_X1    g066(.A(G217), .ZN(new_n253));
  AOI21_X1  g067(.A(new_n253), .B1(G234), .B2(new_n251), .ZN(new_n254));
  NOR2_X1   g068(.A1(new_n252), .A2(new_n254), .ZN(new_n255));
  INV_X1    g069(.A(KEYINPUT25), .ZN(new_n256));
  AOI21_X1  g070(.A(G902), .B1(new_n247), .B2(new_n249), .ZN(new_n257));
  OAI21_X1  g071(.A(new_n256), .B1(new_n257), .B2(KEYINPUT77), .ZN(new_n258));
  XOR2_X1   g072(.A(new_n254), .B(KEYINPUT71), .Z(new_n259));
  INV_X1    g073(.A(new_n259), .ZN(new_n260));
  AND2_X1   g074(.A1(new_n258), .A2(new_n260), .ZN(new_n261));
  INV_X1    g075(.A(KEYINPUT77), .ZN(new_n262));
  NAND3_X1  g076(.A1(new_n252), .A2(new_n262), .A3(KEYINPUT25), .ZN(new_n263));
  AOI21_X1  g077(.A(new_n255), .B1(new_n261), .B2(new_n263), .ZN(new_n264));
  INV_X1    g078(.A(G143), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n265), .A2(G146), .ZN(new_n266));
  NAND2_X1  g080(.A1(new_n214), .A2(G143), .ZN(new_n267));
  AND4_X1   g081(.A1(KEYINPUT0), .A2(new_n266), .A3(new_n267), .A4(G128), .ZN(new_n268));
  INV_X1    g082(.A(KEYINPUT64), .ZN(new_n269));
  XNOR2_X1  g083(.A(G143), .B(G146), .ZN(new_n270));
  XNOR2_X1  g084(.A(KEYINPUT0), .B(G128), .ZN(new_n271));
  OAI21_X1  g085(.A(new_n269), .B1(new_n270), .B2(new_n271), .ZN(new_n272));
  NAND2_X1  g086(.A1(new_n266), .A2(new_n267), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n190), .A2(KEYINPUT0), .ZN(new_n274));
  INV_X1    g088(.A(KEYINPUT0), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n275), .A2(G128), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n274), .A2(new_n276), .ZN(new_n277));
  NAND3_X1  g091(.A1(new_n273), .A2(new_n277), .A3(KEYINPUT64), .ZN(new_n278));
  AOI21_X1  g092(.A(new_n268), .B1(new_n272), .B2(new_n278), .ZN(new_n279));
  INV_X1    g093(.A(G131), .ZN(new_n280));
  INV_X1    g094(.A(KEYINPUT67), .ZN(new_n281));
  INV_X1    g095(.A(G137), .ZN(new_n282));
  AND2_X1   g096(.A1(KEYINPUT66), .A2(G134), .ZN(new_n283));
  NOR2_X1   g097(.A1(KEYINPUT66), .A2(G134), .ZN(new_n284));
  OAI21_X1  g098(.A(new_n282), .B1(new_n283), .B2(new_n284), .ZN(new_n285));
  XNOR2_X1  g099(.A(KEYINPUT65), .B(KEYINPUT11), .ZN(new_n286));
  AOI21_X1  g100(.A(new_n281), .B1(new_n285), .B2(new_n286), .ZN(new_n287));
  NAND3_X1  g101(.A1(new_n282), .A2(KEYINPUT11), .A3(G134), .ZN(new_n288));
  INV_X1    g102(.A(KEYINPUT66), .ZN(new_n289));
  INV_X1    g103(.A(G134), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n289), .A2(new_n290), .ZN(new_n291));
  NAND2_X1  g105(.A1(KEYINPUT66), .A2(G134), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n291), .A2(new_n292), .ZN(new_n293));
  OAI21_X1  g107(.A(new_n288), .B1(new_n293), .B2(new_n282), .ZN(new_n294));
  NOR2_X1   g108(.A1(new_n287), .A2(new_n294), .ZN(new_n295));
  NAND3_X1  g109(.A1(new_n285), .A2(new_n281), .A3(new_n286), .ZN(new_n296));
  AOI21_X1  g110(.A(new_n280), .B1(new_n295), .B2(new_n296), .ZN(new_n297));
  AOI21_X1  g111(.A(G137), .B1(new_n291), .B2(new_n292), .ZN(new_n298));
  AND2_X1   g112(.A1(KEYINPUT65), .A2(KEYINPUT11), .ZN(new_n299));
  NOR2_X1   g113(.A1(KEYINPUT65), .A2(KEYINPUT11), .ZN(new_n300));
  NOR2_X1   g114(.A1(new_n299), .A2(new_n300), .ZN(new_n301));
  OAI21_X1  g115(.A(KEYINPUT67), .B1(new_n298), .B2(new_n301), .ZN(new_n302));
  INV_X1    g116(.A(new_n288), .ZN(new_n303));
  NOR2_X1   g117(.A1(new_n283), .A2(new_n284), .ZN(new_n304));
  AOI21_X1  g118(.A(new_n303), .B1(new_n304), .B2(G137), .ZN(new_n305));
  NAND4_X1  g119(.A1(new_n302), .A2(new_n296), .A3(new_n305), .A4(new_n280), .ZN(new_n306));
  INV_X1    g120(.A(new_n306), .ZN(new_n307));
  OAI21_X1  g121(.A(new_n279), .B1(new_n297), .B2(new_n307), .ZN(new_n308));
  OAI21_X1  g122(.A(new_n285), .B1(G134), .B2(new_n282), .ZN(new_n309));
  NOR2_X1   g123(.A1(new_n214), .A2(G143), .ZN(new_n310));
  AOI22_X1  g124(.A1(new_n273), .A2(new_n190), .B1(KEYINPUT1), .B2(new_n310), .ZN(new_n311));
  NOR2_X1   g125(.A1(new_n190), .A2(KEYINPUT1), .ZN(new_n312));
  NAND3_X1  g126(.A1(new_n312), .A2(new_n266), .A3(new_n267), .ZN(new_n313));
  AOI22_X1  g127(.A1(G131), .A2(new_n309), .B1(new_n311), .B2(new_n313), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n314), .A2(new_n306), .ZN(new_n315));
  NAND3_X1  g129(.A1(new_n308), .A2(KEYINPUT30), .A3(new_n315), .ZN(new_n316));
  INV_X1    g130(.A(KEYINPUT30), .ZN(new_n317));
  INV_X1    g131(.A(new_n268), .ZN(new_n318));
  NOR3_X1   g132(.A1(new_n270), .A2(new_n271), .A3(new_n269), .ZN(new_n319));
  AOI21_X1  g133(.A(KEYINPUT64), .B1(new_n273), .B2(new_n277), .ZN(new_n320));
  OAI21_X1  g134(.A(new_n318), .B1(new_n319), .B2(new_n320), .ZN(new_n321));
  NAND3_X1  g135(.A1(new_n302), .A2(new_n296), .A3(new_n305), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n322), .A2(G131), .ZN(new_n323));
  AOI21_X1  g137(.A(new_n321), .B1(new_n323), .B2(new_n306), .ZN(new_n324));
  INV_X1    g138(.A(new_n315), .ZN(new_n325));
  OAI21_X1  g139(.A(new_n317), .B1(new_n324), .B2(new_n325), .ZN(new_n326));
  XNOR2_X1  g140(.A(G116), .B(G119), .ZN(new_n327));
  INV_X1    g141(.A(new_n327), .ZN(new_n328));
  OR2_X1    g142(.A1(KEYINPUT2), .A2(G113), .ZN(new_n329));
  NAND2_X1  g143(.A1(KEYINPUT2), .A2(G113), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n329), .A2(new_n330), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n328), .A2(new_n331), .ZN(new_n332));
  NAND3_X1  g146(.A1(new_n327), .A2(new_n329), .A3(new_n330), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n332), .A2(new_n333), .ZN(new_n334));
  NAND3_X1  g148(.A1(new_n316), .A2(new_n326), .A3(new_n334), .ZN(new_n335));
  INV_X1    g149(.A(G237), .ZN(new_n336));
  NAND3_X1  g150(.A1(new_n336), .A2(new_n237), .A3(G210), .ZN(new_n337));
  XOR2_X1   g151(.A(new_n337), .B(KEYINPUT27), .Z(new_n338));
  XNOR2_X1  g152(.A(new_n338), .B(KEYINPUT26), .ZN(new_n339));
  INV_X1    g153(.A(G101), .ZN(new_n340));
  XNOR2_X1  g154(.A(new_n339), .B(new_n340), .ZN(new_n341));
  INV_X1    g155(.A(new_n341), .ZN(new_n342));
  INV_X1    g156(.A(KEYINPUT29), .ZN(new_n343));
  INV_X1    g157(.A(new_n334), .ZN(new_n344));
  NAND3_X1  g158(.A1(new_n308), .A2(new_n344), .A3(new_n315), .ZN(new_n345));
  NAND4_X1  g159(.A1(new_n335), .A2(new_n342), .A3(new_n343), .A4(new_n345), .ZN(new_n346));
  AND2_X1   g160(.A1(new_n346), .A2(new_n251), .ZN(new_n347));
  INV_X1    g161(.A(KEYINPUT28), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n345), .A2(new_n348), .ZN(new_n349));
  OAI21_X1  g163(.A(new_n334), .B1(new_n324), .B2(new_n325), .ZN(new_n350));
  INV_X1    g164(.A(KEYINPUT68), .ZN(new_n351));
  AND3_X1   g165(.A1(new_n345), .A2(new_n350), .A3(new_n351), .ZN(new_n352));
  OAI21_X1  g166(.A(KEYINPUT28), .B1(new_n350), .B2(new_n351), .ZN(new_n353));
  OAI211_X1 g167(.A(new_n343), .B(new_n349), .C1(new_n352), .C2(new_n353), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n354), .A2(new_n341), .ZN(new_n355));
  INV_X1    g169(.A(KEYINPUT70), .ZN(new_n356));
  AND3_X1   g170(.A1(new_n345), .A2(new_n356), .A3(new_n348), .ZN(new_n357));
  AOI21_X1  g171(.A(new_n356), .B1(new_n345), .B2(new_n348), .ZN(new_n358));
  NOR2_X1   g172(.A1(new_n357), .A2(new_n358), .ZN(new_n359));
  INV_X1    g173(.A(KEYINPUT69), .ZN(new_n360));
  NAND3_X1  g174(.A1(new_n345), .A2(new_n350), .A3(new_n360), .ZN(new_n361));
  NAND4_X1  g175(.A1(new_n308), .A2(KEYINPUT69), .A3(new_n344), .A4(new_n315), .ZN(new_n362));
  NAND3_X1  g176(.A1(new_n361), .A2(new_n362), .A3(KEYINPUT28), .ZN(new_n363));
  AOI21_X1  g177(.A(new_n343), .B1(new_n359), .B2(new_n363), .ZN(new_n364));
  OAI21_X1  g178(.A(new_n347), .B1(new_n355), .B2(new_n364), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n365), .A2(G472), .ZN(new_n366));
  NOR2_X1   g180(.A1(G472), .A2(G902), .ZN(new_n367));
  NAND3_X1  g181(.A1(new_n335), .A2(new_n345), .A3(new_n341), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n368), .A2(KEYINPUT31), .ZN(new_n369));
  INV_X1    g183(.A(KEYINPUT31), .ZN(new_n370));
  NAND4_X1  g184(.A1(new_n335), .A2(new_n370), .A3(new_n345), .A4(new_n341), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n369), .A2(new_n371), .ZN(new_n372));
  AOI21_X1  g186(.A(new_n344), .B1(new_n308), .B2(new_n315), .ZN(new_n373));
  AOI21_X1  g187(.A(new_n348), .B1(new_n373), .B2(KEYINPUT68), .ZN(new_n374));
  NAND3_X1  g188(.A1(new_n345), .A2(new_n350), .A3(new_n351), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n374), .A2(new_n375), .ZN(new_n376));
  AOI21_X1  g190(.A(new_n341), .B1(new_n376), .B2(new_n349), .ZN(new_n377));
  OAI21_X1  g191(.A(new_n367), .B1(new_n372), .B2(new_n377), .ZN(new_n378));
  INV_X1    g192(.A(KEYINPUT32), .ZN(new_n379));
  NAND2_X1  g193(.A1(new_n378), .A2(new_n379), .ZN(new_n380));
  AOI22_X1  g194(.A1(new_n374), .A2(new_n375), .B1(new_n348), .B2(new_n345), .ZN(new_n381));
  OAI211_X1 g195(.A(new_n369), .B(new_n371), .C1(new_n381), .C2(new_n341), .ZN(new_n382));
  NAND3_X1  g196(.A1(new_n382), .A2(KEYINPUT32), .A3(new_n367), .ZN(new_n383));
  NAND3_X1  g197(.A1(new_n366), .A2(new_n380), .A3(new_n383), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n264), .A2(new_n384), .ZN(new_n385));
  INV_X1    g199(.A(KEYINPUT78), .ZN(new_n386));
  NAND2_X1  g200(.A1(new_n385), .A2(new_n386), .ZN(new_n387));
  NAND3_X1  g201(.A1(new_n264), .A2(new_n384), .A3(KEYINPUT78), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n387), .A2(new_n388), .ZN(new_n389));
  NAND3_X1  g203(.A1(new_n321), .A2(KEYINPUT85), .A3(new_n217), .ZN(new_n390));
  INV_X1    g204(.A(KEYINPUT85), .ZN(new_n391));
  OAI21_X1  g205(.A(new_n391), .B1(new_n279), .B2(new_n198), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n273), .A2(new_n190), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n310), .A2(KEYINPUT1), .ZN(new_n394));
  NAND4_X1  g208(.A1(new_n393), .A2(new_n198), .A3(new_n313), .A4(new_n394), .ZN(new_n395));
  NAND3_X1  g209(.A1(new_n390), .A2(new_n392), .A3(new_n395), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n237), .A2(G224), .ZN(new_n397));
  XNOR2_X1  g211(.A(new_n396), .B(new_n397), .ZN(new_n398));
  XNOR2_X1  g212(.A(G110), .B(G122), .ZN(new_n399));
  XNOR2_X1  g213(.A(new_n399), .B(KEYINPUT84), .ZN(new_n400));
  INV_X1    g214(.A(KEYINPUT79), .ZN(new_n401));
  INV_X1    g215(.A(G107), .ZN(new_n402));
  NAND3_X1  g216(.A1(new_n401), .A2(new_n402), .A3(G104), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n403), .A2(KEYINPUT3), .ZN(new_n404));
  NOR2_X1   g218(.A1(new_n402), .A2(G104), .ZN(new_n405));
  INV_X1    g219(.A(new_n405), .ZN(new_n406));
  INV_X1    g220(.A(KEYINPUT3), .ZN(new_n407));
  NAND4_X1  g221(.A1(new_n401), .A2(new_n407), .A3(new_n402), .A4(G104), .ZN(new_n408));
  NAND4_X1  g222(.A1(new_n404), .A2(new_n340), .A3(new_n406), .A4(new_n408), .ZN(new_n409));
  INV_X1    g223(.A(G104), .ZN(new_n410));
  NOR2_X1   g224(.A1(new_n410), .A2(G107), .ZN(new_n411));
  OAI21_X1  g225(.A(G101), .B1(new_n411), .B2(new_n405), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n409), .A2(new_n412), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n413), .A2(KEYINPUT81), .ZN(new_n414));
  INV_X1    g228(.A(KEYINPUT81), .ZN(new_n415));
  NAND3_X1  g229(.A1(new_n409), .A2(new_n415), .A3(new_n412), .ZN(new_n416));
  NAND2_X1  g230(.A1(new_n414), .A2(new_n416), .ZN(new_n417));
  AND2_X1   g231(.A1(G116), .A2(G119), .ZN(new_n418));
  NOR2_X1   g232(.A1(G116), .A2(G119), .ZN(new_n419));
  OAI21_X1  g233(.A(KEYINPUT5), .B1(new_n418), .B2(new_n419), .ZN(new_n420));
  INV_X1    g234(.A(G116), .ZN(new_n421));
  OR3_X1    g235(.A1(new_n421), .A2(KEYINPUT5), .A3(G119), .ZN(new_n422));
  NAND3_X1  g236(.A1(new_n420), .A2(new_n422), .A3(G113), .ZN(new_n423));
  NAND3_X1  g237(.A1(new_n417), .A2(new_n333), .A3(new_n423), .ZN(new_n424));
  INV_X1    g238(.A(KEYINPUT4), .ZN(new_n425));
  INV_X1    g239(.A(new_n404), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n406), .A2(new_n408), .ZN(new_n427));
  OAI211_X1 g241(.A(new_n425), .B(G101), .C1(new_n426), .C2(new_n427), .ZN(new_n428));
  NAND2_X1  g242(.A1(new_n428), .A2(new_n334), .ZN(new_n429));
  INV_X1    g243(.A(KEYINPUT80), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n409), .A2(KEYINPUT4), .ZN(new_n431));
  NOR3_X1   g245(.A1(new_n410), .A2(KEYINPUT79), .A3(G107), .ZN(new_n432));
  AOI21_X1  g246(.A(new_n405), .B1(new_n432), .B2(new_n407), .ZN(new_n433));
  AOI21_X1  g247(.A(new_n340), .B1(new_n433), .B2(new_n404), .ZN(new_n434));
  OAI21_X1  g248(.A(new_n430), .B1(new_n431), .B2(new_n434), .ZN(new_n435));
  OAI21_X1  g249(.A(G101), .B1(new_n426), .B2(new_n427), .ZN(new_n436));
  NAND4_X1  g250(.A1(new_n436), .A2(KEYINPUT80), .A3(KEYINPUT4), .A4(new_n409), .ZN(new_n437));
  AOI21_X1  g251(.A(new_n429), .B1(new_n435), .B2(new_n437), .ZN(new_n438));
  OAI21_X1  g252(.A(new_n424), .B1(new_n438), .B2(KEYINPUT83), .ZN(new_n439));
  INV_X1    g253(.A(KEYINPUT83), .ZN(new_n440));
  AOI211_X1 g254(.A(new_n440), .B(new_n429), .C1(new_n435), .C2(new_n437), .ZN(new_n441));
  OAI21_X1  g255(.A(new_n400), .B1(new_n439), .B2(new_n441), .ZN(new_n442));
  INV_X1    g256(.A(new_n399), .ZN(new_n443));
  NOR3_X1   g257(.A1(new_n439), .A2(new_n441), .A3(new_n443), .ZN(new_n444));
  INV_X1    g258(.A(KEYINPUT6), .ZN(new_n445));
  OAI21_X1  g259(.A(new_n442), .B1(new_n444), .B2(new_n445), .ZN(new_n446));
  AND2_X1   g260(.A1(new_n435), .A2(new_n437), .ZN(new_n447));
  OAI21_X1  g261(.A(new_n440), .B1(new_n447), .B2(new_n429), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n438), .A2(KEYINPUT83), .ZN(new_n449));
  NAND3_X1  g263(.A1(new_n448), .A2(new_n449), .A3(new_n424), .ZN(new_n450));
  NAND3_X1  g264(.A1(new_n450), .A2(KEYINPUT6), .A3(new_n400), .ZN(new_n451));
  AOI21_X1  g265(.A(new_n398), .B1(new_n446), .B2(new_n451), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n423), .A2(new_n333), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n413), .A2(new_n453), .ZN(new_n454));
  NAND4_X1  g268(.A1(new_n409), .A2(new_n423), .A3(new_n333), .A4(new_n412), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n454), .A2(new_n455), .ZN(new_n456));
  XOR2_X1   g270(.A(new_n399), .B(KEYINPUT8), .Z(new_n457));
  INV_X1    g271(.A(new_n457), .ZN(new_n458));
  AOI21_X1  g272(.A(KEYINPUT86), .B1(new_n456), .B2(new_n458), .ZN(new_n459));
  INV_X1    g273(.A(KEYINPUT86), .ZN(new_n460));
  AOI211_X1 g274(.A(new_n460), .B(new_n457), .C1(new_n454), .C2(new_n455), .ZN(new_n461));
  NOR2_X1   g275(.A1(new_n459), .A2(new_n461), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n397), .A2(KEYINPUT7), .ZN(new_n463));
  INV_X1    g277(.A(new_n463), .ZN(new_n464));
  NAND4_X1  g278(.A1(new_n390), .A2(new_n392), .A3(new_n395), .A4(new_n464), .ZN(new_n465));
  NAND2_X1  g279(.A1(new_n395), .A2(KEYINPUT87), .ZN(new_n466));
  INV_X1    g280(.A(KEYINPUT87), .ZN(new_n467));
  NAND4_X1  g281(.A1(new_n311), .A2(new_n467), .A3(new_n198), .A4(new_n313), .ZN(new_n468));
  OAI211_X1 g282(.A(new_n466), .B(new_n468), .C1(new_n279), .C2(new_n198), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n469), .A2(new_n463), .ZN(new_n470));
  NAND2_X1  g284(.A1(new_n465), .A2(new_n470), .ZN(new_n471));
  OAI21_X1  g285(.A(KEYINPUT88), .B1(new_n462), .B2(new_n471), .ZN(new_n472));
  NAND4_X1  g286(.A1(new_n448), .A2(new_n449), .A3(new_n424), .A4(new_n399), .ZN(new_n473));
  AND4_X1   g287(.A1(new_n409), .A2(new_n423), .A3(new_n333), .A4(new_n412), .ZN(new_n474));
  AOI22_X1  g288(.A1(new_n409), .A2(new_n412), .B1(new_n423), .B2(new_n333), .ZN(new_n475));
  OAI21_X1  g289(.A(new_n458), .B1(new_n474), .B2(new_n475), .ZN(new_n476));
  NAND2_X1  g290(.A1(new_n476), .A2(new_n460), .ZN(new_n477));
  NAND3_X1  g291(.A1(new_n456), .A2(KEYINPUT86), .A3(new_n458), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  INV_X1    g293(.A(KEYINPUT88), .ZN(new_n480));
  NAND4_X1  g294(.A1(new_n479), .A2(new_n480), .A3(new_n465), .A4(new_n470), .ZN(new_n481));
  NAND3_X1  g295(.A1(new_n472), .A2(new_n473), .A3(new_n481), .ZN(new_n482));
  NAND2_X1  g296(.A1(new_n482), .A2(new_n251), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n483), .A2(KEYINPUT89), .ZN(new_n484));
  INV_X1    g298(.A(KEYINPUT89), .ZN(new_n485));
  NAND3_X1  g299(.A1(new_n482), .A2(new_n485), .A3(new_n251), .ZN(new_n486));
  AOI21_X1  g300(.A(new_n452), .B1(new_n484), .B2(new_n486), .ZN(new_n487));
  OAI21_X1  g301(.A(G210), .B1(G237), .B2(G902), .ZN(new_n488));
  XOR2_X1   g302(.A(new_n488), .B(KEYINPUT90), .Z(new_n489));
  INV_X1    g303(.A(new_n489), .ZN(new_n490));
  OAI21_X1  g304(.A(KEYINPUT91), .B1(new_n487), .B2(new_n490), .ZN(new_n491));
  INV_X1    g305(.A(new_n398), .ZN(new_n492));
  AOI22_X1  g306(.A1(KEYINPUT6), .A2(new_n473), .B1(new_n450), .B2(new_n400), .ZN(new_n493));
  INV_X1    g307(.A(new_n451), .ZN(new_n494));
  OAI21_X1  g308(.A(new_n492), .B1(new_n493), .B2(new_n494), .ZN(new_n495));
  AND3_X1   g309(.A1(new_n482), .A2(new_n485), .A3(new_n251), .ZN(new_n496));
  AOI21_X1  g310(.A(new_n485), .B1(new_n482), .B2(new_n251), .ZN(new_n497));
  OAI211_X1 g311(.A(new_n495), .B(new_n490), .C1(new_n496), .C2(new_n497), .ZN(new_n498));
  OAI21_X1  g312(.A(new_n495), .B1(new_n496), .B2(new_n497), .ZN(new_n499));
  INV_X1    g313(.A(KEYINPUT91), .ZN(new_n500));
  NAND3_X1  g314(.A1(new_n499), .A2(new_n500), .A3(new_n489), .ZN(new_n501));
  NAND3_X1  g315(.A1(new_n491), .A2(new_n498), .A3(new_n501), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n435), .A2(new_n437), .ZN(new_n503));
  NAND3_X1  g317(.A1(new_n503), .A2(new_n279), .A3(new_n428), .ZN(new_n504));
  INV_X1    g318(.A(KEYINPUT10), .ZN(new_n505));
  AOI21_X1  g319(.A(new_n505), .B1(new_n311), .B2(new_n313), .ZN(new_n506));
  OAI211_X1 g320(.A(new_n313), .B(new_n394), .C1(G128), .C2(new_n270), .ZN(new_n507));
  NAND3_X1  g321(.A1(new_n507), .A2(new_n409), .A3(new_n412), .ZN(new_n508));
  AOI22_X1  g322(.A1(new_n417), .A2(new_n506), .B1(new_n505), .B2(new_n508), .ZN(new_n509));
  NAND2_X1  g323(.A1(new_n323), .A2(new_n306), .ZN(new_n510));
  INV_X1    g324(.A(new_n510), .ZN(new_n511));
  NAND3_X1  g325(.A1(new_n504), .A2(new_n509), .A3(new_n511), .ZN(new_n512));
  AND3_X1   g326(.A1(new_n409), .A2(new_n415), .A3(new_n412), .ZN(new_n513));
  AOI21_X1  g327(.A(new_n415), .B1(new_n409), .B2(new_n412), .ZN(new_n514));
  OAI21_X1  g328(.A(new_n506), .B1(new_n513), .B2(new_n514), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n508), .A2(new_n505), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  NAND2_X1  g331(.A1(new_n279), .A2(new_n428), .ZN(new_n518));
  AOI21_X1  g332(.A(new_n518), .B1(new_n435), .B2(new_n437), .ZN(new_n519));
  OAI21_X1  g333(.A(new_n510), .B1(new_n517), .B2(new_n519), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n512), .A2(new_n520), .ZN(new_n521));
  XNOR2_X1  g335(.A(G110), .B(G140), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n237), .A2(G227), .ZN(new_n523));
  XOR2_X1   g337(.A(new_n522), .B(new_n523), .Z(new_n524));
  NAND2_X1  g338(.A1(new_n521), .A2(new_n524), .ZN(new_n525));
  AOI21_X1  g339(.A(new_n507), .B1(new_n409), .B2(new_n412), .ZN(new_n526));
  AOI21_X1  g340(.A(new_n526), .B1(KEYINPUT82), .B2(new_n508), .ZN(new_n527));
  AND4_X1   g341(.A1(KEYINPUT82), .A2(new_n413), .A3(new_n313), .A4(new_n311), .ZN(new_n528));
  OAI21_X1  g342(.A(new_n510), .B1(new_n527), .B2(new_n528), .ZN(new_n529));
  NAND2_X1  g343(.A1(new_n529), .A2(KEYINPUT12), .ZN(new_n530));
  INV_X1    g344(.A(new_n524), .ZN(new_n531));
  INV_X1    g345(.A(KEYINPUT12), .ZN(new_n532));
  OAI211_X1 g346(.A(new_n510), .B(new_n532), .C1(new_n527), .C2(new_n528), .ZN(new_n533));
  NAND4_X1  g347(.A1(new_n530), .A2(new_n512), .A3(new_n531), .A4(new_n533), .ZN(new_n534));
  NAND2_X1  g348(.A1(new_n525), .A2(new_n534), .ZN(new_n535));
  INV_X1    g349(.A(G469), .ZN(new_n536));
  NAND3_X1  g350(.A1(new_n535), .A2(new_n536), .A3(new_n251), .ZN(new_n537));
  NOR2_X1   g351(.A1(new_n536), .A2(new_n251), .ZN(new_n538));
  INV_X1    g352(.A(new_n538), .ZN(new_n539));
  NAND3_X1  g353(.A1(new_n530), .A2(new_n512), .A3(new_n533), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n540), .A2(new_n524), .ZN(new_n541));
  NAND3_X1  g355(.A1(new_n512), .A2(new_n520), .A3(new_n531), .ZN(new_n542));
  NAND3_X1  g356(.A1(new_n541), .A2(G469), .A3(new_n542), .ZN(new_n543));
  NAND3_X1  g357(.A1(new_n537), .A2(new_n539), .A3(new_n543), .ZN(new_n544));
  XNOR2_X1  g358(.A(KEYINPUT9), .B(G234), .ZN(new_n545));
  OAI21_X1  g359(.A(G221), .B1(new_n545), .B2(G902), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n544), .A2(new_n546), .ZN(new_n547));
  NOR2_X1   g361(.A1(G475), .A2(G902), .ZN(new_n548));
  INV_X1    g362(.A(KEYINPUT92), .ZN(new_n549));
  XNOR2_X1  g363(.A(G113), .B(G122), .ZN(new_n550));
  XNOR2_X1  g364(.A(new_n550), .B(G104), .ZN(new_n551));
  INV_X1    g365(.A(new_n551), .ZN(new_n552));
  NAND3_X1  g366(.A1(new_n336), .A2(new_n237), .A3(G214), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n553), .A2(new_n265), .ZN(new_n554));
  NAND4_X1  g368(.A1(new_n336), .A2(new_n237), .A3(G143), .A4(G214), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n556), .A2(G131), .ZN(new_n557));
  INV_X1    g371(.A(KEYINPUT17), .ZN(new_n558));
  NAND3_X1  g372(.A1(new_n554), .A2(new_n280), .A3(new_n555), .ZN(new_n559));
  NAND3_X1  g373(.A1(new_n557), .A2(new_n558), .A3(new_n559), .ZN(new_n560));
  NAND3_X1  g374(.A1(new_n556), .A2(KEYINPUT17), .A3(G131), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n560), .A2(new_n561), .ZN(new_n562));
  NOR3_X1   g376(.A1(new_n242), .A2(new_n224), .A3(new_n562), .ZN(new_n563));
  NAND2_X1  g377(.A1(KEYINPUT18), .A2(G131), .ZN(new_n564));
  XOR2_X1   g378(.A(new_n556), .B(new_n564), .Z(new_n565));
  NAND2_X1  g379(.A1(new_n218), .A2(G146), .ZN(new_n566));
  AND2_X1   g380(.A1(new_n233), .A2(new_n566), .ZN(new_n567));
  NOR2_X1   g381(.A1(new_n565), .A2(new_n567), .ZN(new_n568));
  OAI21_X1  g382(.A(new_n552), .B1(new_n563), .B2(new_n568), .ZN(new_n569));
  OAI21_X1  g383(.A(new_n551), .B1(new_n565), .B2(new_n567), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n211), .A2(KEYINPUT19), .ZN(new_n571));
  OAI21_X1  g385(.A(new_n571), .B1(KEYINPUT19), .B2(new_n232), .ZN(new_n572));
  AOI22_X1  g386(.A1(new_n572), .A2(new_n214), .B1(new_n557), .B2(new_n559), .ZN(new_n573));
  AOI21_X1  g387(.A(new_n570), .B1(new_n573), .B2(new_n222), .ZN(new_n574));
  INV_X1    g388(.A(new_n574), .ZN(new_n575));
  AOI21_X1  g389(.A(new_n549), .B1(new_n569), .B2(new_n575), .ZN(new_n576));
  INV_X1    g390(.A(new_n562), .ZN(new_n577));
  NAND3_X1  g391(.A1(new_n215), .A2(new_n222), .A3(new_n577), .ZN(new_n578));
  INV_X1    g392(.A(new_n568), .ZN(new_n579));
  AOI21_X1  g393(.A(new_n551), .B1(new_n578), .B2(new_n579), .ZN(new_n580));
  NOR3_X1   g394(.A1(new_n580), .A2(new_n574), .A3(KEYINPUT92), .ZN(new_n581));
  OAI211_X1 g395(.A(KEYINPUT20), .B(new_n548), .C1(new_n576), .C2(new_n581), .ZN(new_n582));
  NAND3_X1  g396(.A1(new_n569), .A2(new_n548), .A3(new_n575), .ZN(new_n583));
  INV_X1    g397(.A(KEYINPUT20), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n578), .A2(new_n579), .ZN(new_n586));
  NAND2_X1  g400(.A1(new_n551), .A2(KEYINPUT94), .ZN(new_n587));
  AOI21_X1  g401(.A(G902), .B1(new_n586), .B2(new_n587), .ZN(new_n588));
  OAI21_X1  g402(.A(new_n588), .B1(new_n586), .B2(new_n587), .ZN(new_n589));
  XOR2_X1   g403(.A(KEYINPUT93), .B(G475), .Z(new_n590));
  NAND2_X1  g404(.A1(new_n589), .A2(new_n590), .ZN(new_n591));
  NAND3_X1  g405(.A1(new_n582), .A2(new_n585), .A3(new_n591), .ZN(new_n592));
  INV_X1    g406(.A(G952), .ZN(new_n593));
  NOR2_X1   g407(.A1(new_n593), .A2(G953), .ZN(new_n594));
  INV_X1    g408(.A(G234), .ZN(new_n595));
  OAI21_X1  g409(.A(new_n594), .B1(new_n595), .B2(new_n336), .ZN(new_n596));
  INV_X1    g410(.A(new_n596), .ZN(new_n597));
  AOI211_X1 g411(.A(new_n251), .B(new_n237), .C1(G234), .C2(G237), .ZN(new_n598));
  XNOR2_X1  g412(.A(KEYINPUT21), .B(G898), .ZN(new_n599));
  AOI21_X1  g413(.A(new_n597), .B1(new_n598), .B2(new_n599), .ZN(new_n600));
  XOR2_X1   g414(.A(G116), .B(G122), .Z(new_n601));
  NAND2_X1  g415(.A1(new_n601), .A2(G107), .ZN(new_n602));
  XNOR2_X1  g416(.A(G116), .B(G122), .ZN(new_n603));
  NAND2_X1  g417(.A1(new_n603), .A2(new_n402), .ZN(new_n604));
  NAND2_X1  g418(.A1(new_n602), .A2(new_n604), .ZN(new_n605));
  NAND2_X1  g419(.A1(new_n265), .A2(G128), .ZN(new_n606));
  NAND2_X1  g420(.A1(new_n190), .A2(G143), .ZN(new_n607));
  NAND3_X1  g421(.A1(new_n606), .A2(new_n607), .A3(KEYINPUT13), .ZN(new_n608));
  OAI211_X1 g422(.A(new_n608), .B(G134), .C1(KEYINPUT13), .C2(new_n606), .ZN(new_n609));
  NAND3_X1  g423(.A1(new_n304), .A2(new_n606), .A3(new_n607), .ZN(new_n610));
  NAND3_X1  g424(.A1(new_n605), .A2(new_n609), .A3(new_n610), .ZN(new_n611));
  NAND2_X1  g425(.A1(new_n606), .A2(new_n607), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n612), .A2(new_n293), .ZN(new_n613));
  NAND2_X1  g427(.A1(new_n610), .A2(new_n613), .ZN(new_n614));
  NAND3_X1  g428(.A1(new_n421), .A2(KEYINPUT14), .A3(G122), .ZN(new_n615));
  OAI211_X1 g429(.A(G107), .B(new_n615), .C1(new_n601), .C2(KEYINPUT14), .ZN(new_n616));
  NAND3_X1  g430(.A1(new_n614), .A2(new_n616), .A3(new_n604), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n611), .A2(new_n617), .ZN(new_n618));
  NOR3_X1   g432(.A1(new_n545), .A2(new_n253), .A3(G953), .ZN(new_n619));
  INV_X1    g433(.A(new_n619), .ZN(new_n620));
  NOR2_X1   g434(.A1(new_n618), .A2(new_n620), .ZN(new_n621));
  AOI21_X1  g435(.A(new_n619), .B1(new_n611), .B2(new_n617), .ZN(new_n622));
  OR2_X1    g436(.A1(new_n621), .A2(new_n622), .ZN(new_n623));
  INV_X1    g437(.A(G478), .ZN(new_n624));
  OR2_X1    g438(.A1(new_n624), .A2(KEYINPUT15), .ZN(new_n625));
  NAND3_X1  g439(.A1(new_n623), .A2(new_n251), .A3(new_n625), .ZN(new_n626));
  OAI21_X1  g440(.A(new_n251), .B1(new_n621), .B2(new_n622), .ZN(new_n627));
  INV_X1    g441(.A(KEYINPUT95), .ZN(new_n628));
  NAND2_X1  g442(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  OAI211_X1 g443(.A(KEYINPUT95), .B(new_n251), .C1(new_n621), .C2(new_n622), .ZN(new_n630));
  AOI21_X1  g444(.A(new_n625), .B1(new_n629), .B2(new_n630), .ZN(new_n631));
  INV_X1    g445(.A(KEYINPUT96), .ZN(new_n632));
  OAI21_X1  g446(.A(new_n626), .B1(new_n631), .B2(new_n632), .ZN(new_n633));
  AOI211_X1 g447(.A(KEYINPUT96), .B(new_n625), .C1(new_n629), .C2(new_n630), .ZN(new_n634));
  OR2_X1    g448(.A1(new_n633), .A2(new_n634), .ZN(new_n635));
  NOR4_X1   g449(.A1(new_n547), .A2(new_n592), .A3(new_n600), .A4(new_n635), .ZN(new_n636));
  OAI21_X1  g450(.A(G214), .B1(G237), .B2(G902), .ZN(new_n637));
  NAND3_X1  g451(.A1(new_n502), .A2(new_n636), .A3(new_n637), .ZN(new_n638));
  INV_X1    g452(.A(new_n638), .ZN(new_n639));
  NAND2_X1  g453(.A1(new_n389), .A2(new_n639), .ZN(new_n640));
  XNOR2_X1  g454(.A(new_n640), .B(G101), .ZN(G3));
  INV_X1    g455(.A(new_n637), .ZN(new_n642));
  NAND2_X1  g456(.A1(new_n499), .A2(new_n489), .ZN(new_n643));
  AOI21_X1  g457(.A(new_n642), .B1(new_n643), .B2(new_n498), .ZN(new_n644));
  INV_X1    g458(.A(new_n592), .ZN(new_n645));
  XNOR2_X1  g459(.A(new_n623), .B(KEYINPUT33), .ZN(new_n646));
  NAND3_X1  g460(.A1(new_n646), .A2(G478), .A3(new_n251), .ZN(new_n647));
  AND2_X1   g461(.A1(new_n629), .A2(new_n630), .ZN(new_n648));
  OAI21_X1  g462(.A(new_n647), .B1(new_n648), .B2(G478), .ZN(new_n649));
  INV_X1    g463(.A(new_n649), .ZN(new_n650));
  NOR2_X1   g464(.A1(new_n645), .A2(new_n650), .ZN(new_n651));
  INV_X1    g465(.A(new_n600), .ZN(new_n652));
  NAND3_X1  g466(.A1(new_n644), .A2(new_n651), .A3(new_n652), .ZN(new_n653));
  INV_X1    g467(.A(G472), .ZN(new_n654));
  NOR2_X1   g468(.A1(new_n654), .A2(KEYINPUT97), .ZN(new_n655));
  INV_X1    g469(.A(new_n655), .ZN(new_n656));
  NAND3_X1  g470(.A1(new_n382), .A2(new_n251), .A3(new_n656), .ZN(new_n657));
  INV_X1    g471(.A(new_n657), .ZN(new_n658));
  AOI21_X1  g472(.A(new_n656), .B1(new_n382), .B2(new_n251), .ZN(new_n659));
  NOR2_X1   g473(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  INV_X1    g474(.A(new_n546), .ZN(new_n661));
  AOI21_X1  g475(.A(G902), .B1(new_n525), .B2(new_n534), .ZN(new_n662));
  AOI21_X1  g476(.A(new_n538), .B1(new_n662), .B2(new_n536), .ZN(new_n663));
  AOI21_X1  g477(.A(new_n661), .B1(new_n663), .B2(new_n543), .ZN(new_n664));
  NAND3_X1  g478(.A1(new_n264), .A2(new_n660), .A3(new_n664), .ZN(new_n665));
  NOR2_X1   g479(.A1(new_n653), .A2(new_n665), .ZN(new_n666));
  XNOR2_X1  g480(.A(KEYINPUT34), .B(G104), .ZN(new_n667));
  XNOR2_X1  g481(.A(new_n666), .B(new_n667), .ZN(G6));
  NAND2_X1  g482(.A1(new_n582), .A2(new_n591), .ZN(new_n669));
  INV_X1    g483(.A(new_n548), .ZN(new_n670));
  NAND3_X1  g484(.A1(new_n569), .A2(new_n549), .A3(new_n575), .ZN(new_n671));
  OAI21_X1  g485(.A(KEYINPUT92), .B1(new_n580), .B2(new_n574), .ZN(new_n672));
  AOI21_X1  g486(.A(new_n670), .B1(new_n671), .B2(new_n672), .ZN(new_n673));
  NOR2_X1   g487(.A1(new_n673), .A2(KEYINPUT20), .ZN(new_n674));
  NOR2_X1   g488(.A1(new_n633), .A2(new_n634), .ZN(new_n675));
  NOR3_X1   g489(.A1(new_n669), .A2(new_n674), .A3(new_n675), .ZN(new_n676));
  NAND3_X1  g490(.A1(new_n644), .A2(new_n652), .A3(new_n676), .ZN(new_n677));
  NOR2_X1   g491(.A1(new_n677), .A2(new_n665), .ZN(new_n678));
  XNOR2_X1  g492(.A(KEYINPUT35), .B(G107), .ZN(new_n679));
  XNOR2_X1  g493(.A(new_n678), .B(new_n679), .ZN(G9));
  NAND3_X1  g494(.A1(new_n263), .A2(new_n258), .A3(new_n260), .ZN(new_n681));
  NOR2_X1   g495(.A1(new_n241), .A2(KEYINPUT36), .ZN(new_n682));
  XNOR2_X1  g496(.A(new_n248), .B(new_n682), .ZN(new_n683));
  OAI211_X1 g497(.A(new_n683), .B(new_n251), .C1(new_n253), .C2(G234), .ZN(new_n684));
  NAND2_X1  g498(.A1(new_n681), .A2(new_n684), .ZN(new_n685));
  INV_X1    g499(.A(KEYINPUT98), .ZN(new_n686));
  NAND2_X1  g500(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  NAND3_X1  g501(.A1(new_n681), .A2(KEYINPUT98), .A3(new_n684), .ZN(new_n688));
  NAND3_X1  g502(.A1(new_n687), .A2(new_n660), .A3(new_n688), .ZN(new_n689));
  NOR2_X1   g503(.A1(new_n638), .A2(new_n689), .ZN(new_n690));
  XNOR2_X1  g504(.A(KEYINPUT37), .B(G110), .ZN(new_n691));
  XNOR2_X1  g505(.A(new_n690), .B(new_n691), .ZN(G12));
  NAND3_X1  g506(.A1(new_n687), .A2(new_n384), .A3(new_n688), .ZN(new_n693));
  AOI22_X1  g507(.A1(new_n673), .A2(KEYINPUT20), .B1(new_n589), .B2(new_n590), .ZN(new_n694));
  NAND2_X1  g508(.A1(new_n671), .A2(new_n672), .ZN(new_n695));
  NAND2_X1  g509(.A1(new_n695), .A2(new_n548), .ZN(new_n696));
  NAND2_X1  g510(.A1(new_n696), .A2(new_n584), .ZN(new_n697));
  INV_X1    g511(.A(G900), .ZN(new_n698));
  NAND2_X1  g512(.A1(new_n598), .A2(new_n698), .ZN(new_n699));
  NAND2_X1  g513(.A1(new_n699), .A2(new_n596), .ZN(new_n700));
  NAND4_X1  g514(.A1(new_n694), .A2(new_n635), .A3(new_n697), .A4(new_n700), .ZN(new_n701));
  INV_X1    g515(.A(new_n701), .ZN(new_n702));
  NAND3_X1  g516(.A1(new_n644), .A2(new_n664), .A3(new_n702), .ZN(new_n703));
  NOR2_X1   g517(.A1(new_n693), .A2(new_n703), .ZN(new_n704));
  XNOR2_X1  g518(.A(new_n704), .B(new_n190), .ZN(G30));
  OR2_X1    g519(.A1(new_n502), .A2(KEYINPUT38), .ZN(new_n706));
  NAND2_X1  g520(.A1(new_n502), .A2(KEYINPUT38), .ZN(new_n707));
  NAND2_X1  g521(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  XNOR2_X1  g522(.A(new_n700), .B(KEYINPUT99), .ZN(new_n709));
  XNOR2_X1  g523(.A(new_n709), .B(KEYINPUT39), .ZN(new_n710));
  NOR2_X1   g524(.A1(new_n547), .A2(new_n710), .ZN(new_n711));
  XNOR2_X1  g525(.A(new_n711), .B(KEYINPUT40), .ZN(new_n712));
  AND3_X1   g526(.A1(new_n382), .A2(KEYINPUT32), .A3(new_n367), .ZN(new_n713));
  AOI21_X1  g527(.A(KEYINPUT32), .B1(new_n382), .B2(new_n367), .ZN(new_n714));
  NOR2_X1   g528(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  NAND2_X1  g529(.A1(new_n335), .A2(new_n345), .ZN(new_n716));
  NAND2_X1  g530(.A1(new_n716), .A2(new_n341), .ZN(new_n717));
  NAND2_X1  g531(.A1(new_n717), .A2(new_n251), .ZN(new_n718));
  AOI21_X1  g532(.A(new_n341), .B1(new_n361), .B2(new_n362), .ZN(new_n719));
  OAI21_X1  g533(.A(G472), .B1(new_n718), .B2(new_n719), .ZN(new_n720));
  AOI21_X1  g534(.A(new_n685), .B1(new_n715), .B2(new_n720), .ZN(new_n721));
  NOR2_X1   g535(.A1(new_n645), .A2(new_n675), .ZN(new_n722));
  AND3_X1   g536(.A1(new_n721), .A2(new_n637), .A3(new_n722), .ZN(new_n723));
  NAND3_X1  g537(.A1(new_n708), .A2(new_n712), .A3(new_n723), .ZN(new_n724));
  XNOR2_X1  g538(.A(new_n724), .B(G143), .ZN(G45));
  AND3_X1   g539(.A1(new_n687), .A2(new_n384), .A3(new_n688), .ZN(new_n726));
  NAND2_X1  g540(.A1(new_n643), .A2(new_n498), .ZN(new_n727));
  NAND3_X1  g541(.A1(new_n727), .A2(new_n637), .A3(new_n664), .ZN(new_n728));
  NAND3_X1  g542(.A1(new_n592), .A2(new_n649), .A3(new_n700), .ZN(new_n729));
  NAND2_X1  g543(.A1(new_n729), .A2(KEYINPUT100), .ZN(new_n730));
  INV_X1    g544(.A(KEYINPUT100), .ZN(new_n731));
  NAND4_X1  g545(.A1(new_n592), .A2(new_n649), .A3(new_n731), .A4(new_n700), .ZN(new_n732));
  NAND2_X1  g546(.A1(new_n730), .A2(new_n732), .ZN(new_n733));
  NOR2_X1   g547(.A1(new_n728), .A2(new_n733), .ZN(new_n734));
  NAND3_X1  g548(.A1(new_n726), .A2(new_n734), .A3(KEYINPUT101), .ZN(new_n735));
  INV_X1    g549(.A(KEYINPUT101), .ZN(new_n736));
  NAND4_X1  g550(.A1(new_n644), .A2(new_n664), .A3(new_n732), .A4(new_n730), .ZN(new_n737));
  OAI21_X1  g551(.A(new_n736), .B1(new_n737), .B2(new_n693), .ZN(new_n738));
  NAND2_X1  g552(.A1(new_n735), .A2(new_n738), .ZN(new_n739));
  XNOR2_X1  g553(.A(new_n739), .B(G146), .ZN(G48));
  INV_X1    g554(.A(new_n653), .ZN(new_n741));
  INV_X1    g555(.A(KEYINPUT103), .ZN(new_n742));
  INV_X1    g556(.A(new_n255), .ZN(new_n743));
  NAND2_X1  g557(.A1(new_n681), .A2(new_n743), .ZN(new_n744));
  AOI21_X1  g558(.A(new_n744), .B1(new_n715), .B2(new_n366), .ZN(new_n745));
  NOR2_X1   g559(.A1(new_n662), .A2(new_n536), .ZN(new_n746));
  AOI211_X1 g560(.A(G469), .B(G902), .C1(new_n525), .C2(new_n534), .ZN(new_n747));
  NOR2_X1   g561(.A1(new_n746), .A2(new_n747), .ZN(new_n748));
  AOI21_X1  g562(.A(KEYINPUT102), .B1(new_n748), .B2(new_n546), .ZN(new_n749));
  INV_X1    g563(.A(KEYINPUT102), .ZN(new_n750));
  NOR4_X1   g564(.A1(new_n746), .A2(new_n747), .A3(new_n750), .A4(new_n661), .ZN(new_n751));
  NOR2_X1   g565(.A1(new_n749), .A2(new_n751), .ZN(new_n752));
  NAND4_X1  g566(.A1(new_n741), .A2(new_n742), .A3(new_n745), .A4(new_n752), .ZN(new_n753));
  NAND3_X1  g567(.A1(new_n752), .A2(new_n384), .A3(new_n264), .ZN(new_n754));
  OAI21_X1  g568(.A(KEYINPUT103), .B1(new_n754), .B2(new_n653), .ZN(new_n755));
  NAND2_X1  g569(.A1(new_n753), .A2(new_n755), .ZN(new_n756));
  XNOR2_X1  g570(.A(new_n756), .B(KEYINPUT41), .ZN(new_n757));
  XNOR2_X1  g571(.A(new_n757), .B(G113), .ZN(G15));
  AOI211_X1 g572(.A(new_n642), .B(new_n600), .C1(new_n643), .C2(new_n498), .ZN(new_n759));
  NAND4_X1  g573(.A1(new_n745), .A2(new_n759), .A3(new_n676), .A4(new_n752), .ZN(new_n760));
  XOR2_X1   g574(.A(KEYINPUT104), .B(G116), .Z(new_n761));
  XNOR2_X1  g575(.A(new_n760), .B(new_n761), .ZN(G18));
  NOR3_X1   g576(.A1(new_n592), .A2(new_n635), .A3(new_n600), .ZN(new_n763));
  NAND3_X1  g577(.A1(new_n752), .A2(new_n763), .A3(new_n644), .ZN(new_n764));
  NOR2_X1   g578(.A1(new_n764), .A2(new_n693), .ZN(new_n765));
  XOR2_X1   g579(.A(new_n765), .B(G119), .Z(G21));
  AND3_X1   g580(.A1(new_n727), .A2(new_n637), .A3(new_n722), .ZN(new_n767));
  AOI21_X1  g581(.A(new_n341), .B1(new_n359), .B2(new_n363), .ZN(new_n768));
  OAI21_X1  g582(.A(new_n367), .B1(new_n372), .B2(new_n768), .ZN(new_n769));
  INV_X1    g583(.A(KEYINPUT105), .ZN(new_n770));
  NAND2_X1  g584(.A1(new_n769), .A2(new_n770), .ZN(new_n771));
  OAI21_X1  g585(.A(new_n251), .B1(new_n372), .B2(new_n377), .ZN(new_n772));
  NAND2_X1  g586(.A1(new_n772), .A2(G472), .ZN(new_n773));
  OAI211_X1 g587(.A(KEYINPUT105), .B(new_n367), .C1(new_n372), .C2(new_n768), .ZN(new_n774));
  NAND3_X1  g588(.A1(new_n771), .A2(new_n773), .A3(new_n774), .ZN(new_n775));
  NOR2_X1   g589(.A1(new_n775), .A2(new_n744), .ZN(new_n776));
  NOR3_X1   g590(.A1(new_n749), .A2(new_n751), .A3(new_n600), .ZN(new_n777));
  NAND3_X1  g591(.A1(new_n767), .A2(new_n776), .A3(new_n777), .ZN(new_n778));
  XNOR2_X1  g592(.A(new_n778), .B(G122), .ZN(G24));
  INV_X1    g593(.A(new_n775), .ZN(new_n780));
  NAND4_X1  g594(.A1(new_n780), .A2(new_n685), .A3(new_n732), .A4(new_n730), .ZN(new_n781));
  NAND2_X1  g595(.A1(new_n752), .A2(new_n644), .ZN(new_n782));
  NOR2_X1   g596(.A1(new_n781), .A2(new_n782), .ZN(new_n783));
  XNOR2_X1  g597(.A(new_n783), .B(new_n202), .ZN(G27));
  AOI21_X1  g598(.A(new_n642), .B1(new_n487), .B2(new_n490), .ZN(new_n785));
  NAND2_X1  g599(.A1(new_n541), .A2(new_n542), .ZN(new_n786));
  INV_X1    g600(.A(KEYINPUT106), .ZN(new_n787));
  NAND2_X1  g601(.A1(new_n786), .A2(new_n787), .ZN(new_n788));
  NAND2_X1  g602(.A1(new_n542), .A2(KEYINPUT106), .ZN(new_n789));
  NAND3_X1  g603(.A1(new_n788), .A2(G469), .A3(new_n789), .ZN(new_n790));
  AOI21_X1  g604(.A(new_n661), .B1(new_n790), .B2(new_n663), .ZN(new_n791));
  AND4_X1   g605(.A1(new_n491), .A2(new_n785), .A3(new_n501), .A4(new_n791), .ZN(new_n792));
  AND3_X1   g606(.A1(new_n730), .A2(KEYINPUT42), .A3(new_n732), .ZN(new_n793));
  INV_X1    g607(.A(KEYINPUT107), .ZN(new_n794));
  OAI21_X1  g608(.A(new_n794), .B1(new_n713), .B2(new_n714), .ZN(new_n795));
  NAND3_X1  g609(.A1(new_n380), .A2(KEYINPUT107), .A3(new_n383), .ZN(new_n796));
  NAND3_X1  g610(.A1(new_n795), .A2(new_n366), .A3(new_n796), .ZN(new_n797));
  NAND4_X1  g611(.A1(new_n792), .A2(new_n793), .A3(new_n264), .A4(new_n797), .ZN(new_n798));
  NAND4_X1  g612(.A1(new_n491), .A2(new_n785), .A3(new_n501), .A4(new_n791), .ZN(new_n799));
  NOR3_X1   g613(.A1(new_n799), .A2(new_n385), .A3(new_n733), .ZN(new_n800));
  OAI21_X1  g614(.A(new_n798), .B1(new_n800), .B2(KEYINPUT42), .ZN(new_n801));
  INV_X1    g615(.A(KEYINPUT108), .ZN(new_n802));
  NAND2_X1  g616(.A1(new_n801), .A2(new_n802), .ZN(new_n803));
  OAI211_X1 g617(.A(new_n798), .B(KEYINPUT108), .C1(new_n800), .C2(KEYINPUT42), .ZN(new_n804));
  AND2_X1   g618(.A1(new_n803), .A2(new_n804), .ZN(new_n805));
  XNOR2_X1  g619(.A(new_n805), .B(G131), .ZN(G33));
  INV_X1    g620(.A(KEYINPUT109), .ZN(new_n807));
  XNOR2_X1  g621(.A(new_n701), .B(new_n807), .ZN(new_n808));
  NAND3_X1  g622(.A1(new_n792), .A2(new_n808), .A3(new_n745), .ZN(new_n809));
  NAND2_X1  g623(.A1(new_n809), .A2(KEYINPUT110), .ZN(new_n810));
  INV_X1    g624(.A(KEYINPUT110), .ZN(new_n811));
  NAND4_X1  g625(.A1(new_n792), .A2(new_n808), .A3(new_n811), .A4(new_n745), .ZN(new_n812));
  NAND2_X1  g626(.A1(new_n810), .A2(new_n812), .ZN(new_n813));
  XNOR2_X1  g627(.A(new_n813), .B(G134), .ZN(G36));
  NAND3_X1  g628(.A1(new_n788), .A2(KEYINPUT45), .A3(new_n789), .ZN(new_n815));
  INV_X1    g629(.A(KEYINPUT45), .ZN(new_n816));
  AOI21_X1  g630(.A(new_n536), .B1(new_n786), .B2(new_n816), .ZN(new_n817));
  NAND2_X1  g631(.A1(new_n815), .A2(new_n817), .ZN(new_n818));
  NAND2_X1  g632(.A1(new_n818), .A2(new_n539), .ZN(new_n819));
  INV_X1    g633(.A(KEYINPUT46), .ZN(new_n820));
  AOI21_X1  g634(.A(new_n747), .B1(new_n819), .B2(new_n820), .ZN(new_n821));
  OAI21_X1  g635(.A(new_n821), .B1(new_n820), .B2(new_n819), .ZN(new_n822));
  NAND2_X1  g636(.A1(new_n822), .A2(new_n546), .ZN(new_n823));
  OR2_X1    g637(.A1(new_n823), .A2(new_n710), .ZN(new_n824));
  INV_X1    g638(.A(new_n824), .ZN(new_n825));
  AND3_X1   g639(.A1(new_n491), .A2(new_n785), .A3(new_n501), .ZN(new_n826));
  AOI21_X1  g640(.A(KEYINPUT111), .B1(new_n645), .B2(new_n649), .ZN(new_n827));
  XOR2_X1   g641(.A(new_n827), .B(KEYINPUT43), .Z(new_n828));
  INV_X1    g642(.A(new_n685), .ZN(new_n829));
  NOR2_X1   g643(.A1(new_n829), .A2(new_n660), .ZN(new_n830));
  NAND2_X1  g644(.A1(new_n828), .A2(new_n830), .ZN(new_n831));
  AND2_X1   g645(.A1(new_n831), .A2(KEYINPUT44), .ZN(new_n832));
  NOR2_X1   g646(.A1(new_n831), .A2(KEYINPUT44), .ZN(new_n833));
  OAI211_X1 g647(.A(new_n825), .B(new_n826), .C1(new_n832), .C2(new_n833), .ZN(new_n834));
  XNOR2_X1  g648(.A(new_n834), .B(KEYINPUT112), .ZN(new_n835));
  XNOR2_X1  g649(.A(new_n835), .B(new_n282), .ZN(G39));
  INV_X1    g650(.A(KEYINPUT47), .ZN(new_n837));
  NAND3_X1  g651(.A1(new_n822), .A2(new_n837), .A3(new_n546), .ZN(new_n838));
  INV_X1    g652(.A(new_n838), .ZN(new_n839));
  AOI21_X1  g653(.A(new_n837), .B1(new_n822), .B2(new_n546), .ZN(new_n840));
  NOR2_X1   g654(.A1(new_n839), .A2(new_n840), .ZN(new_n841));
  NOR3_X1   g655(.A1(new_n733), .A2(new_n384), .A3(new_n264), .ZN(new_n842));
  NAND3_X1  g656(.A1(new_n841), .A2(new_n826), .A3(new_n842), .ZN(new_n843));
  XNOR2_X1  g657(.A(new_n843), .B(KEYINPUT113), .ZN(new_n844));
  XNOR2_X1  g658(.A(new_n844), .B(new_n201), .ZN(G42));
  NOR3_X1   g659(.A1(new_n749), .A2(new_n751), .A3(new_n596), .ZN(new_n846));
  AND2_X1   g660(.A1(new_n826), .A2(new_n846), .ZN(new_n847));
  AND4_X1   g661(.A1(new_n264), .A2(new_n847), .A3(new_n828), .A4(new_n797), .ZN(new_n848));
  INV_X1    g662(.A(KEYINPUT48), .ZN(new_n849));
  XNOR2_X1  g663(.A(new_n848), .B(new_n849), .ZN(new_n850));
  NOR3_X1   g664(.A1(new_n775), .A2(new_n744), .A3(new_n596), .ZN(new_n851));
  NAND2_X1  g665(.A1(new_n828), .A2(new_n851), .ZN(new_n852));
  OAI21_X1  g666(.A(new_n594), .B1(new_n852), .B2(new_n782), .ZN(new_n853));
  NAND3_X1  g667(.A1(new_n380), .A2(new_n383), .A3(new_n720), .ZN(new_n854));
  NOR2_X1   g668(.A1(new_n854), .A2(new_n744), .ZN(new_n855));
  AND3_X1   g669(.A1(new_n847), .A2(new_n651), .A3(new_n855), .ZN(new_n856));
  OR3_X1    g670(.A1(new_n853), .A2(KEYINPUT124), .A3(new_n856), .ZN(new_n857));
  OAI21_X1  g671(.A(KEYINPUT124), .B1(new_n853), .B2(new_n856), .ZN(new_n858));
  AND3_X1   g672(.A1(new_n850), .A2(new_n857), .A3(new_n858), .ZN(new_n859));
  INV_X1    g673(.A(KEYINPUT121), .ZN(new_n860));
  NAND4_X1  g674(.A1(new_n828), .A2(new_n851), .A3(new_n707), .A4(new_n706), .ZN(new_n861));
  NAND2_X1  g675(.A1(new_n752), .A2(new_n642), .ZN(new_n862));
  XNOR2_X1  g676(.A(new_n862), .B(KEYINPUT120), .ZN(new_n863));
  OAI21_X1  g677(.A(new_n860), .B1(new_n861), .B2(new_n863), .ZN(new_n864));
  INV_X1    g678(.A(KEYINPUT50), .ZN(new_n865));
  OR2_X1    g679(.A1(new_n864), .A2(new_n865), .ZN(new_n866));
  NAND4_X1  g680(.A1(new_n847), .A2(new_n828), .A3(new_n685), .A4(new_n780), .ZN(new_n867));
  NAND4_X1  g681(.A1(new_n847), .A2(new_n645), .A3(new_n650), .A4(new_n855), .ZN(new_n868));
  NAND2_X1  g682(.A1(new_n867), .A2(new_n868), .ZN(new_n869));
  XNOR2_X1  g683(.A(new_n748), .B(KEYINPUT114), .ZN(new_n870));
  INV_X1    g684(.A(KEYINPUT119), .ZN(new_n871));
  AOI21_X1  g685(.A(new_n546), .B1(new_n870), .B2(new_n871), .ZN(new_n872));
  OAI21_X1  g686(.A(new_n872), .B1(new_n871), .B2(new_n870), .ZN(new_n873));
  OAI21_X1  g687(.A(new_n873), .B1(new_n839), .B2(new_n840), .ZN(new_n874));
  AND3_X1   g688(.A1(new_n828), .A2(new_n826), .A3(new_n851), .ZN(new_n875));
  AOI21_X1  g689(.A(new_n869), .B1(new_n874), .B2(new_n875), .ZN(new_n876));
  NAND2_X1  g690(.A1(new_n864), .A2(new_n865), .ZN(new_n877));
  AND3_X1   g691(.A1(new_n866), .A2(new_n876), .A3(new_n877), .ZN(new_n878));
  OAI21_X1  g692(.A(new_n859), .B1(new_n878), .B2(KEYINPUT51), .ZN(new_n879));
  XNOR2_X1  g693(.A(new_n869), .B(KEYINPUT122), .ZN(new_n880));
  NAND3_X1  g694(.A1(new_n880), .A2(new_n866), .A3(new_n877), .ZN(new_n881));
  NAND2_X1  g695(.A1(new_n881), .A2(KEYINPUT123), .ZN(new_n882));
  INV_X1    g696(.A(KEYINPUT123), .ZN(new_n883));
  NAND4_X1  g697(.A1(new_n880), .A2(new_n883), .A3(new_n866), .A4(new_n877), .ZN(new_n884));
  NAND2_X1  g698(.A1(new_n882), .A2(new_n884), .ZN(new_n885));
  INV_X1    g699(.A(KEYINPUT51), .ZN(new_n886));
  AOI21_X1  g700(.A(new_n886), .B1(new_n874), .B2(new_n875), .ZN(new_n887));
  AOI21_X1  g701(.A(new_n879), .B1(new_n885), .B2(new_n887), .ZN(new_n888));
  OAI22_X1  g702(.A1(new_n693), .A2(new_n764), .B1(new_n754), .B2(new_n677), .ZN(new_n889));
  INV_X1    g703(.A(new_n778), .ZN(new_n890));
  NOR2_X1   g704(.A1(new_n889), .A2(new_n890), .ZN(new_n891));
  AND3_X1   g705(.A1(new_n502), .A2(new_n637), .A3(new_n651), .ZN(new_n892));
  NAND3_X1  g706(.A1(new_n681), .A2(new_n664), .A3(new_n743), .ZN(new_n893));
  NAND2_X1  g707(.A1(new_n772), .A2(new_n655), .ZN(new_n894));
  NAND2_X1  g708(.A1(new_n894), .A2(new_n657), .ZN(new_n895));
  NOR3_X1   g709(.A1(new_n893), .A2(new_n895), .A3(new_n600), .ZN(new_n896));
  AOI22_X1  g710(.A1(new_n389), .A2(new_n639), .B1(new_n892), .B2(new_n896), .ZN(new_n897));
  AND3_X1   g711(.A1(new_n891), .A2(new_n897), .A3(new_n756), .ZN(new_n898));
  NOR2_X1   g712(.A1(new_n592), .A2(new_n675), .ZN(new_n899));
  NAND3_X1  g713(.A1(new_n502), .A2(new_n637), .A3(new_n899), .ZN(new_n900));
  NAND4_X1  g714(.A1(new_n264), .A2(new_n660), .A3(new_n664), .A4(new_n652), .ZN(new_n901));
  OAI22_X1  g715(.A1(new_n638), .A2(new_n689), .B1(new_n900), .B2(new_n901), .ZN(new_n902));
  INV_X1    g716(.A(KEYINPUT115), .ZN(new_n903));
  NAND2_X1  g717(.A1(new_n902), .A2(new_n903), .ZN(new_n904));
  NAND4_X1  g718(.A1(new_n896), .A2(new_n637), .A3(new_n502), .A4(new_n899), .ZN(new_n905));
  OAI211_X1 g719(.A(new_n905), .B(KEYINPUT115), .C1(new_n638), .C2(new_n689), .ZN(new_n906));
  NAND2_X1  g720(.A1(new_n904), .A2(new_n906), .ZN(new_n907));
  NOR2_X1   g721(.A1(new_n781), .A2(new_n799), .ZN(new_n908));
  INV_X1    g722(.A(new_n700), .ZN(new_n909));
  NOR3_X1   g723(.A1(new_n633), .A2(new_n634), .A3(new_n909), .ZN(new_n910));
  NAND3_X1  g724(.A1(new_n694), .A2(new_n697), .A3(new_n910), .ZN(new_n911));
  NOR2_X1   g725(.A1(new_n911), .A2(new_n547), .ZN(new_n912));
  NAND4_X1  g726(.A1(new_n912), .A2(new_n491), .A3(new_n501), .A4(new_n785), .ZN(new_n913));
  INV_X1    g727(.A(new_n913), .ZN(new_n914));
  INV_X1    g728(.A(KEYINPUT116), .ZN(new_n915));
  NAND3_X1  g729(.A1(new_n726), .A2(new_n914), .A3(new_n915), .ZN(new_n916));
  OAI21_X1  g730(.A(KEYINPUT116), .B1(new_n693), .B2(new_n913), .ZN(new_n917));
  AOI21_X1  g731(.A(new_n908), .B1(new_n916), .B2(new_n917), .ZN(new_n918));
  AND2_X1   g732(.A1(new_n918), .A2(new_n813), .ZN(new_n919));
  NAND4_X1  g733(.A1(new_n805), .A2(new_n898), .A3(new_n907), .A4(new_n919), .ZN(new_n920));
  OAI22_X1  g734(.A1(new_n781), .A2(new_n782), .B1(new_n693), .B2(new_n703), .ZN(new_n921));
  AOI21_X1  g735(.A(new_n921), .B1(new_n738), .B2(new_n735), .ZN(new_n922));
  INV_X1    g736(.A(KEYINPUT118), .ZN(new_n923));
  AOI211_X1 g737(.A(new_n661), .B(new_n909), .C1(new_n790), .C2(new_n663), .ZN(new_n924));
  NAND4_X1  g738(.A1(new_n767), .A2(new_n721), .A3(new_n923), .A4(new_n924), .ZN(new_n925));
  NAND3_X1  g739(.A1(new_n829), .A2(new_n924), .A3(new_n854), .ZN(new_n926));
  NAND2_X1  g740(.A1(new_n644), .A2(new_n722), .ZN(new_n927));
  OAI21_X1  g741(.A(KEYINPUT118), .B1(new_n926), .B2(new_n927), .ZN(new_n928));
  NAND2_X1  g742(.A1(new_n925), .A2(new_n928), .ZN(new_n929));
  AOI21_X1  g743(.A(KEYINPUT52), .B1(new_n922), .B2(new_n929), .ZN(new_n930));
  INV_X1    g744(.A(new_n921), .ZN(new_n931));
  AND4_X1   g745(.A1(KEYINPUT52), .A2(new_n739), .A3(new_n929), .A4(new_n931), .ZN(new_n932));
  NOR2_X1   g746(.A1(new_n930), .A2(new_n932), .ZN(new_n933));
  OAI21_X1  g747(.A(KEYINPUT53), .B1(new_n920), .B2(new_n933), .ZN(new_n934));
  NAND4_X1  g748(.A1(new_n896), .A2(new_n637), .A3(new_n502), .A4(new_n651), .ZN(new_n935));
  AND3_X1   g749(.A1(new_n264), .A2(new_n384), .A3(KEYINPUT78), .ZN(new_n936));
  AOI21_X1  g750(.A(KEYINPUT78), .B1(new_n264), .B2(new_n384), .ZN(new_n937));
  NOR2_X1   g751(.A1(new_n936), .A2(new_n937), .ZN(new_n938));
  OAI21_X1  g752(.A(new_n935), .B1(new_n938), .B2(new_n638), .ZN(new_n939));
  OAI211_X1 g753(.A(new_n778), .B(new_n760), .C1(new_n693), .C2(new_n764), .ZN(new_n940));
  NOR2_X1   g754(.A1(new_n939), .A2(new_n940), .ZN(new_n941));
  NAND3_X1  g755(.A1(new_n941), .A2(new_n907), .A3(new_n756), .ZN(new_n942));
  NAND4_X1  g756(.A1(new_n803), .A2(new_n804), .A3(new_n813), .A4(new_n918), .ZN(new_n943));
  NOR2_X1   g757(.A1(new_n942), .A2(new_n943), .ZN(new_n944));
  NAND3_X1  g758(.A1(new_n739), .A2(new_n931), .A3(new_n929), .ZN(new_n945));
  INV_X1    g759(.A(KEYINPUT52), .ZN(new_n946));
  NAND2_X1  g760(.A1(new_n945), .A2(new_n946), .ZN(new_n947));
  AND2_X1   g761(.A1(new_n921), .A2(KEYINPUT117), .ZN(new_n948));
  NOR2_X1   g762(.A1(new_n921), .A2(KEYINPUT117), .ZN(new_n949));
  NOR2_X1   g763(.A1(new_n948), .A2(new_n949), .ZN(new_n950));
  NAND3_X1  g764(.A1(new_n739), .A2(KEYINPUT52), .A3(new_n929), .ZN(new_n951));
  OAI21_X1  g765(.A(new_n947), .B1(new_n950), .B2(new_n951), .ZN(new_n952));
  INV_X1    g766(.A(KEYINPUT53), .ZN(new_n953));
  NAND3_X1  g767(.A1(new_n944), .A2(new_n952), .A3(new_n953), .ZN(new_n954));
  NAND3_X1  g768(.A1(new_n934), .A2(KEYINPUT54), .A3(new_n954), .ZN(new_n955));
  OAI21_X1  g769(.A(new_n953), .B1(new_n920), .B2(new_n933), .ZN(new_n956));
  NAND4_X1  g770(.A1(new_n918), .A2(new_n813), .A3(KEYINPUT53), .A4(new_n801), .ZN(new_n957));
  NOR2_X1   g771(.A1(new_n942), .A2(new_n957), .ZN(new_n958));
  AOI21_X1  g772(.A(KEYINPUT54), .B1(new_n958), .B2(new_n952), .ZN(new_n959));
  NAND2_X1  g773(.A1(new_n956), .A2(new_n959), .ZN(new_n960));
  AND3_X1   g774(.A1(new_n888), .A2(new_n955), .A3(new_n960), .ZN(new_n961));
  NOR2_X1   g775(.A1(G952), .A2(G953), .ZN(new_n962));
  NOR4_X1   g776(.A1(new_n592), .A2(new_n650), .A3(new_n642), .A4(new_n661), .ZN(new_n963));
  INV_X1    g777(.A(KEYINPUT49), .ZN(new_n964));
  OAI21_X1  g778(.A(new_n963), .B1(new_n870), .B2(new_n964), .ZN(new_n965));
  AOI21_X1  g779(.A(new_n965), .B1(new_n964), .B2(new_n870), .ZN(new_n966));
  NAND2_X1  g780(.A1(new_n966), .A2(new_n855), .ZN(new_n967));
  OAI22_X1  g781(.A1(new_n961), .A2(new_n962), .B1(new_n708), .B2(new_n967), .ZN(G75));
  NAND2_X1  g782(.A1(new_n958), .A2(new_n952), .ZN(new_n969));
  AOI21_X1  g783(.A(new_n251), .B1(new_n956), .B2(new_n969), .ZN(new_n970));
  NAND2_X1  g784(.A1(new_n970), .A2(new_n489), .ZN(new_n971));
  INV_X1    g785(.A(KEYINPUT56), .ZN(new_n972));
  NOR3_X1   g786(.A1(new_n493), .A2(new_n494), .A3(new_n492), .ZN(new_n973));
  NOR2_X1   g787(.A1(new_n973), .A2(new_n452), .ZN(new_n974));
  XNOR2_X1  g788(.A(new_n974), .B(KEYINPUT55), .ZN(new_n975));
  AND3_X1   g789(.A1(new_n971), .A2(new_n972), .A3(new_n975), .ZN(new_n976));
  AOI21_X1  g790(.A(new_n975), .B1(new_n971), .B2(new_n972), .ZN(new_n977));
  NOR2_X1   g791(.A1(new_n237), .A2(G952), .ZN(new_n978));
  NOR3_X1   g792(.A1(new_n976), .A2(new_n977), .A3(new_n978), .ZN(G51));
  NAND3_X1  g793(.A1(new_n922), .A2(KEYINPUT52), .A3(new_n929), .ZN(new_n980));
  NAND2_X1  g794(.A1(new_n947), .A2(new_n980), .ZN(new_n981));
  AOI21_X1  g795(.A(KEYINPUT53), .B1(new_n944), .B2(new_n981), .ZN(new_n982));
  INV_X1    g796(.A(KEYINPUT54), .ZN(new_n983));
  AND2_X1   g797(.A1(new_n801), .A2(KEYINPUT53), .ZN(new_n984));
  NAND4_X1  g798(.A1(new_n898), .A2(new_n919), .A3(new_n907), .A4(new_n984), .ZN(new_n985));
  AND3_X1   g799(.A1(new_n739), .A2(KEYINPUT52), .A3(new_n929), .ZN(new_n986));
  XNOR2_X1  g800(.A(new_n921), .B(KEYINPUT117), .ZN(new_n987));
  AOI22_X1  g801(.A1(new_n986), .A2(new_n987), .B1(new_n945), .B2(new_n946), .ZN(new_n988));
  OAI21_X1  g802(.A(new_n983), .B1(new_n985), .B2(new_n988), .ZN(new_n989));
  OAI21_X1  g803(.A(KEYINPUT125), .B1(new_n982), .B2(new_n989), .ZN(new_n990));
  NOR2_X1   g804(.A1(new_n985), .A2(new_n988), .ZN(new_n991));
  OAI21_X1  g805(.A(KEYINPUT54), .B1(new_n982), .B2(new_n991), .ZN(new_n992));
  INV_X1    g806(.A(KEYINPUT125), .ZN(new_n993));
  NAND3_X1  g807(.A1(new_n956), .A2(new_n959), .A3(new_n993), .ZN(new_n994));
  NAND3_X1  g808(.A1(new_n990), .A2(new_n992), .A3(new_n994), .ZN(new_n995));
  XNOR2_X1  g809(.A(new_n538), .B(KEYINPUT57), .ZN(new_n996));
  NAND2_X1  g810(.A1(new_n995), .A2(new_n996), .ZN(new_n997));
  NAND2_X1  g811(.A1(new_n997), .A2(new_n535), .ZN(new_n998));
  NAND3_X1  g812(.A1(new_n970), .A2(new_n815), .A3(new_n817), .ZN(new_n999));
  AOI21_X1  g813(.A(new_n978), .B1(new_n998), .B2(new_n999), .ZN(G54));
  NAND2_X1  g814(.A1(KEYINPUT58), .A2(G475), .ZN(new_n1001));
  XOR2_X1   g815(.A(new_n1001), .B(KEYINPUT126), .Z(new_n1002));
  AND3_X1   g816(.A1(new_n970), .A2(new_n695), .A3(new_n1002), .ZN(new_n1003));
  AOI21_X1  g817(.A(new_n695), .B1(new_n970), .B2(new_n1002), .ZN(new_n1004));
  NOR3_X1   g818(.A1(new_n1003), .A2(new_n1004), .A3(new_n978), .ZN(G60));
  INV_X1    g819(.A(new_n978), .ZN(new_n1006));
  NAND2_X1  g820(.A1(G478), .A2(G902), .ZN(new_n1007));
  XOR2_X1   g821(.A(new_n1007), .B(KEYINPUT59), .Z(new_n1008));
  AOI21_X1  g822(.A(new_n1008), .B1(new_n955), .B2(new_n960), .ZN(new_n1009));
  OAI21_X1  g823(.A(new_n1006), .B1(new_n1009), .B2(new_n646), .ZN(new_n1010));
  INV_X1    g824(.A(new_n1008), .ZN(new_n1011));
  AND2_X1   g825(.A1(new_n646), .A2(new_n1011), .ZN(new_n1012));
  AOI21_X1  g826(.A(new_n1010), .B1(new_n995), .B2(new_n1012), .ZN(G63));
  NAND2_X1  g827(.A1(G217), .A2(G902), .ZN(new_n1014));
  XNOR2_X1  g828(.A(new_n1014), .B(KEYINPUT60), .ZN(new_n1015));
  AOI21_X1  g829(.A(new_n1015), .B1(new_n956), .B2(new_n969), .ZN(new_n1016));
  NAND2_X1  g830(.A1(new_n1016), .A2(new_n683), .ZN(new_n1017));
  OAI211_X1 g831(.A(new_n1017), .B(new_n1006), .C1(new_n250), .C2(new_n1016), .ZN(new_n1018));
  INV_X1    g832(.A(KEYINPUT61), .ZN(new_n1019));
  NAND2_X1  g833(.A1(new_n1018), .A2(new_n1019), .ZN(new_n1020));
  OR2_X1    g834(.A1(new_n1016), .A2(new_n250), .ZN(new_n1021));
  NAND4_X1  g835(.A1(new_n1021), .A2(KEYINPUT61), .A3(new_n1006), .A4(new_n1017), .ZN(new_n1022));
  NAND2_X1  g836(.A1(new_n1020), .A2(new_n1022), .ZN(G66));
  NAND2_X1  g837(.A1(G224), .A2(G953), .ZN(new_n1024));
  OAI22_X1  g838(.A1(new_n942), .A2(G953), .B1(new_n599), .B2(new_n1024), .ZN(new_n1025));
  OAI211_X1 g839(.A(new_n446), .B(new_n451), .C1(G898), .C2(new_n237), .ZN(new_n1026));
  XOR2_X1   g840(.A(new_n1025), .B(new_n1026), .Z(G69));
  NAND4_X1  g841(.A1(new_n825), .A2(new_n264), .A3(new_n767), .A4(new_n797), .ZN(new_n1028));
  AND4_X1   g842(.A1(new_n813), .A2(new_n834), .A3(new_n843), .A4(new_n1028), .ZN(new_n1029));
  AND2_X1   g843(.A1(new_n987), .A2(new_n739), .ZN(new_n1030));
  NAND4_X1  g844(.A1(new_n1029), .A2(new_n237), .A3(new_n805), .A4(new_n1030), .ZN(new_n1031));
  NAND2_X1  g845(.A1(G900), .A2(G953), .ZN(new_n1032));
  NAND2_X1  g846(.A1(new_n1031), .A2(new_n1032), .ZN(new_n1033));
  NAND2_X1  g847(.A1(G227), .A2(G900), .ZN(new_n1034));
  NAND2_X1  g848(.A1(new_n316), .A2(new_n326), .ZN(new_n1035));
  XNOR2_X1  g849(.A(new_n572), .B(KEYINPUT127), .ZN(new_n1036));
  XNOR2_X1  g850(.A(new_n1035), .B(new_n1036), .ZN(new_n1037));
  AND4_X1   g851(.A1(G953), .A2(new_n1033), .A3(new_n1034), .A4(new_n1037), .ZN(new_n1038));
  INV_X1    g852(.A(new_n1037), .ZN(new_n1039));
  AOI21_X1  g853(.A(new_n1039), .B1(new_n1031), .B2(new_n1032), .ZN(new_n1040));
  NAND2_X1  g854(.A1(new_n1039), .A2(new_n237), .ZN(new_n1041));
  OR2_X1    g855(.A1(new_n651), .A2(new_n899), .ZN(new_n1042));
  NAND4_X1  g856(.A1(new_n389), .A2(new_n711), .A3(new_n826), .A4(new_n1042), .ZN(new_n1043));
  NAND3_X1  g857(.A1(new_n834), .A2(new_n843), .A3(new_n1043), .ZN(new_n1044));
  NAND2_X1  g858(.A1(new_n1030), .A2(new_n724), .ZN(new_n1045));
  AOI21_X1  g859(.A(new_n1044), .B1(new_n1045), .B2(KEYINPUT62), .ZN(new_n1046));
  OR2_X1    g860(.A1(new_n1045), .A2(KEYINPUT62), .ZN(new_n1047));
  AOI21_X1  g861(.A(new_n1041), .B1(new_n1046), .B2(new_n1047), .ZN(new_n1048));
  AOI21_X1  g862(.A(new_n237), .B1(G227), .B2(G900), .ZN(new_n1049));
  NOR3_X1   g863(.A1(new_n1040), .A2(new_n1048), .A3(new_n1049), .ZN(new_n1050));
  NOR2_X1   g864(.A1(new_n1038), .A2(new_n1050), .ZN(G72));
  NAND2_X1  g865(.A1(G472), .A2(G902), .ZN(new_n1052));
  XOR2_X1   g866(.A(new_n1052), .B(KEYINPUT63), .Z(new_n1053));
  NAND2_X1  g867(.A1(new_n1046), .A2(new_n1047), .ZN(new_n1054));
  OAI21_X1  g868(.A(new_n1053), .B1(new_n1054), .B2(new_n942), .ZN(new_n1055));
  INV_X1    g869(.A(new_n717), .ZN(new_n1056));
  NAND2_X1  g870(.A1(new_n1055), .A2(new_n1056), .ZN(new_n1057));
  NAND3_X1  g871(.A1(new_n1029), .A2(new_n805), .A3(new_n1030), .ZN(new_n1058));
  OAI21_X1  g872(.A(new_n1053), .B1(new_n1058), .B2(new_n942), .ZN(new_n1059));
  NOR2_X1   g873(.A1(new_n716), .A2(new_n341), .ZN(new_n1060));
  AOI21_X1  g874(.A(new_n978), .B1(new_n1059), .B2(new_n1060), .ZN(new_n1061));
  OAI21_X1  g875(.A(new_n1053), .B1(new_n716), .B2(new_n341), .ZN(new_n1062));
  NOR2_X1   g876(.A1(new_n1056), .A2(new_n1062), .ZN(new_n1063));
  NAND3_X1  g877(.A1(new_n934), .A2(new_n954), .A3(new_n1063), .ZN(new_n1064));
  AND3_X1   g878(.A1(new_n1057), .A2(new_n1061), .A3(new_n1064), .ZN(G57));
endmodule


