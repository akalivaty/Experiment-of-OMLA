

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
         n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598,
         n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609,
         n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620,
         n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631,
         n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642,
         n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653,
         n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664,
         n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675,
         n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686,
         n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697,
         n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708,
         n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719,
         n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, n730,
         n731, n732, n733, n734, n735, n736, n737, n738, n739, n740, n741,
         n742, n743, n744, n745, n746, n747, n748, n749, n750, n751, n752,
         n753, n754, n755, n756, n757, n758, n759, n760, n761, n762, n763,
         n764, n765, n766, n767, n768, n769, n770, n771, n772, n773, n774,
         n775, n776, n777, n778, n779, n780, n781, n782, n783, n784, n785,
         n786, n787, n788, n789, n790, n791, n792, n793, n794, n795, n796,
         n797, n798, n799, n800, n801, n802, n803, n804, n805, n806, n807,
         n808, n809, n810, n811, n812, n813, n814, n815, n816, n817, n818,
         n819, n820, n821, n822, n823, n824, n825, n826, n827, n828, n829,
         n830, n831, n832, n833, n834, n835, n836, n837, n838, n839, n840,
         n841, n842, n843, n844, n845, n846, n847, n848, n849, n850, n851,
         n852, n853, n854, n855, n856, n857, n858, n859, n860, n861, n862,
         n863, n864, n865, n866, n867, n868, n869, n870, n871, n872, n873,
         n874, n875, n876, n877, n878, n879, n880, n881, n882, n883, n884,
         n885, n886, n887, n888, n889, n890, n891, n892, n893, n894, n895,
         n896, n897, n898, n899, n900, n901, n902, n903, n904, n905, n906,
         n907, n908, n909, n910, n911, n912, n913, n914, n915, n916, n917,
         n918, n919, n920, n921, n922, n923, n924, n925, n926, n927, n928,
         n929, n930, n931, n932, n933, n934, n935, n936, n937, n938, n939,
         n940, n941, n942, n943, n944, n945, n946, n947, n948, n949, n950,
         n951, n952, n953, n954, n955, n956, n957, n958, n959, n960, n961,
         n962, n963, n964, n965, n966, n967, n968, n969, n970, n971, n972,
         n973, n974, n975, n976, n977, n978, n979, n980, n981, n982, n983,
         n984, n985, n986, n987, n988, n989, n990, n991, n992, n993, n994,
         n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
         n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
         n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
         n1025, n1026, n1027;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NOR2_X1 U552 ( .A1(n683), .A2(n938), .ZN(n685) );
  NAND2_X1 U553 ( .A1(n682), .A2(n518), .ZN(n683) );
  OR2_X1 U554 ( .A1(n690), .A2(n691), .ZN(n689) );
  NAND2_X1 U555 ( .A1(n724), .A2(G1341), .ZN(n518) );
  NAND2_X1 U556 ( .A1(n801), .A2(n800), .ZN(n519) );
  OR2_X1 U557 ( .A1(n787), .A2(n786), .ZN(n520) );
  XOR2_X1 U558 ( .A(KEYINPUT97), .B(n722), .Z(n521) );
  INV_X1 U559 ( .A(KEYINPUT26), .ZN(n680) );
  INV_X1 U560 ( .A(KEYINPUT64), .ZN(n684) );
  NAND2_X1 U561 ( .A1(n679), .A2(n756), .ZN(n724) );
  NOR2_X1 U562 ( .A1(G2105), .A2(G2104), .ZN(n522) );
  NOR2_X1 U563 ( .A1(n539), .A2(n538), .ZN(G160) );
  XOR2_X2 U564 ( .A(KEYINPUT17), .B(n522), .Z(n879) );
  NAND2_X1 U565 ( .A1(n879), .A2(G138), .ZN(n524) );
  AND2_X1 U566 ( .A1(G2105), .A2(G2104), .ZN(n887) );
  NAND2_X1 U567 ( .A1(n887), .A2(G114), .ZN(n523) );
  NAND2_X1 U568 ( .A1(n524), .A2(n523), .ZN(n532) );
  INV_X1 U569 ( .A(G2104), .ZN(n525) );
  AND2_X1 U570 ( .A1(n525), .A2(G2105), .ZN(n885) );
  NAND2_X1 U571 ( .A1(G126), .A2(n885), .ZN(n526) );
  XNOR2_X1 U572 ( .A(n526), .B(KEYINPUT86), .ZN(n530) );
  INV_X1 U573 ( .A(G2104), .ZN(n527) );
  NOR2_X4 U574 ( .A1(G2105), .A2(n527), .ZN(n881) );
  NAND2_X1 U575 ( .A1(G102), .A2(n881), .ZN(n528) );
  XOR2_X1 U576 ( .A(n528), .B(KEYINPUT87), .Z(n529) );
  NAND2_X1 U577 ( .A1(n530), .A2(n529), .ZN(n531) );
  NOR2_X1 U578 ( .A1(n532), .A2(n531), .ZN(G164) );
  NAND2_X1 U579 ( .A1(G101), .A2(n881), .ZN(n533) );
  XOR2_X1 U580 ( .A(KEYINPUT23), .B(n533), .Z(n535) );
  NAND2_X1 U581 ( .A1(n887), .A2(G113), .ZN(n534) );
  NAND2_X1 U582 ( .A1(n535), .A2(n534), .ZN(n539) );
  NAND2_X1 U583 ( .A1(G125), .A2(n885), .ZN(n537) );
  NAND2_X1 U584 ( .A1(G137), .A2(n879), .ZN(n536) );
  NAND2_X1 U585 ( .A1(n537), .A2(n536), .ZN(n538) );
  INV_X1 U586 ( .A(G651), .ZN(n544) );
  NOR2_X1 U587 ( .A1(G543), .A2(n544), .ZN(n540) );
  XOR2_X1 U588 ( .A(KEYINPUT1), .B(n540), .Z(n643) );
  NAND2_X1 U589 ( .A1(G64), .A2(n643), .ZN(n543) );
  XOR2_X1 U590 ( .A(KEYINPUT0), .B(G543), .Z(n621) );
  NOR2_X1 U591 ( .A1(G651), .A2(n621), .ZN(n541) );
  XOR2_X1 U592 ( .A(KEYINPUT65), .B(n541), .Z(n644) );
  NAND2_X1 U593 ( .A1(G52), .A2(n644), .ZN(n542) );
  NAND2_X1 U594 ( .A1(n543), .A2(n542), .ZN(n549) );
  NOR2_X1 U595 ( .A1(G651), .A2(G543), .ZN(n647) );
  NAND2_X1 U596 ( .A1(G90), .A2(n647), .ZN(n546) );
  NOR2_X1 U597 ( .A1(n621), .A2(n544), .ZN(n641) );
  NAND2_X1 U598 ( .A1(G77), .A2(n641), .ZN(n545) );
  NAND2_X1 U599 ( .A1(n546), .A2(n545), .ZN(n547) );
  XOR2_X1 U600 ( .A(KEYINPUT9), .B(n547), .Z(n548) );
  NOR2_X1 U601 ( .A1(n549), .A2(n548), .ZN(G171) );
  AND2_X1 U602 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U603 ( .A(G132), .ZN(G219) );
  INV_X1 U604 ( .A(G108), .ZN(G238) );
  NAND2_X1 U605 ( .A1(G7), .A2(G661), .ZN(n550) );
  XNOR2_X1 U606 ( .A(n550), .B(KEYINPUT68), .ZN(n551) );
  XNOR2_X1 U607 ( .A(KEYINPUT10), .B(n551), .ZN(G223) );
  INV_X1 U608 ( .A(G223), .ZN(n827) );
  NAND2_X1 U609 ( .A1(n827), .A2(G567), .ZN(n552) );
  XOR2_X1 U610 ( .A(KEYINPUT11), .B(n552), .Z(G234) );
  NAND2_X1 U611 ( .A1(n647), .A2(G81), .ZN(n553) );
  XNOR2_X1 U612 ( .A(n553), .B(KEYINPUT12), .ZN(n555) );
  NAND2_X1 U613 ( .A1(G68), .A2(n641), .ZN(n554) );
  NAND2_X1 U614 ( .A1(n555), .A2(n554), .ZN(n556) );
  XOR2_X1 U615 ( .A(KEYINPUT13), .B(n556), .Z(n560) );
  NAND2_X1 U616 ( .A1(G56), .A2(n643), .ZN(n557) );
  XNOR2_X1 U617 ( .A(n557), .B(KEYINPUT69), .ZN(n558) );
  XNOR2_X1 U618 ( .A(n558), .B(KEYINPUT14), .ZN(n559) );
  NOR2_X1 U619 ( .A1(n560), .A2(n559), .ZN(n562) );
  NAND2_X1 U620 ( .A1(n644), .A2(G43), .ZN(n561) );
  NAND2_X1 U621 ( .A1(n562), .A2(n561), .ZN(n938) );
  INV_X1 U622 ( .A(G860), .ZN(n593) );
  OR2_X1 U623 ( .A1(n938), .A2(n593), .ZN(G153) );
  INV_X1 U624 ( .A(G171), .ZN(G301) );
  NAND2_X1 U625 ( .A1(G66), .A2(n643), .ZN(n564) );
  NAND2_X1 U626 ( .A1(G54), .A2(n644), .ZN(n563) );
  NAND2_X1 U627 ( .A1(n564), .A2(n563), .ZN(n568) );
  NAND2_X1 U628 ( .A1(G92), .A2(n647), .ZN(n566) );
  NAND2_X1 U629 ( .A1(G79), .A2(n641), .ZN(n565) );
  NAND2_X1 U630 ( .A1(n566), .A2(n565), .ZN(n567) );
  NOR2_X1 U631 ( .A1(n568), .A2(n567), .ZN(n569) );
  XNOR2_X1 U632 ( .A(n569), .B(KEYINPUT15), .ZN(n690) );
  INV_X1 U633 ( .A(G868), .ZN(n662) );
  NAND2_X1 U634 ( .A1(n690), .A2(n662), .ZN(n570) );
  XNOR2_X1 U635 ( .A(n570), .B(KEYINPUT70), .ZN(n572) );
  NAND2_X1 U636 ( .A1(G868), .A2(G301), .ZN(n571) );
  NAND2_X1 U637 ( .A1(n572), .A2(n571), .ZN(G284) );
  NAND2_X1 U638 ( .A1(G63), .A2(n643), .ZN(n574) );
  NAND2_X1 U639 ( .A1(G51), .A2(n644), .ZN(n573) );
  NAND2_X1 U640 ( .A1(n574), .A2(n573), .ZN(n575) );
  XNOR2_X1 U641 ( .A(KEYINPUT6), .B(n575), .ZN(n581) );
  NAND2_X1 U642 ( .A1(n647), .A2(G89), .ZN(n576) );
  XNOR2_X1 U643 ( .A(n576), .B(KEYINPUT4), .ZN(n578) );
  NAND2_X1 U644 ( .A1(G76), .A2(n641), .ZN(n577) );
  NAND2_X1 U645 ( .A1(n578), .A2(n577), .ZN(n579) );
  XOR2_X1 U646 ( .A(n579), .B(KEYINPUT5), .Z(n580) );
  NOR2_X1 U647 ( .A1(n581), .A2(n580), .ZN(n582) );
  XOR2_X1 U648 ( .A(KEYINPUT71), .B(n582), .Z(n583) );
  XOR2_X1 U649 ( .A(KEYINPUT7), .B(n583), .Z(G168) );
  XOR2_X1 U650 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U651 ( .A1(G65), .A2(n643), .ZN(n585) );
  NAND2_X1 U652 ( .A1(G53), .A2(n644), .ZN(n584) );
  NAND2_X1 U653 ( .A1(n585), .A2(n584), .ZN(n586) );
  XOR2_X1 U654 ( .A(KEYINPUT66), .B(n586), .Z(n590) );
  NAND2_X1 U655 ( .A1(G91), .A2(n647), .ZN(n588) );
  NAND2_X1 U656 ( .A1(G78), .A2(n641), .ZN(n587) );
  AND2_X1 U657 ( .A1(n588), .A2(n587), .ZN(n589) );
  NAND2_X1 U658 ( .A1(n590), .A2(n589), .ZN(G299) );
  NOR2_X1 U659 ( .A1(G286), .A2(n662), .ZN(n592) );
  NOR2_X1 U660 ( .A1(G868), .A2(G299), .ZN(n591) );
  NOR2_X1 U661 ( .A1(n592), .A2(n591), .ZN(G297) );
  NAND2_X1 U662 ( .A1(n593), .A2(G559), .ZN(n594) );
  INV_X1 U663 ( .A(n690), .ZN(n937) );
  NAND2_X1 U664 ( .A1(n594), .A2(n937), .ZN(n595) );
  XNOR2_X1 U665 ( .A(n595), .B(KEYINPUT16), .ZN(G148) );
  NAND2_X1 U666 ( .A1(n937), .A2(G868), .ZN(n596) );
  NOR2_X1 U667 ( .A1(G559), .A2(n596), .ZN(n597) );
  XNOR2_X1 U668 ( .A(n597), .B(KEYINPUT72), .ZN(n599) );
  NOR2_X1 U669 ( .A1(n938), .A2(G868), .ZN(n598) );
  NOR2_X1 U670 ( .A1(n599), .A2(n598), .ZN(G282) );
  NAND2_X1 U671 ( .A1(G99), .A2(n881), .ZN(n601) );
  NAND2_X1 U672 ( .A1(G111), .A2(n887), .ZN(n600) );
  NAND2_X1 U673 ( .A1(n601), .A2(n600), .ZN(n602) );
  XNOR2_X1 U674 ( .A(n602), .B(KEYINPUT73), .ZN(n604) );
  NAND2_X1 U675 ( .A1(G135), .A2(n879), .ZN(n603) );
  NAND2_X1 U676 ( .A1(n604), .A2(n603), .ZN(n607) );
  NAND2_X1 U677 ( .A1(n885), .A2(G123), .ZN(n605) );
  XOR2_X1 U678 ( .A(KEYINPUT18), .B(n605), .Z(n606) );
  NOR2_X1 U679 ( .A1(n607), .A2(n606), .ZN(n1002) );
  XNOR2_X1 U680 ( .A(n1002), .B(G2096), .ZN(n609) );
  INV_X1 U681 ( .A(G2100), .ZN(n608) );
  NAND2_X1 U682 ( .A1(n609), .A2(n608), .ZN(G156) );
  NAND2_X1 U683 ( .A1(G75), .A2(n641), .ZN(n610) );
  XNOR2_X1 U684 ( .A(n610), .B(KEYINPUT82), .ZN(n617) );
  NAND2_X1 U685 ( .A1(G62), .A2(n643), .ZN(n612) );
  NAND2_X1 U686 ( .A1(G50), .A2(n644), .ZN(n611) );
  NAND2_X1 U687 ( .A1(n612), .A2(n611), .ZN(n615) );
  NAND2_X1 U688 ( .A1(G88), .A2(n647), .ZN(n613) );
  XNOR2_X1 U689 ( .A(KEYINPUT81), .B(n613), .ZN(n614) );
  NOR2_X1 U690 ( .A1(n615), .A2(n614), .ZN(n616) );
  NAND2_X1 U691 ( .A1(n617), .A2(n616), .ZN(G303) );
  INV_X1 U692 ( .A(G303), .ZN(G166) );
  NAND2_X1 U693 ( .A1(G49), .A2(n644), .ZN(n619) );
  NAND2_X1 U694 ( .A1(G74), .A2(G651), .ZN(n618) );
  NAND2_X1 U695 ( .A1(n619), .A2(n618), .ZN(n620) );
  NOR2_X1 U696 ( .A1(n643), .A2(n620), .ZN(n623) );
  NAND2_X1 U697 ( .A1(n621), .A2(G87), .ZN(n622) );
  NAND2_X1 U698 ( .A1(n623), .A2(n622), .ZN(G288) );
  NAND2_X1 U699 ( .A1(G86), .A2(n647), .ZN(n625) );
  NAND2_X1 U700 ( .A1(G48), .A2(n644), .ZN(n624) );
  NAND2_X1 U701 ( .A1(n625), .A2(n624), .ZN(n628) );
  NAND2_X1 U702 ( .A1(n643), .A2(G61), .ZN(n626) );
  XOR2_X1 U703 ( .A(KEYINPUT78), .B(n626), .Z(n627) );
  NOR2_X1 U704 ( .A1(n628), .A2(n627), .ZN(n632) );
  XOR2_X1 U705 ( .A(KEYINPUT79), .B(KEYINPUT2), .Z(n630) );
  NAND2_X1 U706 ( .A1(G73), .A2(n641), .ZN(n629) );
  XNOR2_X1 U707 ( .A(n630), .B(n629), .ZN(n631) );
  NAND2_X1 U708 ( .A1(n632), .A2(n631), .ZN(n633) );
  XNOR2_X1 U709 ( .A(n633), .B(KEYINPUT80), .ZN(G305) );
  AND2_X1 U710 ( .A1(n643), .A2(G60), .ZN(n637) );
  NAND2_X1 U711 ( .A1(G85), .A2(n647), .ZN(n635) );
  NAND2_X1 U712 ( .A1(G72), .A2(n641), .ZN(n634) );
  NAND2_X1 U713 ( .A1(n635), .A2(n634), .ZN(n636) );
  NOR2_X1 U714 ( .A1(n637), .A2(n636), .ZN(n639) );
  NAND2_X1 U715 ( .A1(n644), .A2(G47), .ZN(n638) );
  NAND2_X1 U716 ( .A1(n639), .A2(n638), .ZN(G290) );
  NAND2_X1 U717 ( .A1(G559), .A2(n937), .ZN(n640) );
  XNOR2_X1 U718 ( .A(n640), .B(KEYINPUT74), .ZN(n833) );
  NAND2_X1 U719 ( .A1(G80), .A2(n641), .ZN(n642) );
  XNOR2_X1 U720 ( .A(n642), .B(KEYINPUT76), .ZN(n652) );
  NAND2_X1 U721 ( .A1(G67), .A2(n643), .ZN(n646) );
  NAND2_X1 U722 ( .A1(G55), .A2(n644), .ZN(n645) );
  NAND2_X1 U723 ( .A1(n646), .A2(n645), .ZN(n650) );
  NAND2_X1 U724 ( .A1(G93), .A2(n647), .ZN(n648) );
  XNOR2_X1 U725 ( .A(KEYINPUT75), .B(n648), .ZN(n649) );
  NOR2_X1 U726 ( .A1(n650), .A2(n649), .ZN(n651) );
  NAND2_X1 U727 ( .A1(n652), .A2(n651), .ZN(n653) );
  XOR2_X1 U728 ( .A(KEYINPUT77), .B(n653), .Z(n835) );
  XOR2_X1 U729 ( .A(KEYINPUT83), .B(KEYINPUT19), .Z(n654) );
  XNOR2_X1 U730 ( .A(G288), .B(n654), .ZN(n655) );
  XOR2_X1 U731 ( .A(n835), .B(n655), .Z(n657) );
  XNOR2_X1 U732 ( .A(n938), .B(G305), .ZN(n656) );
  XNOR2_X1 U733 ( .A(n657), .B(n656), .ZN(n658) );
  XNOR2_X1 U734 ( .A(G166), .B(n658), .ZN(n660) );
  INV_X1 U735 ( .A(G299), .ZN(n700) );
  XNOR2_X1 U736 ( .A(G290), .B(n700), .ZN(n659) );
  XNOR2_X1 U737 ( .A(n660), .B(n659), .ZN(n903) );
  XNOR2_X1 U738 ( .A(n833), .B(n903), .ZN(n661) );
  NAND2_X1 U739 ( .A1(n661), .A2(G868), .ZN(n664) );
  NAND2_X1 U740 ( .A1(n662), .A2(n835), .ZN(n663) );
  NAND2_X1 U741 ( .A1(n664), .A2(n663), .ZN(G295) );
  NAND2_X1 U742 ( .A1(G2078), .A2(G2084), .ZN(n665) );
  XOR2_X1 U743 ( .A(KEYINPUT20), .B(n665), .Z(n666) );
  NAND2_X1 U744 ( .A1(G2090), .A2(n666), .ZN(n667) );
  XNOR2_X1 U745 ( .A(KEYINPUT21), .B(n667), .ZN(n668) );
  NAND2_X1 U746 ( .A1(n668), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U747 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  XNOR2_X1 U748 ( .A(KEYINPUT67), .B(G82), .ZN(G220) );
  NAND2_X1 U749 ( .A1(G120), .A2(G69), .ZN(n669) );
  XNOR2_X1 U750 ( .A(KEYINPUT84), .B(n669), .ZN(n670) );
  NOR2_X1 U751 ( .A1(G238), .A2(n670), .ZN(n671) );
  NAND2_X1 U752 ( .A1(G57), .A2(n671), .ZN(n831) );
  NAND2_X1 U753 ( .A1(n831), .A2(G567), .ZN(n676) );
  NOR2_X1 U754 ( .A1(G219), .A2(G220), .ZN(n672) );
  XOR2_X1 U755 ( .A(KEYINPUT22), .B(n672), .Z(n673) );
  NOR2_X1 U756 ( .A1(G218), .A2(n673), .ZN(n674) );
  NAND2_X1 U757 ( .A1(G96), .A2(n674), .ZN(n832) );
  NAND2_X1 U758 ( .A1(n832), .A2(G2106), .ZN(n675) );
  NAND2_X1 U759 ( .A1(n676), .A2(n675), .ZN(n837) );
  NAND2_X1 U760 ( .A1(G661), .A2(G483), .ZN(n677) );
  XOR2_X1 U761 ( .A(KEYINPUT85), .B(n677), .Z(n678) );
  NOR2_X1 U762 ( .A1(n837), .A2(n678), .ZN(n830) );
  NAND2_X1 U763 ( .A1(n830), .A2(G36), .ZN(G176) );
  AND2_X1 U764 ( .A1(G160), .A2(G40), .ZN(n679) );
  NOR2_X2 U765 ( .A1(G164), .A2(G1384), .ZN(n756) );
  INV_X1 U766 ( .A(G1996), .ZN(n809) );
  NOR2_X1 U767 ( .A1(n724), .A2(n809), .ZN(n681) );
  XNOR2_X1 U768 ( .A(n681), .B(n680), .ZN(n682) );
  XNOR2_X1 U769 ( .A(n685), .B(n684), .ZN(n691) );
  NOR2_X1 U770 ( .A1(G2067), .A2(n724), .ZN(n687) );
  INV_X1 U771 ( .A(n724), .ZN(n705) );
  NOR2_X1 U772 ( .A1(n705), .A2(G1348), .ZN(n686) );
  NOR2_X1 U773 ( .A1(n687), .A2(n686), .ZN(n688) );
  NAND2_X1 U774 ( .A1(n689), .A2(n688), .ZN(n693) );
  NAND2_X1 U775 ( .A1(n691), .A2(n690), .ZN(n692) );
  NAND2_X1 U776 ( .A1(n693), .A2(n692), .ZN(n698) );
  NAND2_X1 U777 ( .A1(n705), .A2(G2072), .ZN(n694) );
  XNOR2_X1 U778 ( .A(n694), .B(KEYINPUT27), .ZN(n696) );
  INV_X1 U779 ( .A(G1956), .ZN(n953) );
  NOR2_X1 U780 ( .A1(n953), .A2(n705), .ZN(n695) );
  NOR2_X1 U781 ( .A1(n696), .A2(n695), .ZN(n699) );
  NAND2_X1 U782 ( .A1(n700), .A2(n699), .ZN(n697) );
  NAND2_X1 U783 ( .A1(n698), .A2(n697), .ZN(n703) );
  NOR2_X1 U784 ( .A1(n700), .A2(n699), .ZN(n701) );
  XOR2_X1 U785 ( .A(n701), .B(KEYINPUT28), .Z(n702) );
  NAND2_X1 U786 ( .A1(n703), .A2(n702), .ZN(n704) );
  XOR2_X1 U787 ( .A(KEYINPUT29), .B(n704), .Z(n711) );
  XOR2_X1 U788 ( .A(G2078), .B(KEYINPUT25), .Z(n975) );
  NOR2_X1 U789 ( .A1(n975), .A2(n724), .ZN(n707) );
  NOR2_X1 U790 ( .A1(n705), .A2(G1961), .ZN(n706) );
  NOR2_X1 U791 ( .A1(n707), .A2(n706), .ZN(n708) );
  XNOR2_X1 U792 ( .A(KEYINPUT95), .B(n708), .ZN(n716) );
  NAND2_X1 U793 ( .A1(G171), .A2(n716), .ZN(n709) );
  XNOR2_X1 U794 ( .A(n709), .B(KEYINPUT96), .ZN(n710) );
  NAND2_X1 U795 ( .A1(n711), .A2(n710), .ZN(n721) );
  NAND2_X1 U796 ( .A1(G8), .A2(n724), .ZN(n797) );
  NOR2_X1 U797 ( .A1(G1966), .A2(n797), .ZN(n735) );
  NOR2_X1 U798 ( .A1(G2084), .A2(n724), .ZN(n712) );
  XOR2_X1 U799 ( .A(KEYINPUT94), .B(n712), .Z(n731) );
  NAND2_X1 U800 ( .A1(G8), .A2(n731), .ZN(n713) );
  NOR2_X1 U801 ( .A1(n735), .A2(n713), .ZN(n714) );
  XOR2_X1 U802 ( .A(KEYINPUT30), .B(n714), .Z(n715) );
  NOR2_X1 U803 ( .A1(G168), .A2(n715), .ZN(n718) );
  NOR2_X1 U804 ( .A1(G171), .A2(n716), .ZN(n717) );
  NOR2_X1 U805 ( .A1(n718), .A2(n717), .ZN(n719) );
  XOR2_X1 U806 ( .A(KEYINPUT31), .B(n719), .Z(n720) );
  NAND2_X1 U807 ( .A1(n721), .A2(n720), .ZN(n733) );
  NAND2_X1 U808 ( .A1(G286), .A2(n733), .ZN(n722) );
  NOR2_X1 U809 ( .A1(G1971), .A2(n797), .ZN(n723) );
  XNOR2_X1 U810 ( .A(n723), .B(KEYINPUT98), .ZN(n726) );
  NOR2_X1 U811 ( .A1(n724), .A2(G2090), .ZN(n725) );
  NOR2_X1 U812 ( .A1(n726), .A2(n725), .ZN(n727) );
  NAND2_X1 U813 ( .A1(G303), .A2(n727), .ZN(n728) );
  NAND2_X1 U814 ( .A1(n521), .A2(n728), .ZN(n729) );
  NAND2_X1 U815 ( .A1(n729), .A2(G8), .ZN(n730) );
  XNOR2_X1 U816 ( .A(n730), .B(KEYINPUT32), .ZN(n790) );
  INV_X1 U817 ( .A(n731), .ZN(n732) );
  NAND2_X1 U818 ( .A1(n732), .A2(G8), .ZN(n737) );
  INV_X1 U819 ( .A(n733), .ZN(n734) );
  NOR2_X1 U820 ( .A1(n735), .A2(n734), .ZN(n736) );
  NAND2_X1 U821 ( .A1(n737), .A2(n736), .ZN(n789) );
  INV_X1 U822 ( .A(n797), .ZN(n739) );
  NAND2_X1 U823 ( .A1(G288), .A2(G1976), .ZN(n738) );
  XOR2_X1 U824 ( .A(KEYINPUT99), .B(n738), .Z(n925) );
  AND2_X1 U825 ( .A1(n739), .A2(n925), .ZN(n740) );
  NOR2_X1 U826 ( .A1(KEYINPUT33), .A2(n740), .ZN(n744) );
  NOR2_X1 U827 ( .A1(G1976), .A2(G288), .ZN(n748) );
  NAND2_X1 U828 ( .A1(KEYINPUT33), .A2(n748), .ZN(n741) );
  NOR2_X1 U829 ( .A1(n797), .A2(n741), .ZN(n742) );
  XNOR2_X1 U830 ( .A(n742), .B(KEYINPUT100), .ZN(n743) );
  NOR2_X1 U831 ( .A1(n744), .A2(n743), .ZN(n746) );
  AND2_X1 U832 ( .A1(n789), .A2(n746), .ZN(n745) );
  NAND2_X1 U833 ( .A1(n790), .A2(n745), .ZN(n753) );
  INV_X1 U834 ( .A(n746), .ZN(n751) );
  NOR2_X1 U835 ( .A1(G1971), .A2(G303), .ZN(n747) );
  NOR2_X1 U836 ( .A1(n748), .A2(n747), .ZN(n928) );
  INV_X1 U837 ( .A(KEYINPUT33), .ZN(n749) );
  AND2_X1 U838 ( .A1(n928), .A2(n749), .ZN(n750) );
  OR2_X1 U839 ( .A1(n751), .A2(n750), .ZN(n752) );
  NAND2_X1 U840 ( .A1(n753), .A2(n752), .ZN(n754) );
  XNOR2_X1 U841 ( .A(n754), .B(KEYINPUT101), .ZN(n787) );
  XOR2_X1 U842 ( .A(G1981), .B(G305), .Z(n934) );
  INV_X1 U843 ( .A(n934), .ZN(n785) );
  NAND2_X1 U844 ( .A1(G160), .A2(G40), .ZN(n755) );
  NOR2_X1 U845 ( .A1(n756), .A2(n755), .ZN(n822) );
  NAND2_X1 U846 ( .A1(n881), .A2(G105), .ZN(n757) );
  XNOR2_X1 U847 ( .A(n757), .B(KEYINPUT38), .ZN(n759) );
  NAND2_X1 U848 ( .A1(G117), .A2(n887), .ZN(n758) );
  NAND2_X1 U849 ( .A1(n759), .A2(n758), .ZN(n763) );
  NAND2_X1 U850 ( .A1(G129), .A2(n885), .ZN(n761) );
  NAND2_X1 U851 ( .A1(G141), .A2(n879), .ZN(n760) );
  NAND2_X1 U852 ( .A1(n761), .A2(n760), .ZN(n762) );
  NOR2_X1 U853 ( .A1(n763), .A2(n762), .ZN(n866) );
  OR2_X1 U854 ( .A1(n809), .A2(n866), .ZN(n772) );
  NAND2_X1 U855 ( .A1(G95), .A2(n881), .ZN(n765) );
  NAND2_X1 U856 ( .A1(G131), .A2(n879), .ZN(n764) );
  NAND2_X1 U857 ( .A1(n765), .A2(n764), .ZN(n768) );
  NAND2_X1 U858 ( .A1(n887), .A2(G107), .ZN(n766) );
  XOR2_X1 U859 ( .A(KEYINPUT92), .B(n766), .Z(n767) );
  NOR2_X1 U860 ( .A1(n768), .A2(n767), .ZN(n770) );
  NAND2_X1 U861 ( .A1(n885), .A2(G119), .ZN(n769) );
  NAND2_X1 U862 ( .A1(n770), .A2(n769), .ZN(n865) );
  NAND2_X1 U863 ( .A1(G1991), .A2(n865), .ZN(n771) );
  NAND2_X1 U864 ( .A1(n772), .A2(n771), .ZN(n1006) );
  NAND2_X1 U865 ( .A1(n822), .A2(n1006), .ZN(n813) );
  XNOR2_X1 U866 ( .A(G2067), .B(KEYINPUT37), .ZN(n807) );
  NAND2_X1 U867 ( .A1(n885), .A2(G128), .ZN(n773) );
  XNOR2_X1 U868 ( .A(KEYINPUT90), .B(n773), .ZN(n776) );
  NAND2_X1 U869 ( .A1(n887), .A2(G116), .ZN(n774) );
  XOR2_X1 U870 ( .A(KEYINPUT91), .B(n774), .Z(n775) );
  NAND2_X1 U871 ( .A1(n776), .A2(n775), .ZN(n777) );
  XNOR2_X1 U872 ( .A(n777), .B(KEYINPUT35), .ZN(n782) );
  NAND2_X1 U873 ( .A1(G104), .A2(n881), .ZN(n779) );
  NAND2_X1 U874 ( .A1(G140), .A2(n879), .ZN(n778) );
  NAND2_X1 U875 ( .A1(n779), .A2(n778), .ZN(n780) );
  XOR2_X1 U876 ( .A(KEYINPUT34), .B(n780), .Z(n781) );
  NAND2_X1 U877 ( .A1(n782), .A2(n781), .ZN(n783) );
  XOR2_X1 U878 ( .A(n783), .B(KEYINPUT36), .Z(n894) );
  NOR2_X1 U879 ( .A1(n807), .A2(n894), .ZN(n1018) );
  NAND2_X1 U880 ( .A1(n822), .A2(n1018), .ZN(n817) );
  NAND2_X1 U881 ( .A1(n813), .A2(n817), .ZN(n784) );
  XOR2_X1 U882 ( .A(KEYINPUT93), .B(n784), .Z(n788) );
  OR2_X1 U883 ( .A1(n785), .A2(n788), .ZN(n786) );
  INV_X1 U884 ( .A(n788), .ZN(n801) );
  NAND2_X1 U885 ( .A1(n790), .A2(n789), .ZN(n793) );
  NOR2_X1 U886 ( .A1(G2090), .A2(G303), .ZN(n791) );
  NAND2_X1 U887 ( .A1(G8), .A2(n791), .ZN(n792) );
  NAND2_X1 U888 ( .A1(n793), .A2(n792), .ZN(n794) );
  NAND2_X1 U889 ( .A1(n794), .A2(n797), .ZN(n799) );
  NOR2_X1 U890 ( .A1(G1981), .A2(G305), .ZN(n795) );
  XOR2_X1 U891 ( .A(n795), .B(KEYINPUT24), .Z(n796) );
  OR2_X1 U892 ( .A1(n797), .A2(n796), .ZN(n798) );
  NAND2_X1 U893 ( .A1(n799), .A2(n798), .ZN(n800) );
  NAND2_X1 U894 ( .A1(n520), .A2(n519), .ZN(n802) );
  XNOR2_X1 U895 ( .A(n802), .B(KEYINPUT102), .ZN(n806) );
  XNOR2_X1 U896 ( .A(KEYINPUT88), .B(G1986), .ZN(n803) );
  XNOR2_X1 U897 ( .A(n803), .B(G290), .ZN(n927) );
  NAND2_X1 U898 ( .A1(n927), .A2(n822), .ZN(n804) );
  XOR2_X1 U899 ( .A(KEYINPUT89), .B(n804), .Z(n805) );
  NAND2_X1 U900 ( .A1(n806), .A2(n805), .ZN(n825) );
  AND2_X1 U901 ( .A1(n807), .A2(n894), .ZN(n808) );
  XOR2_X1 U902 ( .A(KEYINPUT106), .B(n808), .Z(n1016) );
  NAND2_X1 U903 ( .A1(n866), .A2(n809), .ZN(n998) );
  NOR2_X1 U904 ( .A1(G1986), .A2(G290), .ZN(n810) );
  XNOR2_X1 U905 ( .A(KEYINPUT103), .B(n810), .ZN(n812) );
  NOR2_X1 U906 ( .A1(G1991), .A2(n865), .ZN(n811) );
  XOR2_X1 U907 ( .A(KEYINPUT104), .B(n811), .Z(n1008) );
  NAND2_X1 U908 ( .A1(n812), .A2(n1008), .ZN(n814) );
  NAND2_X1 U909 ( .A1(n814), .A2(n813), .ZN(n815) );
  NAND2_X1 U910 ( .A1(n998), .A2(n815), .ZN(n816) );
  XOR2_X1 U911 ( .A(KEYINPUT39), .B(n816), .Z(n818) );
  NAND2_X1 U912 ( .A1(n818), .A2(n817), .ZN(n819) );
  XOR2_X1 U913 ( .A(KEYINPUT105), .B(n819), .Z(n820) );
  NAND2_X1 U914 ( .A1(n1016), .A2(n820), .ZN(n821) );
  NAND2_X1 U915 ( .A1(n822), .A2(n821), .ZN(n823) );
  XOR2_X1 U916 ( .A(KEYINPUT107), .B(n823), .Z(n824) );
  NAND2_X1 U917 ( .A1(n825), .A2(n824), .ZN(n826) );
  XNOR2_X1 U918 ( .A(KEYINPUT40), .B(n826), .ZN(G329) );
  NAND2_X1 U919 ( .A1(G2106), .A2(n827), .ZN(G217) );
  AND2_X1 U920 ( .A1(G15), .A2(G2), .ZN(n828) );
  NAND2_X1 U921 ( .A1(G661), .A2(n828), .ZN(G259) );
  NAND2_X1 U922 ( .A1(G3), .A2(G1), .ZN(n829) );
  NAND2_X1 U923 ( .A1(n830), .A2(n829), .ZN(G188) );
  XOR2_X1 U924 ( .A(G69), .B(KEYINPUT110), .Z(G235) );
  INV_X1 U926 ( .A(G120), .ZN(G236) );
  INV_X1 U927 ( .A(G96), .ZN(G221) );
  NOR2_X1 U928 ( .A1(n832), .A2(n831), .ZN(G325) );
  INV_X1 U929 ( .A(G325), .ZN(G261) );
  XNOR2_X1 U930 ( .A(n833), .B(n938), .ZN(n834) );
  NOR2_X1 U931 ( .A1(n834), .A2(G860), .ZN(n836) );
  XOR2_X1 U932 ( .A(n836), .B(n835), .Z(G145) );
  INV_X1 U933 ( .A(n837), .ZN(G319) );
  XOR2_X1 U934 ( .A(G2100), .B(G2096), .Z(n839) );
  XNOR2_X1 U935 ( .A(KEYINPUT42), .B(G2678), .ZN(n838) );
  XNOR2_X1 U936 ( .A(n839), .B(n838), .ZN(n843) );
  XOR2_X1 U937 ( .A(KEYINPUT43), .B(G2090), .Z(n841) );
  XNOR2_X1 U938 ( .A(G2067), .B(G2072), .ZN(n840) );
  XNOR2_X1 U939 ( .A(n841), .B(n840), .ZN(n842) );
  XOR2_X1 U940 ( .A(n843), .B(n842), .Z(n845) );
  XNOR2_X1 U941 ( .A(G2078), .B(G2084), .ZN(n844) );
  XNOR2_X1 U942 ( .A(n845), .B(n844), .ZN(G227) );
  XOR2_X1 U943 ( .A(KEYINPUT112), .B(G1991), .Z(n847) );
  XNOR2_X1 U944 ( .A(G1996), .B(G1956), .ZN(n846) );
  XNOR2_X1 U945 ( .A(n847), .B(n846), .ZN(n848) );
  XOR2_X1 U946 ( .A(n848), .B(KEYINPUT41), .Z(n850) );
  XNOR2_X1 U947 ( .A(G1986), .B(G1971), .ZN(n849) );
  XNOR2_X1 U948 ( .A(n850), .B(n849), .ZN(n854) );
  XOR2_X1 U949 ( .A(G1976), .B(G1981), .Z(n852) );
  XNOR2_X1 U950 ( .A(G1966), .B(G1961), .ZN(n851) );
  XNOR2_X1 U951 ( .A(n852), .B(n851), .ZN(n853) );
  XOR2_X1 U952 ( .A(n854), .B(n853), .Z(n856) );
  XNOR2_X1 U953 ( .A(G2474), .B(KEYINPUT111), .ZN(n855) );
  XNOR2_X1 U954 ( .A(n856), .B(n855), .ZN(G229) );
  NAND2_X1 U955 ( .A1(G124), .A2(n885), .ZN(n857) );
  XOR2_X1 U956 ( .A(KEYINPUT113), .B(n857), .Z(n858) );
  XNOR2_X1 U957 ( .A(n858), .B(KEYINPUT44), .ZN(n860) );
  NAND2_X1 U958 ( .A1(G100), .A2(n881), .ZN(n859) );
  NAND2_X1 U959 ( .A1(n860), .A2(n859), .ZN(n864) );
  NAND2_X1 U960 ( .A1(G112), .A2(n887), .ZN(n862) );
  NAND2_X1 U961 ( .A1(G136), .A2(n879), .ZN(n861) );
  NAND2_X1 U962 ( .A1(n862), .A2(n861), .ZN(n863) );
  NOR2_X1 U963 ( .A1(n864), .A2(n863), .ZN(G162) );
  XNOR2_X1 U964 ( .A(n865), .B(G162), .ZN(n868) );
  XNOR2_X1 U965 ( .A(G160), .B(n866), .ZN(n867) );
  XNOR2_X1 U966 ( .A(n868), .B(n867), .ZN(n878) );
  NAND2_X1 U967 ( .A1(G130), .A2(n885), .ZN(n870) );
  NAND2_X1 U968 ( .A1(G118), .A2(n887), .ZN(n869) );
  NAND2_X1 U969 ( .A1(n870), .A2(n869), .ZN(n876) );
  NAND2_X1 U970 ( .A1(n881), .A2(G106), .ZN(n871) );
  XNOR2_X1 U971 ( .A(n871), .B(KEYINPUT114), .ZN(n873) );
  NAND2_X1 U972 ( .A1(G142), .A2(n879), .ZN(n872) );
  NAND2_X1 U973 ( .A1(n873), .A2(n872), .ZN(n874) );
  XOR2_X1 U974 ( .A(KEYINPUT45), .B(n874), .Z(n875) );
  NOR2_X1 U975 ( .A1(n876), .A2(n875), .ZN(n877) );
  XOR2_X1 U976 ( .A(n878), .B(n877), .Z(n896) );
  NAND2_X1 U977 ( .A1(G139), .A2(n879), .ZN(n880) );
  XNOR2_X1 U978 ( .A(n880), .B(KEYINPUT116), .ZN(n884) );
  NAND2_X1 U979 ( .A1(G103), .A2(n881), .ZN(n882) );
  XOR2_X1 U980 ( .A(KEYINPUT115), .B(n882), .Z(n883) );
  NAND2_X1 U981 ( .A1(n884), .A2(n883), .ZN(n893) );
  NAND2_X1 U982 ( .A1(n885), .A2(G127), .ZN(n886) );
  XNOR2_X1 U983 ( .A(KEYINPUT117), .B(n886), .ZN(n890) );
  NAND2_X1 U984 ( .A1(n887), .A2(G115), .ZN(n888) );
  XOR2_X1 U985 ( .A(KEYINPUT118), .B(n888), .Z(n889) );
  NOR2_X1 U986 ( .A1(n890), .A2(n889), .ZN(n891) );
  XNOR2_X1 U987 ( .A(n891), .B(KEYINPUT47), .ZN(n892) );
  NOR2_X1 U988 ( .A1(n893), .A2(n892), .ZN(n1009) );
  XOR2_X1 U989 ( .A(n894), .B(n1009), .Z(n895) );
  XNOR2_X1 U990 ( .A(n896), .B(n895), .ZN(n901) );
  XOR2_X1 U991 ( .A(KEYINPUT119), .B(KEYINPUT46), .Z(n898) );
  XNOR2_X1 U992 ( .A(n1002), .B(KEYINPUT48), .ZN(n897) );
  XNOR2_X1 U993 ( .A(n898), .B(n897), .ZN(n899) );
  XOR2_X1 U994 ( .A(G164), .B(n899), .Z(n900) );
  XNOR2_X1 U995 ( .A(n901), .B(n900), .ZN(n902) );
  NOR2_X1 U996 ( .A1(G37), .A2(n902), .ZN(G395) );
  XOR2_X1 U997 ( .A(n903), .B(G286), .Z(n905) );
  XNOR2_X1 U998 ( .A(n937), .B(G171), .ZN(n904) );
  XNOR2_X1 U999 ( .A(n905), .B(n904), .ZN(n906) );
  NOR2_X1 U1000 ( .A1(G37), .A2(n906), .ZN(G397) );
  XNOR2_X1 U1001 ( .A(G2435), .B(G2443), .ZN(n916) );
  XOR2_X1 U1002 ( .A(G2454), .B(G2430), .Z(n908) );
  XNOR2_X1 U1003 ( .A(G2446), .B(KEYINPUT109), .ZN(n907) );
  XNOR2_X1 U1004 ( .A(n908), .B(n907), .ZN(n912) );
  XOR2_X1 U1005 ( .A(G2451), .B(G2427), .Z(n910) );
  XNOR2_X1 U1006 ( .A(G1348), .B(G1341), .ZN(n909) );
  XNOR2_X1 U1007 ( .A(n910), .B(n909), .ZN(n911) );
  XOR2_X1 U1008 ( .A(n912), .B(n911), .Z(n914) );
  XNOR2_X1 U1009 ( .A(KEYINPUT108), .B(G2438), .ZN(n913) );
  XNOR2_X1 U1010 ( .A(n914), .B(n913), .ZN(n915) );
  XNOR2_X1 U1011 ( .A(n916), .B(n915), .ZN(n917) );
  NAND2_X1 U1012 ( .A1(n917), .A2(G14), .ZN(n923) );
  NAND2_X1 U1013 ( .A1(G319), .A2(n923), .ZN(n920) );
  NOR2_X1 U1014 ( .A1(G227), .A2(G229), .ZN(n918) );
  XNOR2_X1 U1015 ( .A(KEYINPUT49), .B(n918), .ZN(n919) );
  NOR2_X1 U1016 ( .A1(n920), .A2(n919), .ZN(n922) );
  NOR2_X1 U1017 ( .A1(G395), .A2(G397), .ZN(n921) );
  NAND2_X1 U1018 ( .A1(n922), .A2(n921), .ZN(G225) );
  INV_X1 U1019 ( .A(G225), .ZN(G308) );
  INV_X1 U1020 ( .A(G57), .ZN(G237) );
  INV_X1 U1021 ( .A(n923), .ZN(G401) );
  NAND2_X1 U1022 ( .A1(G1971), .A2(G303), .ZN(n924) );
  NAND2_X1 U1023 ( .A1(n925), .A2(n924), .ZN(n926) );
  NOR2_X1 U1024 ( .A1(n927), .A2(n926), .ZN(n933) );
  XNOR2_X1 U1025 ( .A(G171), .B(G1961), .ZN(n929) );
  NAND2_X1 U1026 ( .A1(n929), .A2(n928), .ZN(n931) );
  XNOR2_X1 U1027 ( .A(G1956), .B(G299), .ZN(n930) );
  NOR2_X1 U1028 ( .A1(n931), .A2(n930), .ZN(n932) );
  NAND2_X1 U1029 ( .A1(n933), .A2(n932), .ZN(n944) );
  XNOR2_X1 U1030 ( .A(G1966), .B(G168), .ZN(n935) );
  NAND2_X1 U1031 ( .A1(n935), .A2(n934), .ZN(n936) );
  XNOR2_X1 U1032 ( .A(n936), .B(KEYINPUT57), .ZN(n942) );
  XOR2_X1 U1033 ( .A(G1348), .B(n937), .Z(n940) );
  XNOR2_X1 U1034 ( .A(n938), .B(G1341), .ZN(n939) );
  NOR2_X1 U1035 ( .A1(n940), .A2(n939), .ZN(n941) );
  NAND2_X1 U1036 ( .A1(n942), .A2(n941), .ZN(n943) );
  NOR2_X1 U1037 ( .A1(n944), .A2(n943), .ZN(n945) );
  XOR2_X1 U1038 ( .A(KEYINPUT124), .B(n945), .Z(n947) );
  XNOR2_X1 U1039 ( .A(G16), .B(KEYINPUT56), .ZN(n946) );
  NAND2_X1 U1040 ( .A1(n947), .A2(n946), .ZN(n1026) );
  XNOR2_X1 U1041 ( .A(G16), .B(KEYINPUT125), .ZN(n972) );
  XNOR2_X1 U1042 ( .A(G1348), .B(KEYINPUT59), .ZN(n948) );
  XNOR2_X1 U1043 ( .A(n948), .B(G4), .ZN(n952) );
  XNOR2_X1 U1044 ( .A(G1341), .B(G19), .ZN(n950) );
  XNOR2_X1 U1045 ( .A(G1981), .B(G6), .ZN(n949) );
  NOR2_X1 U1046 ( .A1(n950), .A2(n949), .ZN(n951) );
  NAND2_X1 U1047 ( .A1(n952), .A2(n951), .ZN(n956) );
  XOR2_X1 U1048 ( .A(G20), .B(n953), .Z(n954) );
  XNOR2_X1 U1049 ( .A(KEYINPUT126), .B(n954), .ZN(n955) );
  NOR2_X1 U1050 ( .A1(n956), .A2(n955), .ZN(n957) );
  XNOR2_X1 U1051 ( .A(KEYINPUT60), .B(n957), .ZN(n961) );
  XNOR2_X1 U1052 ( .A(G1966), .B(G21), .ZN(n959) );
  XNOR2_X1 U1053 ( .A(G5), .B(G1961), .ZN(n958) );
  NOR2_X1 U1054 ( .A1(n959), .A2(n958), .ZN(n960) );
  NAND2_X1 U1055 ( .A1(n961), .A2(n960), .ZN(n968) );
  XNOR2_X1 U1056 ( .A(G1971), .B(G22), .ZN(n963) );
  XNOR2_X1 U1057 ( .A(G23), .B(G1976), .ZN(n962) );
  NOR2_X1 U1058 ( .A1(n963), .A2(n962), .ZN(n965) );
  XOR2_X1 U1059 ( .A(G1986), .B(G24), .Z(n964) );
  NAND2_X1 U1060 ( .A1(n965), .A2(n964), .ZN(n966) );
  XNOR2_X1 U1061 ( .A(KEYINPUT58), .B(n966), .ZN(n967) );
  NOR2_X1 U1062 ( .A1(n968), .A2(n967), .ZN(n969) );
  XOR2_X1 U1063 ( .A(n969), .B(KEYINPUT61), .Z(n970) );
  XNOR2_X1 U1064 ( .A(KEYINPUT127), .B(n970), .ZN(n971) );
  NAND2_X1 U1065 ( .A1(n972), .A2(n971), .ZN(n997) );
  INV_X1 U1066 ( .A(G29), .ZN(n1021) );
  XOR2_X1 U1067 ( .A(KEYINPUT55), .B(KEYINPUT122), .Z(n992) );
  XNOR2_X1 U1068 ( .A(G2090), .B(G35), .ZN(n987) );
  XNOR2_X1 U1069 ( .A(KEYINPUT121), .B(G1996), .ZN(n973) );
  XNOR2_X1 U1070 ( .A(n973), .B(G32), .ZN(n979) );
  XOR2_X1 U1071 ( .A(G1991), .B(G25), .Z(n974) );
  NAND2_X1 U1072 ( .A1(n974), .A2(G28), .ZN(n977) );
  XNOR2_X1 U1073 ( .A(G27), .B(n975), .ZN(n976) );
  NOR2_X1 U1074 ( .A1(n977), .A2(n976), .ZN(n978) );
  NAND2_X1 U1075 ( .A1(n979), .A2(n978), .ZN(n984) );
  XNOR2_X1 U1076 ( .A(G2067), .B(G26), .ZN(n981) );
  XNOR2_X1 U1077 ( .A(G2072), .B(G33), .ZN(n980) );
  NOR2_X1 U1078 ( .A1(n981), .A2(n980), .ZN(n982) );
  XOR2_X1 U1079 ( .A(KEYINPUT120), .B(n982), .Z(n983) );
  NOR2_X1 U1080 ( .A1(n984), .A2(n983), .ZN(n985) );
  XNOR2_X1 U1081 ( .A(KEYINPUT53), .B(n985), .ZN(n986) );
  NOR2_X1 U1082 ( .A1(n987), .A2(n986), .ZN(n990) );
  XOR2_X1 U1083 ( .A(G2084), .B(G34), .Z(n988) );
  XNOR2_X1 U1084 ( .A(KEYINPUT54), .B(n988), .ZN(n989) );
  NAND2_X1 U1085 ( .A1(n990), .A2(n989), .ZN(n991) );
  XNOR2_X1 U1086 ( .A(n992), .B(n991), .ZN(n993) );
  NAND2_X1 U1087 ( .A1(n1021), .A2(n993), .ZN(n994) );
  NAND2_X1 U1088 ( .A1(n994), .A2(G11), .ZN(n995) );
  XNOR2_X1 U1089 ( .A(n995), .B(KEYINPUT123), .ZN(n996) );
  NAND2_X1 U1090 ( .A1(n997), .A2(n996), .ZN(n1024) );
  XNOR2_X1 U1091 ( .A(G2090), .B(G162), .ZN(n999) );
  NAND2_X1 U1092 ( .A1(n999), .A2(n998), .ZN(n1000) );
  XNOR2_X1 U1093 ( .A(n1000), .B(KEYINPUT51), .ZN(n1004) );
  XOR2_X1 U1094 ( .A(G2084), .B(G160), .Z(n1001) );
  NOR2_X1 U1095 ( .A1(n1002), .A2(n1001), .ZN(n1003) );
  NAND2_X1 U1096 ( .A1(n1004), .A2(n1003), .ZN(n1005) );
  NOR2_X1 U1097 ( .A1(n1006), .A2(n1005), .ZN(n1007) );
  NAND2_X1 U1098 ( .A1(n1008), .A2(n1007), .ZN(n1014) );
  XOR2_X1 U1099 ( .A(G2072), .B(n1009), .Z(n1011) );
  XOR2_X1 U1100 ( .A(G164), .B(G2078), .Z(n1010) );
  NOR2_X1 U1101 ( .A1(n1011), .A2(n1010), .ZN(n1012) );
  XOR2_X1 U1102 ( .A(KEYINPUT50), .B(n1012), .Z(n1013) );
  NOR2_X1 U1103 ( .A1(n1014), .A2(n1013), .ZN(n1015) );
  NAND2_X1 U1104 ( .A1(n1016), .A2(n1015), .ZN(n1017) );
  NOR2_X1 U1105 ( .A1(n1018), .A2(n1017), .ZN(n1019) );
  XOR2_X1 U1106 ( .A(KEYINPUT52), .B(n1019), .Z(n1020) );
  NOR2_X1 U1107 ( .A1(KEYINPUT55), .A2(n1020), .ZN(n1022) );
  NOR2_X1 U1108 ( .A1(n1022), .A2(n1021), .ZN(n1023) );
  NOR2_X1 U1109 ( .A1(n1024), .A2(n1023), .ZN(n1025) );
  NAND2_X1 U1110 ( .A1(n1026), .A2(n1025), .ZN(n1027) );
  XOR2_X1 U1111 ( .A(KEYINPUT62), .B(n1027), .Z(G311) );
  INV_X1 U1112 ( .A(G311), .ZN(G150) );
endmodule

