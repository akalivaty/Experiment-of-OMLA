

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n350, n351, n352, n353, n354, n355, n356, n357, n358, n359, n360,
         n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, n371,
         n372, n373, n374, n375, n376, n377, n378, n379, n380, n381, n382,
         n383, n384, n385, n386, n387, n388, n389, n390, n391, n392, n393,
         n394, n395, n396, n397, n398, n399, n400, n401, n402, n403, n404,
         n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, n415,
         n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426,
         n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437,
         n438, n439, n440, n441, n442, n443, n444, n445, n446, n447, n448,
         n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, n459,
         n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, n470,
         n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481,
         n482, n483, n484, n485, n486, n487, n488, n489, n490, n491, n492,
         n493, n494, n495, n496, n497, n498, n499, n500, n501, n502, n503,
         n504, n505, n506, n507, n508, n509, n510, n511, n512, n513, n514,
         n515, n516, n517, n518, n519, n520, n521, n522, n523, n524, n525,
         n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536,
         n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547,
         n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558,
         n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569,
         n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580,
         n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591,
         n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602,
         n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, n613,
         n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624,
         n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635,
         n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, n646,
         n647, n648, n649, n650, n651, n652, n653, n654, n655, n656, n657,
         n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668,
         n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679,
         n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690,
         n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701,
         n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712,
         n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723,
         n724, n725, n726, n727, n728, n729, n730, n731, n732;

  NOR2_X1 U371 ( .A1(n551), .A2(n350), .ZN(n399) );
  INV_X1 U372 ( .A(G953), .ZN(n721) );
  XNOR2_X2 U373 ( .A(n459), .B(n458), .ZN(n588) );
  XNOR2_X2 U374 ( .A(n505), .B(KEYINPUT33), .ZN(n678) );
  AND2_X2 U375 ( .A1(n567), .A2(n382), .ZN(n505) );
  NOR2_X2 U376 ( .A1(n551), .A2(n678), .ZN(n506) );
  XNOR2_X2 U377 ( .A(n466), .B(KEYINPUT0), .ZN(n551) );
  AND2_X1 U378 ( .A1(n366), .A2(n365), .ZN(n409) );
  NOR2_X1 U379 ( .A1(n606), .A2(n701), .ZN(n608) );
  XNOR2_X1 U380 ( .A(n411), .B(n410), .ZN(n731) );
  NOR2_X1 U381 ( .A1(n730), .A2(n624), .ZN(n540) );
  XNOR2_X1 U382 ( .A(n579), .B(KEYINPUT42), .ZN(n732) );
  NOR2_X1 U383 ( .A1(n575), .A2(n658), .ZN(n581) );
  NAND2_X1 U384 ( .A1(n416), .A2(n413), .ZN(n658) );
  INV_X1 U385 ( .A(n563), .ZN(n416) );
  XNOR2_X1 U386 ( .A(n495), .B(n494), .ZN(n563) );
  XNOR2_X1 U387 ( .A(n420), .B(G128), .ZN(n468) );
  XNOR2_X1 U388 ( .A(n355), .B(n449), .ZN(n500) );
  XNOR2_X1 U389 ( .A(G104), .B(G110), .ZN(n406) );
  XOR2_X1 U390 ( .A(KEYINPUT69), .B(G140), .Z(n484) );
  XOR2_X1 U391 ( .A(G122), .B(KEYINPUT16), .Z(n450) );
  INV_X1 U392 ( .A(G143), .ZN(n420) );
  NAND2_X1 U393 ( .A1(n393), .A2(n593), .ZN(n392) );
  NOR2_X1 U394 ( .A1(n731), .A2(n732), .ZN(n396) );
  XNOR2_X1 U395 ( .A(n434), .B(G146), .ZN(n478) );
  INV_X1 U396 ( .A(G125), .ZN(n434) );
  XNOR2_X1 U397 ( .A(n446), .B(n445), .ZN(n572) );
  INV_X1 U398 ( .A(KEYINPUT71), .ZN(n445) );
  NOR2_X1 U399 ( .A1(n582), .A2(n448), .ZN(n447) );
  XOR2_X1 U400 ( .A(G475), .B(n519), .Z(n546) );
  OR2_X1 U401 ( .A1(n689), .A2(G902), .ZN(n477) );
  INV_X1 U402 ( .A(n592), .ZN(n384) );
  XNOR2_X1 U403 ( .A(n432), .B(KEYINPUT85), .ZN(n431) );
  XNOR2_X1 U404 ( .A(n492), .B(n491), .ZN(n496) );
  XOR2_X1 U405 ( .A(KEYINPUT20), .B(KEYINPUT93), .Z(n492) );
  NAND2_X1 U406 ( .A1(n496), .A2(G217), .ZN(n493) );
  XNOR2_X1 U407 ( .A(n520), .B(n471), .ZN(n499) );
  XNOR2_X1 U408 ( .A(n470), .B(n469), .ZN(n471) );
  INV_X1 U409 ( .A(G137), .ZN(n469) );
  XNOR2_X1 U410 ( .A(KEYINPUT4), .B(KEYINPUT67), .ZN(n719) );
  XNOR2_X1 U411 ( .A(n473), .B(n376), .ZN(n498) );
  INV_X1 U412 ( .A(G146), .ZN(n376) );
  XNOR2_X1 U413 ( .A(n499), .B(n419), .ZN(n716) );
  INV_X1 U414 ( .A(n484), .ZN(n419) );
  XNOR2_X1 U415 ( .A(n719), .B(n367), .ZN(n473) );
  XNOR2_X1 U416 ( .A(KEYINPUT66), .B(G101), .ZN(n367) );
  NAND2_X1 U417 ( .A1(n387), .A2(n385), .ZN(n598) );
  AND2_X1 U418 ( .A1(n390), .A2(n388), .ZN(n387) );
  INV_X1 U419 ( .A(KEYINPUT96), .ZN(n414) );
  NOR2_X1 U420 ( .A1(n559), .A2(n377), .ZN(n560) );
  NAND2_X1 U421 ( .A1(G953), .A2(n378), .ZN(n377) );
  XNOR2_X1 U422 ( .A(n375), .B(n373), .ZN(n603) );
  XNOR2_X1 U423 ( .A(n374), .B(n500), .ZN(n373) );
  XNOR2_X1 U424 ( .A(n499), .B(n498), .ZN(n375) );
  XNOR2_X1 U425 ( .A(n503), .B(n359), .ZN(n374) );
  NOR2_X1 U426 ( .A1(n573), .A2(n572), .ZN(n574) );
  NAND2_X1 U427 ( .A1(n380), .A2(n379), .ZN(n381) );
  AND2_X1 U428 ( .A1(n584), .A2(n647), .ZN(n379) );
  INV_X1 U429 ( .A(KEYINPUT1), .ZN(n429) );
  XNOR2_X1 U430 ( .A(n488), .B(n489), .ZN(n700) );
  INV_X1 U431 ( .A(KEYINPUT123), .ZN(n443) );
  NAND2_X1 U432 ( .A1(n352), .A2(n384), .ZN(n393) );
  NOR2_X1 U433 ( .A1(G953), .A2(G237), .ZN(n510) );
  NAND2_X1 U434 ( .A1(n636), .A2(n618), .ZN(n427) );
  INV_X1 U435 ( .A(n641), .ZN(n397) );
  NOR2_X1 U436 ( .A1(n644), .A2(KEYINPUT48), .ZN(n435) );
  NOR2_X1 U437 ( .A1(n596), .A2(n436), .ZN(n438) );
  XNOR2_X1 U438 ( .A(n415), .B(n497), .ZN(n661) );
  NAND2_X1 U439 ( .A1(n496), .A2(G221), .ZN(n415) );
  OR2_X1 U440 ( .A1(G237), .A2(G902), .ZN(n457) );
  INV_X1 U441 ( .A(G900), .ZN(n378) );
  NAND2_X1 U442 ( .A1(n462), .A2(G902), .ZN(n559) );
  XNOR2_X1 U443 ( .A(KEYINPUT77), .B(KEYINPUT97), .ZN(n501) );
  AND2_X1 U444 ( .A1(n545), .A2(n616), .ZN(n555) );
  XNOR2_X1 U445 ( .A(KEYINPUT105), .B(n553), .ZN(n554) );
  AND2_X1 U446 ( .A1(n426), .A2(n425), .ZN(n553) );
  INV_X1 U447 ( .A(n651), .ZN(n425) );
  XNOR2_X1 U448 ( .A(n427), .B(KEYINPUT100), .ZN(n426) );
  XOR2_X1 U449 ( .A(G140), .B(G122), .Z(n508) );
  XNOR2_X1 U450 ( .A(G113), .B(G104), .ZN(n507) );
  XNOR2_X1 U451 ( .A(n369), .B(n512), .ZN(n514) );
  XOR2_X1 U452 ( .A(KEYINPUT12), .B(KEYINPUT11), .Z(n512) );
  XNOR2_X1 U453 ( .A(n511), .B(n370), .ZN(n369) );
  INV_X1 U454 ( .A(KEYINPUT101), .ZN(n370) );
  XNOR2_X1 U455 ( .A(G143), .B(G131), .ZN(n513) );
  XNOR2_X1 U456 ( .A(n461), .B(n460), .ZN(n462) );
  NAND2_X1 U457 ( .A1(G234), .A2(G237), .ZN(n460) );
  XOR2_X1 U458 ( .A(KEYINPUT75), .B(KEYINPUT14), .Z(n461) );
  XNOR2_X1 U459 ( .A(n493), .B(n354), .ZN(n494) );
  NOR2_X1 U460 ( .A1(G902), .A2(n700), .ZN(n495) );
  XNOR2_X1 U461 ( .A(n478), .B(n433), .ZN(n715) );
  XNOR2_X1 U462 ( .A(KEYINPUT68), .B(KEYINPUT10), .ZN(n433) );
  XNOR2_X1 U463 ( .A(n468), .B(n467), .ZN(n520) );
  INV_X1 U464 ( .A(G134), .ZN(n467) );
  XNOR2_X1 U465 ( .A(G116), .B(G107), .ZN(n524) );
  XNOR2_X1 U466 ( .A(n418), .B(n417), .ZN(n599) );
  INV_X1 U467 ( .A(KEYINPUT90), .ZN(n417) );
  XNOR2_X1 U468 ( .A(G902), .B(KEYINPUT15), .ZN(n418) );
  XNOR2_X1 U469 ( .A(n498), .B(n368), .ZN(n372) );
  XNOR2_X1 U470 ( .A(n472), .B(n474), .ZN(n368) );
  XNOR2_X1 U471 ( .A(n394), .B(n455), .ZN(n612) );
  XNOR2_X1 U472 ( .A(n710), .B(n395), .ZN(n394) );
  XNOR2_X1 U473 ( .A(n453), .B(n452), .ZN(n454) );
  NAND2_X1 U474 ( .A1(n598), .A2(n358), .ZN(n371) );
  XNOR2_X1 U475 ( .A(n399), .B(n362), .ZN(n538) );
  AND2_X1 U476 ( .A1(n567), .A2(n428), .ZN(n549) );
  INV_X1 U477 ( .A(n658), .ZN(n428) );
  XNOR2_X1 U478 ( .A(n412), .B(KEYINPUT78), .ZN(n380) );
  NOR2_X1 U479 ( .A1(n583), .A2(n582), .ZN(n412) );
  XNOR2_X1 U480 ( .A(n589), .B(KEYINPUT80), .ZN(n625) );
  INV_X1 U481 ( .A(KEYINPUT6), .ZN(n408) );
  XNOR2_X1 U482 ( .A(n603), .B(n602), .ZN(n604) );
  INV_X1 U483 ( .A(KEYINPUT40), .ZN(n410) );
  XNOR2_X1 U484 ( .A(n534), .B(n533), .ZN(n730) );
  XNOR2_X1 U485 ( .A(KEYINPUT86), .B(KEYINPUT35), .ZN(n533) );
  XNOR2_X1 U486 ( .A(n401), .B(n400), .ZN(n729) );
  INV_X1 U487 ( .A(KEYINPUT32), .ZN(n400) );
  NOR2_X1 U488 ( .A1(n538), .A2(n403), .ZN(n401) );
  NAND2_X1 U489 ( .A1(n539), .A2(n567), .ZN(n403) );
  XNOR2_X1 U490 ( .A(n550), .B(KEYINPUT31), .ZN(n636) );
  NOR2_X1 U491 ( .A1(n551), .A2(n667), .ZN(n550) );
  AND2_X1 U492 ( .A1(n543), .A2(n405), .ZN(n624) );
  NOR2_X1 U493 ( .A1(n664), .A2(n416), .ZN(n405) );
  XNOR2_X1 U494 ( .A(n444), .B(n442), .ZN(n441) );
  NAND2_X1 U495 ( .A1(n699), .A2(G217), .ZN(n444) );
  XNOR2_X1 U496 ( .A(n696), .B(n404), .ZN(n698) );
  XNOR2_X1 U497 ( .A(n697), .B(KEYINPUT122), .ZN(n404) );
  INV_X1 U498 ( .A(KEYINPUT60), .ZN(n421) );
  INV_X1 U499 ( .A(G143), .ZN(n383) );
  NAND2_X1 U500 ( .A1(n536), .A2(n413), .ZN(n350) );
  INV_X1 U501 ( .A(n644), .ZN(n439) );
  XOR2_X1 U502 ( .A(n695), .B(n364), .Z(n351) );
  AND2_X1 U503 ( .A1(n591), .A2(n590), .ZN(n352) );
  AND2_X1 U504 ( .A1(G210), .A2(n457), .ZN(n353) );
  XOR2_X1 U505 ( .A(KEYINPUT94), .B(KEYINPUT25), .Z(n354) );
  XOR2_X1 U506 ( .A(G113), .B(G116), .Z(n355) );
  XOR2_X1 U507 ( .A(G472), .B(KEYINPUT99), .Z(n356) );
  XNOR2_X1 U508 ( .A(n661), .B(n414), .ZN(n535) );
  INV_X1 U509 ( .A(n535), .ZN(n413) );
  AND2_X1 U510 ( .A1(n588), .A2(n576), .ZN(n357) );
  AND2_X1 U511 ( .A1(n643), .A2(KEYINPUT2), .ZN(n358) );
  AND2_X1 U512 ( .A1(n510), .A2(G210), .ZN(n359) );
  AND2_X1 U513 ( .A1(n439), .A2(n436), .ZN(n360) );
  XOR2_X1 U514 ( .A(KEYINPUT38), .B(KEYINPUT76), .Z(n361) );
  XOR2_X1 U515 ( .A(KEYINPUT22), .B(KEYINPUT64), .Z(n362) );
  XOR2_X1 U516 ( .A(n612), .B(n611), .Z(n363) );
  NOR2_X1 U517 ( .A1(G952), .A2(n721), .ZN(n701) );
  INV_X1 U518 ( .A(n701), .ZN(n365) );
  XNOR2_X1 U519 ( .A(KEYINPUT59), .B(KEYINPUT89), .ZN(n364) );
  NOR2_X1 U520 ( .A1(n542), .A2(KEYINPUT44), .ZN(n541) );
  XNOR2_X1 U521 ( .A(n613), .B(n363), .ZN(n366) );
  NAND2_X1 U522 ( .A1(n682), .A2(n599), .ZN(n601) );
  NOR2_X2 U523 ( .A1(n706), .A2(n720), .ZN(n600) );
  NOR2_X2 U524 ( .A1(n557), .A2(n556), .ZN(n558) );
  XNOR2_X2 U525 ( .A(n558), .B(KEYINPUT45), .ZN(n706) );
  XNOR2_X1 U526 ( .A(n372), .B(n716), .ZN(n689) );
  NAND2_X1 U527 ( .A1(n598), .A2(n643), .ZN(n720) );
  OR2_X2 U528 ( .A1(n706), .A2(n371), .ZN(n682) );
  NOR2_X1 U529 ( .A1(n389), .A2(n644), .ZN(n437) );
  NAND2_X1 U530 ( .A1(n398), .A2(n397), .ZN(n389) );
  NAND2_X1 U531 ( .A1(n577), .A2(n576), .ZN(n578) );
  NAND2_X1 U532 ( .A1(n577), .A2(n357), .ZN(n589) );
  AND2_X1 U533 ( .A1(n380), .A2(n584), .ZN(n591) );
  XNOR2_X2 U534 ( .A(n381), .B(KEYINPUT39), .ZN(n597) );
  INV_X1 U535 ( .A(n567), .ZN(n657) );
  NOR2_X1 U536 ( .A1(n564), .A2(n658), .ZN(n382) );
  XNOR2_X2 U537 ( .A(n573), .B(n408), .ZN(n564) );
  XNOR2_X2 U538 ( .A(n504), .B(n356), .ZN(n573) );
  XNOR2_X2 U539 ( .A(n575), .B(n429), .ZN(n567) );
  XNOR2_X2 U540 ( .A(n477), .B(n476), .ZN(n575) );
  XNOR2_X1 U541 ( .A(n393), .B(n383), .ZN(n630) );
  NAND2_X1 U542 ( .A1(n437), .A2(n386), .ZN(n385) );
  AND2_X1 U543 ( .A1(n594), .A2(n438), .ZN(n386) );
  NAND2_X1 U544 ( .A1(n389), .A2(n360), .ZN(n388) );
  NAND2_X1 U545 ( .A1(n391), .A2(n435), .ZN(n390) );
  NAND2_X1 U546 ( .A1(n594), .A2(n440), .ZN(n391) );
  NOR2_X1 U547 ( .A1(n431), .A2(n392), .ZN(n430) );
  XNOR2_X1 U548 ( .A(n451), .B(n468), .ZN(n395) );
  XNOR2_X1 U549 ( .A(n396), .B(KEYINPUT46), .ZN(n594) );
  XNOR2_X1 U550 ( .A(n430), .B(KEYINPUT84), .ZN(n398) );
  XNOR2_X1 U551 ( .A(n402), .B(KEYINPUT41), .ZN(n677) );
  NOR2_X1 U552 ( .A1(n652), .A2(n650), .ZN(n402) );
  NOR2_X2 U553 ( .A1(n600), .A2(KEYINPUT2), .ZN(n681) );
  NOR2_X4 U554 ( .A1(n601), .A2(n681), .ZN(n699) );
  NAND2_X1 U555 ( .A1(n540), .A2(n729), .ZN(n542) );
  XNOR2_X2 U556 ( .A(n406), .B(G107), .ZN(n472) );
  XNOR2_X2 U557 ( .A(n407), .B(n500), .ZN(n710) );
  XNOR2_X2 U558 ( .A(n472), .B(n450), .ZN(n407) );
  XNOR2_X1 U559 ( .A(n409), .B(n615), .ZN(G51) );
  NAND2_X1 U560 ( .A1(n647), .A2(n646), .ZN(n571) );
  XNOR2_X1 U561 ( .A(n570), .B(n361), .ZN(n647) );
  NAND2_X1 U562 ( .A1(n597), .A2(n631), .ZN(n411) );
  XNOR2_X1 U563 ( .A(n422), .B(n421), .ZN(G60) );
  NAND2_X1 U564 ( .A1(n423), .A2(n365), .ZN(n422) );
  XNOR2_X1 U565 ( .A(n424), .B(n351), .ZN(n423) );
  NAND2_X1 U566 ( .A1(n699), .A2(G475), .ZN(n424) );
  NAND2_X1 U567 ( .A1(n625), .A2(KEYINPUT47), .ZN(n432) );
  INV_X1 U568 ( .A(KEYINPUT48), .ZN(n436) );
  INV_X1 U569 ( .A(n596), .ZN(n440) );
  NOR2_X1 U570 ( .A1(n441), .A2(n701), .ZN(G66) );
  XNOR2_X1 U571 ( .A(n700), .B(n443), .ZN(n442) );
  NAND2_X1 U572 ( .A1(n563), .A2(n447), .ZN(n446) );
  INV_X1 U573 ( .A(n661), .ZN(n448) );
  INV_X1 U574 ( .A(KEYINPUT17), .ZN(n452) );
  XNOR2_X1 U575 ( .A(n482), .B(n481), .ZN(n483) );
  INV_X1 U576 ( .A(n625), .ZN(n632) );
  INV_X1 U577 ( .A(KEYINPUT63), .ZN(n607) );
  XNOR2_X1 U578 ( .A(G119), .B(KEYINPUT3), .ZN(n449) );
  AND2_X1 U579 ( .A1(G224), .A2(n721), .ZN(n451) );
  XNOR2_X1 U580 ( .A(n478), .B(KEYINPUT18), .ZN(n453) );
  XNOR2_X1 U581 ( .A(n473), .B(n454), .ZN(n455) );
  INV_X1 U582 ( .A(n599), .ZN(n490) );
  NAND2_X1 U583 ( .A1(n612), .A2(n490), .ZN(n456) );
  XNOR2_X2 U584 ( .A(n456), .B(n353), .ZN(n570) );
  NAND2_X1 U585 ( .A1(G214), .A2(n457), .ZN(n646) );
  NAND2_X1 U586 ( .A1(n570), .A2(n646), .ZN(n459) );
  XOR2_X1 U587 ( .A(KEYINPUT19), .B(KEYINPUT65), .Z(n458) );
  NAND2_X1 U588 ( .A1(G952), .A2(n462), .ZN(n676) );
  NOR2_X1 U589 ( .A1(G953), .A2(n676), .ZN(n561) );
  INV_X1 U590 ( .A(G898), .ZN(n704) );
  NAND2_X1 U591 ( .A1(G953), .A2(n704), .ZN(n711) );
  NOR2_X1 U592 ( .A1(n559), .A2(n711), .ZN(n463) );
  NOR2_X1 U593 ( .A1(n561), .A2(n463), .ZN(n464) );
  XNOR2_X1 U594 ( .A(KEYINPUT91), .B(n464), .ZN(n465) );
  NAND2_X1 U595 ( .A1(n588), .A2(n465), .ZN(n466) );
  XNOR2_X1 U596 ( .A(G131), .B(KEYINPUT70), .ZN(n470) );
  AND2_X1 U597 ( .A1(G227), .A2(n721), .ZN(n474) );
  XNOR2_X1 U598 ( .A(G469), .B(KEYINPUT72), .ZN(n475) );
  XNOR2_X1 U599 ( .A(n475), .B(KEYINPUT73), .ZN(n476) );
  XOR2_X1 U600 ( .A(G110), .B(G119), .Z(n480) );
  XNOR2_X1 U601 ( .A(G137), .B(G128), .ZN(n479) );
  XNOR2_X1 U602 ( .A(n480), .B(n479), .ZN(n482) );
  XOR2_X1 U603 ( .A(KEYINPUT23), .B(KEYINPUT24), .Z(n481) );
  XNOR2_X1 U604 ( .A(n715), .B(n483), .ZN(n489) );
  XOR2_X1 U605 ( .A(n484), .B(KEYINPUT92), .Z(n487) );
  NAND2_X1 U606 ( .A1(G234), .A2(n721), .ZN(n485) );
  XOR2_X1 U607 ( .A(KEYINPUT8), .B(n485), .Z(n528) );
  NAND2_X1 U608 ( .A1(G221), .A2(n528), .ZN(n486) );
  XNOR2_X1 U609 ( .A(n487), .B(n486), .ZN(n488) );
  NAND2_X1 U610 ( .A1(G234), .A2(n490), .ZN(n491) );
  XNOR2_X1 U611 ( .A(KEYINPUT95), .B(KEYINPUT21), .ZN(n497) );
  XOR2_X1 U612 ( .A(KEYINPUT98), .B(KEYINPUT5), .Z(n502) );
  XNOR2_X1 U613 ( .A(n502), .B(n501), .ZN(n503) );
  NOR2_X1 U614 ( .A1(G902), .A2(n603), .ZN(n504) );
  XNOR2_X1 U615 ( .A(n506), .B(KEYINPUT34), .ZN(n532) );
  XNOR2_X1 U616 ( .A(KEYINPUT102), .B(KEYINPUT13), .ZN(n518) );
  XNOR2_X1 U617 ( .A(n508), .B(n507), .ZN(n509) );
  XNOR2_X1 U618 ( .A(n715), .B(n509), .ZN(n516) );
  NAND2_X1 U619 ( .A1(G214), .A2(n510), .ZN(n511) );
  XNOR2_X1 U620 ( .A(n514), .B(n513), .ZN(n515) );
  XNOR2_X1 U621 ( .A(n516), .B(n515), .ZN(n695) );
  NOR2_X1 U622 ( .A1(G902), .A2(n695), .ZN(n517) );
  XNOR2_X1 U623 ( .A(n518), .B(n517), .ZN(n519) );
  INV_X1 U624 ( .A(n520), .ZN(n527) );
  XOR2_X1 U625 ( .A(KEYINPUT7), .B(KEYINPUT103), .Z(n522) );
  XNOR2_X1 U626 ( .A(G122), .B(KEYINPUT104), .ZN(n521) );
  XNOR2_X1 U627 ( .A(n522), .B(n521), .ZN(n523) );
  XOR2_X1 U628 ( .A(n523), .B(KEYINPUT9), .Z(n525) );
  XNOR2_X1 U629 ( .A(n525), .B(n524), .ZN(n526) );
  XNOR2_X1 U630 ( .A(n527), .B(n526), .ZN(n530) );
  NAND2_X1 U631 ( .A1(G217), .A2(n528), .ZN(n529) );
  XNOR2_X1 U632 ( .A(n530), .B(n529), .ZN(n697) );
  NOR2_X1 U633 ( .A1(n697), .A2(G902), .ZN(n531) );
  XNOR2_X1 U634 ( .A(n531), .B(G478), .ZN(n548) );
  NOR2_X1 U635 ( .A1(n546), .A2(n548), .ZN(n590) );
  NAND2_X1 U636 ( .A1(n532), .A2(n590), .ZN(n534) );
  INV_X1 U637 ( .A(n573), .ZN(n664) );
  NAND2_X1 U638 ( .A1(n546), .A2(n548), .ZN(n650) );
  INV_X1 U639 ( .A(n650), .ZN(n536) );
  NOR2_X1 U640 ( .A1(n538), .A2(n567), .ZN(n543) );
  XOR2_X1 U641 ( .A(KEYINPUT106), .B(n563), .Z(n660) );
  XNOR2_X1 U642 ( .A(KEYINPUT79), .B(n564), .ZN(n537) );
  NOR2_X1 U643 ( .A1(n660), .A2(n537), .ZN(n539) );
  XNOR2_X1 U644 ( .A(n541), .B(KEYINPUT74), .ZN(n557) );
  NAND2_X1 U645 ( .A1(n542), .A2(KEYINPUT44), .ZN(n545) );
  AND2_X1 U646 ( .A1(n660), .A2(n543), .ZN(n544) );
  NAND2_X1 U647 ( .A1(n544), .A2(n564), .ZN(n616) );
  INV_X1 U648 ( .A(n546), .ZN(n547) );
  NOR2_X1 U649 ( .A1(n548), .A2(n547), .ZN(n626) );
  NAND2_X1 U650 ( .A1(n548), .A2(n547), .ZN(n634) );
  INV_X1 U651 ( .A(n634), .ZN(n631) );
  NOR2_X1 U652 ( .A1(n626), .A2(n631), .ZN(n651) );
  NAND2_X1 U653 ( .A1(n664), .A2(n549), .ZN(n667) );
  NOR2_X1 U654 ( .A1(n664), .A2(n551), .ZN(n552) );
  NAND2_X1 U655 ( .A1(n581), .A2(n552), .ZN(n618) );
  NAND2_X1 U656 ( .A1(n555), .A2(n554), .ZN(n556) );
  NOR2_X1 U657 ( .A1(n561), .A2(n560), .ZN(n562) );
  XOR2_X1 U658 ( .A(KEYINPUT81), .B(n562), .Z(n582) );
  OR2_X1 U659 ( .A1(n572), .A2(n564), .ZN(n565) );
  NOR2_X1 U660 ( .A1(n634), .A2(n565), .ZN(n566) );
  NAND2_X1 U661 ( .A1(n566), .A2(n646), .ZN(n585) );
  NOR2_X1 U662 ( .A1(n567), .A2(n585), .ZN(n568) );
  XNOR2_X1 U663 ( .A(n568), .B(KEYINPUT43), .ZN(n569) );
  NOR2_X1 U664 ( .A1(n384), .A2(n569), .ZN(n644) );
  XNOR2_X1 U665 ( .A(n571), .B(KEYINPUT108), .ZN(n652) );
  XNOR2_X1 U666 ( .A(n574), .B(KEYINPUT28), .ZN(n577) );
  INV_X1 U667 ( .A(n575), .ZN(n576) );
  NOR2_X1 U668 ( .A1(n677), .A2(n578), .ZN(n579) );
  NAND2_X1 U669 ( .A1(n664), .A2(n646), .ZN(n580) );
  XOR2_X1 U670 ( .A(KEYINPUT30), .B(n580), .Z(n584) );
  XNOR2_X1 U671 ( .A(n581), .B(KEYINPUT107), .ZN(n583) );
  INV_X1 U672 ( .A(n570), .ZN(n592) );
  NOR2_X1 U673 ( .A1(n592), .A2(n585), .ZN(n586) );
  XOR2_X1 U674 ( .A(KEYINPUT36), .B(n586), .Z(n587) );
  NOR2_X1 U675 ( .A1(n657), .A2(n587), .ZN(n641) );
  NAND2_X1 U676 ( .A1(n651), .A2(KEYINPUT47), .ZN(n593) );
  OR2_X1 U677 ( .A1(n625), .A2(n651), .ZN(n595) );
  NOR2_X1 U678 ( .A1(KEYINPUT47), .A2(n595), .ZN(n596) );
  NAND2_X1 U679 ( .A1(n597), .A2(n626), .ZN(n643) );
  NAND2_X1 U680 ( .A1(n699), .A2(G472), .ZN(n605) );
  XOR2_X1 U681 ( .A(KEYINPUT109), .B(KEYINPUT62), .Z(n602) );
  XNOR2_X1 U682 ( .A(n605), .B(n604), .ZN(n606) );
  XNOR2_X1 U683 ( .A(n608), .B(n607), .ZN(G57) );
  NAND2_X1 U684 ( .A1(n699), .A2(G210), .ZN(n613) );
  XOR2_X1 U685 ( .A(KEYINPUT55), .B(KEYINPUT54), .Z(n610) );
  XNOR2_X1 U686 ( .A(KEYINPUT88), .B(KEYINPUT83), .ZN(n609) );
  XNOR2_X1 U687 ( .A(n610), .B(n609), .ZN(n611) );
  INV_X1 U688 ( .A(KEYINPUT56), .ZN(n614) );
  XNOR2_X1 U689 ( .A(n614), .B(KEYINPUT87), .ZN(n615) );
  XNOR2_X1 U690 ( .A(G101), .B(n616), .ZN(G3) );
  NOR2_X1 U691 ( .A1(n634), .A2(n618), .ZN(n617) );
  XOR2_X1 U692 ( .A(G104), .B(n617), .Z(G6) );
  INV_X1 U693 ( .A(n626), .ZN(n637) );
  NOR2_X1 U694 ( .A1(n637), .A2(n618), .ZN(n623) );
  XOR2_X1 U695 ( .A(KEYINPUT111), .B(KEYINPUT27), .Z(n620) );
  XNOR2_X1 U696 ( .A(G107), .B(KEYINPUT26), .ZN(n619) );
  XNOR2_X1 U697 ( .A(n620), .B(n619), .ZN(n621) );
  XNOR2_X1 U698 ( .A(KEYINPUT110), .B(n621), .ZN(n622) );
  XNOR2_X1 U699 ( .A(n623), .B(n622), .ZN(G9) );
  XOR2_X1 U700 ( .A(n624), .B(G110), .Z(G12) );
  XOR2_X1 U701 ( .A(KEYINPUT112), .B(KEYINPUT29), .Z(n628) );
  NAND2_X1 U702 ( .A1(n626), .A2(n632), .ZN(n627) );
  XNOR2_X1 U703 ( .A(n628), .B(n627), .ZN(n629) );
  XNOR2_X1 U704 ( .A(G128), .B(n629), .ZN(G30) );
  XNOR2_X1 U705 ( .A(n630), .B(KEYINPUT113), .ZN(G45) );
  NAND2_X1 U706 ( .A1(n632), .A2(n631), .ZN(n633) );
  XNOR2_X1 U707 ( .A(n633), .B(G146), .ZN(G48) );
  NOR2_X1 U708 ( .A1(n634), .A2(n636), .ZN(n635) );
  XOR2_X1 U709 ( .A(G113), .B(n635), .Z(G15) );
  NOR2_X1 U710 ( .A1(n637), .A2(n636), .ZN(n639) );
  XNOR2_X1 U711 ( .A(KEYINPUT114), .B(KEYINPUT115), .ZN(n638) );
  XNOR2_X1 U712 ( .A(n639), .B(n638), .ZN(n640) );
  XNOR2_X1 U713 ( .A(G116), .B(n640), .ZN(G18) );
  XNOR2_X1 U714 ( .A(G125), .B(n641), .ZN(n642) );
  XNOR2_X1 U715 ( .A(n642), .B(KEYINPUT37), .ZN(G27) );
  XNOR2_X1 U716 ( .A(G134), .B(n643), .ZN(G36) );
  XOR2_X1 U717 ( .A(G140), .B(n644), .Z(n645) );
  XNOR2_X1 U718 ( .A(KEYINPUT116), .B(n645), .ZN(G42) );
  NOR2_X1 U719 ( .A1(n647), .A2(n646), .ZN(n648) );
  XOR2_X1 U720 ( .A(KEYINPUT117), .B(n648), .Z(n649) );
  NOR2_X1 U721 ( .A1(n650), .A2(n649), .ZN(n655) );
  NOR2_X1 U722 ( .A1(n652), .A2(n651), .ZN(n653) );
  XNOR2_X1 U723 ( .A(n653), .B(KEYINPUT118), .ZN(n654) );
  NOR2_X1 U724 ( .A1(n655), .A2(n654), .ZN(n656) );
  NOR2_X1 U725 ( .A1(n656), .A2(n678), .ZN(n672) );
  NAND2_X1 U726 ( .A1(n658), .A2(n657), .ZN(n659) );
  XNOR2_X1 U727 ( .A(n659), .B(KEYINPUT50), .ZN(n666) );
  NOR2_X1 U728 ( .A1(n661), .A2(n660), .ZN(n662) );
  XOR2_X1 U729 ( .A(KEYINPUT49), .B(n662), .Z(n663) );
  NOR2_X1 U730 ( .A1(n664), .A2(n663), .ZN(n665) );
  NAND2_X1 U731 ( .A1(n666), .A2(n665), .ZN(n668) );
  NAND2_X1 U732 ( .A1(n668), .A2(n667), .ZN(n669) );
  XNOR2_X1 U733 ( .A(KEYINPUT51), .B(n669), .ZN(n670) );
  NOR2_X1 U734 ( .A1(n670), .A2(n677), .ZN(n671) );
  NOR2_X1 U735 ( .A1(n672), .A2(n671), .ZN(n673) );
  XOR2_X1 U736 ( .A(n673), .B(KEYINPUT119), .Z(n674) );
  XNOR2_X1 U737 ( .A(KEYINPUT52), .B(n674), .ZN(n675) );
  NOR2_X1 U738 ( .A1(n676), .A2(n675), .ZN(n680) );
  NOR2_X1 U739 ( .A1(n678), .A2(n677), .ZN(n679) );
  NOR2_X1 U740 ( .A1(n680), .A2(n679), .ZN(n685) );
  XOR2_X1 U741 ( .A(n681), .B(KEYINPUT82), .Z(n683) );
  NAND2_X1 U742 ( .A1(n683), .A2(n682), .ZN(n684) );
  NAND2_X1 U743 ( .A1(n685), .A2(n684), .ZN(n686) );
  NOR2_X1 U744 ( .A1(G953), .A2(n686), .ZN(n688) );
  XNOR2_X1 U745 ( .A(KEYINPUT53), .B(KEYINPUT120), .ZN(n687) );
  XNOR2_X1 U746 ( .A(n688), .B(n687), .ZN(G75) );
  XOR2_X1 U747 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n691) );
  XNOR2_X1 U748 ( .A(n689), .B(KEYINPUT121), .ZN(n690) );
  XNOR2_X1 U749 ( .A(n691), .B(n690), .ZN(n693) );
  NAND2_X1 U750 ( .A1(n699), .A2(G469), .ZN(n692) );
  XOR2_X1 U751 ( .A(n693), .B(n692), .Z(n694) );
  NOR2_X1 U752 ( .A1(n701), .A2(n694), .ZN(G54) );
  NAND2_X1 U753 ( .A1(n699), .A2(G478), .ZN(n696) );
  NOR2_X1 U754 ( .A1(n701), .A2(n698), .ZN(G63) );
  NAND2_X1 U755 ( .A1(G953), .A2(G224), .ZN(n702) );
  XOR2_X1 U756 ( .A(KEYINPUT61), .B(n702), .Z(n703) );
  NOR2_X1 U757 ( .A1(n704), .A2(n703), .ZN(n705) );
  XNOR2_X1 U758 ( .A(n705), .B(KEYINPUT124), .ZN(n708) );
  NOR2_X1 U759 ( .A1(n706), .A2(G953), .ZN(n707) );
  NOR2_X1 U760 ( .A1(n708), .A2(n707), .ZN(n709) );
  XOR2_X1 U761 ( .A(n709), .B(KEYINPUT125), .Z(n714) );
  XOR2_X1 U762 ( .A(n710), .B(G101), .Z(n712) );
  NAND2_X1 U763 ( .A1(n712), .A2(n711), .ZN(n713) );
  XNOR2_X1 U764 ( .A(n714), .B(n713), .ZN(G69) );
  XOR2_X1 U765 ( .A(n716), .B(n715), .Z(n717) );
  XNOR2_X1 U766 ( .A(KEYINPUT126), .B(n717), .ZN(n718) );
  XNOR2_X1 U767 ( .A(n719), .B(n718), .ZN(n723) );
  XNOR2_X1 U768 ( .A(n723), .B(n720), .ZN(n722) );
  NAND2_X1 U769 ( .A1(n722), .A2(n721), .ZN(n728) );
  XNOR2_X1 U770 ( .A(G227), .B(n723), .ZN(n724) );
  NAND2_X1 U771 ( .A1(n724), .A2(G900), .ZN(n725) );
  XOR2_X1 U772 ( .A(KEYINPUT127), .B(n725), .Z(n726) );
  NAND2_X1 U773 ( .A1(G953), .A2(n726), .ZN(n727) );
  NAND2_X1 U774 ( .A1(n728), .A2(n727), .ZN(G72) );
  XNOR2_X1 U775 ( .A(n729), .B(G119), .ZN(G21) );
  XOR2_X1 U776 ( .A(n730), .B(G122), .Z(G24) );
  XOR2_X1 U777 ( .A(n731), .B(G131), .Z(G33) );
  XOR2_X1 U778 ( .A(n732), .B(G137), .Z(G39) );
endmodule

