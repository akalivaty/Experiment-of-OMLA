//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 1 1 0 0 1 1 1 1 1 0 0 1 0 0 1 0 1 0 0 0 1 0 0 0 0 1 1 0 1 1 1 0 0 1 1 0 1 0 1 1 1 1 1 0 1 0 0 0 1 1 1 1 0 1 1 0 1 1 1 0 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:27:52 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n697, new_n698, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n713, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n723, new_n724, new_n725, new_n726, new_n727, new_n728,
    new_n729, new_n730, new_n731, new_n732, new_n733, new_n734, new_n735,
    new_n736, new_n737, new_n738, new_n739, new_n740, new_n741, new_n743,
    new_n744, new_n745, new_n746, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n764, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n790, new_n791, new_n792, new_n793, new_n794, new_n795, new_n796,
    new_n797, new_n798, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n904, new_n905, new_n906, new_n907, new_n908, new_n909, new_n910,
    new_n911, new_n912, new_n913, new_n914, new_n915, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n930, new_n931, new_n932, new_n933, new_n934,
    new_n935, new_n936, new_n937, new_n938, new_n939, new_n940, new_n941,
    new_n942, new_n943, new_n945, new_n946, new_n947, new_n948, new_n949,
    new_n950, new_n951, new_n952, new_n953, new_n954, new_n955, new_n956,
    new_n957, new_n959, new_n960, new_n961, new_n962, new_n963, new_n964,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n988, new_n989, new_n990, new_n991, new_n992, new_n993, new_n994,
    new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002;
  OR2_X1    g000(.A1(KEYINPUT64), .A2(G143), .ZN(new_n187));
  INV_X1    g001(.A(G146), .ZN(new_n188));
  NAND2_X1  g002(.A1(KEYINPUT64), .A2(G143), .ZN(new_n189));
  NAND3_X1  g003(.A1(new_n187), .A2(new_n188), .A3(new_n189), .ZN(new_n190));
  INV_X1    g004(.A(KEYINPUT65), .ZN(new_n191));
  INV_X1    g005(.A(G143), .ZN(new_n192));
  AOI21_X1  g006(.A(new_n191), .B1(new_n192), .B2(G146), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n190), .A2(new_n193), .ZN(new_n194));
  INV_X1    g008(.A(KEYINPUT0), .ZN(new_n195));
  INV_X1    g009(.A(G128), .ZN(new_n196));
  NOR2_X1   g010(.A1(new_n195), .A2(new_n196), .ZN(new_n197));
  INV_X1    g011(.A(new_n197), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n195), .A2(new_n196), .ZN(new_n199));
  NAND4_X1  g013(.A1(new_n187), .A2(new_n191), .A3(new_n188), .A4(new_n189), .ZN(new_n200));
  NAND4_X1  g014(.A1(new_n194), .A2(new_n198), .A3(new_n199), .A4(new_n200), .ZN(new_n201));
  NAND2_X1  g015(.A1(KEYINPUT75), .A2(G125), .ZN(new_n202));
  INV_X1    g016(.A(new_n202), .ZN(new_n203));
  NOR2_X1   g017(.A1(KEYINPUT75), .A2(G125), .ZN(new_n204));
  NOR2_X1   g018(.A1(new_n203), .A2(new_n204), .ZN(new_n205));
  INV_X1    g019(.A(KEYINPUT67), .ZN(new_n206));
  XNOR2_X1  g020(.A(KEYINPUT64), .B(G143), .ZN(new_n207));
  OAI21_X1  g021(.A(KEYINPUT66), .B1(new_n192), .B2(G146), .ZN(new_n208));
  INV_X1    g022(.A(KEYINPUT66), .ZN(new_n209));
  NAND3_X1  g023(.A1(new_n209), .A2(new_n188), .A3(G143), .ZN(new_n210));
  AOI22_X1  g024(.A1(new_n207), .A2(G146), .B1(new_n208), .B2(new_n210), .ZN(new_n211));
  AOI21_X1  g025(.A(new_n206), .B1(new_n211), .B2(new_n197), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n208), .A2(new_n210), .ZN(new_n213));
  AND2_X1   g027(.A1(KEYINPUT64), .A2(G143), .ZN(new_n214));
  NOR2_X1   g028(.A1(KEYINPUT64), .A2(G143), .ZN(new_n215));
  OAI21_X1  g029(.A(G146), .B1(new_n214), .B2(new_n215), .ZN(new_n216));
  NAND4_X1  g030(.A1(new_n213), .A2(new_n216), .A3(new_n206), .A4(new_n197), .ZN(new_n217));
  INV_X1    g031(.A(new_n217), .ZN(new_n218));
  OAI211_X1 g032(.A(new_n201), .B(new_n205), .C1(new_n212), .C2(new_n218), .ZN(new_n219));
  OAI21_X1  g033(.A(KEYINPUT1), .B1(new_n192), .B2(G146), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n220), .A2(G128), .ZN(new_n221));
  NOR3_X1   g035(.A1(new_n214), .A2(new_n215), .A3(G146), .ZN(new_n222));
  INV_X1    g036(.A(new_n193), .ZN(new_n223));
  OAI211_X1 g037(.A(new_n200), .B(new_n221), .C1(new_n222), .C2(new_n223), .ZN(new_n224));
  INV_X1    g038(.A(KEYINPUT1), .ZN(new_n225));
  NAND4_X1  g039(.A1(new_n213), .A2(new_n216), .A3(new_n225), .A4(G128), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n224), .A2(new_n226), .ZN(new_n227));
  OAI21_X1  g041(.A(new_n227), .B1(new_n204), .B2(new_n203), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n219), .A2(new_n228), .ZN(new_n229));
  INV_X1    g043(.A(G224), .ZN(new_n230));
  NOR2_X1   g044(.A1(new_n230), .A2(G953), .ZN(new_n231));
  INV_X1    g045(.A(new_n231), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n229), .A2(new_n232), .ZN(new_n233));
  NAND3_X1  g047(.A1(new_n219), .A2(new_n228), .A3(new_n231), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n233), .A2(new_n234), .ZN(new_n235));
  XNOR2_X1  g049(.A(KEYINPUT2), .B(G113), .ZN(new_n236));
  INV_X1    g050(.A(G119), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n237), .A2(G116), .ZN(new_n238));
  INV_X1    g052(.A(G116), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n239), .A2(G119), .ZN(new_n240));
  AND3_X1   g054(.A1(new_n238), .A2(new_n240), .A3(KEYINPUT69), .ZN(new_n241));
  AOI21_X1  g055(.A(KEYINPUT69), .B1(new_n238), .B2(new_n240), .ZN(new_n242));
  OAI21_X1  g056(.A(new_n236), .B1(new_n241), .B2(new_n242), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n238), .A2(new_n240), .ZN(new_n244));
  OR2_X1    g058(.A1(new_n244), .A2(new_n236), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n243), .A2(new_n245), .ZN(new_n246));
  INV_X1    g060(.A(G104), .ZN(new_n247));
  OAI21_X1  g061(.A(KEYINPUT3), .B1(new_n247), .B2(G107), .ZN(new_n248));
  INV_X1    g062(.A(KEYINPUT3), .ZN(new_n249));
  INV_X1    g063(.A(G107), .ZN(new_n250));
  NAND3_X1  g064(.A1(new_n249), .A2(new_n250), .A3(G104), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n247), .A2(G107), .ZN(new_n252));
  NAND3_X1  g066(.A1(new_n248), .A2(new_n251), .A3(new_n252), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n253), .A2(G101), .ZN(new_n254));
  XNOR2_X1  g068(.A(KEYINPUT78), .B(G101), .ZN(new_n255));
  NAND4_X1  g069(.A1(new_n255), .A2(new_n252), .A3(new_n248), .A4(new_n251), .ZN(new_n256));
  NAND3_X1  g070(.A1(new_n254), .A2(KEYINPUT4), .A3(new_n256), .ZN(new_n257));
  INV_X1    g071(.A(KEYINPUT4), .ZN(new_n258));
  NAND3_X1  g072(.A1(new_n253), .A2(new_n258), .A3(G101), .ZN(new_n259));
  NAND3_X1  g073(.A1(new_n246), .A2(new_n257), .A3(new_n259), .ZN(new_n260));
  INV_X1    g074(.A(KEYINPUT69), .ZN(new_n261));
  NOR2_X1   g075(.A1(new_n239), .A2(G119), .ZN(new_n262));
  NOR2_X1   g076(.A1(new_n237), .A2(G116), .ZN(new_n263));
  OAI21_X1  g077(.A(new_n261), .B1(new_n262), .B2(new_n263), .ZN(new_n264));
  NAND3_X1  g078(.A1(new_n238), .A2(new_n240), .A3(KEYINPUT69), .ZN(new_n265));
  NAND3_X1  g079(.A1(new_n264), .A2(KEYINPUT5), .A3(new_n265), .ZN(new_n266));
  INV_X1    g080(.A(G113), .ZN(new_n267));
  INV_X1    g081(.A(KEYINPUT5), .ZN(new_n268));
  AOI21_X1  g082(.A(new_n267), .B1(new_n262), .B2(new_n268), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n266), .A2(new_n269), .ZN(new_n270));
  AND3_X1   g084(.A1(new_n248), .A2(new_n251), .A3(new_n252), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n250), .A2(G104), .ZN(new_n272));
  NAND2_X1  g086(.A1(new_n252), .A2(new_n272), .ZN(new_n273));
  AOI22_X1  g087(.A1(new_n271), .A2(new_n255), .B1(G101), .B2(new_n273), .ZN(new_n274));
  NAND3_X1  g088(.A1(new_n270), .A2(new_n245), .A3(new_n274), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n260), .A2(new_n275), .ZN(new_n276));
  XNOR2_X1  g090(.A(G110), .B(G122), .ZN(new_n277));
  INV_X1    g091(.A(new_n277), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n276), .A2(new_n278), .ZN(new_n279));
  NAND3_X1  g093(.A1(new_n260), .A2(new_n275), .A3(new_n277), .ZN(new_n280));
  NAND3_X1  g094(.A1(new_n279), .A2(KEYINPUT6), .A3(new_n280), .ZN(new_n281));
  INV_X1    g095(.A(KEYINPUT80), .ZN(new_n282));
  INV_X1    g096(.A(KEYINPUT6), .ZN(new_n283));
  AND4_X1   g097(.A1(new_n282), .A2(new_n276), .A3(new_n283), .A4(new_n278), .ZN(new_n284));
  AOI21_X1  g098(.A(new_n277), .B1(new_n260), .B2(new_n275), .ZN(new_n285));
  AOI21_X1  g099(.A(new_n282), .B1(new_n285), .B2(new_n283), .ZN(new_n286));
  OAI211_X1 g100(.A(new_n235), .B(new_n281), .C1(new_n284), .C2(new_n286), .ZN(new_n287));
  INV_X1    g101(.A(G902), .ZN(new_n288));
  INV_X1    g102(.A(KEYINPUT7), .ZN(new_n289));
  NAND3_X1  g103(.A1(new_n219), .A2(new_n228), .A3(new_n289), .ZN(new_n290));
  AND2_X1   g104(.A1(new_n290), .A2(new_n280), .ZN(new_n291));
  NAND3_X1  g105(.A1(new_n229), .A2(KEYINPUT7), .A3(new_n232), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n273), .A2(G101), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n256), .A2(new_n293), .ZN(new_n294));
  NAND3_X1  g108(.A1(new_n270), .A2(new_n245), .A3(new_n294), .ZN(new_n295));
  XNOR2_X1  g109(.A(new_n277), .B(KEYINPUT8), .ZN(new_n296));
  OAI21_X1  g110(.A(new_n269), .B1(new_n268), .B2(new_n244), .ZN(new_n297));
  AND2_X1   g111(.A1(new_n297), .A2(new_n245), .ZN(new_n298));
  OAI211_X1 g112(.A(new_n295), .B(new_n296), .C1(new_n294), .C2(new_n298), .ZN(new_n299));
  NAND4_X1  g113(.A1(new_n291), .A2(new_n292), .A3(new_n299), .A4(new_n234), .ZN(new_n300));
  NAND3_X1  g114(.A1(new_n287), .A2(new_n288), .A3(new_n300), .ZN(new_n301));
  OAI21_X1  g115(.A(G210), .B1(G237), .B2(G902), .ZN(new_n302));
  XNOR2_X1  g116(.A(new_n302), .B(KEYINPUT81), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n301), .A2(new_n303), .ZN(new_n304));
  NAND4_X1  g118(.A1(new_n287), .A2(new_n288), .A3(new_n300), .A4(new_n302), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n304), .A2(new_n305), .ZN(new_n306));
  OAI21_X1  g120(.A(G214), .B1(G237), .B2(G902), .ZN(new_n307));
  INV_X1    g121(.A(G953), .ZN(new_n308));
  AND2_X1   g122(.A1(new_n308), .A2(G952), .ZN(new_n309));
  NAND2_X1  g123(.A1(G234), .A2(G237), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n309), .A2(new_n310), .ZN(new_n311));
  INV_X1    g125(.A(new_n311), .ZN(new_n312));
  XOR2_X1   g126(.A(KEYINPUT21), .B(G898), .Z(new_n313));
  INV_X1    g127(.A(new_n313), .ZN(new_n314));
  NAND3_X1  g128(.A1(new_n310), .A2(G902), .A3(G953), .ZN(new_n315));
  INV_X1    g129(.A(new_n315), .ZN(new_n316));
  AOI21_X1  g130(.A(new_n312), .B1(new_n314), .B2(new_n316), .ZN(new_n317));
  INV_X1    g131(.A(new_n317), .ZN(new_n318));
  NAND3_X1  g132(.A1(new_n306), .A2(new_n307), .A3(new_n318), .ZN(new_n319));
  INV_X1    g133(.A(G469), .ZN(new_n320));
  AOI21_X1  g134(.A(new_n196), .B1(new_n190), .B2(KEYINPUT1), .ZN(new_n321));
  OAI21_X1  g135(.A(new_n226), .B1(new_n321), .B2(new_n211), .ZN(new_n322));
  AOI21_X1  g136(.A(KEYINPUT10), .B1(new_n322), .B2(new_n274), .ZN(new_n323));
  INV_X1    g137(.A(new_n323), .ZN(new_n324));
  NAND3_X1  g138(.A1(new_n213), .A2(new_n216), .A3(new_n197), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n325), .A2(KEYINPUT67), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n326), .A2(new_n217), .ZN(new_n327));
  NAND4_X1  g141(.A1(new_n327), .A2(new_n201), .A3(new_n257), .A4(new_n259), .ZN(new_n328));
  INV_X1    g142(.A(KEYINPUT11), .ZN(new_n329));
  INV_X1    g143(.A(G134), .ZN(new_n330));
  OAI21_X1  g144(.A(new_n329), .B1(new_n330), .B2(G137), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n330), .A2(G137), .ZN(new_n332));
  INV_X1    g146(.A(G137), .ZN(new_n333));
  NAND3_X1  g147(.A1(new_n333), .A2(KEYINPUT11), .A3(G134), .ZN(new_n334));
  NAND3_X1  g148(.A1(new_n331), .A2(new_n332), .A3(new_n334), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n335), .A2(G131), .ZN(new_n336));
  INV_X1    g150(.A(G131), .ZN(new_n337));
  NAND4_X1  g151(.A1(new_n331), .A2(new_n334), .A3(new_n337), .A4(new_n332), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n336), .A2(new_n338), .ZN(new_n339));
  INV_X1    g153(.A(new_n339), .ZN(new_n340));
  NAND3_X1  g154(.A1(new_n227), .A2(KEYINPUT10), .A3(new_n274), .ZN(new_n341));
  NAND4_X1  g155(.A1(new_n324), .A2(new_n328), .A3(new_n340), .A4(new_n341), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n322), .A2(new_n274), .ZN(new_n343));
  NAND3_X1  g157(.A1(new_n294), .A2(new_n224), .A3(new_n226), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n343), .A2(new_n344), .ZN(new_n345));
  AOI21_X1  g159(.A(KEYINPUT12), .B1(new_n345), .B2(new_n339), .ZN(new_n346));
  INV_X1    g160(.A(KEYINPUT12), .ZN(new_n347));
  AOI211_X1 g161(.A(new_n347), .B(new_n340), .C1(new_n343), .C2(new_n344), .ZN(new_n348));
  OAI21_X1  g162(.A(new_n342), .B1(new_n346), .B2(new_n348), .ZN(new_n349));
  XNOR2_X1  g163(.A(G110), .B(G140), .ZN(new_n350));
  INV_X1    g164(.A(G227), .ZN(new_n351));
  NOR2_X1   g165(.A1(new_n351), .A2(G953), .ZN(new_n352));
  XOR2_X1   g166(.A(new_n350), .B(new_n352), .Z(new_n353));
  INV_X1    g167(.A(new_n353), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n349), .A2(new_n354), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n328), .A2(new_n341), .ZN(new_n356));
  OAI21_X1  g170(.A(new_n339), .B1(new_n356), .B2(new_n323), .ZN(new_n357));
  NAND3_X1  g171(.A1(new_n357), .A2(new_n342), .A3(new_n353), .ZN(new_n358));
  NAND2_X1  g172(.A1(new_n355), .A2(new_n358), .ZN(new_n359));
  AOI21_X1  g173(.A(new_n320), .B1(new_n359), .B2(new_n288), .ZN(new_n360));
  OAI211_X1 g174(.A(new_n342), .B(new_n353), .C1(new_n346), .C2(new_n348), .ZN(new_n361));
  INV_X1    g175(.A(new_n361), .ZN(new_n362));
  AOI21_X1  g176(.A(new_n353), .B1(new_n357), .B2(new_n342), .ZN(new_n363));
  OAI211_X1 g177(.A(new_n320), .B(new_n288), .C1(new_n362), .C2(new_n363), .ZN(new_n364));
  INV_X1    g178(.A(KEYINPUT79), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n364), .A2(new_n365), .ZN(new_n366));
  AND3_X1   g180(.A1(new_n194), .A2(new_n198), .A3(new_n200), .ZN(new_n367));
  AOI22_X1  g181(.A1(new_n367), .A2(new_n199), .B1(new_n326), .B2(new_n217), .ZN(new_n368));
  AND2_X1   g182(.A1(new_n257), .A2(new_n259), .ZN(new_n369));
  AOI21_X1  g183(.A(new_n294), .B1(new_n224), .B2(new_n226), .ZN(new_n370));
  AOI22_X1  g184(.A1(new_n368), .A2(new_n369), .B1(KEYINPUT10), .B2(new_n370), .ZN(new_n371));
  AOI21_X1  g185(.A(new_n340), .B1(new_n371), .B2(new_n324), .ZN(new_n372));
  INV_X1    g186(.A(new_n342), .ZN(new_n373));
  OAI21_X1  g187(.A(new_n354), .B1(new_n372), .B2(new_n373), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n374), .A2(new_n361), .ZN(new_n375));
  NAND4_X1  g189(.A1(new_n375), .A2(KEYINPUT79), .A3(new_n320), .A4(new_n288), .ZN(new_n376));
  AOI21_X1  g190(.A(new_n360), .B1(new_n366), .B2(new_n376), .ZN(new_n377));
  INV_X1    g191(.A(G221), .ZN(new_n378));
  XOR2_X1   g192(.A(KEYINPUT9), .B(G234), .Z(new_n379));
  AOI21_X1  g193(.A(new_n378), .B1(new_n379), .B2(new_n288), .ZN(new_n380));
  NOR3_X1   g194(.A1(new_n319), .A2(new_n377), .A3(new_n380), .ZN(new_n381));
  INV_X1    g195(.A(KEYINPUT87), .ZN(new_n382));
  OAI21_X1  g196(.A(new_n382), .B1(new_n192), .B2(G128), .ZN(new_n383));
  NAND3_X1  g197(.A1(new_n196), .A2(KEYINPUT87), .A3(G143), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n383), .A2(new_n384), .ZN(new_n385));
  OAI21_X1  g199(.A(G128), .B1(new_n214), .B2(new_n215), .ZN(new_n386));
  NAND2_X1  g200(.A1(new_n385), .A2(new_n386), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n387), .A2(G134), .ZN(new_n388));
  NAND3_X1  g202(.A1(new_n385), .A2(new_n386), .A3(new_n330), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n388), .A2(new_n389), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n390), .A2(KEYINPUT90), .ZN(new_n391));
  INV_X1    g205(.A(KEYINPUT14), .ZN(new_n392));
  NAND3_X1  g206(.A1(new_n392), .A2(new_n239), .A3(G122), .ZN(new_n393));
  INV_X1    g207(.A(KEYINPUT91), .ZN(new_n394));
  OR2_X1    g208(.A1(new_n393), .A2(new_n394), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n393), .A2(new_n394), .ZN(new_n396));
  OAI211_X1 g210(.A(new_n395), .B(new_n396), .C1(new_n239), .C2(G122), .ZN(new_n397));
  AOI21_X1  g211(.A(new_n392), .B1(new_n239), .B2(G122), .ZN(new_n398));
  OAI21_X1  g212(.A(G107), .B1(new_n397), .B2(new_n398), .ZN(new_n399));
  XNOR2_X1  g213(.A(G116), .B(G122), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n400), .A2(new_n250), .ZN(new_n401));
  INV_X1    g215(.A(KEYINPUT90), .ZN(new_n402));
  NAND3_X1  g216(.A1(new_n388), .A2(new_n402), .A3(new_n389), .ZN(new_n403));
  NAND4_X1  g217(.A1(new_n391), .A2(new_n399), .A3(new_n401), .A4(new_n403), .ZN(new_n404));
  AOI21_X1  g218(.A(new_n196), .B1(new_n187), .B2(new_n189), .ZN(new_n405));
  XNOR2_X1  g219(.A(KEYINPUT86), .B(KEYINPUT13), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n405), .A2(new_n406), .ZN(new_n407));
  XOR2_X1   g221(.A(KEYINPUT86), .B(KEYINPUT13), .Z(new_n408));
  NAND2_X1  g222(.A1(new_n408), .A2(new_n386), .ZN(new_n409));
  NAND3_X1  g223(.A1(new_n407), .A2(new_n409), .A3(new_n385), .ZN(new_n410));
  INV_X1    g224(.A(KEYINPUT88), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n389), .A2(new_n411), .ZN(new_n412));
  NAND4_X1  g226(.A1(new_n385), .A2(new_n386), .A3(KEYINPUT88), .A4(new_n330), .ZN(new_n413));
  AOI22_X1  g227(.A1(G134), .A2(new_n410), .B1(new_n412), .B2(new_n413), .ZN(new_n414));
  XNOR2_X1  g228(.A(new_n400), .B(new_n250), .ZN(new_n415));
  AOI21_X1  g229(.A(KEYINPUT89), .B1(new_n414), .B2(new_n415), .ZN(new_n416));
  NAND2_X1  g230(.A1(new_n412), .A2(new_n413), .ZN(new_n417));
  OAI21_X1  g231(.A(new_n385), .B1(new_n405), .B2(new_n406), .ZN(new_n418));
  NOR2_X1   g232(.A1(new_n408), .A2(new_n386), .ZN(new_n419));
  OAI21_X1  g233(.A(G134), .B1(new_n418), .B2(new_n419), .ZN(new_n420));
  AND4_X1   g234(.A1(KEYINPUT89), .A2(new_n417), .A3(new_n415), .A4(new_n420), .ZN(new_n421));
  OAI21_X1  g235(.A(new_n404), .B1(new_n416), .B2(new_n421), .ZN(new_n422));
  NAND3_X1  g236(.A1(new_n379), .A2(G217), .A3(new_n308), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n422), .A2(new_n423), .ZN(new_n424));
  INV_X1    g238(.A(new_n423), .ZN(new_n425));
  OAI211_X1 g239(.A(new_n404), .B(new_n425), .C1(new_n416), .C2(new_n421), .ZN(new_n426));
  NAND3_X1  g240(.A1(new_n424), .A2(KEYINPUT92), .A3(new_n426), .ZN(new_n427));
  INV_X1    g241(.A(new_n422), .ZN(new_n428));
  INV_X1    g242(.A(KEYINPUT92), .ZN(new_n429));
  NAND3_X1  g243(.A1(new_n428), .A2(new_n429), .A3(new_n425), .ZN(new_n430));
  NAND3_X1  g244(.A1(new_n427), .A2(new_n288), .A3(new_n430), .ZN(new_n431));
  INV_X1    g245(.A(KEYINPUT93), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n431), .A2(new_n432), .ZN(new_n433));
  NAND4_X1  g247(.A1(new_n427), .A2(new_n430), .A3(KEYINPUT93), .A4(new_n288), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n433), .A2(new_n434), .ZN(new_n435));
  INV_X1    g249(.A(G478), .ZN(new_n436));
  NOR2_X1   g250(.A1(new_n436), .A2(KEYINPUT15), .ZN(new_n437));
  NAND2_X1  g251(.A1(new_n435), .A2(new_n437), .ZN(new_n438));
  INV_X1    g252(.A(KEYINPUT94), .ZN(new_n439));
  NOR2_X1   g253(.A1(new_n431), .A2(new_n437), .ZN(new_n440));
  INV_X1    g254(.A(new_n440), .ZN(new_n441));
  NAND3_X1  g255(.A1(new_n438), .A2(new_n439), .A3(new_n441), .ZN(new_n442));
  INV_X1    g256(.A(G214), .ZN(new_n443));
  NOR3_X1   g257(.A1(new_n443), .A2(G237), .A3(G953), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n444), .A2(new_n192), .ZN(new_n445));
  OAI21_X1  g259(.A(new_n445), .B1(new_n207), .B2(new_n444), .ZN(new_n446));
  INV_X1    g260(.A(KEYINPUT18), .ZN(new_n447));
  NOR3_X1   g261(.A1(new_n446), .A2(new_n447), .A3(new_n337), .ZN(new_n448));
  INV_X1    g262(.A(KEYINPUT82), .ZN(new_n449));
  XNOR2_X1  g263(.A(new_n448), .B(new_n449), .ZN(new_n450));
  AND2_X1   g264(.A1(G125), .A2(G140), .ZN(new_n451));
  NOR2_X1   g265(.A1(G125), .A2(G140), .ZN(new_n452));
  NOR2_X1   g266(.A1(new_n451), .A2(new_n452), .ZN(new_n453));
  NOR2_X1   g267(.A1(new_n453), .A2(G146), .ZN(new_n454));
  XNOR2_X1  g268(.A(new_n454), .B(KEYINPUT76), .ZN(new_n455));
  INV_X1    g269(.A(G140), .ZN(new_n456));
  NOR3_X1   g270(.A1(new_n203), .A2(new_n204), .A3(new_n456), .ZN(new_n457));
  NOR2_X1   g271(.A1(new_n457), .A2(new_n452), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n458), .A2(G146), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n455), .A2(new_n459), .ZN(new_n460));
  OAI21_X1  g274(.A(new_n446), .B1(new_n447), .B2(new_n337), .ZN(new_n461));
  INV_X1    g275(.A(KEYINPUT83), .ZN(new_n462));
  XNOR2_X1  g276(.A(new_n461), .B(new_n462), .ZN(new_n463));
  NAND3_X1  g277(.A1(new_n450), .A2(new_n460), .A3(new_n463), .ZN(new_n464));
  XNOR2_X1  g278(.A(G113), .B(G122), .ZN(new_n465));
  XNOR2_X1  g279(.A(new_n465), .B(new_n247), .ZN(new_n466));
  OAI21_X1  g280(.A(KEYINPUT16), .B1(new_n457), .B2(new_n452), .ZN(new_n467));
  NOR4_X1   g281(.A1(new_n203), .A2(new_n204), .A3(KEYINPUT16), .A4(G140), .ZN(new_n468));
  INV_X1    g282(.A(new_n468), .ZN(new_n469));
  AOI21_X1  g283(.A(G146), .B1(new_n467), .B2(new_n469), .ZN(new_n470));
  INV_X1    g284(.A(KEYINPUT16), .ZN(new_n471));
  OR2_X1    g285(.A1(KEYINPUT75), .A2(G125), .ZN(new_n472));
  NAND3_X1  g286(.A1(new_n472), .A2(G140), .A3(new_n202), .ZN(new_n473));
  INV_X1    g287(.A(new_n452), .ZN(new_n474));
  AOI21_X1  g288(.A(new_n471), .B1(new_n473), .B2(new_n474), .ZN(new_n475));
  NOR3_X1   g289(.A1(new_n475), .A2(new_n188), .A3(new_n468), .ZN(new_n476));
  NOR2_X1   g290(.A1(new_n470), .A2(new_n476), .ZN(new_n477));
  NOR2_X1   g291(.A1(new_n446), .A2(new_n337), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n478), .A2(KEYINPUT17), .ZN(new_n479));
  XNOR2_X1  g293(.A(new_n446), .B(new_n337), .ZN(new_n480));
  OAI211_X1 g294(.A(new_n477), .B(new_n479), .C1(KEYINPUT17), .C2(new_n480), .ZN(new_n481));
  NAND3_X1  g295(.A1(new_n464), .A2(new_n466), .A3(new_n481), .ZN(new_n482));
  INV_X1    g296(.A(new_n482), .ZN(new_n483));
  AOI21_X1  g297(.A(new_n466), .B1(new_n464), .B2(new_n481), .ZN(new_n484));
  OAI21_X1  g298(.A(new_n288), .B1(new_n483), .B2(new_n484), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n485), .A2(G475), .ZN(new_n486));
  NAND3_X1  g300(.A1(new_n467), .A2(G146), .A3(new_n469), .ZN(new_n487));
  NAND2_X1  g301(.A1(new_n458), .A2(KEYINPUT19), .ZN(new_n488));
  NOR2_X1   g302(.A1(new_n453), .A2(KEYINPUT19), .ZN(new_n489));
  OAI21_X1  g303(.A(new_n488), .B1(KEYINPUT84), .B2(new_n489), .ZN(new_n490));
  OAI21_X1  g304(.A(new_n490), .B1(KEYINPUT84), .B2(new_n488), .ZN(new_n491));
  OAI211_X1 g305(.A(new_n487), .B(new_n480), .C1(new_n491), .C2(G146), .ZN(new_n492));
  AND2_X1   g306(.A1(new_n464), .A2(new_n492), .ZN(new_n493));
  OAI21_X1  g307(.A(new_n482), .B1(new_n493), .B2(new_n466), .ZN(new_n494));
  INV_X1    g308(.A(KEYINPUT20), .ZN(new_n495));
  INV_X1    g309(.A(G475), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n496), .A2(new_n288), .ZN(new_n497));
  XNOR2_X1  g311(.A(new_n497), .B(KEYINPUT85), .ZN(new_n498));
  NAND3_X1  g312(.A1(new_n494), .A2(new_n495), .A3(new_n498), .ZN(new_n499));
  INV_X1    g313(.A(new_n499), .ZN(new_n500));
  AOI21_X1  g314(.A(new_n495), .B1(new_n494), .B2(new_n498), .ZN(new_n501));
  OAI21_X1  g315(.A(new_n486), .B1(new_n500), .B2(new_n501), .ZN(new_n502));
  INV_X1    g316(.A(new_n502), .ZN(new_n503));
  INV_X1    g317(.A(new_n437), .ZN(new_n504));
  AOI21_X1  g318(.A(new_n504), .B1(new_n433), .B2(new_n434), .ZN(new_n505));
  OAI21_X1  g319(.A(KEYINPUT94), .B1(new_n505), .B2(new_n440), .ZN(new_n506));
  NAND4_X1  g320(.A1(new_n381), .A2(new_n442), .A3(new_n503), .A4(new_n506), .ZN(new_n507));
  OAI211_X1 g321(.A(new_n339), .B(new_n201), .C1(new_n212), .C2(new_n218), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n508), .A2(KEYINPUT68), .ZN(new_n509));
  INV_X1    g323(.A(new_n332), .ZN(new_n510));
  NOR2_X1   g324(.A1(new_n330), .A2(G137), .ZN(new_n511));
  OAI21_X1  g325(.A(G131), .B1(new_n510), .B2(new_n511), .ZN(new_n512));
  NAND3_X1  g326(.A1(new_n227), .A2(new_n338), .A3(new_n512), .ZN(new_n513));
  INV_X1    g327(.A(KEYINPUT68), .ZN(new_n514));
  NAND4_X1  g328(.A1(new_n327), .A2(new_n514), .A3(new_n339), .A4(new_n201), .ZN(new_n515));
  NAND3_X1  g329(.A1(new_n509), .A2(new_n513), .A3(new_n515), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n516), .A2(new_n246), .ZN(new_n517));
  INV_X1    g331(.A(new_n246), .ZN(new_n518));
  NAND3_X1  g332(.A1(new_n508), .A2(new_n513), .A3(new_n518), .ZN(new_n519));
  INV_X1    g333(.A(new_n519), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n520), .A2(KEYINPUT28), .ZN(new_n521));
  INV_X1    g335(.A(KEYINPUT28), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n519), .A2(new_n522), .ZN(new_n523));
  AND3_X1   g337(.A1(new_n517), .A2(new_n521), .A3(new_n523), .ZN(new_n524));
  XOR2_X1   g338(.A(KEYINPUT70), .B(KEYINPUT27), .Z(new_n525));
  INV_X1    g339(.A(G210), .ZN(new_n526));
  NOR3_X1   g340(.A1(new_n526), .A2(G237), .A3(G953), .ZN(new_n527));
  XNOR2_X1  g341(.A(new_n525), .B(new_n527), .ZN(new_n528));
  XNOR2_X1  g342(.A(KEYINPUT26), .B(G101), .ZN(new_n529));
  XNOR2_X1  g343(.A(new_n528), .B(new_n529), .ZN(new_n530));
  AOI21_X1  g344(.A(KEYINPUT29), .B1(new_n524), .B2(new_n530), .ZN(new_n531));
  INV_X1    g345(.A(new_n530), .ZN(new_n532));
  NAND3_X1  g346(.A1(new_n508), .A2(new_n513), .A3(KEYINPUT30), .ZN(new_n533));
  INV_X1    g347(.A(new_n533), .ZN(new_n534));
  INV_X1    g348(.A(KEYINPUT30), .ZN(new_n535));
  AOI211_X1 g349(.A(new_n518), .B(new_n534), .C1(new_n516), .C2(new_n535), .ZN(new_n536));
  OAI21_X1  g350(.A(new_n532), .B1(new_n536), .B2(new_n520), .ZN(new_n537));
  AOI21_X1  g351(.A(G902), .B1(new_n531), .B2(new_n537), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n508), .A2(new_n513), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n539), .A2(new_n246), .ZN(new_n540));
  NAND3_X1  g354(.A1(new_n540), .A2(KEYINPUT71), .A3(new_n519), .ZN(new_n541));
  INV_X1    g355(.A(KEYINPUT71), .ZN(new_n542));
  NAND3_X1  g356(.A1(new_n539), .A2(new_n542), .A3(new_n246), .ZN(new_n543));
  NAND3_X1  g357(.A1(new_n541), .A2(KEYINPUT28), .A3(new_n543), .ZN(new_n544));
  NAND2_X1  g358(.A1(new_n544), .A2(new_n523), .ZN(new_n545));
  NAND2_X1  g359(.A1(new_n545), .A2(KEYINPUT72), .ZN(new_n546));
  INV_X1    g360(.A(KEYINPUT72), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n544), .A2(new_n547), .ZN(new_n548));
  NAND4_X1  g362(.A1(new_n546), .A2(KEYINPUT29), .A3(new_n530), .A4(new_n548), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n538), .A2(new_n549), .ZN(new_n550));
  NAND2_X1  g364(.A1(new_n550), .A2(G472), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n516), .A2(new_n535), .ZN(new_n552));
  NAND3_X1  g366(.A1(new_n552), .A2(new_n246), .A3(new_n533), .ZN(new_n553));
  NAND3_X1  g367(.A1(new_n553), .A2(new_n530), .A3(new_n519), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n554), .A2(KEYINPUT31), .ZN(new_n555));
  NAND3_X1  g369(.A1(new_n517), .A2(new_n521), .A3(new_n523), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n556), .A2(new_n532), .ZN(new_n557));
  INV_X1    g371(.A(KEYINPUT31), .ZN(new_n558));
  NAND4_X1  g372(.A1(new_n553), .A2(new_n558), .A3(new_n530), .A4(new_n519), .ZN(new_n559));
  NAND3_X1  g373(.A1(new_n555), .A2(new_n557), .A3(new_n559), .ZN(new_n560));
  NOR2_X1   g374(.A1(G472), .A2(G902), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n560), .A2(new_n561), .ZN(new_n562));
  INV_X1    g376(.A(KEYINPUT32), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  NAND3_X1  g378(.A1(new_n560), .A2(KEYINPUT32), .A3(new_n561), .ZN(new_n565));
  NAND3_X1  g379(.A1(new_n551), .A2(new_n564), .A3(new_n565), .ZN(new_n566));
  NAND3_X1  g380(.A1(new_n308), .A2(G221), .A3(G234), .ZN(new_n567));
  XNOR2_X1  g381(.A(new_n567), .B(KEYINPUT22), .ZN(new_n568));
  XNOR2_X1  g382(.A(new_n568), .B(new_n333), .ZN(new_n569));
  XOR2_X1   g383(.A(KEYINPUT24), .B(G110), .Z(new_n570));
  XNOR2_X1  g384(.A(G119), .B(G128), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n570), .A2(new_n571), .ZN(new_n572));
  INV_X1    g386(.A(KEYINPUT23), .ZN(new_n573));
  OAI21_X1  g387(.A(new_n573), .B1(new_n237), .B2(G128), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n237), .A2(G128), .ZN(new_n575));
  NAND3_X1  g389(.A1(new_n196), .A2(KEYINPUT23), .A3(G119), .ZN(new_n576));
  NAND3_X1  g390(.A1(new_n574), .A2(new_n575), .A3(new_n576), .ZN(new_n577));
  NAND2_X1  g391(.A1(new_n577), .A2(G110), .ZN(new_n578));
  NAND2_X1  g392(.A1(new_n578), .A2(KEYINPUT74), .ZN(new_n579));
  INV_X1    g393(.A(KEYINPUT74), .ZN(new_n580));
  NAND3_X1  g394(.A1(new_n577), .A2(new_n580), .A3(G110), .ZN(new_n581));
  NAND2_X1  g395(.A1(new_n579), .A2(new_n581), .ZN(new_n582));
  OAI211_X1 g396(.A(new_n572), .B(new_n582), .C1(new_n470), .C2(new_n476), .ZN(new_n583));
  INV_X1    g397(.A(KEYINPUT77), .ZN(new_n584));
  OAI22_X1  g398(.A1(new_n577), .A2(G110), .B1(new_n570), .B2(new_n571), .ZN(new_n585));
  NAND3_X1  g399(.A1(new_n455), .A2(new_n487), .A3(new_n585), .ZN(new_n586));
  AND3_X1   g400(.A1(new_n583), .A2(new_n584), .A3(new_n586), .ZN(new_n587));
  AOI21_X1  g401(.A(new_n584), .B1(new_n583), .B2(new_n586), .ZN(new_n588));
  OAI21_X1  g402(.A(new_n569), .B1(new_n587), .B2(new_n588), .ZN(new_n589));
  INV_X1    g403(.A(new_n569), .ZN(new_n590));
  NAND3_X1  g404(.A1(new_n583), .A2(new_n586), .A3(new_n590), .ZN(new_n591));
  NAND3_X1  g405(.A1(new_n589), .A2(new_n288), .A3(new_n591), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n592), .A2(KEYINPUT25), .ZN(new_n593));
  INV_X1    g407(.A(G234), .ZN(new_n594));
  OAI21_X1  g408(.A(G217), .B1(new_n594), .B2(G902), .ZN(new_n595));
  XNOR2_X1  g409(.A(new_n595), .B(KEYINPUT73), .ZN(new_n596));
  INV_X1    g410(.A(new_n596), .ZN(new_n597));
  INV_X1    g411(.A(KEYINPUT25), .ZN(new_n598));
  NAND4_X1  g412(.A1(new_n589), .A2(new_n598), .A3(new_n288), .A4(new_n591), .ZN(new_n599));
  NAND3_X1  g413(.A1(new_n593), .A2(new_n597), .A3(new_n599), .ZN(new_n600));
  NOR2_X1   g414(.A1(new_n597), .A2(G902), .ZN(new_n601));
  NAND3_X1  g415(.A1(new_n589), .A2(new_n591), .A3(new_n601), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n600), .A2(new_n602), .ZN(new_n603));
  INV_X1    g417(.A(new_n603), .ZN(new_n604));
  NAND2_X1  g418(.A1(new_n566), .A2(new_n604), .ZN(new_n605));
  NOR2_X1   g419(.A1(new_n507), .A2(new_n605), .ZN(new_n606));
  XNOR2_X1  g420(.A(new_n606), .B(new_n255), .ZN(G3));
  XNOR2_X1  g421(.A(KEYINPUT96), .B(KEYINPUT33), .ZN(new_n608));
  INV_X1    g422(.A(new_n608), .ZN(new_n609));
  NAND3_X1  g423(.A1(new_n427), .A2(new_n430), .A3(new_n609), .ZN(new_n610));
  NAND3_X1  g424(.A1(new_n424), .A2(KEYINPUT33), .A3(new_n426), .ZN(new_n611));
  AND2_X1   g425(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  INV_X1    g426(.A(KEYINPUT97), .ZN(new_n613));
  NAND4_X1  g427(.A1(new_n612), .A2(new_n613), .A3(G478), .A4(new_n288), .ZN(new_n614));
  NAND2_X1  g428(.A1(new_n435), .A2(new_n436), .ZN(new_n615));
  NAND4_X1  g429(.A1(new_n610), .A2(G478), .A3(new_n288), .A4(new_n611), .ZN(new_n616));
  NAND2_X1  g430(.A1(new_n616), .A2(KEYINPUT97), .ZN(new_n617));
  NAND3_X1  g431(.A1(new_n614), .A2(new_n615), .A3(new_n617), .ZN(new_n618));
  NAND2_X1  g432(.A1(new_n618), .A2(new_n502), .ZN(new_n619));
  INV_X1    g433(.A(KEYINPUT95), .ZN(new_n620));
  INV_X1    g434(.A(new_n302), .ZN(new_n621));
  NAND2_X1  g435(.A1(new_n301), .A2(new_n621), .ZN(new_n622));
  NAND2_X1  g436(.A1(new_n622), .A2(new_n305), .ZN(new_n623));
  AOI21_X1  g437(.A(new_n620), .B1(new_n623), .B2(new_n307), .ZN(new_n624));
  INV_X1    g438(.A(new_n624), .ZN(new_n625));
  INV_X1    g439(.A(new_n307), .ZN(new_n626));
  AOI211_X1 g440(.A(KEYINPUT95), .B(new_n626), .C1(new_n622), .C2(new_n305), .ZN(new_n627));
  INV_X1    g441(.A(new_n627), .ZN(new_n628));
  NAND3_X1  g442(.A1(new_n625), .A2(new_n628), .A3(new_n318), .ZN(new_n629));
  OAI21_X1  g443(.A(KEYINPUT98), .B1(new_n619), .B2(new_n629), .ZN(new_n630));
  NOR3_X1   g444(.A1(new_n624), .A2(new_n627), .A3(new_n317), .ZN(new_n631));
  INV_X1    g445(.A(KEYINPUT98), .ZN(new_n632));
  NAND4_X1  g446(.A1(new_n631), .A2(new_n632), .A3(new_n502), .A4(new_n618), .ZN(new_n633));
  NAND2_X1  g447(.A1(new_n630), .A2(new_n633), .ZN(new_n634));
  NAND2_X1  g448(.A1(new_n560), .A2(new_n288), .ZN(new_n635));
  AOI22_X1  g449(.A1(new_n635), .A2(G472), .B1(new_n560), .B2(new_n561), .ZN(new_n636));
  NOR3_X1   g450(.A1(new_n377), .A2(new_n603), .A3(new_n380), .ZN(new_n637));
  NAND2_X1  g451(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  INV_X1    g452(.A(new_n638), .ZN(new_n639));
  NAND2_X1  g453(.A1(new_n634), .A2(new_n639), .ZN(new_n640));
  XOR2_X1   g454(.A(KEYINPUT34), .B(G104), .Z(new_n641));
  XNOR2_X1  g455(.A(new_n640), .B(new_n641), .ZN(G6));
  NAND2_X1  g456(.A1(new_n442), .A2(new_n506), .ZN(new_n643));
  INV_X1    g457(.A(new_n501), .ZN(new_n644));
  NAND3_X1  g458(.A1(new_n644), .A2(KEYINPUT99), .A3(new_n499), .ZN(new_n645));
  OR2_X1    g459(.A1(new_n499), .A2(KEYINPUT99), .ZN(new_n646));
  AND3_X1   g460(.A1(new_n645), .A2(new_n486), .A3(new_n646), .ZN(new_n647));
  AND3_X1   g461(.A1(new_n643), .A2(new_n631), .A3(new_n647), .ZN(new_n648));
  NAND2_X1  g462(.A1(new_n648), .A2(new_n639), .ZN(new_n649));
  XOR2_X1   g463(.A(KEYINPUT35), .B(G107), .Z(new_n650));
  XNOR2_X1  g464(.A(new_n649), .B(new_n650), .ZN(G9));
  NOR2_X1   g465(.A1(new_n587), .A2(new_n588), .ZN(new_n652));
  NOR2_X1   g466(.A1(new_n569), .A2(KEYINPUT36), .ZN(new_n653));
  XOR2_X1   g467(.A(new_n652), .B(new_n653), .Z(new_n654));
  NAND2_X1  g468(.A1(new_n654), .A2(new_n601), .ZN(new_n655));
  NAND2_X1  g469(.A1(new_n655), .A2(new_n600), .ZN(new_n656));
  NAND2_X1  g470(.A1(new_n656), .A2(KEYINPUT100), .ZN(new_n657));
  INV_X1    g471(.A(KEYINPUT100), .ZN(new_n658));
  NAND3_X1  g472(.A1(new_n655), .A2(new_n658), .A3(new_n600), .ZN(new_n659));
  NAND2_X1  g473(.A1(new_n657), .A2(new_n659), .ZN(new_n660));
  NAND2_X1  g474(.A1(new_n660), .A2(new_n636), .ZN(new_n661));
  NOR2_X1   g475(.A1(new_n507), .A2(new_n661), .ZN(new_n662));
  XNOR2_X1  g476(.A(new_n662), .B(KEYINPUT37), .ZN(new_n663));
  XNOR2_X1  g477(.A(new_n663), .B(G110), .ZN(G12));
  NOR2_X1   g478(.A1(new_n377), .A2(new_n380), .ZN(new_n665));
  AND2_X1   g479(.A1(new_n566), .A2(new_n665), .ZN(new_n666));
  NOR2_X1   g480(.A1(new_n624), .A2(new_n627), .ZN(new_n667));
  NAND2_X1  g481(.A1(new_n660), .A2(new_n667), .ZN(new_n668));
  INV_X1    g482(.A(new_n668), .ZN(new_n669));
  OR2_X1    g483(.A1(new_n315), .A2(G900), .ZN(new_n670));
  NAND2_X1  g484(.A1(new_n670), .A2(new_n311), .ZN(new_n671));
  NAND4_X1  g485(.A1(new_n645), .A2(new_n646), .A3(new_n486), .A4(new_n671), .ZN(new_n672));
  AOI21_X1  g486(.A(new_n672), .B1(new_n442), .B2(new_n506), .ZN(new_n673));
  NAND3_X1  g487(.A1(new_n666), .A2(new_n669), .A3(new_n673), .ZN(new_n674));
  XNOR2_X1  g488(.A(new_n674), .B(G128), .ZN(G30));
  INV_X1    g489(.A(new_n656), .ZN(new_n676));
  AND4_X1   g490(.A1(new_n502), .A2(new_n643), .A3(new_n307), .A4(new_n676), .ZN(new_n677));
  XNOR2_X1  g491(.A(new_n677), .B(KEYINPUT102), .ZN(new_n678));
  AND2_X1   g492(.A1(new_n564), .A2(new_n565), .ZN(new_n679));
  NAND3_X1  g493(.A1(new_n541), .A2(new_n532), .A3(new_n543), .ZN(new_n680));
  OR2_X1    g494(.A1(new_n680), .A2(KEYINPUT101), .ZN(new_n681));
  NAND2_X1  g495(.A1(new_n681), .A2(new_n554), .ZN(new_n682));
  AOI21_X1  g496(.A(new_n682), .B1(KEYINPUT101), .B2(new_n680), .ZN(new_n683));
  OAI21_X1  g497(.A(G472), .B1(new_n683), .B2(G902), .ZN(new_n684));
  NAND2_X1  g498(.A1(new_n679), .A2(new_n684), .ZN(new_n685));
  XOR2_X1   g499(.A(new_n306), .B(KEYINPUT38), .Z(new_n686));
  INV_X1    g500(.A(new_n686), .ZN(new_n687));
  NAND3_X1  g501(.A1(new_n678), .A2(new_n685), .A3(new_n687), .ZN(new_n688));
  INV_X1    g502(.A(KEYINPUT103), .ZN(new_n689));
  OR2_X1    g503(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  NAND2_X1  g504(.A1(new_n688), .A2(new_n689), .ZN(new_n691));
  XOR2_X1   g505(.A(new_n671), .B(KEYINPUT39), .Z(new_n692));
  OR3_X1    g506(.A1(new_n377), .A2(new_n380), .A3(new_n692), .ZN(new_n693));
  XOR2_X1   g507(.A(new_n693), .B(KEYINPUT40), .Z(new_n694));
  NAND3_X1  g508(.A1(new_n690), .A2(new_n691), .A3(new_n694), .ZN(new_n695));
  XOR2_X1   g509(.A(new_n695), .B(new_n207), .Z(G45));
  AND3_X1   g510(.A1(new_n618), .A2(new_n502), .A3(new_n671), .ZN(new_n697));
  NAND3_X1  g511(.A1(new_n666), .A2(new_n669), .A3(new_n697), .ZN(new_n698));
  XNOR2_X1  g512(.A(new_n698), .B(G146), .ZN(G48));
  INV_X1    g513(.A(KEYINPUT104), .ZN(new_n700));
  NAND2_X1  g514(.A1(new_n366), .A2(new_n376), .ZN(new_n701));
  NAND2_X1  g515(.A1(new_n375), .A2(new_n288), .ZN(new_n702));
  NAND2_X1  g516(.A1(new_n702), .A2(G469), .ZN(new_n703));
  NAND2_X1  g517(.A1(new_n701), .A2(new_n703), .ZN(new_n704));
  NOR2_X1   g518(.A1(new_n704), .A2(new_n380), .ZN(new_n705));
  NAND3_X1  g519(.A1(new_n566), .A2(new_n604), .A3(new_n705), .ZN(new_n706));
  INV_X1    g520(.A(new_n706), .ZN(new_n707));
  AOI21_X1  g521(.A(new_n700), .B1(new_n634), .B2(new_n707), .ZN(new_n708));
  AOI211_X1 g522(.A(KEYINPUT104), .B(new_n706), .C1(new_n630), .C2(new_n633), .ZN(new_n709));
  NOR2_X1   g523(.A1(new_n708), .A2(new_n709), .ZN(new_n710));
  XNOR2_X1  g524(.A(new_n710), .B(KEYINPUT41), .ZN(new_n711));
  XNOR2_X1  g525(.A(new_n711), .B(new_n267), .ZN(G15));
  NAND2_X1  g526(.A1(new_n648), .A2(new_n707), .ZN(new_n713));
  XNOR2_X1  g527(.A(new_n713), .B(G116), .ZN(G18));
  INV_X1    g528(.A(new_n704), .ZN(new_n715));
  INV_X1    g529(.A(new_n380), .ZN(new_n716));
  NAND2_X1  g530(.A1(new_n715), .A2(new_n716), .ZN(new_n717));
  NOR2_X1   g531(.A1(new_n717), .A2(new_n317), .ZN(new_n718));
  AND2_X1   g532(.A1(new_n718), .A2(new_n566), .ZN(new_n719));
  NOR3_X1   g533(.A1(new_n668), .A2(new_n643), .A3(new_n502), .ZN(new_n720));
  NAND2_X1  g534(.A1(new_n719), .A2(new_n720), .ZN(new_n721));
  XNOR2_X1  g535(.A(new_n721), .B(G119), .ZN(G21));
  AOI21_X1  g536(.A(new_n439), .B1(new_n438), .B2(new_n441), .ZN(new_n723));
  NOR3_X1   g537(.A1(new_n505), .A2(KEYINPUT94), .A3(new_n440), .ZN(new_n724));
  OAI211_X1 g538(.A(new_n502), .B(new_n667), .C1(new_n723), .C2(new_n724), .ZN(new_n725));
  INV_X1    g539(.A(KEYINPUT105), .ZN(new_n726));
  NAND2_X1  g540(.A1(new_n725), .A2(new_n726), .ZN(new_n727));
  NAND4_X1  g541(.A1(new_n643), .A2(KEYINPUT105), .A3(new_n502), .A4(new_n667), .ZN(new_n728));
  NAND2_X1  g542(.A1(new_n727), .A2(new_n728), .ZN(new_n729));
  NAND2_X1  g543(.A1(new_n546), .A2(new_n548), .ZN(new_n730));
  NAND2_X1  g544(.A1(new_n730), .A2(new_n532), .ZN(new_n731));
  AND2_X1   g545(.A1(new_n555), .A2(new_n559), .ZN(new_n732));
  AOI211_X1 g546(.A(G472), .B(G902), .C1(new_n731), .C2(new_n732), .ZN(new_n733));
  NAND2_X1  g547(.A1(new_n635), .A2(G472), .ZN(new_n734));
  INV_X1    g548(.A(new_n734), .ZN(new_n735));
  NOR3_X1   g549(.A1(new_n733), .A2(new_n735), .A3(new_n603), .ZN(new_n736));
  NAND3_X1  g550(.A1(new_n729), .A2(new_n718), .A3(new_n736), .ZN(new_n737));
  NAND2_X1  g551(.A1(new_n737), .A2(KEYINPUT106), .ZN(new_n738));
  INV_X1    g552(.A(KEYINPUT106), .ZN(new_n739));
  NAND4_X1  g553(.A1(new_n729), .A2(new_n739), .A3(new_n718), .A4(new_n736), .ZN(new_n740));
  NAND2_X1  g554(.A1(new_n738), .A2(new_n740), .ZN(new_n741));
  XNOR2_X1  g555(.A(new_n741), .B(G122), .ZN(G24));
  NOR3_X1   g556(.A1(new_n733), .A2(new_n735), .A3(new_n676), .ZN(new_n743));
  AND2_X1   g557(.A1(new_n667), .A2(new_n705), .ZN(new_n744));
  NAND3_X1  g558(.A1(new_n743), .A2(new_n697), .A3(new_n744), .ZN(new_n745));
  XNOR2_X1  g559(.A(KEYINPUT107), .B(G125), .ZN(new_n746));
  XNOR2_X1  g560(.A(new_n745), .B(new_n746), .ZN(G27));
  INV_X1    g561(.A(KEYINPUT42), .ZN(new_n748));
  INV_X1    g562(.A(KEYINPUT108), .ZN(new_n749));
  NAND3_X1  g563(.A1(new_n749), .A2(new_n288), .A3(G469), .ZN(new_n750));
  OAI22_X1  g564(.A1(new_n360), .A2(new_n749), .B1(new_n359), .B2(new_n750), .ZN(new_n751));
  AOI21_X1  g565(.A(new_n306), .B1(new_n751), .B2(new_n701), .ZN(new_n752));
  NOR2_X1   g566(.A1(new_n380), .A2(new_n626), .ZN(new_n753));
  AND2_X1   g567(.A1(new_n752), .A2(new_n753), .ZN(new_n754));
  NAND3_X1  g568(.A1(new_n754), .A2(new_n566), .A3(new_n604), .ZN(new_n755));
  XNOR2_X1  g569(.A(new_n616), .B(new_n613), .ZN(new_n756));
  AOI21_X1  g570(.A(new_n503), .B1(new_n756), .B2(new_n615), .ZN(new_n757));
  NAND2_X1  g571(.A1(new_n757), .A2(new_n671), .ZN(new_n758));
  OAI21_X1  g572(.A(new_n748), .B1(new_n755), .B2(new_n758), .ZN(new_n759));
  AND2_X1   g573(.A1(new_n566), .A2(new_n604), .ZN(new_n760));
  NAND4_X1  g574(.A1(new_n760), .A2(KEYINPUT42), .A3(new_n697), .A4(new_n754), .ZN(new_n761));
  NAND2_X1  g575(.A1(new_n759), .A2(new_n761), .ZN(new_n762));
  XNOR2_X1  g576(.A(new_n762), .B(G131), .ZN(G33));
  NAND3_X1  g577(.A1(new_n760), .A2(new_n673), .A3(new_n754), .ZN(new_n764));
  XNOR2_X1  g578(.A(new_n764), .B(G134), .ZN(G36));
  NAND2_X1  g579(.A1(new_n618), .A2(new_n503), .ZN(new_n766));
  AOI21_X1  g580(.A(KEYINPUT43), .B1(new_n503), .B2(KEYINPUT109), .ZN(new_n767));
  NOR2_X1   g581(.A1(new_n766), .A2(new_n767), .ZN(new_n768));
  INV_X1    g582(.A(new_n768), .ZN(new_n769));
  NAND2_X1  g583(.A1(new_n766), .A2(new_n767), .ZN(new_n770));
  NAND2_X1  g584(.A1(new_n769), .A2(new_n770), .ZN(new_n771));
  INV_X1    g585(.A(new_n636), .ZN(new_n772));
  NAND3_X1  g586(.A1(new_n771), .A2(new_n772), .A3(new_n656), .ZN(new_n773));
  INV_X1    g587(.A(KEYINPUT44), .ZN(new_n774));
  NAND2_X1  g588(.A1(new_n773), .A2(new_n774), .ZN(new_n775));
  XNOR2_X1  g589(.A(new_n359), .B(KEYINPUT45), .ZN(new_n776));
  NAND2_X1  g590(.A1(new_n776), .A2(G469), .ZN(new_n777));
  NAND2_X1  g591(.A1(G469), .A2(G902), .ZN(new_n778));
  NAND2_X1  g592(.A1(new_n777), .A2(new_n778), .ZN(new_n779));
  INV_X1    g593(.A(KEYINPUT46), .ZN(new_n780));
  NOR2_X1   g594(.A1(new_n779), .A2(new_n780), .ZN(new_n781));
  INV_X1    g595(.A(new_n701), .ZN(new_n782));
  AOI21_X1  g596(.A(KEYINPUT46), .B1(new_n777), .B2(new_n778), .ZN(new_n783));
  NOR3_X1   g597(.A1(new_n781), .A2(new_n782), .A3(new_n783), .ZN(new_n784));
  NOR3_X1   g598(.A1(new_n784), .A2(new_n380), .A3(new_n692), .ZN(new_n785));
  NOR2_X1   g599(.A1(new_n306), .A2(new_n626), .ZN(new_n786));
  NAND4_X1  g600(.A1(new_n771), .A2(KEYINPUT44), .A3(new_n772), .A4(new_n656), .ZN(new_n787));
  NAND4_X1  g601(.A1(new_n775), .A2(new_n785), .A3(new_n786), .A4(new_n787), .ZN(new_n788));
  XNOR2_X1  g602(.A(new_n788), .B(G137), .ZN(G39));
  INV_X1    g603(.A(new_n786), .ZN(new_n790));
  NOR4_X1   g604(.A1(new_n758), .A2(new_n566), .A3(new_n604), .A4(new_n790), .ZN(new_n791));
  INV_X1    g605(.A(KEYINPUT110), .ZN(new_n792));
  OR2_X1    g606(.A1(new_n791), .A2(new_n792), .ZN(new_n793));
  OAI21_X1  g607(.A(KEYINPUT47), .B1(new_n784), .B2(new_n380), .ZN(new_n794));
  OR3_X1    g608(.A1(new_n784), .A2(KEYINPUT47), .A3(new_n380), .ZN(new_n795));
  NAND2_X1  g609(.A1(new_n791), .A2(new_n792), .ZN(new_n796));
  NAND4_X1  g610(.A1(new_n793), .A2(new_n794), .A3(new_n795), .A4(new_n796), .ZN(new_n797));
  XNOR2_X1  g611(.A(new_n797), .B(KEYINPUT111), .ZN(new_n798));
  XNOR2_X1  g612(.A(new_n798), .B(new_n456), .ZN(G42));
  INV_X1    g613(.A(new_n770), .ZN(new_n800));
  OAI211_X1 g614(.A(new_n312), .B(new_n736), .C1(new_n800), .C2(new_n768), .ZN(new_n801));
  NOR2_X1   g615(.A1(new_n801), .A2(new_n307), .ZN(new_n802));
  NOR2_X1   g616(.A1(new_n687), .A2(new_n717), .ZN(new_n803));
  AND3_X1   g617(.A1(new_n802), .A2(KEYINPUT50), .A3(new_n803), .ZN(new_n804));
  AOI21_X1  g618(.A(KEYINPUT50), .B1(new_n802), .B2(new_n803), .ZN(new_n805));
  OR2_X1    g619(.A1(new_n804), .A2(new_n805), .ZN(new_n806));
  AOI21_X1  g620(.A(new_n311), .B1(new_n769), .B2(new_n770), .ZN(new_n807));
  NOR2_X1   g621(.A1(new_n717), .A2(new_n790), .ZN(new_n808));
  NAND3_X1  g622(.A1(new_n807), .A2(new_n743), .A3(new_n808), .ZN(new_n809));
  INV_X1    g623(.A(new_n685), .ZN(new_n810));
  NOR2_X1   g624(.A1(new_n603), .A2(new_n311), .ZN(new_n811));
  NAND3_X1  g625(.A1(new_n810), .A2(new_n808), .A3(new_n811), .ZN(new_n812));
  INV_X1    g626(.A(KEYINPUT118), .ZN(new_n813));
  XNOR2_X1  g627(.A(new_n812), .B(new_n813), .ZN(new_n814));
  NOR2_X1   g628(.A1(new_n814), .A2(new_n502), .ZN(new_n815));
  INV_X1    g629(.A(new_n618), .ZN(new_n816));
  INV_X1    g630(.A(new_n801), .ZN(new_n817));
  NAND2_X1  g631(.A1(new_n795), .A2(new_n794), .ZN(new_n818));
  NAND2_X1  g632(.A1(new_n715), .A2(new_n380), .ZN(new_n819));
  AOI21_X1  g633(.A(new_n790), .B1(new_n818), .B2(new_n819), .ZN(new_n820));
  AOI22_X1  g634(.A1(new_n815), .A2(new_n816), .B1(new_n817), .B2(new_n820), .ZN(new_n821));
  NAND3_X1  g635(.A1(new_n806), .A2(new_n809), .A3(new_n821), .ZN(new_n822));
  INV_X1    g636(.A(KEYINPUT51), .ZN(new_n823));
  NAND2_X1  g637(.A1(new_n822), .A2(new_n823), .ZN(new_n824));
  INV_X1    g638(.A(KEYINPUT119), .ZN(new_n825));
  NAND2_X1  g639(.A1(new_n309), .A2(new_n825), .ZN(new_n826));
  NAND4_X1  g640(.A1(new_n806), .A2(new_n821), .A3(KEYINPUT51), .A4(new_n809), .ZN(new_n827));
  NAND2_X1  g641(.A1(new_n817), .A2(new_n744), .ZN(new_n828));
  OAI221_X1 g642(.A(new_n828), .B1(new_n825), .B2(new_n309), .C1(new_n814), .C2(new_n619), .ZN(new_n829));
  NAND3_X1  g643(.A1(new_n807), .A2(new_n760), .A3(new_n808), .ZN(new_n830));
  NAND2_X1  g644(.A1(new_n830), .A2(KEYINPUT48), .ZN(new_n831));
  OR2_X1    g645(.A1(new_n830), .A2(KEYINPUT48), .ZN(new_n832));
  AOI21_X1  g646(.A(new_n829), .B1(new_n831), .B2(new_n832), .ZN(new_n833));
  NAND4_X1  g647(.A1(new_n824), .A2(new_n826), .A3(new_n827), .A4(new_n833), .ZN(new_n834));
  XNOR2_X1  g648(.A(new_n834), .B(KEYINPUT120), .ZN(new_n835));
  INV_X1    g649(.A(KEYINPUT117), .ZN(new_n836));
  AND3_X1   g650(.A1(new_n698), .A2(new_n674), .A3(new_n745), .ZN(new_n837));
  AOI21_X1  g651(.A(new_n380), .B1(new_n311), .B2(new_n670), .ZN(new_n838));
  AOI21_X1  g652(.A(new_n656), .B1(new_n701), .B2(new_n751), .ZN(new_n839));
  NAND4_X1  g653(.A1(new_n729), .A2(new_n685), .A3(new_n838), .A4(new_n839), .ZN(new_n840));
  INV_X1    g654(.A(KEYINPUT52), .ZN(new_n841));
  AND3_X1   g655(.A1(new_n837), .A2(new_n840), .A3(new_n841), .ZN(new_n842));
  AOI21_X1  g656(.A(new_n841), .B1(new_n837), .B2(new_n840), .ZN(new_n843));
  NOR2_X1   g657(.A1(new_n842), .A2(new_n843), .ZN(new_n844));
  AOI22_X1  g658(.A1(new_n719), .A2(new_n720), .B1(new_n648), .B2(new_n707), .ZN(new_n845));
  OAI21_X1  g659(.A(new_n845), .B1(new_n708), .B2(new_n709), .ZN(new_n846));
  AOI21_X1  g660(.A(new_n846), .B1(new_n740), .B2(new_n738), .ZN(new_n847));
  AOI21_X1  g661(.A(new_n502), .B1(new_n438), .B2(new_n441), .ZN(new_n848));
  INV_X1    g662(.A(new_n319), .ZN(new_n849));
  NAND4_X1  g663(.A1(new_n848), .A2(new_n636), .A3(new_n637), .A4(new_n849), .ZN(new_n850));
  OAI21_X1  g664(.A(new_n850), .B1(new_n507), .B2(new_n661), .ZN(new_n851));
  INV_X1    g665(.A(KEYINPUT113), .ZN(new_n852));
  NAND2_X1  g666(.A1(new_n851), .A2(new_n852), .ZN(new_n853));
  AND4_X1   g667(.A1(new_n503), .A2(new_n381), .A3(new_n506), .A4(new_n442), .ZN(new_n854));
  AND3_X1   g668(.A1(new_n636), .A2(new_n637), .A3(new_n849), .ZN(new_n855));
  AOI22_X1  g669(.A1(new_n854), .A2(new_n760), .B1(new_n757), .B2(new_n855), .ZN(new_n856));
  OAI211_X1 g670(.A(KEYINPUT113), .B(new_n850), .C1(new_n507), .C2(new_n661), .ZN(new_n857));
  NAND3_X1  g671(.A1(new_n853), .A2(new_n856), .A3(new_n857), .ZN(new_n858));
  INV_X1    g672(.A(KEYINPUT114), .ZN(new_n859));
  NAND2_X1  g673(.A1(new_n858), .A2(new_n859), .ZN(new_n860));
  NAND4_X1  g674(.A1(new_n853), .A2(new_n856), .A3(KEYINPUT114), .A4(new_n857), .ZN(new_n861));
  NAND2_X1  g675(.A1(new_n860), .A2(new_n861), .ZN(new_n862));
  NAND2_X1  g676(.A1(new_n566), .A2(new_n665), .ZN(new_n863));
  NAND3_X1  g677(.A1(new_n660), .A2(new_n438), .A3(new_n441), .ZN(new_n864));
  OR4_X1    g678(.A1(new_n863), .A2(new_n864), .A3(new_n672), .A4(new_n790), .ZN(new_n865));
  NAND3_X1  g679(.A1(new_n743), .A2(new_n697), .A3(new_n754), .ZN(new_n866));
  AND4_X1   g680(.A1(new_n762), .A2(new_n764), .A3(new_n865), .A4(new_n866), .ZN(new_n867));
  NAND4_X1  g681(.A1(new_n844), .A2(new_n847), .A3(new_n862), .A4(new_n867), .ZN(new_n868));
  INV_X1    g682(.A(KEYINPUT53), .ZN(new_n869));
  OAI21_X1  g683(.A(new_n836), .B1(new_n868), .B2(new_n869), .ZN(new_n870));
  INV_X1    g684(.A(KEYINPUT54), .ZN(new_n871));
  XNOR2_X1  g685(.A(KEYINPUT116), .B(KEYINPUT53), .ZN(new_n872));
  INV_X1    g686(.A(new_n872), .ZN(new_n873));
  NAND2_X1  g687(.A1(new_n868), .A2(new_n873), .ZN(new_n874));
  NAND2_X1  g688(.A1(new_n721), .A2(new_n713), .ZN(new_n875));
  NAND2_X1  g689(.A1(new_n634), .A2(new_n707), .ZN(new_n876));
  NAND2_X1  g690(.A1(new_n876), .A2(KEYINPUT104), .ZN(new_n877));
  NAND3_X1  g691(.A1(new_n634), .A2(new_n700), .A3(new_n707), .ZN(new_n878));
  AOI21_X1  g692(.A(new_n875), .B1(new_n877), .B2(new_n878), .ZN(new_n879));
  NAND4_X1  g693(.A1(new_n862), .A2(new_n741), .A3(new_n879), .A4(new_n867), .ZN(new_n880));
  INV_X1    g694(.A(new_n880), .ZN(new_n881));
  NAND4_X1  g695(.A1(new_n881), .A2(KEYINPUT117), .A3(KEYINPUT53), .A4(new_n844), .ZN(new_n882));
  NAND4_X1  g696(.A1(new_n870), .A2(new_n871), .A3(new_n874), .A4(new_n882), .ZN(new_n883));
  NAND2_X1  g697(.A1(new_n880), .A2(KEYINPUT115), .ZN(new_n884));
  INV_X1    g698(.A(KEYINPUT115), .ZN(new_n885));
  NAND4_X1  g699(.A1(new_n847), .A2(new_n885), .A3(new_n862), .A4(new_n867), .ZN(new_n886));
  NAND3_X1  g700(.A1(new_n884), .A2(new_n886), .A3(new_n844), .ZN(new_n887));
  NAND2_X1  g701(.A1(new_n837), .A2(new_n840), .ZN(new_n888));
  NAND2_X1  g702(.A1(new_n888), .A2(KEYINPUT52), .ZN(new_n889));
  NAND3_X1  g703(.A1(new_n837), .A2(new_n840), .A3(new_n841), .ZN(new_n890));
  NAND2_X1  g704(.A1(new_n889), .A2(new_n890), .ZN(new_n891));
  NOR2_X1   g705(.A1(new_n880), .A2(new_n891), .ZN(new_n892));
  AOI22_X1  g706(.A1(new_n887), .A2(new_n869), .B1(new_n892), .B2(new_n872), .ZN(new_n893));
  OAI21_X1  g707(.A(new_n883), .B1(new_n893), .B2(new_n871), .ZN(new_n894));
  OAI22_X1  g708(.A1(new_n835), .A2(new_n894), .B1(G952), .B2(G953), .ZN(new_n895));
  INV_X1    g709(.A(KEYINPUT49), .ZN(new_n896));
  OAI21_X1  g710(.A(new_n686), .B1(new_n715), .B2(new_n896), .ZN(new_n897));
  AOI21_X1  g711(.A(new_n897), .B1(new_n896), .B2(new_n715), .ZN(new_n898));
  INV_X1    g712(.A(new_n766), .ZN(new_n899));
  NAND2_X1  g713(.A1(new_n604), .A2(new_n753), .ZN(new_n900));
  XNOR2_X1  g714(.A(new_n900), .B(KEYINPUT112), .ZN(new_n901));
  NAND4_X1  g715(.A1(new_n898), .A2(new_n810), .A3(new_n899), .A4(new_n901), .ZN(new_n902));
  NAND2_X1  g716(.A1(new_n895), .A2(new_n902), .ZN(G75));
  NOR2_X1   g717(.A1(new_n308), .A2(G952), .ZN(new_n904));
  XOR2_X1   g718(.A(new_n904), .B(KEYINPUT121), .Z(new_n905));
  NAND3_X1  g719(.A1(new_n870), .A2(new_n874), .A3(new_n882), .ZN(new_n906));
  NAND3_X1  g720(.A1(new_n906), .A2(G902), .A3(new_n303), .ZN(new_n907));
  OAI21_X1  g721(.A(new_n281), .B1(new_n284), .B2(new_n286), .ZN(new_n908));
  XOR2_X1   g722(.A(new_n908), .B(new_n235), .Z(new_n909));
  XNOR2_X1  g723(.A(new_n909), .B(KEYINPUT55), .ZN(new_n910));
  NOR2_X1   g724(.A1(new_n910), .A2(KEYINPUT56), .ZN(new_n911));
  AND2_X1   g725(.A1(new_n907), .A2(new_n911), .ZN(new_n912));
  INV_X1    g726(.A(KEYINPUT56), .ZN(new_n913));
  NAND2_X1  g727(.A1(new_n906), .A2(G902), .ZN(new_n914));
  OAI21_X1  g728(.A(new_n913), .B1(new_n914), .B2(new_n526), .ZN(new_n915));
  AOI211_X1 g729(.A(new_n905), .B(new_n912), .C1(new_n910), .C2(new_n915), .ZN(G51));
  NAND2_X1  g730(.A1(new_n906), .A2(KEYINPUT54), .ZN(new_n917));
  NAND2_X1  g731(.A1(new_n917), .A2(new_n883), .ZN(new_n918));
  INV_X1    g732(.A(new_n918), .ZN(new_n919));
  XNOR2_X1  g733(.A(new_n778), .B(KEYINPUT57), .ZN(new_n920));
  OAI21_X1  g734(.A(new_n375), .B1(new_n919), .B2(new_n920), .ZN(new_n921));
  OR2_X1    g735(.A1(new_n914), .A2(new_n777), .ZN(new_n922));
  AOI21_X1  g736(.A(new_n904), .B1(new_n921), .B2(new_n922), .ZN(G54));
  INV_X1    g737(.A(KEYINPUT58), .ZN(new_n924));
  NOR2_X1   g738(.A1(new_n914), .A2(new_n924), .ZN(new_n925));
  AOI21_X1  g739(.A(new_n494), .B1(new_n925), .B2(G475), .ZN(new_n926));
  INV_X1    g740(.A(new_n494), .ZN(new_n927));
  NOR4_X1   g741(.A1(new_n914), .A2(new_n924), .A3(new_n496), .A4(new_n927), .ZN(new_n928));
  NOR3_X1   g742(.A1(new_n926), .A2(new_n904), .A3(new_n928), .ZN(G60));
  NAND2_X1  g743(.A1(G478), .A2(G902), .ZN(new_n930));
  XNOR2_X1  g744(.A(new_n930), .B(KEYINPUT59), .ZN(new_n931));
  AOI21_X1  g745(.A(KEYINPUT117), .B1(new_n892), .B2(KEYINPUT53), .ZN(new_n932));
  NOR4_X1   g746(.A1(new_n880), .A2(new_n891), .A3(new_n836), .A4(new_n869), .ZN(new_n933));
  NOR2_X1   g747(.A1(new_n932), .A2(new_n933), .ZN(new_n934));
  AOI21_X1  g748(.A(new_n871), .B1(new_n934), .B2(new_n874), .ZN(new_n935));
  INV_X1    g749(.A(new_n883), .ZN(new_n936));
  OAI211_X1 g750(.A(new_n612), .B(new_n931), .C1(new_n935), .C2(new_n936), .ZN(new_n937));
  INV_X1    g751(.A(KEYINPUT122), .ZN(new_n938));
  NAND2_X1  g752(.A1(new_n937), .A2(new_n938), .ZN(new_n939));
  NAND2_X1  g753(.A1(new_n894), .A2(new_n931), .ZN(new_n940));
  INV_X1    g754(.A(new_n612), .ZN(new_n941));
  AOI21_X1  g755(.A(new_n905), .B1(new_n940), .B2(new_n941), .ZN(new_n942));
  NAND4_X1  g756(.A1(new_n918), .A2(KEYINPUT122), .A3(new_n612), .A4(new_n931), .ZN(new_n943));
  AND3_X1   g757(.A1(new_n939), .A2(new_n942), .A3(new_n943), .ZN(G63));
  NAND2_X1  g758(.A1(G217), .A2(G902), .ZN(new_n945));
  XOR2_X1   g759(.A(new_n945), .B(KEYINPUT60), .Z(new_n946));
  NAND2_X1  g760(.A1(new_n906), .A2(new_n946), .ZN(new_n947));
  NAND2_X1  g761(.A1(new_n589), .A2(new_n591), .ZN(new_n948));
  AOI21_X1  g762(.A(new_n905), .B1(new_n947), .B2(new_n948), .ZN(new_n949));
  NAND3_X1  g763(.A1(new_n906), .A2(new_n654), .A3(new_n946), .ZN(new_n950));
  INV_X1    g764(.A(KEYINPUT123), .ZN(new_n951));
  NAND2_X1  g765(.A1(new_n950), .A2(new_n951), .ZN(new_n952));
  NAND4_X1  g766(.A1(new_n906), .A2(KEYINPUT123), .A3(new_n654), .A4(new_n946), .ZN(new_n953));
  NAND3_X1  g767(.A1(new_n949), .A2(new_n952), .A3(new_n953), .ZN(new_n954));
  INV_X1    g768(.A(KEYINPUT61), .ZN(new_n955));
  NAND2_X1  g769(.A1(new_n954), .A2(new_n955), .ZN(new_n956));
  NAND4_X1  g770(.A1(new_n949), .A2(new_n952), .A3(KEYINPUT61), .A4(new_n953), .ZN(new_n957));
  NAND2_X1  g771(.A1(new_n956), .A2(new_n957), .ZN(G66));
  OAI21_X1  g772(.A(G953), .B1(new_n314), .B2(new_n230), .ZN(new_n959));
  NAND2_X1  g773(.A1(new_n847), .A2(new_n862), .ZN(new_n960));
  INV_X1    g774(.A(new_n960), .ZN(new_n961));
  OAI21_X1  g775(.A(new_n959), .B1(new_n961), .B2(G953), .ZN(new_n962));
  OAI21_X1  g776(.A(new_n908), .B1(G898), .B2(new_n308), .ZN(new_n963));
  XNOR2_X1  g777(.A(new_n963), .B(KEYINPUT124), .ZN(new_n964));
  XNOR2_X1  g778(.A(new_n962), .B(new_n964), .ZN(G69));
  NAND2_X1  g779(.A1(new_n552), .A2(new_n533), .ZN(new_n966));
  XNOR2_X1  g780(.A(new_n966), .B(new_n491), .ZN(new_n967));
  OAI21_X1  g781(.A(G900), .B1(new_n967), .B2(G227), .ZN(new_n968));
  AOI211_X1 g782(.A(new_n308), .B(new_n968), .C1(G227), .C2(new_n967), .ZN(new_n969));
  NAND2_X1  g783(.A1(new_n695), .A2(new_n837), .ZN(new_n970));
  INV_X1    g784(.A(KEYINPUT62), .ZN(new_n971));
  XNOR2_X1  g785(.A(new_n970), .B(new_n971), .ZN(new_n972));
  OAI21_X1  g786(.A(new_n760), .B1(new_n757), .B2(new_n848), .ZN(new_n973));
  NOR3_X1   g787(.A1(new_n973), .A2(new_n693), .A3(new_n790), .ZN(new_n974));
  XNOR2_X1  g788(.A(new_n974), .B(KEYINPUT125), .ZN(new_n975));
  AND2_X1   g789(.A1(new_n975), .A2(new_n788), .ZN(new_n976));
  NAND3_X1  g790(.A1(new_n972), .A2(new_n976), .A3(new_n797), .ZN(new_n977));
  INV_X1    g791(.A(new_n967), .ZN(new_n978));
  AOI21_X1  g792(.A(G953), .B1(new_n977), .B2(new_n978), .ZN(new_n979));
  NAND3_X1  g793(.A1(new_n775), .A2(new_n786), .A3(new_n787), .ZN(new_n980));
  NAND2_X1  g794(.A1(new_n729), .A2(new_n760), .ZN(new_n981));
  NAND2_X1  g795(.A1(new_n980), .A2(new_n981), .ZN(new_n982));
  NAND2_X1  g796(.A1(new_n982), .A2(new_n785), .ZN(new_n983));
  AND2_X1   g797(.A1(new_n797), .A2(new_n837), .ZN(new_n984));
  NAND4_X1  g798(.A1(new_n983), .A2(new_n762), .A3(new_n764), .A4(new_n984), .ZN(new_n985));
  OR2_X1    g799(.A1(new_n985), .A2(new_n978), .ZN(new_n986));
  AOI21_X1  g800(.A(new_n969), .B1(new_n979), .B2(new_n986), .ZN(G72));
  NAND2_X1  g801(.A1(G472), .A2(G902), .ZN(new_n988));
  XOR2_X1   g802(.A(new_n988), .B(KEYINPUT63), .Z(new_n989));
  OAI21_X1  g803(.A(new_n989), .B1(new_n985), .B2(new_n960), .ZN(new_n990));
  NOR2_X1   g804(.A1(new_n536), .A2(new_n520), .ZN(new_n991));
  INV_X1    g805(.A(new_n991), .ZN(new_n992));
  NOR2_X1   g806(.A1(new_n992), .A2(new_n530), .ZN(new_n993));
  AOI21_X1  g807(.A(new_n904), .B1(new_n990), .B2(new_n993), .ZN(new_n994));
  XOR2_X1   g808(.A(new_n994), .B(KEYINPUT126), .Z(new_n995));
  NAND2_X1  g809(.A1(new_n992), .A2(new_n530), .ZN(new_n996));
  NAND4_X1  g810(.A1(new_n972), .A2(new_n976), .A3(new_n797), .A4(new_n961), .ZN(new_n997));
  AOI21_X1  g811(.A(new_n996), .B1(new_n997), .B2(new_n989), .ZN(new_n998));
  INV_X1    g812(.A(new_n993), .ZN(new_n999));
  NAND3_X1  g813(.A1(new_n999), .A2(new_n989), .A3(new_n996), .ZN(new_n1000));
  XOR2_X1   g814(.A(new_n1000), .B(KEYINPUT127), .Z(new_n1001));
  NOR2_X1   g815(.A1(new_n893), .A2(new_n1001), .ZN(new_n1002));
  NOR3_X1   g816(.A1(new_n995), .A2(new_n998), .A3(new_n1002), .ZN(G57));
endmodule


