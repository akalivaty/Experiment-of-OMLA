//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 1 0 1 0 0 0 1 1 0 0 0 1 1 0 0 1 0 0 0 1 1 0 1 0 1 1 0 0 0 1 1 0 1 1 1 1 0 0 0 0 1 1 1 0 0 0 1 1 0 1 1 1 1 1 0 1 0 1 1 1 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:26:30 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n713, new_n714, new_n715, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n733,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n744, new_n745, new_n746, new_n747, new_n748, new_n749,
    new_n750, new_n751, new_n752, new_n753, new_n755, new_n756, new_n757,
    new_n758, new_n759, new_n760, new_n761, new_n762, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n775, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n806, new_n807, new_n808, new_n809, new_n810,
    new_n811, new_n812, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n948, new_n949, new_n950, new_n951, new_n952,
    new_n953, new_n954, new_n955, new_n956, new_n957, new_n958, new_n959,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n978, new_n979, new_n980, new_n981, new_n982, new_n983,
    new_n984, new_n985, new_n986, new_n988, new_n989, new_n990, new_n991,
    new_n992, new_n993, new_n994, new_n995, new_n996, new_n997, new_n999,
    new_n1000, new_n1001, new_n1002, new_n1003, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1017, new_n1018,
    new_n1019, new_n1020, new_n1021, new_n1022, new_n1023, new_n1024,
    new_n1025, new_n1026, new_n1027, new_n1028, new_n1029, new_n1030,
    new_n1031, new_n1032, new_n1033, new_n1034, new_n1036, new_n1037,
    new_n1038, new_n1039, new_n1040, new_n1041, new_n1042, new_n1043,
    new_n1044, new_n1045, new_n1046, new_n1047;
  INV_X1    g000(.A(KEYINPUT73), .ZN(new_n187));
  XNOR2_X1  g001(.A(KEYINPUT22), .B(G137), .ZN(new_n188));
  INV_X1    g002(.A(G953), .ZN(new_n189));
  AND3_X1   g003(.A1(new_n189), .A2(G221), .A3(G234), .ZN(new_n190));
  XOR2_X1   g004(.A(new_n188), .B(new_n190), .Z(new_n191));
  INV_X1    g005(.A(new_n191), .ZN(new_n192));
  INV_X1    g006(.A(KEYINPUT16), .ZN(new_n193));
  INV_X1    g007(.A(G140), .ZN(new_n194));
  NAND3_X1  g008(.A1(new_n193), .A2(new_n194), .A3(G125), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n194), .A2(G125), .ZN(new_n196));
  INV_X1    g010(.A(G125), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n197), .A2(G140), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n196), .A2(new_n198), .ZN(new_n199));
  OAI21_X1  g013(.A(new_n195), .B1(new_n199), .B2(new_n193), .ZN(new_n200));
  INV_X1    g014(.A(G146), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n200), .A2(new_n201), .ZN(new_n202));
  OAI211_X1 g016(.A(G146), .B(new_n195), .C1(new_n199), .C2(new_n193), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n202), .A2(new_n203), .ZN(new_n204));
  NAND2_X1  g018(.A1(KEYINPUT64), .A2(G128), .ZN(new_n205));
  INV_X1    g019(.A(new_n205), .ZN(new_n206));
  NOR2_X1   g020(.A1(KEYINPUT64), .A2(G128), .ZN(new_n207));
  OAI21_X1  g021(.A(G119), .B1(new_n206), .B2(new_n207), .ZN(new_n208));
  INV_X1    g022(.A(G128), .ZN(new_n209));
  NOR2_X1   g023(.A1(new_n209), .A2(G119), .ZN(new_n210));
  INV_X1    g024(.A(new_n210), .ZN(new_n211));
  NAND3_X1  g025(.A1(new_n208), .A2(KEYINPUT23), .A3(new_n211), .ZN(new_n212));
  INV_X1    g026(.A(G119), .ZN(new_n213));
  OR3_X1    g027(.A1(new_n213), .A2(KEYINPUT23), .A3(G128), .ZN(new_n214));
  NAND3_X1  g028(.A1(new_n212), .A2(G110), .A3(new_n214), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n204), .A2(new_n215), .ZN(new_n216));
  XOR2_X1   g030(.A(KEYINPUT24), .B(G110), .Z(new_n217));
  OR2_X1    g031(.A1(KEYINPUT64), .A2(G128), .ZN(new_n218));
  AOI21_X1  g032(.A(new_n213), .B1(new_n218), .B2(new_n205), .ZN(new_n219));
  NOR3_X1   g033(.A1(new_n219), .A2(KEYINPUT70), .A3(new_n210), .ZN(new_n220));
  INV_X1    g034(.A(KEYINPUT70), .ZN(new_n221));
  AOI21_X1  g035(.A(new_n221), .B1(new_n208), .B2(new_n211), .ZN(new_n222));
  OAI21_X1  g036(.A(new_n217), .B1(new_n220), .B2(new_n222), .ZN(new_n223));
  INV_X1    g037(.A(KEYINPUT71), .ZN(new_n224));
  NAND2_X1  g038(.A1(new_n223), .A2(new_n224), .ZN(new_n225));
  OAI21_X1  g039(.A(KEYINPUT70), .B1(new_n219), .B2(new_n210), .ZN(new_n226));
  NAND3_X1  g040(.A1(new_n208), .A2(new_n221), .A3(new_n211), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n226), .A2(new_n227), .ZN(new_n228));
  NAND3_X1  g042(.A1(new_n228), .A2(KEYINPUT71), .A3(new_n217), .ZN(new_n229));
  AOI21_X1  g043(.A(new_n216), .B1(new_n225), .B2(new_n229), .ZN(new_n230));
  INV_X1    g044(.A(new_n199), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n231), .A2(new_n201), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n232), .A2(new_n203), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n212), .A2(new_n214), .ZN(new_n234));
  INV_X1    g048(.A(G110), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n234), .A2(new_n235), .ZN(new_n236));
  INV_X1    g050(.A(new_n217), .ZN(new_n237));
  NAND3_X1  g051(.A1(new_n226), .A2(new_n237), .A3(new_n227), .ZN(new_n238));
  AOI21_X1  g052(.A(new_n233), .B1(new_n236), .B2(new_n238), .ZN(new_n239));
  OAI21_X1  g053(.A(new_n192), .B1(new_n230), .B2(new_n239), .ZN(new_n240));
  AOI21_X1  g054(.A(KEYINPUT71), .B1(new_n228), .B2(new_n217), .ZN(new_n241));
  AOI211_X1 g055(.A(new_n224), .B(new_n237), .C1(new_n226), .C2(new_n227), .ZN(new_n242));
  OAI211_X1 g056(.A(new_n204), .B(new_n215), .C1(new_n241), .C2(new_n242), .ZN(new_n243));
  INV_X1    g057(.A(new_n239), .ZN(new_n244));
  NAND3_X1  g058(.A1(new_n243), .A2(new_n244), .A3(new_n191), .ZN(new_n245));
  INV_X1    g059(.A(G902), .ZN(new_n246));
  NAND3_X1  g060(.A1(new_n240), .A2(new_n245), .A3(new_n246), .ZN(new_n247));
  INV_X1    g061(.A(KEYINPUT25), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n247), .A2(new_n248), .ZN(new_n249));
  NAND4_X1  g063(.A1(new_n240), .A2(new_n245), .A3(KEYINPUT25), .A4(new_n246), .ZN(new_n250));
  AND3_X1   g064(.A1(new_n249), .A2(KEYINPUT72), .A3(new_n250), .ZN(new_n251));
  INV_X1    g065(.A(KEYINPUT72), .ZN(new_n252));
  NAND3_X1  g066(.A1(new_n247), .A2(new_n252), .A3(new_n248), .ZN(new_n253));
  INV_X1    g067(.A(G217), .ZN(new_n254));
  AOI21_X1  g068(.A(new_n254), .B1(G234), .B2(new_n246), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n253), .A2(new_n255), .ZN(new_n256));
  OAI21_X1  g070(.A(new_n187), .B1(new_n251), .B2(new_n256), .ZN(new_n257));
  NAND3_X1  g071(.A1(new_n249), .A2(KEYINPUT72), .A3(new_n250), .ZN(new_n258));
  NAND4_X1  g072(.A1(new_n258), .A2(KEYINPUT73), .A3(new_n255), .A4(new_n253), .ZN(new_n259));
  NOR2_X1   g073(.A1(new_n255), .A2(G902), .ZN(new_n260));
  NAND3_X1  g074(.A1(new_n240), .A2(new_n245), .A3(new_n260), .ZN(new_n261));
  NAND3_X1  g075(.A1(new_n257), .A2(new_n259), .A3(new_n261), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n262), .A2(KEYINPUT74), .ZN(new_n263));
  INV_X1    g077(.A(KEYINPUT74), .ZN(new_n264));
  NAND4_X1  g078(.A1(new_n257), .A2(new_n264), .A3(new_n259), .A4(new_n261), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n263), .A2(new_n265), .ZN(new_n266));
  NAND2_X1  g080(.A1(new_n201), .A2(G143), .ZN(new_n267));
  INV_X1    g081(.A(G143), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n268), .A2(G146), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n267), .A2(new_n269), .ZN(new_n270));
  NAND2_X1  g084(.A1(KEYINPUT0), .A2(G128), .ZN(new_n271));
  OR2_X1    g085(.A1(KEYINPUT0), .A2(G128), .ZN(new_n272));
  NAND3_X1  g086(.A1(new_n270), .A2(new_n271), .A3(new_n272), .ZN(new_n273));
  XNOR2_X1  g087(.A(G143), .B(G146), .ZN(new_n274));
  NAND3_X1  g088(.A1(new_n274), .A2(KEYINPUT0), .A3(G128), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n273), .A2(new_n275), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n276), .A2(G125), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n218), .A2(new_n205), .ZN(new_n278));
  INV_X1    g092(.A(KEYINPUT1), .ZN(new_n279));
  AOI21_X1  g093(.A(new_n279), .B1(G143), .B2(new_n201), .ZN(new_n280));
  OAI21_X1  g094(.A(new_n270), .B1(new_n278), .B2(new_n280), .ZN(new_n281));
  NAND3_X1  g095(.A1(new_n274), .A2(new_n279), .A3(G128), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n281), .A2(new_n282), .ZN(new_n283));
  OAI21_X1  g097(.A(new_n277), .B1(G125), .B2(new_n283), .ZN(new_n284));
  AND2_X1   g098(.A1(new_n189), .A2(G224), .ZN(new_n285));
  XNOR2_X1  g099(.A(new_n284), .B(new_n285), .ZN(new_n286));
  NOR2_X1   g100(.A1(KEYINPUT2), .A2(G113), .ZN(new_n287));
  NAND2_X1  g101(.A1(KEYINPUT2), .A2(G113), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n288), .A2(KEYINPUT65), .ZN(new_n289));
  INV_X1    g103(.A(KEYINPUT65), .ZN(new_n290));
  NAND3_X1  g104(.A1(new_n290), .A2(KEYINPUT2), .A3(G113), .ZN(new_n291));
  AOI21_X1  g105(.A(new_n287), .B1(new_n289), .B2(new_n291), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n213), .A2(G116), .ZN(new_n293));
  INV_X1    g107(.A(G116), .ZN(new_n294));
  NAND2_X1  g108(.A1(new_n294), .A2(G119), .ZN(new_n295));
  NAND3_X1  g109(.A1(new_n292), .A2(new_n293), .A3(new_n295), .ZN(new_n296));
  INV_X1    g110(.A(KEYINPUT66), .ZN(new_n297));
  AND3_X1   g111(.A1(new_n293), .A2(new_n295), .A3(new_n297), .ZN(new_n298));
  AOI21_X1  g112(.A(new_n297), .B1(new_n293), .B2(new_n295), .ZN(new_n299));
  NOR2_X1   g113(.A1(new_n298), .A2(new_n299), .ZN(new_n300));
  OAI21_X1  g114(.A(new_n296), .B1(new_n300), .B2(new_n292), .ZN(new_n301));
  INV_X1    g115(.A(KEYINPUT4), .ZN(new_n302));
  INV_X1    g116(.A(G107), .ZN(new_n303));
  NOR2_X1   g117(.A1(new_n303), .A2(G104), .ZN(new_n304));
  INV_X1    g118(.A(KEYINPUT3), .ZN(new_n305));
  INV_X1    g119(.A(G104), .ZN(new_n306));
  OAI21_X1  g120(.A(new_n305), .B1(new_n306), .B2(G107), .ZN(new_n307));
  NAND3_X1  g121(.A1(new_n303), .A2(KEYINPUT3), .A3(G104), .ZN(new_n308));
  AOI21_X1  g122(.A(new_n304), .B1(new_n307), .B2(new_n308), .ZN(new_n309));
  INV_X1    g123(.A(G101), .ZN(new_n310));
  AOI21_X1  g124(.A(new_n302), .B1(new_n309), .B2(new_n310), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n306), .A2(G107), .ZN(new_n312));
  AND3_X1   g126(.A1(new_n303), .A2(KEYINPUT3), .A3(G104), .ZN(new_n313));
  AOI21_X1  g127(.A(KEYINPUT3), .B1(new_n303), .B2(G104), .ZN(new_n314));
  OAI21_X1  g128(.A(new_n312), .B1(new_n313), .B2(new_n314), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n315), .A2(G101), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n311), .A2(new_n316), .ZN(new_n317));
  NAND3_X1  g131(.A1(new_n315), .A2(new_n302), .A3(G101), .ZN(new_n318));
  NAND3_X1  g132(.A1(new_n301), .A2(new_n317), .A3(new_n318), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n303), .A2(G104), .ZN(new_n320));
  AOI21_X1  g134(.A(new_n310), .B1(new_n312), .B2(new_n320), .ZN(new_n321));
  AOI21_X1  g135(.A(new_n321), .B1(new_n309), .B2(new_n310), .ZN(new_n322));
  INV_X1    g136(.A(KEYINPUT5), .ZN(new_n323));
  NOR3_X1   g137(.A1(new_n298), .A2(new_n299), .A3(new_n323), .ZN(new_n324));
  OAI21_X1  g138(.A(G113), .B1(new_n293), .B2(KEYINPUT5), .ZN(new_n325));
  OAI211_X1 g139(.A(new_n296), .B(new_n322), .C1(new_n324), .C2(new_n325), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n319), .A2(new_n326), .ZN(new_n327));
  XNOR2_X1  g141(.A(G110), .B(G122), .ZN(new_n328));
  INV_X1    g142(.A(new_n328), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n327), .A2(new_n329), .ZN(new_n330));
  INV_X1    g144(.A(KEYINPUT81), .ZN(new_n331));
  NOR2_X1   g145(.A1(new_n330), .A2(new_n331), .ZN(new_n332));
  NAND3_X1  g146(.A1(new_n319), .A2(new_n326), .A3(new_n328), .ZN(new_n333));
  INV_X1    g147(.A(KEYINPUT80), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n333), .A2(new_n334), .ZN(new_n335));
  NAND4_X1  g149(.A1(new_n319), .A2(new_n326), .A3(KEYINPUT80), .A4(new_n328), .ZN(new_n336));
  NAND3_X1  g150(.A1(new_n335), .A2(new_n330), .A3(new_n336), .ZN(new_n337));
  AOI21_X1  g151(.A(new_n332), .B1(new_n337), .B2(KEYINPUT6), .ZN(new_n338));
  INV_X1    g152(.A(KEYINPUT6), .ZN(new_n339));
  NOR3_X1   g153(.A1(new_n330), .A2(new_n331), .A3(new_n339), .ZN(new_n340));
  OAI21_X1  g154(.A(new_n286), .B1(new_n338), .B2(new_n340), .ZN(new_n341));
  XOR2_X1   g155(.A(new_n328), .B(KEYINPUT8), .Z(new_n342));
  AND3_X1   g156(.A1(new_n293), .A2(new_n295), .A3(KEYINPUT5), .ZN(new_n343));
  OAI21_X1  g157(.A(new_n296), .B1(new_n325), .B2(new_n343), .ZN(new_n344));
  AOI21_X1  g158(.A(new_n342), .B1(new_n344), .B2(new_n322), .ZN(new_n345));
  OAI21_X1  g159(.A(new_n296), .B1(new_n324), .B2(new_n325), .ZN(new_n346));
  OAI21_X1  g160(.A(new_n345), .B1(new_n346), .B2(new_n322), .ZN(new_n347));
  OR2_X1    g161(.A1(new_n284), .A2(new_n285), .ZN(new_n348));
  INV_X1    g162(.A(KEYINPUT7), .ZN(new_n349));
  OAI21_X1  g163(.A(new_n347), .B1(new_n348), .B2(new_n349), .ZN(new_n350));
  OAI21_X1  g164(.A(new_n284), .B1(new_n349), .B2(new_n285), .ZN(new_n351));
  AND2_X1   g165(.A1(new_n351), .A2(KEYINPUT82), .ZN(new_n352));
  NOR2_X1   g166(.A1(new_n351), .A2(KEYINPUT82), .ZN(new_n353));
  NOR3_X1   g167(.A1(new_n350), .A2(new_n352), .A3(new_n353), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n335), .A2(new_n336), .ZN(new_n355));
  AOI21_X1  g169(.A(G902), .B1(new_n354), .B2(new_n355), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n341), .A2(new_n356), .ZN(new_n357));
  OAI21_X1  g171(.A(G210), .B1(G237), .B2(G902), .ZN(new_n358));
  INV_X1    g172(.A(new_n358), .ZN(new_n359));
  NAND2_X1  g173(.A1(new_n357), .A2(new_n359), .ZN(new_n360));
  NAND3_X1  g174(.A1(new_n341), .A2(new_n358), .A3(new_n356), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n360), .A2(new_n361), .ZN(new_n362));
  OAI21_X1  g176(.A(G214), .B1(G237), .B2(G902), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n362), .A2(new_n363), .ZN(new_n364));
  INV_X1    g178(.A(KEYINPUT89), .ZN(new_n365));
  OAI21_X1  g179(.A(KEYINPUT85), .B1(new_n209), .B2(G143), .ZN(new_n366));
  INV_X1    g180(.A(KEYINPUT85), .ZN(new_n367));
  NAND3_X1  g181(.A1(new_n367), .A2(new_n268), .A3(G128), .ZN(new_n368));
  NAND3_X1  g182(.A1(new_n366), .A2(new_n368), .A3(KEYINPUT13), .ZN(new_n369));
  XOR2_X1   g183(.A(new_n369), .B(KEYINPUT87), .Z(new_n370));
  NAND2_X1  g184(.A1(new_n278), .A2(G143), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n371), .A2(KEYINPUT86), .ZN(new_n372));
  INV_X1    g186(.A(KEYINPUT86), .ZN(new_n373));
  NAND3_X1  g187(.A1(new_n278), .A2(new_n373), .A3(G143), .ZN(new_n374));
  INV_X1    g188(.A(KEYINPUT13), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n366), .A2(new_n368), .ZN(new_n376));
  AOI22_X1  g190(.A1(new_n372), .A2(new_n374), .B1(new_n375), .B2(new_n376), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n370), .A2(new_n377), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n378), .A2(G134), .ZN(new_n379));
  XOR2_X1   g193(.A(G116), .B(G122), .Z(new_n380));
  XNOR2_X1  g194(.A(new_n380), .B(new_n303), .ZN(new_n381));
  AOI22_X1  g195(.A1(new_n372), .A2(new_n374), .B1(new_n368), .B2(new_n366), .ZN(new_n382));
  INV_X1    g196(.A(G134), .ZN(new_n383));
  AOI21_X1  g197(.A(new_n381), .B1(new_n382), .B2(new_n383), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n379), .A2(new_n384), .ZN(new_n385));
  OR2_X1    g199(.A1(new_n294), .A2(G122), .ZN(new_n386));
  AOI21_X1  g200(.A(new_n303), .B1(new_n386), .B2(KEYINPUT14), .ZN(new_n387));
  XOR2_X1   g201(.A(new_n387), .B(new_n380), .Z(new_n388));
  NAND2_X1  g202(.A1(new_n372), .A2(new_n374), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n389), .A2(new_n376), .ZN(new_n390));
  NOR2_X1   g204(.A1(new_n390), .A2(G134), .ZN(new_n391));
  NOR2_X1   g205(.A1(new_n382), .A2(new_n383), .ZN(new_n392));
  OAI21_X1  g206(.A(new_n388), .B1(new_n391), .B2(new_n392), .ZN(new_n393));
  XOR2_X1   g207(.A(KEYINPUT9), .B(G234), .Z(new_n394));
  NAND3_X1  g208(.A1(new_n394), .A2(G217), .A3(new_n189), .ZN(new_n395));
  INV_X1    g209(.A(new_n395), .ZN(new_n396));
  AND3_X1   g210(.A1(new_n385), .A2(new_n393), .A3(new_n396), .ZN(new_n397));
  AOI21_X1  g211(.A(new_n396), .B1(new_n385), .B2(new_n393), .ZN(new_n398));
  OAI211_X1 g212(.A(KEYINPUT88), .B(new_n246), .C1(new_n397), .C2(new_n398), .ZN(new_n399));
  INV_X1    g213(.A(G478), .ZN(new_n400));
  NOR2_X1   g214(.A1(new_n400), .A2(KEYINPUT15), .ZN(new_n401));
  AND2_X1   g215(.A1(new_n399), .A2(new_n401), .ZN(new_n402));
  NOR2_X1   g216(.A1(new_n399), .A2(new_n401), .ZN(new_n403));
  OAI21_X1  g217(.A(new_n365), .B1(new_n402), .B2(new_n403), .ZN(new_n404));
  INV_X1    g218(.A(G475), .ZN(new_n405));
  INV_X1    g219(.A(G237), .ZN(new_n406));
  NAND3_X1  g220(.A1(new_n406), .A2(new_n189), .A3(G214), .ZN(new_n407));
  XNOR2_X1  g221(.A(new_n407), .B(G143), .ZN(new_n408));
  INV_X1    g222(.A(KEYINPUT18), .ZN(new_n409));
  INV_X1    g223(.A(G131), .ZN(new_n410));
  OAI21_X1  g224(.A(new_n408), .B1(new_n409), .B2(new_n410), .ZN(new_n411));
  XNOR2_X1  g225(.A(new_n407), .B(new_n268), .ZN(new_n412));
  NAND3_X1  g226(.A1(new_n412), .A2(KEYINPUT18), .A3(G131), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n199), .A2(G146), .ZN(new_n414));
  NAND2_X1  g228(.A1(new_n232), .A2(new_n414), .ZN(new_n415));
  NAND3_X1  g229(.A1(new_n411), .A2(new_n413), .A3(new_n415), .ZN(new_n416));
  INV_X1    g230(.A(new_n416), .ZN(new_n417));
  NAND2_X1  g231(.A1(new_n412), .A2(G131), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n408), .A2(new_n410), .ZN(new_n419));
  INV_X1    g233(.A(KEYINPUT17), .ZN(new_n420));
  AND3_X1   g234(.A1(new_n418), .A2(new_n419), .A3(new_n420), .ZN(new_n421));
  INV_X1    g235(.A(new_n421), .ZN(new_n422));
  OAI211_X1 g236(.A(new_n202), .B(new_n203), .C1(new_n418), .C2(new_n420), .ZN(new_n423));
  INV_X1    g237(.A(new_n423), .ZN(new_n424));
  AOI21_X1  g238(.A(new_n417), .B1(new_n422), .B2(new_n424), .ZN(new_n425));
  XNOR2_X1  g239(.A(G113), .B(G122), .ZN(new_n426));
  XNOR2_X1  g240(.A(new_n426), .B(new_n306), .ZN(new_n427));
  XNOR2_X1  g241(.A(new_n425), .B(new_n427), .ZN(new_n428));
  AOI21_X1  g242(.A(new_n405), .B1(new_n428), .B2(new_n246), .ZN(new_n429));
  NOR2_X1   g243(.A1(G475), .A2(G902), .ZN(new_n430));
  INV_X1    g244(.A(new_n430), .ZN(new_n431));
  AND2_X1   g245(.A1(new_n418), .A2(new_n419), .ZN(new_n432));
  OR2_X1    g246(.A1(new_n199), .A2(KEYINPUT19), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n199), .A2(KEYINPUT19), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n433), .A2(new_n434), .ZN(new_n435));
  OAI21_X1  g249(.A(new_n203), .B1(new_n435), .B2(G146), .ZN(new_n436));
  OAI21_X1  g250(.A(new_n416), .B1(new_n432), .B2(new_n436), .ZN(new_n437));
  INV_X1    g251(.A(new_n427), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n437), .A2(new_n438), .ZN(new_n439));
  OAI211_X1 g253(.A(new_n427), .B(new_n416), .C1(new_n421), .C2(new_n423), .ZN(new_n440));
  AOI211_X1 g254(.A(KEYINPUT20), .B(new_n431), .C1(new_n439), .C2(new_n440), .ZN(new_n441));
  INV_X1    g255(.A(KEYINPUT84), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n439), .A2(new_n440), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n443), .A2(new_n430), .ZN(new_n444));
  XOR2_X1   g258(.A(KEYINPUT83), .B(KEYINPUT20), .Z(new_n445));
  AOI22_X1  g259(.A1(new_n441), .A2(new_n442), .B1(new_n444), .B2(new_n445), .ZN(new_n446));
  OAI21_X1  g260(.A(KEYINPUT84), .B1(new_n444), .B2(KEYINPUT20), .ZN(new_n447));
  AOI21_X1  g261(.A(new_n429), .B1(new_n446), .B2(new_n447), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n399), .A2(new_n401), .ZN(new_n449));
  AOI21_X1  g263(.A(new_n383), .B1(new_n370), .B2(new_n377), .ZN(new_n450));
  NOR3_X1   g264(.A1(new_n450), .A2(new_n391), .A3(new_n381), .ZN(new_n451));
  INV_X1    g265(.A(new_n388), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n390), .A2(G134), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n382), .A2(new_n383), .ZN(new_n454));
  AOI21_X1  g268(.A(new_n452), .B1(new_n453), .B2(new_n454), .ZN(new_n455));
  OAI21_X1  g269(.A(new_n395), .B1(new_n451), .B2(new_n455), .ZN(new_n456));
  NAND3_X1  g270(.A1(new_n385), .A2(new_n393), .A3(new_n396), .ZN(new_n457));
  NAND2_X1  g271(.A1(new_n456), .A2(new_n457), .ZN(new_n458));
  INV_X1    g272(.A(new_n401), .ZN(new_n459));
  NAND4_X1  g273(.A1(new_n458), .A2(KEYINPUT88), .A3(new_n246), .A4(new_n459), .ZN(new_n460));
  NAND3_X1  g274(.A1(new_n449), .A2(new_n460), .A3(KEYINPUT89), .ZN(new_n461));
  INV_X1    g275(.A(G952), .ZN(new_n462));
  AOI211_X1 g276(.A(G953), .B(new_n462), .C1(G234), .C2(G237), .ZN(new_n463));
  XOR2_X1   g277(.A(KEYINPUT21), .B(G898), .Z(new_n464));
  INV_X1    g278(.A(new_n464), .ZN(new_n465));
  AOI211_X1 g279(.A(new_n246), .B(new_n189), .C1(G234), .C2(G237), .ZN(new_n466));
  AOI21_X1  g280(.A(new_n463), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  INV_X1    g281(.A(new_n467), .ZN(new_n468));
  NAND4_X1  g282(.A1(new_n404), .A2(new_n448), .A3(new_n461), .A4(new_n468), .ZN(new_n469));
  NOR2_X1   g283(.A1(new_n364), .A2(new_n469), .ZN(new_n470));
  INV_X1    g284(.A(new_n276), .ZN(new_n471));
  INV_X1    g285(.A(KEYINPUT11), .ZN(new_n472));
  OAI21_X1  g286(.A(new_n472), .B1(new_n383), .B2(G137), .ZN(new_n473));
  INV_X1    g287(.A(G137), .ZN(new_n474));
  NAND3_X1  g288(.A1(new_n474), .A2(KEYINPUT11), .A3(G134), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n383), .A2(G137), .ZN(new_n476));
  NAND3_X1  g290(.A1(new_n473), .A2(new_n475), .A3(new_n476), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n477), .A2(G131), .ZN(new_n478));
  NAND4_X1  g292(.A1(new_n473), .A2(new_n475), .A3(new_n410), .A4(new_n476), .ZN(new_n479));
  AND3_X1   g293(.A1(new_n478), .A2(KEYINPUT67), .A3(new_n479), .ZN(new_n480));
  AOI21_X1  g294(.A(KEYINPUT67), .B1(new_n478), .B2(new_n479), .ZN(new_n481));
  OAI21_X1  g295(.A(new_n471), .B1(new_n480), .B2(new_n481), .ZN(new_n482));
  INV_X1    g296(.A(new_n476), .ZN(new_n483));
  NOR2_X1   g297(.A1(new_n383), .A2(G137), .ZN(new_n484));
  OAI21_X1  g298(.A(G131), .B1(new_n483), .B2(new_n484), .ZN(new_n485));
  NAND3_X1  g299(.A1(new_n283), .A2(new_n479), .A3(new_n485), .ZN(new_n486));
  AND2_X1   g300(.A1(new_n482), .A2(new_n486), .ZN(new_n487));
  INV_X1    g301(.A(new_n301), .ZN(new_n488));
  NAND3_X1  g302(.A1(new_n487), .A2(KEYINPUT28), .A3(new_n488), .ZN(new_n489));
  NAND3_X1  g303(.A1(new_n482), .A2(new_n488), .A3(new_n486), .ZN(new_n490));
  INV_X1    g304(.A(KEYINPUT28), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  AND2_X1   g306(.A1(new_n489), .A2(new_n492), .ZN(new_n493));
  NAND3_X1  g307(.A1(new_n406), .A2(new_n189), .A3(G210), .ZN(new_n494));
  XNOR2_X1  g308(.A(new_n494), .B(G101), .ZN(new_n495));
  XNOR2_X1  g309(.A(KEYINPUT26), .B(KEYINPUT27), .ZN(new_n496));
  XNOR2_X1  g310(.A(new_n495), .B(new_n496), .ZN(new_n497));
  NOR2_X1   g311(.A1(new_n487), .A2(new_n488), .ZN(new_n498));
  INV_X1    g312(.A(new_n498), .ZN(new_n499));
  NAND4_X1  g313(.A1(new_n493), .A2(KEYINPUT29), .A3(new_n497), .A4(new_n499), .ZN(new_n500));
  AOI21_X1  g314(.A(G902), .B1(new_n500), .B2(KEYINPUT69), .ZN(new_n501));
  OAI21_X1  g315(.A(new_n501), .B1(KEYINPUT69), .B2(new_n500), .ZN(new_n502));
  NAND3_X1  g316(.A1(new_n482), .A2(KEYINPUT30), .A3(new_n486), .ZN(new_n503));
  AND2_X1   g317(.A1(new_n478), .A2(new_n479), .ZN(new_n504));
  OAI21_X1  g318(.A(new_n486), .B1(new_n504), .B2(new_n276), .ZN(new_n505));
  INV_X1    g319(.A(KEYINPUT30), .ZN(new_n506));
  NAND2_X1  g320(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  NAND3_X1  g321(.A1(new_n503), .A2(new_n507), .A3(new_n301), .ZN(new_n508));
  AND2_X1   g322(.A1(new_n508), .A2(new_n490), .ZN(new_n509));
  INV_X1    g323(.A(new_n497), .ZN(new_n510));
  NAND2_X1  g324(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n505), .A2(new_n301), .ZN(new_n512));
  NAND3_X1  g326(.A1(new_n489), .A2(new_n512), .A3(new_n492), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n513), .A2(new_n497), .ZN(new_n514));
  AOI21_X1  g328(.A(KEYINPUT29), .B1(new_n511), .B2(new_n514), .ZN(new_n515));
  OAI21_X1  g329(.A(G472), .B1(new_n502), .B2(new_n515), .ZN(new_n516));
  NAND3_X1  g330(.A1(new_n508), .A2(new_n490), .A3(new_n497), .ZN(new_n517));
  INV_X1    g331(.A(KEYINPUT31), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  NAND4_X1  g333(.A1(new_n508), .A2(KEYINPUT31), .A3(new_n490), .A4(new_n497), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n513), .A2(new_n510), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  INV_X1    g337(.A(KEYINPUT68), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  NAND3_X1  g339(.A1(new_n521), .A2(new_n522), .A3(KEYINPUT68), .ZN(new_n526));
  NOR2_X1   g340(.A1(G472), .A2(G902), .ZN(new_n527));
  NAND3_X1  g341(.A1(new_n525), .A2(new_n526), .A3(new_n527), .ZN(new_n528));
  INV_X1    g342(.A(KEYINPUT32), .ZN(new_n529));
  NAND2_X1  g343(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  NAND4_X1  g344(.A1(new_n525), .A2(KEYINPUT32), .A3(new_n526), .A4(new_n527), .ZN(new_n531));
  NAND3_X1  g345(.A1(new_n516), .A2(new_n530), .A3(new_n531), .ZN(new_n532));
  INV_X1    g346(.A(G221), .ZN(new_n533));
  AOI21_X1  g347(.A(new_n533), .B1(new_n394), .B2(new_n246), .ZN(new_n534));
  INV_X1    g348(.A(G469), .ZN(new_n535));
  INV_X1    g349(.A(KEYINPUT10), .ZN(new_n536));
  AND4_X1   g350(.A1(new_n279), .A2(new_n267), .A3(new_n269), .A4(G128), .ZN(new_n537));
  OAI21_X1  g351(.A(KEYINPUT1), .B1(new_n268), .B2(G146), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n538), .A2(KEYINPUT76), .ZN(new_n539));
  INV_X1    g353(.A(KEYINPUT76), .ZN(new_n540));
  OAI211_X1 g354(.A(new_n540), .B(KEYINPUT1), .C1(new_n268), .C2(G146), .ZN(new_n541));
  NAND3_X1  g355(.A1(new_n539), .A2(G128), .A3(new_n541), .ZN(new_n542));
  AOI21_X1  g356(.A(new_n537), .B1(new_n542), .B2(new_n270), .ZN(new_n543));
  OAI211_X1 g357(.A(new_n310), .B(new_n312), .C1(new_n313), .C2(new_n314), .ZN(new_n544));
  INV_X1    g358(.A(new_n321), .ZN(new_n545));
  NAND2_X1  g359(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  NOR3_X1   g360(.A1(new_n543), .A2(KEYINPUT77), .A3(new_n546), .ZN(new_n547));
  INV_X1    g361(.A(KEYINPUT77), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n541), .A2(G128), .ZN(new_n549));
  AOI21_X1  g363(.A(new_n540), .B1(new_n267), .B2(KEYINPUT1), .ZN(new_n550));
  OAI21_X1  g364(.A(new_n270), .B1(new_n549), .B2(new_n550), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n551), .A2(new_n282), .ZN(new_n552));
  AOI21_X1  g366(.A(new_n548), .B1(new_n552), .B2(new_n322), .ZN(new_n553));
  OAI21_X1  g367(.A(new_n536), .B1(new_n547), .B2(new_n553), .ZN(new_n554));
  INV_X1    g368(.A(KEYINPUT78), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  AND3_X1   g370(.A1(new_n283), .A2(KEYINPUT10), .A3(new_n322), .ZN(new_n557));
  NAND3_X1  g371(.A1(new_n317), .A2(new_n471), .A3(new_n318), .ZN(new_n558));
  INV_X1    g372(.A(KEYINPUT75), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  NAND4_X1  g374(.A1(new_n317), .A2(KEYINPUT75), .A3(new_n471), .A4(new_n318), .ZN(new_n561));
  AOI21_X1  g375(.A(new_n557), .B1(new_n560), .B2(new_n561), .ZN(new_n562));
  NOR2_X1   g376(.A1(new_n480), .A2(new_n481), .ZN(new_n563));
  OAI211_X1 g377(.A(KEYINPUT78), .B(new_n536), .C1(new_n547), .C2(new_n553), .ZN(new_n564));
  NAND4_X1  g378(.A1(new_n556), .A2(new_n562), .A3(new_n563), .A4(new_n564), .ZN(new_n565));
  XNOR2_X1  g379(.A(G110), .B(G140), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n189), .A2(G227), .ZN(new_n567));
  XNOR2_X1  g381(.A(new_n566), .B(new_n567), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n565), .A2(new_n568), .ZN(new_n569));
  INV_X1    g383(.A(KEYINPUT79), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n569), .A2(new_n570), .ZN(new_n571));
  NAND3_X1  g385(.A1(new_n565), .A2(KEYINPUT79), .A3(new_n568), .ZN(new_n572));
  INV_X1    g386(.A(KEYINPUT12), .ZN(new_n573));
  NOR2_X1   g387(.A1(new_n283), .A2(new_n322), .ZN(new_n574));
  OAI21_X1  g388(.A(KEYINPUT77), .B1(new_n543), .B2(new_n546), .ZN(new_n575));
  NAND3_X1  g389(.A1(new_n552), .A2(new_n548), .A3(new_n322), .ZN(new_n576));
  AOI21_X1  g390(.A(new_n574), .B1(new_n575), .B2(new_n576), .ZN(new_n577));
  OAI21_X1  g391(.A(new_n573), .B1(new_n577), .B2(new_n563), .ZN(new_n578));
  NOR2_X1   g392(.A1(new_n504), .A2(new_n573), .ZN(new_n579));
  NOR2_X1   g393(.A1(new_n547), .A2(new_n553), .ZN(new_n580));
  OAI21_X1  g394(.A(new_n579), .B1(new_n580), .B2(new_n574), .ZN(new_n581));
  NAND2_X1  g395(.A1(new_n578), .A2(new_n581), .ZN(new_n582));
  AND3_X1   g396(.A1(new_n571), .A2(new_n572), .A3(new_n582), .ZN(new_n583));
  NAND3_X1  g397(.A1(new_n556), .A2(new_n564), .A3(new_n562), .ZN(new_n584));
  INV_X1    g398(.A(new_n563), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n584), .A2(new_n585), .ZN(new_n586));
  AOI21_X1  g400(.A(new_n568), .B1(new_n586), .B2(new_n565), .ZN(new_n587));
  OAI211_X1 g401(.A(new_n535), .B(new_n246), .C1(new_n583), .C2(new_n587), .ZN(new_n588));
  NOR2_X1   g402(.A1(new_n535), .A2(new_n246), .ZN(new_n589));
  NAND3_X1  g403(.A1(new_n586), .A2(new_n565), .A3(new_n568), .ZN(new_n590));
  NAND2_X1  g404(.A1(new_n565), .A2(new_n582), .ZN(new_n591));
  INV_X1    g405(.A(new_n568), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  NAND2_X1  g407(.A1(new_n590), .A2(new_n593), .ZN(new_n594));
  INV_X1    g408(.A(new_n594), .ZN(new_n595));
  AOI21_X1  g409(.A(new_n589), .B1(new_n595), .B2(G469), .ZN(new_n596));
  AOI21_X1  g410(.A(new_n534), .B1(new_n588), .B2(new_n596), .ZN(new_n597));
  NAND4_X1  g411(.A1(new_n266), .A2(new_n470), .A3(new_n532), .A4(new_n597), .ZN(new_n598));
  XNOR2_X1  g412(.A(new_n598), .B(G101), .ZN(G3));
  INV_X1    g413(.A(KEYINPUT91), .ZN(new_n600));
  NAND3_X1  g414(.A1(new_n525), .A2(new_n246), .A3(new_n526), .ZN(new_n601));
  INV_X1    g415(.A(KEYINPUT90), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n601), .A2(new_n602), .ZN(new_n603));
  NAND4_X1  g417(.A1(new_n525), .A2(KEYINPUT90), .A3(new_n246), .A4(new_n526), .ZN(new_n604));
  NAND3_X1  g418(.A1(new_n603), .A2(G472), .A3(new_n604), .ZN(new_n605));
  AOI21_X1  g419(.A(new_n600), .B1(new_n605), .B2(new_n528), .ZN(new_n606));
  NAND2_X1  g420(.A1(new_n588), .A2(new_n596), .ZN(new_n607));
  INV_X1    g421(.A(new_n534), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  INV_X1    g423(.A(G472), .ZN(new_n610));
  AOI21_X1  g424(.A(new_n610), .B1(new_n601), .B2(new_n602), .ZN(new_n611));
  AOI21_X1  g425(.A(KEYINPUT91), .B1(new_n611), .B2(new_n604), .ZN(new_n612));
  NOR3_X1   g426(.A1(new_n606), .A2(new_n609), .A3(new_n612), .ZN(new_n613));
  INV_X1    g427(.A(KEYINPUT92), .ZN(new_n614));
  NAND3_X1  g428(.A1(new_n360), .A2(new_n614), .A3(new_n361), .ZN(new_n615));
  NAND4_X1  g429(.A1(new_n341), .A2(new_n356), .A3(KEYINPUT92), .A4(new_n358), .ZN(new_n616));
  NAND2_X1  g430(.A1(new_n616), .A2(new_n363), .ZN(new_n617));
  INV_X1    g431(.A(new_n617), .ZN(new_n618));
  NAND2_X1  g432(.A1(new_n615), .A2(new_n618), .ZN(new_n619));
  NOR2_X1   g433(.A1(new_n425), .A2(new_n427), .ZN(new_n620));
  INV_X1    g434(.A(new_n440), .ZN(new_n621));
  OAI21_X1  g435(.A(new_n246), .B1(new_n620), .B2(new_n621), .ZN(new_n622));
  NAND2_X1  g436(.A1(new_n622), .A2(G475), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n444), .A2(new_n445), .ZN(new_n624));
  INV_X1    g438(.A(KEYINPUT20), .ZN(new_n625));
  NAND4_X1  g439(.A1(new_n443), .A2(new_n442), .A3(new_n625), .A4(new_n430), .ZN(new_n626));
  NAND2_X1  g440(.A1(new_n624), .A2(new_n626), .ZN(new_n627));
  NOR2_X1   g441(.A1(new_n441), .A2(new_n442), .ZN(new_n628));
  OAI21_X1  g442(.A(new_n623), .B1(new_n627), .B2(new_n628), .ZN(new_n629));
  INV_X1    g443(.A(KEYINPUT33), .ZN(new_n630));
  AOI21_X1  g444(.A(new_n630), .B1(new_n395), .B2(KEYINPUT93), .ZN(new_n631));
  INV_X1    g445(.A(new_n631), .ZN(new_n632));
  OAI21_X1  g446(.A(new_n632), .B1(new_n397), .B2(new_n398), .ZN(new_n633));
  NAND3_X1  g447(.A1(new_n456), .A2(new_n457), .A3(new_n631), .ZN(new_n634));
  NOR2_X1   g448(.A1(new_n400), .A2(G902), .ZN(new_n635));
  NAND3_X1  g449(.A1(new_n633), .A2(new_n634), .A3(new_n635), .ZN(new_n636));
  OAI21_X1  g450(.A(new_n246), .B1(new_n397), .B2(new_n398), .ZN(new_n637));
  NAND2_X1  g451(.A1(new_n637), .A2(new_n400), .ZN(new_n638));
  NAND2_X1  g452(.A1(new_n636), .A2(new_n638), .ZN(new_n639));
  NAND2_X1  g453(.A1(new_n629), .A2(new_n639), .ZN(new_n640));
  NOR3_X1   g454(.A1(new_n619), .A2(new_n467), .A3(new_n640), .ZN(new_n641));
  NAND3_X1  g455(.A1(new_n613), .A2(new_n266), .A3(new_n641), .ZN(new_n642));
  XNOR2_X1  g456(.A(new_n642), .B(KEYINPUT94), .ZN(new_n643));
  XNOR2_X1  g457(.A(KEYINPUT34), .B(G104), .ZN(new_n644));
  XNOR2_X1  g458(.A(new_n643), .B(new_n644), .ZN(G6));
  AND3_X1   g459(.A1(new_n341), .A2(new_n358), .A3(new_n356), .ZN(new_n646));
  AOI21_X1  g460(.A(new_n358), .B1(new_n341), .B2(new_n356), .ZN(new_n647));
  NOR2_X1   g461(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  AOI21_X1  g462(.A(new_n617), .B1(new_n648), .B2(new_n614), .ZN(new_n649));
  OR2_X1    g463(.A1(new_n444), .A2(new_n445), .ZN(new_n650));
  AOI21_X1  g464(.A(new_n429), .B1(new_n624), .B2(new_n650), .ZN(new_n651));
  INV_X1    g465(.A(new_n651), .ZN(new_n652));
  AOI21_X1  g466(.A(new_n652), .B1(new_n404), .B2(new_n461), .ZN(new_n653));
  AND3_X1   g467(.A1(new_n649), .A2(new_n653), .A3(new_n468), .ZN(new_n654));
  NAND3_X1  g468(.A1(new_n613), .A2(new_n266), .A3(new_n654), .ZN(new_n655));
  XOR2_X1   g469(.A(KEYINPUT35), .B(G107), .Z(new_n656));
  XNOR2_X1  g470(.A(new_n655), .B(new_n656), .ZN(G9));
  NAND2_X1  g471(.A1(new_n605), .A2(new_n600), .ZN(new_n658));
  INV_X1    g472(.A(new_n528), .ZN(new_n659));
  AOI21_X1  g473(.A(new_n659), .B1(new_n611), .B2(new_n604), .ZN(new_n660));
  OAI211_X1 g474(.A(new_n658), .B(new_n597), .C1(new_n660), .C2(new_n600), .ZN(new_n661));
  NAND2_X1  g475(.A1(new_n243), .A2(new_n244), .ZN(new_n662));
  OR2_X1    g476(.A1(new_n192), .A2(KEYINPUT36), .ZN(new_n663));
  OR2_X1    g477(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  NAND2_X1  g478(.A1(new_n662), .A2(new_n663), .ZN(new_n665));
  NAND3_X1  g479(.A1(new_n664), .A2(new_n260), .A3(new_n665), .ZN(new_n666));
  XNOR2_X1  g480(.A(new_n666), .B(KEYINPUT95), .ZN(new_n667));
  NAND3_X1  g481(.A1(new_n257), .A2(new_n259), .A3(new_n667), .ZN(new_n668));
  NAND2_X1  g482(.A1(new_n668), .A2(KEYINPUT96), .ZN(new_n669));
  INV_X1    g483(.A(KEYINPUT96), .ZN(new_n670));
  NAND4_X1  g484(.A1(new_n257), .A2(new_n670), .A3(new_n259), .A4(new_n667), .ZN(new_n671));
  NAND2_X1  g485(.A1(new_n669), .A2(new_n671), .ZN(new_n672));
  NAND2_X1  g486(.A1(new_n672), .A2(new_n470), .ZN(new_n673));
  NOR2_X1   g487(.A1(new_n661), .A2(new_n673), .ZN(new_n674));
  XNOR2_X1  g488(.A(KEYINPUT37), .B(G110), .ZN(new_n675));
  XNOR2_X1  g489(.A(new_n674), .B(new_n675), .ZN(G12));
  NOR2_X1   g490(.A1(new_n609), .A2(new_n619), .ZN(new_n677));
  INV_X1    g491(.A(G900), .ZN(new_n678));
  NAND2_X1  g492(.A1(new_n466), .A2(new_n678), .ZN(new_n679));
  INV_X1    g493(.A(new_n463), .ZN(new_n680));
  NAND2_X1  g494(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  AND3_X1   g495(.A1(new_n449), .A2(KEYINPUT89), .A3(new_n460), .ZN(new_n682));
  AOI21_X1  g496(.A(KEYINPUT89), .B1(new_n449), .B2(new_n460), .ZN(new_n683));
  OAI211_X1 g497(.A(new_n651), .B(new_n681), .C1(new_n682), .C2(new_n683), .ZN(new_n684));
  XNOR2_X1  g498(.A(new_n684), .B(KEYINPUT97), .ZN(new_n685));
  NAND4_X1  g499(.A1(new_n677), .A2(new_n685), .A3(new_n532), .A4(new_n672), .ZN(new_n686));
  XNOR2_X1  g500(.A(new_n686), .B(G128), .ZN(G30));
  NOR2_X1   g501(.A1(new_n509), .A2(new_n510), .ZN(new_n688));
  NAND2_X1  g502(.A1(new_n490), .A2(new_n510), .ZN(new_n689));
  OAI21_X1  g503(.A(new_n246), .B1(new_n498), .B2(new_n689), .ZN(new_n690));
  OAI21_X1  g504(.A(G472), .B1(new_n688), .B2(new_n690), .ZN(new_n691));
  NAND3_X1  g505(.A1(new_n530), .A2(new_n531), .A3(new_n691), .ZN(new_n692));
  INV_X1    g506(.A(new_n668), .ZN(new_n693));
  NAND2_X1  g507(.A1(new_n692), .A2(new_n693), .ZN(new_n694));
  INV_X1    g508(.A(new_n694), .ZN(new_n695));
  INV_X1    g509(.A(KEYINPUT99), .ZN(new_n696));
  XNOR2_X1  g510(.A(KEYINPUT98), .B(KEYINPUT38), .ZN(new_n697));
  XNOR2_X1  g511(.A(new_n362), .B(new_n697), .ZN(new_n698));
  AOI21_X1  g512(.A(new_n448), .B1(new_n404), .B2(new_n461), .ZN(new_n699));
  INV_X1    g513(.A(new_n699), .ZN(new_n700));
  INV_X1    g514(.A(new_n363), .ZN(new_n701));
  NOR2_X1   g515(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  NAND4_X1  g516(.A1(new_n695), .A2(new_n696), .A3(new_n698), .A4(new_n702), .ZN(new_n703));
  NAND2_X1  g517(.A1(new_n702), .A2(new_n698), .ZN(new_n704));
  OAI21_X1  g518(.A(KEYINPUT99), .B1(new_n704), .B2(new_n694), .ZN(new_n705));
  XOR2_X1   g519(.A(new_n681), .B(KEYINPUT39), .Z(new_n706));
  INV_X1    g520(.A(new_n706), .ZN(new_n707));
  NAND2_X1  g521(.A1(new_n597), .A2(new_n707), .ZN(new_n708));
  INV_X1    g522(.A(KEYINPUT40), .ZN(new_n709));
  XNOR2_X1  g523(.A(new_n708), .B(new_n709), .ZN(new_n710));
  NAND3_X1  g524(.A1(new_n703), .A2(new_n705), .A3(new_n710), .ZN(new_n711));
  XNOR2_X1  g525(.A(new_n711), .B(G143), .ZN(G45));
  NAND3_X1  g526(.A1(new_n629), .A2(new_n639), .A3(new_n681), .ZN(new_n713));
  INV_X1    g527(.A(new_n713), .ZN(new_n714));
  NAND4_X1  g528(.A1(new_n677), .A2(new_n532), .A3(new_n672), .A4(new_n714), .ZN(new_n715));
  XNOR2_X1  g529(.A(new_n715), .B(G146), .ZN(G48));
  AOI22_X1  g530(.A1(new_n569), .A2(new_n570), .B1(new_n578), .B2(new_n581), .ZN(new_n717));
  AOI21_X1  g531(.A(new_n587), .B1(new_n717), .B2(new_n572), .ZN(new_n718));
  OAI21_X1  g532(.A(G469), .B1(new_n718), .B2(G902), .ZN(new_n719));
  NAND3_X1  g533(.A1(new_n719), .A2(new_n588), .A3(new_n608), .ZN(new_n720));
  INV_X1    g534(.A(KEYINPUT100), .ZN(new_n721));
  NAND2_X1  g535(.A1(new_n720), .A2(new_n721), .ZN(new_n722));
  NAND4_X1  g536(.A1(new_n719), .A2(new_n588), .A3(KEYINPUT100), .A4(new_n608), .ZN(new_n723));
  NAND2_X1  g537(.A1(new_n722), .A2(new_n723), .ZN(new_n724));
  NAND4_X1  g538(.A1(new_n724), .A2(new_n532), .A3(new_n266), .A4(new_n641), .ZN(new_n725));
  NAND2_X1  g539(.A1(new_n725), .A2(KEYINPUT101), .ZN(new_n726));
  AND2_X1   g540(.A1(new_n266), .A2(new_n532), .ZN(new_n727));
  INV_X1    g541(.A(KEYINPUT101), .ZN(new_n728));
  NAND4_X1  g542(.A1(new_n727), .A2(new_n728), .A3(new_n641), .A4(new_n724), .ZN(new_n729));
  NAND2_X1  g543(.A1(new_n726), .A2(new_n729), .ZN(new_n730));
  XNOR2_X1  g544(.A(KEYINPUT41), .B(G113), .ZN(new_n731));
  XNOR2_X1  g545(.A(new_n730), .B(new_n731), .ZN(G15));
  NAND3_X1  g546(.A1(new_n727), .A2(new_n654), .A3(new_n724), .ZN(new_n733));
  XNOR2_X1  g547(.A(new_n733), .B(G116), .ZN(G18));
  AND3_X1   g548(.A1(new_n719), .A2(new_n588), .A3(new_n608), .ZN(new_n735));
  INV_X1    g549(.A(KEYINPUT102), .ZN(new_n736));
  NAND3_X1  g550(.A1(new_n735), .A2(new_n736), .A3(new_n649), .ZN(new_n737));
  OAI21_X1  g551(.A(KEYINPUT102), .B1(new_n720), .B2(new_n619), .ZN(new_n738));
  NAND2_X1  g552(.A1(new_n737), .A2(new_n738), .ZN(new_n739));
  INV_X1    g553(.A(new_n469), .ZN(new_n740));
  AND3_X1   g554(.A1(new_n672), .A2(new_n532), .A3(new_n740), .ZN(new_n741));
  NAND2_X1  g555(.A1(new_n739), .A2(new_n741), .ZN(new_n742));
  XNOR2_X1  g556(.A(new_n742), .B(G119), .ZN(G21));
  NAND3_X1  g557(.A1(new_n649), .A2(new_n468), .A3(new_n699), .ZN(new_n744));
  AND3_X1   g558(.A1(new_n257), .A2(new_n259), .A3(new_n261), .ZN(new_n745));
  NAND2_X1  g559(.A1(new_n601), .A2(G472), .ZN(new_n746));
  XOR2_X1   g560(.A(new_n527), .B(KEYINPUT103), .Z(new_n747));
  INV_X1    g561(.A(new_n521), .ZN(new_n748));
  AOI21_X1  g562(.A(new_n497), .B1(new_n493), .B2(new_n499), .ZN(new_n749));
  OAI21_X1  g563(.A(new_n747), .B1(new_n748), .B2(new_n749), .ZN(new_n750));
  NAND3_X1  g564(.A1(new_n745), .A2(new_n746), .A3(new_n750), .ZN(new_n751));
  NOR2_X1   g565(.A1(new_n744), .A2(new_n751), .ZN(new_n752));
  NAND2_X1  g566(.A1(new_n752), .A2(new_n724), .ZN(new_n753));
  XNOR2_X1  g567(.A(new_n753), .B(G122), .ZN(G24));
  NAND3_X1  g568(.A1(new_n746), .A2(new_n668), .A3(new_n750), .ZN(new_n755));
  NAND2_X1  g569(.A1(new_n713), .A2(KEYINPUT104), .ZN(new_n756));
  INV_X1    g570(.A(KEYINPUT104), .ZN(new_n757));
  NAND4_X1  g571(.A1(new_n629), .A2(new_n639), .A3(new_n757), .A4(new_n681), .ZN(new_n758));
  AOI21_X1  g572(.A(new_n755), .B1(new_n756), .B2(new_n758), .ZN(new_n759));
  AOI21_X1  g573(.A(new_n736), .B1(new_n735), .B2(new_n649), .ZN(new_n760));
  NOR3_X1   g574(.A1(new_n720), .A2(new_n619), .A3(KEYINPUT102), .ZN(new_n761));
  OAI21_X1  g575(.A(new_n759), .B1(new_n760), .B2(new_n761), .ZN(new_n762));
  XNOR2_X1  g576(.A(new_n762), .B(G125), .ZN(G27));
  INV_X1    g577(.A(KEYINPUT42), .ZN(new_n764));
  NAND2_X1  g578(.A1(new_n756), .A2(new_n758), .ZN(new_n765));
  NAND2_X1  g579(.A1(new_n648), .A2(new_n363), .ZN(new_n766));
  NOR2_X1   g580(.A1(new_n609), .A2(new_n766), .ZN(new_n767));
  NAND4_X1  g581(.A1(new_n727), .A2(new_n764), .A3(new_n765), .A4(new_n767), .ZN(new_n768));
  NAND2_X1  g582(.A1(new_n532), .A2(new_n745), .ZN(new_n769));
  INV_X1    g583(.A(new_n766), .ZN(new_n770));
  NAND3_X1  g584(.A1(new_n770), .A2(new_n597), .A3(new_n765), .ZN(new_n771));
  OAI21_X1  g585(.A(KEYINPUT42), .B1(new_n769), .B2(new_n771), .ZN(new_n772));
  NAND2_X1  g586(.A1(new_n768), .A2(new_n772), .ZN(new_n773));
  XNOR2_X1  g587(.A(new_n773), .B(new_n410), .ZN(G33));
  NAND3_X1  g588(.A1(new_n727), .A2(new_n685), .A3(new_n767), .ZN(new_n775));
  XNOR2_X1  g589(.A(new_n775), .B(G134), .ZN(G36));
  INV_X1    g590(.A(KEYINPUT45), .ZN(new_n777));
  AOI21_X1  g591(.A(new_n535), .B1(new_n594), .B2(new_n777), .ZN(new_n778));
  NAND3_X1  g592(.A1(new_n590), .A2(new_n593), .A3(KEYINPUT45), .ZN(new_n779));
  NAND2_X1  g593(.A1(new_n779), .A2(KEYINPUT105), .ZN(new_n780));
  INV_X1    g594(.A(KEYINPUT105), .ZN(new_n781));
  NAND4_X1  g595(.A1(new_n590), .A2(new_n593), .A3(new_n781), .A4(KEYINPUT45), .ZN(new_n782));
  NAND3_X1  g596(.A1(new_n778), .A2(new_n780), .A3(new_n782), .ZN(new_n783));
  NAND2_X1  g597(.A1(new_n783), .A2(KEYINPUT106), .ZN(new_n784));
  INV_X1    g598(.A(KEYINPUT106), .ZN(new_n785));
  NAND4_X1  g599(.A1(new_n778), .A2(new_n780), .A3(new_n785), .A4(new_n782), .ZN(new_n786));
  NAND2_X1  g600(.A1(new_n784), .A2(new_n786), .ZN(new_n787));
  INV_X1    g601(.A(new_n589), .ZN(new_n788));
  NAND3_X1  g602(.A1(new_n787), .A2(KEYINPUT46), .A3(new_n788), .ZN(new_n789));
  NAND2_X1  g603(.A1(new_n789), .A2(new_n588), .ZN(new_n790));
  AOI21_X1  g604(.A(new_n589), .B1(new_n784), .B2(new_n786), .ZN(new_n791));
  NOR2_X1   g605(.A1(new_n791), .A2(KEYINPUT46), .ZN(new_n792));
  OAI21_X1  g606(.A(new_n608), .B1(new_n790), .B2(new_n792), .ZN(new_n793));
  NOR2_X1   g607(.A1(new_n793), .A2(new_n706), .ZN(new_n794));
  NAND2_X1  g608(.A1(new_n448), .A2(new_n639), .ZN(new_n795));
  INV_X1    g609(.A(KEYINPUT107), .ZN(new_n796));
  NOR2_X1   g610(.A1(new_n796), .A2(KEYINPUT43), .ZN(new_n797));
  NAND2_X1  g611(.A1(new_n795), .A2(new_n797), .ZN(new_n798));
  AOI22_X1  g612(.A1(new_n448), .A2(new_n639), .B1(new_n796), .B2(KEYINPUT43), .ZN(new_n799));
  OAI21_X1  g613(.A(new_n798), .B1(new_n799), .B2(new_n797), .ZN(new_n800));
  OAI211_X1 g614(.A(new_n668), .B(new_n800), .C1(new_n606), .C2(new_n612), .ZN(new_n801));
  INV_X1    g615(.A(KEYINPUT44), .ZN(new_n802));
  AOI21_X1  g616(.A(new_n766), .B1(new_n801), .B2(new_n802), .ZN(new_n803));
  OAI211_X1 g617(.A(new_n794), .B(new_n803), .C1(new_n802), .C2(new_n801), .ZN(new_n804));
  XNOR2_X1  g618(.A(new_n804), .B(G137), .ZN(G39));
  XOR2_X1   g619(.A(KEYINPUT108), .B(KEYINPUT47), .Z(new_n806));
  INV_X1    g620(.A(new_n806), .ZN(new_n807));
  NAND2_X1  g621(.A1(new_n793), .A2(new_n807), .ZN(new_n808));
  NAND2_X1  g622(.A1(KEYINPUT108), .A2(KEYINPUT47), .ZN(new_n809));
  OAI211_X1 g623(.A(new_n608), .B(new_n809), .C1(new_n790), .C2(new_n792), .ZN(new_n810));
  NOR4_X1   g624(.A1(new_n266), .A2(new_n532), .A3(new_n713), .A4(new_n766), .ZN(new_n811));
  NAND3_X1  g625(.A1(new_n808), .A2(new_n810), .A3(new_n811), .ZN(new_n812));
  XNOR2_X1  g626(.A(new_n812), .B(G140), .ZN(G42));
  INV_X1    g627(.A(KEYINPUT54), .ZN(new_n814));
  INV_X1    g628(.A(KEYINPUT53), .ZN(new_n815));
  NAND3_X1  g629(.A1(new_n742), .A2(new_n733), .A3(new_n753), .ZN(new_n816));
  AOI21_X1  g630(.A(new_n816), .B1(new_n729), .B2(new_n726), .ZN(new_n817));
  NAND3_X1  g631(.A1(new_n768), .A2(new_n772), .A3(new_n775), .ZN(new_n818));
  AND2_X1   g632(.A1(new_n672), .A2(new_n532), .ZN(new_n819));
  NOR2_X1   g633(.A1(new_n402), .A2(new_n403), .ZN(new_n820));
  INV_X1    g634(.A(new_n681), .ZN(new_n821));
  NOR2_X1   g635(.A1(new_n652), .A2(new_n821), .ZN(new_n822));
  NAND4_X1  g636(.A1(new_n819), .A2(new_n820), .A3(new_n767), .A4(new_n822), .ZN(new_n823));
  OAI21_X1  g637(.A(KEYINPUT111), .B1(new_n771), .B2(new_n755), .ZN(new_n824));
  NAND2_X1  g638(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  NOR3_X1   g639(.A1(new_n771), .A2(KEYINPUT111), .A3(new_n755), .ZN(new_n826));
  NOR3_X1   g640(.A1(new_n818), .A2(new_n825), .A3(new_n826), .ZN(new_n827));
  INV_X1    g641(.A(new_n266), .ZN(new_n828));
  OAI21_X1  g642(.A(new_n640), .B1(new_n820), .B2(new_n629), .ZN(new_n829));
  NAND2_X1  g643(.A1(new_n829), .A2(new_n468), .ZN(new_n830));
  NOR2_X1   g644(.A1(new_n830), .A2(new_n364), .ZN(new_n831));
  INV_X1    g645(.A(new_n831), .ZN(new_n832));
  NOR3_X1   g646(.A1(new_n661), .A2(new_n828), .A3(new_n832), .ZN(new_n833));
  OAI21_X1  g647(.A(new_n598), .B1(new_n661), .B2(new_n673), .ZN(new_n834));
  NOR3_X1   g648(.A1(new_n833), .A2(new_n834), .A3(KEYINPUT110), .ZN(new_n835));
  INV_X1    g649(.A(KEYINPUT110), .ZN(new_n836));
  INV_X1    g650(.A(new_n598), .ZN(new_n837));
  INV_X1    g651(.A(new_n673), .ZN(new_n838));
  AOI21_X1  g652(.A(new_n837), .B1(new_n613), .B2(new_n838), .ZN(new_n839));
  NAND3_X1  g653(.A1(new_n613), .A2(new_n266), .A3(new_n831), .ZN(new_n840));
  AOI21_X1  g654(.A(new_n836), .B1(new_n839), .B2(new_n840), .ZN(new_n841));
  OAI211_X1 g655(.A(new_n817), .B(new_n827), .C1(new_n835), .C2(new_n841), .ZN(new_n842));
  NOR2_X1   g656(.A1(new_n609), .A2(new_n821), .ZN(new_n843));
  NOR2_X1   g657(.A1(new_n700), .A2(new_n619), .ZN(new_n844));
  NAND4_X1  g658(.A1(new_n843), .A2(new_n844), .A3(new_n693), .A4(new_n692), .ZN(new_n845));
  NAND4_X1  g659(.A1(new_n762), .A2(new_n686), .A3(new_n845), .A4(new_n715), .ZN(new_n846));
  INV_X1    g660(.A(KEYINPUT52), .ZN(new_n847));
  NAND2_X1  g661(.A1(new_n846), .A2(new_n847), .ZN(new_n848));
  OAI211_X1 g662(.A(new_n819), .B(new_n677), .C1(new_n685), .C2(new_n714), .ZN(new_n849));
  NAND4_X1  g663(.A1(new_n849), .A2(KEYINPUT52), .A3(new_n762), .A4(new_n845), .ZN(new_n850));
  NAND3_X1  g664(.A1(new_n848), .A2(KEYINPUT112), .A3(new_n850), .ZN(new_n851));
  INV_X1    g665(.A(KEYINPUT112), .ZN(new_n852));
  NAND3_X1  g666(.A1(new_n846), .A2(new_n852), .A3(new_n847), .ZN(new_n853));
  NAND2_X1  g667(.A1(new_n851), .A2(new_n853), .ZN(new_n854));
  OAI21_X1  g668(.A(new_n815), .B1(new_n842), .B2(new_n854), .ZN(new_n855));
  AND2_X1   g669(.A1(new_n733), .A2(new_n753), .ZN(new_n856));
  NAND3_X1  g670(.A1(new_n730), .A2(new_n856), .A3(new_n742), .ZN(new_n857));
  OAI21_X1  g671(.A(KEYINPUT110), .B1(new_n833), .B2(new_n834), .ZN(new_n858));
  NAND3_X1  g672(.A1(new_n839), .A2(new_n836), .A3(new_n840), .ZN(new_n859));
  AOI21_X1  g673(.A(new_n857), .B1(new_n858), .B2(new_n859), .ZN(new_n860));
  NAND2_X1  g674(.A1(new_n848), .A2(new_n850), .ZN(new_n861));
  NAND4_X1  g675(.A1(new_n860), .A2(KEYINPUT53), .A3(new_n827), .A4(new_n861), .ZN(new_n862));
  AOI21_X1  g676(.A(new_n814), .B1(new_n855), .B2(new_n862), .ZN(new_n863));
  NAND2_X1  g677(.A1(new_n859), .A2(new_n858), .ZN(new_n864));
  NAND4_X1  g678(.A1(new_n864), .A2(new_n817), .A3(new_n827), .A4(new_n861), .ZN(new_n865));
  AND2_X1   g679(.A1(new_n865), .A2(new_n815), .ZN(new_n866));
  NOR3_X1   g680(.A1(new_n842), .A2(new_n854), .A3(new_n815), .ZN(new_n867));
  NOR2_X1   g681(.A1(new_n866), .A2(new_n867), .ZN(new_n868));
  XNOR2_X1  g682(.A(KEYINPUT113), .B(KEYINPUT54), .ZN(new_n869));
  INV_X1    g683(.A(new_n869), .ZN(new_n870));
  AOI21_X1  g684(.A(new_n863), .B1(new_n868), .B2(new_n870), .ZN(new_n871));
  NOR2_X1   g685(.A1(new_n828), .A2(new_n680), .ZN(new_n872));
  AND3_X1   g686(.A1(new_n530), .A2(new_n531), .A3(new_n691), .ZN(new_n873));
  NOR2_X1   g687(.A1(new_n720), .A2(new_n766), .ZN(new_n874));
  AND3_X1   g688(.A1(new_n872), .A2(new_n873), .A3(new_n874), .ZN(new_n875));
  NOR2_X1   g689(.A1(new_n629), .A2(new_n639), .ZN(new_n876));
  NAND3_X1  g690(.A1(new_n875), .A2(KEYINPUT116), .A3(new_n876), .ZN(new_n877));
  NAND3_X1  g691(.A1(new_n874), .A2(new_n463), .A3(new_n800), .ZN(new_n878));
  NOR2_X1   g692(.A1(new_n878), .A2(new_n755), .ZN(new_n879));
  NAND4_X1  g693(.A1(new_n872), .A2(new_n873), .A3(new_n874), .A4(new_n876), .ZN(new_n880));
  INV_X1    g694(.A(KEYINPUT116), .ZN(new_n881));
  AOI21_X1  g695(.A(new_n879), .B1(new_n880), .B2(new_n881), .ZN(new_n882));
  NAND2_X1  g696(.A1(new_n877), .A2(new_n882), .ZN(new_n883));
  NOR3_X1   g697(.A1(new_n698), .A2(new_n363), .A3(new_n720), .ZN(new_n884));
  NAND2_X1  g698(.A1(new_n800), .A2(new_n463), .ZN(new_n885));
  NOR2_X1   g699(.A1(new_n885), .A2(new_n751), .ZN(new_n886));
  AOI21_X1  g700(.A(KEYINPUT50), .B1(new_n884), .B2(new_n886), .ZN(new_n887));
  INV_X1    g701(.A(new_n887), .ZN(new_n888));
  NAND3_X1  g702(.A1(new_n884), .A2(new_n886), .A3(KEYINPUT50), .ZN(new_n889));
  AOI22_X1  g703(.A1(new_n883), .A2(KEYINPUT117), .B1(new_n888), .B2(new_n889), .ZN(new_n890));
  NAND2_X1  g704(.A1(new_n886), .A2(new_n770), .ZN(new_n891));
  INV_X1    g705(.A(KEYINPUT114), .ZN(new_n892));
  XNOR2_X1  g706(.A(new_n891), .B(new_n892), .ZN(new_n893));
  INV_X1    g707(.A(new_n893), .ZN(new_n894));
  NAND2_X1  g708(.A1(new_n719), .A2(new_n588), .ZN(new_n895));
  NOR2_X1   g709(.A1(new_n895), .A2(new_n608), .ZN(new_n896));
  AOI21_X1  g710(.A(new_n896), .B1(new_n808), .B2(new_n810), .ZN(new_n897));
  OAI21_X1  g711(.A(new_n894), .B1(new_n897), .B2(KEYINPUT118), .ZN(new_n898));
  INV_X1    g712(.A(KEYINPUT118), .ZN(new_n899));
  AOI211_X1 g713(.A(new_n899), .B(new_n896), .C1(new_n808), .C2(new_n810), .ZN(new_n900));
  OAI21_X1  g714(.A(new_n890), .B1(new_n898), .B2(new_n900), .ZN(new_n901));
  INV_X1    g715(.A(new_n883), .ZN(new_n902));
  INV_X1    g716(.A(KEYINPUT51), .ZN(new_n903));
  OR2_X1    g717(.A1(new_n903), .A2(KEYINPUT117), .ZN(new_n904));
  OR2_X1    g718(.A1(new_n791), .A2(KEYINPUT46), .ZN(new_n905));
  INV_X1    g719(.A(new_n588), .ZN(new_n906));
  AOI21_X1  g720(.A(new_n906), .B1(new_n791), .B2(KEYINPUT46), .ZN(new_n907));
  AOI21_X1  g721(.A(new_n534), .B1(new_n905), .B2(new_n907), .ZN(new_n908));
  OAI21_X1  g722(.A(new_n810), .B1(new_n908), .B2(new_n806), .ZN(new_n909));
  INV_X1    g723(.A(new_n896), .ZN(new_n910));
  AOI21_X1  g724(.A(new_n893), .B1(new_n909), .B2(new_n910), .ZN(new_n911));
  NAND3_X1  g725(.A1(new_n888), .A2(new_n889), .A3(KEYINPUT115), .ZN(new_n912));
  INV_X1    g726(.A(KEYINPUT115), .ZN(new_n913));
  INV_X1    g727(.A(new_n889), .ZN(new_n914));
  OAI21_X1  g728(.A(new_n913), .B1(new_n914), .B2(new_n887), .ZN(new_n915));
  NAND3_X1  g729(.A1(new_n912), .A2(new_n915), .A3(new_n903), .ZN(new_n916));
  OAI21_X1  g730(.A(new_n904), .B1(new_n911), .B2(new_n916), .ZN(new_n917));
  AOI22_X1  g731(.A1(new_n901), .A2(KEYINPUT51), .B1(new_n902), .B2(new_n917), .ZN(new_n918));
  NOR2_X1   g732(.A1(new_n878), .A2(new_n769), .ZN(new_n919));
  XOR2_X1   g733(.A(new_n919), .B(KEYINPUT48), .Z(new_n920));
  NAND3_X1  g734(.A1(new_n875), .A2(new_n629), .A3(new_n639), .ZN(new_n921));
  AOI211_X1 g735(.A(new_n462), .B(G953), .C1(new_n739), .C2(new_n886), .ZN(new_n922));
  NAND3_X1  g736(.A1(new_n920), .A2(new_n921), .A3(new_n922), .ZN(new_n923));
  OAI21_X1  g737(.A(KEYINPUT119), .B1(new_n918), .B2(new_n923), .ZN(new_n924));
  INV_X1    g738(.A(KEYINPUT119), .ZN(new_n925));
  INV_X1    g739(.A(new_n923), .ZN(new_n926));
  AND2_X1   g740(.A1(new_n917), .A2(new_n902), .ZN(new_n927));
  NAND2_X1  g741(.A1(new_n909), .A2(new_n910), .ZN(new_n928));
  NAND2_X1  g742(.A1(new_n928), .A2(new_n899), .ZN(new_n929));
  NAND2_X1  g743(.A1(new_n897), .A2(KEYINPUT118), .ZN(new_n930));
  NAND3_X1  g744(.A1(new_n929), .A2(new_n930), .A3(new_n894), .ZN(new_n931));
  AOI21_X1  g745(.A(new_n903), .B1(new_n931), .B2(new_n890), .ZN(new_n932));
  OAI211_X1 g746(.A(new_n925), .B(new_n926), .C1(new_n927), .C2(new_n932), .ZN(new_n933));
  NAND3_X1  g747(.A1(new_n871), .A2(new_n924), .A3(new_n933), .ZN(new_n934));
  NAND2_X1  g748(.A1(new_n462), .A2(new_n189), .ZN(new_n935));
  NAND2_X1  g749(.A1(new_n934), .A2(new_n935), .ZN(new_n936));
  NOR3_X1   g750(.A1(new_n795), .A2(new_n534), .A3(new_n701), .ZN(new_n937));
  INV_X1    g751(.A(new_n895), .ZN(new_n938));
  INV_X1    g752(.A(KEYINPUT49), .ZN(new_n939));
  OAI211_X1 g753(.A(new_n745), .B(new_n937), .C1(new_n938), .C2(new_n939), .ZN(new_n940));
  INV_X1    g754(.A(KEYINPUT109), .ZN(new_n941));
  OR2_X1    g755(.A1(new_n940), .A2(new_n941), .ZN(new_n942));
  NAND2_X1  g756(.A1(new_n940), .A2(new_n941), .ZN(new_n943));
  NAND2_X1  g757(.A1(new_n938), .A2(new_n939), .ZN(new_n944));
  NOR2_X1   g758(.A1(new_n698), .A2(new_n692), .ZN(new_n945));
  NAND4_X1  g759(.A1(new_n942), .A2(new_n943), .A3(new_n944), .A4(new_n945), .ZN(new_n946));
  NAND2_X1  g760(.A1(new_n936), .A2(new_n946), .ZN(G75));
  AND2_X1   g761(.A1(new_n851), .A2(new_n853), .ZN(new_n948));
  NAND4_X1  g762(.A1(new_n948), .A2(KEYINPUT53), .A3(new_n860), .A4(new_n827), .ZN(new_n949));
  NAND2_X1  g763(.A1(new_n865), .A2(new_n815), .ZN(new_n950));
  NAND2_X1  g764(.A1(new_n949), .A2(new_n950), .ZN(new_n951));
  NAND3_X1  g765(.A1(new_n951), .A2(G210), .A3(G902), .ZN(new_n952));
  INV_X1    g766(.A(KEYINPUT56), .ZN(new_n953));
  NOR2_X1   g767(.A1(new_n338), .A2(new_n340), .ZN(new_n954));
  XNOR2_X1  g768(.A(new_n954), .B(new_n286), .ZN(new_n955));
  XNOR2_X1  g769(.A(new_n955), .B(KEYINPUT55), .ZN(new_n956));
  AND3_X1   g770(.A1(new_n952), .A2(new_n953), .A3(new_n956), .ZN(new_n957));
  AOI21_X1  g771(.A(new_n956), .B1(new_n952), .B2(new_n953), .ZN(new_n958));
  NOR2_X1   g772(.A1(new_n189), .A2(G952), .ZN(new_n959));
  NOR3_X1   g773(.A1(new_n957), .A2(new_n958), .A3(new_n959), .ZN(G51));
  XNOR2_X1  g774(.A(new_n589), .B(KEYINPUT120), .ZN(new_n961));
  XOR2_X1   g775(.A(new_n961), .B(KEYINPUT57), .Z(new_n962));
  NOR2_X1   g776(.A1(new_n951), .A2(new_n869), .ZN(new_n963));
  AOI21_X1  g777(.A(new_n870), .B1(new_n949), .B2(new_n950), .ZN(new_n964));
  OAI21_X1  g778(.A(new_n962), .B1(new_n963), .B2(new_n964), .ZN(new_n965));
  INV_X1    g779(.A(new_n718), .ZN(new_n966));
  NAND2_X1  g780(.A1(new_n965), .A2(new_n966), .ZN(new_n967));
  NAND2_X1  g781(.A1(new_n951), .A2(G902), .ZN(new_n968));
  OR2_X1    g782(.A1(new_n968), .A2(new_n787), .ZN(new_n969));
  AOI21_X1  g783(.A(new_n959), .B1(new_n967), .B2(new_n969), .ZN(G54));
  INV_X1    g784(.A(new_n443), .ZN(new_n971));
  NAND2_X1  g785(.A1(KEYINPUT58), .A2(G475), .ZN(new_n972));
  OAI21_X1  g786(.A(new_n971), .B1(new_n968), .B2(new_n972), .ZN(new_n973));
  INV_X1    g787(.A(new_n959), .ZN(new_n974));
  NAND2_X1  g788(.A1(new_n973), .A2(new_n974), .ZN(new_n975));
  NOR3_X1   g789(.A1(new_n968), .A2(new_n971), .A3(new_n972), .ZN(new_n976));
  NOR2_X1   g790(.A1(new_n975), .A2(new_n976), .ZN(G60));
  AND2_X1   g791(.A1(new_n633), .A2(new_n634), .ZN(new_n978));
  NAND2_X1  g792(.A1(G478), .A2(G902), .ZN(new_n979));
  XNOR2_X1  g793(.A(new_n979), .B(KEYINPUT59), .ZN(new_n980));
  OAI211_X1 g794(.A(new_n978), .B(new_n980), .C1(new_n963), .C2(new_n964), .ZN(new_n981));
  NAND2_X1  g795(.A1(new_n981), .A2(new_n974), .ZN(new_n982));
  NAND2_X1  g796(.A1(new_n855), .A2(new_n862), .ZN(new_n983));
  NAND2_X1  g797(.A1(new_n983), .A2(KEYINPUT54), .ZN(new_n984));
  OAI21_X1  g798(.A(new_n984), .B1(new_n869), .B2(new_n951), .ZN(new_n985));
  AOI21_X1  g799(.A(new_n978), .B1(new_n985), .B2(new_n980), .ZN(new_n986));
  NOR2_X1   g800(.A1(new_n982), .A2(new_n986), .ZN(G63));
  NAND2_X1  g801(.A1(new_n240), .A2(new_n245), .ZN(new_n988));
  NAND2_X1  g802(.A1(G217), .A2(G902), .ZN(new_n989));
  XNOR2_X1  g803(.A(new_n989), .B(KEYINPUT60), .ZN(new_n990));
  OAI21_X1  g804(.A(new_n988), .B1(new_n868), .B2(new_n990), .ZN(new_n991));
  INV_X1    g805(.A(new_n990), .ZN(new_n992));
  NAND4_X1  g806(.A1(new_n951), .A2(new_n664), .A3(new_n665), .A4(new_n992), .ZN(new_n993));
  NAND3_X1  g807(.A1(new_n991), .A2(new_n974), .A3(new_n993), .ZN(new_n994));
  INV_X1    g808(.A(KEYINPUT61), .ZN(new_n995));
  NAND2_X1  g809(.A1(new_n994), .A2(new_n995), .ZN(new_n996));
  NAND4_X1  g810(.A1(new_n991), .A2(new_n993), .A3(KEYINPUT61), .A4(new_n974), .ZN(new_n997));
  NAND2_X1  g811(.A1(new_n996), .A2(new_n997), .ZN(G66));
  AOI21_X1  g812(.A(new_n189), .B1(new_n464), .B2(G224), .ZN(new_n999));
  INV_X1    g813(.A(new_n860), .ZN(new_n1000));
  AOI21_X1  g814(.A(new_n999), .B1(new_n1000), .B2(new_n189), .ZN(new_n1001));
  XNOR2_X1  g815(.A(new_n1001), .B(KEYINPUT121), .ZN(new_n1002));
  OAI21_X1  g816(.A(new_n954), .B1(G898), .B2(new_n189), .ZN(new_n1003));
  XOR2_X1   g817(.A(new_n1002), .B(new_n1003), .Z(G69));
  NAND2_X1  g818(.A1(new_n503), .A2(new_n507), .ZN(new_n1005));
  XOR2_X1   g819(.A(new_n435), .B(KEYINPUT122), .Z(new_n1006));
  XNOR2_X1  g820(.A(new_n1005), .B(new_n1006), .ZN(new_n1007));
  NAND2_X1  g821(.A1(G900), .A2(G953), .ZN(new_n1008));
  INV_X1    g822(.A(new_n818), .ZN(new_n1009));
  AND2_X1   g823(.A1(new_n849), .A2(new_n762), .ZN(new_n1010));
  AND2_X1   g824(.A1(new_n1009), .A2(new_n1010), .ZN(new_n1011));
  NAND4_X1  g825(.A1(new_n794), .A2(new_n532), .A3(new_n745), .A4(new_n844), .ZN(new_n1012));
  NAND4_X1  g826(.A1(new_n804), .A2(new_n1011), .A3(new_n1012), .A4(new_n812), .ZN(new_n1013));
  OAI211_X1 g827(.A(new_n1007), .B(new_n1008), .C1(new_n1013), .C2(G953), .ZN(new_n1014));
  NAND3_X1  g828(.A1(new_n711), .A2(new_n762), .A3(new_n849), .ZN(new_n1015));
  XNOR2_X1  g829(.A(KEYINPUT123), .B(KEYINPUT62), .ZN(new_n1016));
  NAND2_X1  g830(.A1(new_n1015), .A2(new_n1016), .ZN(new_n1017));
  NAND2_X1  g831(.A1(KEYINPUT123), .A2(KEYINPUT62), .ZN(new_n1018));
  NAND3_X1  g832(.A1(new_n1010), .A2(new_n711), .A3(new_n1018), .ZN(new_n1019));
  INV_X1    g833(.A(new_n708), .ZN(new_n1020));
  NAND4_X1  g834(.A1(new_n727), .A2(new_n1020), .A3(new_n770), .A4(new_n829), .ZN(new_n1021));
  AND3_X1   g835(.A1(new_n1017), .A2(new_n1019), .A3(new_n1021), .ZN(new_n1022));
  INV_X1    g836(.A(KEYINPUT124), .ZN(new_n1023));
  NAND4_X1  g837(.A1(new_n1022), .A2(new_n1023), .A3(new_n804), .A4(new_n812), .ZN(new_n1024));
  NAND3_X1  g838(.A1(new_n1017), .A2(new_n1019), .A3(new_n1021), .ZN(new_n1025));
  NAND2_X1  g839(.A1(new_n804), .A2(new_n812), .ZN(new_n1026));
  OAI21_X1  g840(.A(KEYINPUT124), .B1(new_n1025), .B2(new_n1026), .ZN(new_n1027));
  AOI21_X1  g841(.A(G953), .B1(new_n1024), .B2(new_n1027), .ZN(new_n1028));
  OAI21_X1  g842(.A(new_n1014), .B1(new_n1028), .B2(new_n1007), .ZN(new_n1029));
  AOI21_X1  g843(.A(new_n189), .B1(G227), .B2(G900), .ZN(new_n1030));
  INV_X1    g844(.A(KEYINPUT125), .ZN(new_n1031));
  AOI21_X1  g845(.A(new_n1030), .B1(new_n1014), .B2(new_n1031), .ZN(new_n1032));
  AND2_X1   g846(.A1(new_n1029), .A2(new_n1032), .ZN(new_n1033));
  NOR2_X1   g847(.A1(new_n1029), .A2(new_n1032), .ZN(new_n1034));
  NOR2_X1   g848(.A1(new_n1033), .A2(new_n1034), .ZN(G72));
  INV_X1    g849(.A(new_n688), .ZN(new_n1036));
  NAND2_X1  g850(.A1(G472), .A2(G902), .ZN(new_n1037));
  XOR2_X1   g851(.A(new_n1037), .B(KEYINPUT63), .Z(new_n1038));
  NAND4_X1  g852(.A1(new_n983), .A2(new_n511), .A3(new_n1036), .A4(new_n1038), .ZN(new_n1039));
  OAI21_X1  g853(.A(new_n1038), .B1(new_n1000), .B2(new_n1013), .ZN(new_n1040));
  XNOR2_X1  g854(.A(new_n511), .B(KEYINPUT127), .ZN(new_n1041));
  AOI21_X1  g855(.A(new_n959), .B1(new_n1040), .B2(new_n1041), .ZN(new_n1042));
  NAND2_X1  g856(.A1(new_n1039), .A2(new_n1042), .ZN(new_n1043));
  NAND3_X1  g857(.A1(new_n1024), .A2(new_n1027), .A3(new_n860), .ZN(new_n1044));
  AOI21_X1  g858(.A(new_n1036), .B1(new_n1044), .B2(new_n1038), .ZN(new_n1045));
  OR2_X1    g859(.A1(new_n1045), .A2(KEYINPUT126), .ZN(new_n1046));
  NAND2_X1  g860(.A1(new_n1045), .A2(KEYINPUT126), .ZN(new_n1047));
  AOI21_X1  g861(.A(new_n1043), .B1(new_n1046), .B2(new_n1047), .ZN(G57));
endmodule


