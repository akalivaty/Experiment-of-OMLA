//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 0 1 1 0 1 0 1 0 1 0 0 0 0 1 0 0 1 0 1 0 1 0 1 0 0 0 0 0 0 1 0 0 0 0 0 0 0 0 0 1 0 1 0 0 1 0 0 0 1 0 1 0 0 1 1 0 0 1 1 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:19:55 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n689, new_n690, new_n691, new_n692,
    new_n693, new_n694, new_n695, new_n696, new_n697, new_n698, new_n700,
    new_n701, new_n702, new_n704, new_n705, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n730, new_n731,
    new_n732, new_n733, new_n734, new_n735, new_n737, new_n738, new_n739,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n764, new_n765, new_n766, new_n767, new_n769, new_n770,
    new_n771, new_n773, new_n774, new_n775, new_n776, new_n778, new_n779,
    new_n781, new_n782, new_n783, new_n784, new_n785, new_n786, new_n787,
    new_n788, new_n789, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n805, new_n806, new_n807, new_n808, new_n809, new_n810,
    new_n811, new_n812, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n878, new_n879, new_n881, new_n882, new_n883, new_n884,
    new_n886, new_n887, new_n888, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n927, new_n928, new_n930, new_n931,
    new_n932, new_n934, new_n935, new_n936, new_n937, new_n938, new_n940,
    new_n941, new_n943, new_n944, new_n945, new_n946, new_n947, new_n948,
    new_n950, new_n951, new_n952, new_n953, new_n954, new_n955, new_n956,
    new_n957, new_n958, new_n959, new_n960, new_n961, new_n962, new_n964,
    new_n965, new_n966, new_n967, new_n968, new_n969, new_n970, new_n971,
    new_n972, new_n973, new_n974, new_n975, new_n976, new_n977, new_n978,
    new_n979, new_n980, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n988, new_n989, new_n990, new_n991, new_n992, new_n993, new_n995,
    new_n996;
  AND2_X1   g000(.A1(KEYINPUT85), .A2(G29gat), .ZN(new_n202));
  NOR2_X1   g001(.A1(KEYINPUT85), .A2(G29gat), .ZN(new_n203));
  NOR2_X1   g002(.A1(new_n202), .A2(new_n203), .ZN(new_n204));
  AOI21_X1  g003(.A(KEYINPUT86), .B1(new_n204), .B2(G36gat), .ZN(new_n205));
  INV_X1    g004(.A(KEYINPUT86), .ZN(new_n206));
  INV_X1    g005(.A(G36gat), .ZN(new_n207));
  NOR4_X1   g006(.A1(new_n202), .A2(new_n203), .A3(new_n206), .A4(new_n207), .ZN(new_n208));
  OAI21_X1  g007(.A(KEYINPUT88), .B1(new_n205), .B2(new_n208), .ZN(new_n209));
  INV_X1    g008(.A(new_n203), .ZN(new_n210));
  NAND2_X1  g009(.A1(KEYINPUT85), .A2(G29gat), .ZN(new_n211));
  NAND3_X1  g010(.A1(new_n210), .A2(G36gat), .A3(new_n211), .ZN(new_n212));
  NAND2_X1  g011(.A1(new_n212), .A2(new_n206), .ZN(new_n213));
  NAND3_X1  g012(.A1(new_n204), .A2(KEYINPUT86), .A3(G36gat), .ZN(new_n214));
  INV_X1    g013(.A(KEYINPUT88), .ZN(new_n215));
  NAND3_X1  g014(.A1(new_n213), .A2(new_n214), .A3(new_n215), .ZN(new_n216));
  OAI21_X1  g015(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n217));
  INV_X1    g016(.A(KEYINPUT87), .ZN(new_n218));
  NAND2_X1  g017(.A1(new_n217), .A2(new_n218), .ZN(new_n219));
  INV_X1    g018(.A(KEYINPUT14), .ZN(new_n220));
  INV_X1    g019(.A(G29gat), .ZN(new_n221));
  NAND3_X1  g020(.A1(new_n220), .A2(new_n221), .A3(new_n207), .ZN(new_n222));
  XNOR2_X1  g021(.A(new_n219), .B(new_n222), .ZN(new_n223));
  NAND3_X1  g022(.A1(new_n209), .A2(new_n216), .A3(new_n223), .ZN(new_n224));
  XNOR2_X1  g023(.A(G43gat), .B(G50gat), .ZN(new_n225));
  NAND2_X1  g024(.A1(new_n225), .A2(KEYINPUT15), .ZN(new_n226));
  NAND2_X1  g025(.A1(new_n224), .A2(new_n226), .ZN(new_n227));
  NOR3_X1   g026(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n228));
  INV_X1    g027(.A(KEYINPUT84), .ZN(new_n229));
  XNOR2_X1  g028(.A(new_n228), .B(new_n229), .ZN(new_n230));
  INV_X1    g029(.A(KEYINPUT83), .ZN(new_n231));
  XNOR2_X1  g030(.A(new_n217), .B(new_n231), .ZN(new_n232));
  AOI21_X1  g031(.A(new_n226), .B1(new_n230), .B2(new_n232), .ZN(new_n233));
  NOR2_X1   g032(.A1(new_n205), .A2(new_n208), .ZN(new_n234));
  NAND2_X1  g033(.A1(new_n233), .A2(new_n234), .ZN(new_n235));
  NOR2_X1   g034(.A1(new_n225), .A2(KEYINPUT15), .ZN(new_n236));
  INV_X1    g035(.A(new_n236), .ZN(new_n237));
  NAND3_X1  g036(.A1(new_n227), .A2(new_n235), .A3(new_n237), .ZN(new_n238));
  INV_X1    g037(.A(G15gat), .ZN(new_n239));
  INV_X1    g038(.A(G22gat), .ZN(new_n240));
  NAND2_X1  g039(.A1(new_n239), .A2(new_n240), .ZN(new_n241));
  NAND2_X1  g040(.A1(G15gat), .A2(G22gat), .ZN(new_n242));
  AOI21_X1  g041(.A(KEYINPUT16), .B1(new_n241), .B2(new_n242), .ZN(new_n243));
  OR3_X1    g042(.A1(new_n243), .A2(G1gat), .A3(G8gat), .ZN(new_n244));
  AOI21_X1  g043(.A(KEYINPUT90), .B1(new_n241), .B2(new_n242), .ZN(new_n245));
  OAI21_X1  g044(.A(G8gat), .B1(new_n243), .B2(G1gat), .ZN(new_n246));
  AND3_X1   g045(.A1(new_n244), .A2(new_n245), .A3(new_n246), .ZN(new_n247));
  AOI21_X1  g046(.A(new_n245), .B1(new_n244), .B2(new_n246), .ZN(new_n248));
  NOR2_X1   g047(.A1(new_n247), .A2(new_n248), .ZN(new_n249));
  INV_X1    g048(.A(new_n249), .ZN(new_n250));
  AOI21_X1  g049(.A(KEYINPUT92), .B1(new_n238), .B2(new_n250), .ZN(new_n251));
  AOI221_X4 g050(.A(new_n236), .B1(new_n233), .B2(new_n234), .C1(new_n224), .C2(new_n226), .ZN(new_n252));
  NAND2_X1  g051(.A1(new_n252), .A2(new_n249), .ZN(new_n253));
  NAND2_X1  g052(.A1(new_n251), .A2(new_n253), .ZN(new_n254));
  NAND3_X1  g053(.A1(new_n252), .A2(KEYINPUT92), .A3(new_n249), .ZN(new_n255));
  AND2_X1   g054(.A1(new_n254), .A2(new_n255), .ZN(new_n256));
  NAND2_X1  g055(.A1(G229gat), .A2(G233gat), .ZN(new_n257));
  XNOR2_X1  g056(.A(new_n257), .B(KEYINPUT13), .ZN(new_n258));
  INV_X1    g057(.A(new_n258), .ZN(new_n259));
  INV_X1    g058(.A(KEYINPUT18), .ZN(new_n260));
  XNOR2_X1  g059(.A(KEYINPUT89), .B(KEYINPUT17), .ZN(new_n261));
  NAND4_X1  g060(.A1(new_n227), .A2(new_n235), .A3(new_n237), .A4(new_n261), .ZN(new_n262));
  INV_X1    g061(.A(KEYINPUT17), .ZN(new_n263));
  OAI211_X1 g062(.A(new_n250), .B(new_n262), .C1(new_n252), .C2(new_n263), .ZN(new_n264));
  NAND3_X1  g063(.A1(new_n264), .A2(new_n257), .A3(new_n253), .ZN(new_n265));
  AOI22_X1  g064(.A1(new_n256), .A2(new_n259), .B1(new_n260), .B2(new_n265), .ZN(new_n266));
  NAND4_X1  g065(.A1(new_n264), .A2(KEYINPUT18), .A3(new_n257), .A4(new_n253), .ZN(new_n267));
  NAND2_X1  g066(.A1(new_n267), .A2(KEYINPUT91), .ZN(new_n268));
  OR2_X1    g067(.A1(new_n267), .A2(KEYINPUT91), .ZN(new_n269));
  NAND3_X1  g068(.A1(new_n266), .A2(new_n268), .A3(new_n269), .ZN(new_n270));
  XNOR2_X1  g069(.A(G113gat), .B(G141gat), .ZN(new_n271));
  INV_X1    g070(.A(G197gat), .ZN(new_n272));
  XNOR2_X1  g071(.A(new_n271), .B(new_n272), .ZN(new_n273));
  XNOR2_X1  g072(.A(KEYINPUT11), .B(G169gat), .ZN(new_n274));
  XNOR2_X1  g073(.A(new_n273), .B(new_n274), .ZN(new_n275));
  XOR2_X1   g074(.A(KEYINPUT82), .B(KEYINPUT12), .Z(new_n276));
  XOR2_X1   g075(.A(new_n275), .B(new_n276), .Z(new_n277));
  INV_X1    g076(.A(new_n277), .ZN(new_n278));
  NAND2_X1  g077(.A1(new_n270), .A2(new_n278), .ZN(new_n279));
  INV_X1    g078(.A(KEYINPUT91), .ZN(new_n280));
  XNOR2_X1  g079(.A(new_n267), .B(new_n280), .ZN(new_n281));
  NAND3_X1  g080(.A1(new_n281), .A2(new_n277), .A3(new_n266), .ZN(new_n282));
  NAND2_X1  g081(.A1(new_n279), .A2(new_n282), .ZN(new_n283));
  INV_X1    g082(.A(new_n283), .ZN(new_n284));
  INV_X1    g083(.A(KEYINPUT35), .ZN(new_n285));
  NAND2_X1  g084(.A1(G227gat), .A2(G233gat), .ZN(new_n286));
  INV_X1    g085(.A(new_n286), .ZN(new_n287));
  NAND2_X1  g086(.A1(G183gat), .A2(G190gat), .ZN(new_n288));
  NAND2_X1  g087(.A1(new_n288), .A2(KEYINPUT24), .ZN(new_n289));
  INV_X1    g088(.A(KEYINPUT24), .ZN(new_n290));
  NAND3_X1  g089(.A1(new_n290), .A2(G183gat), .A3(G190gat), .ZN(new_n291));
  NAND2_X1  g090(.A1(new_n289), .A2(new_n291), .ZN(new_n292));
  INV_X1    g091(.A(G183gat), .ZN(new_n293));
  INV_X1    g092(.A(G190gat), .ZN(new_n294));
  NAND2_X1  g093(.A1(new_n293), .A2(new_n294), .ZN(new_n295));
  NAND2_X1  g094(.A1(new_n292), .A2(new_n295), .ZN(new_n296));
  NAND2_X1  g095(.A1(G169gat), .A2(G176gat), .ZN(new_n297));
  OR3_X1    g096(.A1(KEYINPUT23), .A2(G169gat), .A3(G176gat), .ZN(new_n298));
  OAI21_X1  g097(.A(KEYINPUT23), .B1(G169gat), .B2(G176gat), .ZN(new_n299));
  NAND2_X1  g098(.A1(new_n298), .A2(new_n299), .ZN(new_n300));
  NAND4_X1  g099(.A1(new_n296), .A2(KEYINPUT25), .A3(new_n297), .A4(new_n300), .ZN(new_n301));
  NAND2_X1  g100(.A1(new_n301), .A2(KEYINPUT64), .ZN(new_n302));
  NAND3_X1  g101(.A1(new_n296), .A2(new_n297), .A3(new_n300), .ZN(new_n303));
  INV_X1    g102(.A(KEYINPUT25), .ZN(new_n304));
  NAND2_X1  g103(.A1(new_n303), .A2(new_n304), .ZN(new_n305));
  NAND2_X1  g104(.A1(new_n302), .A2(new_n305), .ZN(new_n306));
  NAND3_X1  g105(.A1(new_n303), .A2(KEYINPUT64), .A3(new_n304), .ZN(new_n307));
  NAND2_X1  g106(.A1(new_n306), .A2(new_n307), .ZN(new_n308));
  INV_X1    g107(.A(G120gat), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n309), .A2(G113gat), .ZN(new_n310));
  INV_X1    g109(.A(G113gat), .ZN(new_n311));
  NAND2_X1  g110(.A1(new_n311), .A2(G120gat), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n310), .A2(new_n312), .ZN(new_n313));
  INV_X1    g112(.A(KEYINPUT1), .ZN(new_n314));
  NAND2_X1  g113(.A1(new_n313), .A2(new_n314), .ZN(new_n315));
  XNOR2_X1  g114(.A(KEYINPUT65), .B(G127gat), .ZN(new_n316));
  NAND2_X1  g115(.A1(new_n316), .A2(G134gat), .ZN(new_n317));
  OAI211_X1 g116(.A(new_n315), .B(new_n317), .C1(G127gat), .C2(G134gat), .ZN(new_n318));
  XNOR2_X1  g117(.A(G127gat), .B(G134gat), .ZN(new_n319));
  OR2_X1    g118(.A1(KEYINPUT66), .A2(G113gat), .ZN(new_n320));
  NAND2_X1  g119(.A1(KEYINPUT66), .A2(G113gat), .ZN(new_n321));
  AOI21_X1  g120(.A(new_n309), .B1(new_n320), .B2(new_n321), .ZN(new_n322));
  INV_X1    g121(.A(new_n310), .ZN(new_n323));
  OAI211_X1 g122(.A(new_n314), .B(new_n319), .C1(new_n322), .C2(new_n323), .ZN(new_n324));
  AND2_X1   g123(.A1(new_n318), .A2(new_n324), .ZN(new_n325));
  AND2_X1   g124(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n326));
  NOR2_X1   g125(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n327));
  OAI21_X1  g126(.A(new_n294), .B1(new_n326), .B2(new_n327), .ZN(new_n328));
  INV_X1    g127(.A(KEYINPUT28), .ZN(new_n329));
  XNOR2_X1  g128(.A(new_n328), .B(new_n329), .ZN(new_n330));
  AOI21_X1  g129(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n331));
  OAI21_X1  g130(.A(new_n331), .B1(G169gat), .B2(G176gat), .ZN(new_n332));
  INV_X1    g131(.A(G169gat), .ZN(new_n333));
  INV_X1    g132(.A(G176gat), .ZN(new_n334));
  NAND3_X1  g133(.A1(new_n333), .A2(new_n334), .A3(KEYINPUT26), .ZN(new_n335));
  NAND4_X1  g134(.A1(new_n330), .A2(new_n332), .A3(new_n335), .A4(new_n288), .ZN(new_n336));
  AND3_X1   g135(.A1(new_n308), .A2(new_n325), .A3(new_n336), .ZN(new_n337));
  AOI21_X1  g136(.A(new_n325), .B1(new_n308), .B2(new_n336), .ZN(new_n338));
  OAI21_X1  g137(.A(new_n287), .B1(new_n337), .B2(new_n338), .ZN(new_n339));
  NAND2_X1  g138(.A1(new_n339), .A2(KEYINPUT32), .ZN(new_n340));
  INV_X1    g139(.A(KEYINPUT33), .ZN(new_n341));
  NAND2_X1  g140(.A1(new_n339), .A2(new_n341), .ZN(new_n342));
  XNOR2_X1  g141(.A(G15gat), .B(G43gat), .ZN(new_n343));
  XNOR2_X1  g142(.A(G71gat), .B(G99gat), .ZN(new_n344));
  XOR2_X1   g143(.A(new_n343), .B(new_n344), .Z(new_n345));
  NAND3_X1  g144(.A1(new_n340), .A2(new_n342), .A3(new_n345), .ZN(new_n346));
  INV_X1    g145(.A(new_n345), .ZN(new_n347));
  OAI211_X1 g146(.A(new_n339), .B(KEYINPUT32), .C1(new_n341), .C2(new_n347), .ZN(new_n348));
  AOI22_X1  g147(.A1(new_n292), .A2(new_n295), .B1(G169gat), .B2(G176gat), .ZN(new_n349));
  AOI21_X1  g148(.A(KEYINPUT25), .B1(new_n349), .B2(new_n300), .ZN(new_n350));
  AOI21_X1  g149(.A(new_n350), .B1(KEYINPUT64), .B2(new_n301), .ZN(new_n351));
  INV_X1    g150(.A(new_n307), .ZN(new_n352));
  OAI21_X1  g151(.A(new_n336), .B1(new_n351), .B2(new_n352), .ZN(new_n353));
  NAND2_X1  g152(.A1(new_n318), .A2(new_n324), .ZN(new_n354));
  NAND2_X1  g153(.A1(new_n353), .A2(new_n354), .ZN(new_n355));
  NAND3_X1  g154(.A1(new_n308), .A2(new_n325), .A3(new_n336), .ZN(new_n356));
  NAND3_X1  g155(.A1(new_n355), .A2(new_n286), .A3(new_n356), .ZN(new_n357));
  INV_X1    g156(.A(KEYINPUT34), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n357), .A2(new_n358), .ZN(new_n359));
  NAND4_X1  g158(.A1(new_n355), .A2(KEYINPUT34), .A3(new_n286), .A4(new_n356), .ZN(new_n360));
  NAND2_X1  g159(.A1(new_n359), .A2(new_n360), .ZN(new_n361));
  NAND3_X1  g160(.A1(new_n346), .A2(new_n348), .A3(new_n361), .ZN(new_n362));
  NAND2_X1  g161(.A1(new_n362), .A2(KEYINPUT68), .ZN(new_n363));
  INV_X1    g162(.A(KEYINPUT68), .ZN(new_n364));
  NAND4_X1  g163(.A1(new_n346), .A2(new_n364), .A3(new_n348), .A4(new_n361), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n363), .A2(new_n365), .ZN(new_n366));
  XNOR2_X1  g165(.A(G78gat), .B(G106gat), .ZN(new_n367));
  XNOR2_X1  g166(.A(KEYINPUT31), .B(G50gat), .ZN(new_n368));
  XNOR2_X1  g167(.A(new_n367), .B(new_n368), .ZN(new_n369));
  INV_X1    g168(.A(new_n369), .ZN(new_n370));
  NAND2_X1  g169(.A1(G155gat), .A2(G162gat), .ZN(new_n371));
  INV_X1    g170(.A(G155gat), .ZN(new_n372));
  INV_X1    g171(.A(G162gat), .ZN(new_n373));
  NAND2_X1  g172(.A1(new_n372), .A2(new_n373), .ZN(new_n374));
  XNOR2_X1  g173(.A(G141gat), .B(G148gat), .ZN(new_n375));
  OAI211_X1 g174(.A(new_n371), .B(new_n374), .C1(new_n375), .C2(KEYINPUT2), .ZN(new_n376));
  NAND2_X1  g175(.A1(new_n376), .A2(KEYINPUT75), .ZN(new_n377));
  OAI21_X1  g176(.A(new_n371), .B1(new_n374), .B2(KEYINPUT2), .ZN(new_n378));
  INV_X1    g177(.A(G141gat), .ZN(new_n379));
  NOR2_X1   g178(.A1(new_n379), .A2(G148gat), .ZN(new_n380));
  INV_X1    g179(.A(G148gat), .ZN(new_n381));
  NOR2_X1   g180(.A1(new_n381), .A2(G141gat), .ZN(new_n382));
  OAI21_X1  g181(.A(new_n378), .B1(new_n380), .B2(new_n382), .ZN(new_n383));
  INV_X1    g182(.A(KEYINPUT2), .ZN(new_n384));
  OAI21_X1  g183(.A(new_n384), .B1(new_n380), .B2(new_n382), .ZN(new_n385));
  INV_X1    g184(.A(KEYINPUT75), .ZN(new_n386));
  NAND4_X1  g185(.A1(new_n385), .A2(new_n386), .A3(new_n371), .A4(new_n374), .ZN(new_n387));
  AND3_X1   g186(.A1(new_n377), .A2(new_n383), .A3(new_n387), .ZN(new_n388));
  OR2_X1    g187(.A1(KEYINPUT70), .A2(G197gat), .ZN(new_n389));
  NAND2_X1  g188(.A1(KEYINPUT70), .A2(G197gat), .ZN(new_n390));
  NAND3_X1  g189(.A1(new_n389), .A2(G204gat), .A3(new_n390), .ZN(new_n391));
  INV_X1    g190(.A(G204gat), .ZN(new_n392));
  AND2_X1   g191(.A1(KEYINPUT70), .A2(G197gat), .ZN(new_n393));
  NOR2_X1   g192(.A1(KEYINPUT70), .A2(G197gat), .ZN(new_n394));
  OAI21_X1  g193(.A(new_n392), .B1(new_n393), .B2(new_n394), .ZN(new_n395));
  NAND2_X1  g194(.A1(G211gat), .A2(G218gat), .ZN(new_n396));
  INV_X1    g195(.A(KEYINPUT22), .ZN(new_n397));
  AND3_X1   g196(.A1(new_n396), .A2(KEYINPUT71), .A3(new_n397), .ZN(new_n398));
  AOI21_X1  g197(.A(KEYINPUT71), .B1(new_n396), .B2(new_n397), .ZN(new_n399));
  OAI211_X1 g198(.A(new_n391), .B(new_n395), .C1(new_n398), .C2(new_n399), .ZN(new_n400));
  NAND2_X1  g199(.A1(new_n400), .A2(KEYINPUT72), .ZN(new_n401));
  XNOR2_X1  g200(.A(G211gat), .B(G218gat), .ZN(new_n402));
  INV_X1    g201(.A(new_n402), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n401), .A2(new_n403), .ZN(new_n404));
  INV_X1    g203(.A(KEYINPUT29), .ZN(new_n405));
  NAND3_X1  g204(.A1(new_n400), .A2(KEYINPUT72), .A3(new_n402), .ZN(new_n406));
  NAND3_X1  g205(.A1(new_n404), .A2(new_n405), .A3(new_n406), .ZN(new_n407));
  INV_X1    g206(.A(KEYINPUT3), .ZN(new_n408));
  AOI21_X1  g207(.A(new_n388), .B1(new_n407), .B2(new_n408), .ZN(new_n409));
  NAND2_X1  g208(.A1(G228gat), .A2(G233gat), .ZN(new_n410));
  NAND4_X1  g209(.A1(new_n377), .A2(new_n408), .A3(new_n387), .A4(new_n383), .ZN(new_n411));
  AOI22_X1  g210(.A1(new_n405), .A2(new_n411), .B1(new_n404), .B2(new_n406), .ZN(new_n412));
  NOR3_X1   g211(.A1(new_n409), .A2(new_n410), .A3(new_n412), .ZN(new_n413));
  INV_X1    g212(.A(KEYINPUT77), .ZN(new_n414));
  NAND3_X1  g213(.A1(new_n377), .A2(new_n383), .A3(new_n387), .ZN(new_n415));
  AND2_X1   g214(.A1(new_n400), .A2(new_n402), .ZN(new_n416));
  OAI21_X1  g215(.A(new_n405), .B1(new_n400), .B2(new_n402), .ZN(new_n417));
  OAI21_X1  g216(.A(new_n408), .B1(new_n416), .B2(new_n417), .ZN(new_n418));
  NAND2_X1  g217(.A1(new_n411), .A2(new_n405), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n404), .A2(new_n406), .ZN(new_n420));
  AOI22_X1  g219(.A1(new_n415), .A2(new_n418), .B1(new_n419), .B2(new_n420), .ZN(new_n421));
  INV_X1    g220(.A(new_n410), .ZN(new_n422));
  OAI21_X1  g221(.A(new_n414), .B1(new_n421), .B2(new_n422), .ZN(new_n423));
  AND2_X1   g222(.A1(new_n418), .A2(new_n415), .ZN(new_n424));
  OAI211_X1 g223(.A(KEYINPUT77), .B(new_n410), .C1(new_n424), .C2(new_n412), .ZN(new_n425));
  AOI21_X1  g224(.A(new_n413), .B1(new_n423), .B2(new_n425), .ZN(new_n426));
  INV_X1    g225(.A(KEYINPUT79), .ZN(new_n427));
  XNOR2_X1  g226(.A(KEYINPUT78), .B(G22gat), .ZN(new_n428));
  NAND3_X1  g227(.A1(new_n426), .A2(new_n427), .A3(new_n428), .ZN(new_n429));
  OAI21_X1  g228(.A(KEYINPUT79), .B1(new_n426), .B2(new_n428), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n423), .A2(new_n425), .ZN(new_n431));
  INV_X1    g230(.A(new_n413), .ZN(new_n432));
  AND3_X1   g231(.A1(new_n431), .A2(new_n432), .A3(new_n428), .ZN(new_n433));
  OAI211_X1 g232(.A(new_n370), .B(new_n429), .C1(new_n430), .C2(new_n433), .ZN(new_n434));
  NAND2_X1  g233(.A1(new_n431), .A2(new_n432), .ZN(new_n435));
  INV_X1    g234(.A(KEYINPUT80), .ZN(new_n436));
  NAND3_X1  g235(.A1(new_n435), .A2(new_n436), .A3(G22gat), .ZN(new_n437));
  OAI21_X1  g236(.A(KEYINPUT80), .B1(new_n426), .B2(new_n240), .ZN(new_n438));
  NAND2_X1  g237(.A1(new_n426), .A2(new_n428), .ZN(new_n439));
  NAND4_X1  g238(.A1(new_n437), .A2(new_n438), .A3(new_n369), .A4(new_n439), .ZN(new_n440));
  NAND2_X1  g239(.A1(new_n434), .A2(new_n440), .ZN(new_n441));
  INV_X1    g240(.A(KEYINPUT69), .ZN(new_n442));
  INV_X1    g241(.A(new_n361), .ZN(new_n443));
  AOI21_X1  g242(.A(new_n286), .B1(new_n355), .B2(new_n356), .ZN(new_n444));
  OAI21_X1  g243(.A(new_n345), .B1(new_n444), .B2(KEYINPUT33), .ZN(new_n445));
  INV_X1    g244(.A(KEYINPUT32), .ZN(new_n446));
  NOR2_X1   g245(.A1(new_n444), .A2(new_n446), .ZN(new_n447));
  NOR2_X1   g246(.A1(new_n445), .A2(new_n447), .ZN(new_n448));
  INV_X1    g247(.A(new_n348), .ZN(new_n449));
  OAI211_X1 g248(.A(new_n442), .B(new_n443), .C1(new_n448), .C2(new_n449), .ZN(new_n450));
  OAI21_X1  g249(.A(new_n443), .B1(new_n448), .B2(new_n449), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n451), .A2(KEYINPUT69), .ZN(new_n452));
  NAND4_X1  g251(.A1(new_n366), .A2(new_n441), .A3(new_n450), .A4(new_n452), .ZN(new_n453));
  XNOR2_X1  g252(.A(G1gat), .B(G29gat), .ZN(new_n454));
  INV_X1    g253(.A(G85gat), .ZN(new_n455));
  XNOR2_X1  g254(.A(new_n454), .B(new_n455), .ZN(new_n456));
  XNOR2_X1  g255(.A(KEYINPUT0), .B(G57gat), .ZN(new_n457));
  XOR2_X1   g256(.A(new_n456), .B(new_n457), .Z(new_n458));
  INV_X1    g257(.A(KEYINPUT4), .ZN(new_n459));
  NAND3_X1  g258(.A1(new_n388), .A2(new_n459), .A3(new_n325), .ZN(new_n460));
  OAI21_X1  g259(.A(KEYINPUT4), .B1(new_n415), .B2(new_n354), .ZN(new_n461));
  NAND2_X1  g260(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  NAND2_X1  g261(.A1(G225gat), .A2(G233gat), .ZN(new_n463));
  NAND2_X1  g262(.A1(new_n415), .A2(KEYINPUT3), .ZN(new_n464));
  NAND3_X1  g263(.A1(new_n464), .A2(new_n354), .A3(new_n411), .ZN(new_n465));
  NAND3_X1  g264(.A1(new_n462), .A2(new_n463), .A3(new_n465), .ZN(new_n466));
  INV_X1    g265(.A(KEYINPUT5), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  NAND2_X1  g267(.A1(new_n388), .A2(new_n325), .ZN(new_n469));
  NAND2_X1  g268(.A1(new_n415), .A2(new_n354), .ZN(new_n470));
  AOI21_X1  g269(.A(new_n463), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  AOI21_X1  g270(.A(new_n325), .B1(KEYINPUT3), .B2(new_n415), .ZN(new_n472));
  AOI22_X1  g271(.A1(new_n472), .A2(new_n411), .B1(new_n460), .B2(new_n461), .ZN(new_n473));
  AOI21_X1  g272(.A(new_n471), .B1(new_n473), .B2(new_n463), .ZN(new_n474));
  OAI211_X1 g273(.A(new_n458), .B(new_n468), .C1(new_n474), .C2(new_n467), .ZN(new_n475));
  NOR2_X1   g274(.A1(new_n475), .A2(KEYINPUT6), .ZN(new_n476));
  INV_X1    g275(.A(new_n458), .ZN(new_n477));
  INV_X1    g276(.A(new_n471), .ZN(new_n478));
  AOI21_X1  g277(.A(new_n467), .B1(new_n466), .B2(new_n478), .ZN(new_n479));
  AOI21_X1  g278(.A(KEYINPUT5), .B1(new_n473), .B2(new_n463), .ZN(new_n480));
  OAI21_X1  g279(.A(new_n477), .B1(new_n479), .B2(new_n480), .ZN(new_n481));
  NAND2_X1  g280(.A1(new_n481), .A2(KEYINPUT76), .ZN(new_n482));
  INV_X1    g281(.A(KEYINPUT6), .ZN(new_n483));
  INV_X1    g282(.A(KEYINPUT76), .ZN(new_n484));
  OAI211_X1 g283(.A(new_n484), .B(new_n477), .C1(new_n479), .C2(new_n480), .ZN(new_n485));
  NAND3_X1  g284(.A1(new_n482), .A2(new_n483), .A3(new_n485), .ZN(new_n486));
  AOI21_X1  g285(.A(new_n476), .B1(new_n486), .B2(new_n475), .ZN(new_n487));
  INV_X1    g286(.A(KEYINPUT30), .ZN(new_n488));
  XNOR2_X1  g287(.A(G8gat), .B(G36gat), .ZN(new_n489));
  XNOR2_X1  g288(.A(G64gat), .B(G92gat), .ZN(new_n490));
  XNOR2_X1  g289(.A(new_n489), .B(new_n490), .ZN(new_n491));
  NAND2_X1  g290(.A1(G226gat), .A2(G233gat), .ZN(new_n492));
  AND3_X1   g291(.A1(new_n308), .A2(new_n492), .A3(new_n336), .ZN(new_n493));
  AOI21_X1  g292(.A(KEYINPUT29), .B1(G226gat), .B2(G233gat), .ZN(new_n494));
  AOI21_X1  g293(.A(new_n494), .B1(new_n308), .B2(new_n336), .ZN(new_n495));
  OAI21_X1  g294(.A(new_n420), .B1(new_n493), .B2(new_n495), .ZN(new_n496));
  INV_X1    g295(.A(KEYINPUT73), .ZN(new_n497));
  NAND3_X1  g296(.A1(new_n308), .A2(new_n492), .A3(new_n336), .ZN(new_n498));
  INV_X1    g297(.A(new_n420), .ZN(new_n499));
  AND3_X1   g298(.A1(new_n330), .A2(new_n335), .A3(new_n288), .ZN(new_n500));
  AOI22_X1  g299(.A1(new_n306), .A2(new_n307), .B1(new_n500), .B2(new_n332), .ZN(new_n501));
  OAI211_X1 g300(.A(new_n498), .B(new_n499), .C1(new_n501), .C2(new_n494), .ZN(new_n502));
  NAND3_X1  g301(.A1(new_n496), .A2(new_n497), .A3(new_n502), .ZN(new_n503));
  OAI211_X1 g302(.A(KEYINPUT73), .B(new_n420), .C1(new_n493), .C2(new_n495), .ZN(new_n504));
  AOI21_X1  g303(.A(new_n491), .B1(new_n503), .B2(new_n504), .ZN(new_n505));
  INV_X1    g304(.A(KEYINPUT74), .ZN(new_n506));
  NOR2_X1   g305(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  AOI211_X1 g306(.A(KEYINPUT74), .B(new_n491), .C1(new_n503), .C2(new_n504), .ZN(new_n508));
  OAI21_X1  g307(.A(new_n488), .B1(new_n507), .B2(new_n508), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n503), .A2(new_n504), .ZN(new_n510));
  INV_X1    g309(.A(new_n491), .ZN(new_n511));
  NOR2_X1   g310(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  AOI21_X1  g311(.A(new_n512), .B1(KEYINPUT30), .B2(new_n505), .ZN(new_n513));
  NAND3_X1  g312(.A1(new_n487), .A2(new_n509), .A3(new_n513), .ZN(new_n514));
  OAI21_X1  g313(.A(new_n285), .B1(new_n453), .B2(new_n514), .ZN(new_n515));
  AND3_X1   g314(.A1(new_n487), .A2(new_n509), .A3(new_n513), .ZN(new_n516));
  NAND3_X1  g315(.A1(new_n359), .A2(KEYINPUT67), .A3(new_n360), .ZN(new_n517));
  AND3_X1   g316(.A1(new_n346), .A2(new_n348), .A3(new_n517), .ZN(new_n518));
  AOI21_X1  g317(.A(new_n517), .B1(new_n346), .B2(new_n348), .ZN(new_n519));
  NOR2_X1   g318(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  AND3_X1   g319(.A1(new_n441), .A2(new_n520), .A3(KEYINPUT35), .ZN(new_n521));
  NAND2_X1  g320(.A1(new_n516), .A2(new_n521), .ZN(new_n522));
  AND2_X1   g321(.A1(new_n515), .A2(new_n522), .ZN(new_n523));
  NAND3_X1  g322(.A1(new_n366), .A2(new_n450), .A3(new_n452), .ZN(new_n524));
  INV_X1    g323(.A(KEYINPUT36), .ZN(new_n525));
  NAND2_X1  g324(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  NAND2_X1  g325(.A1(new_n520), .A2(KEYINPUT36), .ZN(new_n527));
  NAND2_X1  g326(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  OR3_X1    g327(.A1(new_n473), .A2(KEYINPUT39), .A3(new_n463), .ZN(new_n529));
  NAND3_X1  g328(.A1(new_n469), .A2(new_n463), .A3(new_n470), .ZN(new_n530));
  OAI211_X1 g329(.A(new_n530), .B(KEYINPUT39), .C1(new_n473), .C2(new_n463), .ZN(new_n531));
  NAND3_X1  g330(.A1(new_n529), .A2(new_n477), .A3(new_n531), .ZN(new_n532));
  INV_X1    g331(.A(KEYINPUT40), .ZN(new_n533));
  OR2_X1    g332(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  AND2_X1   g333(.A1(new_n534), .A2(new_n475), .ZN(new_n535));
  NAND2_X1  g334(.A1(new_n532), .A2(new_n533), .ZN(new_n536));
  INV_X1    g335(.A(KEYINPUT81), .ZN(new_n537));
  XNOR2_X1  g336(.A(new_n536), .B(new_n537), .ZN(new_n538));
  NAND2_X1  g337(.A1(new_n510), .A2(new_n511), .ZN(new_n539));
  NAND2_X1  g338(.A1(new_n539), .A2(KEYINPUT74), .ZN(new_n540));
  NAND2_X1  g339(.A1(new_n505), .A2(new_n506), .ZN(new_n541));
  AOI21_X1  g340(.A(KEYINPUT30), .B1(new_n540), .B2(new_n541), .ZN(new_n542));
  NAND2_X1  g341(.A1(new_n505), .A2(KEYINPUT30), .ZN(new_n543));
  OAI21_X1  g342(.A(new_n543), .B1(new_n510), .B2(new_n511), .ZN(new_n544));
  OAI211_X1 g343(.A(new_n535), .B(new_n538), .C1(new_n542), .C2(new_n544), .ZN(new_n545));
  INV_X1    g344(.A(KEYINPUT37), .ZN(new_n546));
  NAND2_X1  g345(.A1(new_n510), .A2(new_n546), .ZN(new_n547));
  NAND3_X1  g346(.A1(new_n503), .A2(KEYINPUT37), .A3(new_n504), .ZN(new_n548));
  NAND4_X1  g347(.A1(new_n547), .A2(KEYINPUT38), .A3(new_n491), .A4(new_n548), .ZN(new_n549));
  AOI21_X1  g348(.A(new_n546), .B1(new_n496), .B2(new_n502), .ZN(new_n550));
  AOI211_X1 g349(.A(new_n511), .B(new_n550), .C1(new_n510), .C2(new_n546), .ZN(new_n551));
  OAI21_X1  g350(.A(new_n549), .B1(new_n551), .B2(KEYINPUT38), .ZN(new_n552));
  NAND2_X1  g351(.A1(new_n485), .A2(new_n483), .ZN(new_n553));
  OAI21_X1  g352(.A(new_n468), .B1(new_n474), .B2(new_n467), .ZN(new_n554));
  AOI21_X1  g353(.A(new_n484), .B1(new_n554), .B2(new_n477), .ZN(new_n555));
  OAI21_X1  g354(.A(new_n475), .B1(new_n553), .B2(new_n555), .ZN(new_n556));
  INV_X1    g355(.A(new_n476), .ZN(new_n557));
  NAND2_X1  g356(.A1(new_n556), .A2(new_n557), .ZN(new_n558));
  NAND2_X1  g357(.A1(new_n540), .A2(new_n541), .ZN(new_n559));
  NAND3_X1  g358(.A1(new_n552), .A2(new_n558), .A3(new_n559), .ZN(new_n560));
  NAND3_X1  g359(.A1(new_n545), .A2(new_n560), .A3(new_n441), .ZN(new_n561));
  INV_X1    g360(.A(new_n441), .ZN(new_n562));
  NAND2_X1  g361(.A1(new_n514), .A2(new_n562), .ZN(new_n563));
  NAND3_X1  g362(.A1(new_n528), .A2(new_n561), .A3(new_n563), .ZN(new_n564));
  AOI21_X1  g363(.A(new_n284), .B1(new_n523), .B2(new_n564), .ZN(new_n565));
  INV_X1    g364(.A(KEYINPUT101), .ZN(new_n566));
  INV_X1    g365(.A(G57gat), .ZN(new_n567));
  OAI21_X1  g366(.A(KEYINPUT94), .B1(new_n567), .B2(G64gat), .ZN(new_n568));
  INV_X1    g367(.A(KEYINPUT94), .ZN(new_n569));
  INV_X1    g368(.A(G64gat), .ZN(new_n570));
  NAND3_X1  g369(.A1(new_n569), .A2(new_n570), .A3(G57gat), .ZN(new_n571));
  NAND2_X1  g370(.A1(new_n567), .A2(G64gat), .ZN(new_n572));
  NAND3_X1  g371(.A1(new_n568), .A2(new_n571), .A3(new_n572), .ZN(new_n573));
  AND2_X1   g372(.A1(G71gat), .A2(G78gat), .ZN(new_n574));
  OR2_X1    g373(.A1(new_n574), .A2(KEYINPUT9), .ZN(new_n575));
  XNOR2_X1  g374(.A(G71gat), .B(G78gat), .ZN(new_n576));
  NAND3_X1  g375(.A1(new_n573), .A2(new_n575), .A3(new_n576), .ZN(new_n577));
  NAND2_X1  g376(.A1(new_n570), .A2(G57gat), .ZN(new_n578));
  INV_X1    g377(.A(KEYINPUT93), .ZN(new_n579));
  AND3_X1   g378(.A1(new_n572), .A2(new_n578), .A3(new_n579), .ZN(new_n580));
  AOI21_X1  g379(.A(new_n579), .B1(new_n572), .B2(new_n578), .ZN(new_n581));
  NOR2_X1   g380(.A1(new_n574), .A2(KEYINPUT9), .ZN(new_n582));
  NOR3_X1   g381(.A1(new_n580), .A2(new_n581), .A3(new_n582), .ZN(new_n583));
  OAI21_X1  g382(.A(new_n577), .B1(new_n583), .B2(new_n576), .ZN(new_n584));
  INV_X1    g383(.A(KEYINPUT21), .ZN(new_n585));
  NAND2_X1  g384(.A1(new_n584), .A2(new_n585), .ZN(new_n586));
  XOR2_X1   g385(.A(new_n586), .B(G211gat), .Z(new_n587));
  INV_X1    g386(.A(new_n587), .ZN(new_n588));
  OAI21_X1  g387(.A(new_n250), .B1(new_n585), .B2(new_n584), .ZN(new_n589));
  XNOR2_X1  g388(.A(new_n589), .B(G183gat), .ZN(new_n590));
  XNOR2_X1  g389(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n591));
  INV_X1    g390(.A(new_n591), .ZN(new_n592));
  NAND2_X1  g391(.A1(new_n590), .A2(new_n592), .ZN(new_n593));
  XNOR2_X1  g392(.A(new_n589), .B(new_n293), .ZN(new_n594));
  NAND2_X1  g393(.A1(new_n594), .A2(new_n591), .ZN(new_n595));
  AOI21_X1  g394(.A(new_n588), .B1(new_n593), .B2(new_n595), .ZN(new_n596));
  INV_X1    g395(.A(new_n596), .ZN(new_n597));
  XNOR2_X1  g396(.A(G127gat), .B(G155gat), .ZN(new_n598));
  NAND2_X1  g397(.A1(G231gat), .A2(G233gat), .ZN(new_n599));
  XNOR2_X1  g398(.A(new_n598), .B(new_n599), .ZN(new_n600));
  NAND3_X1  g399(.A1(new_n593), .A2(new_n595), .A3(new_n588), .ZN(new_n601));
  NAND3_X1  g400(.A1(new_n597), .A2(new_n600), .A3(new_n601), .ZN(new_n602));
  INV_X1    g401(.A(new_n600), .ZN(new_n603));
  INV_X1    g402(.A(new_n601), .ZN(new_n604));
  OAI21_X1  g403(.A(new_n603), .B1(new_n604), .B2(new_n596), .ZN(new_n605));
  NAND2_X1  g404(.A1(new_n602), .A2(new_n605), .ZN(new_n606));
  XOR2_X1   g405(.A(G190gat), .B(G218gat), .Z(new_n607));
  INV_X1    g406(.A(new_n607), .ZN(new_n608));
  NAND2_X1  g407(.A1(new_n608), .A2(KEYINPUT99), .ZN(new_n609));
  INV_X1    g408(.A(KEYINPUT96), .ZN(new_n610));
  NAND2_X1  g409(.A1(new_n610), .A2(KEYINPUT7), .ZN(new_n611));
  AND3_X1   g410(.A1(KEYINPUT97), .A2(G85gat), .A3(G92gat), .ZN(new_n612));
  AOI21_X1  g411(.A(KEYINPUT97), .B1(G85gat), .B2(G92gat), .ZN(new_n613));
  OAI21_X1  g412(.A(new_n611), .B1(new_n612), .B2(new_n613), .ZN(new_n614));
  NAND2_X1  g413(.A1(G85gat), .A2(G92gat), .ZN(new_n615));
  INV_X1    g414(.A(KEYINPUT97), .ZN(new_n616));
  NAND2_X1  g415(.A1(new_n615), .A2(new_n616), .ZN(new_n617));
  INV_X1    g416(.A(KEYINPUT7), .ZN(new_n618));
  NOR2_X1   g417(.A1(new_n618), .A2(KEYINPUT96), .ZN(new_n619));
  NAND3_X1  g418(.A1(KEYINPUT97), .A2(G85gat), .A3(G92gat), .ZN(new_n620));
  NAND3_X1  g419(.A1(new_n617), .A2(new_n619), .A3(new_n620), .ZN(new_n621));
  NAND2_X1  g420(.A1(G99gat), .A2(G106gat), .ZN(new_n622));
  INV_X1    g421(.A(G92gat), .ZN(new_n623));
  AOI22_X1  g422(.A1(KEYINPUT8), .A2(new_n622), .B1(new_n455), .B2(new_n623), .ZN(new_n624));
  NAND3_X1  g423(.A1(new_n614), .A2(new_n621), .A3(new_n624), .ZN(new_n625));
  XNOR2_X1  g424(.A(G99gat), .B(G106gat), .ZN(new_n626));
  INV_X1    g425(.A(new_n626), .ZN(new_n627));
  INV_X1    g426(.A(KEYINPUT98), .ZN(new_n628));
  NAND2_X1  g427(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  NAND2_X1  g428(.A1(new_n626), .A2(KEYINPUT98), .ZN(new_n630));
  AND3_X1   g429(.A1(new_n625), .A2(new_n629), .A3(new_n630), .ZN(new_n631));
  AOI21_X1  g430(.A(new_n629), .B1(new_n625), .B2(new_n630), .ZN(new_n632));
  NOR2_X1   g431(.A1(new_n631), .A2(new_n632), .ZN(new_n633));
  OAI21_X1  g432(.A(new_n609), .B1(new_n238), .B2(new_n633), .ZN(new_n634));
  AND2_X1   g433(.A1(G232gat), .A2(G233gat), .ZN(new_n635));
  AOI21_X1  g434(.A(new_n634), .B1(KEYINPUT41), .B2(new_n635), .ZN(new_n636));
  XOR2_X1   g435(.A(G134gat), .B(G162gat), .Z(new_n637));
  INV_X1    g436(.A(new_n637), .ZN(new_n638));
  OAI211_X1 g437(.A(new_n262), .B(new_n633), .C1(new_n252), .C2(new_n263), .ZN(new_n639));
  AND3_X1   g438(.A1(new_n636), .A2(new_n638), .A3(new_n639), .ZN(new_n640));
  NOR2_X1   g439(.A1(new_n608), .A2(KEYINPUT99), .ZN(new_n641));
  AOI21_X1  g440(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n642));
  XNOR2_X1  g441(.A(new_n641), .B(new_n642), .ZN(new_n643));
  XNOR2_X1  g442(.A(new_n643), .B(KEYINPUT95), .ZN(new_n644));
  INV_X1    g443(.A(new_n644), .ZN(new_n645));
  AOI21_X1  g444(.A(new_n638), .B1(new_n636), .B2(new_n639), .ZN(new_n646));
  OR3_X1    g445(.A1(new_n640), .A2(new_n645), .A3(new_n646), .ZN(new_n647));
  OAI21_X1  g446(.A(new_n645), .B1(new_n640), .B2(new_n646), .ZN(new_n648));
  NAND2_X1  g447(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  INV_X1    g448(.A(new_n649), .ZN(new_n650));
  NAND2_X1  g449(.A1(new_n606), .A2(new_n650), .ZN(new_n651));
  INV_X1    g450(.A(KEYINPUT100), .ZN(new_n652));
  NAND2_X1  g451(.A1(new_n625), .A2(new_n652), .ZN(new_n653));
  NAND2_X1  g452(.A1(new_n653), .A2(new_n627), .ZN(new_n654));
  NOR2_X1   g453(.A1(new_n570), .A2(G57gat), .ZN(new_n655));
  NOR2_X1   g454(.A1(new_n567), .A2(G64gat), .ZN(new_n656));
  OAI21_X1  g455(.A(KEYINPUT93), .B1(new_n655), .B2(new_n656), .ZN(new_n657));
  NAND3_X1  g456(.A1(new_n572), .A2(new_n578), .A3(new_n579), .ZN(new_n658));
  NAND3_X1  g457(.A1(new_n657), .A2(new_n575), .A3(new_n658), .ZN(new_n659));
  INV_X1    g458(.A(new_n576), .ZN(new_n660));
  NAND2_X1  g459(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  NAND3_X1  g460(.A1(new_n625), .A2(new_n652), .A3(new_n626), .ZN(new_n662));
  NAND4_X1  g461(.A1(new_n654), .A2(new_n661), .A3(new_n577), .A4(new_n662), .ZN(new_n663));
  OAI21_X1  g462(.A(new_n584), .B1(new_n631), .B2(new_n632), .ZN(new_n664));
  AOI21_X1  g463(.A(KEYINPUT10), .B1(new_n663), .B2(new_n664), .ZN(new_n665));
  OAI21_X1  g464(.A(KEYINPUT10), .B1(new_n631), .B2(new_n632), .ZN(new_n666));
  NOR2_X1   g465(.A1(new_n666), .A2(new_n584), .ZN(new_n667));
  INV_X1    g466(.A(G230gat), .ZN(new_n668));
  INV_X1    g467(.A(G233gat), .ZN(new_n669));
  OAI22_X1  g468(.A1(new_n665), .A2(new_n667), .B1(new_n668), .B2(new_n669), .ZN(new_n670));
  NOR2_X1   g469(.A1(new_n668), .A2(new_n669), .ZN(new_n671));
  NAND3_X1  g470(.A1(new_n663), .A2(new_n664), .A3(new_n671), .ZN(new_n672));
  NAND2_X1  g471(.A1(new_n670), .A2(new_n672), .ZN(new_n673));
  XNOR2_X1  g472(.A(G120gat), .B(G148gat), .ZN(new_n674));
  XNOR2_X1  g473(.A(G176gat), .B(G204gat), .ZN(new_n675));
  XNOR2_X1  g474(.A(new_n674), .B(new_n675), .ZN(new_n676));
  NAND2_X1  g475(.A1(new_n673), .A2(new_n676), .ZN(new_n677));
  INV_X1    g476(.A(new_n676), .ZN(new_n678));
  NAND3_X1  g477(.A1(new_n670), .A2(new_n672), .A3(new_n678), .ZN(new_n679));
  AND2_X1   g478(.A1(new_n677), .A2(new_n679), .ZN(new_n680));
  INV_X1    g479(.A(new_n680), .ZN(new_n681));
  OAI21_X1  g480(.A(new_n566), .B1(new_n651), .B2(new_n681), .ZN(new_n682));
  NAND4_X1  g481(.A1(new_n606), .A2(KEYINPUT101), .A3(new_n650), .A4(new_n680), .ZN(new_n683));
  AND2_X1   g482(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  NAND2_X1  g483(.A1(new_n565), .A2(new_n684), .ZN(new_n685));
  INV_X1    g484(.A(new_n685), .ZN(new_n686));
  NAND2_X1  g485(.A1(new_n686), .A2(new_n558), .ZN(new_n687));
  XNOR2_X1  g486(.A(new_n687), .B(G1gat), .ZN(G1324gat));
  NOR2_X1   g487(.A1(new_n542), .A2(new_n544), .ZN(new_n689));
  INV_X1    g488(.A(new_n689), .ZN(new_n690));
  NAND2_X1  g489(.A1(new_n686), .A2(new_n690), .ZN(new_n691));
  INV_X1    g490(.A(KEYINPUT42), .ZN(new_n692));
  XNOR2_X1  g491(.A(KEYINPUT16), .B(G8gat), .ZN(new_n693));
  OR3_X1    g492(.A1(new_n691), .A2(new_n692), .A3(new_n693), .ZN(new_n694));
  NAND2_X1  g493(.A1(new_n691), .A2(G8gat), .ZN(new_n695));
  OAI21_X1  g494(.A(new_n692), .B1(new_n691), .B2(new_n693), .ZN(new_n696));
  NAND3_X1  g495(.A1(new_n694), .A2(new_n695), .A3(new_n696), .ZN(new_n697));
  INV_X1    g496(.A(KEYINPUT102), .ZN(new_n698));
  XNOR2_X1  g497(.A(new_n697), .B(new_n698), .ZN(G1325gat));
  NOR3_X1   g498(.A1(new_n685), .A2(new_n239), .A3(new_n528), .ZN(new_n700));
  INV_X1    g499(.A(new_n524), .ZN(new_n701));
  NAND2_X1  g500(.A1(new_n686), .A2(new_n701), .ZN(new_n702));
  AOI21_X1  g501(.A(new_n700), .B1(new_n239), .B2(new_n702), .ZN(G1326gat));
  NOR2_X1   g502(.A1(new_n685), .A2(new_n441), .ZN(new_n704));
  XOR2_X1   g503(.A(KEYINPUT43), .B(G22gat), .Z(new_n705));
  XNOR2_X1  g504(.A(new_n704), .B(new_n705), .ZN(G1327gat));
  NOR3_X1   g505(.A1(new_n606), .A2(new_n650), .A3(new_n681), .ZN(new_n707));
  AND2_X1   g506(.A1(new_n565), .A2(new_n707), .ZN(new_n708));
  OAI211_X1 g507(.A(new_n708), .B(new_n558), .C1(new_n203), .C2(new_n202), .ZN(new_n709));
  XNOR2_X1  g508(.A(new_n709), .B(KEYINPUT45), .ZN(new_n710));
  INV_X1    g509(.A(KEYINPUT44), .ZN(new_n711));
  AOI211_X1 g510(.A(new_n711), .B(new_n650), .C1(new_n523), .C2(new_n564), .ZN(new_n712));
  AND3_X1   g511(.A1(new_n515), .A2(new_n522), .A3(KEYINPUT105), .ZN(new_n713));
  AOI21_X1  g512(.A(KEYINPUT105), .B1(new_n515), .B2(new_n522), .ZN(new_n714));
  OAI21_X1  g513(.A(new_n564), .B1(new_n713), .B2(new_n714), .ZN(new_n715));
  NAND2_X1  g514(.A1(new_n715), .A2(new_n649), .ZN(new_n716));
  AOI21_X1  g515(.A(new_n712), .B1(new_n716), .B2(new_n711), .ZN(new_n717));
  AND3_X1   g516(.A1(new_n281), .A2(new_n277), .A3(new_n266), .ZN(new_n718));
  AOI21_X1  g517(.A(new_n277), .B1(new_n281), .B2(new_n266), .ZN(new_n719));
  OAI21_X1  g518(.A(KEYINPUT103), .B1(new_n718), .B2(new_n719), .ZN(new_n720));
  INV_X1    g519(.A(KEYINPUT103), .ZN(new_n721));
  NAND3_X1  g520(.A1(new_n279), .A2(new_n721), .A3(new_n282), .ZN(new_n722));
  AND2_X1   g521(.A1(new_n720), .A2(new_n722), .ZN(new_n723));
  NOR2_X1   g522(.A1(new_n606), .A2(new_n681), .ZN(new_n724));
  NAND2_X1  g523(.A1(new_n723), .A2(new_n724), .ZN(new_n725));
  XNOR2_X1  g524(.A(new_n725), .B(KEYINPUT104), .ZN(new_n726));
  NAND2_X1  g525(.A1(new_n717), .A2(new_n726), .ZN(new_n727));
  OAI21_X1  g526(.A(new_n204), .B1(new_n727), .B2(new_n487), .ZN(new_n728));
  NAND2_X1  g527(.A1(new_n710), .A2(new_n728), .ZN(G1328gat));
  OAI21_X1  g528(.A(G36gat), .B1(new_n727), .B2(new_n689), .ZN(new_n730));
  NAND3_X1  g529(.A1(new_n708), .A2(new_n207), .A3(new_n690), .ZN(new_n731));
  NAND2_X1  g530(.A1(new_n731), .A2(KEYINPUT46), .ZN(new_n732));
  OR2_X1    g531(.A1(new_n731), .A2(KEYINPUT46), .ZN(new_n733));
  NAND3_X1  g532(.A1(new_n730), .A2(new_n732), .A3(new_n733), .ZN(new_n734));
  INV_X1    g533(.A(KEYINPUT106), .ZN(new_n735));
  XNOR2_X1  g534(.A(new_n734), .B(new_n735), .ZN(G1329gat));
  NAND3_X1  g535(.A1(new_n717), .A2(G43gat), .A3(new_n726), .ZN(new_n737));
  AND2_X1   g536(.A1(new_n708), .A2(new_n701), .ZN(new_n738));
  OAI22_X1  g537(.A1(new_n737), .A2(new_n528), .B1(G43gat), .B2(new_n738), .ZN(new_n739));
  XNOR2_X1  g538(.A(new_n739), .B(KEYINPUT47), .ZN(G1330gat));
  NAND2_X1  g539(.A1(new_n515), .A2(new_n522), .ZN(new_n741));
  INV_X1    g540(.A(KEYINPUT105), .ZN(new_n742));
  NAND2_X1  g541(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  NAND3_X1  g542(.A1(new_n515), .A2(new_n522), .A3(KEYINPUT105), .ZN(new_n744));
  AOI22_X1  g543(.A1(new_n526), .A2(new_n527), .B1(new_n562), .B2(new_n514), .ZN(new_n745));
  AOI22_X1  g544(.A1(new_n743), .A2(new_n744), .B1(new_n561), .B2(new_n745), .ZN(new_n746));
  OAI21_X1  g545(.A(new_n711), .B1(new_n746), .B2(new_n650), .ZN(new_n747));
  INV_X1    g546(.A(new_n712), .ZN(new_n748));
  NAND4_X1  g547(.A1(new_n747), .A2(new_n748), .A3(new_n562), .A4(new_n726), .ZN(new_n749));
  NAND2_X1  g548(.A1(new_n749), .A2(G50gat), .ZN(new_n750));
  INV_X1    g549(.A(G50gat), .ZN(new_n751));
  NAND3_X1  g550(.A1(new_n708), .A2(new_n751), .A3(new_n562), .ZN(new_n752));
  NAND2_X1  g551(.A1(new_n750), .A2(new_n752), .ZN(new_n753));
  XOR2_X1   g552(.A(KEYINPUT107), .B(KEYINPUT48), .Z(new_n754));
  NAND2_X1  g553(.A1(new_n753), .A2(new_n754), .ZN(new_n755));
  NAND2_X1  g554(.A1(new_n749), .A2(KEYINPUT108), .ZN(new_n756));
  INV_X1    g555(.A(KEYINPUT108), .ZN(new_n757));
  NAND4_X1  g556(.A1(new_n717), .A2(new_n757), .A3(new_n562), .A4(new_n726), .ZN(new_n758));
  NAND3_X1  g557(.A1(new_n756), .A2(new_n758), .A3(G50gat), .ZN(new_n759));
  AND2_X1   g558(.A1(new_n752), .A2(KEYINPUT48), .ZN(new_n760));
  AND3_X1   g559(.A1(new_n759), .A2(KEYINPUT109), .A3(new_n760), .ZN(new_n761));
  AOI21_X1  g560(.A(KEYINPUT109), .B1(new_n759), .B2(new_n760), .ZN(new_n762));
  OAI21_X1  g561(.A(new_n755), .B1(new_n761), .B2(new_n762), .ZN(G1331gat));
  NOR3_X1   g562(.A1(new_n723), .A2(new_n651), .A3(new_n680), .ZN(new_n764));
  XOR2_X1   g563(.A(new_n764), .B(KEYINPUT110), .Z(new_n765));
  NOR2_X1   g564(.A1(new_n765), .A2(new_n746), .ZN(new_n766));
  NAND2_X1  g565(.A1(new_n766), .A2(new_n558), .ZN(new_n767));
  XNOR2_X1  g566(.A(new_n767), .B(G57gat), .ZN(G1332gat));
  NAND2_X1  g567(.A1(new_n766), .A2(new_n690), .ZN(new_n769));
  OAI21_X1  g568(.A(new_n769), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n770));
  XOR2_X1   g569(.A(KEYINPUT49), .B(G64gat), .Z(new_n771));
  OAI21_X1  g570(.A(new_n770), .B1(new_n769), .B2(new_n771), .ZN(G1333gat));
  INV_X1    g571(.A(new_n528), .ZN(new_n773));
  AND3_X1   g572(.A1(new_n766), .A2(G71gat), .A3(new_n773), .ZN(new_n774));
  AOI21_X1  g573(.A(G71gat), .B1(new_n766), .B2(new_n701), .ZN(new_n775));
  NOR2_X1   g574(.A1(new_n774), .A2(new_n775), .ZN(new_n776));
  XOR2_X1   g575(.A(new_n776), .B(KEYINPUT50), .Z(G1334gat));
  NAND2_X1  g576(.A1(new_n766), .A2(new_n562), .ZN(new_n778));
  XOR2_X1   g577(.A(KEYINPUT111), .B(G78gat), .Z(new_n779));
  XNOR2_X1  g578(.A(new_n778), .B(new_n779), .ZN(G1335gat));
  NOR2_X1   g579(.A1(new_n723), .A2(new_n606), .ZN(new_n781));
  NAND3_X1  g580(.A1(new_n717), .A2(new_n681), .A3(new_n781), .ZN(new_n782));
  OAI21_X1  g581(.A(G85gat), .B1(new_n782), .B2(new_n487), .ZN(new_n783));
  NAND3_X1  g582(.A1(new_n715), .A2(new_n649), .A3(new_n781), .ZN(new_n784));
  INV_X1    g583(.A(KEYINPUT51), .ZN(new_n785));
  XNOR2_X1  g584(.A(new_n784), .B(new_n785), .ZN(new_n786));
  NAND3_X1  g585(.A1(new_n558), .A2(new_n455), .A3(new_n681), .ZN(new_n787));
  XNOR2_X1  g586(.A(new_n787), .B(KEYINPUT112), .ZN(new_n788));
  NAND2_X1  g587(.A1(new_n786), .A2(new_n788), .ZN(new_n789));
  NAND2_X1  g588(.A1(new_n783), .A2(new_n789), .ZN(G1336gat));
  NAND4_X1  g589(.A1(new_n717), .A2(new_n690), .A3(new_n681), .A4(new_n781), .ZN(new_n791));
  NAND2_X1  g590(.A1(new_n791), .A2(G92gat), .ZN(new_n792));
  NOR3_X1   g591(.A1(new_n689), .A2(G92gat), .A3(new_n680), .ZN(new_n793));
  NAND2_X1  g592(.A1(new_n786), .A2(new_n793), .ZN(new_n794));
  INV_X1    g593(.A(KEYINPUT52), .ZN(new_n795));
  NAND3_X1  g594(.A1(new_n792), .A2(new_n794), .A3(new_n795), .ZN(new_n796));
  XNOR2_X1  g595(.A(KEYINPUT113), .B(KEYINPUT51), .ZN(new_n797));
  NAND2_X1  g596(.A1(new_n784), .A2(new_n797), .ZN(new_n798));
  INV_X1    g597(.A(KEYINPUT114), .ZN(new_n799));
  NAND2_X1  g598(.A1(new_n798), .A2(new_n799), .ZN(new_n800));
  NAND3_X1  g599(.A1(new_n784), .A2(KEYINPUT114), .A3(new_n797), .ZN(new_n801));
  OAI211_X1 g600(.A(new_n800), .B(new_n801), .C1(new_n785), .C2(new_n784), .ZN(new_n802));
  AOI22_X1  g601(.A1(new_n802), .A2(new_n793), .B1(G92gat), .B2(new_n791), .ZN(new_n803));
  OAI21_X1  g602(.A(new_n796), .B1(new_n803), .B2(new_n795), .ZN(G1337gat));
  XOR2_X1   g603(.A(KEYINPUT115), .B(G99gat), .Z(new_n805));
  INV_X1    g604(.A(new_n805), .ZN(new_n806));
  NAND4_X1  g605(.A1(new_n786), .A2(new_n701), .A3(new_n681), .A4(new_n806), .ZN(new_n807));
  OAI21_X1  g606(.A(new_n805), .B1(new_n782), .B2(new_n528), .ZN(new_n808));
  NAND2_X1  g607(.A1(new_n807), .A2(new_n808), .ZN(new_n809));
  NAND2_X1  g608(.A1(new_n809), .A2(KEYINPUT116), .ZN(new_n810));
  INV_X1    g609(.A(KEYINPUT116), .ZN(new_n811));
  NAND3_X1  g610(.A1(new_n807), .A2(new_n808), .A3(new_n811), .ZN(new_n812));
  NAND2_X1  g611(.A1(new_n810), .A2(new_n812), .ZN(G1338gat));
  NAND4_X1  g612(.A1(new_n717), .A2(new_n562), .A3(new_n681), .A4(new_n781), .ZN(new_n814));
  NAND2_X1  g613(.A1(new_n814), .A2(G106gat), .ZN(new_n815));
  NOR3_X1   g614(.A1(new_n441), .A2(G106gat), .A3(new_n680), .ZN(new_n816));
  NAND2_X1  g615(.A1(new_n786), .A2(new_n816), .ZN(new_n817));
  INV_X1    g616(.A(KEYINPUT53), .ZN(new_n818));
  NAND3_X1  g617(.A1(new_n815), .A2(new_n817), .A3(new_n818), .ZN(new_n819));
  AOI22_X1  g618(.A1(new_n802), .A2(new_n816), .B1(G106gat), .B2(new_n814), .ZN(new_n820));
  OAI21_X1  g619(.A(new_n819), .B1(new_n820), .B2(new_n818), .ZN(G1339gat));
  NOR2_X1   g620(.A1(new_n690), .A2(new_n487), .ZN(new_n822));
  INV_X1    g621(.A(new_n822), .ZN(new_n823));
  INV_X1    g622(.A(new_n606), .ZN(new_n824));
  INV_X1    g623(.A(KEYINPUT118), .ZN(new_n825));
  INV_X1    g624(.A(KEYINPUT117), .ZN(new_n826));
  INV_X1    g625(.A(KEYINPUT10), .ZN(new_n827));
  AND3_X1   g626(.A1(new_n625), .A2(new_n652), .A3(new_n626), .ZN(new_n828));
  AOI21_X1  g627(.A(new_n626), .B1(new_n625), .B2(new_n652), .ZN(new_n829));
  NOR3_X1   g628(.A1(new_n584), .A2(new_n828), .A3(new_n829), .ZN(new_n830));
  AND2_X1   g629(.A1(new_n614), .A2(new_n621), .ZN(new_n831));
  NAND4_X1  g630(.A1(new_n831), .A2(new_n628), .A3(new_n627), .A4(new_n624), .ZN(new_n832));
  NAND3_X1  g631(.A1(new_n625), .A2(new_n629), .A3(new_n630), .ZN(new_n833));
  AOI22_X1  g632(.A1(new_n832), .A2(new_n833), .B1(new_n661), .B2(new_n577), .ZN(new_n834));
  OAI21_X1  g633(.A(new_n827), .B1(new_n830), .B2(new_n834), .ZN(new_n835));
  OR2_X1    g634(.A1(new_n666), .A2(new_n584), .ZN(new_n836));
  AOI21_X1  g635(.A(new_n671), .B1(new_n835), .B2(new_n836), .ZN(new_n837));
  INV_X1    g636(.A(KEYINPUT54), .ZN(new_n838));
  AOI21_X1  g637(.A(new_n678), .B1(new_n837), .B2(new_n838), .ZN(new_n839));
  NAND3_X1  g638(.A1(new_n835), .A2(new_n671), .A3(new_n836), .ZN(new_n840));
  NAND3_X1  g639(.A1(new_n670), .A2(new_n840), .A3(KEYINPUT54), .ZN(new_n841));
  NAND2_X1  g640(.A1(new_n839), .A2(new_n841), .ZN(new_n842));
  INV_X1    g641(.A(KEYINPUT55), .ZN(new_n843));
  AOI21_X1  g642(.A(new_n826), .B1(new_n842), .B2(new_n843), .ZN(new_n844));
  AOI211_X1 g643(.A(KEYINPUT117), .B(KEYINPUT55), .C1(new_n839), .C2(new_n841), .ZN(new_n845));
  NOR2_X1   g644(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  NAND3_X1  g645(.A1(new_n839), .A2(KEYINPUT55), .A3(new_n841), .ZN(new_n847));
  AND2_X1   g646(.A1(new_n847), .A2(new_n679), .ZN(new_n848));
  AOI21_X1  g647(.A(new_n825), .B1(new_n846), .B2(new_n848), .ZN(new_n849));
  AND3_X1   g648(.A1(new_n670), .A2(new_n840), .A3(KEYINPUT54), .ZN(new_n850));
  OAI21_X1  g649(.A(new_n676), .B1(new_n670), .B2(KEYINPUT54), .ZN(new_n851));
  OAI21_X1  g650(.A(new_n843), .B1(new_n850), .B2(new_n851), .ZN(new_n852));
  NAND2_X1  g651(.A1(new_n852), .A2(KEYINPUT117), .ZN(new_n853));
  NAND3_X1  g652(.A1(new_n842), .A2(new_n826), .A3(new_n843), .ZN(new_n854));
  AND4_X1   g653(.A1(new_n825), .A2(new_n848), .A3(new_n853), .A4(new_n854), .ZN(new_n855));
  OAI211_X1 g654(.A(new_n720), .B(new_n722), .C1(new_n849), .C2(new_n855), .ZN(new_n856));
  NOR2_X1   g655(.A1(new_n256), .A2(new_n259), .ZN(new_n857));
  AOI21_X1  g656(.A(new_n257), .B1(new_n264), .B2(new_n253), .ZN(new_n858));
  OAI21_X1  g657(.A(new_n275), .B1(new_n857), .B2(new_n858), .ZN(new_n859));
  NAND3_X1  g658(.A1(new_n282), .A2(new_n681), .A3(new_n859), .ZN(new_n860));
  AOI21_X1  g659(.A(new_n649), .B1(new_n856), .B2(new_n860), .ZN(new_n861));
  NOR2_X1   g660(.A1(new_n849), .A2(new_n855), .ZN(new_n862));
  NAND3_X1  g661(.A1(new_n649), .A2(new_n282), .A3(new_n859), .ZN(new_n863));
  NOR2_X1   g662(.A1(new_n862), .A2(new_n863), .ZN(new_n864));
  OAI21_X1  g663(.A(new_n824), .B1(new_n861), .B2(new_n864), .ZN(new_n865));
  NAND2_X1  g664(.A1(new_n720), .A2(new_n722), .ZN(new_n866));
  NAND4_X1  g665(.A1(new_n866), .A2(new_n606), .A3(new_n650), .A4(new_n680), .ZN(new_n867));
  AOI21_X1  g666(.A(new_n823), .B1(new_n865), .B2(new_n867), .ZN(new_n868));
  AND2_X1   g667(.A1(new_n441), .A2(new_n520), .ZN(new_n869));
  NAND2_X1  g668(.A1(new_n868), .A2(new_n869), .ZN(new_n870));
  XOR2_X1   g669(.A(new_n870), .B(KEYINPUT119), .Z(new_n871));
  NAND2_X1  g670(.A1(new_n320), .A2(new_n321), .ZN(new_n872));
  NAND3_X1  g671(.A1(new_n871), .A2(new_n872), .A3(new_n723), .ZN(new_n873));
  INV_X1    g672(.A(new_n453), .ZN(new_n874));
  NAND2_X1  g673(.A1(new_n868), .A2(new_n874), .ZN(new_n875));
  OAI21_X1  g674(.A(G113gat), .B1(new_n875), .B2(new_n284), .ZN(new_n876));
  NAND2_X1  g675(.A1(new_n873), .A2(new_n876), .ZN(G1340gat));
  NAND3_X1  g676(.A1(new_n871), .A2(new_n309), .A3(new_n681), .ZN(new_n878));
  OAI21_X1  g677(.A(G120gat), .B1(new_n875), .B2(new_n680), .ZN(new_n879));
  NAND2_X1  g678(.A1(new_n878), .A2(new_n879), .ZN(G1341gat));
  INV_X1    g679(.A(new_n316), .ZN(new_n881));
  NOR3_X1   g680(.A1(new_n875), .A2(new_n881), .A3(new_n824), .ZN(new_n882));
  XNOR2_X1  g681(.A(new_n882), .B(KEYINPUT120), .ZN(new_n883));
  NAND3_X1  g682(.A1(new_n868), .A2(new_n869), .A3(new_n606), .ZN(new_n884));
  AOI21_X1  g683(.A(new_n883), .B1(new_n881), .B2(new_n884), .ZN(G1342gat));
  NOR3_X1   g684(.A1(new_n870), .A2(G134gat), .A3(new_n650), .ZN(new_n886));
  XNOR2_X1  g685(.A(new_n886), .B(KEYINPUT56), .ZN(new_n887));
  OAI21_X1  g686(.A(G134gat), .B1(new_n875), .B2(new_n650), .ZN(new_n888));
  NAND2_X1  g687(.A1(new_n887), .A2(new_n888), .ZN(G1343gat));
  AOI21_X1  g688(.A(new_n441), .B1(new_n865), .B2(new_n867), .ZN(new_n890));
  NAND2_X1  g689(.A1(new_n822), .A2(new_n528), .ZN(new_n891));
  INV_X1    g690(.A(new_n891), .ZN(new_n892));
  NAND2_X1  g691(.A1(new_n890), .A2(new_n892), .ZN(new_n893));
  NOR3_X1   g692(.A1(new_n893), .A2(G141gat), .A3(new_n284), .ZN(new_n894));
  INV_X1    g693(.A(new_n890), .ZN(new_n895));
  INV_X1    g694(.A(KEYINPUT57), .ZN(new_n896));
  NAND2_X1  g695(.A1(new_n895), .A2(new_n896), .ZN(new_n897));
  NAND3_X1  g696(.A1(new_n283), .A2(new_n848), .A3(new_n852), .ZN(new_n898));
  AOI21_X1  g697(.A(new_n649), .B1(new_n898), .B2(new_n860), .ZN(new_n899));
  OAI21_X1  g698(.A(new_n824), .B1(new_n899), .B2(new_n864), .ZN(new_n900));
  NAND2_X1  g699(.A1(new_n900), .A2(new_n867), .ZN(new_n901));
  NAND3_X1  g700(.A1(new_n901), .A2(KEYINPUT57), .A3(new_n562), .ZN(new_n902));
  AOI21_X1  g701(.A(new_n891), .B1(new_n897), .B2(new_n902), .ZN(new_n903));
  NAND2_X1  g702(.A1(new_n903), .A2(new_n723), .ZN(new_n904));
  AOI21_X1  g703(.A(new_n894), .B1(new_n904), .B2(G141gat), .ZN(new_n905));
  INV_X1    g704(.A(KEYINPUT58), .ZN(new_n906));
  AOI21_X1  g705(.A(new_n379), .B1(new_n903), .B2(new_n283), .ZN(new_n907));
  OR2_X1    g706(.A1(new_n894), .A2(KEYINPUT58), .ZN(new_n908));
  OAI22_X1  g707(.A1(new_n905), .A2(new_n906), .B1(new_n907), .B2(new_n908), .ZN(G1344gat));
  INV_X1    g708(.A(new_n893), .ZN(new_n910));
  NAND3_X1  g709(.A1(new_n910), .A2(new_n381), .A3(new_n681), .ZN(new_n911));
  AOI211_X1 g710(.A(KEYINPUT59), .B(new_n381), .C1(new_n903), .C2(new_n681), .ZN(new_n912));
  INV_X1    g711(.A(KEYINPUT59), .ZN(new_n913));
  OAI21_X1  g712(.A(new_n860), .B1(new_n866), .B2(new_n862), .ZN(new_n914));
  AOI21_X1  g713(.A(new_n864), .B1(new_n914), .B2(new_n650), .ZN(new_n915));
  OAI21_X1  g714(.A(new_n867), .B1(new_n915), .B2(new_n606), .ZN(new_n916));
  AOI21_X1  g715(.A(new_n896), .B1(new_n916), .B2(new_n562), .ZN(new_n917));
  NAND3_X1  g716(.A1(new_n682), .A2(new_n284), .A3(new_n683), .ZN(new_n918));
  NAND2_X1  g717(.A1(new_n846), .A2(new_n848), .ZN(new_n919));
  NOR2_X1   g718(.A1(new_n863), .A2(new_n919), .ZN(new_n920));
  OAI21_X1  g719(.A(new_n824), .B1(new_n899), .B2(new_n920), .ZN(new_n921));
  AOI211_X1 g720(.A(KEYINPUT57), .B(new_n441), .C1(new_n918), .C2(new_n921), .ZN(new_n922));
  NOR2_X1   g721(.A1(new_n917), .A2(new_n922), .ZN(new_n923));
  NAND3_X1  g722(.A1(new_n923), .A2(new_n681), .A3(new_n892), .ZN(new_n924));
  AOI21_X1  g723(.A(new_n913), .B1(new_n924), .B2(G148gat), .ZN(new_n925));
  OAI21_X1  g724(.A(new_n911), .B1(new_n912), .B2(new_n925), .ZN(G1345gat));
  AOI21_X1  g725(.A(G155gat), .B1(new_n910), .B2(new_n606), .ZN(new_n927));
  NOR2_X1   g726(.A1(new_n824), .A2(new_n372), .ZN(new_n928));
  AOI21_X1  g727(.A(new_n927), .B1(new_n903), .B2(new_n928), .ZN(G1346gat));
  NOR3_X1   g728(.A1(new_n893), .A2(G162gat), .A3(new_n650), .ZN(new_n930));
  XNOR2_X1  g729(.A(new_n930), .B(KEYINPUT121), .ZN(new_n931));
  AND2_X1   g730(.A1(new_n903), .A2(new_n649), .ZN(new_n932));
  OAI21_X1  g731(.A(new_n931), .B1(new_n373), .B2(new_n932), .ZN(G1347gat));
  NOR2_X1   g732(.A1(new_n689), .A2(new_n558), .ZN(new_n934));
  AND2_X1   g733(.A1(new_n916), .A2(new_n934), .ZN(new_n935));
  NAND2_X1  g734(.A1(new_n935), .A2(new_n874), .ZN(new_n936));
  OAI21_X1  g735(.A(G169gat), .B1(new_n936), .B2(new_n284), .ZN(new_n937));
  NAND3_X1  g736(.A1(new_n935), .A2(new_n333), .A3(new_n869), .ZN(new_n938));
  OAI21_X1  g737(.A(new_n937), .B1(new_n866), .B2(new_n938), .ZN(G1348gat));
  NOR3_X1   g738(.A1(new_n936), .A2(new_n334), .A3(new_n680), .ZN(new_n940));
  NAND3_X1  g739(.A1(new_n935), .A2(new_n869), .A3(new_n681), .ZN(new_n941));
  AOI21_X1  g740(.A(new_n940), .B1(new_n334), .B2(new_n941), .ZN(G1349gat));
  OAI21_X1  g741(.A(G183gat), .B1(new_n936), .B2(new_n824), .ZN(new_n943));
  NAND2_X1  g742(.A1(new_n935), .A2(new_n869), .ZN(new_n944));
  OAI21_X1  g743(.A(new_n606), .B1(new_n327), .B2(new_n326), .ZN(new_n945));
  OAI21_X1  g744(.A(new_n943), .B1(new_n944), .B2(new_n945), .ZN(new_n946));
  INV_X1    g745(.A(KEYINPUT60), .ZN(new_n947));
  NOR2_X1   g746(.A1(new_n947), .A2(KEYINPUT122), .ZN(new_n948));
  XNOR2_X1  g747(.A(new_n946), .B(new_n948), .ZN(G1350gat));
  NAND4_X1  g748(.A1(new_n916), .A2(new_n874), .A3(new_n649), .A4(new_n934), .ZN(new_n950));
  NAND2_X1  g749(.A1(new_n950), .A2(G190gat), .ZN(new_n951));
  NAND2_X1  g750(.A1(new_n951), .A2(KEYINPUT123), .ZN(new_n952));
  INV_X1    g751(.A(KEYINPUT123), .ZN(new_n953));
  NAND3_X1  g752(.A1(new_n950), .A2(new_n953), .A3(G190gat), .ZN(new_n954));
  NAND3_X1  g753(.A1(new_n952), .A2(KEYINPUT61), .A3(new_n954), .ZN(new_n955));
  NAND4_X1  g754(.A1(new_n935), .A2(new_n294), .A3(new_n869), .A4(new_n649), .ZN(new_n956));
  INV_X1    g755(.A(KEYINPUT61), .ZN(new_n957));
  NAND3_X1  g756(.A1(new_n951), .A2(KEYINPUT123), .A3(new_n957), .ZN(new_n958));
  NAND3_X1  g757(.A1(new_n955), .A2(new_n956), .A3(new_n958), .ZN(new_n959));
  NAND2_X1  g758(.A1(new_n959), .A2(KEYINPUT124), .ZN(new_n960));
  INV_X1    g759(.A(KEYINPUT124), .ZN(new_n961));
  NAND4_X1  g760(.A1(new_n955), .A2(new_n961), .A3(new_n956), .A4(new_n958), .ZN(new_n962));
  NAND2_X1  g761(.A1(new_n960), .A2(new_n962), .ZN(G1351gat));
  INV_X1    g762(.A(KEYINPUT126), .ZN(new_n964));
  OAI21_X1  g763(.A(new_n964), .B1(new_n917), .B2(new_n922), .ZN(new_n965));
  NAND2_X1  g764(.A1(new_n528), .A2(new_n934), .ZN(new_n966));
  INV_X1    g765(.A(new_n966), .ZN(new_n967));
  NAND2_X1  g766(.A1(new_n918), .A2(new_n921), .ZN(new_n968));
  NAND3_X1  g767(.A1(new_n968), .A2(new_n896), .A3(new_n562), .ZN(new_n969));
  OAI211_X1 g768(.A(new_n969), .B(KEYINPUT126), .C1(new_n890), .C2(new_n896), .ZN(new_n970));
  NAND4_X1  g769(.A1(new_n965), .A2(new_n283), .A3(new_n967), .A4(new_n970), .ZN(new_n971));
  NAND2_X1  g770(.A1(new_n971), .A2(G197gat), .ZN(new_n972));
  NOR3_X1   g771(.A1(new_n895), .A2(KEYINPUT125), .A3(new_n966), .ZN(new_n973));
  INV_X1    g772(.A(KEYINPUT125), .ZN(new_n974));
  AOI21_X1  g773(.A(new_n974), .B1(new_n890), .B2(new_n967), .ZN(new_n975));
  OAI211_X1 g774(.A(new_n272), .B(new_n723), .C1(new_n973), .C2(new_n975), .ZN(new_n976));
  NAND2_X1  g775(.A1(new_n972), .A2(new_n976), .ZN(new_n977));
  NAND2_X1  g776(.A1(new_n977), .A2(KEYINPUT127), .ZN(new_n978));
  INV_X1    g777(.A(KEYINPUT127), .ZN(new_n979));
  NAND3_X1  g778(.A1(new_n972), .A2(new_n979), .A3(new_n976), .ZN(new_n980));
  NAND2_X1  g779(.A1(new_n978), .A2(new_n980), .ZN(G1352gat));
  NOR3_X1   g780(.A1(new_n773), .A2(new_n441), .A3(new_n680), .ZN(new_n982));
  NAND3_X1  g781(.A1(new_n935), .A2(new_n392), .A3(new_n982), .ZN(new_n983));
  XOR2_X1   g782(.A(new_n983), .B(KEYINPUT62), .Z(new_n984));
  NAND3_X1  g783(.A1(new_n965), .A2(new_n967), .A3(new_n970), .ZN(new_n985));
  OAI21_X1  g784(.A(G204gat), .B1(new_n985), .B2(new_n680), .ZN(new_n986));
  NAND2_X1  g785(.A1(new_n984), .A2(new_n986), .ZN(G1353gat));
  NAND3_X1  g786(.A1(new_n923), .A2(new_n606), .A3(new_n967), .ZN(new_n988));
  NAND3_X1  g787(.A1(new_n988), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n989));
  INV_X1    g788(.A(new_n989), .ZN(new_n990));
  AOI21_X1  g789(.A(KEYINPUT63), .B1(new_n988), .B2(G211gat), .ZN(new_n991));
  NOR2_X1   g790(.A1(new_n973), .A2(new_n975), .ZN(new_n992));
  OR2_X1    g791(.A1(new_n824), .A2(G211gat), .ZN(new_n993));
  OAI22_X1  g792(.A1(new_n990), .A2(new_n991), .B1(new_n992), .B2(new_n993), .ZN(G1354gat));
  OAI21_X1  g793(.A(G218gat), .B1(new_n985), .B2(new_n650), .ZN(new_n995));
  OR2_X1    g794(.A1(new_n650), .A2(G218gat), .ZN(new_n996));
  OAI21_X1  g795(.A(new_n995), .B1(new_n992), .B2(new_n996), .ZN(G1355gat));
endmodule


