//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 1 0 0 0 0 0 1 0 0 1 1 0 1 0 1 1 0 0 1 0 1 1 1 0 1 1 0 1 0 0 0 1 1 0 1 0 0 1 0 0 0 1 0 0 0 1 1 0 0 1 1 0 1 0 0 0 0 0 1 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:23:53 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n677, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n692, new_n693,
    new_n694, new_n695, new_n696, new_n697, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n713, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n735, new_n736, new_n737, new_n738,
    new_n739, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n749, new_n750, new_n751, new_n752, new_n753, new_n755,
    new_n756, new_n758, new_n759, new_n760, new_n761, new_n762, new_n763,
    new_n764, new_n765, new_n767, new_n768, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n776, new_n777, new_n778, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n801, new_n802, new_n803,
    new_n804, new_n805, new_n806, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n919, new_n920,
    new_n921, new_n922, new_n923, new_n924, new_n925, new_n926, new_n927,
    new_n928, new_n929, new_n930, new_n931, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n939, new_n940, new_n942, new_n943,
    new_n944, new_n945, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n971, new_n972, new_n973,
    new_n974, new_n975, new_n976, new_n977, new_n978, new_n979, new_n980,
    new_n981, new_n982, new_n983, new_n984, new_n985;
  INV_X1    g000(.A(G217), .ZN(new_n187));
  XOR2_X1   g001(.A(KEYINPUT78), .B(G902), .Z(new_n188));
  AOI21_X1  g002(.A(new_n187), .B1(new_n188), .B2(G234), .ZN(new_n189));
  INV_X1    g003(.A(new_n188), .ZN(new_n190));
  INV_X1    g004(.A(G140), .ZN(new_n191));
  NAND2_X1  g005(.A1(new_n191), .A2(G125), .ZN(new_n192));
  INV_X1    g006(.A(G125), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n193), .A2(G140), .ZN(new_n194));
  NAND3_X1  g008(.A1(new_n192), .A2(new_n194), .A3(KEYINPUT16), .ZN(new_n195));
  OR3_X1    g009(.A1(new_n193), .A2(KEYINPUT16), .A3(G140), .ZN(new_n196));
  NAND3_X1  g010(.A1(new_n195), .A2(new_n196), .A3(G146), .ZN(new_n197));
  INV_X1    g011(.A(KEYINPUT80), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n197), .A2(new_n198), .ZN(new_n199));
  NAND4_X1  g013(.A1(new_n195), .A2(new_n196), .A3(KEYINPUT80), .A4(G146), .ZN(new_n200));
  AND2_X1   g014(.A1(new_n195), .A2(new_n196), .ZN(new_n201));
  OAI211_X1 g015(.A(new_n199), .B(new_n200), .C1(G146), .C2(new_n201), .ZN(new_n202));
  INV_X1    g016(.A(KEYINPUT23), .ZN(new_n203));
  INV_X1    g017(.A(G119), .ZN(new_n204));
  OAI21_X1  g018(.A(new_n203), .B1(new_n204), .B2(G128), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n204), .A2(G128), .ZN(new_n206));
  INV_X1    g020(.A(G128), .ZN(new_n207));
  NAND3_X1  g021(.A1(new_n207), .A2(KEYINPUT23), .A3(G119), .ZN(new_n208));
  NAND3_X1  g022(.A1(new_n205), .A2(new_n206), .A3(new_n208), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n209), .A2(G110), .ZN(new_n210));
  XNOR2_X1  g024(.A(KEYINPUT24), .B(G110), .ZN(new_n211));
  OAI21_X1  g025(.A(KEYINPUT79), .B1(new_n204), .B2(G128), .ZN(new_n212));
  INV_X1    g026(.A(KEYINPUT79), .ZN(new_n213));
  NAND3_X1  g027(.A1(new_n213), .A2(new_n207), .A3(G119), .ZN(new_n214));
  NAND3_X1  g028(.A1(new_n212), .A2(new_n214), .A3(new_n206), .ZN(new_n215));
  OAI211_X1 g029(.A(new_n202), .B(new_n210), .C1(new_n211), .C2(new_n215), .ZN(new_n216));
  INV_X1    g030(.A(KEYINPUT82), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n197), .A2(new_n217), .ZN(new_n218));
  NAND4_X1  g032(.A1(new_n195), .A2(new_n196), .A3(KEYINPUT82), .A4(G146), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n218), .A2(new_n219), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n192), .A2(new_n194), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n215), .A2(new_n211), .ZN(new_n222));
  INV_X1    g036(.A(KEYINPUT81), .ZN(new_n223));
  INV_X1    g037(.A(G110), .ZN(new_n224));
  NAND4_X1  g038(.A1(new_n205), .A2(new_n208), .A3(new_n224), .A4(new_n206), .ZN(new_n225));
  AND3_X1   g039(.A1(new_n222), .A2(new_n223), .A3(new_n225), .ZN(new_n226));
  AOI21_X1  g040(.A(new_n223), .B1(new_n222), .B2(new_n225), .ZN(new_n227));
  OAI221_X1 g041(.A(new_n220), .B1(G146), .B2(new_n221), .C1(new_n226), .C2(new_n227), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n216), .A2(new_n228), .ZN(new_n229));
  XNOR2_X1  g043(.A(KEYINPUT22), .B(G137), .ZN(new_n230));
  XNOR2_X1  g044(.A(new_n230), .B(KEYINPUT83), .ZN(new_n231));
  INV_X1    g045(.A(G953), .ZN(new_n232));
  AND3_X1   g046(.A1(new_n232), .A2(G221), .A3(G234), .ZN(new_n233));
  XOR2_X1   g047(.A(new_n231), .B(new_n233), .Z(new_n234));
  INV_X1    g048(.A(new_n234), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n229), .A2(new_n235), .ZN(new_n236));
  NAND3_X1  g050(.A1(new_n216), .A2(new_n228), .A3(new_n234), .ZN(new_n237));
  AOI21_X1  g051(.A(new_n190), .B1(new_n236), .B2(new_n237), .ZN(new_n238));
  INV_X1    g052(.A(KEYINPUT84), .ZN(new_n239));
  NOR3_X1   g053(.A1(new_n238), .A2(new_n239), .A3(KEYINPUT25), .ZN(new_n240));
  INV_X1    g054(.A(KEYINPUT25), .ZN(new_n241));
  INV_X1    g055(.A(new_n237), .ZN(new_n242));
  AOI21_X1  g056(.A(new_n234), .B1(new_n216), .B2(new_n228), .ZN(new_n243));
  OAI21_X1  g057(.A(new_n188), .B1(new_n242), .B2(new_n243), .ZN(new_n244));
  AOI21_X1  g058(.A(new_n241), .B1(new_n244), .B2(KEYINPUT84), .ZN(new_n245));
  OAI21_X1  g059(.A(new_n189), .B1(new_n240), .B2(new_n245), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n236), .A2(new_n237), .ZN(new_n247));
  NOR2_X1   g061(.A1(new_n189), .A2(G902), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n247), .A2(new_n248), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n246), .A2(new_n249), .ZN(new_n250));
  INV_X1    g064(.A(G116), .ZN(new_n251));
  NOR2_X1   g065(.A1(new_n251), .A2(G119), .ZN(new_n252));
  INV_X1    g066(.A(new_n252), .ZN(new_n253));
  AND3_X1   g067(.A1(new_n251), .A2(KEYINPUT68), .A3(G119), .ZN(new_n254));
  AOI21_X1  g068(.A(KEYINPUT68), .B1(new_n251), .B2(G119), .ZN(new_n255));
  OAI21_X1  g069(.A(new_n253), .B1(new_n254), .B2(new_n255), .ZN(new_n256));
  AND2_X1   g070(.A1(KEYINPUT2), .A2(G113), .ZN(new_n257));
  NOR2_X1   g071(.A1(KEYINPUT2), .A2(G113), .ZN(new_n258));
  NOR2_X1   g072(.A1(new_n257), .A2(new_n258), .ZN(new_n259));
  INV_X1    g073(.A(new_n259), .ZN(new_n260));
  AOI21_X1  g074(.A(KEYINPUT69), .B1(new_n256), .B2(new_n260), .ZN(new_n261));
  INV_X1    g075(.A(KEYINPUT68), .ZN(new_n262));
  OAI21_X1  g076(.A(new_n262), .B1(new_n204), .B2(G116), .ZN(new_n263));
  NAND3_X1  g077(.A1(new_n251), .A2(KEYINPUT68), .A3(G119), .ZN(new_n264));
  AOI21_X1  g078(.A(new_n252), .B1(new_n263), .B2(new_n264), .ZN(new_n265));
  INV_X1    g079(.A(KEYINPUT69), .ZN(new_n266));
  NOR3_X1   g080(.A1(new_n265), .A2(new_n266), .A3(new_n259), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n263), .A2(new_n264), .ZN(new_n268));
  AND4_X1   g082(.A1(KEYINPUT70), .A2(new_n268), .A3(new_n259), .A4(new_n253), .ZN(new_n269));
  AOI21_X1  g083(.A(KEYINPUT70), .B1(new_n265), .B2(new_n259), .ZN(new_n270));
  OAI22_X1  g084(.A1(new_n261), .A2(new_n267), .B1(new_n269), .B2(new_n270), .ZN(new_n271));
  INV_X1    g085(.A(KEYINPUT71), .ZN(new_n272));
  NAND2_X1  g086(.A1(new_n271), .A2(new_n272), .ZN(new_n273));
  INV_X1    g087(.A(G143), .ZN(new_n274));
  OAI21_X1  g088(.A(KEYINPUT1), .B1(new_n274), .B2(G146), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n275), .A2(G128), .ZN(new_n276));
  INV_X1    g090(.A(G146), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n277), .A2(G143), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n274), .A2(G146), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n278), .A2(new_n279), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n276), .A2(new_n280), .ZN(new_n281));
  NOR2_X1   g095(.A1(new_n207), .A2(KEYINPUT1), .ZN(new_n282));
  INV_X1    g096(.A(KEYINPUT64), .ZN(new_n283));
  AOI21_X1  g097(.A(new_n283), .B1(new_n274), .B2(G146), .ZN(new_n284));
  NOR3_X1   g098(.A1(new_n277), .A2(KEYINPUT64), .A3(G143), .ZN(new_n285));
  OAI211_X1 g099(.A(new_n278), .B(new_n282), .C1(new_n284), .C2(new_n285), .ZN(new_n286));
  NOR2_X1   g100(.A1(new_n286), .A2(KEYINPUT66), .ZN(new_n287));
  INV_X1    g101(.A(KEYINPUT66), .ZN(new_n288));
  OAI21_X1  g102(.A(KEYINPUT64), .B1(new_n277), .B2(G143), .ZN(new_n289));
  NAND3_X1  g103(.A1(new_n283), .A2(new_n274), .A3(G146), .ZN(new_n290));
  AOI22_X1  g104(.A1(new_n289), .A2(new_n290), .B1(G143), .B2(new_n277), .ZN(new_n291));
  AOI21_X1  g105(.A(new_n288), .B1(new_n291), .B2(new_n282), .ZN(new_n292));
  OAI21_X1  g106(.A(new_n281), .B1(new_n287), .B2(new_n292), .ZN(new_n293));
  INV_X1    g107(.A(KEYINPUT11), .ZN(new_n294));
  INV_X1    g108(.A(G134), .ZN(new_n295));
  OAI21_X1  g109(.A(new_n294), .B1(new_n295), .B2(G137), .ZN(new_n296));
  INV_X1    g110(.A(G137), .ZN(new_n297));
  NAND3_X1  g111(.A1(new_n297), .A2(KEYINPUT11), .A3(G134), .ZN(new_n298));
  INV_X1    g112(.A(G131), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n295), .A2(G137), .ZN(new_n300));
  NAND4_X1  g114(.A1(new_n296), .A2(new_n298), .A3(new_n299), .A4(new_n300), .ZN(new_n301));
  NOR2_X1   g115(.A1(new_n295), .A2(G137), .ZN(new_n302));
  NOR2_X1   g116(.A1(new_n297), .A2(G134), .ZN(new_n303));
  OAI21_X1  g117(.A(G131), .B1(new_n302), .B2(new_n303), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n301), .A2(new_n304), .ZN(new_n305));
  INV_X1    g119(.A(new_n305), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n293), .A2(new_n306), .ZN(new_n307));
  AND2_X1   g121(.A1(KEYINPUT0), .A2(G128), .ZN(new_n308));
  NOR2_X1   g122(.A1(KEYINPUT0), .A2(G128), .ZN(new_n309));
  NOR2_X1   g123(.A1(new_n308), .A2(new_n309), .ZN(new_n310));
  AOI22_X1  g124(.A1(new_n291), .A2(new_n308), .B1(new_n310), .B2(new_n280), .ZN(new_n311));
  NAND3_X1  g125(.A1(new_n296), .A2(new_n300), .A3(new_n298), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n312), .A2(G131), .ZN(new_n313));
  NAND2_X1  g127(.A1(new_n313), .A2(new_n301), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n311), .A2(new_n314), .ZN(new_n315));
  NAND3_X1  g129(.A1(new_n268), .A2(new_n259), .A3(new_n253), .ZN(new_n316));
  INV_X1    g130(.A(KEYINPUT70), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n316), .A2(new_n317), .ZN(new_n318));
  NAND3_X1  g132(.A1(new_n265), .A2(KEYINPUT70), .A3(new_n259), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n318), .A2(new_n319), .ZN(new_n320));
  NAND3_X1  g134(.A1(new_n256), .A2(KEYINPUT69), .A3(new_n260), .ZN(new_n321));
  OAI21_X1  g135(.A(new_n266), .B1(new_n265), .B2(new_n259), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n321), .A2(new_n322), .ZN(new_n323));
  NAND3_X1  g137(.A1(new_n320), .A2(new_n323), .A3(KEYINPUT71), .ZN(new_n324));
  NAND4_X1  g138(.A1(new_n273), .A2(new_n307), .A3(new_n315), .A4(new_n324), .ZN(new_n325));
  INV_X1    g139(.A(KEYINPUT72), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n325), .A2(new_n326), .ZN(new_n327));
  AOI22_X1  g141(.A1(new_n293), .A2(new_n306), .B1(new_n314), .B2(new_n311), .ZN(new_n328));
  NAND4_X1  g142(.A1(new_n328), .A2(KEYINPUT72), .A3(new_n273), .A4(new_n324), .ZN(new_n329));
  XNOR2_X1  g143(.A(KEYINPUT73), .B(KEYINPUT27), .ZN(new_n330));
  XNOR2_X1  g144(.A(new_n330), .B(KEYINPUT74), .ZN(new_n331));
  NOR2_X1   g145(.A1(G237), .A2(G953), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n332), .A2(G210), .ZN(new_n333));
  XNOR2_X1  g147(.A(new_n331), .B(new_n333), .ZN(new_n334));
  XNOR2_X1  g148(.A(KEYINPUT26), .B(G101), .ZN(new_n335));
  XNOR2_X1  g149(.A(new_n334), .B(new_n335), .ZN(new_n336));
  NAND3_X1  g150(.A1(new_n327), .A2(new_n329), .A3(new_n336), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n286), .A2(KEYINPUT66), .ZN(new_n338));
  NAND3_X1  g152(.A1(new_n291), .A2(new_n288), .A3(new_n282), .ZN(new_n339));
  AOI22_X1  g153(.A1(new_n338), .A2(new_n339), .B1(new_n280), .B2(new_n276), .ZN(new_n340));
  OAI211_X1 g154(.A(KEYINPUT30), .B(new_n315), .C1(new_n340), .C2(new_n305), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n341), .A2(new_n271), .ZN(new_n342));
  INV_X1    g156(.A(KEYINPUT65), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n305), .A2(new_n343), .ZN(new_n344));
  NAND3_X1  g158(.A1(new_n301), .A2(new_n304), .A3(KEYINPUT65), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n344), .A2(new_n345), .ZN(new_n346));
  OAI21_X1  g160(.A(KEYINPUT67), .B1(new_n340), .B2(new_n346), .ZN(new_n347));
  INV_X1    g161(.A(KEYINPUT67), .ZN(new_n348));
  AND3_X1   g162(.A1(new_n301), .A2(new_n304), .A3(KEYINPUT65), .ZN(new_n349));
  AOI21_X1  g163(.A(KEYINPUT65), .B1(new_n301), .B2(new_n304), .ZN(new_n350));
  NOR2_X1   g164(.A1(new_n349), .A2(new_n350), .ZN(new_n351));
  NAND3_X1  g165(.A1(new_n293), .A2(new_n348), .A3(new_n351), .ZN(new_n352));
  NAND3_X1  g166(.A1(new_n347), .A2(new_n352), .A3(new_n315), .ZN(new_n353));
  INV_X1    g167(.A(KEYINPUT30), .ZN(new_n354));
  AOI21_X1  g168(.A(new_n342), .B1(new_n353), .B2(new_n354), .ZN(new_n355));
  OAI21_X1  g169(.A(KEYINPUT31), .B1(new_n337), .B2(new_n355), .ZN(new_n356));
  NOR3_X1   g170(.A1(new_n337), .A2(KEYINPUT31), .A3(new_n355), .ZN(new_n357));
  INV_X1    g171(.A(KEYINPUT75), .ZN(new_n358));
  OAI21_X1  g172(.A(new_n356), .B1(new_n357), .B2(new_n358), .ZN(new_n359));
  AND2_X1   g173(.A1(new_n327), .A2(new_n329), .ZN(new_n360));
  INV_X1    g174(.A(new_n355), .ZN(new_n361));
  NAND3_X1  g175(.A1(new_n360), .A2(new_n361), .A3(new_n336), .ZN(new_n362));
  NAND3_X1  g176(.A1(new_n362), .A2(KEYINPUT75), .A3(KEYINPUT31), .ZN(new_n363));
  INV_X1    g177(.A(KEYINPUT76), .ZN(new_n364));
  NAND2_X1  g178(.A1(new_n353), .A2(new_n271), .ZN(new_n365));
  NAND3_X1  g179(.A1(new_n327), .A2(new_n365), .A3(new_n329), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n366), .A2(KEYINPUT28), .ZN(new_n367));
  INV_X1    g181(.A(KEYINPUT28), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n325), .A2(new_n368), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n367), .A2(new_n369), .ZN(new_n370));
  INV_X1    g184(.A(new_n336), .ZN(new_n371));
  AOI21_X1  g185(.A(new_n364), .B1(new_n370), .B2(new_n371), .ZN(new_n372));
  INV_X1    g186(.A(new_n369), .ZN(new_n373));
  AOI21_X1  g187(.A(new_n373), .B1(new_n366), .B2(KEYINPUT28), .ZN(new_n374));
  NOR3_X1   g188(.A1(new_n374), .A2(KEYINPUT76), .A3(new_n336), .ZN(new_n375));
  OAI211_X1 g189(.A(new_n359), .B(new_n363), .C1(new_n372), .C2(new_n375), .ZN(new_n376));
  NOR2_X1   g190(.A1(G472), .A2(G902), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n376), .A2(new_n377), .ZN(new_n378));
  INV_X1    g192(.A(KEYINPUT32), .ZN(new_n379));
  NAND2_X1  g193(.A1(new_n378), .A2(new_n379), .ZN(new_n380));
  INV_X1    g194(.A(new_n377), .ZN(new_n381));
  NOR2_X1   g195(.A1(new_n381), .A2(new_n379), .ZN(new_n382));
  NAND3_X1  g196(.A1(new_n327), .A2(new_n329), .A3(KEYINPUT77), .ZN(new_n383));
  AND2_X1   g197(.A1(new_n273), .A2(new_n324), .ZN(new_n384));
  OR2_X1    g198(.A1(new_n384), .A2(new_n328), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n383), .A2(new_n385), .ZN(new_n386));
  AOI21_X1  g200(.A(KEYINPUT77), .B1(new_n327), .B2(new_n329), .ZN(new_n387));
  OAI21_X1  g201(.A(KEYINPUT28), .B1(new_n386), .B2(new_n387), .ZN(new_n388));
  NAND4_X1  g202(.A1(new_n388), .A2(KEYINPUT29), .A3(new_n369), .A4(new_n336), .ZN(new_n389));
  NAND3_X1  g203(.A1(new_n367), .A2(new_n369), .A3(new_n336), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n360), .A2(new_n361), .ZN(new_n391));
  NAND2_X1  g205(.A1(new_n391), .A2(new_n371), .ZN(new_n392));
  INV_X1    g206(.A(KEYINPUT29), .ZN(new_n393));
  NAND3_X1  g207(.A1(new_n390), .A2(new_n392), .A3(new_n393), .ZN(new_n394));
  NAND3_X1  g208(.A1(new_n389), .A2(new_n394), .A3(new_n188), .ZN(new_n395));
  AOI22_X1  g209(.A1(new_n376), .A2(new_n382), .B1(new_n395), .B2(G472), .ZN(new_n396));
  AOI21_X1  g210(.A(new_n250), .B1(new_n380), .B2(new_n396), .ZN(new_n397));
  OAI21_X1  g211(.A(G214), .B1(G237), .B2(G902), .ZN(new_n398));
  INV_X1    g212(.A(KEYINPUT6), .ZN(new_n399));
  INV_X1    g213(.A(G104), .ZN(new_n400));
  NOR2_X1   g214(.A1(new_n400), .A2(KEYINPUT3), .ZN(new_n401));
  OR2_X1    g215(.A1(KEYINPUT87), .A2(G107), .ZN(new_n402));
  NAND2_X1  g216(.A1(KEYINPUT87), .A2(G107), .ZN(new_n403));
  AND3_X1   g217(.A1(new_n401), .A2(new_n402), .A3(new_n403), .ZN(new_n404));
  OAI21_X1  g218(.A(KEYINPUT3), .B1(new_n400), .B2(G107), .ZN(new_n405));
  INV_X1    g219(.A(KEYINPUT88), .ZN(new_n406));
  INV_X1    g220(.A(G107), .ZN(new_n407));
  OAI21_X1  g221(.A(new_n406), .B1(new_n407), .B2(G104), .ZN(new_n408));
  NAND3_X1  g222(.A1(new_n400), .A2(KEYINPUT88), .A3(G107), .ZN(new_n409));
  NAND3_X1  g223(.A1(new_n405), .A2(new_n408), .A3(new_n409), .ZN(new_n410));
  OAI21_X1  g224(.A(G101), .B1(new_n404), .B2(new_n410), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n400), .A2(G107), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n407), .A2(G104), .ZN(new_n413));
  AOI22_X1  g227(.A1(new_n406), .A2(new_n412), .B1(new_n413), .B2(KEYINPUT3), .ZN(new_n414));
  INV_X1    g228(.A(G101), .ZN(new_n415));
  NAND3_X1  g229(.A1(new_n401), .A2(new_n402), .A3(new_n403), .ZN(new_n416));
  NAND4_X1  g230(.A1(new_n414), .A2(new_n415), .A3(new_n416), .A4(new_n409), .ZN(new_n417));
  NAND3_X1  g231(.A1(new_n411), .A2(new_n417), .A3(KEYINPUT4), .ZN(new_n418));
  INV_X1    g232(.A(KEYINPUT4), .ZN(new_n419));
  OAI211_X1 g233(.A(new_n419), .B(G101), .C1(new_n404), .C2(new_n410), .ZN(new_n420));
  NAND3_X1  g234(.A1(new_n271), .A2(new_n418), .A3(new_n420), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n265), .A2(KEYINPUT5), .ZN(new_n422));
  INV_X1    g236(.A(G113), .ZN(new_n423));
  INV_X1    g237(.A(KEYINPUT5), .ZN(new_n424));
  AOI21_X1  g238(.A(new_n423), .B1(new_n252), .B2(new_n424), .ZN(new_n425));
  AOI22_X1  g239(.A1(new_n318), .A2(new_n319), .B1(new_n422), .B2(new_n425), .ZN(new_n426));
  AOI21_X1  g240(.A(G104), .B1(new_n402), .B2(new_n403), .ZN(new_n427));
  INV_X1    g241(.A(new_n413), .ZN(new_n428));
  OAI21_X1  g242(.A(G101), .B1(new_n427), .B2(new_n428), .ZN(new_n429));
  AND2_X1   g243(.A1(new_n417), .A2(new_n429), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n426), .A2(new_n430), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n421), .A2(new_n431), .ZN(new_n432));
  XNOR2_X1  g246(.A(G110), .B(G122), .ZN(new_n433));
  XNOR2_X1  g247(.A(new_n433), .B(KEYINPUT93), .ZN(new_n434));
  INV_X1    g248(.A(new_n434), .ZN(new_n435));
  AOI21_X1  g249(.A(new_n399), .B1(new_n432), .B2(new_n435), .ZN(new_n436));
  INV_X1    g250(.A(new_n410), .ZN(new_n437));
  AOI21_X1  g251(.A(new_n415), .B1(new_n437), .B2(new_n416), .ZN(new_n438));
  AOI22_X1  g252(.A1(new_n320), .A2(new_n323), .B1(new_n419), .B2(new_n438), .ZN(new_n439));
  AOI22_X1  g253(.A1(new_n439), .A2(new_n418), .B1(new_n430), .B2(new_n426), .ZN(new_n440));
  AOI21_X1  g254(.A(KEYINPUT94), .B1(new_n440), .B2(new_n434), .ZN(new_n441));
  NAND4_X1  g255(.A1(new_n421), .A2(KEYINPUT94), .A3(new_n434), .A4(new_n431), .ZN(new_n442));
  INV_X1    g256(.A(new_n442), .ZN(new_n443));
  OAI21_X1  g257(.A(new_n436), .B1(new_n441), .B2(new_n443), .ZN(new_n444));
  AOI211_X1 g258(.A(KEYINPUT6), .B(new_n434), .C1(new_n421), .C2(new_n431), .ZN(new_n445));
  INV_X1    g259(.A(new_n445), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n338), .A2(new_n339), .ZN(new_n447));
  NAND3_X1  g261(.A1(new_n447), .A2(new_n193), .A3(new_n281), .ZN(new_n448));
  OR2_X1    g262(.A1(new_n311), .A2(new_n193), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n448), .A2(new_n449), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n232), .A2(G224), .ZN(new_n451));
  XNOR2_X1  g265(.A(new_n450), .B(new_n451), .ZN(new_n452));
  INV_X1    g266(.A(new_n452), .ZN(new_n453));
  NAND3_X1  g267(.A1(new_n444), .A2(new_n446), .A3(new_n453), .ZN(new_n454));
  OAI21_X1  g268(.A(G210), .B1(G237), .B2(G902), .ZN(new_n455));
  XOR2_X1   g269(.A(new_n434), .B(KEYINPUT8), .Z(new_n456));
  OR2_X1    g270(.A1(new_n426), .A2(new_n430), .ZN(new_n457));
  AOI21_X1  g271(.A(new_n456), .B1(new_n457), .B2(new_n431), .ZN(new_n458));
  AND4_X1   g272(.A1(KEYINPUT7), .A2(new_n448), .A3(new_n451), .A4(new_n449), .ZN(new_n459));
  AOI22_X1  g273(.A1(new_n448), .A2(new_n449), .B1(KEYINPUT7), .B2(new_n451), .ZN(new_n460));
  NOR3_X1   g274(.A1(new_n458), .A2(new_n459), .A3(new_n460), .ZN(new_n461));
  NAND3_X1  g275(.A1(new_n421), .A2(new_n434), .A3(new_n431), .ZN(new_n462));
  INV_X1    g276(.A(KEYINPUT94), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n464), .A2(new_n442), .ZN(new_n465));
  AOI21_X1  g279(.A(G902), .B1(new_n461), .B2(new_n465), .ZN(new_n466));
  AND3_X1   g280(.A1(new_n454), .A2(new_n455), .A3(new_n466), .ZN(new_n467));
  AOI21_X1  g281(.A(new_n455), .B1(new_n454), .B2(new_n466), .ZN(new_n468));
  OAI21_X1  g282(.A(new_n398), .B1(new_n467), .B2(new_n468), .ZN(new_n469));
  INV_X1    g283(.A(KEYINPUT95), .ZN(new_n470));
  NAND2_X1  g284(.A1(new_n469), .A2(new_n470), .ZN(new_n471));
  INV_X1    g285(.A(new_n455), .ZN(new_n472));
  AOI211_X1 g286(.A(new_n445), .B(new_n452), .C1(new_n465), .C2(new_n436), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n461), .A2(new_n465), .ZN(new_n474));
  INV_X1    g288(.A(G902), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n474), .A2(new_n475), .ZN(new_n476));
  OAI21_X1  g290(.A(new_n472), .B1(new_n473), .B2(new_n476), .ZN(new_n477));
  NAND3_X1  g291(.A1(new_n454), .A2(new_n455), .A3(new_n466), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  NAND3_X1  g293(.A1(new_n479), .A2(KEYINPUT95), .A3(new_n398), .ZN(new_n480));
  NAND2_X1  g294(.A1(new_n471), .A2(new_n480), .ZN(new_n481));
  NOR2_X1   g295(.A1(G475), .A2(G902), .ZN(new_n482));
  INV_X1    g296(.A(G237), .ZN(new_n483));
  NAND3_X1  g297(.A1(new_n483), .A2(new_n232), .A3(G214), .ZN(new_n484));
  NOR2_X1   g298(.A1(KEYINPUT96), .A2(G143), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n484), .A2(new_n485), .ZN(new_n486));
  OAI211_X1 g300(.A(new_n332), .B(G214), .C1(KEYINPUT96), .C2(G143), .ZN(new_n487));
  NAND2_X1  g301(.A1(new_n486), .A2(new_n487), .ZN(new_n488));
  NAND2_X1  g302(.A1(new_n488), .A2(G131), .ZN(new_n489));
  INV_X1    g303(.A(KEYINPUT17), .ZN(new_n490));
  NAND3_X1  g304(.A1(new_n486), .A2(new_n487), .A3(new_n299), .ZN(new_n491));
  NAND3_X1  g305(.A1(new_n489), .A2(new_n490), .A3(new_n491), .ZN(new_n492));
  AOI21_X1  g306(.A(G146), .B1(new_n195), .B2(new_n196), .ZN(new_n493));
  AND3_X1   g307(.A1(new_n195), .A2(G146), .A3(new_n196), .ZN(new_n494));
  AOI21_X1  g308(.A(new_n493), .B1(new_n494), .B2(KEYINPUT80), .ZN(new_n495));
  NAND3_X1  g309(.A1(new_n488), .A2(KEYINPUT17), .A3(G131), .ZN(new_n496));
  NAND4_X1  g310(.A1(new_n492), .A2(new_n495), .A3(new_n199), .A4(new_n496), .ZN(new_n497));
  XNOR2_X1  g311(.A(G113), .B(G122), .ZN(new_n498));
  XNOR2_X1  g312(.A(new_n498), .B(new_n400), .ZN(new_n499));
  NAND3_X1  g313(.A1(new_n488), .A2(KEYINPUT18), .A3(G131), .ZN(new_n500));
  XNOR2_X1  g314(.A(new_n221), .B(G146), .ZN(new_n501));
  NAND2_X1  g315(.A1(KEYINPUT18), .A2(G131), .ZN(new_n502));
  NAND3_X1  g316(.A1(new_n486), .A2(new_n487), .A3(new_n502), .ZN(new_n503));
  NAND3_X1  g317(.A1(new_n500), .A2(new_n501), .A3(new_n503), .ZN(new_n504));
  AND3_X1   g318(.A1(new_n497), .A2(new_n499), .A3(new_n504), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n489), .A2(new_n491), .ZN(new_n506));
  AND3_X1   g320(.A1(new_n192), .A2(new_n194), .A3(KEYINPUT19), .ZN(new_n507));
  AOI21_X1  g321(.A(KEYINPUT19), .B1(new_n192), .B2(new_n194), .ZN(new_n508));
  NOR2_X1   g322(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  OAI211_X1 g323(.A(new_n220), .B(new_n506), .C1(G146), .C2(new_n509), .ZN(new_n510));
  AOI21_X1  g324(.A(new_n499), .B1(new_n510), .B2(new_n504), .ZN(new_n511));
  OAI21_X1  g325(.A(new_n482), .B1(new_n505), .B2(new_n511), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n510), .A2(new_n504), .ZN(new_n513));
  INV_X1    g327(.A(new_n499), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  NAND3_X1  g329(.A1(new_n497), .A2(new_n499), .A3(new_n504), .ZN(new_n516));
  AOI21_X1  g330(.A(KEYINPUT97), .B1(new_n515), .B2(new_n516), .ZN(new_n517));
  OAI21_X1  g331(.A(new_n512), .B1(new_n517), .B2(KEYINPUT20), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n515), .A2(new_n516), .ZN(new_n519));
  INV_X1    g333(.A(KEYINPUT20), .ZN(new_n520));
  NAND4_X1  g334(.A1(new_n519), .A2(KEYINPUT97), .A3(new_n520), .A4(new_n482), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n518), .A2(new_n521), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n492), .A2(new_n496), .ZN(new_n523));
  OAI21_X1  g337(.A(new_n504), .B1(new_n523), .B2(new_n202), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n524), .A2(new_n514), .ZN(new_n525));
  AOI21_X1  g339(.A(G902), .B1(new_n525), .B2(new_n516), .ZN(new_n526));
  INV_X1    g340(.A(KEYINPUT99), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  AOI21_X1  g342(.A(new_n499), .B1(new_n497), .B2(new_n504), .ZN(new_n529));
  OAI21_X1  g343(.A(new_n475), .B1(new_n505), .B2(new_n529), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n530), .A2(KEYINPUT99), .ZN(new_n531));
  XNOR2_X1  g345(.A(KEYINPUT98), .B(G475), .ZN(new_n532));
  NAND3_X1  g346(.A1(new_n528), .A2(new_n531), .A3(new_n532), .ZN(new_n533));
  AND2_X1   g347(.A1(new_n522), .A2(new_n533), .ZN(new_n534));
  NAND2_X1  g348(.A1(new_n232), .A2(G952), .ZN(new_n535));
  AOI21_X1  g349(.A(new_n535), .B1(G234), .B2(G237), .ZN(new_n536));
  AOI211_X1 g350(.A(new_n232), .B(new_n188), .C1(G234), .C2(G237), .ZN(new_n537));
  XNOR2_X1  g351(.A(KEYINPUT21), .B(G898), .ZN(new_n538));
  AOI21_X1  g352(.A(new_n536), .B1(new_n537), .B2(new_n538), .ZN(new_n539));
  INV_X1    g353(.A(new_n539), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n534), .A2(new_n540), .ZN(new_n541));
  XNOR2_X1  g355(.A(G128), .B(G143), .ZN(new_n542));
  XNOR2_X1  g356(.A(new_n542), .B(new_n295), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n402), .A2(new_n403), .ZN(new_n544));
  INV_X1    g358(.A(G122), .ZN(new_n545));
  NAND2_X1  g359(.A1(new_n545), .A2(G116), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n251), .A2(G122), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n546), .A2(new_n547), .ZN(new_n548));
  OR2_X1    g362(.A1(new_n544), .A2(new_n548), .ZN(new_n549));
  OAI21_X1  g363(.A(new_n546), .B1(new_n547), .B2(KEYINPUT14), .ZN(new_n550));
  INV_X1    g364(.A(KEYINPUT100), .ZN(new_n551));
  NAND3_X1  g365(.A1(new_n547), .A2(new_n551), .A3(KEYINPUT14), .ZN(new_n552));
  OAI21_X1  g366(.A(KEYINPUT14), .B1(new_n545), .B2(G116), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n553), .A2(KEYINPUT100), .ZN(new_n554));
  AOI21_X1  g368(.A(new_n550), .B1(new_n552), .B2(new_n554), .ZN(new_n555));
  OAI211_X1 g369(.A(new_n543), .B(new_n549), .C1(new_n407), .C2(new_n555), .ZN(new_n556));
  XNOR2_X1  g370(.A(new_n544), .B(new_n548), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n542), .A2(KEYINPUT13), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n274), .A2(G128), .ZN(new_n559));
  OAI211_X1 g373(.A(new_n558), .B(G134), .C1(KEYINPUT13), .C2(new_n559), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n542), .A2(new_n295), .ZN(new_n561));
  NAND3_X1  g375(.A1(new_n557), .A2(new_n560), .A3(new_n561), .ZN(new_n562));
  XNOR2_X1  g376(.A(KEYINPUT9), .B(G234), .ZN(new_n563));
  NOR3_X1   g377(.A1(new_n563), .A2(new_n187), .A3(G953), .ZN(new_n564));
  AND3_X1   g378(.A1(new_n556), .A2(new_n562), .A3(new_n564), .ZN(new_n565));
  AOI21_X1  g379(.A(new_n564), .B1(new_n556), .B2(new_n562), .ZN(new_n566));
  OAI21_X1  g380(.A(new_n188), .B1(new_n565), .B2(new_n566), .ZN(new_n567));
  INV_X1    g381(.A(KEYINPUT15), .ZN(new_n568));
  NAND3_X1  g382(.A1(new_n567), .A2(new_n568), .A3(G478), .ZN(new_n569));
  INV_X1    g383(.A(G478), .ZN(new_n570));
  OAI221_X1 g384(.A(new_n188), .B1(KEYINPUT15), .B2(new_n570), .C1(new_n565), .C2(new_n566), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n569), .A2(new_n571), .ZN(new_n572));
  NOR2_X1   g386(.A1(new_n541), .A2(new_n572), .ZN(new_n573));
  INV_X1    g387(.A(G469), .ZN(new_n574));
  XNOR2_X1  g388(.A(G110), .B(G140), .ZN(new_n575));
  XNOR2_X1  g389(.A(new_n575), .B(KEYINPUT86), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n232), .A2(G227), .ZN(new_n577));
  XNOR2_X1  g391(.A(new_n576), .B(new_n577), .ZN(new_n578));
  INV_X1    g392(.A(KEYINPUT89), .ZN(new_n579));
  AND3_X1   g393(.A1(new_n411), .A2(new_n417), .A3(KEYINPUT4), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n420), .A2(new_n311), .ZN(new_n581));
  OAI21_X1  g395(.A(new_n579), .B1(new_n580), .B2(new_n581), .ZN(new_n582));
  NAND4_X1  g396(.A1(new_n418), .A2(KEYINPUT89), .A3(new_n311), .A4(new_n420), .ZN(new_n583));
  NAND2_X1  g397(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n417), .A2(new_n429), .ZN(new_n585));
  OAI21_X1  g399(.A(KEYINPUT10), .B1(new_n340), .B2(new_n585), .ZN(new_n586));
  INV_X1    g400(.A(new_n291), .ZN(new_n587));
  INV_X1    g401(.A(KEYINPUT90), .ZN(new_n588));
  NAND2_X1  g402(.A1(new_n275), .A2(new_n588), .ZN(new_n589));
  NAND3_X1  g403(.A1(new_n278), .A2(KEYINPUT90), .A3(KEYINPUT1), .ZN(new_n590));
  NAND3_X1  g404(.A1(new_n589), .A2(G128), .A3(new_n590), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n587), .A2(new_n591), .ZN(new_n592));
  OAI21_X1  g406(.A(new_n592), .B1(new_n287), .B2(new_n292), .ZN(new_n593));
  INV_X1    g407(.A(KEYINPUT10), .ZN(new_n594));
  NAND3_X1  g408(.A1(new_n593), .A2(new_n594), .A3(new_n430), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n586), .A2(new_n595), .ZN(new_n596));
  INV_X1    g410(.A(new_n314), .ZN(new_n597));
  NAND3_X1  g411(.A1(new_n584), .A2(new_n596), .A3(new_n597), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n598), .A2(KEYINPUT91), .ZN(new_n599));
  INV_X1    g413(.A(KEYINPUT91), .ZN(new_n600));
  NAND4_X1  g414(.A1(new_n584), .A2(new_n596), .A3(new_n600), .A4(new_n597), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n599), .A2(new_n601), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n584), .A2(new_n596), .ZN(new_n603));
  NAND2_X1  g417(.A1(new_n603), .A2(KEYINPUT92), .ZN(new_n604));
  INV_X1    g418(.A(KEYINPUT92), .ZN(new_n605));
  NAND3_X1  g419(.A1(new_n584), .A2(new_n596), .A3(new_n605), .ZN(new_n606));
  NAND3_X1  g420(.A1(new_n604), .A2(new_n606), .A3(new_n314), .ZN(new_n607));
  AOI21_X1  g421(.A(new_n578), .B1(new_n602), .B2(new_n607), .ZN(new_n608));
  INV_X1    g422(.A(new_n578), .ZN(new_n609));
  NOR2_X1   g423(.A1(new_n293), .A2(new_n430), .ZN(new_n610));
  AOI21_X1  g424(.A(new_n585), .B1(new_n447), .B2(new_n592), .ZN(new_n611));
  OAI211_X1 g425(.A(KEYINPUT12), .B(new_n314), .C1(new_n610), .C2(new_n611), .ZN(new_n612));
  OAI21_X1  g426(.A(new_n314), .B1(new_n610), .B2(new_n611), .ZN(new_n613));
  INV_X1    g427(.A(KEYINPUT12), .ZN(new_n614));
  NAND2_X1  g428(.A1(new_n613), .A2(new_n614), .ZN(new_n615));
  AOI221_X4 g429(.A(new_n609), .B1(new_n612), .B2(new_n615), .C1(new_n599), .C2(new_n601), .ZN(new_n616));
  OAI211_X1 g430(.A(new_n574), .B(new_n188), .C1(new_n608), .C2(new_n616), .ZN(new_n617));
  NAND2_X1  g431(.A1(G469), .A2(G902), .ZN(new_n618));
  NAND2_X1  g432(.A1(new_n615), .A2(new_n612), .ZN(new_n619));
  NAND2_X1  g433(.A1(new_n602), .A2(new_n619), .ZN(new_n620));
  NAND2_X1  g434(.A1(new_n620), .A2(new_n609), .ZN(new_n621));
  AOI21_X1  g435(.A(new_n609), .B1(new_n599), .B2(new_n601), .ZN(new_n622));
  NAND2_X1  g436(.A1(new_n622), .A2(new_n607), .ZN(new_n623));
  NAND3_X1  g437(.A1(new_n621), .A2(G469), .A3(new_n623), .ZN(new_n624));
  NAND3_X1  g438(.A1(new_n617), .A2(new_n618), .A3(new_n624), .ZN(new_n625));
  OAI21_X1  g439(.A(G221), .B1(new_n563), .B2(G902), .ZN(new_n626));
  XNOR2_X1  g440(.A(new_n626), .B(KEYINPUT85), .ZN(new_n627));
  INV_X1    g441(.A(new_n627), .ZN(new_n628));
  NAND3_X1  g442(.A1(new_n573), .A2(new_n625), .A3(new_n628), .ZN(new_n629));
  NOR2_X1   g443(.A1(new_n481), .A2(new_n629), .ZN(new_n630));
  NAND2_X1  g444(.A1(new_n397), .A2(new_n630), .ZN(new_n631));
  XNOR2_X1  g445(.A(new_n631), .B(G101), .ZN(G3));
  INV_X1    g446(.A(KEYINPUT101), .ZN(new_n633));
  AND2_X1   g447(.A1(new_n359), .A2(new_n363), .ZN(new_n634));
  NAND3_X1  g448(.A1(new_n370), .A2(new_n364), .A3(new_n371), .ZN(new_n635));
  OAI21_X1  g449(.A(KEYINPUT76), .B1(new_n374), .B2(new_n336), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n635), .A2(new_n636), .ZN(new_n637));
  AOI21_X1  g451(.A(new_n190), .B1(new_n634), .B2(new_n637), .ZN(new_n638));
  INV_X1    g452(.A(G472), .ZN(new_n639));
  OAI21_X1  g453(.A(new_n378), .B1(new_n638), .B2(new_n639), .ZN(new_n640));
  INV_X1    g454(.A(new_n250), .ZN(new_n641));
  NAND3_X1  g455(.A1(new_n625), .A2(new_n641), .A3(new_n628), .ZN(new_n642));
  OAI21_X1  g456(.A(new_n633), .B1(new_n640), .B2(new_n642), .ZN(new_n643));
  INV_X1    g457(.A(new_n642), .ZN(new_n644));
  NAND2_X1  g458(.A1(new_n376), .A2(new_n188), .ZN(new_n645));
  NAND2_X1  g459(.A1(new_n645), .A2(G472), .ZN(new_n646));
  NAND4_X1  g460(.A1(new_n644), .A2(KEYINPUT101), .A3(new_n646), .A4(new_n378), .ZN(new_n647));
  NAND2_X1  g461(.A1(new_n643), .A2(new_n647), .ZN(new_n648));
  INV_X1    g462(.A(new_n648), .ZN(new_n649));
  INV_X1    g463(.A(new_n398), .ZN(new_n650));
  AOI21_X1  g464(.A(new_n650), .B1(new_n477), .B2(new_n478), .ZN(new_n651));
  INV_X1    g465(.A(KEYINPUT33), .ZN(new_n652));
  OR3_X1    g466(.A1(new_n565), .A2(new_n566), .A3(new_n652), .ZN(new_n653));
  OAI21_X1  g467(.A(new_n652), .B1(new_n565), .B2(new_n566), .ZN(new_n654));
  NAND4_X1  g468(.A1(new_n653), .A2(G478), .A3(new_n188), .A4(new_n654), .ZN(new_n655));
  NAND2_X1  g469(.A1(new_n567), .A2(new_n570), .ZN(new_n656));
  NAND2_X1  g470(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  INV_X1    g471(.A(new_n657), .ZN(new_n658));
  NOR2_X1   g472(.A1(new_n534), .A2(new_n658), .ZN(new_n659));
  NAND4_X1  g473(.A1(new_n649), .A2(new_n651), .A3(new_n540), .A4(new_n659), .ZN(new_n660));
  XNOR2_X1  g474(.A(new_n660), .B(KEYINPUT34), .ZN(new_n661));
  XNOR2_X1  g475(.A(new_n661), .B(new_n400), .ZN(G6));
  INV_X1    g476(.A(KEYINPUT102), .ZN(new_n663));
  NAND3_X1  g477(.A1(new_n512), .A2(new_n663), .A3(new_n520), .ZN(new_n664));
  NAND2_X1  g478(.A1(KEYINPUT102), .A2(KEYINPUT20), .ZN(new_n665));
  NAND2_X1  g479(.A1(new_n663), .A2(new_n520), .ZN(new_n666));
  NAND4_X1  g480(.A1(new_n519), .A2(new_n482), .A3(new_n665), .A4(new_n666), .ZN(new_n667));
  AND3_X1   g481(.A1(new_n664), .A2(new_n572), .A3(new_n667), .ZN(new_n668));
  INV_X1    g482(.A(KEYINPUT103), .ZN(new_n669));
  OAI21_X1  g483(.A(new_n532), .B1(new_n526), .B2(new_n527), .ZN(new_n670));
  NOR2_X1   g484(.A1(new_n530), .A2(KEYINPUT99), .ZN(new_n671));
  OAI21_X1  g485(.A(new_n669), .B1(new_n670), .B2(new_n671), .ZN(new_n672));
  NAND4_X1  g486(.A1(new_n528), .A2(new_n531), .A3(KEYINPUT103), .A4(new_n532), .ZN(new_n673));
  AND3_X1   g487(.A1(new_n668), .A2(new_n672), .A3(new_n673), .ZN(new_n674));
  NAND4_X1  g488(.A1(new_n479), .A2(new_n398), .A3(new_n674), .A4(new_n540), .ZN(new_n675));
  NOR2_X1   g489(.A1(new_n648), .A2(new_n675), .ZN(new_n676));
  XNOR2_X1  g490(.A(KEYINPUT35), .B(G107), .ZN(new_n677));
  XNOR2_X1  g491(.A(new_n676), .B(new_n677), .ZN(G9));
  INV_X1    g492(.A(KEYINPUT105), .ZN(new_n679));
  NOR2_X1   g493(.A1(new_n234), .A2(KEYINPUT36), .ZN(new_n680));
  XNOR2_X1  g494(.A(new_n229), .B(new_n680), .ZN(new_n681));
  NAND2_X1  g495(.A1(new_n681), .A2(new_n248), .ZN(new_n682));
  NAND3_X1  g496(.A1(new_n246), .A2(KEYINPUT104), .A3(new_n682), .ZN(new_n683));
  INV_X1    g497(.A(KEYINPUT104), .ZN(new_n684));
  INV_X1    g498(.A(new_n189), .ZN(new_n685));
  OAI21_X1  g499(.A(KEYINPUT25), .B1(new_n238), .B2(new_n239), .ZN(new_n686));
  NAND3_X1  g500(.A1(new_n244), .A2(KEYINPUT84), .A3(new_n241), .ZN(new_n687));
  AOI21_X1  g501(.A(new_n685), .B1(new_n686), .B2(new_n687), .ZN(new_n688));
  INV_X1    g502(.A(new_n682), .ZN(new_n689));
  OAI21_X1  g503(.A(new_n684), .B1(new_n688), .B2(new_n689), .ZN(new_n690));
  NAND2_X1  g504(.A1(new_n683), .A2(new_n690), .ZN(new_n691));
  INV_X1    g505(.A(new_n691), .ZN(new_n692));
  OAI21_X1  g506(.A(new_n679), .B1(new_n640), .B2(new_n692), .ZN(new_n693));
  NAND4_X1  g507(.A1(new_n646), .A2(KEYINPUT105), .A3(new_n378), .A4(new_n691), .ZN(new_n694));
  NAND3_X1  g508(.A1(new_n693), .A2(new_n630), .A3(new_n694), .ZN(new_n695));
  XNOR2_X1  g509(.A(new_n695), .B(KEYINPUT106), .ZN(new_n696));
  XNOR2_X1  g510(.A(KEYINPUT37), .B(G110), .ZN(new_n697));
  XNOR2_X1  g511(.A(new_n696), .B(new_n697), .ZN(G12));
  NAND2_X1  g512(.A1(new_n376), .A2(new_n382), .ZN(new_n699));
  NAND2_X1  g513(.A1(new_n395), .A2(G472), .ZN(new_n700));
  AOI21_X1  g514(.A(new_n381), .B1(new_n634), .B2(new_n637), .ZN(new_n701));
  OAI211_X1 g515(.A(new_n699), .B(new_n700), .C1(new_n701), .C2(KEYINPUT32), .ZN(new_n702));
  INV_X1    g516(.A(KEYINPUT107), .ZN(new_n703));
  INV_X1    g517(.A(G900), .ZN(new_n704));
  AOI21_X1  g518(.A(new_n536), .B1(new_n537), .B2(new_n704), .ZN(new_n705));
  INV_X1    g519(.A(new_n705), .ZN(new_n706));
  NAND2_X1  g520(.A1(new_n674), .A2(new_n706), .ZN(new_n707));
  OAI21_X1  g521(.A(new_n703), .B1(new_n707), .B2(new_n469), .ZN(new_n708));
  NAND4_X1  g522(.A1(new_n651), .A2(KEYINPUT107), .A3(new_n674), .A4(new_n706), .ZN(new_n709));
  NAND2_X1  g523(.A1(new_n708), .A2(new_n709), .ZN(new_n710));
  NAND3_X1  g524(.A1(new_n691), .A2(new_n625), .A3(new_n628), .ZN(new_n711));
  INV_X1    g525(.A(new_n711), .ZN(new_n712));
  NAND3_X1  g526(.A1(new_n702), .A2(new_n710), .A3(new_n712), .ZN(new_n713));
  XNOR2_X1  g527(.A(new_n713), .B(G128), .ZN(G30));
  NAND2_X1  g528(.A1(new_n391), .A2(new_n336), .ZN(new_n715));
  OR2_X1    g529(.A1(new_n386), .A2(new_n387), .ZN(new_n716));
  OAI211_X1 g530(.A(new_n475), .B(new_n715), .C1(new_n716), .C2(new_n336), .ZN(new_n717));
  NAND2_X1  g531(.A1(new_n717), .A2(G472), .ZN(new_n718));
  OAI211_X1 g532(.A(new_n699), .B(new_n718), .C1(new_n701), .C2(KEYINPUT32), .ZN(new_n719));
  INV_X1    g533(.A(KEYINPUT108), .ZN(new_n720));
  XNOR2_X1  g534(.A(new_n719), .B(new_n720), .ZN(new_n721));
  XOR2_X1   g535(.A(new_n705), .B(KEYINPUT39), .Z(new_n722));
  NAND3_X1  g536(.A1(new_n625), .A2(new_n628), .A3(new_n722), .ZN(new_n723));
  XOR2_X1   g537(.A(new_n723), .B(KEYINPUT40), .Z(new_n724));
  XNOR2_X1  g538(.A(new_n479), .B(KEYINPUT38), .ZN(new_n725));
  INV_X1    g539(.A(new_n572), .ZN(new_n726));
  AOI21_X1  g540(.A(new_n726), .B1(new_n522), .B2(new_n533), .ZN(new_n727));
  NAND2_X1  g541(.A1(new_n727), .A2(new_n398), .ZN(new_n728));
  NOR2_X1   g542(.A1(new_n691), .A2(new_n728), .ZN(new_n729));
  NAND4_X1  g543(.A1(new_n721), .A2(new_n724), .A3(new_n725), .A4(new_n729), .ZN(new_n730));
  OR2_X1    g544(.A1(new_n730), .A2(KEYINPUT109), .ZN(new_n731));
  NAND2_X1  g545(.A1(new_n730), .A2(KEYINPUT109), .ZN(new_n732));
  NAND2_X1  g546(.A1(new_n731), .A2(new_n732), .ZN(new_n733));
  XNOR2_X1  g547(.A(new_n733), .B(new_n274), .ZN(G45));
  NOR3_X1   g548(.A1(new_n534), .A2(new_n658), .A3(new_n705), .ZN(new_n735));
  NAND2_X1  g549(.A1(new_n735), .A2(new_n651), .ZN(new_n736));
  INV_X1    g550(.A(new_n736), .ZN(new_n737));
  NAND3_X1  g551(.A1(new_n702), .A2(new_n712), .A3(new_n737), .ZN(new_n738));
  XOR2_X1   g552(.A(KEYINPUT110), .B(G146), .Z(new_n739));
  XNOR2_X1  g553(.A(new_n738), .B(new_n739), .ZN(G48));
  NAND2_X1  g554(.A1(new_n602), .A2(new_n607), .ZN(new_n741));
  AOI22_X1  g555(.A1(new_n741), .A2(new_n609), .B1(new_n619), .B2(new_n622), .ZN(new_n742));
  OAI21_X1  g556(.A(G469), .B1(new_n742), .B2(new_n190), .ZN(new_n743));
  AND4_X1   g557(.A1(new_n651), .A2(new_n743), .A3(new_n626), .A4(new_n617), .ZN(new_n744));
  AND3_X1   g558(.A1(new_n744), .A2(new_n540), .A3(new_n659), .ZN(new_n745));
  NAND2_X1  g559(.A1(new_n745), .A2(new_n397), .ZN(new_n746));
  XNOR2_X1  g560(.A(new_n746), .B(KEYINPUT41), .ZN(new_n747));
  XNOR2_X1  g561(.A(new_n747), .B(G113), .ZN(G15));
  NAND3_X1  g562(.A1(new_n743), .A2(new_n626), .A3(new_n617), .ZN(new_n749));
  NOR2_X1   g563(.A1(new_n749), .A2(new_n675), .ZN(new_n750));
  NAND2_X1  g564(.A1(new_n699), .A2(new_n700), .ZN(new_n751));
  AOI21_X1  g565(.A(KEYINPUT32), .B1(new_n376), .B2(new_n377), .ZN(new_n752));
  OAI211_X1 g566(.A(new_n750), .B(new_n641), .C1(new_n751), .C2(new_n752), .ZN(new_n753));
  XNOR2_X1  g567(.A(new_n753), .B(G116), .ZN(G18));
  AND2_X1   g568(.A1(new_n691), .A2(new_n573), .ZN(new_n755));
  OAI211_X1 g569(.A(new_n744), .B(new_n755), .C1(new_n751), .C2(new_n752), .ZN(new_n756));
  XNOR2_X1  g570(.A(new_n756), .B(G119), .ZN(G21));
  NAND4_X1  g571(.A1(new_n479), .A2(new_n398), .A3(new_n727), .A4(new_n540), .ZN(new_n758));
  NOR2_X1   g572(.A1(new_n749), .A2(new_n758), .ZN(new_n759));
  XOR2_X1   g573(.A(new_n362), .B(KEYINPUT31), .Z(new_n760));
  NAND2_X1  g574(.A1(new_n388), .A2(new_n369), .ZN(new_n761));
  NAND2_X1  g575(.A1(new_n761), .A2(new_n371), .ZN(new_n762));
  AOI21_X1  g576(.A(new_n381), .B1(new_n760), .B2(new_n762), .ZN(new_n763));
  INV_X1    g577(.A(new_n763), .ZN(new_n764));
  NAND4_X1  g578(.A1(new_n759), .A2(new_n646), .A3(new_n641), .A4(new_n764), .ZN(new_n765));
  XNOR2_X1  g579(.A(new_n765), .B(G122), .ZN(G24));
  NOR2_X1   g580(.A1(new_n749), .A2(new_n736), .ZN(new_n767));
  NAND4_X1  g581(.A1(new_n767), .A2(new_n646), .A3(new_n691), .A4(new_n764), .ZN(new_n768));
  XNOR2_X1  g582(.A(new_n768), .B(G125), .ZN(G27));
  NOR3_X1   g583(.A1(new_n467), .A2(new_n468), .A3(new_n650), .ZN(new_n770));
  AND4_X1   g584(.A1(new_n626), .A2(new_n625), .A3(new_n735), .A4(new_n770), .ZN(new_n771));
  AOI21_X1  g585(.A(KEYINPUT42), .B1(new_n397), .B2(new_n771), .ZN(new_n772));
  AND4_X1   g586(.A1(KEYINPUT42), .A2(new_n702), .A3(new_n771), .A4(new_n641), .ZN(new_n773));
  OR2_X1    g587(.A1(new_n772), .A2(new_n773), .ZN(new_n774));
  XNOR2_X1  g588(.A(new_n774), .B(G131), .ZN(G33));
  NAND3_X1  g589(.A1(new_n625), .A2(new_n626), .A3(new_n770), .ZN(new_n776));
  NOR2_X1   g590(.A1(new_n776), .A2(new_n707), .ZN(new_n777));
  NAND2_X1  g591(.A1(new_n397), .A2(new_n777), .ZN(new_n778));
  XNOR2_X1  g592(.A(new_n778), .B(G134), .ZN(G36));
  INV_X1    g593(.A(new_n626), .ZN(new_n780));
  NAND2_X1  g594(.A1(new_n621), .A2(new_n623), .ZN(new_n781));
  INV_X1    g595(.A(KEYINPUT45), .ZN(new_n782));
  AOI21_X1  g596(.A(new_n574), .B1(new_n781), .B2(new_n782), .ZN(new_n783));
  OAI21_X1  g597(.A(new_n783), .B1(new_n782), .B2(new_n781), .ZN(new_n784));
  AOI21_X1  g598(.A(KEYINPUT46), .B1(new_n784), .B2(new_n618), .ZN(new_n785));
  INV_X1    g599(.A(new_n617), .ZN(new_n786));
  NOR2_X1   g600(.A1(new_n785), .A2(new_n786), .ZN(new_n787));
  NAND3_X1  g601(.A1(new_n784), .A2(KEYINPUT46), .A3(new_n618), .ZN(new_n788));
  AOI21_X1  g602(.A(new_n780), .B1(new_n787), .B2(new_n788), .ZN(new_n789));
  AND2_X1   g603(.A1(new_n789), .A2(new_n722), .ZN(new_n790));
  NAND2_X1  g604(.A1(new_n534), .A2(new_n657), .ZN(new_n791));
  XNOR2_X1  g605(.A(new_n791), .B(KEYINPUT43), .ZN(new_n792));
  NOR2_X1   g606(.A1(new_n792), .A2(new_n692), .ZN(new_n793));
  NAND3_X1  g607(.A1(new_n793), .A2(KEYINPUT44), .A3(new_n640), .ZN(new_n794));
  XNOR2_X1  g608(.A(new_n794), .B(KEYINPUT111), .ZN(new_n795));
  AOI21_X1  g609(.A(KEYINPUT44), .B1(new_n793), .B2(new_n640), .ZN(new_n796));
  INV_X1    g610(.A(new_n770), .ZN(new_n797));
  NOR2_X1   g611(.A1(new_n796), .A2(new_n797), .ZN(new_n798));
  NAND3_X1  g612(.A1(new_n790), .A2(new_n795), .A3(new_n798), .ZN(new_n799));
  XNOR2_X1  g613(.A(new_n799), .B(G137), .ZN(G39));
  INV_X1    g614(.A(KEYINPUT47), .ZN(new_n801));
  OR2_X1    g615(.A1(new_n789), .A2(new_n801), .ZN(new_n802));
  NAND2_X1  g616(.A1(new_n789), .A2(new_n801), .ZN(new_n803));
  NAND3_X1  g617(.A1(new_n770), .A2(new_n250), .A3(new_n735), .ZN(new_n804));
  NOR2_X1   g618(.A1(new_n702), .A2(new_n804), .ZN(new_n805));
  NAND3_X1  g619(.A1(new_n802), .A2(new_n803), .A3(new_n805), .ZN(new_n806));
  XNOR2_X1  g620(.A(new_n806), .B(G140), .ZN(G42));
  INV_X1    g621(.A(new_n721), .ZN(new_n808));
  NOR2_X1   g622(.A1(new_n749), .A2(new_n797), .ZN(new_n809));
  NAND4_X1  g623(.A1(new_n808), .A2(new_n641), .A3(new_n536), .A4(new_n809), .ZN(new_n810));
  OR2_X1    g624(.A1(new_n810), .A2(KEYINPUT115), .ZN(new_n811));
  NAND2_X1  g625(.A1(new_n810), .A2(KEYINPUT115), .ZN(new_n812));
  NAND4_X1  g626(.A1(new_n811), .A2(new_n534), .A3(new_n658), .A4(new_n812), .ZN(new_n813));
  INV_X1    g627(.A(new_n536), .ZN(new_n814));
  NOR2_X1   g628(.A1(new_n792), .A2(new_n814), .ZN(new_n815));
  AND4_X1   g629(.A1(new_n641), .A2(new_n815), .A3(new_n646), .A4(new_n764), .ZN(new_n816));
  AND2_X1   g630(.A1(new_n802), .A2(new_n803), .ZN(new_n817));
  AND2_X1   g631(.A1(new_n743), .A2(new_n617), .ZN(new_n818));
  AND2_X1   g632(.A1(new_n818), .A2(new_n627), .ZN(new_n819));
  OAI211_X1 g633(.A(new_n770), .B(new_n816), .C1(new_n817), .C2(new_n819), .ZN(new_n820));
  AOI21_X1  g634(.A(new_n639), .B1(new_n376), .B2(new_n188), .ZN(new_n821));
  NOR3_X1   g635(.A1(new_n821), .A2(new_n692), .A3(new_n763), .ZN(new_n822));
  AND3_X1   g636(.A1(new_n822), .A2(new_n815), .A3(new_n809), .ZN(new_n823));
  NOR3_X1   g637(.A1(new_n725), .A2(new_n398), .A3(new_n749), .ZN(new_n824));
  NAND2_X1  g638(.A1(new_n816), .A2(new_n824), .ZN(new_n825));
  INV_X1    g639(.A(KEYINPUT50), .ZN(new_n826));
  NAND2_X1  g640(.A1(new_n825), .A2(new_n826), .ZN(new_n827));
  NAND3_X1  g641(.A1(new_n816), .A2(KEYINPUT50), .A3(new_n824), .ZN(new_n828));
  AOI21_X1  g642(.A(new_n823), .B1(new_n827), .B2(new_n828), .ZN(new_n829));
  NAND3_X1  g643(.A1(new_n813), .A2(new_n820), .A3(new_n829), .ZN(new_n830));
  INV_X1    g644(.A(KEYINPUT51), .ZN(new_n831));
  NAND2_X1  g645(.A1(new_n830), .A2(new_n831), .ZN(new_n832));
  NAND4_X1  g646(.A1(new_n813), .A2(new_n820), .A3(KEYINPUT51), .A4(new_n829), .ZN(new_n833));
  NAND3_X1  g647(.A1(new_n811), .A2(new_n659), .A3(new_n812), .ZN(new_n834));
  NAND3_X1  g648(.A1(new_n397), .A2(new_n815), .A3(new_n809), .ZN(new_n835));
  XOR2_X1   g649(.A(new_n835), .B(KEYINPUT48), .Z(new_n836));
  AOI211_X1 g650(.A(new_n535), .B(new_n836), .C1(new_n744), .C2(new_n816), .ZN(new_n837));
  NAND4_X1  g651(.A1(new_n832), .A2(new_n833), .A3(new_n834), .A4(new_n837), .ZN(new_n838));
  AND3_X1   g652(.A1(new_n753), .A2(new_n756), .A3(new_n765), .ZN(new_n839));
  NOR2_X1   g653(.A1(new_n541), .A2(new_n726), .ZN(new_n840));
  NAND3_X1  g654(.A1(new_n471), .A2(new_n480), .A3(new_n840), .ZN(new_n841));
  INV_X1    g655(.A(KEYINPUT112), .ZN(new_n842));
  NAND2_X1  g656(.A1(new_n841), .A2(new_n842), .ZN(new_n843));
  NAND4_X1  g657(.A1(new_n471), .A2(KEYINPUT112), .A3(new_n480), .A4(new_n840), .ZN(new_n844));
  NAND4_X1  g658(.A1(new_n471), .A2(new_n480), .A3(new_n540), .A4(new_n659), .ZN(new_n845));
  NAND3_X1  g659(.A1(new_n843), .A2(new_n844), .A3(new_n845), .ZN(new_n846));
  NAND3_X1  g660(.A1(new_n846), .A2(new_n643), .A3(new_n647), .ZN(new_n847));
  OAI21_X1  g661(.A(new_n397), .B1(new_n745), .B2(new_n630), .ZN(new_n848));
  AND4_X1   g662(.A1(new_n695), .A2(new_n839), .A3(new_n847), .A4(new_n848), .ZN(new_n849));
  AOI21_X1  g663(.A(new_n711), .B1(new_n380), .B2(new_n396), .ZN(new_n850));
  AOI22_X1  g664(.A1(new_n850), .A2(new_n710), .B1(new_n822), .B2(new_n767), .ZN(new_n851));
  AOI21_X1  g665(.A(new_n728), .B1(new_n477), .B2(new_n478), .ZN(new_n852));
  NOR4_X1   g666(.A1(new_n688), .A2(new_n780), .A3(new_n689), .A4(new_n705), .ZN(new_n853));
  AND3_X1   g667(.A1(new_n852), .A2(new_n625), .A3(new_n853), .ZN(new_n854));
  NAND2_X1  g668(.A1(new_n719), .A2(new_n854), .ZN(new_n855));
  NAND4_X1  g669(.A1(new_n851), .A2(KEYINPUT52), .A3(new_n738), .A4(new_n855), .ZN(new_n856));
  NAND4_X1  g670(.A1(new_n713), .A2(new_n738), .A3(new_n768), .A4(new_n855), .ZN(new_n857));
  INV_X1    g671(.A(KEYINPUT52), .ZN(new_n858));
  NAND2_X1  g672(.A1(new_n857), .A2(new_n858), .ZN(new_n859));
  NAND2_X1  g673(.A1(new_n856), .A2(new_n859), .ZN(new_n860));
  AND4_X1   g674(.A1(new_n726), .A2(new_n664), .A3(new_n667), .A4(new_n706), .ZN(new_n861));
  AND4_X1   g675(.A1(new_n672), .A2(new_n770), .A3(new_n673), .A4(new_n861), .ZN(new_n862));
  AOI22_X1  g676(.A1(new_n850), .A2(new_n862), .B1(new_n822), .B2(new_n771), .ZN(new_n863));
  OAI211_X1 g677(.A(new_n863), .B(new_n778), .C1(new_n772), .C2(new_n773), .ZN(new_n864));
  INV_X1    g678(.A(new_n864), .ZN(new_n865));
  NAND3_X1  g679(.A1(new_n849), .A2(new_n860), .A3(new_n865), .ZN(new_n866));
  INV_X1    g680(.A(KEYINPUT53), .ZN(new_n867));
  NAND2_X1  g681(.A1(new_n866), .A2(new_n867), .ZN(new_n868));
  INV_X1    g682(.A(KEYINPUT54), .ZN(new_n869));
  NAND4_X1  g683(.A1(new_n849), .A2(new_n860), .A3(new_n865), .A4(KEYINPUT53), .ZN(new_n870));
  NAND3_X1  g684(.A1(new_n868), .A2(new_n869), .A3(new_n870), .ZN(new_n871));
  INV_X1    g685(.A(KEYINPUT114), .ZN(new_n872));
  NAND2_X1  g686(.A1(new_n871), .A2(new_n872), .ZN(new_n873));
  NAND4_X1  g687(.A1(new_n868), .A2(KEYINPUT114), .A3(new_n869), .A4(new_n870), .ZN(new_n874));
  NAND2_X1  g688(.A1(new_n873), .A2(new_n874), .ZN(new_n875));
  AOI21_X1  g689(.A(KEYINPUT113), .B1(new_n868), .B2(new_n870), .ZN(new_n876));
  INV_X1    g690(.A(KEYINPUT113), .ZN(new_n877));
  AOI21_X1  g691(.A(new_n877), .B1(new_n866), .B2(new_n867), .ZN(new_n878));
  OAI21_X1  g692(.A(KEYINPUT54), .B1(new_n876), .B2(new_n878), .ZN(new_n879));
  NAND2_X1  g693(.A1(new_n875), .A2(new_n879), .ZN(new_n880));
  OAI22_X1  g694(.A1(new_n838), .A2(new_n880), .B1(G952), .B2(G953), .ZN(new_n881));
  XOR2_X1   g695(.A(new_n818), .B(KEYINPUT49), .Z(new_n882));
  NAND3_X1  g696(.A1(new_n641), .A2(new_n398), .A3(new_n628), .ZN(new_n883));
  OR4_X1    g697(.A1(new_n725), .A2(new_n882), .A3(new_n791), .A4(new_n883), .ZN(new_n884));
  OAI21_X1  g698(.A(new_n881), .B1(new_n721), .B2(new_n884), .ZN(G75));
  NOR2_X1   g699(.A1(new_n232), .A2(G952), .ZN(new_n886));
  INV_X1    g700(.A(new_n886), .ZN(new_n887));
  NAND2_X1  g701(.A1(new_n868), .A2(new_n870), .ZN(new_n888));
  NAND2_X1  g702(.A1(new_n888), .A2(new_n190), .ZN(new_n889));
  NOR2_X1   g703(.A1(new_n889), .A2(new_n455), .ZN(new_n890));
  NAND2_X1  g704(.A1(new_n444), .A2(new_n446), .ZN(new_n891));
  NAND2_X1  g705(.A1(new_n891), .A2(new_n452), .ZN(new_n892));
  NAND2_X1  g706(.A1(new_n892), .A2(new_n454), .ZN(new_n893));
  XNOR2_X1  g707(.A(new_n893), .B(KEYINPUT55), .ZN(new_n894));
  OR2_X1    g708(.A1(new_n894), .A2(KEYINPUT56), .ZN(new_n895));
  OAI21_X1  g709(.A(new_n887), .B1(new_n890), .B2(new_n895), .ZN(new_n896));
  OR2_X1    g710(.A1(new_n890), .A2(KEYINPUT116), .ZN(new_n897));
  INV_X1    g711(.A(KEYINPUT56), .ZN(new_n898));
  NAND2_X1  g712(.A1(new_n890), .A2(KEYINPUT116), .ZN(new_n899));
  NAND3_X1  g713(.A1(new_n897), .A2(new_n898), .A3(new_n899), .ZN(new_n900));
  AOI21_X1  g714(.A(new_n896), .B1(new_n900), .B2(new_n894), .ZN(G51));
  NAND2_X1  g715(.A1(new_n888), .A2(KEYINPUT54), .ZN(new_n902));
  NAND2_X1  g716(.A1(new_n902), .A2(new_n871), .ZN(new_n903));
  XNOR2_X1  g717(.A(new_n618), .B(KEYINPUT117), .ZN(new_n904));
  XNOR2_X1  g718(.A(new_n904), .B(KEYINPUT57), .ZN(new_n905));
  AOI21_X1  g719(.A(new_n742), .B1(new_n903), .B2(new_n905), .ZN(new_n906));
  NOR2_X1   g720(.A1(new_n889), .A2(new_n784), .ZN(new_n907));
  OAI21_X1  g721(.A(new_n887), .B1(new_n906), .B2(new_n907), .ZN(new_n908));
  INV_X1    g722(.A(KEYINPUT118), .ZN(new_n909));
  NAND2_X1  g723(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  OAI211_X1 g724(.A(KEYINPUT118), .B(new_n887), .C1(new_n906), .C2(new_n907), .ZN(new_n911));
  NAND2_X1  g725(.A1(new_n910), .A2(new_n911), .ZN(G54));
  INV_X1    g726(.A(new_n519), .ZN(new_n913));
  NAND2_X1  g727(.A1(KEYINPUT58), .A2(G475), .ZN(new_n914));
  OR3_X1    g728(.A1(new_n889), .A2(new_n913), .A3(new_n914), .ZN(new_n915));
  OAI21_X1  g729(.A(new_n913), .B1(new_n889), .B2(new_n914), .ZN(new_n916));
  NAND3_X1  g730(.A1(new_n915), .A2(new_n887), .A3(new_n916), .ZN(new_n917));
  XNOR2_X1  g731(.A(new_n917), .B(KEYINPUT119), .ZN(G60));
  NAND2_X1  g732(.A1(new_n653), .A2(new_n654), .ZN(new_n919));
  XNOR2_X1  g733(.A(new_n919), .B(KEYINPUT120), .ZN(new_n920));
  XNOR2_X1  g734(.A(KEYINPUT121), .B(KEYINPUT59), .ZN(new_n921));
  NOR2_X1   g735(.A1(new_n570), .A2(new_n475), .ZN(new_n922));
  XNOR2_X1  g736(.A(new_n921), .B(new_n922), .ZN(new_n923));
  AND2_X1   g737(.A1(new_n920), .A2(new_n923), .ZN(new_n924));
  AOI21_X1  g738(.A(new_n886), .B1(new_n903), .B2(new_n924), .ZN(new_n925));
  INV_X1    g739(.A(new_n923), .ZN(new_n926));
  AOI21_X1  g740(.A(new_n926), .B1(new_n875), .B2(new_n879), .ZN(new_n927));
  OAI21_X1  g741(.A(new_n925), .B1(new_n927), .B2(new_n920), .ZN(new_n928));
  NAND2_X1  g742(.A1(new_n928), .A2(KEYINPUT122), .ZN(new_n929));
  INV_X1    g743(.A(KEYINPUT122), .ZN(new_n930));
  OAI211_X1 g744(.A(new_n930), .B(new_n925), .C1(new_n927), .C2(new_n920), .ZN(new_n931));
  NAND2_X1  g745(.A1(new_n929), .A2(new_n931), .ZN(G63));
  NAND2_X1  g746(.A1(G217), .A2(G902), .ZN(new_n933));
  XNOR2_X1  g747(.A(new_n933), .B(KEYINPUT60), .ZN(new_n934));
  AOI21_X1  g748(.A(new_n934), .B1(new_n868), .B2(new_n870), .ZN(new_n935));
  XOR2_X1   g749(.A(new_n681), .B(KEYINPUT123), .Z(new_n936));
  NAND2_X1  g750(.A1(new_n935), .A2(new_n936), .ZN(new_n937));
  OAI211_X1 g751(.A(new_n937), .B(new_n887), .C1(new_n247), .C2(new_n935), .ZN(new_n938));
  INV_X1    g752(.A(KEYINPUT124), .ZN(new_n939));
  AOI21_X1  g753(.A(KEYINPUT61), .B1(new_n937), .B2(new_n939), .ZN(new_n940));
  XNOR2_X1  g754(.A(new_n938), .B(new_n940), .ZN(G66));
  NAND2_X1  g755(.A1(G224), .A2(G953), .ZN(new_n942));
  NOR2_X1   g756(.A1(new_n538), .A2(new_n942), .ZN(new_n943));
  AOI21_X1  g757(.A(new_n943), .B1(new_n849), .B2(new_n232), .ZN(new_n944));
  OAI21_X1  g758(.A(new_n891), .B1(G898), .B2(new_n232), .ZN(new_n945));
  XNOR2_X1  g759(.A(new_n944), .B(new_n945), .ZN(G69));
  NAND2_X1  g760(.A1(new_n353), .A2(new_n354), .ZN(new_n947));
  NAND2_X1  g761(.A1(new_n947), .A2(new_n341), .ZN(new_n948));
  XNOR2_X1  g762(.A(new_n948), .B(new_n509), .ZN(new_n949));
  AND2_X1   g763(.A1(new_n851), .A2(new_n738), .ZN(new_n950));
  AND3_X1   g764(.A1(new_n950), .A2(new_n774), .A3(new_n778), .ZN(new_n951));
  NAND3_X1  g765(.A1(new_n790), .A2(new_n397), .A3(new_n852), .ZN(new_n952));
  AND4_X1   g766(.A1(new_n799), .A2(new_n951), .A3(new_n806), .A4(new_n952), .ZN(new_n953));
  NOR2_X1   g767(.A1(new_n953), .A2(G953), .ZN(new_n954));
  NAND2_X1  g768(.A1(new_n704), .A2(G953), .ZN(new_n955));
  XNOR2_X1  g769(.A(new_n955), .B(KEYINPUT125), .ZN(new_n956));
  OAI21_X1  g770(.A(new_n949), .B1(new_n954), .B2(new_n956), .ZN(new_n957));
  AOI21_X1  g771(.A(new_n659), .B1(new_n572), .B2(new_n534), .ZN(new_n958));
  NOR3_X1   g772(.A1(new_n723), .A2(new_n797), .A3(new_n958), .ZN(new_n959));
  NAND2_X1  g773(.A1(new_n397), .A2(new_n959), .ZN(new_n960));
  AND3_X1   g774(.A1(new_n806), .A2(new_n799), .A3(new_n960), .ZN(new_n961));
  INV_X1    g775(.A(KEYINPUT62), .ZN(new_n962));
  NAND4_X1  g776(.A1(new_n731), .A2(new_n962), .A3(new_n732), .A4(new_n950), .ZN(new_n963));
  AND2_X1   g777(.A1(new_n961), .A2(new_n963), .ZN(new_n964));
  NAND3_X1  g778(.A1(new_n731), .A2(new_n732), .A3(new_n950), .ZN(new_n965));
  NAND2_X1  g779(.A1(new_n965), .A2(KEYINPUT62), .ZN(new_n966));
  AOI21_X1  g780(.A(G953), .B1(new_n964), .B2(new_n966), .ZN(new_n967));
  OAI21_X1  g781(.A(new_n957), .B1(new_n967), .B2(new_n949), .ZN(new_n968));
  AOI21_X1  g782(.A(new_n232), .B1(G227), .B2(G900), .ZN(new_n969));
  XNOR2_X1  g783(.A(new_n968), .B(new_n969), .ZN(G72));
  NOR2_X1   g784(.A1(new_n876), .A2(new_n878), .ZN(new_n971));
  NOR2_X1   g785(.A1(new_n391), .A2(new_n336), .ZN(new_n972));
  INV_X1    g786(.A(new_n972), .ZN(new_n973));
  NAND2_X1  g787(.A1(G472), .A2(G902), .ZN(new_n974));
  XOR2_X1   g788(.A(new_n974), .B(KEYINPUT63), .Z(new_n975));
  NAND3_X1  g789(.A1(new_n973), .A2(new_n715), .A3(new_n975), .ZN(new_n976));
  NOR2_X1   g790(.A1(new_n971), .A2(new_n976), .ZN(new_n977));
  INV_X1    g791(.A(new_n975), .ZN(new_n978));
  AOI21_X1  g792(.A(new_n978), .B1(new_n953), .B2(new_n849), .ZN(new_n979));
  OAI21_X1  g793(.A(new_n887), .B1(new_n979), .B2(new_n973), .ZN(new_n980));
  NAND4_X1  g794(.A1(new_n966), .A2(new_n961), .A3(new_n849), .A4(new_n963), .ZN(new_n981));
  AOI21_X1  g795(.A(new_n715), .B1(new_n981), .B2(new_n975), .ZN(new_n982));
  OR4_X1    g796(.A1(KEYINPUT126), .A2(new_n977), .A3(new_n980), .A4(new_n982), .ZN(new_n983));
  OR2_X1    g797(.A1(new_n980), .A2(new_n982), .ZN(new_n984));
  OAI21_X1  g798(.A(KEYINPUT126), .B1(new_n984), .B2(new_n977), .ZN(new_n985));
  NAND2_X1  g799(.A1(new_n983), .A2(new_n985), .ZN(G57));
endmodule


