

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359,
         n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370,
         n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381,
         n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392,
         n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403,
         n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414,
         n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425,
         n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436,
         n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447,
         n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458,
         n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469,
         n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480,
         n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491,
         n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502,
         n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n513,
         n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
         n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
         n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590,
         n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601,
         n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612,
         n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623,
         n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634,
         n635, n636, n637, n638, n639, n640, n641, n642, n643, n644, n645,
         n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, n656,
         n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n667,
         n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678,
         n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689,
         n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700,
         n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711,
         n712, n713, n714, n715, n716, n717, n718, n719, n720, n721, n722,
         n723, n724, n725, n726, n727, n728, n729, n730, n731, n732, n733,
         n734, n735, n736, n737, n738, n739, n740, n741, n742, n743, n744,
         n745, n746, n747, n748, n749, n750, n751, n752, n753, n754, n755,
         n756, n757, n758, n759, n760, n761, n762, n763, n764, n765, n766;

  BUF_X1 U371 ( .A(n721), .Z(n730) );
  XNOR2_X1 U372 ( .A(n555), .B(KEYINPUT1), .ZN(n537) );
  INV_X1 U373 ( .A(G953), .ZN(n754) );
  NOR2_X2 U374 ( .A1(n678), .A2(n576), .ZN(n683) );
  XNOR2_X2 U375 ( .A(n583), .B(KEYINPUT42), .ZN(n765) );
  XNOR2_X2 U376 ( .A(n486), .B(n485), .ZN(n576) );
  XNOR2_X2 U377 ( .A(n491), .B(n441), .ZN(n722) );
  XNOR2_X2 U378 ( .A(n750), .B(G146), .ZN(n491) );
  INV_X2 U379 ( .A(G143), .ZN(n437) );
  XNOR2_X1 U380 ( .A(n440), .B(n438), .ZN(n763) );
  BUF_X1 U381 ( .A(n537), .Z(n351) );
  NOR2_X1 U382 ( .A1(n578), .A2(n594), .ZN(n579) );
  NAND2_X1 U383 ( .A1(n372), .A2(n369), .ZN(n762) );
  NAND2_X1 U384 ( .A1(n371), .A2(n370), .ZN(n369) );
  NOR2_X1 U385 ( .A1(n376), .A2(n763), .ZN(n368) );
  AND2_X1 U386 ( .A1(n374), .A2(n373), .ZN(n372) );
  NAND2_X1 U387 ( .A1(n400), .A2(n398), .ZN(n698) );
  XNOR2_X1 U388 ( .A(n542), .B(n541), .ZN(n548) );
  NOR2_X1 U389 ( .A1(n402), .A2(n401), .ZN(n400) );
  NAND2_X1 U390 ( .A1(n422), .A2(n428), .ZN(n401) );
  NAND2_X1 U391 ( .A1(n537), .A2(n683), .ZN(n487) );
  NAND2_X1 U392 ( .A1(n412), .A2(n409), .ZN(n603) );
  AND2_X1 U393 ( .A1(n364), .A2(n363), .ZN(n362) );
  AND2_X1 U394 ( .A1(n414), .A2(n413), .ZN(n412) );
  XNOR2_X1 U395 ( .A(n716), .B(n715), .ZN(n718) );
  OR2_X1 U396 ( .A1(n633), .A2(G902), .ZN(n450) );
  XNOR2_X1 U397 ( .A(KEYINPUT67), .B(G101), .ZN(n465) );
  XNOR2_X1 U398 ( .A(G137), .B(G140), .ZN(n474) );
  XNOR2_X1 U399 ( .A(n502), .B(n501), .ZN(n349) );
  XNOR2_X1 U400 ( .A(n502), .B(n501), .ZN(n666) );
  XNOR2_X1 U401 ( .A(n566), .B(n565), .ZN(n350) );
  XNOR2_X1 U402 ( .A(n566), .B(n565), .ZN(n737) );
  NOR2_X1 U403 ( .A1(n736), .A2(n636), .ZN(n639) );
  INV_X1 U404 ( .A(G107), .ZN(n417) );
  XNOR2_X1 U405 ( .A(G104), .B(G110), .ZN(n418) );
  XNOR2_X1 U406 ( .A(n505), .B(KEYINPUT10), .ZN(n475) );
  XNOR2_X1 U407 ( .A(n614), .B(KEYINPUT110), .ZN(n392) );
  XNOR2_X1 U408 ( .A(n534), .B(n535), .ZN(n552) );
  NAND2_X1 U409 ( .A1(n365), .A2(G902), .ZN(n363) );
  NAND2_X1 U410 ( .A1(n420), .A2(n467), .ZN(n419) );
  NAND2_X1 U411 ( .A1(n488), .A2(n466), .ZN(n420) );
  NAND2_X1 U412 ( .A1(n603), .A2(n582), .ZN(n598) );
  XNOR2_X1 U413 ( .A(KEYINPUT82), .B(KEYINPUT36), .ZN(n599) );
  NAND2_X1 U414 ( .A1(n574), .A2(n573), .ZN(n601) );
  NOR2_X1 U415 ( .A1(n575), .A2(n572), .ZN(n574) );
  NAND2_X1 U416 ( .A1(n611), .A2(n379), .ZN(n612) );
  XNOR2_X1 U417 ( .A(n586), .B(n452), .ZN(n611) );
  INV_X1 U418 ( .A(KEYINPUT69), .ZN(n380) );
  NAND2_X1 U419 ( .A1(n670), .A2(n431), .ZN(n430) );
  NAND2_X1 U420 ( .A1(n668), .A2(KEYINPUT109), .ZN(n434) );
  XNOR2_X1 U421 ( .A(KEYINPUT4), .B(KEYINPUT17), .ZN(n436) );
  XOR2_X1 U422 ( .A(KEYINPUT73), .B(KEYINPUT34), .Z(n524) );
  XNOR2_X1 U423 ( .A(n512), .B(n381), .ZN(n744) );
  XNOR2_X1 U424 ( .A(n382), .B(G122), .ZN(n381) );
  INV_X1 U425 ( .A(KEYINPUT16), .ZN(n382) );
  XNOR2_X1 U426 ( .A(n447), .B(n446), .ZN(n529) );
  INV_X1 U427 ( .A(KEYINPUT8), .ZN(n446) );
  NAND2_X1 U428 ( .A1(n754), .A2(G234), .ZN(n447) );
  XNOR2_X1 U429 ( .A(n476), .B(n395), .ZN(n394) );
  XNOR2_X1 U430 ( .A(G119), .B(KEYINPUT89), .ZN(n476) );
  XNOR2_X1 U431 ( .A(KEYINPUT23), .B(KEYINPUT24), .ZN(n395) );
  INV_X1 U432 ( .A(KEYINPUT88), .ZN(n477) );
  XNOR2_X1 U433 ( .A(G128), .B(G110), .ZN(n478) );
  XNOR2_X1 U434 ( .A(n475), .B(n474), .ZN(n751) );
  XNOR2_X1 U435 ( .A(G116), .B(KEYINPUT9), .ZN(n526) );
  XNOR2_X1 U436 ( .A(n528), .B(n527), .ZN(n405) );
  XNOR2_X1 U437 ( .A(G107), .B(G122), .ZN(n527) );
  XNOR2_X1 U438 ( .A(n461), .B(n460), .ZN(n462) );
  NAND2_X1 U439 ( .A1(n709), .A2(n623), .ZN(n624) );
  NAND2_X1 U440 ( .A1(n389), .A2(n355), .ZN(n388) );
  INV_X1 U441 ( .A(n599), .ZN(n387) );
  NAND2_X1 U442 ( .A1(n602), .A2(n375), .ZN(n373) );
  NAND2_X1 U443 ( .A1(n411), .A2(n410), .ZN(n409) );
  AND2_X1 U444 ( .A1(n515), .A2(n503), .ZN(n410) );
  XNOR2_X1 U445 ( .A(n445), .B(n444), .ZN(n553) );
  INV_X1 U446 ( .A(G478), .ZN(n444) );
  XNOR2_X1 U447 ( .A(n397), .B(n396), .ZN(n573) );
  INV_X1 U448 ( .A(KEYINPUT92), .ZN(n396) );
  XNOR2_X1 U449 ( .A(n504), .B(n442), .ZN(n441) );
  XNOR2_X1 U450 ( .A(n468), .B(n443), .ZN(n442) );
  NOR2_X1 U451 ( .A1(G952), .A2(n754), .ZN(n736) );
  INV_X1 U452 ( .A(KEYINPUT78), .ZN(n378) );
  NOR2_X1 U453 ( .A1(G953), .A2(G237), .ZN(n494) );
  NAND2_X1 U454 ( .A1(n427), .A2(n433), .ZN(n432) );
  NAND2_X1 U455 ( .A1(n470), .A2(n361), .ZN(n360) );
  INV_X1 U456 ( .A(G902), .ZN(n361) );
  XOR2_X1 U457 ( .A(KEYINPUT75), .B(G137), .Z(n489) );
  XOR2_X1 U458 ( .A(G122), .B(G104), .Z(n454) );
  XNOR2_X1 U459 ( .A(G113), .B(G140), .ZN(n453) );
  XNOR2_X1 U460 ( .A(n459), .B(n458), .ZN(n460) );
  INV_X1 U461 ( .A(KEYINPUT12), .ZN(n458) );
  XNOR2_X1 U462 ( .A(G131), .B(G143), .ZN(n459) );
  INV_X1 U463 ( .A(KEYINPUT72), .ZN(n466) );
  XNOR2_X1 U464 ( .A(G131), .B(KEYINPUT4), .ZN(n464) );
  INV_X1 U465 ( .A(n664), .ZN(n408) );
  NAND2_X1 U466 ( .A1(n538), .A2(KEYINPUT41), .ZN(n428) );
  AND2_X1 U467 ( .A1(n432), .A2(KEYINPUT41), .ZN(n399) );
  NOR2_X1 U468 ( .A1(n430), .A2(n426), .ZN(n425) );
  XNOR2_X1 U469 ( .A(n617), .B(n567), .ZN(n667) );
  INV_X1 U470 ( .A(KEYINPUT38), .ZN(n567) );
  NAND2_X1 U471 ( .A1(n415), .A2(n623), .ZN(n413) );
  XNOR2_X1 U472 ( .A(n622), .B(KEYINPUT80), .ZN(n752) );
  INV_X1 U473 ( .A(KEYINPUT45), .ZN(n565) );
  XNOR2_X1 U474 ( .A(n474), .B(KEYINPUT87), .ZN(n443) );
  XNOR2_X1 U475 ( .A(n513), .B(n416), .ZN(n714) );
  NAND2_X1 U476 ( .A1(n752), .A2(n702), .ZN(n709) );
  INV_X1 U477 ( .A(n603), .ZN(n617) );
  XNOR2_X1 U478 ( .A(n449), .B(n448), .ZN(n584) );
  INV_X1 U479 ( .A(KEYINPUT39), .ZN(n448) );
  NOR2_X1 U480 ( .A1(n601), .A2(n667), .ZN(n449) );
  XNOR2_X1 U481 ( .A(n598), .B(KEYINPUT19), .ZN(n588) );
  XNOR2_X1 U482 ( .A(n552), .B(KEYINPUT99), .ZN(n554) );
  OR2_X1 U483 ( .A1(n554), .A2(n553), .ZN(n595) );
  XNOR2_X1 U484 ( .A(n751), .B(n393), .ZN(n481) );
  XNOR2_X1 U485 ( .A(n479), .B(n394), .ZN(n393) );
  XNOR2_X1 U486 ( .A(n404), .B(n403), .ZN(n728) );
  XNOR2_X1 U487 ( .A(n530), .B(n405), .ZN(n404) );
  NAND2_X1 U488 ( .A1(n721), .A2(G475), .ZN(n626) );
  AND2_X1 U489 ( .A1(n600), .A2(n391), .ZN(n390) );
  NOR2_X1 U490 ( .A1(n602), .A2(n375), .ZN(n370) );
  XNOR2_X1 U491 ( .A(n439), .B(KEYINPUT32), .ZN(n438) );
  OR2_X2 U492 ( .A1(n548), .A2(n547), .ZN(n440) );
  INV_X1 U493 ( .A(KEYINPUT64), .ZN(n439) );
  NOR2_X1 U494 ( .A1(n601), .A2(n602), .ZN(n604) );
  INV_X1 U495 ( .A(n595), .ZN(n655) );
  XNOR2_X1 U496 ( .A(n725), .B(n724), .ZN(n726) );
  XNOR2_X1 U497 ( .A(n722), .B(n723), .ZN(n724) );
  XNOR2_X1 U498 ( .A(n419), .B(n742), .ZN(n504) );
  XOR2_X1 U499 ( .A(n526), .B(KEYINPUT7), .Z(n352) );
  NOR2_X1 U500 ( .A1(n553), .A2(n552), .ZN(n670) );
  AND2_X1 U501 ( .A1(n408), .A2(n764), .ZN(n353) );
  NAND2_X2 U502 ( .A1(n362), .A2(n359), .ZN(n555) );
  OR2_X1 U503 ( .A1(n671), .A2(n562), .ZN(n354) );
  OR2_X1 U504 ( .A1(n598), .A2(n599), .ZN(n355) );
  AND2_X1 U505 ( .A1(n421), .A2(n434), .ZN(n356) );
  OR2_X1 U506 ( .A1(n430), .A2(n434), .ZN(n357) );
  NAND2_X1 U507 ( .A1(n385), .A2(n390), .ZN(n662) );
  XOR2_X1 U508 ( .A(KEYINPUT66), .B(KEYINPUT0), .Z(n358) );
  XNOR2_X1 U509 ( .A(n418), .B(n417), .ZN(n742) );
  OR2_X1 U510 ( .A1(n722), .A2(n360), .ZN(n359) );
  NAND2_X1 U511 ( .A1(n722), .A2(n365), .ZN(n364) );
  INV_X1 U512 ( .A(n470), .ZN(n365) );
  XNOR2_X2 U513 ( .A(n366), .B(n464), .ZN(n750) );
  XNOR2_X1 U514 ( .A(n352), .B(n366), .ZN(n403) );
  XNOR2_X2 U515 ( .A(n406), .B(G134), .ZN(n366) );
  XNOR2_X1 U516 ( .A(n367), .B(n407), .ZN(n564) );
  NAND2_X1 U517 ( .A1(n368), .A2(n762), .ZN(n367) );
  INV_X1 U518 ( .A(n536), .ZN(n371) );
  NAND2_X1 U519 ( .A1(n536), .A2(n375), .ZN(n374) );
  INV_X1 U520 ( .A(KEYINPUT35), .ZN(n375) );
  INV_X1 U521 ( .A(n648), .ZN(n376) );
  NAND2_X1 U522 ( .A1(n377), .A2(n593), .ZN(n609) );
  XNOR2_X1 U523 ( .A(n589), .B(n378), .ZN(n377) );
  XNOR2_X1 U524 ( .A(n610), .B(n380), .ZN(n379) );
  NOR2_X1 U525 ( .A1(n628), .A2(n736), .ZN(n631) );
  NAND2_X1 U526 ( .A1(n383), .A2(n353), .ZN(n622) );
  XNOR2_X1 U527 ( .A(n612), .B(n384), .ZN(n383) );
  INV_X1 U528 ( .A(KEYINPUT48), .ZN(n384) );
  NAND2_X1 U529 ( .A1(n388), .A2(n386), .ZN(n385) );
  NAND2_X1 U530 ( .A1(n392), .A2(n387), .ZN(n386) );
  INV_X1 U531 ( .A(n392), .ZN(n389) );
  NAND2_X1 U532 ( .A1(n598), .A2(n599), .ZN(n391) );
  XNOR2_X2 U533 ( .A(G146), .B(G125), .ZN(n505) );
  NAND2_X1 U534 ( .A1(n683), .A2(n555), .ZN(n397) );
  NAND2_X1 U535 ( .A1(n698), .A2(n587), .ZN(n583) );
  NAND2_X1 U536 ( .A1(n399), .A2(n356), .ZN(n398) );
  NAND2_X1 U537 ( .A1(n429), .A2(n357), .ZN(n402) );
  XNOR2_X1 U538 ( .A(n406), .B(n436), .ZN(n509) );
  XNOR2_X2 U539 ( .A(n437), .B(G128), .ZN(n406) );
  INV_X1 U540 ( .A(KEYINPUT44), .ZN(n407) );
  INV_X1 U541 ( .A(n714), .ZN(n411) );
  NAND2_X1 U542 ( .A1(n714), .A2(n415), .ZN(n414) );
  INV_X1 U543 ( .A(n515), .ZN(n415) );
  INV_X1 U544 ( .A(n744), .ZN(n416) );
  INV_X1 U545 ( .A(n465), .ZN(n488) );
  INV_X1 U546 ( .A(n667), .ZN(n427) );
  NAND2_X1 U547 ( .A1(n667), .A2(KEYINPUT109), .ZN(n421) );
  NAND2_X1 U548 ( .A1(n423), .A2(n667), .ZN(n422) );
  NOR2_X1 U549 ( .A1(n430), .A2(n424), .ZN(n423) );
  INV_X1 U550 ( .A(KEYINPUT109), .ZN(n424) );
  NAND2_X1 U551 ( .A1(n427), .A2(n425), .ZN(n429) );
  INV_X1 U552 ( .A(n433), .ZN(n426) );
  NAND2_X1 U553 ( .A1(n356), .A2(n432), .ZN(n673) );
  INV_X1 U554 ( .A(KEYINPUT41), .ZN(n431) );
  NOR2_X1 U555 ( .A1(n668), .A2(KEYINPUT109), .ZN(n433) );
  XNOR2_X2 U556 ( .A(n435), .B(n358), .ZN(n559) );
  NAND2_X1 U557 ( .A1(n588), .A2(n523), .ZN(n435) );
  NOR2_X1 U558 ( .A1(n728), .A2(G902), .ZN(n445) );
  NAND2_X1 U559 ( .A1(n584), .A2(n655), .ZN(n585) );
  XNOR2_X2 U560 ( .A(n450), .B(G472), .ZN(n570) );
  XNOR2_X1 U561 ( .A(n491), .B(n451), .ZN(n633) );
  XNOR2_X1 U562 ( .A(n498), .B(n490), .ZN(n451) );
  NOR2_X2 U563 ( .A1(n620), .A2(n702), .ZN(n704) );
  XNOR2_X1 U564 ( .A(KEYINPUT46), .B(KEYINPUT81), .ZN(n452) );
  XNOR2_X1 U565 ( .A(n508), .B(n507), .ZN(n510) );
  XNOR2_X1 U566 ( .A(n489), .B(n488), .ZN(n490) );
  XNOR2_X1 U567 ( .A(n478), .B(n477), .ZN(n479) );
  XNOR2_X1 U568 ( .A(n469), .B(G469), .ZN(n470) );
  XNOR2_X1 U569 ( .A(n514), .B(KEYINPUT86), .ZN(n515) );
  INV_X1 U570 ( .A(n576), .ZN(n543) );
  XNOR2_X1 U571 ( .A(n732), .B(n731), .ZN(n733) );
  XNOR2_X1 U572 ( .A(n637), .B(KEYINPUT83), .ZN(n638) );
  XNOR2_X1 U573 ( .A(n734), .B(n733), .ZN(n735) );
  XNOR2_X1 U574 ( .A(n454), .B(n453), .ZN(n455) );
  XNOR2_X1 U575 ( .A(n475), .B(n455), .ZN(n463) );
  XOR2_X1 U576 ( .A(KEYINPUT96), .B(KEYINPUT11), .Z(n457) );
  NAND2_X1 U577 ( .A1(G214), .A2(n494), .ZN(n456) );
  XNOR2_X1 U578 ( .A(n457), .B(n456), .ZN(n461) );
  XNOR2_X1 U579 ( .A(n463), .B(n462), .ZN(n533) );
  XOR2_X1 U580 ( .A(n533), .B(KEYINPUT59), .Z(n627) );
  NAND2_X1 U581 ( .A1(n465), .A2(KEYINPUT72), .ZN(n467) );
  AND2_X1 U582 ( .A1(G227), .A2(n754), .ZN(n468) );
  XNOR2_X1 U583 ( .A(KEYINPUT70), .B(KEYINPUT71), .ZN(n469) );
  XOR2_X1 U584 ( .A(KEYINPUT91), .B(KEYINPUT21), .Z(n473) );
  XNOR2_X1 U585 ( .A(G902), .B(KEYINPUT15), .ZN(n503) );
  NAND2_X1 U586 ( .A1(G234), .A2(n503), .ZN(n471) );
  XNOR2_X1 U587 ( .A(KEYINPUT20), .B(n471), .ZN(n482) );
  NAND2_X1 U588 ( .A1(n482), .A2(G221), .ZN(n472) );
  XNOR2_X1 U589 ( .A(n473), .B(n472), .ZN(n678) );
  NAND2_X1 U590 ( .A1(G221), .A2(n529), .ZN(n480) );
  XNOR2_X1 U591 ( .A(n481), .B(n480), .ZN(n732) );
  NOR2_X1 U592 ( .A1(n732), .A2(G902), .ZN(n486) );
  XOR2_X1 U593 ( .A(KEYINPUT90), .B(KEYINPUT25), .Z(n484) );
  NAND2_X1 U594 ( .A1(n482), .A2(G217), .ZN(n483) );
  XNOR2_X1 U595 ( .A(n484), .B(n483), .ZN(n485) );
  XNOR2_X2 U596 ( .A(n487), .B(KEYINPUT74), .ZN(n557) );
  XNOR2_X1 U597 ( .A(n557), .B(KEYINPUT105), .ZN(n500) );
  XNOR2_X1 U598 ( .A(KEYINPUT102), .B(KEYINPUT6), .ZN(n499) );
  XOR2_X1 U599 ( .A(G119), .B(KEYINPUT3), .Z(n493) );
  XNOR2_X1 U600 ( .A(G116), .B(G113), .ZN(n492) );
  XNOR2_X1 U601 ( .A(n493), .B(n492), .ZN(n512) );
  XOR2_X1 U602 ( .A(KEYINPUT93), .B(KEYINPUT5), .Z(n496) );
  NAND2_X1 U603 ( .A1(n494), .A2(G210), .ZN(n495) );
  XNOR2_X1 U604 ( .A(n496), .B(n495), .ZN(n497) );
  XNOR2_X1 U605 ( .A(n512), .B(n497), .ZN(n498) );
  XOR2_X1 U606 ( .A(n499), .B(n570), .Z(n596) );
  NAND2_X1 U607 ( .A1(n500), .A2(n596), .ZN(n502) );
  XNOR2_X1 U608 ( .A(KEYINPUT33), .B(KEYINPUT106), .ZN(n501) );
  INV_X1 U609 ( .A(n503), .ZN(n623) );
  XNOR2_X1 U610 ( .A(KEYINPUT76), .B(KEYINPUT18), .ZN(n506) );
  XNOR2_X1 U611 ( .A(n506), .B(n505), .ZN(n508) );
  NAND2_X1 U612 ( .A1(n754), .A2(G224), .ZN(n507) );
  XNOR2_X1 U613 ( .A(n510), .B(n509), .ZN(n511) );
  XNOR2_X1 U614 ( .A(n504), .B(n511), .ZN(n513) );
  OR2_X1 U615 ( .A1(G237), .A2(G902), .ZN(n516) );
  NAND2_X1 U616 ( .A1(G210), .A2(n516), .ZN(n514) );
  NAND2_X1 U617 ( .A1(G214), .A2(n516), .ZN(n582) );
  AND2_X1 U618 ( .A1(G953), .A2(G898), .ZN(n522) );
  NAND2_X1 U619 ( .A1(G234), .A2(G237), .ZN(n517) );
  XNOR2_X1 U620 ( .A(n517), .B(KEYINPUT14), .ZN(n665) );
  OR2_X1 U621 ( .A1(n754), .A2(G902), .ZN(n518) );
  NAND2_X1 U622 ( .A1(n665), .A2(n518), .ZN(n520) );
  NOR2_X1 U623 ( .A1(G953), .A2(G952), .ZN(n519) );
  NOR2_X1 U624 ( .A1(n520), .A2(n519), .ZN(n569) );
  INV_X1 U625 ( .A(n569), .ZN(n521) );
  NOR2_X1 U626 ( .A1(n522), .A2(n521), .ZN(n523) );
  NAND2_X1 U627 ( .A1(n666), .A2(n559), .ZN(n525) );
  XNOR2_X1 U628 ( .A(n525), .B(n524), .ZN(n536) );
  XOR2_X1 U629 ( .A(KEYINPUT101), .B(KEYINPUT100), .Z(n528) );
  NAND2_X1 U630 ( .A1(G217), .A2(n529), .ZN(n530) );
  XOR2_X1 U631 ( .A(KEYINPUT97), .B(KEYINPUT13), .Z(n532) );
  XNOR2_X1 U632 ( .A(KEYINPUT98), .B(G475), .ZN(n531) );
  XNOR2_X1 U633 ( .A(n532), .B(n531), .ZN(n535) );
  NOR2_X1 U634 ( .A1(G902), .A2(n533), .ZN(n534) );
  NAND2_X1 U635 ( .A1(n553), .A2(n552), .ZN(n602) );
  INV_X1 U636 ( .A(n670), .ZN(n538) );
  NOR2_X1 U637 ( .A1(n678), .A2(n538), .ZN(n539) );
  XOR2_X1 U638 ( .A(KEYINPUT103), .B(n539), .Z(n540) );
  AND2_X2 U639 ( .A1(n540), .A2(n559), .ZN(n542) );
  XNOR2_X1 U640 ( .A(KEYINPUT65), .B(KEYINPUT22), .ZN(n541) );
  NOR2_X1 U641 ( .A1(n351), .A2(n548), .ZN(n551) );
  INV_X1 U642 ( .A(n570), .ZN(n578) );
  NOR2_X1 U643 ( .A1(n570), .A2(n543), .ZN(n544) );
  NAND2_X1 U644 ( .A1(n551), .A2(n544), .ZN(n648) );
  XOR2_X1 U645 ( .A(KEYINPUT85), .B(n351), .Z(n600) );
  INV_X1 U646 ( .A(n600), .ZN(n546) );
  XOR2_X1 U647 ( .A(n576), .B(KEYINPUT104), .Z(n549) );
  OR2_X1 U648 ( .A1(n596), .A2(n549), .ZN(n545) );
  OR2_X1 U649 ( .A1(n546), .A2(n545), .ZN(n547) );
  INV_X1 U650 ( .A(n549), .ZN(n679) );
  NOR2_X1 U651 ( .A1(n679), .A2(n596), .ZN(n550) );
  NAND2_X1 U652 ( .A1(n551), .A2(n550), .ZN(n640) );
  AND2_X1 U653 ( .A1(n554), .A2(n553), .ZN(n658) );
  NOR2_X1 U654 ( .A1(n655), .A2(n658), .ZN(n671) );
  INV_X1 U655 ( .A(n555), .ZN(n581) );
  NAND2_X1 U656 ( .A1(n559), .A2(n573), .ZN(n556) );
  NOR2_X1 U657 ( .A1(n570), .A2(n556), .ZN(n645) );
  XOR2_X1 U658 ( .A(KEYINPUT31), .B(KEYINPUT95), .Z(n561) );
  NOR2_X1 U659 ( .A1(n557), .A2(n578), .ZN(n558) );
  XNOR2_X1 U660 ( .A(n558), .B(KEYINPUT94), .ZN(n689) );
  NAND2_X1 U661 ( .A1(n559), .A2(n689), .ZN(n560) );
  XNOR2_X1 U662 ( .A(n561), .B(n560), .ZN(n657) );
  NOR2_X1 U663 ( .A1(n645), .A2(n657), .ZN(n562) );
  AND2_X1 U664 ( .A1(n640), .A2(n354), .ZN(n563) );
  NAND2_X1 U665 ( .A1(n564), .A2(n563), .ZN(n566) );
  NAND2_X1 U666 ( .A1(G953), .A2(G900), .ZN(n568) );
  NAND2_X1 U667 ( .A1(n569), .A2(n568), .ZN(n575) );
  NAND2_X1 U668 ( .A1(n570), .A2(n582), .ZN(n571) );
  XNOR2_X1 U669 ( .A(KEYINPUT30), .B(n571), .ZN(n572) );
  AND2_X1 U670 ( .A1(n658), .A2(n584), .ZN(n664) );
  NOR2_X1 U671 ( .A1(n678), .A2(n575), .ZN(n577) );
  NAND2_X1 U672 ( .A1(n577), .A2(n576), .ZN(n594) );
  XOR2_X1 U673 ( .A(KEYINPUT28), .B(n579), .Z(n580) );
  NOR2_X1 U674 ( .A1(n581), .A2(n580), .ZN(n587) );
  INV_X1 U675 ( .A(n582), .ZN(n668) );
  XNOR2_X1 U676 ( .A(n585), .B(KEYINPUT40), .ZN(n766) );
  NAND2_X1 U677 ( .A1(n765), .A2(n766), .ZN(n586) );
  AND2_X1 U678 ( .A1(n587), .A2(n588), .ZN(n653) );
  INV_X1 U679 ( .A(KEYINPUT47), .ZN(n590) );
  NOR2_X1 U680 ( .A1(n653), .A2(n590), .ZN(n589) );
  XOR2_X1 U681 ( .A(KEYINPUT68), .B(n590), .Z(n591) );
  NOR2_X1 U682 ( .A1(n671), .A2(n591), .ZN(n592) );
  NAND2_X1 U683 ( .A1(n653), .A2(n592), .ZN(n593) );
  NOR2_X1 U684 ( .A1(n595), .A2(n594), .ZN(n597) );
  NAND2_X1 U685 ( .A1(n597), .A2(n596), .ZN(n614) );
  NAND2_X1 U686 ( .A1(KEYINPUT47), .A2(n671), .ZN(n605) );
  NAND2_X1 U687 ( .A1(n604), .A2(n603), .ZN(n652) );
  NAND2_X1 U688 ( .A1(n605), .A2(n652), .ZN(n606) );
  XNOR2_X1 U689 ( .A(n606), .B(KEYINPUT77), .ZN(n607) );
  NAND2_X1 U690 ( .A1(n662), .A2(n607), .ZN(n608) );
  NOR2_X1 U691 ( .A1(n609), .A2(n608), .ZN(n610) );
  OR2_X1 U692 ( .A1(n351), .A2(n668), .ZN(n613) );
  NOR2_X1 U693 ( .A1(n614), .A2(n613), .ZN(n616) );
  XNOR2_X1 U694 ( .A(KEYINPUT107), .B(KEYINPUT43), .ZN(n615) );
  XNOR2_X1 U695 ( .A(n616), .B(n615), .ZN(n618) );
  NAND2_X1 U696 ( .A1(n618), .A2(n617), .ZN(n619) );
  XNOR2_X1 U697 ( .A(n619), .B(KEYINPUT108), .ZN(n764) );
  NOR2_X2 U698 ( .A1(n737), .A2(n622), .ZN(n620) );
  INV_X1 U699 ( .A(KEYINPUT2), .ZN(n702) );
  NOR2_X1 U700 ( .A1(KEYINPUT2), .A2(n350), .ZN(n621) );
  NOR2_X1 U701 ( .A1(n704), .A2(n621), .ZN(n625) );
  NOR2_X4 U702 ( .A1(n625), .A2(n624), .ZN(n721) );
  XNOR2_X1 U703 ( .A(n627), .B(n626), .ZN(n628) );
  INV_X1 U704 ( .A(KEYINPUT123), .ZN(n629) );
  XNOR2_X1 U705 ( .A(n629), .B(KEYINPUT60), .ZN(n630) );
  XNOR2_X1 U706 ( .A(n631), .B(n630), .ZN(G60) );
  NAND2_X1 U707 ( .A1(n721), .A2(G472), .ZN(n635) );
  XOR2_X1 U708 ( .A(KEYINPUT62), .B(KEYINPUT111), .Z(n632) );
  XNOR2_X1 U709 ( .A(n633), .B(n632), .ZN(n634) );
  XNOR2_X1 U710 ( .A(n635), .B(n634), .ZN(n636) );
  XNOR2_X1 U711 ( .A(KEYINPUT63), .B(KEYINPUT112), .ZN(n637) );
  XNOR2_X1 U712 ( .A(n639), .B(n638), .ZN(G57) );
  XNOR2_X1 U713 ( .A(G101), .B(n640), .ZN(G3) );
  NAND2_X1 U714 ( .A1(n655), .A2(n645), .ZN(n641) );
  XNOR2_X1 U715 ( .A(n641), .B(G104), .ZN(G6) );
  XOR2_X1 U716 ( .A(KEYINPUT114), .B(KEYINPUT27), .Z(n643) );
  XNOR2_X1 U717 ( .A(G107), .B(KEYINPUT26), .ZN(n642) );
  XNOR2_X1 U718 ( .A(n643), .B(n642), .ZN(n644) );
  XOR2_X1 U719 ( .A(KEYINPUT113), .B(n644), .Z(n647) );
  NAND2_X1 U720 ( .A1(n645), .A2(n658), .ZN(n646) );
  XNOR2_X1 U721 ( .A(n647), .B(n646), .ZN(G9) );
  XNOR2_X1 U722 ( .A(n648), .B(G110), .ZN(G12) );
  XOR2_X1 U723 ( .A(KEYINPUT115), .B(KEYINPUT29), .Z(n650) );
  NAND2_X1 U724 ( .A1(n653), .A2(n658), .ZN(n649) );
  XNOR2_X1 U725 ( .A(n650), .B(n649), .ZN(n651) );
  XOR2_X1 U726 ( .A(G128), .B(n651), .Z(G30) );
  XNOR2_X1 U727 ( .A(G143), .B(n652), .ZN(G45) );
  NAND2_X1 U728 ( .A1(n655), .A2(n653), .ZN(n654) );
  XNOR2_X1 U729 ( .A(n654), .B(G146), .ZN(G48) );
  NAND2_X1 U730 ( .A1(n655), .A2(n657), .ZN(n656) );
  XNOR2_X1 U731 ( .A(n656), .B(G113), .ZN(G15) );
  NAND2_X1 U732 ( .A1(n658), .A2(n657), .ZN(n659) );
  XNOR2_X1 U733 ( .A(n659), .B(G116), .ZN(G18) );
  XOR2_X1 U734 ( .A(KEYINPUT116), .B(KEYINPUT117), .Z(n661) );
  XNOR2_X1 U735 ( .A(G125), .B(KEYINPUT37), .ZN(n660) );
  XNOR2_X1 U736 ( .A(n661), .B(n660), .ZN(n663) );
  XOR2_X1 U737 ( .A(n663), .B(n662), .Z(G27) );
  XOR2_X1 U738 ( .A(G134), .B(n664), .Z(G36) );
  NAND2_X1 U739 ( .A1(G952), .A2(n665), .ZN(n696) );
  NAND2_X1 U740 ( .A1(n668), .A2(n667), .ZN(n669) );
  NAND2_X1 U741 ( .A1(n670), .A2(n669), .ZN(n675) );
  INV_X1 U742 ( .A(n671), .ZN(n672) );
  NAND2_X1 U743 ( .A1(n673), .A2(n672), .ZN(n674) );
  NAND2_X1 U744 ( .A1(n675), .A2(n674), .ZN(n676) );
  NAND2_X1 U745 ( .A1(n349), .A2(n676), .ZN(n677) );
  XNOR2_X1 U746 ( .A(n677), .B(KEYINPUT120), .ZN(n693) );
  NAND2_X1 U747 ( .A1(n679), .A2(n678), .ZN(n680) );
  XNOR2_X1 U748 ( .A(KEYINPUT49), .B(n680), .ZN(n681) );
  NOR2_X1 U749 ( .A1(n570), .A2(n681), .ZN(n682) );
  XOR2_X1 U750 ( .A(KEYINPUT118), .B(n682), .Z(n686) );
  NOR2_X1 U751 ( .A1(n351), .A2(n683), .ZN(n684) );
  XNOR2_X1 U752 ( .A(KEYINPUT50), .B(n684), .ZN(n685) );
  NOR2_X1 U753 ( .A1(n686), .A2(n685), .ZN(n687) );
  XOR2_X1 U754 ( .A(KEYINPUT119), .B(n687), .Z(n688) );
  NOR2_X1 U755 ( .A1(n689), .A2(n688), .ZN(n690) );
  XNOR2_X1 U756 ( .A(KEYINPUT51), .B(n690), .ZN(n691) );
  NAND2_X1 U757 ( .A1(n691), .A2(n698), .ZN(n692) );
  NAND2_X1 U758 ( .A1(n693), .A2(n692), .ZN(n694) );
  XOR2_X1 U759 ( .A(KEYINPUT52), .B(n694), .Z(n695) );
  NOR2_X1 U760 ( .A1(n696), .A2(n695), .ZN(n697) );
  XNOR2_X1 U761 ( .A(n697), .B(KEYINPUT121), .ZN(n700) );
  NAND2_X1 U762 ( .A1(n698), .A2(n349), .ZN(n699) );
  NAND2_X1 U763 ( .A1(n700), .A2(n699), .ZN(n701) );
  XOR2_X1 U764 ( .A(KEYINPUT122), .B(n701), .Z(n711) );
  INV_X1 U765 ( .A(KEYINPUT79), .ZN(n705) );
  XOR2_X1 U766 ( .A(n705), .B(n350), .Z(n703) );
  NAND2_X1 U767 ( .A1(n703), .A2(n702), .ZN(n707) );
  NAND2_X1 U768 ( .A1(n705), .A2(n704), .ZN(n706) );
  NAND2_X1 U769 ( .A1(n707), .A2(n706), .ZN(n708) );
  NAND2_X1 U770 ( .A1(n709), .A2(n708), .ZN(n710) );
  NAND2_X1 U771 ( .A1(n711), .A2(n710), .ZN(n712) );
  NOR2_X1 U772 ( .A1(n712), .A2(G953), .ZN(n713) );
  XNOR2_X1 U773 ( .A(n713), .B(KEYINPUT53), .ZN(G75) );
  XOR2_X1 U774 ( .A(KEYINPUT54), .B(KEYINPUT55), .Z(n716) );
  XNOR2_X1 U775 ( .A(n714), .B(KEYINPUT84), .ZN(n715) );
  NAND2_X1 U776 ( .A1(n721), .A2(G210), .ZN(n717) );
  XNOR2_X1 U777 ( .A(n718), .B(n717), .ZN(n719) );
  NOR2_X1 U778 ( .A1(n719), .A2(n736), .ZN(n720) );
  XNOR2_X1 U779 ( .A(n720), .B(KEYINPUT56), .ZN(G51) );
  NAND2_X1 U780 ( .A1(n730), .A2(G469), .ZN(n725) );
  XOR2_X1 U781 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n723) );
  NOR2_X1 U782 ( .A1(n736), .A2(n726), .ZN(G54) );
  NAND2_X1 U783 ( .A1(G478), .A2(n730), .ZN(n727) );
  XNOR2_X1 U784 ( .A(n728), .B(n727), .ZN(n729) );
  NOR2_X1 U785 ( .A1(n736), .A2(n729), .ZN(G63) );
  NAND2_X1 U786 ( .A1(n730), .A2(G217), .ZN(n734) );
  XOR2_X1 U787 ( .A(KEYINPUT124), .B(KEYINPUT125), .Z(n731) );
  NOR2_X1 U788 ( .A1(n736), .A2(n735), .ZN(G66) );
  OR2_X1 U789 ( .A1(G953), .A2(n350), .ZN(n741) );
  NAND2_X1 U790 ( .A1(G953), .A2(G224), .ZN(n738) );
  XNOR2_X1 U791 ( .A(KEYINPUT61), .B(n738), .ZN(n739) );
  NAND2_X1 U792 ( .A1(n739), .A2(G898), .ZN(n740) );
  NAND2_X1 U793 ( .A1(n741), .A2(n740), .ZN(n748) );
  XOR2_X1 U794 ( .A(G101), .B(n742), .Z(n743) );
  XNOR2_X1 U795 ( .A(n744), .B(n743), .ZN(n746) );
  NOR2_X1 U796 ( .A1(G898), .A2(n754), .ZN(n745) );
  NOR2_X1 U797 ( .A1(n746), .A2(n745), .ZN(n747) );
  XNOR2_X1 U798 ( .A(n748), .B(n747), .ZN(n749) );
  XNOR2_X1 U799 ( .A(KEYINPUT126), .B(n749), .ZN(G69) );
  XNOR2_X1 U800 ( .A(n750), .B(n751), .ZN(n756) );
  INV_X1 U801 ( .A(n756), .ZN(n753) );
  XOR2_X1 U802 ( .A(n753), .B(n752), .Z(n755) );
  NAND2_X1 U803 ( .A1(n755), .A2(n754), .ZN(n761) );
  XOR2_X1 U804 ( .A(n756), .B(G227), .Z(n757) );
  XNOR2_X1 U805 ( .A(n757), .B(KEYINPUT127), .ZN(n758) );
  NAND2_X1 U806 ( .A1(n758), .A2(G900), .ZN(n759) );
  NAND2_X1 U807 ( .A1(n759), .A2(G953), .ZN(n760) );
  NAND2_X1 U808 ( .A1(n761), .A2(n760), .ZN(G72) );
  XNOR2_X1 U809 ( .A(n762), .B(G122), .ZN(G24) );
  XOR2_X1 U810 ( .A(n763), .B(G119), .Z(G21) );
  XNOR2_X1 U811 ( .A(G140), .B(n764), .ZN(G42) );
  XNOR2_X1 U812 ( .A(n765), .B(G137), .ZN(G39) );
  XNOR2_X1 U813 ( .A(G131), .B(n766), .ZN(G33) );
endmodule

