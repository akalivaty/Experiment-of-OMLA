//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 1 0 1 0 1 0 0 0 1 0 0 1 1 1 1 1 0 0 1 1 0 1 0 1 0 0 1 0 1 0 1 1 1 0 0 0 1 1 1 1 1 0 0 0 0 0 0 0 1 1 0 1 0 0 0 0 1 0 0 1 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:33:39 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n442, new_n444, new_n448, new_n452, new_n453, new_n454, new_n455,
    new_n458, new_n459, new_n460, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n527, new_n528, new_n529, new_n530, new_n531, new_n532,
    new_n533, new_n534, new_n535, new_n536, new_n537, new_n538, new_n539,
    new_n540, new_n541, new_n542, new_n543, new_n544, new_n545, new_n546,
    new_n547, new_n550, new_n551, new_n552, new_n553, new_n554, new_n556,
    new_n557, new_n558, new_n559, new_n560, new_n561, new_n564, new_n565,
    new_n566, new_n568, new_n569, new_n570, new_n571, new_n572, new_n573,
    new_n574, new_n575, new_n579, new_n580, new_n582, new_n583, new_n584,
    new_n585, new_n586, new_n587, new_n588, new_n589, new_n590, new_n591,
    new_n592, new_n593, new_n594, new_n595, new_n596, new_n597, new_n599,
    new_n600, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n624, new_n625, new_n628, new_n630, new_n631, new_n632, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1197, new_n1198, new_n1199, new_n1200, new_n1201, new_n1202;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  XNOR2_X1  g008(.A(KEYINPUT64), .B(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  XNOR2_X1  g011(.A(KEYINPUT65), .B(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  AND2_X1   g016(.A1(G2072), .A2(G2078), .ZN(new_n442));
  NAND3_X1  g017(.A1(new_n442), .A2(G2084), .A3(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(new_n444));
  XNOR2_X1  g019(.A(new_n444), .B(KEYINPUT66), .ZN(G259));
  BUF_X1    g020(.A(G452), .Z(G391));
  AND2_X1   g021(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g022(.A1(G7), .A2(G661), .ZN(new_n448));
  XOR2_X1   g023(.A(new_n448), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g024(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g025(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g026(.A1(G218), .A2(G220), .A3(G221), .A4(G219), .ZN(new_n452));
  XNOR2_X1  g027(.A(KEYINPUT67), .B(KEYINPUT2), .ZN(new_n453));
  XNOR2_X1  g028(.A(new_n452), .B(new_n453), .ZN(new_n454));
  NAND4_X1  g029(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n455));
  NOR2_X1   g030(.A1(new_n454), .A2(new_n455), .ZN(G325));
  INV_X1    g031(.A(G325), .ZN(G261));
  NAND2_X1  g032(.A1(new_n454), .A2(G2106), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n455), .A2(G567), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  INV_X1    g035(.A(new_n460), .ZN(G319));
  INV_X1    g036(.A(G2105), .ZN(new_n462));
  INV_X1    g037(.A(KEYINPUT68), .ZN(new_n463));
  AND2_X1   g038(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n464));
  NOR2_X1   g039(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n465));
  OAI21_X1  g040(.A(new_n463), .B1(new_n464), .B2(new_n465), .ZN(new_n466));
  INV_X1    g041(.A(KEYINPUT3), .ZN(new_n467));
  INV_X1    g042(.A(G2104), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  NAND2_X1  g044(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n470));
  NAND3_X1  g045(.A1(new_n469), .A2(KEYINPUT68), .A3(new_n470), .ZN(new_n471));
  NAND3_X1  g046(.A1(new_n466), .A2(new_n471), .A3(G125), .ZN(new_n472));
  NAND2_X1  g047(.A1(G113), .A2(G2104), .ZN(new_n473));
  AOI21_X1  g048(.A(new_n462), .B1(new_n472), .B2(new_n473), .ZN(new_n474));
  NOR2_X1   g049(.A1(new_n468), .A2(G2105), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n475), .A2(G101), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n469), .A2(new_n470), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n477), .A2(new_n462), .ZN(new_n478));
  INV_X1    g053(.A(G137), .ZN(new_n479));
  OAI21_X1  g054(.A(new_n476), .B1(new_n478), .B2(new_n479), .ZN(new_n480));
  NOR2_X1   g055(.A1(new_n474), .A2(new_n480), .ZN(G160));
  NAND2_X1  g056(.A1(new_n477), .A2(G2105), .ZN(new_n482));
  INV_X1    g057(.A(new_n482), .ZN(new_n483));
  NAND2_X1  g058(.A1(new_n483), .A2(G124), .ZN(new_n484));
  NOR2_X1   g059(.A1(new_n462), .A2(G112), .ZN(new_n485));
  OAI21_X1  g060(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n486));
  OAI21_X1  g061(.A(new_n484), .B1(new_n485), .B2(new_n486), .ZN(new_n487));
  NOR2_X1   g062(.A1(new_n464), .A2(new_n465), .ZN(new_n488));
  NOR2_X1   g063(.A1(new_n488), .A2(G2105), .ZN(new_n489));
  AOI21_X1  g064(.A(new_n487), .B1(G136), .B2(new_n489), .ZN(new_n490));
  XOR2_X1   g065(.A(new_n490), .B(KEYINPUT69), .Z(G162));
  OR2_X1    g066(.A1(G102), .A2(G2105), .ZN(new_n492));
  INV_X1    g067(.A(KEYINPUT70), .ZN(new_n493));
  INV_X1    g068(.A(G114), .ZN(new_n494));
  AOI21_X1  g069(.A(new_n493), .B1(new_n494), .B2(G2105), .ZN(new_n495));
  NOR3_X1   g070(.A1(new_n462), .A2(KEYINPUT70), .A3(G114), .ZN(new_n496));
  OAI211_X1 g071(.A(G2104), .B(new_n492), .C1(new_n495), .C2(new_n496), .ZN(new_n497));
  NAND3_X1  g072(.A1(new_n477), .A2(G126), .A3(G2105), .ZN(new_n498));
  NAND2_X1  g073(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  INV_X1    g074(.A(G138), .ZN(new_n500));
  NOR3_X1   g075(.A1(new_n500), .A2(KEYINPUT4), .A3(G2105), .ZN(new_n501));
  NAND3_X1  g076(.A1(new_n466), .A2(new_n471), .A3(new_n501), .ZN(new_n502));
  OAI211_X1 g077(.A(G138), .B(new_n462), .C1(new_n464), .C2(new_n465), .ZN(new_n503));
  AOI22_X1  g078(.A1(new_n502), .A2(KEYINPUT71), .B1(KEYINPUT4), .B2(new_n503), .ZN(new_n504));
  INV_X1    g079(.A(KEYINPUT71), .ZN(new_n505));
  NAND4_X1  g080(.A1(new_n466), .A2(new_n471), .A3(new_n505), .A4(new_n501), .ZN(new_n506));
  AOI21_X1  g081(.A(new_n499), .B1(new_n504), .B2(new_n506), .ZN(G164));
  INV_X1    g082(.A(G543), .ZN(new_n508));
  INV_X1    g083(.A(KEYINPUT5), .ZN(new_n509));
  OAI21_X1  g084(.A(new_n508), .B1(new_n509), .B2(KEYINPUT72), .ZN(new_n510));
  INV_X1    g085(.A(KEYINPUT72), .ZN(new_n511));
  NAND3_X1  g086(.A1(new_n511), .A2(KEYINPUT5), .A3(G543), .ZN(new_n512));
  NAND2_X1  g087(.A1(new_n510), .A2(new_n512), .ZN(new_n513));
  AOI22_X1  g088(.A1(new_n513), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n514));
  INV_X1    g089(.A(G651), .ZN(new_n515));
  NOR2_X1   g090(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  INV_X1    g091(.A(KEYINPUT6), .ZN(new_n517));
  NAND2_X1  g092(.A1(new_n517), .A2(new_n515), .ZN(new_n518));
  NAND2_X1  g093(.A1(KEYINPUT6), .A2(G651), .ZN(new_n519));
  AOI21_X1  g094(.A(new_n508), .B1(new_n518), .B2(new_n519), .ZN(new_n520));
  NAND2_X1  g095(.A1(new_n520), .A2(G50), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n518), .A2(new_n519), .ZN(new_n522));
  NAND2_X1  g097(.A1(new_n513), .A2(new_n522), .ZN(new_n523));
  INV_X1    g098(.A(G88), .ZN(new_n524));
  OAI21_X1  g099(.A(new_n521), .B1(new_n523), .B2(new_n524), .ZN(new_n525));
  NOR2_X1   g100(.A1(new_n516), .A2(new_n525), .ZN(G166));
  AND2_X1   g101(.A1(G63), .A2(G651), .ZN(new_n527));
  NAND2_X1  g102(.A1(new_n513), .A2(new_n527), .ZN(new_n528));
  INV_X1    g103(.A(new_n519), .ZN(new_n529));
  NOR2_X1   g104(.A1(KEYINPUT6), .A2(G651), .ZN(new_n530));
  OAI211_X1 g105(.A(G51), .B(G543), .C1(new_n529), .C2(new_n530), .ZN(new_n531));
  NAND2_X1  g106(.A1(new_n528), .A2(new_n531), .ZN(new_n532));
  INV_X1    g107(.A(KEYINPUT73), .ZN(new_n533));
  NAND2_X1  g108(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  NAND3_X1  g109(.A1(new_n528), .A2(KEYINPUT73), .A3(new_n531), .ZN(new_n535));
  AOI22_X1  g110(.A1(new_n510), .A2(new_n512), .B1(new_n518), .B2(new_n519), .ZN(new_n536));
  XOR2_X1   g111(.A(KEYINPUT75), .B(G89), .Z(new_n537));
  NAND2_X1  g112(.A1(new_n536), .A2(new_n537), .ZN(new_n538));
  NAND3_X1  g113(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n539));
  NAND2_X1  g114(.A1(new_n539), .A2(KEYINPUT74), .ZN(new_n540));
  INV_X1    g115(.A(KEYINPUT74), .ZN(new_n541));
  NAND4_X1  g116(.A1(new_n541), .A2(G76), .A3(G543), .A4(G651), .ZN(new_n542));
  NAND2_X1  g117(.A1(new_n540), .A2(new_n542), .ZN(new_n543));
  NAND2_X1  g118(.A1(new_n543), .A2(KEYINPUT7), .ZN(new_n544));
  INV_X1    g119(.A(KEYINPUT7), .ZN(new_n545));
  NAND3_X1  g120(.A1(new_n540), .A2(new_n545), .A3(new_n542), .ZN(new_n546));
  NAND2_X1  g121(.A1(new_n544), .A2(new_n546), .ZN(new_n547));
  NAND4_X1  g122(.A1(new_n534), .A2(new_n535), .A3(new_n538), .A4(new_n547), .ZN(G286));
  INV_X1    g123(.A(G286), .ZN(G168));
  AOI22_X1  g124(.A1(new_n513), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n550));
  NOR2_X1   g125(.A1(new_n550), .A2(new_n515), .ZN(new_n551));
  NAND2_X1  g126(.A1(new_n520), .A2(G52), .ZN(new_n552));
  INV_X1    g127(.A(G90), .ZN(new_n553));
  OAI21_X1  g128(.A(new_n552), .B1(new_n523), .B2(new_n553), .ZN(new_n554));
  NOR2_X1   g129(.A1(new_n551), .A2(new_n554), .ZN(G171));
  XOR2_X1   g130(.A(KEYINPUT76), .B(G43), .Z(new_n556));
  AOI22_X1  g131(.A1(new_n536), .A2(G81), .B1(new_n520), .B2(new_n556), .ZN(new_n557));
  INV_X1    g132(.A(new_n557), .ZN(new_n558));
  AOI22_X1  g133(.A1(new_n513), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n559));
  NOR2_X1   g134(.A1(new_n559), .A2(new_n515), .ZN(new_n560));
  NOR2_X1   g135(.A1(new_n558), .A2(new_n560), .ZN(new_n561));
  NAND2_X1  g136(.A1(new_n561), .A2(G860), .ZN(G153));
  NAND4_X1  g137(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g138(.A1(G1), .A2(G3), .ZN(new_n564));
  XNOR2_X1  g139(.A(new_n564), .B(KEYINPUT8), .ZN(new_n565));
  NAND4_X1  g140(.A1(G319), .A2(G483), .A3(G661), .A4(new_n565), .ZN(new_n566));
  XNOR2_X1  g141(.A(new_n566), .B(KEYINPUT77), .ZN(G188));
  NAND2_X1  g142(.A1(new_n520), .A2(G53), .ZN(new_n568));
  XNOR2_X1  g143(.A(new_n568), .B(KEYINPUT9), .ZN(new_n569));
  XNOR2_X1  g144(.A(KEYINPUT79), .B(G65), .ZN(new_n570));
  AND2_X1   g145(.A1(new_n513), .A2(new_n570), .ZN(new_n571));
  NAND2_X1  g146(.A1(G78), .A2(G543), .ZN(new_n572));
  XOR2_X1   g147(.A(new_n572), .B(KEYINPUT78), .Z(new_n573));
  OAI21_X1  g148(.A(G651), .B1(new_n571), .B2(new_n573), .ZN(new_n574));
  NAND2_X1  g149(.A1(new_n536), .A2(G91), .ZN(new_n575));
  NAND3_X1  g150(.A1(new_n569), .A2(new_n574), .A3(new_n575), .ZN(G299));
  OAI221_X1 g151(.A(new_n552), .B1(new_n523), .B2(new_n553), .C1(new_n550), .C2(new_n515), .ZN(G301));
  INV_X1    g152(.A(G166), .ZN(G303));
  AOI22_X1  g153(.A1(new_n536), .A2(G87), .B1(new_n520), .B2(G49), .ZN(new_n579));
  OAI21_X1  g154(.A(G651), .B1(new_n513), .B2(G74), .ZN(new_n580));
  NAND2_X1  g155(.A1(new_n579), .A2(new_n580), .ZN(G288));
  INV_X1    g156(.A(G61), .ZN(new_n582));
  AOI21_X1  g157(.A(new_n582), .B1(new_n510), .B2(new_n512), .ZN(new_n583));
  INV_X1    g158(.A(KEYINPUT80), .ZN(new_n584));
  INV_X1    g159(.A(G73), .ZN(new_n585));
  OAI21_X1  g160(.A(new_n584), .B1(new_n585), .B2(new_n508), .ZN(new_n586));
  NAND3_X1  g161(.A1(KEYINPUT80), .A2(G73), .A3(G543), .ZN(new_n587));
  NAND2_X1  g162(.A1(new_n586), .A2(new_n587), .ZN(new_n588));
  OAI21_X1  g163(.A(G651), .B1(new_n583), .B2(new_n588), .ZN(new_n589));
  NAND2_X1  g164(.A1(new_n589), .A2(KEYINPUT81), .ZN(new_n590));
  INV_X1    g165(.A(KEYINPUT81), .ZN(new_n591));
  OAI211_X1 g166(.A(new_n591), .B(G651), .C1(new_n583), .C2(new_n588), .ZN(new_n592));
  NAND2_X1  g167(.A1(new_n590), .A2(new_n592), .ZN(new_n593));
  NAND3_X1  g168(.A1(new_n513), .A2(G86), .A3(new_n522), .ZN(new_n594));
  NAND2_X1  g169(.A1(new_n520), .A2(G48), .ZN(new_n595));
  NAND2_X1  g170(.A1(new_n594), .A2(new_n595), .ZN(new_n596));
  INV_X1    g171(.A(new_n596), .ZN(new_n597));
  NAND2_X1  g172(.A1(new_n593), .A2(new_n597), .ZN(G305));
  AOI22_X1  g173(.A1(new_n536), .A2(G85), .B1(new_n520), .B2(G47), .ZN(new_n599));
  AOI22_X1  g174(.A1(new_n513), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n600));
  OAI21_X1  g175(.A(new_n599), .B1(new_n515), .B2(new_n600), .ZN(G290));
  NAND2_X1  g176(.A1(G301), .A2(G868), .ZN(new_n602));
  INV_X1    g177(.A(KEYINPUT82), .ZN(new_n603));
  AOI21_X1  g178(.A(new_n603), .B1(new_n536), .B2(G92), .ZN(new_n604));
  INV_X1    g179(.A(new_n604), .ZN(new_n605));
  NAND3_X1  g180(.A1(new_n536), .A2(new_n603), .A3(G92), .ZN(new_n606));
  NAND3_X1  g181(.A1(new_n605), .A2(KEYINPUT10), .A3(new_n606), .ZN(new_n607));
  INV_X1    g182(.A(KEYINPUT10), .ZN(new_n608));
  INV_X1    g183(.A(new_n606), .ZN(new_n609));
  OAI21_X1  g184(.A(new_n608), .B1(new_n609), .B2(new_n604), .ZN(new_n610));
  INV_X1    g185(.A(G66), .ZN(new_n611));
  AOI21_X1  g186(.A(new_n611), .B1(new_n510), .B2(new_n512), .ZN(new_n612));
  AND2_X1   g187(.A1(G79), .A2(G543), .ZN(new_n613));
  OAI21_X1  g188(.A(G651), .B1(new_n612), .B2(new_n613), .ZN(new_n614));
  NAND2_X1  g189(.A1(new_n520), .A2(G54), .ZN(new_n615));
  NAND2_X1  g190(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  NOR2_X1   g191(.A1(new_n616), .A2(KEYINPUT83), .ZN(new_n617));
  INV_X1    g192(.A(KEYINPUT83), .ZN(new_n618));
  AOI21_X1  g193(.A(new_n618), .B1(new_n614), .B2(new_n615), .ZN(new_n619));
  OAI211_X1 g194(.A(new_n607), .B(new_n610), .C1(new_n617), .C2(new_n619), .ZN(new_n620));
  INV_X1    g195(.A(new_n620), .ZN(new_n621));
  OAI21_X1  g196(.A(new_n602), .B1(new_n621), .B2(G868), .ZN(G321));
  XNOR2_X1  g197(.A(G321), .B(KEYINPUT84), .ZN(G284));
  NAND2_X1  g198(.A1(G286), .A2(G868), .ZN(new_n624));
  AND3_X1   g199(.A1(new_n569), .A2(new_n574), .A3(new_n575), .ZN(new_n625));
  OAI21_X1  g200(.A(new_n624), .B1(new_n625), .B2(G868), .ZN(G297));
  OAI21_X1  g201(.A(new_n624), .B1(new_n625), .B2(G868), .ZN(G280));
  INV_X1    g202(.A(G559), .ZN(new_n628));
  OAI21_X1  g203(.A(new_n621), .B1(new_n628), .B2(G860), .ZN(G148));
  NOR2_X1   g204(.A1(new_n620), .A2(G559), .ZN(new_n630));
  INV_X1    g205(.A(new_n630), .ZN(new_n631));
  NAND2_X1  g206(.A1(new_n631), .A2(G868), .ZN(new_n632));
  OAI21_X1  g207(.A(new_n632), .B1(G868), .B2(new_n561), .ZN(G323));
  XNOR2_X1  g208(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g209(.A1(new_n483), .A2(G123), .ZN(new_n635));
  NAND2_X1  g210(.A1(new_n489), .A2(G135), .ZN(new_n636));
  NOR2_X1   g211(.A1(new_n462), .A2(G111), .ZN(new_n637));
  OAI21_X1  g212(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n638));
  OAI211_X1 g213(.A(new_n635), .B(new_n636), .C1(new_n637), .C2(new_n638), .ZN(new_n639));
  XNOR2_X1  g214(.A(new_n639), .B(KEYINPUT85), .ZN(new_n640));
  XOR2_X1   g215(.A(new_n640), .B(G2096), .Z(new_n641));
  AND2_X1   g216(.A1(new_n466), .A2(new_n471), .ZN(new_n642));
  NAND2_X1  g217(.A1(new_n642), .A2(new_n475), .ZN(new_n643));
  XNOR2_X1  g218(.A(new_n643), .B(KEYINPUT12), .ZN(new_n644));
  XNOR2_X1  g219(.A(new_n644), .B(KEYINPUT13), .ZN(new_n645));
  INV_X1    g220(.A(G2100), .ZN(new_n646));
  OR2_X1    g221(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  NAND2_X1  g222(.A1(new_n645), .A2(new_n646), .ZN(new_n648));
  NAND3_X1  g223(.A1(new_n641), .A2(new_n647), .A3(new_n648), .ZN(G156));
  XOR2_X1   g224(.A(G2451), .B(G2454), .Z(new_n650));
  XNOR2_X1  g225(.A(new_n650), .B(KEYINPUT16), .ZN(new_n651));
  XNOR2_X1  g226(.A(G1341), .B(G1348), .ZN(new_n652));
  XNOR2_X1  g227(.A(new_n652), .B(KEYINPUT87), .ZN(new_n653));
  XOR2_X1   g228(.A(new_n651), .B(new_n653), .Z(new_n654));
  INV_X1    g229(.A(KEYINPUT14), .ZN(new_n655));
  XNOR2_X1  g230(.A(KEYINPUT15), .B(G2435), .ZN(new_n656));
  XNOR2_X1  g231(.A(KEYINPUT86), .B(G2438), .ZN(new_n657));
  XNOR2_X1  g232(.A(new_n656), .B(new_n657), .ZN(new_n658));
  XOR2_X1   g233(.A(G2427), .B(G2430), .Z(new_n659));
  AOI21_X1  g234(.A(new_n655), .B1(new_n658), .B2(new_n659), .ZN(new_n660));
  OAI21_X1  g235(.A(new_n660), .B1(new_n659), .B2(new_n658), .ZN(new_n661));
  XNOR2_X1  g236(.A(new_n654), .B(new_n661), .ZN(new_n662));
  INV_X1    g237(.A(new_n662), .ZN(new_n663));
  XNOR2_X1  g238(.A(G2443), .B(G2446), .ZN(new_n664));
  INV_X1    g239(.A(new_n664), .ZN(new_n665));
  OAI21_X1  g240(.A(G14), .B1(new_n663), .B2(new_n665), .ZN(new_n666));
  AOI21_X1  g241(.A(new_n666), .B1(new_n665), .B2(new_n663), .ZN(G401));
  XNOR2_X1  g242(.A(G2067), .B(G2678), .ZN(new_n668));
  XNOR2_X1  g243(.A(G2072), .B(G2078), .ZN(new_n669));
  INV_X1    g244(.A(KEYINPUT88), .ZN(new_n670));
  AOI21_X1  g245(.A(new_n668), .B1(new_n669), .B2(new_n670), .ZN(new_n671));
  OAI21_X1  g246(.A(new_n671), .B1(new_n670), .B2(new_n669), .ZN(new_n672));
  XOR2_X1   g247(.A(G2084), .B(G2090), .Z(new_n673));
  INV_X1    g248(.A(new_n673), .ZN(new_n674));
  XOR2_X1   g249(.A(new_n669), .B(KEYINPUT17), .Z(new_n675));
  INV_X1    g250(.A(new_n668), .ZN(new_n676));
  OAI211_X1 g251(.A(new_n672), .B(new_n674), .C1(new_n675), .C2(new_n676), .ZN(new_n677));
  XNOR2_X1  g252(.A(new_n677), .B(KEYINPUT89), .ZN(new_n678));
  NAND3_X1  g253(.A1(new_n673), .A2(new_n669), .A3(new_n668), .ZN(new_n679));
  XOR2_X1   g254(.A(new_n679), .B(KEYINPUT18), .Z(new_n680));
  NAND3_X1  g255(.A1(new_n675), .A2(new_n676), .A3(new_n673), .ZN(new_n681));
  NAND3_X1  g256(.A1(new_n678), .A2(new_n680), .A3(new_n681), .ZN(new_n682));
  XNOR2_X1  g257(.A(new_n682), .B(new_n646), .ZN(new_n683));
  XNOR2_X1  g258(.A(KEYINPUT90), .B(G2096), .ZN(new_n684));
  XNOR2_X1  g259(.A(new_n683), .B(new_n684), .ZN(new_n685));
  INV_X1    g260(.A(new_n685), .ZN(G227));
  XNOR2_X1  g261(.A(G1971), .B(G1976), .ZN(new_n687));
  INV_X1    g262(.A(KEYINPUT19), .ZN(new_n688));
  XNOR2_X1  g263(.A(new_n687), .B(new_n688), .ZN(new_n689));
  XOR2_X1   g264(.A(G1956), .B(G2474), .Z(new_n690));
  XOR2_X1   g265(.A(G1961), .B(G1966), .Z(new_n691));
  AND2_X1   g266(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  NAND2_X1  g267(.A1(new_n689), .A2(new_n692), .ZN(new_n693));
  XNOR2_X1  g268(.A(new_n693), .B(KEYINPUT20), .ZN(new_n694));
  NOR2_X1   g269(.A1(new_n690), .A2(new_n691), .ZN(new_n695));
  NOR3_X1   g270(.A1(new_n689), .A2(new_n692), .A3(new_n695), .ZN(new_n696));
  AOI21_X1  g271(.A(new_n696), .B1(new_n689), .B2(new_n695), .ZN(new_n697));
  AND2_X1   g272(.A1(new_n694), .A2(new_n697), .ZN(new_n698));
  XNOR2_X1  g273(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n699));
  XNOR2_X1  g274(.A(new_n698), .B(new_n699), .ZN(new_n700));
  XNOR2_X1  g275(.A(G1991), .B(G1996), .ZN(new_n701));
  XNOR2_X1  g276(.A(new_n700), .B(new_n701), .ZN(new_n702));
  XNOR2_X1  g277(.A(G1981), .B(G1986), .ZN(new_n703));
  XNOR2_X1  g278(.A(new_n702), .B(new_n703), .ZN(new_n704));
  INV_X1    g279(.A(new_n704), .ZN(G229));
  XNOR2_X1  g280(.A(KEYINPUT31), .B(G11), .ZN(new_n706));
  XOR2_X1   g281(.A(new_n706), .B(KEYINPUT101), .Z(new_n707));
  INV_X1    g282(.A(G28), .ZN(new_n708));
  NOR2_X1   g283(.A1(new_n708), .A2(KEYINPUT30), .ZN(new_n709));
  INV_X1    g284(.A(G29), .ZN(new_n710));
  INV_X1    g285(.A(KEYINPUT30), .ZN(new_n711));
  OAI21_X1  g286(.A(new_n710), .B1(new_n711), .B2(G28), .ZN(new_n712));
  OR2_X1    g287(.A1(new_n710), .A2(KEYINPUT91), .ZN(new_n713));
  NAND2_X1  g288(.A1(new_n710), .A2(KEYINPUT91), .ZN(new_n714));
  NAND2_X1  g289(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  INV_X1    g290(.A(new_n715), .ZN(new_n716));
  OAI221_X1 g291(.A(new_n707), .B1(new_n709), .B2(new_n712), .C1(new_n640), .C2(new_n716), .ZN(new_n717));
  NAND2_X1  g292(.A1(new_n710), .A2(G32), .ZN(new_n718));
  NAND3_X1  g293(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n719));
  XOR2_X1   g294(.A(new_n719), .B(KEYINPUT26), .Z(new_n720));
  INV_X1    g295(.A(G129), .ZN(new_n721));
  OAI21_X1  g296(.A(new_n720), .B1(new_n482), .B2(new_n721), .ZN(new_n722));
  NAND2_X1  g297(.A1(new_n475), .A2(G105), .ZN(new_n723));
  INV_X1    g298(.A(G141), .ZN(new_n724));
  OAI21_X1  g299(.A(new_n723), .B1(new_n478), .B2(new_n724), .ZN(new_n725));
  OR2_X1    g300(.A1(new_n722), .A2(new_n725), .ZN(new_n726));
  INV_X1    g301(.A(new_n726), .ZN(new_n727));
  OAI21_X1  g302(.A(new_n718), .B1(new_n727), .B2(new_n710), .ZN(new_n728));
  XNOR2_X1  g303(.A(new_n728), .B(KEYINPUT100), .ZN(new_n729));
  XNOR2_X1  g304(.A(KEYINPUT27), .B(G1996), .ZN(new_n730));
  NOR2_X1   g305(.A1(new_n729), .A2(new_n730), .ZN(new_n731));
  INV_X1    g306(.A(G16), .ZN(new_n732));
  NAND2_X1  g307(.A1(new_n732), .A2(G5), .ZN(new_n733));
  OAI21_X1  g308(.A(new_n733), .B1(G171), .B2(new_n732), .ZN(new_n734));
  AOI211_X1 g309(.A(new_n717), .B(new_n731), .C1(G1961), .C2(new_n734), .ZN(new_n735));
  INV_X1    g310(.A(KEYINPUT24), .ZN(new_n736));
  NAND2_X1  g311(.A1(new_n736), .A2(G34), .ZN(new_n737));
  OAI21_X1  g312(.A(new_n716), .B1(new_n736), .B2(G34), .ZN(new_n738));
  INV_X1    g313(.A(KEYINPUT99), .ZN(new_n739));
  OAI21_X1  g314(.A(new_n737), .B1(new_n738), .B2(new_n739), .ZN(new_n740));
  AOI21_X1  g315(.A(new_n740), .B1(new_n739), .B2(new_n738), .ZN(new_n741));
  AOI21_X1  g316(.A(new_n741), .B1(G160), .B2(G29), .ZN(new_n742));
  AOI22_X1  g317(.A1(new_n729), .A2(new_n730), .B1(G2084), .B2(new_n742), .ZN(new_n743));
  NAND2_X1  g318(.A1(new_n732), .A2(G21), .ZN(new_n744));
  OAI21_X1  g319(.A(new_n744), .B1(G168), .B2(new_n732), .ZN(new_n745));
  INV_X1    g320(.A(G1966), .ZN(new_n746));
  XNOR2_X1  g321(.A(new_n745), .B(new_n746), .ZN(new_n747));
  XOR2_X1   g322(.A(KEYINPUT92), .B(G16), .Z(new_n748));
  INV_X1    g323(.A(new_n748), .ZN(new_n749));
  NAND2_X1  g324(.A1(new_n561), .A2(new_n749), .ZN(new_n750));
  OAI21_X1  g325(.A(new_n750), .B1(G19), .B2(new_n749), .ZN(new_n751));
  INV_X1    g326(.A(G1341), .ZN(new_n752));
  OAI22_X1  g327(.A1(new_n751), .A2(new_n752), .B1(new_n734), .B2(G1961), .ZN(new_n753));
  NAND2_X1  g328(.A1(new_n716), .A2(G26), .ZN(new_n754));
  XNOR2_X1  g329(.A(new_n754), .B(KEYINPUT28), .ZN(new_n755));
  AOI22_X1  g330(.A1(new_n483), .A2(G128), .B1(new_n489), .B2(G140), .ZN(new_n756));
  NOR2_X1   g331(.A1(G104), .A2(G2105), .ZN(new_n757));
  INV_X1    g332(.A(KEYINPUT95), .ZN(new_n758));
  XNOR2_X1  g333(.A(new_n757), .B(new_n758), .ZN(new_n759));
  OAI21_X1  g334(.A(G2104), .B1(new_n462), .B2(G116), .ZN(new_n760));
  OR2_X1    g335(.A1(new_n759), .A2(new_n760), .ZN(new_n761));
  AND2_X1   g336(.A1(new_n756), .A2(new_n761), .ZN(new_n762));
  OAI21_X1  g337(.A(new_n755), .B1(new_n762), .B2(new_n710), .ZN(new_n763));
  XNOR2_X1  g338(.A(new_n763), .B(G2067), .ZN(new_n764));
  AOI211_X1 g339(.A(new_n753), .B(new_n764), .C1(new_n752), .C2(new_n751), .ZN(new_n765));
  NAND4_X1  g340(.A1(new_n735), .A2(new_n743), .A3(new_n747), .A4(new_n765), .ZN(new_n766));
  NAND2_X1  g341(.A1(new_n642), .A2(G127), .ZN(new_n767));
  NAND2_X1  g342(.A1(G115), .A2(G2104), .ZN(new_n768));
  AOI21_X1  g343(.A(new_n462), .B1(new_n767), .B2(new_n768), .ZN(new_n769));
  XNOR2_X1  g344(.A(KEYINPUT96), .B(KEYINPUT25), .ZN(new_n770));
  AND3_X1   g345(.A1(new_n462), .A2(G103), .A3(G2104), .ZN(new_n771));
  XNOR2_X1  g346(.A(new_n770), .B(new_n771), .ZN(new_n772));
  INV_X1    g347(.A(G139), .ZN(new_n773));
  OAI21_X1  g348(.A(new_n772), .B1(new_n773), .B2(new_n478), .ZN(new_n774));
  OR3_X1    g349(.A1(new_n769), .A2(KEYINPUT97), .A3(new_n774), .ZN(new_n775));
  OAI21_X1  g350(.A(KEYINPUT97), .B1(new_n769), .B2(new_n774), .ZN(new_n776));
  NAND2_X1  g351(.A1(new_n775), .A2(new_n776), .ZN(new_n777));
  MUX2_X1   g352(.A(G33), .B(new_n777), .S(G29), .Z(new_n778));
  XNOR2_X1  g353(.A(KEYINPUT98), .B(G2072), .ZN(new_n779));
  XNOR2_X1  g354(.A(new_n778), .B(new_n779), .ZN(new_n780));
  NAND2_X1  g355(.A1(new_n748), .A2(G20), .ZN(new_n781));
  XOR2_X1   g356(.A(new_n781), .B(KEYINPUT23), .Z(new_n782));
  AOI21_X1  g357(.A(new_n782), .B1(G299), .B2(G16), .ZN(new_n783));
  XNOR2_X1  g358(.A(new_n783), .B(G1956), .ZN(new_n784));
  NOR2_X1   g359(.A1(new_n742), .A2(G2084), .ZN(new_n785));
  OAI21_X1  g360(.A(new_n784), .B1(KEYINPUT102), .B2(new_n785), .ZN(new_n786));
  NOR2_X1   g361(.A1(new_n715), .A2(G35), .ZN(new_n787));
  AOI21_X1  g362(.A(new_n787), .B1(G162), .B2(new_n715), .ZN(new_n788));
  XNOR2_X1  g363(.A(KEYINPUT104), .B(KEYINPUT29), .ZN(new_n789));
  INV_X1    g364(.A(G2090), .ZN(new_n790));
  XNOR2_X1  g365(.A(new_n789), .B(new_n790), .ZN(new_n791));
  XNOR2_X1  g366(.A(new_n788), .B(new_n791), .ZN(new_n792));
  NAND2_X1  g367(.A1(new_n785), .A2(KEYINPUT102), .ZN(new_n793));
  NAND2_X1  g368(.A1(new_n792), .A2(new_n793), .ZN(new_n794));
  NOR4_X1   g369(.A1(new_n766), .A2(new_n780), .A3(new_n786), .A4(new_n794), .ZN(new_n795));
  NAND2_X1  g370(.A1(new_n732), .A2(G6), .ZN(new_n796));
  INV_X1    g371(.A(G305), .ZN(new_n797));
  OAI21_X1  g372(.A(new_n796), .B1(new_n797), .B2(new_n732), .ZN(new_n798));
  XNOR2_X1  g373(.A(KEYINPUT32), .B(G1981), .ZN(new_n799));
  OR2_X1    g374(.A1(new_n798), .A2(new_n799), .ZN(new_n800));
  NAND2_X1  g375(.A1(new_n798), .A2(new_n799), .ZN(new_n801));
  NOR2_X1   g376(.A1(new_n749), .A2(G22), .ZN(new_n802));
  AOI21_X1  g377(.A(new_n802), .B1(G166), .B2(new_n749), .ZN(new_n803));
  INV_X1    g378(.A(G1971), .ZN(new_n804));
  XNOR2_X1  g379(.A(new_n803), .B(new_n804), .ZN(new_n805));
  NAND2_X1  g380(.A1(new_n732), .A2(G23), .ZN(new_n806));
  INV_X1    g381(.A(G288), .ZN(new_n807));
  OAI21_X1  g382(.A(new_n806), .B1(new_n807), .B2(new_n732), .ZN(new_n808));
  XNOR2_X1  g383(.A(KEYINPUT33), .B(G1976), .ZN(new_n809));
  XNOR2_X1  g384(.A(new_n808), .B(new_n809), .ZN(new_n810));
  NAND4_X1  g385(.A1(new_n800), .A2(new_n801), .A3(new_n805), .A4(new_n810), .ZN(new_n811));
  OR2_X1    g386(.A1(new_n811), .A2(KEYINPUT34), .ZN(new_n812));
  NAND2_X1  g387(.A1(new_n811), .A2(KEYINPUT34), .ZN(new_n813));
  NAND2_X1  g388(.A1(new_n748), .A2(G24), .ZN(new_n814));
  XNOR2_X1  g389(.A(new_n814), .B(KEYINPUT93), .ZN(new_n815));
  AOI21_X1  g390(.A(new_n815), .B1(G290), .B2(new_n749), .ZN(new_n816));
  XOR2_X1   g391(.A(new_n816), .B(G1986), .Z(new_n817));
  OR2_X1    g392(.A1(G95), .A2(G2105), .ZN(new_n818));
  OAI211_X1 g393(.A(new_n818), .B(G2104), .C1(G107), .C2(new_n462), .ZN(new_n819));
  INV_X1    g394(.A(G131), .ZN(new_n820));
  INV_X1    g395(.A(G119), .ZN(new_n821));
  OAI221_X1 g396(.A(new_n819), .B1(new_n478), .B2(new_n820), .C1(new_n821), .C2(new_n482), .ZN(new_n822));
  MUX2_X1   g397(.A(G25), .B(new_n822), .S(new_n715), .Z(new_n823));
  XNOR2_X1  g398(.A(KEYINPUT35), .B(G1991), .ZN(new_n824));
  XNOR2_X1  g399(.A(new_n823), .B(new_n824), .ZN(new_n825));
  NOR2_X1   g400(.A1(new_n817), .A2(new_n825), .ZN(new_n826));
  NAND3_X1  g401(.A1(new_n812), .A2(new_n813), .A3(new_n826), .ZN(new_n827));
  INV_X1    g402(.A(new_n827), .ZN(new_n828));
  NAND3_X1  g403(.A1(new_n828), .A2(KEYINPUT94), .A3(KEYINPUT36), .ZN(new_n829));
  XOR2_X1   g404(.A(KEYINPUT94), .B(KEYINPUT36), .Z(new_n830));
  NAND2_X1  g405(.A1(new_n827), .A2(new_n830), .ZN(new_n831));
  NAND2_X1  g406(.A1(new_n621), .A2(G16), .ZN(new_n832));
  OAI21_X1  g407(.A(new_n832), .B1(G4), .B2(G16), .ZN(new_n833));
  INV_X1    g408(.A(G1348), .ZN(new_n834));
  OR2_X1    g409(.A1(new_n833), .A2(new_n834), .ZN(new_n835));
  NAND2_X1  g410(.A1(new_n716), .A2(G27), .ZN(new_n836));
  XOR2_X1   g411(.A(new_n836), .B(KEYINPUT103), .Z(new_n837));
  NAND2_X1  g412(.A1(new_n502), .A2(KEYINPUT71), .ZN(new_n838));
  NAND2_X1  g413(.A1(new_n503), .A2(KEYINPUT4), .ZN(new_n839));
  NAND3_X1  g414(.A1(new_n838), .A2(new_n506), .A3(new_n839), .ZN(new_n840));
  INV_X1    g415(.A(new_n499), .ZN(new_n841));
  NAND2_X1  g416(.A1(new_n840), .A2(new_n841), .ZN(new_n842));
  AOI21_X1  g417(.A(new_n837), .B1(new_n842), .B2(new_n715), .ZN(new_n843));
  XNOR2_X1  g418(.A(new_n843), .B(G2078), .ZN(new_n844));
  NAND2_X1  g419(.A1(new_n833), .A2(new_n834), .ZN(new_n845));
  AND3_X1   g420(.A1(new_n835), .A2(new_n844), .A3(new_n845), .ZN(new_n846));
  NAND4_X1  g421(.A1(new_n795), .A2(new_n829), .A3(new_n831), .A4(new_n846), .ZN(G150));
  INV_X1    g422(.A(G150), .ZN(G311));
  NAND2_X1  g423(.A1(new_n621), .A2(G559), .ZN(new_n849));
  XNOR2_X1  g424(.A(new_n849), .B(KEYINPUT38), .ZN(new_n850));
  INV_X1    g425(.A(new_n560), .ZN(new_n851));
  AOI22_X1  g426(.A1(new_n513), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n852));
  OR2_X1    g427(.A1(new_n852), .A2(new_n515), .ZN(new_n853));
  NAND2_X1  g428(.A1(new_n520), .A2(G55), .ZN(new_n854));
  INV_X1    g429(.A(G93), .ZN(new_n855));
  OAI21_X1  g430(.A(new_n854), .B1(new_n523), .B2(new_n855), .ZN(new_n856));
  INV_X1    g431(.A(new_n856), .ZN(new_n857));
  NAND4_X1  g432(.A1(new_n851), .A2(new_n853), .A3(new_n557), .A4(new_n857), .ZN(new_n858));
  NOR2_X1   g433(.A1(new_n852), .A2(new_n515), .ZN(new_n859));
  OAI22_X1  g434(.A1(new_n558), .A2(new_n560), .B1(new_n859), .B2(new_n856), .ZN(new_n860));
  NAND2_X1  g435(.A1(new_n858), .A2(new_n860), .ZN(new_n861));
  INV_X1    g436(.A(new_n861), .ZN(new_n862));
  XNOR2_X1  g437(.A(new_n850), .B(new_n862), .ZN(new_n863));
  NOR2_X1   g438(.A1(new_n863), .A2(KEYINPUT39), .ZN(new_n864));
  XOR2_X1   g439(.A(new_n864), .B(KEYINPUT105), .Z(new_n865));
  AOI21_X1  g440(.A(G860), .B1(new_n863), .B2(KEYINPUT39), .ZN(new_n866));
  NAND2_X1  g441(.A1(new_n865), .A2(new_n866), .ZN(new_n867));
  OAI21_X1  g442(.A(G860), .B1(new_n859), .B2(new_n856), .ZN(new_n868));
  XOR2_X1   g443(.A(new_n868), .B(KEYINPUT37), .Z(new_n869));
  NAND2_X1  g444(.A1(new_n867), .A2(new_n869), .ZN(G145));
  INV_X1    g445(.A(KEYINPUT106), .ZN(new_n871));
  OAI21_X1  g446(.A(new_n727), .B1(new_n777), .B2(new_n871), .ZN(new_n872));
  NAND4_X1  g447(.A1(new_n775), .A2(new_n776), .A3(KEYINPUT106), .A4(new_n726), .ZN(new_n873));
  NAND2_X1  g448(.A1(new_n872), .A2(new_n873), .ZN(new_n874));
  NAND2_X1  g449(.A1(new_n483), .A2(G130), .ZN(new_n875));
  OR2_X1    g450(.A1(G106), .A2(G2105), .ZN(new_n876));
  OAI211_X1 g451(.A(new_n876), .B(G2104), .C1(G118), .C2(new_n462), .ZN(new_n877));
  NAND2_X1  g452(.A1(new_n875), .A2(new_n877), .ZN(new_n878));
  AOI21_X1  g453(.A(new_n878), .B1(G142), .B2(new_n489), .ZN(new_n879));
  XNOR2_X1  g454(.A(new_n879), .B(new_n644), .ZN(new_n880));
  INV_X1    g455(.A(new_n880), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n874), .A2(new_n881), .ZN(new_n882));
  XNOR2_X1  g457(.A(new_n762), .B(new_n842), .ZN(new_n883));
  XNOR2_X1  g458(.A(new_n883), .B(new_n822), .ZN(new_n884));
  INV_X1    g459(.A(new_n884), .ZN(new_n885));
  NAND3_X1  g460(.A1(new_n872), .A2(new_n873), .A3(new_n880), .ZN(new_n886));
  NAND3_X1  g461(.A1(new_n882), .A2(new_n885), .A3(new_n886), .ZN(new_n887));
  AND3_X1   g462(.A1(new_n872), .A2(new_n873), .A3(new_n880), .ZN(new_n888));
  AOI21_X1  g463(.A(new_n880), .B1(new_n872), .B2(new_n873), .ZN(new_n889));
  OAI21_X1  g464(.A(new_n884), .B1(new_n888), .B2(new_n889), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n887), .A2(new_n890), .ZN(new_n891));
  XNOR2_X1  g466(.A(new_n640), .B(G160), .ZN(new_n892));
  XNOR2_X1  g467(.A(new_n892), .B(G162), .ZN(new_n893));
  AOI21_X1  g468(.A(G37), .B1(new_n891), .B2(new_n893), .ZN(new_n894));
  INV_X1    g469(.A(new_n893), .ZN(new_n895));
  NAND3_X1  g470(.A1(new_n895), .A2(new_n887), .A3(new_n890), .ZN(new_n896));
  NAND2_X1  g471(.A1(new_n894), .A2(new_n896), .ZN(new_n897));
  INV_X1    g472(.A(KEYINPUT107), .ZN(new_n898));
  NAND2_X1  g473(.A1(new_n897), .A2(new_n898), .ZN(new_n899));
  NAND3_X1  g474(.A1(new_n894), .A2(KEYINPUT107), .A3(new_n896), .ZN(new_n900));
  AND3_X1   g475(.A1(new_n899), .A2(KEYINPUT40), .A3(new_n900), .ZN(new_n901));
  AOI21_X1  g476(.A(KEYINPUT40), .B1(new_n899), .B2(new_n900), .ZN(new_n902));
  NOR2_X1   g477(.A1(new_n901), .A2(new_n902), .ZN(G395));
  INV_X1    g478(.A(KEYINPUT113), .ZN(new_n904));
  NOR2_X1   g479(.A1(new_n859), .A2(new_n856), .ZN(new_n905));
  OAI21_X1  g480(.A(new_n904), .B1(new_n905), .B2(G868), .ZN(new_n906));
  OR2_X1    g481(.A1(G290), .A2(G288), .ZN(new_n907));
  NAND2_X1  g482(.A1(G290), .A2(G288), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n907), .A2(new_n908), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n909), .A2(KEYINPUT110), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n797), .A2(G166), .ZN(new_n911));
  NAND2_X1  g486(.A1(G305), .A2(G303), .ZN(new_n912));
  NAND3_X1  g487(.A1(new_n910), .A2(new_n911), .A3(new_n912), .ZN(new_n913));
  INV_X1    g488(.A(KEYINPUT110), .ZN(new_n914));
  NAND3_X1  g489(.A1(new_n907), .A2(new_n914), .A3(new_n908), .ZN(new_n915));
  INV_X1    g490(.A(new_n915), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n913), .A2(new_n916), .ZN(new_n917));
  NAND4_X1  g492(.A1(new_n910), .A2(new_n915), .A3(new_n911), .A4(new_n912), .ZN(new_n918));
  NAND2_X1  g493(.A1(new_n917), .A2(new_n918), .ZN(new_n919));
  XNOR2_X1  g494(.A(KEYINPUT111), .B(KEYINPUT42), .ZN(new_n920));
  OR2_X1    g495(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n919), .A2(new_n920), .ZN(new_n922));
  NAND2_X1  g497(.A1(new_n921), .A2(new_n922), .ZN(new_n923));
  INV_X1    g498(.A(KEYINPUT112), .ZN(new_n924));
  AND2_X1   g499(.A1(new_n861), .A2(KEYINPUT108), .ZN(new_n925));
  NOR2_X1   g500(.A1(new_n861), .A2(KEYINPUT108), .ZN(new_n926));
  NOR2_X1   g501(.A1(new_n925), .A2(new_n926), .ZN(new_n927));
  NAND2_X1  g502(.A1(new_n927), .A2(new_n630), .ZN(new_n928));
  OAI21_X1  g503(.A(new_n631), .B1(new_n925), .B2(new_n926), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  AND2_X1   g505(.A1(new_n610), .A2(new_n607), .ZN(new_n931));
  XNOR2_X1  g506(.A(new_n616), .B(KEYINPUT83), .ZN(new_n932));
  NAND3_X1  g507(.A1(new_n931), .A2(new_n932), .A3(new_n625), .ZN(new_n933));
  NAND2_X1  g508(.A1(new_n620), .A2(G299), .ZN(new_n934));
  NAND2_X1  g509(.A1(new_n933), .A2(new_n934), .ZN(new_n935));
  INV_X1    g510(.A(new_n935), .ZN(new_n936));
  NOR2_X1   g511(.A1(new_n930), .A2(new_n936), .ZN(new_n937));
  INV_X1    g512(.A(new_n937), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n935), .A2(KEYINPUT41), .ZN(new_n939));
  INV_X1    g514(.A(KEYINPUT109), .ZN(new_n940));
  INV_X1    g515(.A(KEYINPUT41), .ZN(new_n941));
  NAND3_X1  g516(.A1(new_n933), .A2(new_n934), .A3(new_n941), .ZN(new_n942));
  NAND3_X1  g517(.A1(new_n939), .A2(new_n940), .A3(new_n942), .ZN(new_n943));
  NAND3_X1  g518(.A1(new_n936), .A2(KEYINPUT109), .A3(new_n941), .ZN(new_n944));
  NAND2_X1  g519(.A1(new_n943), .A2(new_n944), .ZN(new_n945));
  NAND2_X1  g520(.A1(new_n945), .A2(new_n930), .ZN(new_n946));
  NAND4_X1  g521(.A1(new_n923), .A2(new_n924), .A3(new_n938), .A4(new_n946), .ZN(new_n947));
  AND2_X1   g522(.A1(new_n947), .A2(G868), .ZN(new_n948));
  INV_X1    g523(.A(new_n946), .ZN(new_n949));
  OAI21_X1  g524(.A(KEYINPUT112), .B1(new_n949), .B2(new_n937), .ZN(new_n950));
  NAND3_X1  g525(.A1(new_n938), .A2(new_n924), .A3(new_n946), .ZN(new_n951));
  NAND4_X1  g526(.A1(new_n950), .A2(new_n921), .A3(new_n922), .A4(new_n951), .ZN(new_n952));
  AOI21_X1  g527(.A(new_n906), .B1(new_n948), .B2(new_n952), .ZN(new_n953));
  AND2_X1   g528(.A1(new_n948), .A2(new_n952), .ZN(new_n954));
  AOI21_X1  g529(.A(new_n953), .B1(KEYINPUT113), .B2(new_n954), .ZN(G295));
  AOI21_X1  g530(.A(new_n953), .B1(KEYINPUT113), .B2(new_n954), .ZN(G331));
  NAND2_X1  g531(.A1(G286), .A2(G301), .ZN(new_n957));
  AOI22_X1  g532(.A1(new_n532), .A2(new_n533), .B1(new_n544), .B2(new_n546), .ZN(new_n958));
  AND2_X1   g533(.A1(new_n535), .A2(new_n538), .ZN(new_n959));
  NAND3_X1  g534(.A1(G171), .A2(new_n958), .A3(new_n959), .ZN(new_n960));
  AND4_X1   g535(.A1(new_n860), .A2(new_n957), .A3(new_n960), .A4(new_n858), .ZN(new_n961));
  AOI22_X1  g536(.A1(new_n957), .A2(new_n960), .B1(new_n858), .B2(new_n860), .ZN(new_n962));
  OAI21_X1  g537(.A(KEYINPUT114), .B1(new_n961), .B2(new_n962), .ZN(new_n963));
  INV_X1    g538(.A(KEYINPUT114), .ZN(new_n964));
  AOI21_X1  g539(.A(G171), .B1(new_n959), .B2(new_n958), .ZN(new_n965));
  NOR2_X1   g540(.A1(G286), .A2(G301), .ZN(new_n966));
  OAI21_X1  g541(.A(new_n861), .B1(new_n965), .B2(new_n966), .ZN(new_n967));
  OAI21_X1  g542(.A(new_n964), .B1(new_n967), .B2(new_n862), .ZN(new_n968));
  NAND2_X1  g543(.A1(new_n963), .A2(new_n968), .ZN(new_n969));
  NAND3_X1  g544(.A1(new_n943), .A2(new_n969), .A3(new_n944), .ZN(new_n970));
  NAND4_X1  g545(.A1(new_n957), .A2(new_n960), .A3(new_n860), .A4(new_n858), .ZN(new_n971));
  NAND4_X1  g546(.A1(new_n967), .A2(new_n934), .A3(new_n933), .A4(new_n971), .ZN(new_n972));
  XNOR2_X1  g547(.A(new_n972), .B(KEYINPUT115), .ZN(new_n973));
  NAND2_X1  g548(.A1(new_n970), .A2(new_n973), .ZN(new_n974));
  NOR2_X1   g549(.A1(new_n974), .A2(new_n919), .ZN(new_n975));
  AOI21_X1  g550(.A(G37), .B1(new_n974), .B2(new_n919), .ZN(new_n976));
  AOI21_X1  g551(.A(new_n975), .B1(new_n976), .B2(KEYINPUT116), .ZN(new_n977));
  INV_X1    g552(.A(KEYINPUT116), .ZN(new_n978));
  INV_X1    g553(.A(new_n919), .ZN(new_n979));
  AOI21_X1  g554(.A(new_n979), .B1(new_n970), .B2(new_n973), .ZN(new_n980));
  OAI21_X1  g555(.A(new_n978), .B1(new_n980), .B2(G37), .ZN(new_n981));
  AOI21_X1  g556(.A(KEYINPUT43), .B1(new_n977), .B2(new_n981), .ZN(new_n982));
  INV_X1    g557(.A(KEYINPUT117), .ZN(new_n983));
  NAND2_X1  g558(.A1(new_n942), .A2(new_n983), .ZN(new_n984));
  NAND4_X1  g559(.A1(new_n933), .A2(new_n934), .A3(KEYINPUT117), .A4(new_n941), .ZN(new_n985));
  NAND3_X1  g560(.A1(new_n984), .A2(new_n939), .A3(new_n985), .ZN(new_n986));
  NAND2_X1  g561(.A1(new_n967), .A2(new_n971), .ZN(new_n987));
  NAND2_X1  g562(.A1(new_n986), .A2(new_n987), .ZN(new_n988));
  OR2_X1    g563(.A1(new_n988), .A2(KEYINPUT118), .ZN(new_n989));
  NOR2_X1   g564(.A1(new_n969), .A2(new_n935), .ZN(new_n990));
  AOI21_X1  g565(.A(new_n990), .B1(new_n988), .B2(KEYINPUT118), .ZN(new_n991));
  AOI21_X1  g566(.A(new_n979), .B1(new_n989), .B2(new_n991), .ZN(new_n992));
  INV_X1    g567(.A(KEYINPUT43), .ZN(new_n993));
  INV_X1    g568(.A(G37), .ZN(new_n994));
  OAI21_X1  g569(.A(new_n994), .B1(new_n974), .B2(new_n919), .ZN(new_n995));
  NOR3_X1   g570(.A1(new_n992), .A2(new_n993), .A3(new_n995), .ZN(new_n996));
  OAI21_X1  g571(.A(KEYINPUT44), .B1(new_n982), .B2(new_n996), .ZN(new_n997));
  INV_X1    g572(.A(KEYINPUT44), .ZN(new_n998));
  AOI21_X1  g573(.A(new_n993), .B1(new_n977), .B2(new_n981), .ZN(new_n999));
  NOR3_X1   g574(.A1(new_n992), .A2(KEYINPUT43), .A3(new_n995), .ZN(new_n1000));
  OAI21_X1  g575(.A(new_n998), .B1(new_n999), .B2(new_n1000), .ZN(new_n1001));
  NAND2_X1  g576(.A1(new_n997), .A2(new_n1001), .ZN(G397));
  AOI21_X1  g577(.A(G1384), .B1(new_n840), .B2(new_n841), .ZN(new_n1003));
  INV_X1    g578(.A(KEYINPUT50), .ZN(new_n1004));
  NAND2_X1  g579(.A1(new_n1003), .A2(new_n1004), .ZN(new_n1005));
  OAI21_X1  g580(.A(KEYINPUT50), .B1(G164), .B2(G1384), .ZN(new_n1006));
  INV_X1    g581(.A(G40), .ZN(new_n1007));
  NOR3_X1   g582(.A1(new_n474), .A2(new_n480), .A3(new_n1007), .ZN(new_n1008));
  NAND3_X1  g583(.A1(new_n1005), .A2(new_n1006), .A3(new_n1008), .ZN(new_n1009));
  INV_X1    g584(.A(G1956), .ZN(new_n1010));
  NAND2_X1  g585(.A1(new_n1009), .A2(new_n1010), .ZN(new_n1011));
  INV_X1    g586(.A(new_n1008), .ZN(new_n1012));
  INV_X1    g587(.A(G1384), .ZN(new_n1013));
  NAND2_X1  g588(.A1(new_n842), .A2(new_n1013), .ZN(new_n1014));
  INV_X1    g589(.A(KEYINPUT45), .ZN(new_n1015));
  AOI21_X1  g590(.A(new_n1012), .B1(new_n1014), .B2(new_n1015), .ZN(new_n1016));
  NAND3_X1  g591(.A1(new_n842), .A2(KEYINPUT45), .A3(new_n1013), .ZN(new_n1017));
  XNOR2_X1  g592(.A(KEYINPUT56), .B(G2072), .ZN(new_n1018));
  NAND3_X1  g593(.A1(new_n1016), .A2(new_n1017), .A3(new_n1018), .ZN(new_n1019));
  XNOR2_X1  g594(.A(G299), .B(KEYINPUT57), .ZN(new_n1020));
  INV_X1    g595(.A(new_n1020), .ZN(new_n1021));
  NAND3_X1  g596(.A1(new_n1011), .A2(new_n1019), .A3(new_n1021), .ZN(new_n1022));
  NAND2_X1  g597(.A1(new_n1022), .A2(KEYINPUT122), .ZN(new_n1023));
  INV_X1    g598(.A(KEYINPUT122), .ZN(new_n1024));
  NAND4_X1  g599(.A1(new_n1011), .A2(new_n1019), .A3(new_n1021), .A4(new_n1024), .ZN(new_n1025));
  NAND2_X1  g600(.A1(new_n1023), .A2(new_n1025), .ZN(new_n1026));
  AOI21_X1  g601(.A(new_n1012), .B1(new_n1014), .B2(KEYINPUT50), .ZN(new_n1027));
  AOI21_X1  g602(.A(G1956), .B1(new_n1027), .B2(new_n1005), .ZN(new_n1028));
  OAI21_X1  g603(.A(new_n1015), .B1(G164), .B2(G1384), .ZN(new_n1029));
  AND4_X1   g604(.A1(new_n1008), .A2(new_n1029), .A3(new_n1017), .A4(new_n1018), .ZN(new_n1030));
  OAI21_X1  g605(.A(new_n1020), .B1(new_n1028), .B2(new_n1030), .ZN(new_n1031));
  INV_X1    g606(.A(new_n1031), .ZN(new_n1032));
  NAND2_X1  g607(.A1(new_n1009), .A2(new_n834), .ZN(new_n1033));
  INV_X1    g608(.A(G2067), .ZN(new_n1034));
  NAND3_X1  g609(.A1(new_n1003), .A2(new_n1034), .A3(new_n1008), .ZN(new_n1035));
  AOI21_X1  g610(.A(new_n620), .B1(new_n1033), .B2(new_n1035), .ZN(new_n1036));
  OAI21_X1  g611(.A(new_n1026), .B1(new_n1032), .B2(new_n1036), .ZN(new_n1037));
  NAND3_X1  g612(.A1(new_n1031), .A2(KEYINPUT61), .A3(new_n1022), .ZN(new_n1038));
  NAND2_X1  g613(.A1(new_n1038), .A2(KEYINPUT123), .ZN(new_n1039));
  AND3_X1   g614(.A1(new_n1033), .A2(new_n620), .A3(new_n1035), .ZN(new_n1040));
  OAI21_X1  g615(.A(KEYINPUT60), .B1(new_n1040), .B2(new_n1036), .ZN(new_n1041));
  NOR2_X1   g616(.A1(new_n620), .A2(KEYINPUT60), .ZN(new_n1042));
  AND3_X1   g617(.A1(new_n1033), .A2(new_n1035), .A3(new_n1042), .ZN(new_n1043));
  INV_X1    g618(.A(G1996), .ZN(new_n1044));
  NAND4_X1  g619(.A1(new_n1029), .A2(new_n1017), .A3(new_n1044), .A4(new_n1008), .ZN(new_n1045));
  NAND2_X1  g620(.A1(new_n1003), .A2(new_n1008), .ZN(new_n1046));
  XOR2_X1   g621(.A(KEYINPUT58), .B(G1341), .Z(new_n1047));
  NAND2_X1  g622(.A1(new_n1046), .A2(new_n1047), .ZN(new_n1048));
  NAND2_X1  g623(.A1(new_n1045), .A2(new_n1048), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n1049), .A2(new_n561), .ZN(new_n1050));
  NAND2_X1  g625(.A1(new_n1050), .A2(KEYINPUT59), .ZN(new_n1051));
  INV_X1    g626(.A(KEYINPUT59), .ZN(new_n1052));
  NAND3_X1  g627(.A1(new_n1049), .A2(new_n1052), .A3(new_n561), .ZN(new_n1053));
  AOI21_X1  g628(.A(new_n1043), .B1(new_n1051), .B2(new_n1053), .ZN(new_n1054));
  INV_X1    g629(.A(KEYINPUT123), .ZN(new_n1055));
  NAND4_X1  g630(.A1(new_n1031), .A2(new_n1022), .A3(new_n1055), .A4(KEYINPUT61), .ZN(new_n1056));
  NAND4_X1  g631(.A1(new_n1039), .A2(new_n1041), .A3(new_n1054), .A4(new_n1056), .ZN(new_n1057));
  AOI21_X1  g632(.A(KEYINPUT61), .B1(new_n1026), .B2(new_n1031), .ZN(new_n1058));
  OAI21_X1  g633(.A(new_n1037), .B1(new_n1057), .B2(new_n1058), .ZN(new_n1059));
  INV_X1    g634(.A(G2078), .ZN(new_n1060));
  NAND4_X1  g635(.A1(new_n1029), .A2(new_n1017), .A3(new_n1060), .A4(new_n1008), .ZN(new_n1061));
  INV_X1    g636(.A(KEYINPUT53), .ZN(new_n1062));
  NAND2_X1  g637(.A1(new_n1061), .A2(new_n1062), .ZN(new_n1063));
  INV_X1    g638(.A(G1961), .ZN(new_n1064));
  NAND2_X1  g639(.A1(new_n1009), .A2(new_n1064), .ZN(new_n1065));
  INV_X1    g640(.A(new_n474), .ZN(new_n1066));
  INV_X1    g641(.A(new_n480), .ZN(new_n1067));
  OR2_X1    g642(.A1(KEYINPUT124), .A2(G2078), .ZN(new_n1068));
  NAND2_X1  g643(.A1(KEYINPUT124), .A2(G2078), .ZN(new_n1069));
  AOI21_X1  g644(.A(new_n1062), .B1(new_n1068), .B2(new_n1069), .ZN(new_n1070));
  NAND4_X1  g645(.A1(new_n1066), .A2(G40), .A3(new_n1067), .A4(new_n1070), .ZN(new_n1071));
  AOI21_X1  g646(.A(new_n1071), .B1(new_n1003), .B2(KEYINPUT45), .ZN(new_n1072));
  NOR2_X1   g647(.A1(new_n1014), .A2(KEYINPUT119), .ZN(new_n1073));
  INV_X1    g648(.A(KEYINPUT119), .ZN(new_n1074));
  OAI21_X1  g649(.A(new_n1015), .B1(new_n1003), .B2(new_n1074), .ZN(new_n1075));
  OAI21_X1  g650(.A(new_n1072), .B1(new_n1073), .B2(new_n1075), .ZN(new_n1076));
  NAND3_X1  g651(.A1(new_n1063), .A2(new_n1065), .A3(new_n1076), .ZN(new_n1077));
  INV_X1    g652(.A(KEYINPUT125), .ZN(new_n1078));
  NAND2_X1  g653(.A1(new_n1077), .A2(new_n1078), .ZN(new_n1079));
  NAND4_X1  g654(.A1(new_n1063), .A2(new_n1065), .A3(new_n1076), .A4(KEYINPUT125), .ZN(new_n1080));
  NAND3_X1  g655(.A1(new_n1079), .A2(G171), .A3(new_n1080), .ZN(new_n1081));
  NAND4_X1  g656(.A1(new_n1016), .A2(KEYINPUT53), .A3(new_n1060), .A4(new_n1017), .ZN(new_n1082));
  NAND4_X1  g657(.A1(new_n1082), .A2(new_n1063), .A3(new_n1065), .A4(G301), .ZN(new_n1083));
  AND2_X1   g658(.A1(new_n1083), .A2(KEYINPUT54), .ZN(new_n1084));
  NAND2_X1  g659(.A1(new_n1081), .A2(new_n1084), .ZN(new_n1085));
  OAI21_X1  g660(.A(new_n1008), .B1(new_n1003), .B2(KEYINPUT45), .ZN(new_n1086));
  NOR3_X1   g661(.A1(G164), .A2(new_n1015), .A3(G1384), .ZN(new_n1087));
  OAI21_X1  g662(.A(new_n746), .B1(new_n1086), .B2(new_n1087), .ZN(new_n1088));
  INV_X1    g663(.A(G2084), .ZN(new_n1089));
  NAND4_X1  g664(.A1(new_n1005), .A2(new_n1006), .A3(new_n1089), .A4(new_n1008), .ZN(new_n1090));
  NAND3_X1  g665(.A1(new_n1088), .A2(G168), .A3(new_n1090), .ZN(new_n1091));
  NAND2_X1  g666(.A1(new_n1091), .A2(G8), .ZN(new_n1092));
  AOI21_X1  g667(.A(G168), .B1(new_n1088), .B2(new_n1090), .ZN(new_n1093));
  OAI21_X1  g668(.A(KEYINPUT51), .B1(new_n1092), .B2(new_n1093), .ZN(new_n1094));
  INV_X1    g669(.A(KEYINPUT51), .ZN(new_n1095));
  NAND3_X1  g670(.A1(new_n1091), .A2(new_n1095), .A3(G8), .ZN(new_n1096));
  NAND2_X1  g671(.A1(new_n1094), .A2(new_n1096), .ZN(new_n1097));
  INV_X1    g672(.A(KEYINPUT54), .ZN(new_n1098));
  NOR2_X1   g673(.A1(new_n1077), .A2(G171), .ZN(new_n1099));
  AOI22_X1  g674(.A1(new_n1062), .A2(new_n1061), .B1(new_n1009), .B2(new_n1064), .ZN(new_n1100));
  AOI21_X1  g675(.A(G301), .B1(new_n1100), .B2(new_n1082), .ZN(new_n1101));
  OAI21_X1  g676(.A(new_n1098), .B1(new_n1099), .B2(new_n1101), .ZN(new_n1102));
  NAND2_X1  g677(.A1(new_n807), .A2(G1976), .ZN(new_n1103));
  NAND3_X1  g678(.A1(new_n1046), .A2(G8), .A3(new_n1103), .ZN(new_n1104));
  NAND2_X1  g679(.A1(new_n1104), .A2(KEYINPUT52), .ZN(new_n1105));
  INV_X1    g680(.A(G8), .ZN(new_n1106));
  AOI21_X1  g681(.A(new_n1106), .B1(new_n1003), .B2(new_n1008), .ZN(new_n1107));
  INV_X1    g682(.A(G1976), .ZN(new_n1108));
  AOI21_X1  g683(.A(KEYINPUT52), .B1(G288), .B2(new_n1108), .ZN(new_n1109));
  NAND3_X1  g684(.A1(new_n1107), .A2(new_n1103), .A3(new_n1109), .ZN(new_n1110));
  INV_X1    g685(.A(KEYINPUT49), .ZN(new_n1111));
  AOI211_X1 g686(.A(G1981), .B(new_n596), .C1(new_n590), .C2(new_n592), .ZN(new_n1112));
  INV_X1    g687(.A(G1981), .ZN(new_n1113));
  AOI21_X1  g688(.A(new_n1113), .B1(new_n597), .B2(new_n589), .ZN(new_n1114));
  OAI21_X1  g689(.A(new_n1111), .B1(new_n1112), .B2(new_n1114), .ZN(new_n1115));
  NAND3_X1  g690(.A1(new_n593), .A2(new_n1113), .A3(new_n597), .ZN(new_n1116));
  NAND2_X1  g691(.A1(new_n597), .A2(new_n589), .ZN(new_n1117));
  NAND2_X1  g692(.A1(new_n1117), .A2(G1981), .ZN(new_n1118));
  NAND3_X1  g693(.A1(new_n1116), .A2(KEYINPUT49), .A3(new_n1118), .ZN(new_n1119));
  NAND3_X1  g694(.A1(new_n1115), .A2(new_n1107), .A3(new_n1119), .ZN(new_n1120));
  AND3_X1   g695(.A1(new_n1105), .A2(new_n1110), .A3(new_n1120), .ZN(new_n1121));
  AOI21_X1  g696(.A(KEYINPUT55), .B1(G303), .B2(G8), .ZN(new_n1122));
  INV_X1    g697(.A(KEYINPUT55), .ZN(new_n1123));
  NOR3_X1   g698(.A1(G166), .A2(new_n1123), .A3(new_n1106), .ZN(new_n1124));
  NOR2_X1   g699(.A1(new_n1122), .A2(new_n1124), .ZN(new_n1125));
  INV_X1    g700(.A(new_n1125), .ZN(new_n1126));
  OAI21_X1  g701(.A(new_n804), .B1(new_n1086), .B2(new_n1087), .ZN(new_n1127));
  NAND4_X1  g702(.A1(new_n1005), .A2(new_n1006), .A3(new_n790), .A4(new_n1008), .ZN(new_n1128));
  AOI21_X1  g703(.A(new_n1106), .B1(new_n1127), .B2(new_n1128), .ZN(new_n1129));
  OAI21_X1  g704(.A(new_n1121), .B1(new_n1126), .B2(new_n1129), .ZN(new_n1130));
  AOI211_X1 g705(.A(new_n1106), .B(new_n1125), .C1(new_n1127), .C2(new_n1128), .ZN(new_n1131));
  NOR2_X1   g706(.A1(new_n1130), .A2(new_n1131), .ZN(new_n1132));
  AND4_X1   g707(.A1(new_n1085), .A2(new_n1097), .A3(new_n1102), .A4(new_n1132), .ZN(new_n1133));
  NAND2_X1  g708(.A1(new_n1059), .A2(new_n1133), .ZN(new_n1134));
  NAND2_X1  g709(.A1(new_n1131), .A2(new_n1121), .ZN(new_n1135));
  INV_X1    g710(.A(new_n1107), .ZN(new_n1136));
  NOR2_X1   g711(.A1(G288), .A2(G1976), .ZN(new_n1137));
  AOI21_X1  g712(.A(new_n1112), .B1(new_n1120), .B2(new_n1137), .ZN(new_n1138));
  OAI21_X1  g713(.A(new_n1135), .B1(new_n1136), .B2(new_n1138), .ZN(new_n1139));
  AOI211_X1 g714(.A(new_n1106), .B(G286), .C1(new_n1088), .C2(new_n1090), .ZN(new_n1140));
  NAND3_X1  g715(.A1(new_n1132), .A2(KEYINPUT63), .A3(new_n1140), .ZN(new_n1141));
  OR2_X1    g716(.A1(new_n1129), .A2(new_n1126), .ZN(new_n1142));
  INV_X1    g717(.A(new_n1131), .ZN(new_n1143));
  NAND4_X1  g718(.A1(new_n1142), .A2(new_n1143), .A3(new_n1121), .A4(new_n1140), .ZN(new_n1144));
  INV_X1    g719(.A(KEYINPUT63), .ZN(new_n1145));
  NAND2_X1  g720(.A1(new_n1144), .A2(new_n1145), .ZN(new_n1146));
  AOI21_X1  g721(.A(new_n1139), .B1(new_n1141), .B2(new_n1146), .ZN(new_n1147));
  INV_X1    g722(.A(KEYINPUT126), .ZN(new_n1148));
  NAND3_X1  g723(.A1(new_n1082), .A2(new_n1063), .A3(new_n1065), .ZN(new_n1149));
  NAND2_X1  g724(.A1(new_n1149), .A2(G171), .ZN(new_n1150));
  NOR3_X1   g725(.A1(new_n1130), .A2(new_n1150), .A3(new_n1131), .ZN(new_n1151));
  AND3_X1   g726(.A1(new_n1091), .A2(new_n1095), .A3(G8), .ZN(new_n1152));
  NAND2_X1  g727(.A1(new_n1088), .A2(new_n1090), .ZN(new_n1153));
  NAND2_X1  g728(.A1(new_n1153), .A2(G286), .ZN(new_n1154));
  NAND3_X1  g729(.A1(new_n1154), .A2(G8), .A3(new_n1091), .ZN(new_n1155));
  AOI21_X1  g730(.A(new_n1152), .B1(new_n1155), .B2(KEYINPUT51), .ZN(new_n1156));
  INV_X1    g731(.A(KEYINPUT62), .ZN(new_n1157));
  OAI21_X1  g732(.A(new_n1151), .B1(new_n1156), .B2(new_n1157), .ZN(new_n1158));
  NOR2_X1   g733(.A1(new_n1097), .A2(KEYINPUT62), .ZN(new_n1159));
  OAI21_X1  g734(.A(new_n1148), .B1(new_n1158), .B2(new_n1159), .ZN(new_n1160));
  NAND2_X1  g735(.A1(new_n1156), .A2(new_n1157), .ZN(new_n1161));
  NAND2_X1  g736(.A1(new_n1097), .A2(KEYINPUT62), .ZN(new_n1162));
  NAND4_X1  g737(.A1(new_n1161), .A2(new_n1162), .A3(KEYINPUT126), .A4(new_n1151), .ZN(new_n1163));
  NAND4_X1  g738(.A1(new_n1134), .A2(new_n1147), .A3(new_n1160), .A4(new_n1163), .ZN(new_n1164));
  NOR3_X1   g739(.A1(new_n1073), .A2(new_n1075), .A3(new_n1012), .ZN(new_n1165));
  NAND3_X1  g740(.A1(new_n1165), .A2(new_n1044), .A3(new_n727), .ZN(new_n1166));
  XOR2_X1   g741(.A(new_n1166), .B(KEYINPUT120), .Z(new_n1167));
  XNOR2_X1  g742(.A(new_n762), .B(G2067), .ZN(new_n1168));
  OAI21_X1  g743(.A(new_n1168), .B1(new_n1044), .B2(new_n727), .ZN(new_n1169));
  NAND2_X1  g744(.A1(new_n1165), .A2(new_n1169), .ZN(new_n1170));
  INV_X1    g745(.A(new_n1165), .ZN(new_n1171));
  XNOR2_X1  g746(.A(new_n822), .B(new_n824), .ZN(new_n1172));
  XNOR2_X1  g747(.A(new_n1172), .B(KEYINPUT121), .ZN(new_n1173));
  OAI211_X1 g748(.A(new_n1167), .B(new_n1170), .C1(new_n1171), .C2(new_n1173), .ZN(new_n1174));
  XNOR2_X1  g749(.A(G290), .B(G1986), .ZN(new_n1175));
  AOI21_X1  g750(.A(new_n1174), .B1(new_n1165), .B2(new_n1175), .ZN(new_n1176));
  NAND2_X1  g751(.A1(new_n1164), .A2(new_n1176), .ZN(new_n1177));
  INV_X1    g752(.A(KEYINPUT46), .ZN(new_n1178));
  OAI21_X1  g753(.A(new_n1178), .B1(new_n1171), .B2(G1996), .ZN(new_n1179));
  OR2_X1    g754(.A1(new_n1179), .A2(KEYINPUT127), .ZN(new_n1180));
  NAND2_X1  g755(.A1(new_n1179), .A2(KEYINPUT127), .ZN(new_n1181));
  OAI211_X1 g756(.A(new_n1168), .B(new_n727), .C1(new_n1178), .C2(G1996), .ZN(new_n1182));
  AOI22_X1  g757(.A1(new_n1180), .A2(new_n1181), .B1(new_n1165), .B2(new_n1182), .ZN(new_n1183));
  INV_X1    g758(.A(KEYINPUT47), .ZN(new_n1184));
  AND2_X1   g759(.A1(new_n1183), .A2(new_n1184), .ZN(new_n1185));
  NOR2_X1   g760(.A1(new_n1183), .A2(new_n1184), .ZN(new_n1186));
  NOR3_X1   g761(.A1(new_n1171), .A2(G1986), .A3(G290), .ZN(new_n1187));
  XNOR2_X1  g762(.A(new_n1187), .B(KEYINPUT48), .ZN(new_n1188));
  OAI22_X1  g763(.A1(new_n1185), .A2(new_n1186), .B1(new_n1174), .B2(new_n1188), .ZN(new_n1189));
  NOR2_X1   g764(.A1(new_n822), .A2(new_n824), .ZN(new_n1190));
  NAND3_X1  g765(.A1(new_n1167), .A2(new_n1170), .A3(new_n1190), .ZN(new_n1191));
  NAND2_X1  g766(.A1(new_n762), .A2(new_n1034), .ZN(new_n1192));
  AOI21_X1  g767(.A(new_n1171), .B1(new_n1191), .B2(new_n1192), .ZN(new_n1193));
  NOR2_X1   g768(.A1(new_n1189), .A2(new_n1193), .ZN(new_n1194));
  NAND2_X1  g769(.A1(new_n1177), .A2(new_n1194), .ZN(G329));
  assign    G231 = 1'b0;
  NOR2_X1   g770(.A1(new_n999), .A2(new_n1000), .ZN(new_n1197));
  NOR2_X1   g771(.A1(G401), .A2(new_n460), .ZN(new_n1198));
  AND3_X1   g772(.A1(new_n704), .A2(new_n685), .A3(new_n1198), .ZN(new_n1199));
  INV_X1    g773(.A(new_n900), .ZN(new_n1200));
  AOI21_X1  g774(.A(KEYINPUT107), .B1(new_n894), .B2(new_n896), .ZN(new_n1201));
  OAI21_X1  g775(.A(new_n1199), .B1(new_n1200), .B2(new_n1201), .ZN(new_n1202));
  NOR2_X1   g776(.A1(new_n1197), .A2(new_n1202), .ZN(G308));
  OAI221_X1 g777(.A(new_n1199), .B1(new_n1200), .B2(new_n1201), .C1(new_n999), .C2(new_n1000), .ZN(G225));
endmodule


