

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n523, n524, n525, n526,
         n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537,
         n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548,
         n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559,
         n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570,
         n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581,
         n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592,
         n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603,
         n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614,
         n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625,
         n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636,
         n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647,
         n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658,
         n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669,
         n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680,
         n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691,
         n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702,
         n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713,
         n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724,
         n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735,
         n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746,
         n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757,
         n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768,
         n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, n779,
         n780, n781, n782, n783, n784, n785, n786, n787, n788, n789, n790,
         n791, n792, n793, n794, n795, n796, n797, n798, n799, n800, n801,
         n802, n803, n804, n805, n806, n807, n808, n809, n810, n811, n812,
         n813, n814, n815, n816, n817, n818, n819, n820, n821, n822, n823,
         n824, n825, n826, n827, n828, n829, n830, n831, n832, n833, n834,
         n835, n836, n837, n838, n839, n840, n841, n842, n843, n844, n845,
         n846, n847, n848, n849, n850, n851, n852, n853, n854, n855, n856,
         n857, n858, n859, n860, n861, n862, n863, n864, n865, n866, n867,
         n868, n869, n870, n871, n872, n873, n874, n875, n876, n877, n878,
         n879, n880, n881, n882, n883, n884, n885, n886, n887, n888, n889,
         n890, n891, n892, n893, n894, n895, n896, n897, n898, n899, n900,
         n901, n902, n903, n904, n905, n906, n907, n908, n909, n910, n911,
         n912, n913, n914, n915, n916, n917, n918, n919, n920, n921, n922,
         n923, n924, n925, n926, n927, n928, n929, n930, n931, n932, n933,
         n934, n935, n936, n937, n938, n939, n940, n941, n942, n943, n944,
         n945, n946, n947, n948, n949, n950, n951, n952, n953, n954, n955,
         n956, n957, n958, n959, n960, n961, n962, n963, n964, n965, n966,
         n967, n968, n969, n970, n971, n972, n973, n974, n975, n976, n977,
         n978, n979, n980, n981, n982, n983, n984, n985, n986, n987, n988,
         n989, n990, n991, n992, n993, n994, n995, n996, n997, n998, n999,
         n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009,
         n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019,
         n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029,
         n1030, n1031, n1032;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  AND2_X1 U556 ( .A1(n526), .A2(G2105), .ZN(n887) );
  XNOR2_X1 U557 ( .A(n727), .B(n726), .ZN(n728) );
  NOR2_X1 U558 ( .A1(n813), .A2(n812), .ZN(n523) );
  AND2_X1 U559 ( .A1(n698), .A2(n763), .ZN(n714) );
  NOR2_X1 U560 ( .A1(n705), .A2(n704), .ZN(n706) );
  OR2_X1 U561 ( .A1(n706), .A2(n920), .ZN(n712) );
  XNOR2_X1 U562 ( .A(n731), .B(KEYINPUT30), .ZN(n732) );
  XNOR2_X1 U563 ( .A(n733), .B(n732), .ZN(n734) );
  INV_X1 U564 ( .A(KEYINPUT29), .ZN(n726) );
  NOR2_X1 U565 ( .A1(n737), .A2(n736), .ZN(n738) );
  NAND2_X1 U566 ( .A1(n698), .A2(n763), .ZN(n740) );
  NOR2_X1 U567 ( .A1(G651), .A2(n650), .ZN(n655) );
  XNOR2_X2 U568 ( .A(G2104), .B(KEYINPUT65), .ZN(n526) );
  NOR2_X4 U569 ( .A1(n526), .A2(G2105), .ZN(n892) );
  NAND2_X1 U570 ( .A1(n892), .A2(G101), .ZN(n525) );
  INV_X1 U571 ( .A(KEYINPUT23), .ZN(n524) );
  XNOR2_X1 U572 ( .A(n525), .B(n524), .ZN(n528) );
  NAND2_X1 U573 ( .A1(n887), .A2(G125), .ZN(n527) );
  NAND2_X1 U574 ( .A1(n528), .A2(n527), .ZN(n529) );
  XNOR2_X1 U575 ( .A(n529), .B(KEYINPUT66), .ZN(n534) );
  NOR2_X1 U576 ( .A1(G2105), .A2(G2104), .ZN(n530) );
  XOR2_X1 U577 ( .A(KEYINPUT17), .B(n530), .Z(n891) );
  NAND2_X1 U578 ( .A1(G137), .A2(n891), .ZN(n532) );
  AND2_X1 U579 ( .A1(G2105), .A2(G2104), .ZN(n888) );
  NAND2_X1 U580 ( .A1(G113), .A2(n888), .ZN(n531) );
  NAND2_X1 U581 ( .A1(n532), .A2(n531), .ZN(n533) );
  NOR2_X1 U582 ( .A1(n534), .A2(n533), .ZN(n535) );
  XNOR2_X2 U583 ( .A(n535), .B(KEYINPUT64), .ZN(G160) );
  XOR2_X1 U584 ( .A(G2443), .B(G2446), .Z(n537) );
  XNOR2_X1 U585 ( .A(G2427), .B(G2451), .ZN(n536) );
  XNOR2_X1 U586 ( .A(n537), .B(n536), .ZN(n543) );
  XOR2_X1 U587 ( .A(G2430), .B(G2454), .Z(n539) );
  XNOR2_X1 U588 ( .A(G1341), .B(G1348), .ZN(n538) );
  XNOR2_X1 U589 ( .A(n539), .B(n538), .ZN(n541) );
  XOR2_X1 U590 ( .A(G2435), .B(G2438), .Z(n540) );
  XNOR2_X1 U591 ( .A(n541), .B(n540), .ZN(n542) );
  XOR2_X1 U592 ( .A(n543), .B(n542), .Z(n544) );
  AND2_X1 U593 ( .A1(G14), .A2(n544), .ZN(G401) );
  XOR2_X1 U594 ( .A(KEYINPUT0), .B(G543), .Z(n650) );
  NAND2_X1 U595 ( .A1(G52), .A2(n655), .ZN(n545) );
  XOR2_X1 U596 ( .A(KEYINPUT70), .B(n545), .Z(n555) );
  INV_X1 U597 ( .A(G651), .ZN(n549) );
  NOR2_X1 U598 ( .A1(n650), .A2(n549), .ZN(n653) );
  NAND2_X1 U599 ( .A1(G77), .A2(n653), .ZN(n547) );
  NOR2_X1 U600 ( .A1(G651), .A2(G543), .ZN(n659) );
  NAND2_X1 U601 ( .A1(G90), .A2(n659), .ZN(n546) );
  NAND2_X1 U602 ( .A1(n547), .A2(n546), .ZN(n548) );
  XNOR2_X1 U603 ( .A(n548), .B(KEYINPUT9), .ZN(n553) );
  NOR2_X1 U604 ( .A1(G543), .A2(n549), .ZN(n550) );
  XOR2_X1 U605 ( .A(KEYINPUT68), .B(n550), .Z(n551) );
  XNOR2_X1 U606 ( .A(KEYINPUT1), .B(n551), .ZN(n656) );
  NAND2_X1 U607 ( .A1(G64), .A2(n656), .ZN(n552) );
  NAND2_X1 U608 ( .A1(n553), .A2(n552), .ZN(n554) );
  NOR2_X1 U609 ( .A1(n555), .A2(n554), .ZN(G171) );
  INV_X1 U610 ( .A(G171), .ZN(G301) );
  AND2_X1 U611 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U612 ( .A(G57), .ZN(G237) );
  NAND2_X1 U613 ( .A1(G75), .A2(n653), .ZN(n557) );
  NAND2_X1 U614 ( .A1(G88), .A2(n659), .ZN(n556) );
  NAND2_X1 U615 ( .A1(n557), .A2(n556), .ZN(n558) );
  XOR2_X1 U616 ( .A(KEYINPUT82), .B(n558), .Z(n562) );
  NAND2_X1 U617 ( .A1(n656), .A2(G62), .ZN(n560) );
  NAND2_X1 U618 ( .A1(n655), .A2(G50), .ZN(n559) );
  AND2_X1 U619 ( .A1(n560), .A2(n559), .ZN(n561) );
  NAND2_X1 U620 ( .A1(n562), .A2(n561), .ZN(G303) );
  NAND2_X1 U621 ( .A1(n659), .A2(G89), .ZN(n563) );
  XNOR2_X1 U622 ( .A(n563), .B(KEYINPUT4), .ZN(n565) );
  NAND2_X1 U623 ( .A1(G76), .A2(n653), .ZN(n564) );
  NAND2_X1 U624 ( .A1(n565), .A2(n564), .ZN(n566) );
  XNOR2_X1 U625 ( .A(KEYINPUT5), .B(n566), .ZN(n572) );
  NAND2_X1 U626 ( .A1(G63), .A2(n656), .ZN(n567) );
  XOR2_X1 U627 ( .A(KEYINPUT75), .B(n567), .Z(n569) );
  NAND2_X1 U628 ( .A1(n655), .A2(G51), .ZN(n568) );
  NAND2_X1 U629 ( .A1(n569), .A2(n568), .ZN(n570) );
  XOR2_X1 U630 ( .A(KEYINPUT6), .B(n570), .Z(n571) );
  NAND2_X1 U631 ( .A1(n572), .A2(n571), .ZN(n573) );
  XNOR2_X1 U632 ( .A(KEYINPUT7), .B(n573), .ZN(G168) );
  XOR2_X1 U633 ( .A(G168), .B(KEYINPUT8), .Z(n574) );
  XNOR2_X1 U634 ( .A(KEYINPUT76), .B(n574), .ZN(G286) );
  NAND2_X1 U635 ( .A1(G126), .A2(n887), .ZN(n576) );
  NAND2_X1 U636 ( .A1(G138), .A2(n891), .ZN(n575) );
  NAND2_X1 U637 ( .A1(n576), .A2(n575), .ZN(n580) );
  NAND2_X1 U638 ( .A1(G114), .A2(n888), .ZN(n578) );
  NAND2_X1 U639 ( .A1(G102), .A2(n892), .ZN(n577) );
  NAND2_X1 U640 ( .A1(n578), .A2(n577), .ZN(n579) );
  NOR2_X1 U641 ( .A1(n580), .A2(n579), .ZN(G164) );
  NAND2_X1 U642 ( .A1(G7), .A2(G661), .ZN(n581) );
  XOR2_X1 U643 ( .A(n581), .B(KEYINPUT10), .Z(n837) );
  NAND2_X1 U644 ( .A1(n837), .A2(G567), .ZN(n582) );
  XNOR2_X1 U645 ( .A(n582), .B(KEYINPUT11), .ZN(n583) );
  XNOR2_X1 U646 ( .A(KEYINPUT71), .B(n583), .ZN(G234) );
  NAND2_X1 U647 ( .A1(G81), .A2(n659), .ZN(n584) );
  XNOR2_X1 U648 ( .A(n584), .B(KEYINPUT12), .ZN(n585) );
  XNOR2_X1 U649 ( .A(n585), .B(KEYINPUT72), .ZN(n587) );
  NAND2_X1 U650 ( .A1(G68), .A2(n653), .ZN(n586) );
  NAND2_X1 U651 ( .A1(n587), .A2(n586), .ZN(n588) );
  XNOR2_X1 U652 ( .A(KEYINPUT13), .B(n588), .ZN(n594) );
  NAND2_X1 U653 ( .A1(n656), .A2(G56), .ZN(n589) );
  XOR2_X1 U654 ( .A(KEYINPUT14), .B(n589), .Z(n592) );
  NAND2_X1 U655 ( .A1(G43), .A2(n655), .ZN(n590) );
  XNOR2_X1 U656 ( .A(KEYINPUT73), .B(n590), .ZN(n591) );
  NOR2_X1 U657 ( .A1(n592), .A2(n591), .ZN(n593) );
  NAND2_X1 U658 ( .A1(n594), .A2(n593), .ZN(n704) );
  INV_X1 U659 ( .A(n704), .ZN(n921) );
  NAND2_X1 U660 ( .A1(n921), .A2(G860), .ZN(G153) );
  NAND2_X1 U661 ( .A1(G868), .A2(G301), .ZN(n604) );
  NAND2_X1 U662 ( .A1(G54), .A2(n655), .ZN(n601) );
  NAND2_X1 U663 ( .A1(G92), .A2(n659), .ZN(n596) );
  NAND2_X1 U664 ( .A1(G66), .A2(n656), .ZN(n595) );
  NAND2_X1 U665 ( .A1(n596), .A2(n595), .ZN(n599) );
  NAND2_X1 U666 ( .A1(n653), .A2(G79), .ZN(n597) );
  XOR2_X1 U667 ( .A(KEYINPUT74), .B(n597), .Z(n598) );
  NOR2_X1 U668 ( .A1(n599), .A2(n598), .ZN(n600) );
  NAND2_X1 U669 ( .A1(n601), .A2(n600), .ZN(n602) );
  XNOR2_X1 U670 ( .A(n602), .B(KEYINPUT15), .ZN(n920) );
  OR2_X1 U671 ( .A1(n920), .A2(G868), .ZN(n603) );
  NAND2_X1 U672 ( .A1(n604), .A2(n603), .ZN(G284) );
  NAND2_X1 U673 ( .A1(G868), .A2(G286), .ZN(n612) );
  NAND2_X1 U674 ( .A1(n655), .A2(G53), .ZN(n606) );
  NAND2_X1 U675 ( .A1(G65), .A2(n656), .ZN(n605) );
  NAND2_X1 U676 ( .A1(n606), .A2(n605), .ZN(n610) );
  NAND2_X1 U677 ( .A1(G78), .A2(n653), .ZN(n608) );
  NAND2_X1 U678 ( .A1(G91), .A2(n659), .ZN(n607) );
  NAND2_X1 U679 ( .A1(n608), .A2(n607), .ZN(n609) );
  NOR2_X1 U680 ( .A1(n610), .A2(n609), .ZN(n721) );
  OR2_X1 U681 ( .A1(n721), .A2(G868), .ZN(n611) );
  NAND2_X1 U682 ( .A1(n612), .A2(n611), .ZN(G297) );
  INV_X1 U683 ( .A(n721), .ZN(G299) );
  INV_X1 U684 ( .A(G559), .ZN(n613) );
  NOR2_X1 U685 ( .A1(G860), .A2(n613), .ZN(n614) );
  XNOR2_X1 U686 ( .A(KEYINPUT77), .B(n614), .ZN(n615) );
  NAND2_X1 U687 ( .A1(n615), .A2(n920), .ZN(n616) );
  XNOR2_X1 U688 ( .A(n616), .B(KEYINPUT16), .ZN(n617) );
  XNOR2_X1 U689 ( .A(KEYINPUT78), .B(n617), .ZN(G148) );
  NOR2_X1 U690 ( .A1(G868), .A2(n704), .ZN(n620) );
  NAND2_X1 U691 ( .A1(n920), .A2(G868), .ZN(n618) );
  NOR2_X1 U692 ( .A1(G559), .A2(n618), .ZN(n619) );
  NOR2_X1 U693 ( .A1(n620), .A2(n619), .ZN(G282) );
  NAND2_X1 U694 ( .A1(G111), .A2(n888), .ZN(n622) );
  NAND2_X1 U695 ( .A1(G99), .A2(n892), .ZN(n621) );
  NAND2_X1 U696 ( .A1(n622), .A2(n621), .ZN(n628) );
  NAND2_X1 U697 ( .A1(n887), .A2(G123), .ZN(n623) );
  XNOR2_X1 U698 ( .A(n623), .B(KEYINPUT18), .ZN(n625) );
  NAND2_X1 U699 ( .A1(G135), .A2(n891), .ZN(n624) );
  NAND2_X1 U700 ( .A1(n625), .A2(n624), .ZN(n626) );
  XOR2_X1 U701 ( .A(KEYINPUT79), .B(n626), .Z(n627) );
  NOR2_X1 U702 ( .A1(n628), .A2(n627), .ZN(n953) );
  XNOR2_X1 U703 ( .A(n953), .B(G2096), .ZN(n629) );
  INV_X1 U704 ( .A(G2100), .ZN(n860) );
  NAND2_X1 U705 ( .A1(n629), .A2(n860), .ZN(G156) );
  NAND2_X1 U706 ( .A1(n920), .A2(G559), .ZN(n674) );
  XOR2_X1 U707 ( .A(n921), .B(n674), .Z(n630) );
  NOR2_X1 U708 ( .A1(n630), .A2(G860), .ZN(n637) );
  NAND2_X1 U709 ( .A1(n655), .A2(G55), .ZN(n632) );
  NAND2_X1 U710 ( .A1(G67), .A2(n656), .ZN(n631) );
  NAND2_X1 U711 ( .A1(n632), .A2(n631), .ZN(n636) );
  NAND2_X1 U712 ( .A1(G80), .A2(n653), .ZN(n634) );
  NAND2_X1 U713 ( .A1(G93), .A2(n659), .ZN(n633) );
  NAND2_X1 U714 ( .A1(n634), .A2(n633), .ZN(n635) );
  NOR2_X1 U715 ( .A1(n636), .A2(n635), .ZN(n671) );
  XNOR2_X1 U716 ( .A(n637), .B(n671), .ZN(G145) );
  NAND2_X1 U717 ( .A1(G85), .A2(n659), .ZN(n639) );
  NAND2_X1 U718 ( .A1(G60), .A2(n656), .ZN(n638) );
  NAND2_X1 U719 ( .A1(n639), .A2(n638), .ZN(n642) );
  NAND2_X1 U720 ( .A1(G72), .A2(n653), .ZN(n640) );
  XNOR2_X1 U721 ( .A(KEYINPUT67), .B(n640), .ZN(n641) );
  NOR2_X1 U722 ( .A1(n642), .A2(n641), .ZN(n644) );
  NAND2_X1 U723 ( .A1(n655), .A2(G47), .ZN(n643) );
  NAND2_X1 U724 ( .A1(n644), .A2(n643), .ZN(n645) );
  XOR2_X1 U725 ( .A(KEYINPUT69), .B(n645), .Z(G290) );
  NAND2_X1 U726 ( .A1(G49), .A2(n655), .ZN(n647) );
  NAND2_X1 U727 ( .A1(G74), .A2(G651), .ZN(n646) );
  NAND2_X1 U728 ( .A1(n647), .A2(n646), .ZN(n648) );
  NOR2_X1 U729 ( .A1(n656), .A2(n648), .ZN(n649) );
  XNOR2_X1 U730 ( .A(n649), .B(KEYINPUT80), .ZN(n652) );
  NAND2_X1 U731 ( .A1(G87), .A2(n650), .ZN(n651) );
  NAND2_X1 U732 ( .A1(n652), .A2(n651), .ZN(G288) );
  NAND2_X1 U733 ( .A1(G73), .A2(n653), .ZN(n654) );
  XNOR2_X1 U734 ( .A(n654), .B(KEYINPUT2), .ZN(n664) );
  NAND2_X1 U735 ( .A1(n655), .A2(G48), .ZN(n658) );
  NAND2_X1 U736 ( .A1(G61), .A2(n656), .ZN(n657) );
  NAND2_X1 U737 ( .A1(n658), .A2(n657), .ZN(n662) );
  NAND2_X1 U738 ( .A1(G86), .A2(n659), .ZN(n660) );
  XNOR2_X1 U739 ( .A(KEYINPUT81), .B(n660), .ZN(n661) );
  NOR2_X1 U740 ( .A1(n662), .A2(n661), .ZN(n663) );
  NAND2_X1 U741 ( .A1(n664), .A2(n663), .ZN(G305) );
  NOR2_X1 U742 ( .A1(G868), .A2(n671), .ZN(n665) );
  XOR2_X1 U743 ( .A(n665), .B(KEYINPUT84), .Z(n677) );
  XNOR2_X1 U744 ( .A(KEYINPUT83), .B(KEYINPUT19), .ZN(n667) );
  XOR2_X1 U745 ( .A(G290), .B(G299), .Z(n666) );
  XNOR2_X1 U746 ( .A(n667), .B(n666), .ZN(n670) );
  XOR2_X1 U747 ( .A(G303), .B(n704), .Z(n668) );
  XNOR2_X1 U748 ( .A(n668), .B(G288), .ZN(n669) );
  XNOR2_X1 U749 ( .A(n670), .B(n669), .ZN(n673) );
  XNOR2_X1 U750 ( .A(G305), .B(n671), .ZN(n672) );
  XNOR2_X1 U751 ( .A(n673), .B(n672), .ZN(n910) );
  XOR2_X1 U752 ( .A(n910), .B(n674), .Z(n675) );
  NAND2_X1 U753 ( .A1(G868), .A2(n675), .ZN(n676) );
  NAND2_X1 U754 ( .A1(n677), .A2(n676), .ZN(G295) );
  NAND2_X1 U755 ( .A1(G2084), .A2(G2078), .ZN(n678) );
  XNOR2_X1 U756 ( .A(n678), .B(KEYINPUT20), .ZN(n679) );
  XNOR2_X1 U757 ( .A(KEYINPUT85), .B(n679), .ZN(n680) );
  NAND2_X1 U758 ( .A1(n680), .A2(G2090), .ZN(n681) );
  XNOR2_X1 U759 ( .A(n681), .B(KEYINPUT86), .ZN(n682) );
  XNOR2_X1 U760 ( .A(KEYINPUT21), .B(n682), .ZN(n683) );
  NAND2_X1 U761 ( .A1(n683), .A2(G2072), .ZN(n684) );
  XOR2_X1 U762 ( .A(KEYINPUT87), .B(n684), .Z(G158) );
  XNOR2_X1 U763 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  XOR2_X1 U764 ( .A(KEYINPUT88), .B(KEYINPUT22), .Z(n686) );
  NAND2_X1 U765 ( .A1(G132), .A2(G82), .ZN(n685) );
  XNOR2_X1 U766 ( .A(n686), .B(n685), .ZN(n687) );
  NAND2_X1 U767 ( .A1(n687), .A2(G96), .ZN(n688) );
  NOR2_X1 U768 ( .A1(n688), .A2(G218), .ZN(n689) );
  XNOR2_X1 U769 ( .A(n689), .B(KEYINPUT89), .ZN(n845) );
  NAND2_X1 U770 ( .A1(n845), .A2(G2106), .ZN(n693) );
  NAND2_X1 U771 ( .A1(G120), .A2(G69), .ZN(n690) );
  NOR2_X1 U772 ( .A1(G237), .A2(n690), .ZN(n691) );
  NAND2_X1 U773 ( .A1(G108), .A2(n691), .ZN(n844) );
  NAND2_X1 U774 ( .A1(n844), .A2(G567), .ZN(n692) );
  NAND2_X1 U775 ( .A1(n693), .A2(n692), .ZN(n847) );
  NAND2_X1 U776 ( .A1(G483), .A2(G661), .ZN(n694) );
  NOR2_X1 U777 ( .A1(n847), .A2(n694), .ZN(n841) );
  NAND2_X1 U778 ( .A1(n841), .A2(G36), .ZN(G176) );
  NAND2_X1 U779 ( .A1(G40), .A2(G160), .ZN(n762) );
  XNOR2_X1 U780 ( .A(KEYINPUT93), .B(n762), .ZN(n698) );
  NOR2_X1 U781 ( .A1(G164), .A2(G1384), .ZN(n763) );
  XOR2_X1 U782 ( .A(G2078), .B(KEYINPUT25), .Z(n695) );
  XNOR2_X1 U783 ( .A(KEYINPUT95), .B(n695), .ZN(n981) );
  NOR2_X1 U784 ( .A1(n740), .A2(n981), .ZN(n697) );
  AND2_X1 U785 ( .A1(n740), .A2(G1961), .ZN(n696) );
  NOR2_X1 U786 ( .A1(n697), .A2(n696), .ZN(n735) );
  NAND2_X1 U787 ( .A1(G171), .A2(n735), .ZN(n729) );
  INV_X1 U788 ( .A(KEYINPUT97), .ZN(n703) );
  NAND2_X1 U789 ( .A1(n714), .A2(G1996), .ZN(n699) );
  XNOR2_X1 U790 ( .A(n699), .B(KEYINPUT26), .ZN(n701) );
  NAND2_X1 U791 ( .A1(G1341), .A2(n740), .ZN(n700) );
  NAND2_X1 U792 ( .A1(n701), .A2(n700), .ZN(n702) );
  XNOR2_X1 U793 ( .A(n703), .B(n702), .ZN(n705) );
  NAND2_X1 U794 ( .A1(n920), .A2(n706), .ZN(n710) );
  NOR2_X1 U795 ( .A1(n714), .A2(G1348), .ZN(n708) );
  NOR2_X1 U796 ( .A1(G2067), .A2(n740), .ZN(n707) );
  NOR2_X1 U797 ( .A1(n708), .A2(n707), .ZN(n709) );
  NAND2_X1 U798 ( .A1(n710), .A2(n709), .ZN(n711) );
  NAND2_X1 U799 ( .A1(n712), .A2(n711), .ZN(n713) );
  XNOR2_X1 U800 ( .A(n713), .B(KEYINPUT98), .ZN(n720) );
  NAND2_X1 U801 ( .A1(n714), .A2(G2072), .ZN(n715) );
  XNOR2_X1 U802 ( .A(KEYINPUT27), .B(n715), .ZN(n718) );
  NAND2_X1 U803 ( .A1(G1956), .A2(n740), .ZN(n716) );
  XOR2_X1 U804 ( .A(KEYINPUT96), .B(n716), .Z(n717) );
  NOR2_X1 U805 ( .A1(n718), .A2(n717), .ZN(n722) );
  NAND2_X1 U806 ( .A1(n722), .A2(n721), .ZN(n719) );
  NAND2_X1 U807 ( .A1(n720), .A2(n719), .ZN(n725) );
  NOR2_X1 U808 ( .A1(n722), .A2(n721), .ZN(n723) );
  XOR2_X1 U809 ( .A(n723), .B(KEYINPUT28), .Z(n724) );
  NAND2_X1 U810 ( .A1(n725), .A2(n724), .ZN(n727) );
  NAND2_X1 U811 ( .A1(n729), .A2(n728), .ZN(n753) );
  INV_X1 U812 ( .A(KEYINPUT31), .ZN(n739) );
  NAND2_X1 U813 ( .A1(G8), .A2(n740), .ZN(n813) );
  NOR2_X1 U814 ( .A1(G1966), .A2(n813), .ZN(n755) );
  NOR2_X1 U815 ( .A1(G2084), .A2(n740), .ZN(n751) );
  NOR2_X1 U816 ( .A1(n755), .A2(n751), .ZN(n730) );
  NAND2_X1 U817 ( .A1(G8), .A2(n730), .ZN(n733) );
  INV_X1 U818 ( .A(KEYINPUT99), .ZN(n731) );
  NOR2_X1 U819 ( .A1(G168), .A2(n734), .ZN(n737) );
  NOR2_X1 U820 ( .A1(G171), .A2(n735), .ZN(n736) );
  XNOR2_X1 U821 ( .A(n739), .B(n738), .ZN(n752) );
  NOR2_X1 U822 ( .A1(G1971), .A2(n813), .ZN(n742) );
  NOR2_X1 U823 ( .A1(G2090), .A2(n740), .ZN(n741) );
  NOR2_X1 U824 ( .A1(n742), .A2(n741), .ZN(n743) );
  NAND2_X1 U825 ( .A1(n743), .A2(G303), .ZN(n745) );
  AND2_X1 U826 ( .A1(n752), .A2(n745), .ZN(n744) );
  NAND2_X1 U827 ( .A1(n753), .A2(n744), .ZN(n748) );
  INV_X1 U828 ( .A(n745), .ZN(n746) );
  OR2_X1 U829 ( .A1(n746), .A2(G286), .ZN(n747) );
  AND2_X1 U830 ( .A1(n748), .A2(n747), .ZN(n749) );
  NAND2_X1 U831 ( .A1(G8), .A2(n749), .ZN(n750) );
  XNOR2_X1 U832 ( .A(n750), .B(KEYINPUT32), .ZN(n759) );
  NAND2_X1 U833 ( .A1(G8), .A2(n751), .ZN(n757) );
  AND2_X1 U834 ( .A1(n753), .A2(n752), .ZN(n754) );
  NOR2_X1 U835 ( .A1(n755), .A2(n754), .ZN(n756) );
  NAND2_X1 U836 ( .A1(n757), .A2(n756), .ZN(n758) );
  NAND2_X1 U837 ( .A1(n759), .A2(n758), .ZN(n809) );
  NOR2_X1 U838 ( .A1(G2090), .A2(G303), .ZN(n760) );
  NAND2_X1 U839 ( .A1(G8), .A2(n760), .ZN(n761) );
  NAND2_X1 U840 ( .A1(n809), .A2(n761), .ZN(n793) );
  NOR2_X1 U841 ( .A1(n763), .A2(n762), .ZN(n831) );
  NAND2_X1 U842 ( .A1(G140), .A2(n891), .ZN(n765) );
  NAND2_X1 U843 ( .A1(G104), .A2(n892), .ZN(n764) );
  NAND2_X1 U844 ( .A1(n765), .A2(n764), .ZN(n766) );
  XNOR2_X1 U845 ( .A(KEYINPUT34), .B(n766), .ZN(n771) );
  NAND2_X1 U846 ( .A1(G128), .A2(n887), .ZN(n768) );
  NAND2_X1 U847 ( .A1(G116), .A2(n888), .ZN(n767) );
  NAND2_X1 U848 ( .A1(n768), .A2(n767), .ZN(n769) );
  XOR2_X1 U849 ( .A(KEYINPUT35), .B(n769), .Z(n770) );
  NOR2_X1 U850 ( .A1(n771), .A2(n770), .ZN(n772) );
  XNOR2_X1 U851 ( .A(KEYINPUT36), .B(n772), .ZN(n884) );
  XNOR2_X1 U852 ( .A(G2067), .B(KEYINPUT37), .ZN(n829) );
  NOR2_X1 U853 ( .A1(n884), .A2(n829), .ZN(n948) );
  NAND2_X1 U854 ( .A1(n831), .A2(n948), .ZN(n773) );
  XNOR2_X1 U855 ( .A(KEYINPUT90), .B(n773), .ZN(n827) );
  NAND2_X1 U856 ( .A1(G131), .A2(n891), .ZN(n774) );
  XNOR2_X1 U857 ( .A(n774), .B(KEYINPUT92), .ZN(n781) );
  NAND2_X1 U858 ( .A1(G119), .A2(n887), .ZN(n776) );
  NAND2_X1 U859 ( .A1(G95), .A2(n892), .ZN(n775) );
  NAND2_X1 U860 ( .A1(n776), .A2(n775), .ZN(n779) );
  NAND2_X1 U861 ( .A1(G107), .A2(n888), .ZN(n777) );
  XNOR2_X1 U862 ( .A(KEYINPUT91), .B(n777), .ZN(n778) );
  NOR2_X1 U863 ( .A1(n779), .A2(n778), .ZN(n780) );
  NAND2_X1 U864 ( .A1(n781), .A2(n780), .ZN(n900) );
  AND2_X1 U865 ( .A1(n900), .A2(G1991), .ZN(n790) );
  NAND2_X1 U866 ( .A1(G141), .A2(n891), .ZN(n783) );
  NAND2_X1 U867 ( .A1(G117), .A2(n888), .ZN(n782) );
  NAND2_X1 U868 ( .A1(n783), .A2(n782), .ZN(n786) );
  NAND2_X1 U869 ( .A1(n892), .A2(G105), .ZN(n784) );
  XOR2_X1 U870 ( .A(KEYINPUT38), .B(n784), .Z(n785) );
  NOR2_X1 U871 ( .A1(n786), .A2(n785), .ZN(n788) );
  NAND2_X1 U872 ( .A1(n887), .A2(G129), .ZN(n787) );
  NAND2_X1 U873 ( .A1(n788), .A2(n787), .ZN(n901) );
  AND2_X1 U874 ( .A1(G1996), .A2(n901), .ZN(n789) );
  NOR2_X1 U875 ( .A1(n790), .A2(n789), .ZN(n946) );
  INV_X1 U876 ( .A(n831), .ZN(n819) );
  NOR2_X1 U877 ( .A1(n946), .A2(n819), .ZN(n824) );
  INV_X1 U878 ( .A(n824), .ZN(n791) );
  AND2_X1 U879 ( .A1(n827), .A2(n791), .ZN(n801) );
  AND2_X1 U880 ( .A1(n813), .A2(n801), .ZN(n792) );
  AND2_X1 U881 ( .A1(n793), .A2(n792), .ZN(n806) );
  NOR2_X1 U882 ( .A1(G1981), .A2(G305), .ZN(n794) );
  XOR2_X1 U883 ( .A(n794), .B(KEYINPUT94), .Z(n795) );
  XNOR2_X1 U884 ( .A(KEYINPUT24), .B(n795), .ZN(n796) );
  NOR2_X1 U885 ( .A1(n813), .A2(n796), .ZN(n797) );
  NAND2_X1 U886 ( .A1(n801), .A2(n797), .ZN(n804) );
  NOR2_X1 U887 ( .A1(G1976), .A2(G288), .ZN(n808) );
  NAND2_X1 U888 ( .A1(n808), .A2(KEYINPUT33), .ZN(n798) );
  NOR2_X1 U889 ( .A1(n798), .A2(n813), .ZN(n800) );
  XOR2_X1 U890 ( .A(G1981), .B(G305), .Z(n924) );
  INV_X1 U891 ( .A(n924), .ZN(n799) );
  NOR2_X1 U892 ( .A1(n800), .A2(n799), .ZN(n802) );
  AND2_X1 U893 ( .A1(n802), .A2(n801), .ZN(n814) );
  NAND2_X1 U894 ( .A1(n814), .A2(KEYINPUT33), .ZN(n803) );
  NAND2_X1 U895 ( .A1(n804), .A2(n803), .ZN(n805) );
  NOR2_X1 U896 ( .A1(n806), .A2(n805), .ZN(n818) );
  NOR2_X1 U897 ( .A1(G1971), .A2(G303), .ZN(n807) );
  NOR2_X1 U898 ( .A1(n808), .A2(n807), .ZN(n927) );
  NAND2_X1 U899 ( .A1(n809), .A2(n927), .ZN(n810) );
  XNOR2_X1 U900 ( .A(n810), .B(KEYINPUT100), .ZN(n816) );
  NAND2_X1 U901 ( .A1(G288), .A2(G1976), .ZN(n811) );
  XOR2_X1 U902 ( .A(KEYINPUT101), .B(n811), .Z(n934) );
  INV_X1 U903 ( .A(n934), .ZN(n812) );
  AND2_X1 U904 ( .A1(n523), .A2(n814), .ZN(n815) );
  NAND2_X1 U905 ( .A1(n816), .A2(n815), .ZN(n817) );
  NAND2_X1 U906 ( .A1(n818), .A2(n817), .ZN(n821) );
  XOR2_X1 U907 ( .A(G1986), .B(G290), .Z(n928) );
  OR2_X1 U908 ( .A1(n928), .A2(n819), .ZN(n820) );
  NAND2_X1 U909 ( .A1(n821), .A2(n820), .ZN(n834) );
  NOR2_X1 U910 ( .A1(G1996), .A2(n901), .ZN(n951) );
  NOR2_X1 U911 ( .A1(G1986), .A2(G290), .ZN(n822) );
  NOR2_X1 U912 ( .A1(G1991), .A2(n900), .ZN(n954) );
  NOR2_X1 U913 ( .A1(n822), .A2(n954), .ZN(n823) );
  NOR2_X1 U914 ( .A1(n824), .A2(n823), .ZN(n825) );
  NOR2_X1 U915 ( .A1(n951), .A2(n825), .ZN(n826) );
  XNOR2_X1 U916 ( .A(n826), .B(KEYINPUT39), .ZN(n828) );
  NAND2_X1 U917 ( .A1(n828), .A2(n827), .ZN(n830) );
  NAND2_X1 U918 ( .A1(n884), .A2(n829), .ZN(n945) );
  NAND2_X1 U919 ( .A1(n830), .A2(n945), .ZN(n832) );
  NAND2_X1 U920 ( .A1(n832), .A2(n831), .ZN(n833) );
  NAND2_X1 U921 ( .A1(n834), .A2(n833), .ZN(n835) );
  XNOR2_X1 U922 ( .A(KEYINPUT40), .B(n835), .ZN(G329) );
  NAND2_X1 U923 ( .A1(n837), .A2(G2106), .ZN(n836) );
  XNOR2_X1 U924 ( .A(n836), .B(KEYINPUT102), .ZN(G217) );
  INV_X1 U925 ( .A(n837), .ZN(G223) );
  NAND2_X1 U926 ( .A1(G15), .A2(G2), .ZN(n839) );
  INV_X1 U927 ( .A(G661), .ZN(n838) );
  NOR2_X1 U928 ( .A1(n839), .A2(n838), .ZN(n840) );
  XNOR2_X1 U929 ( .A(n840), .B(KEYINPUT103), .ZN(G259) );
  NAND2_X1 U930 ( .A1(G1), .A2(G3), .ZN(n842) );
  NAND2_X1 U931 ( .A1(n842), .A2(n841), .ZN(n843) );
  XNOR2_X1 U932 ( .A(n843), .B(KEYINPUT104), .ZN(G188) );
  XNOR2_X1 U933 ( .A(G69), .B(KEYINPUT105), .ZN(G235) );
  INV_X1 U935 ( .A(G132), .ZN(G219) );
  INV_X1 U936 ( .A(G120), .ZN(G236) );
  INV_X1 U937 ( .A(G96), .ZN(G221) );
  INV_X1 U938 ( .A(G82), .ZN(G220) );
  NOR2_X1 U939 ( .A1(n845), .A2(n844), .ZN(n846) );
  XOR2_X1 U940 ( .A(n846), .B(KEYINPUT106), .Z(G261) );
  INV_X1 U941 ( .A(G261), .ZN(G325) );
  INV_X1 U942 ( .A(n847), .ZN(G319) );
  XNOR2_X1 U943 ( .A(G1961), .B(KEYINPUT41), .ZN(n857) );
  XOR2_X1 U944 ( .A(G1976), .B(G1981), .Z(n849) );
  XNOR2_X1 U945 ( .A(G1966), .B(G1956), .ZN(n848) );
  XNOR2_X1 U946 ( .A(n849), .B(n848), .ZN(n853) );
  XOR2_X1 U947 ( .A(G1971), .B(G1986), .Z(n851) );
  XNOR2_X1 U948 ( .A(G1996), .B(G1991), .ZN(n850) );
  XNOR2_X1 U949 ( .A(n851), .B(n850), .ZN(n852) );
  XOR2_X1 U950 ( .A(n853), .B(n852), .Z(n855) );
  XNOR2_X1 U951 ( .A(KEYINPUT108), .B(G2474), .ZN(n854) );
  XNOR2_X1 U952 ( .A(n855), .B(n854), .ZN(n856) );
  XNOR2_X1 U953 ( .A(n857), .B(n856), .ZN(G229) );
  XOR2_X1 U954 ( .A(G2678), .B(G2084), .Z(n859) );
  XNOR2_X1 U955 ( .A(G2067), .B(G2072), .ZN(n858) );
  XNOR2_X1 U956 ( .A(n859), .B(n858), .ZN(n861) );
  XNOR2_X1 U957 ( .A(n861), .B(n860), .ZN(n863) );
  XNOR2_X1 U958 ( .A(G2078), .B(G2090), .ZN(n862) );
  XNOR2_X1 U959 ( .A(n863), .B(n862), .ZN(n867) );
  XOR2_X1 U960 ( .A(G2096), .B(KEYINPUT107), .Z(n865) );
  XNOR2_X1 U961 ( .A(KEYINPUT42), .B(KEYINPUT43), .ZN(n864) );
  XNOR2_X1 U962 ( .A(n865), .B(n864), .ZN(n866) );
  XOR2_X1 U963 ( .A(n867), .B(n866), .Z(G227) );
  NAND2_X1 U964 ( .A1(G124), .A2(n887), .ZN(n868) );
  XNOR2_X1 U965 ( .A(n868), .B(KEYINPUT44), .ZN(n871) );
  NAND2_X1 U966 ( .A1(G100), .A2(n892), .ZN(n869) );
  XOR2_X1 U967 ( .A(KEYINPUT109), .B(n869), .Z(n870) );
  NAND2_X1 U968 ( .A1(n871), .A2(n870), .ZN(n875) );
  NAND2_X1 U969 ( .A1(G136), .A2(n891), .ZN(n873) );
  NAND2_X1 U970 ( .A1(G112), .A2(n888), .ZN(n872) );
  NAND2_X1 U971 ( .A1(n873), .A2(n872), .ZN(n874) );
  NOR2_X1 U972 ( .A1(n875), .A2(n874), .ZN(G162) );
  XNOR2_X1 U973 ( .A(KEYINPUT46), .B(KEYINPUT48), .ZN(n886) );
  NAND2_X1 U974 ( .A1(G139), .A2(n891), .ZN(n877) );
  NAND2_X1 U975 ( .A1(G103), .A2(n892), .ZN(n876) );
  NAND2_X1 U976 ( .A1(n877), .A2(n876), .ZN(n878) );
  XOR2_X1 U977 ( .A(KEYINPUT111), .B(n878), .Z(n883) );
  NAND2_X1 U978 ( .A1(G127), .A2(n887), .ZN(n880) );
  NAND2_X1 U979 ( .A1(G115), .A2(n888), .ZN(n879) );
  NAND2_X1 U980 ( .A1(n880), .A2(n879), .ZN(n881) );
  XOR2_X1 U981 ( .A(KEYINPUT47), .B(n881), .Z(n882) );
  NOR2_X1 U982 ( .A1(n883), .A2(n882), .ZN(n963) );
  XNOR2_X1 U983 ( .A(n884), .B(n963), .ZN(n885) );
  XNOR2_X1 U984 ( .A(n886), .B(n885), .ZN(n905) );
  NAND2_X1 U985 ( .A1(G130), .A2(n887), .ZN(n890) );
  NAND2_X1 U986 ( .A1(G118), .A2(n888), .ZN(n889) );
  NAND2_X1 U987 ( .A1(n890), .A2(n889), .ZN(n898) );
  NAND2_X1 U988 ( .A1(G142), .A2(n891), .ZN(n894) );
  NAND2_X1 U989 ( .A1(G106), .A2(n892), .ZN(n893) );
  NAND2_X1 U990 ( .A1(n894), .A2(n893), .ZN(n895) );
  XOR2_X1 U991 ( .A(KEYINPUT45), .B(n895), .Z(n896) );
  XNOR2_X1 U992 ( .A(KEYINPUT110), .B(n896), .ZN(n897) );
  NOR2_X1 U993 ( .A1(n898), .A2(n897), .ZN(n899) );
  XOR2_X1 U994 ( .A(n899), .B(G162), .Z(n903) );
  XNOR2_X1 U995 ( .A(n901), .B(n900), .ZN(n902) );
  XNOR2_X1 U996 ( .A(n903), .B(n902), .ZN(n904) );
  XOR2_X1 U997 ( .A(n905), .B(n904), .Z(n907) );
  XNOR2_X1 U998 ( .A(G164), .B(n953), .ZN(n906) );
  XNOR2_X1 U999 ( .A(n907), .B(n906), .ZN(n908) );
  XNOR2_X1 U1000 ( .A(n908), .B(G160), .ZN(n909) );
  NOR2_X1 U1001 ( .A1(G37), .A2(n909), .ZN(G395) );
  XNOR2_X1 U1002 ( .A(G286), .B(n910), .ZN(n912) );
  XOR2_X1 U1003 ( .A(G301), .B(n920), .Z(n911) );
  XNOR2_X1 U1004 ( .A(n912), .B(n911), .ZN(n913) );
  NOR2_X1 U1005 ( .A1(G37), .A2(n913), .ZN(G397) );
  NOR2_X1 U1006 ( .A1(G229), .A2(G227), .ZN(n914) );
  XOR2_X1 U1007 ( .A(KEYINPUT49), .B(n914), .Z(n915) );
  NAND2_X1 U1008 ( .A1(G319), .A2(n915), .ZN(n916) );
  NOR2_X1 U1009 ( .A1(G401), .A2(n916), .ZN(n917) );
  XNOR2_X1 U1010 ( .A(KEYINPUT112), .B(n917), .ZN(n919) );
  NOR2_X1 U1011 ( .A1(G395), .A2(G397), .ZN(n918) );
  NAND2_X1 U1012 ( .A1(n919), .A2(n918), .ZN(G225) );
  INV_X1 U1013 ( .A(G225), .ZN(G308) );
  INV_X1 U1014 ( .A(G303), .ZN(G166) );
  INV_X1 U1015 ( .A(G108), .ZN(G238) );
  INV_X1 U1016 ( .A(G16), .ZN(n942) );
  XNOR2_X1 U1017 ( .A(n920), .B(G1348), .ZN(n923) );
  XNOR2_X1 U1018 ( .A(G1341), .B(n921), .ZN(n922) );
  NAND2_X1 U1019 ( .A1(n923), .A2(n922), .ZN(n941) );
  XNOR2_X1 U1020 ( .A(G1966), .B(G168), .ZN(n925) );
  NAND2_X1 U1021 ( .A1(n925), .A2(n924), .ZN(n926) );
  XNOR2_X1 U1022 ( .A(n926), .B(KEYINPUT57), .ZN(n939) );
  NAND2_X1 U1023 ( .A1(n928), .A2(n927), .ZN(n937) );
  XOR2_X1 U1024 ( .A(G301), .B(G1961), .Z(n929) );
  XNOR2_X1 U1025 ( .A(n929), .B(KEYINPUT123), .ZN(n933) );
  XOR2_X1 U1026 ( .A(G299), .B(G1956), .Z(n931) );
  NAND2_X1 U1027 ( .A1(G1971), .A2(G303), .ZN(n930) );
  NAND2_X1 U1028 ( .A1(n931), .A2(n930), .ZN(n932) );
  NOR2_X1 U1029 ( .A1(n933), .A2(n932), .ZN(n935) );
  NAND2_X1 U1030 ( .A1(n935), .A2(n934), .ZN(n936) );
  NOR2_X1 U1031 ( .A1(n937), .A2(n936), .ZN(n938) );
  NAND2_X1 U1032 ( .A1(n939), .A2(n938), .ZN(n940) );
  NOR2_X1 U1033 ( .A1(n941), .A2(n940), .ZN(n1024) );
  NOR2_X1 U1034 ( .A1(n942), .A2(n1024), .ZN(n943) );
  NAND2_X1 U1035 ( .A1(KEYINPUT56), .A2(n943), .ZN(n944) );
  NAND2_X1 U1036 ( .A1(G11), .A2(n944), .ZN(n975) );
  NAND2_X1 U1037 ( .A1(n946), .A2(n945), .ZN(n947) );
  NOR2_X1 U1038 ( .A1(n948), .A2(n947), .ZN(n962) );
  XNOR2_X1 U1039 ( .A(G2090), .B(G162), .ZN(n949) );
  XNOR2_X1 U1040 ( .A(n949), .B(KEYINPUT115), .ZN(n950) );
  NOR2_X1 U1041 ( .A1(n951), .A2(n950), .ZN(n952) );
  XOR2_X1 U1042 ( .A(KEYINPUT51), .B(n952), .Z(n957) );
  NOR2_X1 U1043 ( .A1(n954), .A2(n953), .ZN(n955) );
  XNOR2_X1 U1044 ( .A(KEYINPUT114), .B(n955), .ZN(n956) );
  NAND2_X1 U1045 ( .A1(n957), .A2(n956), .ZN(n960) );
  XNOR2_X1 U1046 ( .A(G2084), .B(G160), .ZN(n958) );
  XNOR2_X1 U1047 ( .A(KEYINPUT113), .B(n958), .ZN(n959) );
  NOR2_X1 U1048 ( .A1(n960), .A2(n959), .ZN(n961) );
  NAND2_X1 U1049 ( .A1(n962), .A2(n961), .ZN(n968) );
  XOR2_X1 U1050 ( .A(G2072), .B(n963), .Z(n965) );
  XOR2_X1 U1051 ( .A(G164), .B(G2078), .Z(n964) );
  NOR2_X1 U1052 ( .A1(n965), .A2(n964), .ZN(n966) );
  XOR2_X1 U1053 ( .A(KEYINPUT50), .B(n966), .Z(n967) );
  NOR2_X1 U1054 ( .A1(n968), .A2(n967), .ZN(n969) );
  XNOR2_X1 U1055 ( .A(KEYINPUT52), .B(n969), .ZN(n970) );
  XNOR2_X1 U1056 ( .A(n970), .B(KEYINPUT116), .ZN(n971) );
  INV_X1 U1057 ( .A(KEYINPUT55), .ZN(n998) );
  NAND2_X1 U1058 ( .A1(n971), .A2(n998), .ZN(n972) );
  NAND2_X1 U1059 ( .A1(G29), .A2(n972), .ZN(n973) );
  XNOR2_X1 U1060 ( .A(KEYINPUT117), .B(n973), .ZN(n974) );
  NOR2_X1 U1061 ( .A1(n975), .A2(n974), .ZN(n1031) );
  XNOR2_X1 U1062 ( .A(G2084), .B(KEYINPUT54), .ZN(n976) );
  XNOR2_X1 U1063 ( .A(n976), .B(G34), .ZN(n996) );
  XNOR2_X1 U1064 ( .A(G2090), .B(G35), .ZN(n993) );
  XNOR2_X1 U1065 ( .A(G2072), .B(G33), .ZN(n977) );
  XNOR2_X1 U1066 ( .A(n977), .B(KEYINPUT118), .ZN(n979) );
  XNOR2_X1 U1067 ( .A(G26), .B(G2067), .ZN(n978) );
  NOR2_X1 U1068 ( .A1(n979), .A2(n978), .ZN(n980) );
  XOR2_X1 U1069 ( .A(KEYINPUT119), .B(n980), .Z(n986) );
  XOR2_X1 U1070 ( .A(n981), .B(G27), .Z(n983) );
  XNOR2_X1 U1071 ( .A(G1996), .B(G32), .ZN(n982) );
  NOR2_X1 U1072 ( .A1(n983), .A2(n982), .ZN(n984) );
  XNOR2_X1 U1073 ( .A(KEYINPUT120), .B(n984), .ZN(n985) );
  NAND2_X1 U1074 ( .A1(n986), .A2(n985), .ZN(n987) );
  XNOR2_X1 U1075 ( .A(KEYINPUT121), .B(n987), .ZN(n988) );
  NAND2_X1 U1076 ( .A1(n988), .A2(G28), .ZN(n990) );
  XNOR2_X1 U1077 ( .A(G25), .B(G1991), .ZN(n989) );
  NOR2_X1 U1078 ( .A1(n990), .A2(n989), .ZN(n991) );
  XNOR2_X1 U1079 ( .A(KEYINPUT53), .B(n991), .ZN(n992) );
  NOR2_X1 U1080 ( .A1(n993), .A2(n992), .ZN(n994) );
  XOR2_X1 U1081 ( .A(KEYINPUT122), .B(n994), .Z(n995) );
  NOR2_X1 U1082 ( .A1(n996), .A2(n995), .ZN(n997) );
  XNOR2_X1 U1083 ( .A(n998), .B(n997), .ZN(n999) );
  NOR2_X1 U1084 ( .A1(G29), .A2(n999), .ZN(n1029) );
  XNOR2_X1 U1085 ( .A(G1971), .B(G22), .ZN(n1001) );
  XNOR2_X1 U1086 ( .A(G23), .B(G1976), .ZN(n1000) );
  NOR2_X1 U1087 ( .A1(n1001), .A2(n1000), .ZN(n1002) );
  XOR2_X1 U1088 ( .A(KEYINPUT126), .B(n1002), .Z(n1004) );
  XNOR2_X1 U1089 ( .A(G1986), .B(G24), .ZN(n1003) );
  NOR2_X1 U1090 ( .A1(n1004), .A2(n1003), .ZN(n1005) );
  XNOR2_X1 U1091 ( .A(n1005), .B(KEYINPUT58), .ZN(n1006) );
  XNOR2_X1 U1092 ( .A(n1006), .B(KEYINPUT127), .ZN(n1022) );
  XOR2_X1 U1093 ( .A(G1966), .B(G21), .Z(n1017) );
  XOR2_X1 U1094 ( .A(G1348), .B(KEYINPUT59), .Z(n1007) );
  XNOR2_X1 U1095 ( .A(G4), .B(n1007), .ZN(n1009) );
  XNOR2_X1 U1096 ( .A(G6), .B(G1981), .ZN(n1008) );
  NOR2_X1 U1097 ( .A1(n1009), .A2(n1008), .ZN(n1013) );
  XNOR2_X1 U1098 ( .A(G1956), .B(G20), .ZN(n1011) );
  XNOR2_X1 U1099 ( .A(G19), .B(G1341), .ZN(n1010) );
  NOR2_X1 U1100 ( .A1(n1011), .A2(n1010), .ZN(n1012) );
  NAND2_X1 U1101 ( .A1(n1013), .A2(n1012), .ZN(n1014) );
  XOR2_X1 U1102 ( .A(KEYINPUT124), .B(n1014), .Z(n1015) );
  XNOR2_X1 U1103 ( .A(n1015), .B(KEYINPUT60), .ZN(n1016) );
  NAND2_X1 U1104 ( .A1(n1017), .A2(n1016), .ZN(n1019) );
  XNOR2_X1 U1105 ( .A(G5), .B(G1961), .ZN(n1018) );
  NOR2_X1 U1106 ( .A1(n1019), .A2(n1018), .ZN(n1020) );
  XNOR2_X1 U1107 ( .A(n1020), .B(KEYINPUT125), .ZN(n1021) );
  NOR2_X1 U1108 ( .A1(n1022), .A2(n1021), .ZN(n1023) );
  XNOR2_X1 U1109 ( .A(n1023), .B(KEYINPUT61), .ZN(n1026) );
  NOR2_X1 U1110 ( .A1(KEYINPUT56), .A2(n1024), .ZN(n1025) );
  NOR2_X1 U1111 ( .A1(n1026), .A2(n1025), .ZN(n1027) );
  NOR2_X1 U1112 ( .A1(G16), .A2(n1027), .ZN(n1028) );
  NOR2_X1 U1113 ( .A1(n1029), .A2(n1028), .ZN(n1030) );
  NAND2_X1 U1114 ( .A1(n1031), .A2(n1030), .ZN(n1032) );
  XNOR2_X1 U1115 ( .A(KEYINPUT62), .B(n1032), .ZN(G150) );
  INV_X1 U1116 ( .A(G150), .ZN(G311) );
endmodule

