

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, n371,
         n372, n373, n374, n375, n376, n377, n378, n379, n380, n381, n382,
         n383, n384, n385, n386, n387, n388, n389, n390, n391, n392, n393,
         n394, n395, n396, n397, n398, n399, n400, n401, n403, n404, n405,
         n406, n407, n408, n409, n410, n411, n412, n413, n414, n415, n416,
         n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, n427,
         n428, n429, n430, n431, n432, n433, n435, n436, n437, n438, n439,
         n440, n441, n442, n443, n444, n445, n446, n447, n448, n449, n450,
         n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, n461,
         n462, n463, n464, n465, n466, n467, n468, n469, n470, n471, n472,
         n473, n474, n475, n476, n477, n478, n479, n480, n481, n482, n483,
         n484, n485, n486, n487, n488, n489, n490, n491, n492, n493, n494,
         n495, n496, n497, n498, n499, n500, n501, n502, n503, n504, n505,
         n506, n507, n508, n509, n510, n511, n512, n513, n514, n515, n516,
         n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527,
         n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538,
         n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549,
         n550, n551, n552, n553, n555, n556, n557, n558, n559, n560, n561,
         n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572,
         n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583,
         n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594,
         n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605,
         n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616,
         n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627,
         n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, n638,
         n639, n640, n641, n642, n643, n644, n645, n646, n647, n648, n649,
         n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, n660,
         n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, n671,
         n672, n673, n674, n675, n676, n677, n678, n679, n680, n681, n682,
         n683, n684, n685, n686, n687, n688, n689, n690, n691, n692, n693,
         n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, n704,
         n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n715,
         n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726,
         n727, n728, n729, n730, n731, n732, n733, n734, n735, n736, n737,
         n738, n739, n740, n741, n742, n743, n744, n745, n746, n747, n748,
         n749, n750, n751, n752, n753, n754, n755, n756, n757, n758, n759,
         n760, n761, n762, n763, n764, n765, n766, n767, n768, n769, n770,
         n771, n772;

  INV_X1 U382 ( .A(n401), .ZN(n362) );
  NOR2_X1 U383 ( .A1(n772), .A2(n767), .ZN(n593) );
  XNOR2_X1 U384 ( .A(n588), .B(n393), .ZN(n772) );
  NOR2_X1 U385 ( .A1(n472), .A2(n699), .ZN(n677) );
  NOR2_X1 U386 ( .A1(n688), .A2(n683), .ZN(n587) );
  AND2_X1 U387 ( .A1(n618), .A2(n617), .ZN(n619) );
  NAND2_X1 U388 ( .A1(n416), .A2(n419), .ZN(n580) );
  XNOR2_X1 U389 ( .A(n461), .B(n544), .ZN(n756) );
  NAND2_X1 U390 ( .A1(n432), .A2(n431), .ZN(n430) );
  XOR2_X1 U391 ( .A(KEYINPUT66), .B(G131), .Z(n513) );
  XNOR2_X1 U392 ( .A(n363), .B(n747), .ZN(n723) );
  XNOR2_X1 U393 ( .A(G143), .B(G128), .ZN(n512) );
  INV_X2 U394 ( .A(G953), .ZN(n750) );
  XNOR2_X2 U395 ( .A(n361), .B(n377), .ZN(n742) );
  NAND2_X1 U396 ( .A1(n435), .A2(n641), .ZN(n361) );
  XNOR2_X2 U397 ( .A(n576), .B(n455), .ZN(n626) );
  NOR2_X1 U398 ( .A1(n721), .A2(n722), .ZN(n382) );
  INV_X1 U399 ( .A(n580), .ZN(n442) );
  NOR2_X2 U400 ( .A1(n597), .A2(n765), .ZN(n645) );
  OR2_X2 U401 ( .A1(n742), .A2(n362), .ZN(n405) );
  XNOR2_X1 U402 ( .A(n404), .B(n470), .ZN(n363) );
  NAND2_X2 U403 ( .A1(n661), .A2(n601), .ZN(n463) );
  NAND2_X2 U404 ( .A1(n420), .A2(n417), .ZN(n661) );
  XNOR2_X2 U405 ( .A(n400), .B(KEYINPUT88), .ZN(n636) );
  XOR2_X1 U406 ( .A(KEYINPUT24), .B(G110), .Z(n518) );
  NOR2_X1 U407 ( .A1(n699), .A2(n403), .ZN(n630) );
  AND2_X4 U408 ( .A1(n454), .A2(n452), .ZN(n737) );
  NOR2_X2 U409 ( .A1(n720), .A2(n555), .ZN(n452) );
  BUF_X2 U410 ( .A(n602), .Z(n364) );
  XNOR2_X1 U411 ( .A(n536), .B(n408), .ZN(n602) );
  NOR2_X2 U412 ( .A1(n769), .A2(n766), .ZN(n400) );
  XNOR2_X1 U413 ( .A(n562), .B(n561), .ZN(n589) );
  XNOR2_X1 U414 ( .A(n445), .B(n444), .ZN(n694) );
  XNOR2_X1 U415 ( .A(n372), .B(n529), .ZN(n551) );
  XNOR2_X1 U416 ( .A(n512), .B(KEYINPUT4), .ZN(n544) );
  NAND2_X1 U417 ( .A1(n411), .A2(n410), .ZN(n541) );
  XNOR2_X2 U418 ( .A(n463), .B(n462), .ZN(n611) );
  XNOR2_X1 U419 ( .A(n385), .B(KEYINPUT47), .ZN(n582) );
  XNOR2_X1 U420 ( .A(n593), .B(n376), .ZN(n594) );
  OR2_X1 U421 ( .A1(G902), .A2(G237), .ZN(n556) );
  NOR2_X1 U422 ( .A1(G953), .A2(G237), .ZN(n531) );
  XNOR2_X1 U423 ( .A(G116), .B(KEYINPUT68), .ZN(n529) );
  XNOR2_X1 U424 ( .A(n513), .B(G134), .ZN(n461) );
  XNOR2_X1 U425 ( .A(n544), .B(n471), .ZN(n470) );
  XNOR2_X1 U426 ( .A(n409), .B(n547), .ZN(n404) );
  AND2_X1 U427 ( .A1(n626), .A2(n456), .ZN(n618) );
  INV_X1 U428 ( .A(n698), .ZN(n456) );
  XNOR2_X1 U429 ( .A(n525), .B(KEYINPUT25), .ZN(n444) );
  OR2_X1 U430 ( .A1(n739), .A2(G902), .ZN(n445) );
  NOR2_X1 U431 ( .A1(n730), .A2(G902), .ZN(n514) );
  NAND2_X1 U432 ( .A1(n560), .A2(n585), .ZN(n562) );
  XNOR2_X1 U433 ( .A(KEYINPUT73), .B(G472), .ZN(n408) );
  NAND2_X1 U434 ( .A1(n737), .A2(G472), .ZN(n415) );
  XNOR2_X1 U435 ( .A(n448), .B(G146), .ZN(n540) );
  INV_X1 U436 ( .A(G125), .ZN(n448) );
  XNOR2_X1 U437 ( .A(n541), .B(n542), .ZN(n409) );
  AND2_X1 U438 ( .A1(n686), .A2(n426), .ZN(n425) );
  XNOR2_X1 U439 ( .A(G113), .B(G104), .ZN(n552) );
  INV_X1 U440 ( .A(KEYINPUT87), .ZN(n433) );
  AND2_X1 U441 ( .A1(n635), .A2(n375), .ZN(n435) );
  XNOR2_X1 U442 ( .A(n540), .B(n447), .ZN(n515) );
  INV_X1 U443 ( .A(KEYINPUT10), .ZN(n447) );
  XOR2_X1 U444 ( .A(KEYINPUT65), .B(G101), .Z(n545) );
  XOR2_X1 U445 ( .A(G137), .B(G140), .Z(n516) );
  NAND2_X1 U446 ( .A1(n365), .A2(n643), .ZN(n431) );
  INV_X1 U447 ( .A(KEYINPUT19), .ZN(n426) );
  NAND2_X1 U448 ( .A1(n694), .A2(n608), .ZN(n698) );
  INV_X1 U449 ( .A(KEYINPUT0), .ZN(n462) );
  XNOR2_X1 U450 ( .A(n551), .B(n407), .ZN(n533) );
  XNOR2_X1 U451 ( .A(G128), .B(G119), .ZN(n517) );
  XNOR2_X1 U452 ( .A(n515), .B(n446), .ZN(n755) );
  INV_X1 U453 ( .A(n516), .ZN(n446) );
  AND2_X1 U454 ( .A1(n520), .A2(G221), .ZN(n521) );
  XNOR2_X1 U455 ( .A(n500), .B(n495), .ZN(n384) );
  XNOR2_X1 U456 ( .A(G116), .B(G134), .ZN(n493) );
  XNOR2_X1 U457 ( .A(n557), .B(n558), .ZN(n590) );
  NAND2_X1 U458 ( .A1(n618), .A2(n364), .ZN(n706) );
  AND2_X1 U459 ( .A1(n406), .A2(n366), .ZN(n662) );
  XNOR2_X1 U460 ( .A(n575), .B(KEYINPUT28), .ZN(n406) );
  AND2_X1 U461 ( .A1(n574), .A2(n573), .ZN(n575) );
  XNOR2_X1 U462 ( .A(n486), .B(n398), .ZN(n585) );
  XNOR2_X1 U463 ( .A(n487), .B(n399), .ZN(n398) );
  INV_X1 U464 ( .A(KEYINPUT13), .ZN(n399) );
  BUF_X1 U465 ( .A(n694), .Z(n403) );
  INV_X1 U466 ( .A(KEYINPUT1), .ZN(n455) );
  NAND2_X1 U467 ( .A1(n395), .A2(n394), .ZN(n465) );
  INV_X1 U468 ( .A(n617), .ZN(n394) );
  INV_X1 U469 ( .A(KEYINPUT86), .ZN(n383) );
  INV_X1 U470 ( .A(KEYINPUT75), .ZN(n437) );
  XOR2_X1 U471 ( .A(KEYINPUT96), .B(KEYINPUT99), .Z(n476) );
  XNOR2_X1 U472 ( .A(KEYINPUT11), .B(KEYINPUT12), .ZN(n475) );
  XNOR2_X1 U473 ( .A(KEYINPUT18), .B(KEYINPUT17), .ZN(n546) );
  XNOR2_X1 U474 ( .A(KEYINPUT90), .B(KEYINPUT77), .ZN(n543) );
  NAND2_X1 U475 ( .A1(n429), .A2(n555), .ZN(n428) );
  INV_X1 U476 ( .A(n365), .ZN(n429) );
  XNOR2_X1 U477 ( .A(n530), .B(G113), .ZN(n407) );
  XOR2_X1 U478 ( .A(KEYINPUT5), .B(G137), .Z(n530) );
  INV_X1 U479 ( .A(KEYINPUT101), .ZN(n499) );
  XOR2_X1 U480 ( .A(KEYINPUT100), .B(KEYINPUT7), .Z(n494) );
  XOR2_X1 U481 ( .A(G143), .B(KEYINPUT98), .Z(n480) );
  NAND2_X1 U482 ( .A1(n507), .A2(n508), .ZN(n411) );
  XNOR2_X1 U483 ( .A(n442), .B(KEYINPUT38), .ZN(n685) );
  NAND2_X1 U484 ( .A1(n424), .A2(n423), .ZN(n422) );
  OR2_X1 U485 ( .A1(n686), .A2(n426), .ZN(n423) );
  AND2_X1 U486 ( .A1(n427), .A2(n425), .ZN(n421) );
  INV_X1 U487 ( .A(n427), .ZN(n419) );
  AND2_X1 U488 ( .A1(n602), .A2(n374), .ZN(n573) );
  XNOR2_X1 U489 ( .A(n551), .B(n550), .ZN(n553) );
  XOR2_X1 U490 ( .A(KEYINPUT74), .B(KEYINPUT16), .Z(n548) );
  INV_X1 U491 ( .A(KEYINPUT84), .ZN(n397) );
  XNOR2_X1 U492 ( .A(n756), .B(n370), .ZN(n535) );
  INV_X1 U493 ( .A(n545), .ZN(n511) );
  INV_X1 U494 ( .A(n541), .ZN(n460) );
  XNOR2_X1 U495 ( .A(n516), .B(n368), .ZN(n509) );
  AND2_X1 U496 ( .A1(n443), .A2(n539), .ZN(n579) );
  AND2_X1 U497 ( .A1(n605), .A2(n374), .ZN(n443) );
  NAND2_X1 U498 ( .A1(n419), .A2(n418), .ZN(n417) );
  NOR2_X1 U499 ( .A1(n422), .A2(n421), .ZN(n420) );
  NOR2_X1 U500 ( .A1(n430), .A2(n426), .ZN(n418) );
  NOR2_X1 U501 ( .A1(n698), .A2(n576), .ZN(n605) );
  NAND2_X1 U502 ( .A1(G953), .A2(G900), .ZN(n761) );
  XNOR2_X1 U503 ( .A(n391), .B(n523), .ZN(n739) );
  XNOR2_X1 U504 ( .A(n521), .B(n522), .ZN(n391) );
  XNOR2_X1 U505 ( .A(n390), .B(n498), .ZN(n735) );
  XNOR2_X1 U506 ( .A(n384), .B(n496), .ZN(n390) );
  XNOR2_X1 U507 ( .A(n535), .B(n457), .ZN(n730) );
  XNOR2_X1 U508 ( .A(n459), .B(n458), .ZN(n457) );
  XNOR2_X1 U509 ( .A(n510), .B(KEYINPUT76), .ZN(n458) );
  XNOR2_X1 U510 ( .A(n509), .B(n460), .ZN(n459) );
  INV_X1 U511 ( .A(KEYINPUT42), .ZN(n393) );
  XNOR2_X1 U512 ( .A(KEYINPUT78), .B(KEYINPUT35), .ZN(n449) );
  INV_X1 U513 ( .A(KEYINPUT31), .ZN(n386) );
  INV_X1 U514 ( .A(KEYINPUT108), .ZN(n563) );
  AND2_X1 U515 ( .A1(n579), .A2(n441), .ZN(n667) );
  NOR2_X1 U516 ( .A1(n623), .A2(n442), .ZN(n441) );
  XNOR2_X1 U517 ( .A(n629), .B(KEYINPUT107), .ZN(n766) );
  NOR2_X1 U518 ( .A1(n585), .A2(n560), .ZN(n674) );
  NOR2_X1 U519 ( .A1(n626), .A2(n613), .ZN(n655) );
  NAND2_X1 U520 ( .A1(n414), .A2(n413), .ZN(n412) );
  XNOR2_X1 U521 ( .A(n415), .B(n654), .ZN(n414) );
  INV_X1 U522 ( .A(KEYINPUT56), .ZN(n466) );
  INV_X1 U523 ( .A(KEYINPUT53), .ZN(n379) );
  XNOR2_X1 U524 ( .A(n382), .B(KEYINPUT122), .ZN(n381) );
  AND2_X1 U525 ( .A1(G210), .A2(n556), .ZN(n365) );
  XNOR2_X1 U526 ( .A(n576), .B(KEYINPUT111), .ZN(n366) );
  XOR2_X1 U527 ( .A(KEYINPUT106), .B(n630), .Z(n367) );
  XOR2_X1 U528 ( .A(G104), .B(G107), .Z(n368) );
  NOR2_X1 U529 ( .A1(n675), .A2(n657), .ZN(n369) );
  XNOR2_X1 U530 ( .A(n511), .B(G146), .ZN(n370) );
  XOR2_X1 U531 ( .A(KEYINPUT80), .B(n644), .Z(n371) );
  XOR2_X1 U532 ( .A(G119), .B(KEYINPUT3), .Z(n372) );
  XNOR2_X1 U533 ( .A(n450), .B(n449), .ZN(n770) );
  AND2_X1 U534 ( .A1(n616), .A2(n615), .ZN(n373) );
  AND2_X1 U535 ( .A1(n600), .A2(n761), .ZN(n374) );
  AND2_X1 U536 ( .A1(n634), .A2(n373), .ZN(n375) );
  XNOR2_X1 U537 ( .A(KEYINPUT64), .B(KEYINPUT46), .ZN(n376) );
  XNOR2_X1 U538 ( .A(G902), .B(KEYINPUT15), .ZN(n555) );
  XOR2_X1 U539 ( .A(KEYINPUT45), .B(KEYINPUT85), .Z(n377) );
  XOR2_X1 U540 ( .A(KEYINPUT91), .B(KEYINPUT63), .Z(n378) );
  INV_X1 U541 ( .A(n741), .ZN(n413) );
  XNOR2_X1 U542 ( .A(n380), .B(n379), .ZN(G75) );
  NAND2_X1 U543 ( .A1(n381), .A2(n750), .ZN(n380) );
  NAND2_X1 U544 ( .A1(n723), .A2(n365), .ZN(n432) );
  XNOR2_X1 U545 ( .A(n612), .B(KEYINPUT22), .ZN(n625) );
  NAND2_X1 U546 ( .A1(n637), .A2(n383), .ZN(n634) );
  NAND2_X1 U547 ( .A1(n430), .A2(n425), .ZN(n424) );
  NAND2_X1 U548 ( .A1(n578), .A2(n662), .ZN(n385) );
  XNOR2_X1 U549 ( .A(n603), .B(n386), .ZN(n675) );
  XNOR2_X1 U550 ( .A(n387), .B(n651), .ZN(G60) );
  NOR2_X2 U551 ( .A1(n649), .A2(n741), .ZN(n387) );
  XNOR2_X2 U552 ( .A(n464), .B(KEYINPUT32), .ZN(n769) );
  INV_X1 U553 ( .A(n625), .ZN(n395) );
  XNOR2_X1 U554 ( .A(n388), .B(KEYINPUT124), .ZN(G54) );
  NOR2_X2 U555 ( .A1(n733), .A2(n741), .ZN(n388) );
  XNOR2_X1 U556 ( .A(n389), .B(KEYINPUT67), .ZN(n595) );
  NAND2_X1 U557 ( .A1(n436), .A2(n392), .ZN(n389) );
  OR2_X2 U558 ( .A1(n719), .A2(KEYINPUT2), .ZN(n440) );
  NOR2_X1 U559 ( .A1(n582), .A2(n581), .ZN(n583) );
  NAND2_X1 U560 ( .A1(n611), .A2(n610), .ZN(n612) );
  INV_X1 U561 ( .A(KEYINPUT2), .ZN(n401) );
  NOR2_X2 U562 ( .A1(n465), .A2(n367), .ZN(n464) );
  XNOR2_X1 U563 ( .A(n622), .B(n621), .ZN(n451) );
  XNOR2_X1 U564 ( .A(n636), .B(n433), .ZN(n640) );
  NAND2_X1 U565 ( .A1(n590), .A2(n589), .ZN(n591) );
  INV_X1 U566 ( .A(n677), .ZN(n392) );
  NAND2_X1 U567 ( .A1(n685), .A2(n686), .ZN(n683) );
  INV_X1 U568 ( .A(n465), .ZN(n631) );
  NOR2_X1 U569 ( .A1(n438), .A2(n396), .ZN(n721) );
  NAND2_X1 U570 ( .A1(n440), .A2(n439), .ZN(n396) );
  XNOR2_X2 U571 ( .A(n598), .B(n397), .ZN(n719) );
  XNOR2_X1 U572 ( .A(n405), .B(KEYINPUT83), .ZN(n438) );
  NAND2_X1 U573 ( .A1(n636), .A2(n632), .ZN(n633) );
  NAND2_X1 U574 ( .A1(n451), .A2(n624), .ZN(n450) );
  NAND2_X1 U575 ( .A1(n645), .A2(n771), .ZN(n598) );
  XNOR2_X1 U576 ( .A(n587), .B(n586), .ZN(n679) );
  XNOR2_X1 U577 ( .A(n412), .B(n378), .ZN(G57) );
  NAND2_X1 U578 ( .A1(n749), .A2(KEYINPUT70), .ZN(n410) );
  INV_X1 U579 ( .A(n430), .ZN(n416) );
  NOR2_X1 U580 ( .A1(n723), .A2(n428), .ZN(n427) );
  NAND2_X1 U581 ( .A1(n719), .A2(n742), .ZN(n642) );
  XNOR2_X1 U582 ( .A(n583), .B(n437), .ZN(n436) );
  INV_X1 U583 ( .A(n720), .ZN(n439) );
  AND2_X2 U584 ( .A1(n742), .A2(n453), .ZN(n720) );
  AND2_X1 U585 ( .A1(n645), .A2(n371), .ZN(n453) );
  NAND2_X1 U586 ( .A1(n642), .A2(n401), .ZN(n454) );
  INV_X1 U587 ( .A(n626), .ZN(n699) );
  XNOR2_X2 U588 ( .A(n514), .B(G469), .ZN(n576) );
  INV_X1 U589 ( .A(n611), .ZN(n620) );
  XNOR2_X1 U590 ( .A(n467), .B(n466), .ZN(G51) );
  NAND2_X1 U591 ( .A1(n468), .A2(n413), .ZN(n467) );
  XNOR2_X1 U592 ( .A(n469), .B(n728), .ZN(n468) );
  NAND2_X1 U593 ( .A1(n737), .A2(G210), .ZN(n469) );
  XNOR2_X1 U594 ( .A(n540), .B(n543), .ZN(n471) );
  XNOR2_X1 U595 ( .A(n732), .B(n731), .ZN(n733) );
  XOR2_X1 U596 ( .A(n572), .B(KEYINPUT36), .Z(n472) );
  XNOR2_X1 U597 ( .A(n473), .B(G122), .ZN(n474) );
  NAND2_X1 U598 ( .A1(n595), .A2(n594), .ZN(n596) );
  XNOR2_X1 U599 ( .A(n552), .B(n474), .ZN(n478) );
  XNOR2_X1 U600 ( .A(n596), .B(KEYINPUT48), .ZN(n597) );
  XNOR2_X1 U601 ( .A(n533), .B(n532), .ZN(n534) );
  XNOR2_X1 U602 ( .A(n549), .B(n548), .ZN(n550) );
  XNOR2_X1 U603 ( .A(n483), .B(n515), .ZN(n484) );
  NOR2_X1 U604 ( .A1(n688), .A2(n609), .ZN(n610) );
  XNOR2_X1 U605 ( .A(n535), .B(n534), .ZN(n652) );
  XNOR2_X1 U606 ( .A(n485), .B(n484), .ZN(n646) );
  XNOR2_X1 U607 ( .A(KEYINPUT113), .B(KEYINPUT41), .ZN(n586) );
  INV_X1 U608 ( .A(KEYINPUT104), .ZN(n561) );
  XNOR2_X1 U609 ( .A(KEYINPUT103), .B(G478), .ZN(n501) );
  XNOR2_X1 U610 ( .A(n730), .B(n729), .ZN(n731) );
  XNOR2_X1 U611 ( .A(n502), .B(n501), .ZN(n584) );
  NOR2_X1 U612 ( .A1(G952), .A2(n750), .ZN(n741) );
  INV_X1 U613 ( .A(G475), .ZN(n487) );
  INV_X1 U614 ( .A(KEYINPUT97), .ZN(n473) );
  XNOR2_X1 U615 ( .A(n476), .B(n475), .ZN(n477) );
  XNOR2_X1 U616 ( .A(n477), .B(n478), .ZN(n482) );
  NAND2_X1 U617 ( .A1(G214), .A2(n531), .ZN(n479) );
  XNOR2_X1 U618 ( .A(n480), .B(n479), .ZN(n481) );
  XNOR2_X1 U619 ( .A(n482), .B(n481), .ZN(n485) );
  XOR2_X1 U620 ( .A(n513), .B(G140), .Z(n483) );
  NOR2_X1 U621 ( .A1(G902), .A2(n646), .ZN(n486) );
  INV_X1 U622 ( .A(n512), .ZN(n488) );
  NAND2_X1 U623 ( .A1(n488), .A2(KEYINPUT9), .ZN(n491) );
  INV_X1 U624 ( .A(KEYINPUT9), .ZN(n489) );
  NAND2_X1 U625 ( .A1(n512), .A2(n489), .ZN(n490) );
  NAND2_X1 U626 ( .A1(n491), .A2(n490), .ZN(n492) );
  XNOR2_X1 U627 ( .A(n492), .B(KEYINPUT102), .ZN(n496) );
  XNOR2_X1 U628 ( .A(n494), .B(n493), .ZN(n495) );
  NAND2_X1 U629 ( .A1(n750), .A2(G234), .ZN(n497) );
  XOR2_X1 U630 ( .A(KEYINPUT8), .B(n497), .Z(n520) );
  AND2_X1 U631 ( .A1(G217), .A2(n520), .ZN(n498) );
  XOR2_X1 U632 ( .A(G122), .B(G107), .Z(n549) );
  XNOR2_X1 U633 ( .A(n549), .B(n499), .ZN(n500) );
  NOR2_X1 U634 ( .A1(G902), .A2(n735), .ZN(n502) );
  INV_X1 U635 ( .A(n584), .ZN(n560) );
  XOR2_X1 U636 ( .A(KEYINPUT71), .B(KEYINPUT39), .Z(n558) );
  NAND2_X1 U637 ( .A1(G234), .A2(G237), .ZN(n503) );
  XNOR2_X1 U638 ( .A(KEYINPUT14), .B(n503), .ZN(n681) );
  OR2_X1 U639 ( .A1(n750), .A2(G902), .ZN(n504) );
  NAND2_X1 U640 ( .A1(n681), .A2(n504), .ZN(n506) );
  NOR2_X1 U641 ( .A1(G953), .A2(G952), .ZN(n505) );
  NOR2_X1 U642 ( .A1(n506), .A2(n505), .ZN(n600) );
  XNOR2_X2 U643 ( .A(KEYINPUT92), .B(G110), .ZN(n749) );
  INV_X1 U644 ( .A(KEYINPUT70), .ZN(n508) );
  INV_X1 U645 ( .A(n749), .ZN(n507) );
  NAND2_X1 U646 ( .A1(G227), .A2(n750), .ZN(n510) );
  XNOR2_X1 U647 ( .A(n755), .B(KEYINPUT23), .ZN(n523) );
  XNOR2_X1 U648 ( .A(n518), .B(n517), .ZN(n519) );
  XOR2_X1 U649 ( .A(n519), .B(KEYINPUT69), .Z(n522) );
  NAND2_X1 U650 ( .A1(G234), .A2(n555), .ZN(n524) );
  XNOR2_X1 U651 ( .A(KEYINPUT20), .B(n524), .ZN(n526) );
  AND2_X1 U652 ( .A1(G217), .A2(n526), .ZN(n525) );
  XOR2_X1 U653 ( .A(KEYINPUT93), .B(KEYINPUT21), .Z(n528) );
  NAND2_X1 U654 ( .A1(n526), .A2(G221), .ZN(n527) );
  XNOR2_X1 U655 ( .A(n528), .B(n527), .ZN(n695) );
  XOR2_X1 U656 ( .A(n695), .B(KEYINPUT94), .Z(n608) );
  XOR2_X1 U657 ( .A(KEYINPUT30), .B(KEYINPUT110), .Z(n538) );
  NAND2_X1 U658 ( .A1(n531), .A2(G210), .ZN(n532) );
  NOR2_X1 U659 ( .A1(G902), .A2(n652), .ZN(n536) );
  NAND2_X1 U660 ( .A1(G214), .A2(n556), .ZN(n686) );
  NAND2_X1 U661 ( .A1(n364), .A2(n686), .ZN(n537) );
  XNOR2_X1 U662 ( .A(n538), .B(n537), .ZN(n539) );
  NAND2_X1 U663 ( .A1(G224), .A2(n750), .ZN(n542) );
  XOR2_X1 U664 ( .A(n546), .B(n545), .Z(n547) );
  XNOR2_X1 U665 ( .A(n553), .B(n552), .ZN(n747) );
  INV_X1 U666 ( .A(n555), .ZN(n643) );
  NAND2_X1 U667 ( .A1(n579), .A2(n685), .ZN(n557) );
  NAND2_X1 U668 ( .A1(n674), .A2(n590), .ZN(n559) );
  XNOR2_X1 U669 ( .A(n559), .B(KEYINPUT114), .ZN(n771) );
  XNOR2_X1 U670 ( .A(n589), .B(n563), .ZN(n669) );
  XNOR2_X1 U671 ( .A(KEYINPUT105), .B(KEYINPUT6), .ZN(n564) );
  XNOR2_X1 U672 ( .A(n564), .B(n364), .ZN(n617) );
  AND2_X1 U673 ( .A1(n374), .A2(n686), .ZN(n565) );
  NOR2_X1 U674 ( .A1(n695), .A2(n694), .ZN(n574) );
  AND2_X1 U675 ( .A1(n565), .A2(n574), .ZN(n566) );
  NAND2_X1 U676 ( .A1(n617), .A2(n566), .ZN(n567) );
  NOR2_X1 U677 ( .A1(n669), .A2(n567), .ZN(n571) );
  NAND2_X1 U678 ( .A1(n699), .A2(n571), .ZN(n568) );
  XNOR2_X1 U679 ( .A(n568), .B(KEYINPUT43), .ZN(n569) );
  NAND2_X1 U680 ( .A1(n569), .A2(n442), .ZN(n570) );
  XNOR2_X1 U681 ( .A(KEYINPUT109), .B(n570), .ZN(n765) );
  AND2_X1 U682 ( .A1(n571), .A2(n580), .ZN(n572) );
  INV_X1 U683 ( .A(n674), .ZN(n663) );
  INV_X1 U684 ( .A(n589), .ZN(n577) );
  NAND2_X1 U685 ( .A1(n663), .A2(n577), .ZN(n682) );
  AND2_X1 U686 ( .A1(n661), .A2(n682), .ZN(n578) );
  NAND2_X1 U687 ( .A1(n585), .A2(n584), .ZN(n623) );
  XNOR2_X1 U688 ( .A(n667), .B(KEYINPUT82), .ZN(n581) );
  OR2_X1 U689 ( .A1(n585), .A2(n584), .ZN(n688) );
  NAND2_X1 U690 ( .A1(n662), .A2(n679), .ZN(n588) );
  XOR2_X1 U691 ( .A(KEYINPUT112), .B(KEYINPUT40), .Z(n592) );
  XNOR2_X1 U692 ( .A(n592), .B(n591), .ZN(n767) );
  NAND2_X1 U693 ( .A1(G898), .A2(G953), .ZN(n599) );
  AND2_X1 U694 ( .A1(n600), .A2(n599), .ZN(n601) );
  NOR2_X1 U695 ( .A1(n620), .A2(n706), .ZN(n603) );
  INV_X1 U696 ( .A(n364), .ZN(n604) );
  NAND2_X1 U697 ( .A1(n605), .A2(n604), .ZN(n606) );
  NOR2_X1 U698 ( .A1(n620), .A2(n606), .ZN(n657) );
  XNOR2_X1 U699 ( .A(KEYINPUT95), .B(n369), .ZN(n607) );
  NAND2_X1 U700 ( .A1(n607), .A2(n682), .ZN(n616) );
  INV_X1 U701 ( .A(n608), .ZN(n609) );
  NAND2_X1 U702 ( .A1(n631), .A2(n403), .ZN(n613) );
  NOR2_X1 U703 ( .A1(KEYINPUT44), .A2(KEYINPUT86), .ZN(n614) );
  NOR2_X1 U704 ( .A1(n655), .A2(n614), .ZN(n615) );
  XNOR2_X1 U705 ( .A(n619), .B(KEYINPUT33), .ZN(n693) );
  NOR2_X1 U706 ( .A1(n620), .A2(n693), .ZN(n622) );
  XNOR2_X1 U707 ( .A(KEYINPUT72), .B(KEYINPUT34), .ZN(n621) );
  XNOR2_X1 U708 ( .A(n623), .B(KEYINPUT79), .ZN(n624) );
  NAND2_X1 U709 ( .A1(n770), .A2(KEYINPUT86), .ZN(n632) );
  NOR2_X1 U710 ( .A1(n625), .A2(n403), .ZN(n628) );
  NOR2_X1 U711 ( .A1(n626), .A2(n364), .ZN(n627) );
  NAND2_X1 U712 ( .A1(n628), .A2(n627), .ZN(n629) );
  NAND2_X1 U713 ( .A1(n633), .A2(KEYINPUT44), .ZN(n635) );
  INV_X1 U714 ( .A(KEYINPUT44), .ZN(n638) );
  INV_X1 U715 ( .A(n770), .ZN(n637) );
  AND2_X1 U716 ( .A1(n638), .A2(n637), .ZN(n639) );
  NAND2_X1 U717 ( .A1(n640), .A2(n639), .ZN(n641) );
  NAND2_X1 U718 ( .A1(n771), .A2(KEYINPUT2), .ZN(n644) );
  NAND2_X1 U719 ( .A1(n737), .A2(G475), .ZN(n648) );
  XOR2_X1 U720 ( .A(n646), .B(KEYINPUT59), .Z(n647) );
  XNOR2_X1 U721 ( .A(n648), .B(n647), .ZN(n649) );
  INV_X1 U722 ( .A(KEYINPUT125), .ZN(n650) );
  XNOR2_X1 U723 ( .A(n650), .B(KEYINPUT60), .ZN(n651) );
  XNOR2_X1 U724 ( .A(n652), .B(KEYINPUT62), .ZN(n653) );
  XNOR2_X1 U725 ( .A(n653), .B(KEYINPUT115), .ZN(n654) );
  XOR2_X1 U726 ( .A(G101), .B(n655), .Z(G3) );
  INV_X1 U727 ( .A(n669), .ZN(n672) );
  NAND2_X1 U728 ( .A1(n657), .A2(n672), .ZN(n656) );
  XNOR2_X1 U729 ( .A(n656), .B(G104), .ZN(G6) );
  XOR2_X1 U730 ( .A(KEYINPUT27), .B(KEYINPUT26), .Z(n659) );
  NAND2_X1 U731 ( .A1(n657), .A2(n674), .ZN(n658) );
  XNOR2_X1 U732 ( .A(n659), .B(n658), .ZN(n660) );
  XNOR2_X1 U733 ( .A(G107), .B(n660), .ZN(G9) );
  NAND2_X1 U734 ( .A1(n662), .A2(n661), .ZN(n668) );
  NOR2_X1 U735 ( .A1(n663), .A2(n668), .ZN(n665) );
  XNOR2_X1 U736 ( .A(KEYINPUT116), .B(KEYINPUT29), .ZN(n664) );
  XNOR2_X1 U737 ( .A(n665), .B(n664), .ZN(n666) );
  XNOR2_X1 U738 ( .A(G128), .B(n666), .ZN(G30) );
  XOR2_X1 U739 ( .A(G143), .B(n667), .Z(G45) );
  NOR2_X1 U740 ( .A1(n669), .A2(n668), .ZN(n671) );
  XNOR2_X1 U741 ( .A(G146), .B(KEYINPUT117), .ZN(n670) );
  XNOR2_X1 U742 ( .A(n671), .B(n670), .ZN(G48) );
  NAND2_X1 U743 ( .A1(n675), .A2(n672), .ZN(n673) );
  XNOR2_X1 U744 ( .A(n673), .B(G113), .ZN(G15) );
  NAND2_X1 U745 ( .A1(n675), .A2(n674), .ZN(n676) );
  XNOR2_X1 U746 ( .A(n676), .B(G116), .ZN(G18) );
  XNOR2_X1 U747 ( .A(G125), .B(n677), .ZN(n678) );
  XNOR2_X1 U748 ( .A(n678), .B(KEYINPUT37), .ZN(G27) );
  INV_X1 U749 ( .A(n679), .ZN(n709) );
  NOR2_X1 U750 ( .A1(n709), .A2(n693), .ZN(n680) );
  XNOR2_X1 U751 ( .A(n680), .B(KEYINPUT121), .ZN(n718) );
  INV_X1 U752 ( .A(n681), .ZN(n715) );
  INV_X1 U753 ( .A(n682), .ZN(n684) );
  NOR2_X1 U754 ( .A1(n684), .A2(n683), .ZN(n690) );
  NOR2_X1 U755 ( .A1(n686), .A2(n685), .ZN(n687) );
  NOR2_X1 U756 ( .A1(n688), .A2(n687), .ZN(n689) );
  NOR2_X1 U757 ( .A1(n690), .A2(n689), .ZN(n691) );
  XOR2_X1 U758 ( .A(KEYINPUT119), .B(n691), .Z(n692) );
  NOR2_X1 U759 ( .A1(n693), .A2(n692), .ZN(n711) );
  INV_X1 U760 ( .A(n403), .ZN(n696) );
  NAND2_X1 U761 ( .A1(n696), .A2(n695), .ZN(n697) );
  XOR2_X1 U762 ( .A(KEYINPUT49), .B(n697), .Z(n704) );
  XOR2_X1 U763 ( .A(KEYINPUT50), .B(KEYINPUT118), .Z(n701) );
  NAND2_X1 U764 ( .A1(n699), .A2(n698), .ZN(n700) );
  XNOR2_X1 U765 ( .A(n701), .B(n700), .ZN(n702) );
  NOR2_X1 U766 ( .A1(n702), .A2(n364), .ZN(n703) );
  NAND2_X1 U767 ( .A1(n704), .A2(n703), .ZN(n705) );
  NAND2_X1 U768 ( .A1(n706), .A2(n705), .ZN(n707) );
  XNOR2_X1 U769 ( .A(KEYINPUT51), .B(n707), .ZN(n708) );
  NOR2_X1 U770 ( .A1(n709), .A2(n708), .ZN(n710) );
  NOR2_X1 U771 ( .A1(n711), .A2(n710), .ZN(n712) );
  XNOR2_X1 U772 ( .A(n712), .B(KEYINPUT120), .ZN(n713) );
  XNOR2_X1 U773 ( .A(KEYINPUT52), .B(n713), .ZN(n714) );
  NOR2_X1 U774 ( .A1(n715), .A2(n714), .ZN(n716) );
  NAND2_X1 U775 ( .A1(n716), .A2(G952), .ZN(n717) );
  NAND2_X1 U776 ( .A1(n718), .A2(n717), .ZN(n722) );
  INV_X1 U777 ( .A(n719), .ZN(n757) );
  XNOR2_X1 U778 ( .A(KEYINPUT89), .B(KEYINPUT55), .ZN(n725) );
  XNOR2_X1 U779 ( .A(n723), .B(KEYINPUT81), .ZN(n724) );
  XNOR2_X1 U780 ( .A(n725), .B(n724), .ZN(n727) );
  XOR2_X1 U781 ( .A(KEYINPUT123), .B(KEYINPUT54), .Z(n726) );
  XNOR2_X1 U782 ( .A(n727), .B(n726), .ZN(n728) );
  NAND2_X1 U783 ( .A1(n737), .A2(G469), .ZN(n732) );
  XOR2_X1 U784 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n729) );
  NAND2_X1 U785 ( .A1(G478), .A2(n737), .ZN(n734) );
  XNOR2_X1 U786 ( .A(n735), .B(n734), .ZN(n736) );
  NOR2_X1 U787 ( .A1(n741), .A2(n736), .ZN(G63) );
  NAND2_X1 U788 ( .A1(G217), .A2(n737), .ZN(n738) );
  XNOR2_X1 U789 ( .A(n739), .B(n738), .ZN(n740) );
  NOR2_X1 U790 ( .A1(n741), .A2(n740), .ZN(G66) );
  NAND2_X1 U791 ( .A1(n750), .A2(n742), .ZN(n746) );
  NAND2_X1 U792 ( .A1(G953), .A2(G224), .ZN(n743) );
  XNOR2_X1 U793 ( .A(KEYINPUT61), .B(n743), .ZN(n744) );
  NAND2_X1 U794 ( .A1(n744), .A2(G898), .ZN(n745) );
  NAND2_X1 U795 ( .A1(n746), .A2(n745), .ZN(n754) );
  XOR2_X1 U796 ( .A(n747), .B(G101), .Z(n748) );
  XNOR2_X1 U797 ( .A(n749), .B(n748), .ZN(n752) );
  NOR2_X1 U798 ( .A1(G898), .A2(n750), .ZN(n751) );
  NOR2_X1 U799 ( .A1(n752), .A2(n751), .ZN(n753) );
  XNOR2_X1 U800 ( .A(n754), .B(n753), .ZN(G69) );
  XOR2_X1 U801 ( .A(n756), .B(n755), .Z(n759) );
  XOR2_X1 U802 ( .A(n759), .B(n757), .Z(n758) );
  NOR2_X1 U803 ( .A1(G953), .A2(n758), .ZN(n763) );
  XNOR2_X1 U804 ( .A(n759), .B(G227), .ZN(n760) );
  NOR2_X1 U805 ( .A1(n761), .A2(n760), .ZN(n762) );
  NOR2_X1 U806 ( .A1(n763), .A2(n762), .ZN(n764) );
  XNOR2_X1 U807 ( .A(KEYINPUT126), .B(n764), .ZN(G72) );
  XOR2_X1 U808 ( .A(G140), .B(n765), .Z(G42) );
  XOR2_X1 U809 ( .A(G110), .B(n766), .Z(G12) );
  XNOR2_X1 U810 ( .A(G131), .B(n767), .ZN(n768) );
  XNOR2_X1 U811 ( .A(n768), .B(KEYINPUT127), .ZN(G33) );
  XOR2_X1 U812 ( .A(n769), .B(G119), .Z(G21) );
  XOR2_X1 U813 ( .A(G122), .B(n770), .Z(G24) );
  XNOR2_X1 U814 ( .A(G134), .B(n771), .ZN(G36) );
  XOR2_X1 U815 ( .A(n772), .B(G137), .Z(G39) );
endmodule

