//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 0 0 0 1 0 0 1 0 0 0 0 1 0 1 1 0 1 1 1 0 0 0 0 1 1 1 1 0 0 0 0 0 1 0 0 0 0 1 0 0 0 1 0 1 0 0 0 1 1 0 0 0 1 1 1 0 0 0 0 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:17:11 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n705, new_n706, new_n707, new_n708, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n750, new_n751, new_n752, new_n754, new_n755, new_n756, new_n757,
    new_n758, new_n759, new_n760, new_n762, new_n764, new_n765, new_n766,
    new_n767, new_n768, new_n769, new_n770, new_n771, new_n772, new_n773,
    new_n774, new_n775, new_n776, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n788, new_n789,
    new_n790, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n843, new_n844, new_n846, new_n847, new_n848, new_n849,
    new_n851, new_n852, new_n853, new_n854, new_n855, new_n856, new_n857,
    new_n858, new_n859, new_n860, new_n861, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n907, new_n908, new_n910,
    new_n911, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n922, new_n923, new_n924, new_n926, new_n927,
    new_n928, new_n929, new_n930, new_n931, new_n932, new_n933, new_n935,
    new_n936, new_n937, new_n938, new_n939, new_n940, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n948, new_n949, new_n950,
    new_n952, new_n953, new_n954, new_n956, new_n957, new_n958, new_n959,
    new_n960, new_n962, new_n963, new_n964, new_n965, new_n966;
  INV_X1    g000(.A(KEYINPUT14), .ZN(new_n202));
  INV_X1    g001(.A(G29gat), .ZN(new_n203));
  INV_X1    g002(.A(G36gat), .ZN(new_n204));
  NAND3_X1  g003(.A1(new_n202), .A2(new_n203), .A3(new_n204), .ZN(new_n205));
  OAI21_X1  g004(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n206));
  NAND2_X1  g005(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  XNOR2_X1  g006(.A(new_n207), .B(KEYINPUT91), .ZN(new_n208));
  XOR2_X1   g007(.A(G43gat), .B(G50gat), .Z(new_n209));
  INV_X1    g008(.A(KEYINPUT15), .ZN(new_n210));
  NOR2_X1   g009(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  INV_X1    g010(.A(new_n211), .ZN(new_n212));
  NAND2_X1  g011(.A1(G29gat), .A2(G36gat), .ZN(new_n213));
  NAND2_X1  g012(.A1(new_n209), .A2(new_n210), .ZN(new_n214));
  NAND4_X1  g013(.A1(new_n208), .A2(new_n212), .A3(new_n213), .A4(new_n214), .ZN(new_n215));
  INV_X1    g014(.A(new_n205), .ZN(new_n216));
  AND2_X1   g015(.A1(new_n216), .A2(KEYINPUT90), .ZN(new_n217));
  OAI21_X1  g016(.A(new_n206), .B1(new_n216), .B2(KEYINPUT90), .ZN(new_n218));
  OAI21_X1  g017(.A(new_n213), .B1(new_n217), .B2(new_n218), .ZN(new_n219));
  NAND2_X1  g018(.A1(new_n219), .A2(new_n211), .ZN(new_n220));
  AND2_X1   g019(.A1(new_n215), .A2(new_n220), .ZN(new_n221));
  NAND2_X1  g020(.A1(new_n221), .A2(KEYINPUT17), .ZN(new_n222));
  XNOR2_X1  g021(.A(G15gat), .B(G22gat), .ZN(new_n223));
  INV_X1    g022(.A(G1gat), .ZN(new_n224));
  NAND3_X1  g023(.A1(new_n223), .A2(KEYINPUT16), .A3(new_n224), .ZN(new_n225));
  OR2_X1    g024(.A1(KEYINPUT92), .A2(G8gat), .ZN(new_n226));
  OAI211_X1 g025(.A(new_n225), .B(new_n226), .C1(new_n224), .C2(new_n223), .ZN(new_n227));
  NAND2_X1  g026(.A1(KEYINPUT92), .A2(G8gat), .ZN(new_n228));
  XOR2_X1   g027(.A(new_n227), .B(new_n228), .Z(new_n229));
  NAND2_X1  g028(.A1(new_n215), .A2(new_n220), .ZN(new_n230));
  INV_X1    g029(.A(KEYINPUT17), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n230), .A2(new_n231), .ZN(new_n232));
  NAND3_X1  g031(.A1(new_n222), .A2(new_n229), .A3(new_n232), .ZN(new_n233));
  NAND2_X1  g032(.A1(G229gat), .A2(G233gat), .ZN(new_n234));
  OR2_X1    g033(.A1(new_n229), .A2(new_n221), .ZN(new_n235));
  NAND3_X1  g034(.A1(new_n233), .A2(new_n234), .A3(new_n235), .ZN(new_n236));
  INV_X1    g035(.A(KEYINPUT18), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n236), .A2(new_n237), .ZN(new_n238));
  XNOR2_X1  g037(.A(new_n229), .B(new_n221), .ZN(new_n239));
  XOR2_X1   g038(.A(new_n234), .B(KEYINPUT13), .Z(new_n240));
  NAND2_X1  g039(.A1(new_n239), .A2(new_n240), .ZN(new_n241));
  NAND4_X1  g040(.A1(new_n233), .A2(new_n235), .A3(KEYINPUT18), .A4(new_n234), .ZN(new_n242));
  NAND3_X1  g041(.A1(new_n238), .A2(new_n241), .A3(new_n242), .ZN(new_n243));
  XNOR2_X1  g042(.A(G113gat), .B(G141gat), .ZN(new_n244));
  XNOR2_X1  g043(.A(KEYINPUT89), .B(G197gat), .ZN(new_n245));
  XNOR2_X1  g044(.A(new_n244), .B(new_n245), .ZN(new_n246));
  XOR2_X1   g045(.A(KEYINPUT11), .B(G169gat), .Z(new_n247));
  XNOR2_X1  g046(.A(new_n246), .B(new_n247), .ZN(new_n248));
  XNOR2_X1  g047(.A(new_n248), .B(KEYINPUT12), .ZN(new_n249));
  INV_X1    g048(.A(new_n249), .ZN(new_n250));
  NAND2_X1  g049(.A1(new_n243), .A2(new_n250), .ZN(new_n251));
  NAND4_X1  g050(.A1(new_n238), .A2(new_n241), .A3(new_n242), .A4(new_n249), .ZN(new_n252));
  NAND2_X1  g051(.A1(new_n251), .A2(new_n252), .ZN(new_n253));
  INV_X1    g052(.A(KEYINPUT93), .ZN(new_n254));
  NAND2_X1  g053(.A1(new_n253), .A2(new_n254), .ZN(new_n255));
  NAND3_X1  g054(.A1(new_n251), .A2(KEYINPUT93), .A3(new_n252), .ZN(new_n256));
  NAND2_X1  g055(.A1(new_n255), .A2(new_n256), .ZN(new_n257));
  INV_X1    g056(.A(new_n257), .ZN(new_n258));
  INV_X1    g057(.A(KEYINPUT73), .ZN(new_n259));
  NAND2_X1  g058(.A1(G227gat), .A2(G233gat), .ZN(new_n260));
  INV_X1    g059(.A(new_n260), .ZN(new_n261));
  OAI21_X1  g060(.A(KEYINPUT34), .B1(new_n261), .B2(KEYINPUT72), .ZN(new_n262));
  INV_X1    g061(.A(G183gat), .ZN(new_n263));
  NAND2_X1  g062(.A1(new_n263), .A2(KEYINPUT27), .ZN(new_n264));
  INV_X1    g063(.A(KEYINPUT27), .ZN(new_n265));
  NAND2_X1  g064(.A1(new_n265), .A2(G183gat), .ZN(new_n266));
  INV_X1    g065(.A(G190gat), .ZN(new_n267));
  NAND3_X1  g066(.A1(new_n264), .A2(new_n266), .A3(new_n267), .ZN(new_n268));
  INV_X1    g067(.A(KEYINPUT67), .ZN(new_n269));
  XNOR2_X1  g068(.A(KEYINPUT66), .B(KEYINPUT28), .ZN(new_n270));
  NAND3_X1  g069(.A1(new_n268), .A2(new_n269), .A3(new_n270), .ZN(new_n271));
  XNOR2_X1  g070(.A(KEYINPUT27), .B(G183gat), .ZN(new_n272));
  NAND3_X1  g071(.A1(new_n272), .A2(KEYINPUT28), .A3(new_n267), .ZN(new_n273));
  NAND2_X1  g072(.A1(new_n271), .A2(new_n273), .ZN(new_n274));
  AOI21_X1  g073(.A(new_n269), .B1(new_n268), .B2(new_n270), .ZN(new_n275));
  OAI21_X1  g074(.A(KEYINPUT68), .B1(new_n274), .B2(new_n275), .ZN(new_n276));
  NAND2_X1  g075(.A1(new_n268), .A2(new_n270), .ZN(new_n277));
  NAND2_X1  g076(.A1(new_n277), .A2(KEYINPUT67), .ZN(new_n278));
  INV_X1    g077(.A(KEYINPUT68), .ZN(new_n279));
  NAND4_X1  g078(.A1(new_n278), .A2(new_n279), .A3(new_n273), .A4(new_n271), .ZN(new_n280));
  NOR2_X1   g079(.A1(G169gat), .A2(G176gat), .ZN(new_n281));
  NAND2_X1  g080(.A1(new_n281), .A2(KEYINPUT26), .ZN(new_n282));
  OAI21_X1  g081(.A(new_n282), .B1(new_n263), .B2(new_n267), .ZN(new_n283));
  NAND2_X1  g082(.A1(G169gat), .A2(G176gat), .ZN(new_n284));
  INV_X1    g083(.A(KEYINPUT26), .ZN(new_n285));
  NAND2_X1  g084(.A1(new_n284), .A2(new_n285), .ZN(new_n286));
  NOR2_X1   g085(.A1(new_n286), .A2(new_n281), .ZN(new_n287));
  NOR2_X1   g086(.A1(new_n283), .A2(new_n287), .ZN(new_n288));
  NAND3_X1  g087(.A1(new_n276), .A2(new_n280), .A3(new_n288), .ZN(new_n289));
  OR2_X1    g088(.A1(new_n281), .A2(KEYINPUT23), .ZN(new_n290));
  NAND2_X1  g089(.A1(new_n281), .A2(KEYINPUT23), .ZN(new_n291));
  NAND3_X1  g090(.A1(new_n290), .A2(new_n291), .A3(new_n284), .ZN(new_n292));
  INV_X1    g091(.A(KEYINPUT25), .ZN(new_n293));
  NOR2_X1   g092(.A1(new_n292), .A2(new_n293), .ZN(new_n294));
  NAND3_X1  g093(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n295));
  INV_X1    g094(.A(KEYINPUT64), .ZN(new_n296));
  NAND2_X1  g095(.A1(new_n295), .A2(new_n296), .ZN(new_n297));
  NAND4_X1  g096(.A1(KEYINPUT64), .A2(KEYINPUT24), .A3(G183gat), .A4(G190gat), .ZN(new_n298));
  NAND2_X1  g097(.A1(new_n297), .A2(new_n298), .ZN(new_n299));
  OAI21_X1  g098(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n300));
  OAI21_X1  g099(.A(new_n300), .B1(new_n263), .B2(new_n267), .ZN(new_n301));
  AND3_X1   g100(.A1(new_n299), .A2(KEYINPUT65), .A3(new_n301), .ZN(new_n302));
  AOI21_X1  g101(.A(KEYINPUT65), .B1(new_n299), .B2(new_n301), .ZN(new_n303));
  OAI21_X1  g102(.A(new_n294), .B1(new_n302), .B2(new_n303), .ZN(new_n304));
  AND2_X1   g103(.A1(new_n301), .A2(new_n295), .ZN(new_n305));
  OAI21_X1  g104(.A(new_n293), .B1(new_n305), .B2(new_n292), .ZN(new_n306));
  NAND2_X1  g105(.A1(new_n304), .A2(new_n306), .ZN(new_n307));
  XOR2_X1   g106(.A(G113gat), .B(G120gat), .Z(new_n308));
  OR2_X1    g107(.A1(new_n308), .A2(KEYINPUT70), .ZN(new_n309));
  XOR2_X1   g108(.A(G127gat), .B(G134gat), .Z(new_n310));
  INV_X1    g109(.A(G120gat), .ZN(new_n311));
  AND3_X1   g110(.A1(new_n311), .A2(KEYINPUT70), .A3(G113gat), .ZN(new_n312));
  NOR3_X1   g111(.A1(new_n310), .A2(KEYINPUT1), .A3(new_n312), .ZN(new_n313));
  NAND2_X1  g112(.A1(new_n309), .A2(new_n313), .ZN(new_n314));
  INV_X1    g113(.A(KEYINPUT69), .ZN(new_n315));
  INV_X1    g114(.A(KEYINPUT1), .ZN(new_n316));
  NAND2_X1  g115(.A1(new_n308), .A2(new_n316), .ZN(new_n317));
  AOI21_X1  g116(.A(new_n315), .B1(new_n317), .B2(new_n310), .ZN(new_n318));
  XNOR2_X1  g117(.A(G113gat), .B(G120gat), .ZN(new_n319));
  OAI211_X1 g118(.A(new_n310), .B(new_n315), .C1(KEYINPUT1), .C2(new_n319), .ZN(new_n320));
  INV_X1    g119(.A(new_n320), .ZN(new_n321));
  OAI21_X1  g120(.A(new_n314), .B1(new_n318), .B2(new_n321), .ZN(new_n322));
  NAND3_X1  g121(.A1(new_n289), .A2(new_n307), .A3(new_n322), .ZN(new_n323));
  INV_X1    g122(.A(new_n323), .ZN(new_n324));
  AOI21_X1  g123(.A(new_n322), .B1(new_n289), .B2(new_n307), .ZN(new_n325));
  OAI211_X1 g124(.A(new_n260), .B(new_n262), .C1(new_n324), .C2(new_n325), .ZN(new_n326));
  INV_X1    g125(.A(new_n326), .ZN(new_n327));
  NAND2_X1  g126(.A1(new_n289), .A2(new_n307), .ZN(new_n328));
  OAI21_X1  g127(.A(new_n310), .B1(KEYINPUT1), .B2(new_n319), .ZN(new_n329));
  NAND2_X1  g128(.A1(new_n329), .A2(KEYINPUT69), .ZN(new_n330));
  AOI22_X1  g129(.A1(new_n330), .A2(new_n320), .B1(new_n309), .B2(new_n313), .ZN(new_n331));
  NAND2_X1  g130(.A1(new_n328), .A2(new_n331), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n332), .A2(new_n323), .ZN(new_n333));
  AOI21_X1  g132(.A(new_n262), .B1(new_n333), .B2(new_n260), .ZN(new_n334));
  NOR2_X1   g133(.A1(new_n327), .A2(new_n334), .ZN(new_n335));
  NAND3_X1  g134(.A1(new_n332), .A2(new_n261), .A3(new_n323), .ZN(new_n336));
  NAND2_X1  g135(.A1(new_n336), .A2(KEYINPUT32), .ZN(new_n337));
  INV_X1    g136(.A(KEYINPUT33), .ZN(new_n338));
  NAND2_X1  g137(.A1(new_n336), .A2(new_n338), .ZN(new_n339));
  XNOR2_X1  g138(.A(KEYINPUT71), .B(G71gat), .ZN(new_n340));
  XNOR2_X1  g139(.A(new_n340), .B(G99gat), .ZN(new_n341));
  XOR2_X1   g140(.A(G15gat), .B(G43gat), .Z(new_n342));
  XOR2_X1   g141(.A(new_n341), .B(new_n342), .Z(new_n343));
  AND3_X1   g142(.A1(new_n337), .A2(new_n339), .A3(new_n343), .ZN(new_n344));
  INV_X1    g143(.A(new_n343), .ZN(new_n345));
  OAI211_X1 g144(.A(new_n336), .B(KEYINPUT32), .C1(new_n338), .C2(new_n345), .ZN(new_n346));
  INV_X1    g145(.A(new_n346), .ZN(new_n347));
  OAI211_X1 g146(.A(new_n259), .B(new_n335), .C1(new_n344), .C2(new_n347), .ZN(new_n348));
  OAI21_X1  g147(.A(KEYINPUT73), .B1(new_n327), .B2(new_n334), .ZN(new_n349));
  INV_X1    g148(.A(new_n262), .ZN(new_n350));
  NOR2_X1   g149(.A1(new_n324), .A2(new_n325), .ZN(new_n351));
  OAI21_X1  g150(.A(new_n350), .B1(new_n351), .B2(new_n261), .ZN(new_n352));
  NAND3_X1  g151(.A1(new_n352), .A2(new_n259), .A3(new_n326), .ZN(new_n353));
  NAND3_X1  g152(.A1(new_n337), .A2(new_n339), .A3(new_n343), .ZN(new_n354));
  NAND4_X1  g153(.A1(new_n349), .A2(new_n353), .A3(new_n346), .A4(new_n354), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n348), .A2(new_n355), .ZN(new_n356));
  INV_X1    g155(.A(KEYINPUT36), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n356), .A2(new_n357), .ZN(new_n358));
  NAND3_X1  g157(.A1(new_n348), .A2(KEYINPUT36), .A3(new_n355), .ZN(new_n359));
  NAND2_X1  g158(.A1(new_n358), .A2(new_n359), .ZN(new_n360));
  XOR2_X1   g159(.A(G8gat), .B(G36gat), .Z(new_n361));
  XNOR2_X1  g160(.A(new_n361), .B(KEYINPUT76), .ZN(new_n362));
  XNOR2_X1  g161(.A(G64gat), .B(G92gat), .ZN(new_n363));
  XOR2_X1   g162(.A(new_n362), .B(new_n363), .Z(new_n364));
  INV_X1    g163(.A(new_n364), .ZN(new_n365));
  INV_X1    g164(.A(KEYINPUT75), .ZN(new_n366));
  XNOR2_X1  g165(.A(G197gat), .B(G204gat), .ZN(new_n367));
  INV_X1    g166(.A(G211gat), .ZN(new_n368));
  INV_X1    g167(.A(G218gat), .ZN(new_n369));
  NOR2_X1   g168(.A1(new_n368), .A2(new_n369), .ZN(new_n370));
  OAI21_X1  g169(.A(new_n367), .B1(KEYINPUT22), .B2(new_n370), .ZN(new_n371));
  XNOR2_X1  g170(.A(G211gat), .B(G218gat), .ZN(new_n372));
  XNOR2_X1  g171(.A(new_n371), .B(new_n372), .ZN(new_n373));
  NAND2_X1  g172(.A1(G226gat), .A2(G233gat), .ZN(new_n374));
  INV_X1    g173(.A(new_n288), .ZN(new_n375));
  NAND3_X1  g174(.A1(new_n278), .A2(new_n273), .A3(new_n271), .ZN(new_n376));
  AOI21_X1  g175(.A(new_n375), .B1(new_n376), .B2(KEYINPUT68), .ZN(new_n377));
  AOI22_X1  g176(.A1(new_n377), .A2(new_n280), .B1(new_n306), .B2(new_n304), .ZN(new_n378));
  OAI21_X1  g177(.A(new_n374), .B1(new_n378), .B2(KEYINPUT29), .ZN(new_n379));
  AOI21_X1  g178(.A(new_n374), .B1(new_n289), .B2(new_n307), .ZN(new_n380));
  INV_X1    g179(.A(new_n380), .ZN(new_n381));
  AOI21_X1  g180(.A(KEYINPUT74), .B1(new_n379), .B2(new_n381), .ZN(new_n382));
  INV_X1    g181(.A(KEYINPUT74), .ZN(new_n383));
  INV_X1    g182(.A(KEYINPUT29), .ZN(new_n384));
  NAND2_X1  g183(.A1(new_n328), .A2(new_n384), .ZN(new_n385));
  AOI21_X1  g184(.A(new_n383), .B1(new_n385), .B2(new_n374), .ZN(new_n386));
  OAI211_X1 g185(.A(new_n366), .B(new_n373), .C1(new_n382), .C2(new_n386), .ZN(new_n387));
  INV_X1    g186(.A(new_n374), .ZN(new_n388));
  AOI21_X1  g187(.A(KEYINPUT29), .B1(new_n289), .B2(new_n307), .ZN(new_n389));
  OAI21_X1  g188(.A(new_n381), .B1(new_n388), .B2(new_n389), .ZN(new_n390));
  NOR2_X1   g189(.A1(new_n390), .A2(new_n373), .ZN(new_n391));
  INV_X1    g190(.A(new_n391), .ZN(new_n392));
  NAND2_X1  g191(.A1(new_n387), .A2(new_n392), .ZN(new_n393));
  INV_X1    g192(.A(new_n373), .ZN(new_n394));
  AOI21_X1  g193(.A(new_n388), .B1(new_n328), .B2(new_n384), .ZN(new_n395));
  OAI21_X1  g194(.A(new_n383), .B1(new_n395), .B2(new_n380), .ZN(new_n396));
  NAND2_X1  g195(.A1(new_n379), .A2(KEYINPUT74), .ZN(new_n397));
  AOI21_X1  g196(.A(new_n394), .B1(new_n396), .B2(new_n397), .ZN(new_n398));
  NOR2_X1   g197(.A1(new_n398), .A2(new_n366), .ZN(new_n399));
  OAI21_X1  g198(.A(new_n365), .B1(new_n393), .B2(new_n399), .ZN(new_n400));
  AOI21_X1  g199(.A(new_n391), .B1(new_n398), .B2(new_n366), .ZN(new_n401));
  AOI21_X1  g200(.A(new_n386), .B1(new_n390), .B2(new_n383), .ZN(new_n402));
  OAI21_X1  g201(.A(KEYINPUT75), .B1(new_n402), .B2(new_n394), .ZN(new_n403));
  NAND4_X1  g202(.A1(new_n401), .A2(new_n403), .A3(KEYINPUT30), .A4(new_n364), .ZN(new_n404));
  AND2_X1   g203(.A1(new_n400), .A2(new_n404), .ZN(new_n405));
  INV_X1    g204(.A(KEYINPUT5), .ZN(new_n406));
  XNOR2_X1  g205(.A(KEYINPUT80), .B(G141gat), .ZN(new_n407));
  INV_X1    g206(.A(G148gat), .ZN(new_n408));
  NOR2_X1   g207(.A1(new_n407), .A2(new_n408), .ZN(new_n409));
  NAND2_X1  g208(.A1(new_n409), .A2(KEYINPUT81), .ZN(new_n410));
  AOI21_X1  g209(.A(KEYINPUT81), .B1(new_n408), .B2(G141gat), .ZN(new_n411));
  OAI21_X1  g210(.A(new_n411), .B1(new_n407), .B2(new_n408), .ZN(new_n412));
  OR3_X1    g211(.A1(KEYINPUT2), .A2(G155gat), .A3(G162gat), .ZN(new_n413));
  NAND2_X1  g212(.A1(G155gat), .A2(G162gat), .ZN(new_n414));
  NAND2_X1  g213(.A1(new_n413), .A2(new_n414), .ZN(new_n415));
  NAND3_X1  g214(.A1(new_n410), .A2(new_n412), .A3(new_n415), .ZN(new_n416));
  INV_X1    g215(.A(G155gat), .ZN(new_n417));
  INV_X1    g216(.A(G162gat), .ZN(new_n418));
  NAND2_X1  g217(.A1(new_n417), .A2(new_n418), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n419), .A2(new_n414), .ZN(new_n420));
  XOR2_X1   g219(.A(G141gat), .B(G148gat), .Z(new_n421));
  XOR2_X1   g220(.A(KEYINPUT79), .B(KEYINPUT2), .Z(new_n422));
  AOI21_X1  g221(.A(new_n420), .B1(new_n421), .B2(new_n422), .ZN(new_n423));
  INV_X1    g222(.A(new_n423), .ZN(new_n424));
  NAND2_X1  g223(.A1(new_n416), .A2(new_n424), .ZN(new_n425));
  INV_X1    g224(.A(KEYINPUT82), .ZN(new_n426));
  NAND2_X1  g225(.A1(new_n425), .A2(new_n426), .ZN(new_n427));
  AOI22_X1  g226(.A1(new_n409), .A2(KEYINPUT81), .B1(new_n414), .B2(new_n413), .ZN(new_n428));
  AOI21_X1  g227(.A(new_n423), .B1(new_n428), .B2(new_n412), .ZN(new_n429));
  NAND2_X1  g228(.A1(new_n429), .A2(KEYINPUT82), .ZN(new_n430));
  NAND3_X1  g229(.A1(new_n427), .A2(new_n430), .A3(new_n322), .ZN(new_n431));
  NAND2_X1  g230(.A1(new_n331), .A2(new_n429), .ZN(new_n432));
  NAND2_X1  g231(.A1(new_n431), .A2(new_n432), .ZN(new_n433));
  NAND2_X1  g232(.A1(G225gat), .A2(G233gat), .ZN(new_n434));
  INV_X1    g233(.A(new_n434), .ZN(new_n435));
  AOI21_X1  g234(.A(new_n406), .B1(new_n433), .B2(new_n435), .ZN(new_n436));
  NAND3_X1  g235(.A1(new_n427), .A2(new_n430), .A3(KEYINPUT3), .ZN(new_n437));
  INV_X1    g236(.A(KEYINPUT3), .ZN(new_n438));
  AOI21_X1  g237(.A(new_n331), .B1(new_n438), .B2(new_n429), .ZN(new_n439));
  NAND2_X1  g238(.A1(new_n437), .A2(new_n439), .ZN(new_n440));
  INV_X1    g239(.A(KEYINPUT4), .ZN(new_n441));
  OAI21_X1  g240(.A(new_n441), .B1(new_n322), .B2(new_n425), .ZN(new_n442));
  NAND3_X1  g241(.A1(new_n331), .A2(new_n429), .A3(KEYINPUT4), .ZN(new_n443));
  NAND4_X1  g242(.A1(new_n440), .A2(new_n442), .A3(new_n443), .A4(new_n434), .ZN(new_n444));
  NAND2_X1  g243(.A1(new_n436), .A2(new_n444), .ZN(new_n445));
  INV_X1    g244(.A(KEYINPUT83), .ZN(new_n446));
  AND3_X1   g245(.A1(new_n331), .A2(new_n429), .A3(KEYINPUT4), .ZN(new_n447));
  AOI21_X1  g246(.A(KEYINPUT4), .B1(new_n331), .B2(new_n429), .ZN(new_n448));
  OAI21_X1  g247(.A(new_n446), .B1(new_n447), .B2(new_n448), .ZN(new_n449));
  NAND3_X1  g248(.A1(new_n442), .A2(KEYINPUT83), .A3(new_n443), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n449), .A2(new_n450), .ZN(new_n451));
  NAND4_X1  g250(.A1(new_n451), .A2(new_n406), .A3(new_n434), .A4(new_n440), .ZN(new_n452));
  NAND2_X1  g251(.A1(new_n445), .A2(new_n452), .ZN(new_n453));
  XNOR2_X1  g252(.A(G1gat), .B(G29gat), .ZN(new_n454));
  XNOR2_X1  g253(.A(new_n454), .B(KEYINPUT0), .ZN(new_n455));
  XNOR2_X1  g254(.A(G57gat), .B(G85gat), .ZN(new_n456));
  XOR2_X1   g255(.A(new_n455), .B(new_n456), .Z(new_n457));
  INV_X1    g256(.A(new_n457), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n453), .A2(new_n458), .ZN(new_n459));
  INV_X1    g258(.A(KEYINPUT6), .ZN(new_n460));
  NAND3_X1  g259(.A1(new_n445), .A2(new_n452), .A3(new_n457), .ZN(new_n461));
  NAND3_X1  g260(.A1(new_n459), .A2(new_n460), .A3(new_n461), .ZN(new_n462));
  NAND3_X1  g261(.A1(new_n453), .A2(KEYINPUT6), .A3(new_n458), .ZN(new_n463));
  NAND2_X1  g262(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  NAND3_X1  g263(.A1(new_n401), .A2(new_n364), .A3(new_n403), .ZN(new_n465));
  XOR2_X1   g264(.A(KEYINPUT77), .B(KEYINPUT30), .Z(new_n466));
  AND3_X1   g265(.A1(new_n465), .A2(KEYINPUT78), .A3(new_n466), .ZN(new_n467));
  AOI21_X1  g266(.A(KEYINPUT78), .B1(new_n465), .B2(new_n466), .ZN(new_n468));
  OAI211_X1 g267(.A(new_n405), .B(new_n464), .C1(new_n467), .C2(new_n468), .ZN(new_n469));
  XNOR2_X1  g268(.A(KEYINPUT31), .B(G50gat), .ZN(new_n470));
  INV_X1    g269(.A(new_n470), .ZN(new_n471));
  NAND2_X1  g270(.A1(G228gat), .A2(G233gat), .ZN(new_n472));
  OAI21_X1  g271(.A(new_n438), .B1(new_n373), .B2(KEYINPUT29), .ZN(new_n473));
  AND2_X1   g272(.A1(new_n473), .A2(new_n425), .ZN(new_n474));
  NAND2_X1  g273(.A1(new_n429), .A2(new_n438), .ZN(new_n475));
  AOI21_X1  g274(.A(new_n394), .B1(new_n475), .B2(new_n384), .ZN(new_n476));
  OAI21_X1  g275(.A(new_n472), .B1(new_n474), .B2(new_n476), .ZN(new_n477));
  INV_X1    g276(.A(KEYINPUT85), .ZN(new_n478));
  AOI21_X1  g277(.A(new_n478), .B1(new_n475), .B2(new_n384), .ZN(new_n479));
  AOI211_X1 g278(.A(KEYINPUT85), .B(KEYINPUT29), .C1(new_n429), .C2(new_n438), .ZN(new_n480));
  NOR3_X1   g279(.A1(new_n479), .A2(new_n480), .A3(new_n394), .ZN(new_n481));
  NAND3_X1  g280(.A1(new_n427), .A2(new_n473), .A3(new_n430), .ZN(new_n482));
  NAND3_X1  g281(.A1(new_n482), .A2(G228gat), .A3(G233gat), .ZN(new_n483));
  OAI21_X1  g282(.A(new_n477), .B1(new_n481), .B2(new_n483), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n484), .A2(G22gat), .ZN(new_n485));
  XNOR2_X1  g284(.A(G78gat), .B(G106gat), .ZN(new_n486));
  XOR2_X1   g285(.A(new_n486), .B(KEYINPUT84), .Z(new_n487));
  INV_X1    g286(.A(new_n487), .ZN(new_n488));
  INV_X1    g287(.A(G22gat), .ZN(new_n489));
  OAI211_X1 g288(.A(new_n477), .B(new_n489), .C1(new_n481), .C2(new_n483), .ZN(new_n490));
  NAND3_X1  g289(.A1(new_n485), .A2(new_n488), .A3(new_n490), .ZN(new_n491));
  INV_X1    g290(.A(new_n491), .ZN(new_n492));
  AOI21_X1  g291(.A(new_n488), .B1(new_n485), .B2(new_n490), .ZN(new_n493));
  OAI21_X1  g292(.A(new_n471), .B1(new_n492), .B2(new_n493), .ZN(new_n494));
  NAND2_X1  g293(.A1(new_n485), .A2(new_n490), .ZN(new_n495));
  NAND2_X1  g294(.A1(new_n495), .A2(new_n487), .ZN(new_n496));
  NAND3_X1  g295(.A1(new_n496), .A2(new_n470), .A3(new_n491), .ZN(new_n497));
  NAND2_X1  g296(.A1(new_n494), .A2(new_n497), .ZN(new_n498));
  AOI21_X1  g297(.A(new_n360), .B1(new_n469), .B2(new_n498), .ZN(new_n499));
  AND2_X1   g298(.A1(new_n494), .A2(new_n497), .ZN(new_n500));
  NAND2_X1  g299(.A1(new_n400), .A2(new_n404), .ZN(new_n501));
  NAND2_X1  g300(.A1(new_n465), .A2(new_n466), .ZN(new_n502));
  INV_X1    g301(.A(KEYINPUT78), .ZN(new_n503));
  NAND2_X1  g302(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  NAND3_X1  g303(.A1(new_n465), .A2(KEYINPUT78), .A3(new_n466), .ZN(new_n505));
  AOI21_X1  g304(.A(new_n501), .B1(new_n504), .B2(new_n505), .ZN(new_n506));
  INV_X1    g305(.A(KEYINPUT39), .ZN(new_n507));
  AOI22_X1  g306(.A1(new_n449), .A2(new_n450), .B1(new_n437), .B2(new_n439), .ZN(new_n508));
  NOR3_X1   g307(.A1(new_n508), .A2(KEYINPUT86), .A3(new_n434), .ZN(new_n509));
  INV_X1    g308(.A(KEYINPUT86), .ZN(new_n510));
  NOR3_X1   g309(.A1(new_n447), .A2(new_n448), .A3(new_n446), .ZN(new_n511));
  AOI21_X1  g310(.A(KEYINPUT83), .B1(new_n442), .B2(new_n443), .ZN(new_n512));
  OAI21_X1  g311(.A(new_n440), .B1(new_n511), .B2(new_n512), .ZN(new_n513));
  AOI21_X1  g312(.A(new_n510), .B1(new_n513), .B2(new_n435), .ZN(new_n514));
  OAI21_X1  g313(.A(new_n507), .B1(new_n509), .B2(new_n514), .ZN(new_n515));
  NAND3_X1  g314(.A1(new_n431), .A2(new_n432), .A3(new_n434), .ZN(new_n516));
  AND3_X1   g315(.A1(new_n516), .A2(KEYINPUT87), .A3(KEYINPUT39), .ZN(new_n517));
  AOI21_X1  g316(.A(KEYINPUT87), .B1(new_n516), .B2(KEYINPUT39), .ZN(new_n518));
  NOR2_X1   g317(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  OAI21_X1  g318(.A(KEYINPUT86), .B1(new_n508), .B2(new_n434), .ZN(new_n520));
  NAND3_X1  g319(.A1(new_n513), .A2(new_n510), .A3(new_n435), .ZN(new_n521));
  NAND3_X1  g320(.A1(new_n519), .A2(new_n520), .A3(new_n521), .ZN(new_n522));
  NAND3_X1  g321(.A1(new_n515), .A2(new_n457), .A3(new_n522), .ZN(new_n523));
  INV_X1    g322(.A(KEYINPUT40), .ZN(new_n524));
  NAND2_X1  g323(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  NAND4_X1  g324(.A1(new_n515), .A2(KEYINPUT40), .A3(new_n457), .A4(new_n522), .ZN(new_n526));
  NAND3_X1  g325(.A1(new_n525), .A2(new_n459), .A3(new_n526), .ZN(new_n527));
  OAI21_X1  g326(.A(new_n500), .B1(new_n506), .B2(new_n527), .ZN(new_n528));
  INV_X1    g327(.A(new_n464), .ZN(new_n529));
  OAI21_X1  g328(.A(new_n394), .B1(new_n382), .B2(new_n386), .ZN(new_n530));
  INV_X1    g329(.A(KEYINPUT37), .ZN(new_n531));
  INV_X1    g330(.A(new_n390), .ZN(new_n532));
  AOI21_X1  g331(.A(new_n531), .B1(new_n532), .B2(new_n373), .ZN(new_n533));
  AOI211_X1 g332(.A(KEYINPUT38), .B(new_n364), .C1(new_n530), .C2(new_n533), .ZN(new_n534));
  NAND3_X1  g333(.A1(new_n401), .A2(new_n531), .A3(new_n403), .ZN(new_n535));
  NAND2_X1  g334(.A1(new_n534), .A2(new_n535), .ZN(new_n536));
  NAND3_X1  g335(.A1(new_n529), .A2(new_n536), .A3(new_n465), .ZN(new_n537));
  INV_X1    g336(.A(KEYINPUT88), .ZN(new_n538));
  AOI21_X1  g337(.A(new_n531), .B1(new_n401), .B2(new_n403), .ZN(new_n539));
  OAI21_X1  g338(.A(new_n538), .B1(new_n539), .B2(new_n364), .ZN(new_n540));
  OAI21_X1  g339(.A(KEYINPUT37), .B1(new_n393), .B2(new_n399), .ZN(new_n541));
  NAND3_X1  g340(.A1(new_n541), .A2(KEYINPUT88), .A3(new_n365), .ZN(new_n542));
  NAND3_X1  g341(.A1(new_n540), .A2(new_n542), .A3(new_n535), .ZN(new_n543));
  AOI21_X1  g342(.A(new_n537), .B1(new_n543), .B2(KEYINPUT38), .ZN(new_n544));
  OAI21_X1  g343(.A(new_n499), .B1(new_n528), .B2(new_n544), .ZN(new_n545));
  NAND2_X1  g344(.A1(new_n500), .A2(new_n356), .ZN(new_n546));
  OAI21_X1  g345(.A(KEYINPUT35), .B1(new_n546), .B2(new_n469), .ZN(new_n547));
  INV_X1    g346(.A(new_n356), .ZN(new_n548));
  NOR2_X1   g347(.A1(new_n498), .A2(new_n548), .ZN(new_n549));
  INV_X1    g348(.A(KEYINPUT35), .ZN(new_n550));
  NAND4_X1  g349(.A1(new_n506), .A2(new_n549), .A3(new_n550), .A4(new_n464), .ZN(new_n551));
  NAND2_X1  g350(.A1(new_n547), .A2(new_n551), .ZN(new_n552));
  AOI21_X1  g351(.A(new_n258), .B1(new_n545), .B2(new_n552), .ZN(new_n553));
  AOI21_X1  g352(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n554));
  XNOR2_X1  g353(.A(new_n554), .B(KEYINPUT94), .ZN(new_n555));
  XOR2_X1   g354(.A(G57gat), .B(G64gat), .Z(new_n556));
  NAND2_X1  g355(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  XOR2_X1   g356(.A(G71gat), .B(G78gat), .Z(new_n558));
  NAND2_X1  g357(.A1(new_n557), .A2(new_n558), .ZN(new_n559));
  INV_X1    g358(.A(G64gat), .ZN(new_n560));
  NAND2_X1  g359(.A1(new_n560), .A2(G57gat), .ZN(new_n561));
  XOR2_X1   g360(.A(KEYINPUT95), .B(G57gat), .Z(new_n562));
  OAI21_X1  g361(.A(new_n561), .B1(new_n562), .B2(new_n560), .ZN(new_n563));
  INV_X1    g362(.A(new_n558), .ZN(new_n564));
  NAND3_X1  g363(.A1(new_n563), .A2(new_n564), .A3(new_n555), .ZN(new_n565));
  NAND2_X1  g364(.A1(new_n559), .A2(new_n565), .ZN(new_n566));
  INV_X1    g365(.A(KEYINPUT21), .ZN(new_n567));
  NAND2_X1  g366(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  NAND2_X1  g367(.A1(G231gat), .A2(G233gat), .ZN(new_n569));
  XNOR2_X1  g368(.A(new_n568), .B(new_n569), .ZN(new_n570));
  XNOR2_X1  g369(.A(new_n570), .B(G127gat), .ZN(new_n571));
  OAI21_X1  g370(.A(new_n229), .B1(new_n567), .B2(new_n566), .ZN(new_n572));
  OR2_X1    g371(.A1(new_n571), .A2(new_n572), .ZN(new_n573));
  NAND2_X1  g372(.A1(new_n571), .A2(new_n572), .ZN(new_n574));
  NAND2_X1  g373(.A1(new_n573), .A2(new_n574), .ZN(new_n575));
  XNOR2_X1  g374(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n576));
  XNOR2_X1  g375(.A(new_n576), .B(new_n417), .ZN(new_n577));
  XNOR2_X1  g376(.A(G183gat), .B(G211gat), .ZN(new_n578));
  XOR2_X1   g377(.A(new_n577), .B(new_n578), .Z(new_n579));
  INV_X1    g378(.A(new_n579), .ZN(new_n580));
  NAND2_X1  g379(.A1(new_n575), .A2(new_n580), .ZN(new_n581));
  NAND3_X1  g380(.A1(new_n573), .A2(new_n574), .A3(new_n579), .ZN(new_n582));
  NAND2_X1  g381(.A1(new_n581), .A2(new_n582), .ZN(new_n583));
  NAND2_X1  g382(.A1(G85gat), .A2(G92gat), .ZN(new_n584));
  XNOR2_X1  g383(.A(new_n584), .B(KEYINPUT7), .ZN(new_n585));
  NAND2_X1  g384(.A1(G99gat), .A2(G106gat), .ZN(new_n586));
  INV_X1    g385(.A(G85gat), .ZN(new_n587));
  INV_X1    g386(.A(G92gat), .ZN(new_n588));
  AOI22_X1  g387(.A1(KEYINPUT8), .A2(new_n586), .B1(new_n587), .B2(new_n588), .ZN(new_n589));
  NAND2_X1  g388(.A1(new_n585), .A2(new_n589), .ZN(new_n590));
  XOR2_X1   g389(.A(G99gat), .B(G106gat), .Z(new_n591));
  AND2_X1   g390(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  NOR2_X1   g391(.A1(new_n590), .A2(new_n591), .ZN(new_n593));
  NOR2_X1   g392(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  AND2_X1   g393(.A1(G232gat), .A2(G233gat), .ZN(new_n595));
  AOI22_X1  g394(.A1(new_n230), .A2(new_n594), .B1(KEYINPUT41), .B2(new_n595), .ZN(new_n596));
  INV_X1    g395(.A(new_n594), .ZN(new_n597));
  NAND2_X1  g396(.A1(new_n232), .A2(new_n597), .ZN(new_n598));
  NOR2_X1   g397(.A1(new_n230), .A2(new_n231), .ZN(new_n599));
  OAI21_X1  g398(.A(new_n596), .B1(new_n598), .B2(new_n599), .ZN(new_n600));
  XOR2_X1   g399(.A(G190gat), .B(G218gat), .Z(new_n601));
  XNOR2_X1  g400(.A(new_n601), .B(KEYINPUT96), .ZN(new_n602));
  NAND2_X1  g401(.A1(new_n600), .A2(new_n602), .ZN(new_n603));
  INV_X1    g402(.A(KEYINPUT98), .ZN(new_n604));
  NAND2_X1  g403(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  NAND3_X1  g404(.A1(new_n600), .A2(KEYINPUT98), .A3(new_n602), .ZN(new_n606));
  AND2_X1   g405(.A1(new_n605), .A2(new_n606), .ZN(new_n607));
  OR2_X1    g406(.A1(new_n600), .A2(new_n602), .ZN(new_n608));
  AND2_X1   g407(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  NOR2_X1   g408(.A1(new_n595), .A2(KEYINPUT41), .ZN(new_n610));
  XNOR2_X1  g409(.A(new_n610), .B(G134gat), .ZN(new_n611));
  XNOR2_X1  g410(.A(new_n611), .B(new_n418), .ZN(new_n612));
  NAND2_X1  g411(.A1(new_n605), .A2(new_n606), .ZN(new_n613));
  INV_X1    g412(.A(KEYINPUT97), .ZN(new_n614));
  OAI21_X1  g413(.A(new_n612), .B1(new_n613), .B2(new_n614), .ZN(new_n615));
  NAND2_X1  g414(.A1(new_n609), .A2(new_n615), .ZN(new_n616));
  NAND2_X1  g415(.A1(new_n607), .A2(new_n608), .ZN(new_n617));
  NAND2_X1  g416(.A1(new_n607), .A2(KEYINPUT97), .ZN(new_n618));
  NAND3_X1  g417(.A1(new_n617), .A2(new_n618), .A3(new_n612), .ZN(new_n619));
  NAND3_X1  g418(.A1(new_n583), .A2(new_n616), .A3(new_n619), .ZN(new_n620));
  NAND2_X1  g419(.A1(G230gat), .A2(G233gat), .ZN(new_n621));
  XNOR2_X1  g420(.A(new_n621), .B(KEYINPUT102), .ZN(new_n622));
  AND2_X1   g421(.A1(new_n559), .A2(new_n565), .ZN(new_n623));
  INV_X1    g422(.A(KEYINPUT99), .ZN(new_n624));
  AOI21_X1  g423(.A(new_n593), .B1(new_n592), .B2(new_n624), .ZN(new_n625));
  NAND2_X1  g424(.A1(new_n590), .A2(new_n591), .ZN(new_n626));
  NAND2_X1  g425(.A1(new_n626), .A2(KEYINPUT99), .ZN(new_n627));
  NAND3_X1  g426(.A1(new_n623), .A2(new_n625), .A3(new_n627), .ZN(new_n628));
  NAND2_X1  g427(.A1(new_n628), .A2(KEYINPUT100), .ZN(new_n629));
  INV_X1    g428(.A(KEYINPUT10), .ZN(new_n630));
  NAND2_X1  g429(.A1(new_n597), .A2(new_n566), .ZN(new_n631));
  INV_X1    g430(.A(KEYINPUT100), .ZN(new_n632));
  NAND4_X1  g431(.A1(new_n623), .A2(new_n625), .A3(new_n632), .A4(new_n627), .ZN(new_n633));
  NAND4_X1  g432(.A1(new_n629), .A2(new_n630), .A3(new_n631), .A4(new_n633), .ZN(new_n634));
  NAND3_X1  g433(.A1(new_n623), .A2(KEYINPUT10), .A3(new_n594), .ZN(new_n635));
  AOI21_X1  g434(.A(new_n622), .B1(new_n634), .B2(new_n635), .ZN(new_n636));
  INV_X1    g435(.A(new_n621), .ZN(new_n637));
  NAND3_X1  g436(.A1(new_n629), .A2(new_n631), .A3(new_n633), .ZN(new_n638));
  AOI21_X1  g437(.A(new_n636), .B1(new_n637), .B2(new_n638), .ZN(new_n639));
  XNOR2_X1  g438(.A(G120gat), .B(G148gat), .ZN(new_n640));
  XNOR2_X1  g439(.A(G176gat), .B(G204gat), .ZN(new_n641));
  XOR2_X1   g440(.A(new_n640), .B(new_n641), .Z(new_n642));
  OR2_X1    g441(.A1(new_n639), .A2(new_n642), .ZN(new_n643));
  NAND2_X1  g442(.A1(new_n634), .A2(new_n635), .ZN(new_n644));
  NAND2_X1  g443(.A1(new_n644), .A2(KEYINPUT101), .ZN(new_n645));
  INV_X1    g444(.A(KEYINPUT101), .ZN(new_n646));
  NAND3_X1  g445(.A1(new_n634), .A2(new_n646), .A3(new_n635), .ZN(new_n647));
  NAND3_X1  g446(.A1(new_n645), .A2(new_n621), .A3(new_n647), .ZN(new_n648));
  NAND2_X1  g447(.A1(new_n638), .A2(new_n637), .ZN(new_n649));
  NAND3_X1  g448(.A1(new_n648), .A2(new_n649), .A3(new_n642), .ZN(new_n650));
  NAND2_X1  g449(.A1(new_n643), .A2(new_n650), .ZN(new_n651));
  OR3_X1    g450(.A1(new_n620), .A2(KEYINPUT103), .A3(new_n651), .ZN(new_n652));
  OAI21_X1  g451(.A(KEYINPUT103), .B1(new_n620), .B2(new_n651), .ZN(new_n653));
  AND2_X1   g452(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  AND2_X1   g453(.A1(new_n553), .A2(new_n654), .ZN(new_n655));
  NAND2_X1  g454(.A1(new_n655), .A2(new_n529), .ZN(new_n656));
  XNOR2_X1  g455(.A(new_n656), .B(G1gat), .ZN(G1324gat));
  OAI21_X1  g456(.A(new_n405), .B1(new_n467), .B2(new_n468), .ZN(new_n658));
  AND3_X1   g457(.A1(new_n553), .A2(new_n658), .A3(new_n654), .ZN(new_n659));
  XOR2_X1   g458(.A(KEYINPUT16), .B(G8gat), .Z(new_n660));
  NAND2_X1  g459(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  INV_X1    g460(.A(G8gat), .ZN(new_n662));
  OAI21_X1  g461(.A(new_n661), .B1(new_n662), .B2(new_n659), .ZN(new_n663));
  MUX2_X1   g462(.A(new_n661), .B(new_n663), .S(KEYINPUT42), .Z(G1325gat));
  INV_X1    g463(.A(KEYINPUT105), .ZN(new_n665));
  AND3_X1   g464(.A1(new_n348), .A2(KEYINPUT36), .A3(new_n355), .ZN(new_n666));
  AOI21_X1  g465(.A(KEYINPUT36), .B1(new_n348), .B2(new_n355), .ZN(new_n667));
  OAI21_X1  g466(.A(new_n665), .B1(new_n666), .B2(new_n667), .ZN(new_n668));
  NAND3_X1  g467(.A1(new_n358), .A2(KEYINPUT105), .A3(new_n359), .ZN(new_n669));
  NAND2_X1  g468(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  AND3_X1   g469(.A1(new_n655), .A2(G15gat), .A3(new_n670), .ZN(new_n671));
  AOI21_X1  g470(.A(G15gat), .B1(new_n655), .B2(new_n356), .ZN(new_n672));
  OR2_X1    g471(.A1(new_n672), .A2(KEYINPUT104), .ZN(new_n673));
  NAND2_X1  g472(.A1(new_n672), .A2(KEYINPUT104), .ZN(new_n674));
  AOI21_X1  g473(.A(new_n671), .B1(new_n673), .B2(new_n674), .ZN(G1326gat));
  NAND2_X1  g474(.A1(new_n655), .A2(new_n498), .ZN(new_n676));
  NAND2_X1  g475(.A1(new_n676), .A2(KEYINPUT106), .ZN(new_n677));
  INV_X1    g476(.A(KEYINPUT106), .ZN(new_n678));
  NAND3_X1  g477(.A1(new_n655), .A2(new_n678), .A3(new_n498), .ZN(new_n679));
  NAND2_X1  g478(.A1(new_n677), .A2(new_n679), .ZN(new_n680));
  XNOR2_X1  g479(.A(KEYINPUT43), .B(G22gat), .ZN(new_n681));
  INV_X1    g480(.A(new_n681), .ZN(new_n682));
  XNOR2_X1  g481(.A(new_n680), .B(new_n682), .ZN(G1327gat));
  NAND2_X1  g482(.A1(new_n616), .A2(new_n619), .ZN(new_n684));
  INV_X1    g483(.A(new_n583), .ZN(new_n685));
  INV_X1    g484(.A(new_n651), .ZN(new_n686));
  AND4_X1   g485(.A1(new_n553), .A2(new_n684), .A3(new_n685), .A4(new_n686), .ZN(new_n687));
  NAND3_X1  g486(.A1(new_n687), .A2(new_n203), .A3(new_n529), .ZN(new_n688));
  XNOR2_X1  g487(.A(new_n688), .B(KEYINPUT45), .ZN(new_n689));
  NOR2_X1   g488(.A1(new_n528), .A2(new_n544), .ZN(new_n690));
  NAND2_X1  g489(.A1(new_n469), .A2(new_n498), .ZN(new_n691));
  NAND3_X1  g490(.A1(new_n691), .A2(new_n669), .A3(new_n668), .ZN(new_n692));
  OAI21_X1  g491(.A(new_n552), .B1(new_n690), .B2(new_n692), .ZN(new_n693));
  NAND2_X1  g492(.A1(new_n693), .A2(new_n684), .ZN(new_n694));
  INV_X1    g493(.A(KEYINPUT44), .ZN(new_n695));
  NAND2_X1  g494(.A1(new_n545), .A2(new_n552), .ZN(new_n696));
  INV_X1    g495(.A(new_n684), .ZN(new_n697));
  NOR2_X1   g496(.A1(new_n697), .A2(new_n695), .ZN(new_n698));
  AOI22_X1  g497(.A1(new_n694), .A2(new_n695), .B1(new_n696), .B2(new_n698), .ZN(new_n699));
  INV_X1    g498(.A(new_n253), .ZN(new_n700));
  NOR3_X1   g499(.A1(new_n583), .A2(new_n700), .A3(new_n651), .ZN(new_n701));
  AND2_X1   g500(.A1(new_n699), .A2(new_n701), .ZN(new_n702));
  AND2_X1   g501(.A1(new_n702), .A2(new_n529), .ZN(new_n703));
  OAI21_X1  g502(.A(new_n689), .B1(new_n203), .B2(new_n703), .ZN(G1328gat));
  NAND3_X1  g503(.A1(new_n687), .A2(new_n204), .A3(new_n658), .ZN(new_n705));
  XOR2_X1   g504(.A(new_n705), .B(KEYINPUT46), .Z(new_n706));
  NAND2_X1  g505(.A1(new_n702), .A2(new_n658), .ZN(new_n707));
  NAND2_X1  g506(.A1(new_n707), .A2(G36gat), .ZN(new_n708));
  NAND2_X1  g507(.A1(new_n706), .A2(new_n708), .ZN(G1329gat));
  NAND2_X1  g508(.A1(new_n543), .A2(KEYINPUT38), .ZN(new_n710));
  INV_X1    g509(.A(new_n537), .ZN(new_n711));
  NAND2_X1  g510(.A1(new_n710), .A2(new_n711), .ZN(new_n712));
  AND3_X1   g511(.A1(new_n525), .A2(new_n459), .A3(new_n526), .ZN(new_n713));
  AOI21_X1  g512(.A(new_n498), .B1(new_n658), .B2(new_n713), .ZN(new_n714));
  NAND2_X1  g513(.A1(new_n712), .A2(new_n714), .ZN(new_n715));
  AOI21_X1  g514(.A(new_n670), .B1(new_n469), .B2(new_n498), .ZN(new_n716));
  AOI22_X1  g515(.A1(new_n715), .A2(new_n716), .B1(new_n547), .B2(new_n551), .ZN(new_n717));
  OAI21_X1  g516(.A(new_n695), .B1(new_n717), .B2(new_n697), .ZN(new_n718));
  NAND2_X1  g517(.A1(new_n696), .A2(new_n698), .ZN(new_n719));
  NAND4_X1  g518(.A1(new_n718), .A2(new_n670), .A3(new_n719), .A4(new_n701), .ZN(new_n720));
  INV_X1    g519(.A(KEYINPUT107), .ZN(new_n721));
  AND2_X1   g520(.A1(new_n720), .A2(new_n721), .ZN(new_n722));
  NOR2_X1   g521(.A1(new_n720), .A2(new_n721), .ZN(new_n723));
  INV_X1    g522(.A(G43gat), .ZN(new_n724));
  NOR3_X1   g523(.A1(new_n722), .A2(new_n723), .A3(new_n724), .ZN(new_n725));
  NAND3_X1  g524(.A1(new_n687), .A2(new_n724), .A3(new_n356), .ZN(new_n726));
  NAND2_X1  g525(.A1(new_n726), .A2(KEYINPUT47), .ZN(new_n727));
  NAND2_X1  g526(.A1(new_n720), .A2(G43gat), .ZN(new_n728));
  AND2_X1   g527(.A1(new_n728), .A2(new_n726), .ZN(new_n729));
  OAI22_X1  g528(.A1(new_n725), .A2(new_n727), .B1(new_n729), .B2(KEYINPUT47), .ZN(G1330gat));
  NAND4_X1  g529(.A1(new_n718), .A2(new_n498), .A3(new_n719), .A4(new_n701), .ZN(new_n731));
  NAND2_X1  g530(.A1(new_n731), .A2(KEYINPUT108), .ZN(new_n732));
  NAND2_X1  g531(.A1(new_n732), .A2(G50gat), .ZN(new_n733));
  NOR2_X1   g532(.A1(new_n731), .A2(KEYINPUT108), .ZN(new_n734));
  NOR2_X1   g533(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  INV_X1    g534(.A(G50gat), .ZN(new_n736));
  NAND3_X1  g535(.A1(new_n687), .A2(new_n736), .A3(new_n498), .ZN(new_n737));
  NAND2_X1  g536(.A1(new_n737), .A2(KEYINPUT48), .ZN(new_n738));
  NAND2_X1  g537(.A1(new_n731), .A2(G50gat), .ZN(new_n739));
  AND2_X1   g538(.A1(new_n739), .A2(new_n737), .ZN(new_n740));
  OAI22_X1  g539(.A1(new_n735), .A2(new_n738), .B1(KEYINPUT48), .B2(new_n740), .ZN(G1331gat));
  INV_X1    g540(.A(new_n620), .ZN(new_n742));
  NAND3_X1  g541(.A1(new_n742), .A2(new_n700), .A3(new_n651), .ZN(new_n743));
  OR3_X1    g542(.A1(new_n717), .A2(KEYINPUT109), .A3(new_n743), .ZN(new_n744));
  OAI21_X1  g543(.A(KEYINPUT109), .B1(new_n717), .B2(new_n743), .ZN(new_n745));
  NAND2_X1  g544(.A1(new_n744), .A2(new_n745), .ZN(new_n746));
  INV_X1    g545(.A(new_n746), .ZN(new_n747));
  NAND2_X1  g546(.A1(new_n747), .A2(new_n529), .ZN(new_n748));
  XNOR2_X1  g547(.A(new_n748), .B(new_n562), .ZN(G1332gat));
  NAND2_X1  g548(.A1(new_n747), .A2(new_n658), .ZN(new_n750));
  OAI21_X1  g549(.A(new_n750), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n751));
  XOR2_X1   g550(.A(KEYINPUT49), .B(G64gat), .Z(new_n752));
  OAI21_X1  g551(.A(new_n751), .B1(new_n750), .B2(new_n752), .ZN(G1333gat));
  NAND3_X1  g552(.A1(new_n744), .A2(new_n670), .A3(new_n745), .ZN(new_n754));
  NAND2_X1  g553(.A1(new_n754), .A2(G71gat), .ZN(new_n755));
  OR2_X1    g554(.A1(new_n548), .A2(G71gat), .ZN(new_n756));
  OAI21_X1  g555(.A(new_n755), .B1(new_n746), .B2(new_n756), .ZN(new_n757));
  INV_X1    g556(.A(KEYINPUT50), .ZN(new_n758));
  NAND2_X1  g557(.A1(new_n757), .A2(new_n758), .ZN(new_n759));
  OAI211_X1 g558(.A(new_n755), .B(KEYINPUT50), .C1(new_n746), .C2(new_n756), .ZN(new_n760));
  NAND2_X1  g559(.A1(new_n759), .A2(new_n760), .ZN(G1334gat));
  NAND2_X1  g560(.A1(new_n747), .A2(new_n498), .ZN(new_n762));
  XNOR2_X1  g561(.A(new_n762), .B(G78gat), .ZN(G1335gat));
  NAND2_X1  g562(.A1(new_n685), .A2(new_n700), .ZN(new_n764));
  NOR2_X1   g563(.A1(new_n764), .A2(new_n686), .ZN(new_n765));
  AND2_X1   g564(.A1(new_n699), .A2(new_n765), .ZN(new_n766));
  AOI21_X1  g565(.A(new_n587), .B1(new_n766), .B2(new_n529), .ZN(new_n767));
  INV_X1    g566(.A(KEYINPUT51), .ZN(new_n768));
  AOI21_X1  g567(.A(new_n764), .B1(KEYINPUT110), .B2(new_n768), .ZN(new_n769));
  NAND3_X1  g568(.A1(new_n693), .A2(new_n684), .A3(new_n769), .ZN(new_n770));
  NOR2_X1   g569(.A1(new_n768), .A2(KEYINPUT110), .ZN(new_n771));
  NAND2_X1  g570(.A1(new_n770), .A2(new_n771), .ZN(new_n772));
  INV_X1    g571(.A(new_n771), .ZN(new_n773));
  NAND4_X1  g572(.A1(new_n693), .A2(new_n684), .A3(new_n769), .A4(new_n773), .ZN(new_n774));
  NAND3_X1  g573(.A1(new_n772), .A2(new_n651), .A3(new_n774), .ZN(new_n775));
  NOR3_X1   g574(.A1(new_n775), .A2(G85gat), .A3(new_n464), .ZN(new_n776));
  OR2_X1    g575(.A1(new_n767), .A2(new_n776), .ZN(G1336gat));
  NAND4_X1  g576(.A1(new_n718), .A2(new_n658), .A3(new_n719), .A4(new_n765), .ZN(new_n778));
  NAND2_X1  g577(.A1(new_n778), .A2(G92gat), .ZN(new_n779));
  NAND2_X1  g578(.A1(new_n779), .A2(KEYINPUT111), .ZN(new_n780));
  NOR2_X1   g579(.A1(new_n506), .A2(G92gat), .ZN(new_n781));
  NAND4_X1  g580(.A1(new_n772), .A2(new_n651), .A3(new_n774), .A4(new_n781), .ZN(new_n782));
  NAND2_X1  g581(.A1(new_n779), .A2(new_n782), .ZN(new_n783));
  INV_X1    g582(.A(KEYINPUT52), .ZN(new_n784));
  NAND3_X1  g583(.A1(new_n780), .A2(new_n783), .A3(new_n784), .ZN(new_n785));
  OAI211_X1 g584(.A(new_n779), .B(new_n782), .C1(KEYINPUT111), .C2(KEYINPUT52), .ZN(new_n786));
  AND2_X1   g585(.A1(new_n785), .A2(new_n786), .ZN(G1337gat));
  NAND2_X1  g586(.A1(new_n766), .A2(new_n670), .ZN(new_n788));
  NAND2_X1  g587(.A1(new_n788), .A2(G99gat), .ZN(new_n789));
  OR2_X1    g588(.A1(new_n548), .A2(G99gat), .ZN(new_n790));
  OAI21_X1  g589(.A(new_n789), .B1(new_n775), .B2(new_n790), .ZN(G1338gat));
  NOR3_X1   g590(.A1(new_n500), .A2(new_n686), .A3(G106gat), .ZN(new_n792));
  NAND3_X1  g591(.A1(new_n772), .A2(new_n774), .A3(new_n792), .ZN(new_n793));
  INV_X1    g592(.A(KEYINPUT112), .ZN(new_n794));
  NAND2_X1  g593(.A1(new_n793), .A2(new_n794), .ZN(new_n795));
  NAND4_X1  g594(.A1(new_n772), .A2(KEYINPUT112), .A3(new_n774), .A4(new_n792), .ZN(new_n796));
  NAND2_X1  g595(.A1(new_n795), .A2(new_n796), .ZN(new_n797));
  NAND4_X1  g596(.A1(new_n699), .A2(KEYINPUT113), .A3(new_n498), .A4(new_n765), .ZN(new_n798));
  NAND4_X1  g597(.A1(new_n718), .A2(new_n498), .A3(new_n719), .A4(new_n765), .ZN(new_n799));
  INV_X1    g598(.A(KEYINPUT113), .ZN(new_n800));
  NAND2_X1  g599(.A1(new_n799), .A2(new_n800), .ZN(new_n801));
  NAND3_X1  g600(.A1(new_n798), .A2(new_n801), .A3(G106gat), .ZN(new_n802));
  INV_X1    g601(.A(KEYINPUT53), .ZN(new_n803));
  NAND3_X1  g602(.A1(new_n797), .A2(new_n802), .A3(new_n803), .ZN(new_n804));
  NAND2_X1  g603(.A1(new_n799), .A2(G106gat), .ZN(new_n805));
  NAND2_X1  g604(.A1(new_n805), .A2(new_n793), .ZN(new_n806));
  NAND2_X1  g605(.A1(new_n806), .A2(KEYINPUT53), .ZN(new_n807));
  NAND2_X1  g606(.A1(new_n804), .A2(new_n807), .ZN(G1339gat));
  NAND3_X1  g607(.A1(new_n634), .A2(new_n622), .A3(new_n635), .ZN(new_n809));
  XNOR2_X1  g608(.A(new_n809), .B(KEYINPUT114), .ZN(new_n810));
  NAND3_X1  g609(.A1(new_n810), .A2(new_n648), .A3(KEYINPUT54), .ZN(new_n811));
  INV_X1    g610(.A(KEYINPUT54), .ZN(new_n812));
  AOI21_X1  g611(.A(new_n642), .B1(new_n636), .B2(new_n812), .ZN(new_n813));
  NAND2_X1  g612(.A1(new_n811), .A2(new_n813), .ZN(new_n814));
  INV_X1    g613(.A(KEYINPUT55), .ZN(new_n815));
  NAND2_X1  g614(.A1(new_n814), .A2(new_n815), .ZN(new_n816));
  NAND3_X1  g615(.A1(new_n811), .A2(KEYINPUT55), .A3(new_n813), .ZN(new_n817));
  NAND4_X1  g616(.A1(new_n816), .A2(new_n253), .A3(new_n650), .A4(new_n817), .ZN(new_n818));
  NOR2_X1   g617(.A1(new_n239), .A2(new_n240), .ZN(new_n819));
  AOI21_X1  g618(.A(new_n234), .B1(new_n233), .B2(new_n235), .ZN(new_n820));
  OAI21_X1  g619(.A(new_n248), .B1(new_n819), .B2(new_n820), .ZN(new_n821));
  AND2_X1   g620(.A1(new_n252), .A2(new_n821), .ZN(new_n822));
  NAND2_X1  g621(.A1(new_n651), .A2(new_n822), .ZN(new_n823));
  AOI21_X1  g622(.A(new_n684), .B1(new_n818), .B2(new_n823), .ZN(new_n824));
  NAND3_X1  g623(.A1(new_n816), .A2(new_n650), .A3(new_n817), .ZN(new_n825));
  NAND2_X1  g624(.A1(new_n684), .A2(new_n822), .ZN(new_n826));
  NOR2_X1   g625(.A1(new_n825), .A2(new_n826), .ZN(new_n827));
  OAI21_X1  g626(.A(new_n685), .B1(new_n824), .B2(new_n827), .ZN(new_n828));
  NAND3_X1  g627(.A1(new_n742), .A2(new_n700), .A3(new_n686), .ZN(new_n829));
  AOI21_X1  g628(.A(new_n498), .B1(new_n828), .B2(new_n829), .ZN(new_n830));
  NAND2_X1  g629(.A1(new_n506), .A2(new_n529), .ZN(new_n831));
  NOR2_X1   g630(.A1(new_n831), .A2(new_n548), .ZN(new_n832));
  NAND2_X1  g631(.A1(new_n830), .A2(new_n832), .ZN(new_n833));
  INV_X1    g632(.A(G113gat), .ZN(new_n834));
  NOR3_X1   g633(.A1(new_n833), .A2(new_n834), .A3(new_n258), .ZN(new_n835));
  AOI21_X1  g634(.A(new_n464), .B1(new_n828), .B2(new_n829), .ZN(new_n836));
  NAND2_X1  g635(.A1(new_n506), .A2(new_n549), .ZN(new_n837));
  INV_X1    g636(.A(new_n837), .ZN(new_n838));
  NAND2_X1  g637(.A1(new_n836), .A2(new_n838), .ZN(new_n839));
  INV_X1    g638(.A(new_n839), .ZN(new_n840));
  NAND2_X1  g639(.A1(new_n840), .A2(new_n253), .ZN(new_n841));
  AOI21_X1  g640(.A(new_n835), .B1(new_n834), .B2(new_n841), .ZN(G1340gat));
  NOR3_X1   g641(.A1(new_n833), .A2(new_n311), .A3(new_n686), .ZN(new_n843));
  NAND2_X1  g642(.A1(new_n840), .A2(new_n651), .ZN(new_n844));
  AOI21_X1  g643(.A(new_n843), .B1(new_n311), .B2(new_n844), .ZN(G1341gat));
  AOI21_X1  g644(.A(G127gat), .B1(new_n840), .B2(new_n583), .ZN(new_n846));
  NAND4_X1  g645(.A1(new_n830), .A2(G127gat), .A3(new_n583), .A4(new_n832), .ZN(new_n847));
  AND2_X1   g646(.A1(new_n847), .A2(KEYINPUT115), .ZN(new_n848));
  NOR2_X1   g647(.A1(new_n847), .A2(KEYINPUT115), .ZN(new_n849));
  NOR3_X1   g648(.A1(new_n846), .A2(new_n848), .A3(new_n849), .ZN(G1342gat));
  AOI211_X1 g649(.A(G134gat), .B(new_n697), .C1(KEYINPUT116), .C2(KEYINPUT56), .ZN(new_n851));
  NAND3_X1  g650(.A1(new_n836), .A2(new_n838), .A3(new_n851), .ZN(new_n852));
  NOR2_X1   g651(.A1(KEYINPUT116), .A2(KEYINPUT56), .ZN(new_n853));
  XNOR2_X1  g652(.A(new_n852), .B(new_n853), .ZN(new_n854));
  NAND3_X1  g653(.A1(new_n830), .A2(new_n684), .A3(new_n832), .ZN(new_n855));
  AOI21_X1  g654(.A(KEYINPUT117), .B1(new_n855), .B2(G134gat), .ZN(new_n856));
  AND3_X1   g655(.A1(new_n855), .A2(KEYINPUT117), .A3(G134gat), .ZN(new_n857));
  OAI21_X1  g656(.A(new_n854), .B1(new_n856), .B2(new_n857), .ZN(new_n858));
  NAND2_X1  g657(.A1(new_n858), .A2(KEYINPUT118), .ZN(new_n859));
  INV_X1    g658(.A(KEYINPUT118), .ZN(new_n860));
  OAI211_X1 g659(.A(new_n854), .B(new_n860), .C1(new_n856), .C2(new_n857), .ZN(new_n861));
  NAND2_X1  g660(.A1(new_n859), .A2(new_n861), .ZN(G1343gat));
  XNOR2_X1  g661(.A(KEYINPUT121), .B(KEYINPUT58), .ZN(new_n863));
  NOR2_X1   g662(.A1(new_n670), .A2(new_n500), .ZN(new_n864));
  NAND2_X1  g663(.A1(new_n836), .A2(new_n864), .ZN(new_n865));
  OR2_X1    g664(.A1(new_n865), .A2(KEYINPUT120), .ZN(new_n866));
  NAND2_X1  g665(.A1(new_n865), .A2(KEYINPUT120), .ZN(new_n867));
  NAND3_X1  g666(.A1(new_n866), .A2(new_n506), .A3(new_n867), .ZN(new_n868));
  OR2_X1    g667(.A1(new_n258), .A2(G141gat), .ZN(new_n869));
  OAI21_X1  g668(.A(new_n863), .B1(new_n868), .B2(new_n869), .ZN(new_n870));
  NOR2_X1   g669(.A1(new_n831), .A2(new_n670), .ZN(new_n871));
  NAND2_X1  g670(.A1(new_n498), .A2(KEYINPUT57), .ZN(new_n872));
  NAND4_X1  g671(.A1(new_n816), .A2(new_n257), .A3(new_n650), .A4(new_n817), .ZN(new_n873));
  AOI21_X1  g672(.A(new_n684), .B1(new_n873), .B2(new_n823), .ZN(new_n874));
  OAI21_X1  g673(.A(new_n685), .B1(new_n874), .B2(new_n827), .ZN(new_n875));
  AOI21_X1  g674(.A(new_n872), .B1(new_n875), .B2(new_n829), .ZN(new_n876));
  AOI21_X1  g675(.A(new_n500), .B1(new_n828), .B2(new_n829), .ZN(new_n877));
  OAI22_X1  g676(.A1(KEYINPUT119), .A2(new_n876), .B1(new_n877), .B2(KEYINPUT57), .ZN(new_n878));
  AND2_X1   g677(.A1(new_n876), .A2(KEYINPUT119), .ZN(new_n879));
  OAI211_X1 g678(.A(new_n257), .B(new_n871), .C1(new_n878), .C2(new_n879), .ZN(new_n880));
  AND2_X1   g679(.A1(new_n880), .A2(new_n407), .ZN(new_n881));
  NOR3_X1   g680(.A1(new_n865), .A2(new_n658), .A3(new_n869), .ZN(new_n882));
  OAI211_X1 g681(.A(new_n253), .B(new_n871), .C1(new_n878), .C2(new_n879), .ZN(new_n883));
  AOI21_X1  g682(.A(new_n882), .B1(new_n883), .B2(new_n407), .ZN(new_n884));
  INV_X1    g683(.A(KEYINPUT58), .ZN(new_n885));
  OAI22_X1  g684(.A1(new_n870), .A2(new_n881), .B1(new_n884), .B2(new_n885), .ZN(G1344gat));
  INV_X1    g685(.A(KEYINPUT122), .ZN(new_n887));
  NOR3_X1   g686(.A1(new_n831), .A2(new_n670), .A3(new_n686), .ZN(new_n888));
  NAND3_X1  g687(.A1(new_n652), .A2(new_n258), .A3(new_n653), .ZN(new_n889));
  NAND2_X1  g688(.A1(new_n875), .A2(new_n889), .ZN(new_n890));
  AOI21_X1  g689(.A(KEYINPUT57), .B1(new_n890), .B2(new_n498), .ZN(new_n891));
  AOI21_X1  g690(.A(new_n872), .B1(new_n828), .B2(new_n829), .ZN(new_n892));
  OAI211_X1 g691(.A(new_n887), .B(new_n888), .C1(new_n891), .C2(new_n892), .ZN(new_n893));
  NAND2_X1  g692(.A1(new_n893), .A2(G148gat), .ZN(new_n894));
  AND2_X1   g693(.A1(new_n828), .A2(new_n829), .ZN(new_n895));
  AOI21_X1  g694(.A(new_n500), .B1(new_n875), .B2(new_n889), .ZN(new_n896));
  OAI22_X1  g695(.A1(new_n895), .A2(new_n872), .B1(new_n896), .B2(KEYINPUT57), .ZN(new_n897));
  AOI21_X1  g696(.A(new_n887), .B1(new_n897), .B2(new_n888), .ZN(new_n898));
  OAI21_X1  g697(.A(KEYINPUT59), .B1(new_n894), .B2(new_n898), .ZN(new_n899));
  NOR2_X1   g698(.A1(new_n408), .A2(KEYINPUT59), .ZN(new_n900));
  OAI21_X1  g699(.A(new_n871), .B1(new_n878), .B2(new_n879), .ZN(new_n901));
  OAI21_X1  g700(.A(new_n900), .B1(new_n901), .B2(new_n686), .ZN(new_n902));
  NAND2_X1  g701(.A1(new_n899), .A2(new_n902), .ZN(new_n903));
  INV_X1    g702(.A(new_n868), .ZN(new_n904));
  NAND3_X1  g703(.A1(new_n904), .A2(new_n408), .A3(new_n651), .ZN(new_n905));
  NAND2_X1  g704(.A1(new_n903), .A2(new_n905), .ZN(G1345gat));
  OAI21_X1  g705(.A(G155gat), .B1(new_n901), .B2(new_n685), .ZN(new_n907));
  NAND2_X1  g706(.A1(new_n583), .A2(new_n417), .ZN(new_n908));
  OAI21_X1  g707(.A(new_n907), .B1(new_n868), .B2(new_n908), .ZN(G1346gat));
  OR3_X1    g708(.A1(new_n901), .A2(new_n418), .A3(new_n697), .ZN(new_n910));
  OAI21_X1  g709(.A(new_n418), .B1(new_n868), .B2(new_n697), .ZN(new_n911));
  AND2_X1   g710(.A1(new_n910), .A2(new_n911), .ZN(G1347gat));
  NAND2_X1  g711(.A1(new_n658), .A2(new_n464), .ZN(new_n913));
  NOR2_X1   g712(.A1(new_n913), .A2(new_n548), .ZN(new_n914));
  NAND2_X1  g713(.A1(new_n830), .A2(new_n914), .ZN(new_n915));
  INV_X1    g714(.A(G169gat), .ZN(new_n916));
  NOR3_X1   g715(.A1(new_n915), .A2(new_n916), .A3(new_n258), .ZN(new_n917));
  AOI21_X1  g716(.A(new_n529), .B1(new_n828), .B2(new_n829), .ZN(new_n918));
  AND3_X1   g717(.A1(new_n918), .A2(new_n658), .A3(new_n549), .ZN(new_n919));
  NAND2_X1  g718(.A1(new_n919), .A2(new_n253), .ZN(new_n920));
  AOI21_X1  g719(.A(new_n917), .B1(new_n916), .B2(new_n920), .ZN(G1348gat));
  INV_X1    g720(.A(G176gat), .ZN(new_n922));
  NAND3_X1  g721(.A1(new_n919), .A2(new_n922), .A3(new_n651), .ZN(new_n923));
  OAI21_X1  g722(.A(G176gat), .B1(new_n915), .B2(new_n686), .ZN(new_n924));
  NAND2_X1  g723(.A1(new_n923), .A2(new_n924), .ZN(G1349gat));
  OAI21_X1  g724(.A(G183gat), .B1(new_n915), .B2(new_n685), .ZN(new_n926));
  AND2_X1   g725(.A1(new_n583), .A2(new_n272), .ZN(new_n927));
  AND3_X1   g726(.A1(new_n919), .A2(KEYINPUT123), .A3(new_n927), .ZN(new_n928));
  AOI21_X1  g727(.A(KEYINPUT123), .B1(new_n919), .B2(new_n927), .ZN(new_n929));
  OAI21_X1  g728(.A(new_n926), .B1(new_n928), .B2(new_n929), .ZN(new_n930));
  NAND2_X1  g729(.A1(new_n930), .A2(KEYINPUT60), .ZN(new_n931));
  INV_X1    g730(.A(KEYINPUT60), .ZN(new_n932));
  OAI211_X1 g731(.A(new_n932), .B(new_n926), .C1(new_n928), .C2(new_n929), .ZN(new_n933));
  NAND2_X1  g732(.A1(new_n931), .A2(new_n933), .ZN(G1350gat));
  NAND3_X1  g733(.A1(new_n919), .A2(new_n267), .A3(new_n684), .ZN(new_n935));
  NAND3_X1  g734(.A1(new_n830), .A2(new_n684), .A3(new_n914), .ZN(new_n936));
  NOR2_X1   g735(.A1(KEYINPUT124), .A2(KEYINPUT61), .ZN(new_n937));
  AOI21_X1  g736(.A(new_n267), .B1(KEYINPUT124), .B2(KEYINPUT61), .ZN(new_n938));
  AND3_X1   g737(.A1(new_n936), .A2(new_n937), .A3(new_n938), .ZN(new_n939));
  AOI21_X1  g738(.A(new_n937), .B1(new_n936), .B2(new_n938), .ZN(new_n940));
  OAI21_X1  g739(.A(new_n935), .B1(new_n939), .B2(new_n940), .ZN(G1351gat));
  NOR3_X1   g740(.A1(new_n670), .A2(new_n506), .A3(new_n500), .ZN(new_n942));
  NAND2_X1  g741(.A1(new_n918), .A2(new_n942), .ZN(new_n943));
  XNOR2_X1  g742(.A(new_n943), .B(KEYINPUT125), .ZN(new_n944));
  AOI21_X1  g743(.A(G197gat), .B1(new_n944), .B2(new_n253), .ZN(new_n945));
  OR2_X1    g744(.A1(new_n913), .A2(new_n670), .ZN(new_n946));
  XNOR2_X1  g745(.A(new_n946), .B(KEYINPUT126), .ZN(new_n947));
  NAND2_X1  g746(.A1(new_n897), .A2(new_n947), .ZN(new_n948));
  INV_X1    g747(.A(new_n948), .ZN(new_n949));
  AND2_X1   g748(.A1(new_n257), .A2(G197gat), .ZN(new_n950));
  AOI21_X1  g749(.A(new_n945), .B1(new_n949), .B2(new_n950), .ZN(G1352gat));
  NOR3_X1   g750(.A1(new_n943), .A2(G204gat), .A3(new_n686), .ZN(new_n952));
  XNOR2_X1  g751(.A(new_n952), .B(KEYINPUT62), .ZN(new_n953));
  OAI21_X1  g752(.A(G204gat), .B1(new_n948), .B2(new_n686), .ZN(new_n954));
  NAND2_X1  g753(.A1(new_n953), .A2(new_n954), .ZN(G1353gat));
  NAND3_X1  g754(.A1(new_n944), .A2(new_n368), .A3(new_n583), .ZN(new_n956));
  NOR2_X1   g755(.A1(new_n946), .A2(new_n685), .ZN(new_n957));
  NAND2_X1  g756(.A1(new_n897), .A2(new_n957), .ZN(new_n958));
  AND3_X1   g757(.A1(new_n958), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n959));
  AOI21_X1  g758(.A(KEYINPUT63), .B1(new_n958), .B2(G211gat), .ZN(new_n960));
  OAI21_X1  g759(.A(new_n956), .B1(new_n959), .B2(new_n960), .ZN(G1354gat));
  NAND3_X1  g760(.A1(new_n944), .A2(new_n369), .A3(new_n684), .ZN(new_n962));
  NAND2_X1  g761(.A1(new_n948), .A2(KEYINPUT127), .ZN(new_n963));
  INV_X1    g762(.A(KEYINPUT127), .ZN(new_n964));
  NAND3_X1  g763(.A1(new_n897), .A2(new_n964), .A3(new_n947), .ZN(new_n965));
  AND3_X1   g764(.A1(new_n963), .A2(new_n684), .A3(new_n965), .ZN(new_n966));
  OAI21_X1  g765(.A(new_n962), .B1(new_n966), .B2(new_n369), .ZN(G1355gat));
endmodule


