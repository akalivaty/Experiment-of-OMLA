

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n524, n525, n526, n527,
         n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538,
         n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549,
         n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560,
         n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571,
         n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582,
         n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593,
         n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604,
         n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615,
         n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626,
         n627, n628, n629, n630, n631, n632, n633, n634, n635, n636, n637,
         n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, n648,
         n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659,
         n660, n661, n662, n663, n664, n665, n666, n667, n668, n669, n670,
         n671, n672, n673, n674, n675, n676, n677, n678, n679, n680, n681,
         n682, n683, n684, n685, n686, n687, n688, n689, n690, n691, n692,
         n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, n703,
         n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, n714,
         n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, n725,
         n726, n727, n728, n729, n730, n731, n732, n733, n734, n735, n736,
         n737, n738, n739, n740, n741, n742, n743, n744, n745, n746, n747,
         n748, n749, n750, n751, n752, n753, n754, n755, n756, n757, n758,
         n759, n760, n761, n762, n763, n764, n765, n766, n767, n768, n769,
         n770, n771, n772, n773, n774, n775, n776, n777, n778, n779, n780,
         n781, n782, n783, n784, n785, n786, n787, n788, n789, n790, n791,
         n792, n793, n794, n795, n796, n797, n798, n799, n800, n801, n802,
         n803, n804, n805, n806, n807, n808, n809, n810, n811, n812, n813,
         n814, n815, n816, n817, n818, n819, n820, n821, n822, n823, n824,
         n825, n826, n827, n828, n829, n830, n831, n832, n833, n834, n835,
         n836, n837, n838, n839, n840, n841, n842, n843, n844, n845, n846,
         n847, n848, n849, n850, n851, n852, n853, n854, n855, n856, n857,
         n858, n859, n860, n861, n862, n863, n864, n865, n866, n867, n868,
         n869, n870, n871, n872, n873, n874, n875, n876, n877, n878, n879,
         n880, n881, n882, n883, n884, n885, n886, n887, n888, n889, n890,
         n891, n892, n893, n894, n895, n896, n897, n898, n899, n900, n901,
         n902, n903, n904, n905, n906, n907, n908, n909, n910, n911, n912,
         n913, n914, n915, n916, n917, n918, n919, n920, n921, n922, n923,
         n924, n925, n926, n927, n928, n929, n930, n931, n932, n933, n934,
         n935, n936, n937, n938, n939, n940, n941, n942, n943, n944, n945,
         n946, n947, n948, n949, n950, n951, n952, n953, n954, n955, n956,
         n957, n958, n959, n960, n961, n962, n963, n964, n965, n966, n967,
         n968, n969, n970, n971, n972, n973, n974, n975, n976, n977, n978,
         n979, n980, n981, n982, n983, n984, n985, n986, n987, n988, n989,
         n990, n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000,
         n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010,
         n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020,
         n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030,
         n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NOR2_X1 U557 ( .A1(n532), .A2(n531), .ZN(n533) );
  NOR2_X1 U558 ( .A1(n762), .A2(n761), .ZN(n524) );
  XNOR2_X1 U559 ( .A(n528), .B(KEYINPUT23), .ZN(n532) );
  NOR2_X1 U560 ( .A1(G651), .A2(n652), .ZN(n647) );
  XNOR2_X1 U561 ( .A(n538), .B(KEYINPUT66), .ZN(G160) );
  NOR2_X1 U562 ( .A1(G2105), .A2(G2104), .ZN(n525) );
  XOR2_X1 U563 ( .A(KEYINPUT17), .B(n525), .Z(n1001) );
  NAND2_X1 U564 ( .A1(n1001), .A2(G137), .ZN(n526) );
  XOR2_X1 U565 ( .A(KEYINPUT71), .B(n526), .Z(n537) );
  XNOR2_X1 U566 ( .A(G2104), .B(KEYINPUT67), .ZN(n529) );
  NOR2_X2 U567 ( .A1(G2105), .A2(n529), .ZN(n527) );
  XOR2_X2 U568 ( .A(KEYINPUT69), .B(n527), .Z(n1003) );
  NAND2_X1 U569 ( .A1(n1003), .A2(G101), .ZN(n528) );
  AND2_X1 U570 ( .A1(n529), .A2(G2105), .ZN(n997) );
  NAND2_X1 U571 ( .A1(n997), .A2(G125), .ZN(n530) );
  XOR2_X1 U572 ( .A(KEYINPUT68), .B(n530), .Z(n531) );
  XNOR2_X1 U573 ( .A(n533), .B(KEYINPUT70), .ZN(n535) );
  AND2_X1 U574 ( .A1(G2105), .A2(G2104), .ZN(n998) );
  NAND2_X1 U575 ( .A1(G113), .A2(n998), .ZN(n534) );
  AND2_X1 U576 ( .A1(n535), .A2(n534), .ZN(n536) );
  AND2_X1 U577 ( .A1(n537), .A2(n536), .ZN(n538) );
  NOR2_X1 U578 ( .A1(G651), .A2(G543), .ZN(n638) );
  NAND2_X1 U579 ( .A1(G85), .A2(n638), .ZN(n540) );
  XOR2_X1 U580 ( .A(KEYINPUT0), .B(G543), .Z(n652) );
  INV_X1 U581 ( .A(G651), .ZN(n541) );
  NOR2_X1 U582 ( .A1(n652), .A2(n541), .ZN(n641) );
  NAND2_X1 U583 ( .A1(G72), .A2(n641), .ZN(n539) );
  NAND2_X1 U584 ( .A1(n540), .A2(n539), .ZN(n546) );
  NOR2_X1 U585 ( .A1(G543), .A2(n541), .ZN(n542) );
  XOR2_X1 U586 ( .A(KEYINPUT1), .B(n542), .Z(n651) );
  NAND2_X1 U587 ( .A1(G60), .A2(n651), .ZN(n544) );
  NAND2_X1 U588 ( .A1(G47), .A2(n647), .ZN(n543) );
  NAND2_X1 U589 ( .A1(n544), .A2(n543), .ZN(n545) );
  OR2_X1 U590 ( .A1(n546), .A2(n545), .ZN(G290) );
  NAND2_X1 U591 ( .A1(G64), .A2(n651), .ZN(n547) );
  XOR2_X1 U592 ( .A(KEYINPUT72), .B(n547), .Z(n554) );
  NAND2_X1 U593 ( .A1(G90), .A2(n638), .ZN(n549) );
  NAND2_X1 U594 ( .A1(G77), .A2(n641), .ZN(n548) );
  NAND2_X1 U595 ( .A1(n549), .A2(n548), .ZN(n550) );
  XNOR2_X1 U596 ( .A(n550), .B(KEYINPUT9), .ZN(n552) );
  NAND2_X1 U597 ( .A1(G52), .A2(n647), .ZN(n551) );
  NAND2_X1 U598 ( .A1(n552), .A2(n551), .ZN(n553) );
  NOR2_X1 U599 ( .A1(n554), .A2(n553), .ZN(G171) );
  AND2_X1 U600 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U601 ( .A(G132), .ZN(G219) );
  INV_X1 U602 ( .A(G82), .ZN(G220) );
  INV_X1 U603 ( .A(G57), .ZN(G237) );
  INV_X1 U604 ( .A(G120), .ZN(G236) );
  INV_X1 U605 ( .A(G171), .ZN(G301) );
  NAND2_X1 U606 ( .A1(n638), .A2(G89), .ZN(n555) );
  XNOR2_X1 U607 ( .A(n555), .B(KEYINPUT4), .ZN(n557) );
  NAND2_X1 U608 ( .A1(G76), .A2(n641), .ZN(n556) );
  NAND2_X1 U609 ( .A1(n557), .A2(n556), .ZN(n558) );
  XNOR2_X1 U610 ( .A(KEYINPUT5), .B(n558), .ZN(n564) );
  NAND2_X1 U611 ( .A1(n651), .A2(G63), .ZN(n559) );
  XOR2_X1 U612 ( .A(KEYINPUT79), .B(n559), .Z(n561) );
  NAND2_X1 U613 ( .A1(n647), .A2(G51), .ZN(n560) );
  NAND2_X1 U614 ( .A1(n561), .A2(n560), .ZN(n562) );
  XOR2_X1 U615 ( .A(KEYINPUT6), .B(n562), .Z(n563) );
  NAND2_X1 U616 ( .A1(n564), .A2(n563), .ZN(n565) );
  XNOR2_X1 U617 ( .A(KEYINPUT7), .B(n565), .ZN(G168) );
  XOR2_X1 U618 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  XOR2_X1 U619 ( .A(KEYINPUT74), .B(KEYINPUT11), .Z(n568) );
  NAND2_X1 U620 ( .A1(G7), .A2(G661), .ZN(n566) );
  XOR2_X1 U621 ( .A(n566), .B(KEYINPUT10), .Z(n837) );
  NAND2_X1 U622 ( .A1(G567), .A2(n837), .ZN(n567) );
  XNOR2_X1 U623 ( .A(n568), .B(n567), .ZN(G234) );
  NAND2_X1 U624 ( .A1(G81), .A2(n638), .ZN(n569) );
  XNOR2_X1 U625 ( .A(n569), .B(KEYINPUT12), .ZN(n570) );
  XNOR2_X1 U626 ( .A(n570), .B(KEYINPUT76), .ZN(n572) );
  NAND2_X1 U627 ( .A1(G68), .A2(n641), .ZN(n571) );
  NAND2_X1 U628 ( .A1(n572), .A2(n571), .ZN(n573) );
  XOR2_X1 U629 ( .A(KEYINPUT13), .B(n573), .Z(n577) );
  NAND2_X1 U630 ( .A1(G56), .A2(n651), .ZN(n574) );
  XNOR2_X1 U631 ( .A(n574), .B(KEYINPUT14), .ZN(n575) );
  XNOR2_X1 U632 ( .A(n575), .B(KEYINPUT75), .ZN(n576) );
  NOR2_X1 U633 ( .A1(n577), .A2(n576), .ZN(n579) );
  NAND2_X1 U634 ( .A1(n647), .A2(G43), .ZN(n578) );
  NAND2_X1 U635 ( .A1(n579), .A2(n578), .ZN(n1027) );
  INV_X1 U636 ( .A(G860), .ZN(n618) );
  OR2_X1 U637 ( .A1(n1027), .A2(n618), .ZN(G153) );
  NAND2_X1 U638 ( .A1(G79), .A2(n641), .ZN(n581) );
  NAND2_X1 U639 ( .A1(G54), .A2(n647), .ZN(n580) );
  NAND2_X1 U640 ( .A1(n581), .A2(n580), .ZN(n586) );
  NAND2_X1 U641 ( .A1(G92), .A2(n638), .ZN(n583) );
  NAND2_X1 U642 ( .A1(G66), .A2(n651), .ZN(n582) );
  NAND2_X1 U643 ( .A1(n583), .A2(n582), .ZN(n584) );
  XOR2_X1 U644 ( .A(KEYINPUT77), .B(n584), .Z(n585) );
  NOR2_X1 U645 ( .A1(n586), .A2(n585), .ZN(n587) );
  XNOR2_X1 U646 ( .A(KEYINPUT15), .B(n587), .ZN(n712) );
  INV_X1 U647 ( .A(G868), .ZN(n664) );
  NAND2_X1 U648 ( .A1(n712), .A2(n664), .ZN(n588) );
  XNOR2_X1 U649 ( .A(n588), .B(KEYINPUT78), .ZN(n590) );
  NAND2_X1 U650 ( .A1(G868), .A2(G301), .ZN(n589) );
  NAND2_X1 U651 ( .A1(n590), .A2(n589), .ZN(G284) );
  NAND2_X1 U652 ( .A1(G65), .A2(n651), .ZN(n592) );
  NAND2_X1 U653 ( .A1(G53), .A2(n647), .ZN(n591) );
  NAND2_X1 U654 ( .A1(n592), .A2(n591), .ZN(n593) );
  XNOR2_X1 U655 ( .A(KEYINPUT73), .B(n593), .ZN(n597) );
  NAND2_X1 U656 ( .A1(G91), .A2(n638), .ZN(n595) );
  NAND2_X1 U657 ( .A1(G78), .A2(n641), .ZN(n594) );
  AND2_X1 U658 ( .A1(n595), .A2(n594), .ZN(n596) );
  NAND2_X1 U659 ( .A1(n597), .A2(n596), .ZN(G299) );
  NOR2_X1 U660 ( .A1(G868), .A2(G299), .ZN(n598) );
  XNOR2_X1 U661 ( .A(n598), .B(KEYINPUT80), .ZN(n600) );
  NOR2_X1 U662 ( .A1(n664), .A2(G286), .ZN(n599) );
  NOR2_X1 U663 ( .A1(n600), .A2(n599), .ZN(n601) );
  XOR2_X1 U664 ( .A(KEYINPUT81), .B(n601), .Z(G297) );
  NAND2_X1 U665 ( .A1(n618), .A2(G559), .ZN(n602) );
  INV_X1 U666 ( .A(n712), .ZN(n1028) );
  NAND2_X1 U667 ( .A1(n602), .A2(n1028), .ZN(n603) );
  XNOR2_X1 U668 ( .A(n603), .B(KEYINPUT16), .ZN(G148) );
  NAND2_X1 U669 ( .A1(n1028), .A2(G868), .ZN(n604) );
  NOR2_X1 U670 ( .A1(G559), .A2(n604), .ZN(n605) );
  XNOR2_X1 U671 ( .A(n605), .B(KEYINPUT82), .ZN(n607) );
  NOR2_X1 U672 ( .A1(n1027), .A2(G868), .ZN(n606) );
  NOR2_X1 U673 ( .A1(n607), .A2(n606), .ZN(G282) );
  NAND2_X1 U674 ( .A1(G123), .A2(n997), .ZN(n608) );
  XOR2_X1 U675 ( .A(KEYINPUT83), .B(n608), .Z(n609) );
  XNOR2_X1 U676 ( .A(n609), .B(KEYINPUT18), .ZN(n611) );
  NAND2_X1 U677 ( .A1(G111), .A2(n998), .ZN(n610) );
  NAND2_X1 U678 ( .A1(n611), .A2(n610), .ZN(n615) );
  NAND2_X1 U679 ( .A1(G99), .A2(n1003), .ZN(n613) );
  NAND2_X1 U680 ( .A1(G135), .A2(n1001), .ZN(n612) );
  NAND2_X1 U681 ( .A1(n613), .A2(n612), .ZN(n614) );
  NOR2_X1 U682 ( .A1(n615), .A2(n614), .ZN(n1017) );
  XNOR2_X1 U683 ( .A(n1017), .B(G2096), .ZN(n616) );
  INV_X1 U684 ( .A(G2100), .ZN(n978) );
  NAND2_X1 U685 ( .A1(n616), .A2(n978), .ZN(G156) );
  NAND2_X1 U686 ( .A1(G559), .A2(n1028), .ZN(n617) );
  XOR2_X1 U687 ( .A(n1027), .B(n617), .Z(n661) );
  NAND2_X1 U688 ( .A1(n618), .A2(n661), .ZN(n627) );
  NAND2_X1 U689 ( .A1(G93), .A2(n638), .ZN(n620) );
  NAND2_X1 U690 ( .A1(G80), .A2(n641), .ZN(n619) );
  NAND2_X1 U691 ( .A1(n620), .A2(n619), .ZN(n626) );
  NAND2_X1 U692 ( .A1(n647), .A2(G55), .ZN(n621) );
  XNOR2_X1 U693 ( .A(n621), .B(KEYINPUT84), .ZN(n623) );
  NAND2_X1 U694 ( .A1(G67), .A2(n651), .ZN(n622) );
  NAND2_X1 U695 ( .A1(n623), .A2(n622), .ZN(n624) );
  XOR2_X1 U696 ( .A(KEYINPUT85), .B(n624), .Z(n625) );
  NOR2_X1 U697 ( .A1(n626), .A2(n625), .ZN(n663) );
  XOR2_X1 U698 ( .A(n627), .B(n663), .Z(G145) );
  NAND2_X1 U699 ( .A1(G86), .A2(n638), .ZN(n629) );
  NAND2_X1 U700 ( .A1(G61), .A2(n651), .ZN(n628) );
  NAND2_X1 U701 ( .A1(n629), .A2(n628), .ZN(n630) );
  XNOR2_X1 U702 ( .A(KEYINPUT86), .B(n630), .ZN(n634) );
  NAND2_X1 U703 ( .A1(G73), .A2(n641), .ZN(n631) );
  XNOR2_X1 U704 ( .A(n631), .B(KEYINPUT2), .ZN(n632) );
  XNOR2_X1 U705 ( .A(n632), .B(KEYINPUT87), .ZN(n633) );
  NOR2_X1 U706 ( .A1(n634), .A2(n633), .ZN(n635) );
  XNOR2_X1 U707 ( .A(n635), .B(KEYINPUT88), .ZN(n637) );
  NAND2_X1 U708 ( .A1(G48), .A2(n647), .ZN(n636) );
  NAND2_X1 U709 ( .A1(n637), .A2(n636), .ZN(G305) );
  NAND2_X1 U710 ( .A1(G88), .A2(n638), .ZN(n640) );
  NAND2_X1 U711 ( .A1(G62), .A2(n651), .ZN(n639) );
  NAND2_X1 U712 ( .A1(n640), .A2(n639), .ZN(n644) );
  NAND2_X1 U713 ( .A1(G75), .A2(n641), .ZN(n642) );
  XNOR2_X1 U714 ( .A(KEYINPUT89), .B(n642), .ZN(n643) );
  NOR2_X1 U715 ( .A1(n644), .A2(n643), .ZN(n646) );
  NAND2_X1 U716 ( .A1(n647), .A2(G50), .ZN(n645) );
  NAND2_X1 U717 ( .A1(n646), .A2(n645), .ZN(G303) );
  NAND2_X1 U718 ( .A1(G49), .A2(n647), .ZN(n649) );
  NAND2_X1 U719 ( .A1(G74), .A2(G651), .ZN(n648) );
  NAND2_X1 U720 ( .A1(n649), .A2(n648), .ZN(n650) );
  NOR2_X1 U721 ( .A1(n651), .A2(n650), .ZN(n654) );
  NAND2_X1 U722 ( .A1(n652), .A2(G87), .ZN(n653) );
  NAND2_X1 U723 ( .A1(n654), .A2(n653), .ZN(G288) );
  XOR2_X1 U724 ( .A(KEYINPUT19), .B(KEYINPUT90), .Z(n655) );
  XNOR2_X1 U725 ( .A(G288), .B(n655), .ZN(n656) );
  XOR2_X1 U726 ( .A(G303), .B(n656), .Z(n658) );
  XOR2_X1 U727 ( .A(G290), .B(G299), .Z(n657) );
  XNOR2_X1 U728 ( .A(n658), .B(n657), .ZN(n659) );
  XOR2_X1 U729 ( .A(n663), .B(n659), .Z(n660) );
  XNOR2_X1 U730 ( .A(G305), .B(n660), .ZN(n1026) );
  XOR2_X1 U731 ( .A(n1026), .B(n661), .Z(n662) );
  NOR2_X1 U732 ( .A1(n664), .A2(n662), .ZN(n666) );
  AND2_X1 U733 ( .A1(n664), .A2(n663), .ZN(n665) );
  NOR2_X1 U734 ( .A1(n666), .A2(n665), .ZN(G295) );
  NAND2_X1 U735 ( .A1(G2078), .A2(G2084), .ZN(n667) );
  XOR2_X1 U736 ( .A(KEYINPUT20), .B(n667), .Z(n668) );
  NAND2_X1 U737 ( .A1(G2090), .A2(n668), .ZN(n669) );
  XNOR2_X1 U738 ( .A(KEYINPUT21), .B(n669), .ZN(n670) );
  NAND2_X1 U739 ( .A1(n670), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U740 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U741 ( .A1(G236), .A2(G237), .ZN(n671) );
  NAND2_X1 U742 ( .A1(G69), .A2(n671), .ZN(n672) );
  XNOR2_X1 U743 ( .A(KEYINPUT91), .B(n672), .ZN(n673) );
  NAND2_X1 U744 ( .A1(n673), .A2(G108), .ZN(n965) );
  NAND2_X1 U745 ( .A1(n965), .A2(G567), .ZN(n678) );
  NOR2_X1 U746 ( .A1(G220), .A2(G219), .ZN(n674) );
  XOR2_X1 U747 ( .A(KEYINPUT22), .B(n674), .Z(n675) );
  NOR2_X1 U748 ( .A1(G218), .A2(n675), .ZN(n676) );
  NAND2_X1 U749 ( .A1(G96), .A2(n676), .ZN(n964) );
  NAND2_X1 U750 ( .A1(n964), .A2(G2106), .ZN(n677) );
  NAND2_X1 U751 ( .A1(n678), .A2(n677), .ZN(n1038) );
  NAND2_X1 U752 ( .A1(G483), .A2(G661), .ZN(n679) );
  NOR2_X1 U753 ( .A1(n1038), .A2(n679), .ZN(n841) );
  NAND2_X1 U754 ( .A1(n841), .A2(G36), .ZN(G176) );
  NAND2_X1 U755 ( .A1(G138), .A2(n1001), .ZN(n680) );
  XNOR2_X1 U756 ( .A(n680), .B(KEYINPUT92), .ZN(n682) );
  NAND2_X1 U757 ( .A1(n997), .A2(G126), .ZN(n681) );
  NAND2_X1 U758 ( .A1(n682), .A2(n681), .ZN(n686) );
  NAND2_X1 U759 ( .A1(G114), .A2(n998), .ZN(n684) );
  NAND2_X1 U760 ( .A1(G102), .A2(n1003), .ZN(n683) );
  NAND2_X1 U761 ( .A1(n684), .A2(n683), .ZN(n685) );
  NOR2_X1 U762 ( .A1(n686), .A2(n685), .ZN(G164) );
  INV_X1 U763 ( .A(G303), .ZN(G166) );
  NAND2_X1 U764 ( .A1(G40), .A2(G160), .ZN(n783) );
  NOR2_X1 U765 ( .A1(G1384), .A2(G164), .ZN(n687) );
  XOR2_X1 U766 ( .A(n687), .B(KEYINPUT64), .Z(n781) );
  NOR2_X4 U767 ( .A1(n783), .A2(n781), .ZN(n715) );
  INV_X1 U768 ( .A(n715), .ZN(n716) );
  NAND2_X1 U769 ( .A1(G8), .A2(n716), .ZN(n697) );
  NOR2_X1 U770 ( .A1(G1966), .A2(n697), .ZN(n747) );
  NOR2_X1 U771 ( .A1(G2084), .A2(n716), .ZN(n743) );
  NOR2_X1 U772 ( .A1(n747), .A2(n743), .ZN(n688) );
  NAND2_X1 U773 ( .A1(G8), .A2(n688), .ZN(n689) );
  XNOR2_X1 U774 ( .A(KEYINPUT30), .B(n689), .ZN(n690) );
  NOR2_X1 U775 ( .A1(n690), .A2(G168), .ZN(n695) );
  XNOR2_X1 U776 ( .A(G2078), .B(KEYINPUT25), .ZN(n935) );
  NAND2_X1 U777 ( .A1(n715), .A2(n935), .ZN(n691) );
  XOR2_X1 U778 ( .A(KEYINPUT99), .B(n691), .Z(n693) );
  OR2_X1 U779 ( .A1(n715), .A2(G1961), .ZN(n692) );
  NAND2_X1 U780 ( .A1(n693), .A2(n692), .ZN(n734) );
  NOR2_X1 U781 ( .A1(G171), .A2(n734), .ZN(n694) );
  NOR2_X1 U782 ( .A1(n695), .A2(n694), .ZN(n696) );
  XOR2_X1 U783 ( .A(KEYINPUT31), .B(n696), .Z(n744) );
  INV_X1 U784 ( .A(G8), .ZN(n704) );
  BUF_X1 U785 ( .A(n697), .Z(n762) );
  NOR2_X1 U786 ( .A1(G1971), .A2(n762), .ZN(n698) );
  XNOR2_X1 U787 ( .A(KEYINPUT103), .B(n698), .ZN(n702) );
  NOR2_X1 U788 ( .A1(n716), .A2(G2090), .ZN(n699) );
  XNOR2_X1 U789 ( .A(KEYINPUT104), .B(n699), .ZN(n700) );
  NOR2_X1 U790 ( .A1(G166), .A2(n700), .ZN(n701) );
  NAND2_X1 U791 ( .A1(n702), .A2(n701), .ZN(n703) );
  OR2_X1 U792 ( .A1(n704), .A2(n703), .ZN(n738) );
  AND2_X1 U793 ( .A1(n744), .A2(n738), .ZN(n737) );
  INV_X1 U794 ( .A(G299), .ZN(n885) );
  NAND2_X1 U795 ( .A1(n715), .A2(G2072), .ZN(n706) );
  XNOR2_X1 U796 ( .A(KEYINPUT27), .B(KEYINPUT100), .ZN(n705) );
  XNOR2_X1 U797 ( .A(n706), .B(n705), .ZN(n708) );
  XNOR2_X1 U798 ( .A(G1956), .B(KEYINPUT101), .ZN(n916) );
  NOR2_X1 U799 ( .A1(n715), .A2(n916), .ZN(n707) );
  NOR2_X1 U800 ( .A1(n708), .A2(n707), .ZN(n728) );
  NOR2_X1 U801 ( .A1(n885), .A2(n728), .ZN(n709) );
  XOR2_X1 U802 ( .A(n709), .B(KEYINPUT28), .Z(n732) );
  AND2_X1 U803 ( .A1(n715), .A2(G1996), .ZN(n711) );
  XNOR2_X1 U804 ( .A(KEYINPUT65), .B(KEYINPUT26), .ZN(n710) );
  XNOR2_X1 U805 ( .A(n711), .B(n710), .ZN(n723) );
  NAND2_X1 U806 ( .A1(n716), .A2(G1341), .ZN(n722) );
  NOR2_X1 U807 ( .A1(n712), .A2(n1027), .ZN(n713) );
  AND2_X1 U808 ( .A1(n722), .A2(n713), .ZN(n714) );
  NAND2_X1 U809 ( .A1(n723), .A2(n714), .ZN(n720) );
  NOR2_X1 U810 ( .A1(n715), .A2(G1348), .ZN(n718) );
  NOR2_X1 U811 ( .A1(n716), .A2(G2067), .ZN(n717) );
  NOR2_X1 U812 ( .A1(n718), .A2(n717), .ZN(n719) );
  NAND2_X1 U813 ( .A1(n720), .A2(n719), .ZN(n721) );
  XNOR2_X1 U814 ( .A(n721), .B(KEYINPUT102), .ZN(n727) );
  NAND2_X1 U815 ( .A1(n723), .A2(n722), .ZN(n724) );
  NOR2_X1 U816 ( .A1(n1027), .A2(n724), .ZN(n725) );
  OR2_X1 U817 ( .A1(n725), .A2(n1028), .ZN(n726) );
  NAND2_X1 U818 ( .A1(n727), .A2(n726), .ZN(n730) );
  NAND2_X1 U819 ( .A1(n885), .A2(n728), .ZN(n729) );
  NAND2_X1 U820 ( .A1(n730), .A2(n729), .ZN(n731) );
  NAND2_X1 U821 ( .A1(n732), .A2(n731), .ZN(n733) );
  XOR2_X1 U822 ( .A(KEYINPUT29), .B(n733), .Z(n736) );
  NAND2_X1 U823 ( .A1(G171), .A2(n734), .ZN(n735) );
  NAND2_X1 U824 ( .A1(n736), .A2(n735), .ZN(n745) );
  NAND2_X1 U825 ( .A1(n737), .A2(n745), .ZN(n741) );
  INV_X1 U826 ( .A(n738), .ZN(n739) );
  OR2_X1 U827 ( .A1(n739), .A2(G286), .ZN(n740) );
  NAND2_X1 U828 ( .A1(n741), .A2(n740), .ZN(n742) );
  XNOR2_X1 U829 ( .A(n742), .B(KEYINPUT32), .ZN(n760) );
  NAND2_X1 U830 ( .A1(G8), .A2(n743), .ZN(n749) );
  AND2_X1 U831 ( .A1(n745), .A2(n744), .ZN(n746) );
  NOR2_X1 U832 ( .A1(n747), .A2(n746), .ZN(n748) );
  NAND2_X1 U833 ( .A1(n749), .A2(n748), .ZN(n766) );
  NAND2_X1 U834 ( .A1(n760), .A2(n766), .ZN(n756) );
  NOR2_X1 U835 ( .A1(G2090), .A2(G303), .ZN(n750) );
  NAND2_X1 U836 ( .A1(G8), .A2(n750), .ZN(n754) );
  NOR2_X1 U837 ( .A1(G1981), .A2(G305), .ZN(n751) );
  XOR2_X1 U838 ( .A(n751), .B(KEYINPUT24), .Z(n752) );
  NOR2_X1 U839 ( .A1(n762), .A2(n752), .ZN(n757) );
  INV_X1 U840 ( .A(n757), .ZN(n753) );
  AND2_X1 U841 ( .A1(n754), .A2(n753), .ZN(n755) );
  AND2_X1 U842 ( .A1(n756), .A2(n755), .ZN(n759) );
  NOR2_X1 U843 ( .A1(n757), .A2(n762), .ZN(n758) );
  NOR2_X1 U844 ( .A1(n759), .A2(n758), .ZN(n780) );
  XOR2_X1 U845 ( .A(G1981), .B(G305), .Z(n881) );
  AND2_X1 U846 ( .A1(n760), .A2(n881), .ZN(n768) );
  NAND2_X1 U847 ( .A1(G1976), .A2(G288), .ZN(n889) );
  INV_X1 U848 ( .A(n889), .ZN(n761) );
  NOR2_X1 U849 ( .A1(KEYINPUT33), .A2(n524), .ZN(n765) );
  NOR2_X1 U850 ( .A1(G1976), .A2(G288), .ZN(n771) );
  NAND2_X1 U851 ( .A1(n771), .A2(KEYINPUT33), .ZN(n763) );
  NOR2_X1 U852 ( .A1(n763), .A2(n762), .ZN(n764) );
  NOR2_X1 U853 ( .A1(n765), .A2(n764), .ZN(n769) );
  AND2_X1 U854 ( .A1(n766), .A2(n769), .ZN(n767) );
  NAND2_X1 U855 ( .A1(n768), .A2(n767), .ZN(n778) );
  INV_X1 U856 ( .A(n881), .ZN(n776) );
  INV_X1 U857 ( .A(n769), .ZN(n774) );
  NOR2_X1 U858 ( .A1(G1971), .A2(G303), .ZN(n770) );
  NOR2_X1 U859 ( .A1(n771), .A2(n770), .ZN(n893) );
  INV_X1 U860 ( .A(KEYINPUT33), .ZN(n772) );
  AND2_X1 U861 ( .A1(n893), .A2(n772), .ZN(n773) );
  OR2_X1 U862 ( .A1(n774), .A2(n773), .ZN(n775) );
  OR2_X1 U863 ( .A1(n776), .A2(n775), .ZN(n777) );
  NAND2_X1 U864 ( .A1(n778), .A2(n777), .ZN(n779) );
  OR2_X1 U865 ( .A1(n780), .A2(n779), .ZN(n818) );
  XNOR2_X1 U866 ( .A(G1986), .B(G290), .ZN(n895) );
  INV_X1 U867 ( .A(n781), .ZN(n782) );
  NOR2_X1 U868 ( .A1(n783), .A2(n782), .ZN(n784) );
  XNOR2_X1 U869 ( .A(KEYINPUT93), .B(n784), .ZN(n815) );
  INV_X1 U870 ( .A(n815), .ZN(n828) );
  NAND2_X1 U871 ( .A1(n895), .A2(n828), .ZN(n795) );
  NAND2_X1 U872 ( .A1(n1003), .A2(G104), .ZN(n785) );
  XNOR2_X1 U873 ( .A(n785), .B(KEYINPUT94), .ZN(n787) );
  NAND2_X1 U874 ( .A1(G140), .A2(n1001), .ZN(n786) );
  NAND2_X1 U875 ( .A1(n787), .A2(n786), .ZN(n788) );
  XNOR2_X1 U876 ( .A(KEYINPUT34), .B(n788), .ZN(n793) );
  NAND2_X1 U877 ( .A1(G128), .A2(n997), .ZN(n790) );
  NAND2_X1 U878 ( .A1(G116), .A2(n998), .ZN(n789) );
  NAND2_X1 U879 ( .A1(n790), .A2(n789), .ZN(n791) );
  XOR2_X1 U880 ( .A(KEYINPUT35), .B(n791), .Z(n792) );
  NOR2_X1 U881 ( .A1(n793), .A2(n792), .ZN(n794) );
  XOR2_X1 U882 ( .A(KEYINPUT36), .B(n794), .Z(n1022) );
  XOR2_X1 U883 ( .A(G2067), .B(KEYINPUT37), .Z(n827) );
  AND2_X1 U884 ( .A1(n1022), .A2(n827), .ZN(n852) );
  NAND2_X1 U885 ( .A1(n852), .A2(n828), .ZN(n819) );
  NAND2_X1 U886 ( .A1(n795), .A2(n819), .ZN(n816) );
  NAND2_X1 U887 ( .A1(G105), .A2(n1003), .ZN(n796) );
  XNOR2_X1 U888 ( .A(n796), .B(KEYINPUT38), .ZN(n803) );
  NAND2_X1 U889 ( .A1(G129), .A2(n997), .ZN(n798) );
  NAND2_X1 U890 ( .A1(G141), .A2(n1001), .ZN(n797) );
  NAND2_X1 U891 ( .A1(n798), .A2(n797), .ZN(n801) );
  NAND2_X1 U892 ( .A1(G117), .A2(n998), .ZN(n799) );
  XNOR2_X1 U893 ( .A(KEYINPUT97), .B(n799), .ZN(n800) );
  NOR2_X1 U894 ( .A1(n801), .A2(n800), .ZN(n802) );
  NAND2_X1 U895 ( .A1(n803), .A2(n802), .ZN(n1012) );
  NAND2_X1 U896 ( .A1(G1996), .A2(n1012), .ZN(n813) );
  NAND2_X1 U897 ( .A1(n1003), .A2(G95), .ZN(n804) );
  XOR2_X1 U898 ( .A(KEYINPUT95), .B(n804), .Z(n806) );
  NAND2_X1 U899 ( .A1(n1001), .A2(G131), .ZN(n805) );
  NAND2_X1 U900 ( .A1(n806), .A2(n805), .ZN(n807) );
  XOR2_X1 U901 ( .A(KEYINPUT96), .B(n807), .Z(n811) );
  NAND2_X1 U902 ( .A1(G119), .A2(n997), .ZN(n809) );
  NAND2_X1 U903 ( .A1(G107), .A2(n998), .ZN(n808) );
  AND2_X1 U904 ( .A1(n809), .A2(n808), .ZN(n810) );
  NAND2_X1 U905 ( .A1(n811), .A2(n810), .ZN(n1019) );
  NAND2_X1 U906 ( .A1(G1991), .A2(n1019), .ZN(n812) );
  NAND2_X1 U907 ( .A1(n813), .A2(n812), .ZN(n814) );
  XOR2_X1 U908 ( .A(KEYINPUT98), .B(n814), .Z(n874) );
  NOR2_X1 U909 ( .A1(n815), .A2(n874), .ZN(n822) );
  NOR2_X1 U910 ( .A1(n816), .A2(n822), .ZN(n817) );
  NAND2_X1 U911 ( .A1(n818), .A2(n817), .ZN(n834) );
  INV_X1 U912 ( .A(n819), .ZN(n832) );
  NOR2_X1 U913 ( .A1(G1996), .A2(n1012), .ZN(n854) );
  NOR2_X1 U914 ( .A1(G1986), .A2(G290), .ZN(n820) );
  NOR2_X1 U915 ( .A1(G1991), .A2(n1019), .ZN(n868) );
  NOR2_X1 U916 ( .A1(n820), .A2(n868), .ZN(n821) );
  NOR2_X1 U917 ( .A1(n822), .A2(n821), .ZN(n823) );
  XOR2_X1 U918 ( .A(KEYINPUT105), .B(n823), .Z(n824) );
  NOR2_X1 U919 ( .A1(n854), .A2(n824), .ZN(n825) );
  XNOR2_X1 U920 ( .A(KEYINPUT39), .B(n825), .ZN(n826) );
  NAND2_X1 U921 ( .A1(n826), .A2(n828), .ZN(n830) );
  NOR2_X1 U922 ( .A1(n1022), .A2(n827), .ZN(n851) );
  NAND2_X1 U923 ( .A1(n851), .A2(n828), .ZN(n829) );
  AND2_X1 U924 ( .A1(n830), .A2(n829), .ZN(n831) );
  OR2_X1 U925 ( .A1(n832), .A2(n831), .ZN(n833) );
  NAND2_X1 U926 ( .A1(n834), .A2(n833), .ZN(n836) );
  XNOR2_X1 U927 ( .A(KEYINPUT106), .B(KEYINPUT40), .ZN(n835) );
  XNOR2_X1 U928 ( .A(n836), .B(n835), .ZN(G329) );
  NAND2_X1 U929 ( .A1(G2106), .A2(n837), .ZN(G217) );
  INV_X1 U930 ( .A(n837), .ZN(G223) );
  AND2_X1 U931 ( .A1(G15), .A2(G2), .ZN(n838) );
  NAND2_X1 U932 ( .A1(G661), .A2(n838), .ZN(G259) );
  NAND2_X1 U933 ( .A1(G3), .A2(G1), .ZN(n839) );
  XOR2_X1 U934 ( .A(KEYINPUT109), .B(n839), .Z(n840) );
  NAND2_X1 U935 ( .A1(n841), .A2(n840), .ZN(n842) );
  XNOR2_X1 U936 ( .A(KEYINPUT110), .B(n842), .ZN(G188) );
  NAND2_X1 U938 ( .A1(G124), .A2(n997), .ZN(n843) );
  XNOR2_X1 U939 ( .A(n843), .B(KEYINPUT44), .ZN(n846) );
  NAND2_X1 U940 ( .A1(G112), .A2(n998), .ZN(n844) );
  XOR2_X1 U941 ( .A(KEYINPUT113), .B(n844), .Z(n845) );
  NAND2_X1 U942 ( .A1(n846), .A2(n845), .ZN(n850) );
  NAND2_X1 U943 ( .A1(G100), .A2(n1003), .ZN(n848) );
  NAND2_X1 U944 ( .A1(G136), .A2(n1001), .ZN(n847) );
  NAND2_X1 U945 ( .A1(n848), .A2(n847), .ZN(n849) );
  NOR2_X1 U946 ( .A1(n850), .A2(n849), .ZN(G162) );
  NOR2_X1 U947 ( .A1(n852), .A2(n851), .ZN(n873) );
  XOR2_X1 U948 ( .A(G2090), .B(G162), .Z(n853) );
  NOR2_X1 U949 ( .A1(n854), .A2(n853), .ZN(n855) );
  XOR2_X1 U950 ( .A(KEYINPUT51), .B(n855), .Z(n870) );
  NAND2_X1 U951 ( .A1(G103), .A2(n1003), .ZN(n857) );
  NAND2_X1 U952 ( .A1(G139), .A2(n1001), .ZN(n856) );
  NAND2_X1 U953 ( .A1(n857), .A2(n856), .ZN(n863) );
  NAND2_X1 U954 ( .A1(n998), .A2(G115), .ZN(n858) );
  XOR2_X1 U955 ( .A(KEYINPUT115), .B(n858), .Z(n860) );
  NAND2_X1 U956 ( .A1(n997), .A2(G127), .ZN(n859) );
  NAND2_X1 U957 ( .A1(n860), .A2(n859), .ZN(n861) );
  XOR2_X1 U958 ( .A(KEYINPUT47), .B(n861), .Z(n862) );
  NOR2_X1 U959 ( .A1(n863), .A2(n862), .ZN(n1010) );
  XOR2_X1 U960 ( .A(G2072), .B(n1010), .Z(n865) );
  XOR2_X1 U961 ( .A(G164), .B(G2078), .Z(n864) );
  NOR2_X1 U962 ( .A1(n865), .A2(n864), .ZN(n866) );
  XOR2_X1 U963 ( .A(KEYINPUT50), .B(n866), .Z(n867) );
  NOR2_X1 U964 ( .A1(n868), .A2(n867), .ZN(n869) );
  NAND2_X1 U965 ( .A1(n870), .A2(n869), .ZN(n871) );
  NOR2_X1 U966 ( .A1(n1017), .A2(n871), .ZN(n872) );
  NAND2_X1 U967 ( .A1(n873), .A2(n872), .ZN(n877) );
  XNOR2_X1 U968 ( .A(G2084), .B(G160), .ZN(n875) );
  NAND2_X1 U969 ( .A1(n875), .A2(n874), .ZN(n876) );
  NOR2_X1 U970 ( .A1(n877), .A2(n876), .ZN(n878) );
  XNOR2_X1 U971 ( .A(KEYINPUT52), .B(n878), .ZN(n879) );
  INV_X1 U972 ( .A(KEYINPUT55), .ZN(n954) );
  NAND2_X1 U973 ( .A1(n879), .A2(n954), .ZN(n880) );
  NAND2_X1 U974 ( .A1(n880), .A2(G29), .ZN(n962) );
  INV_X1 U975 ( .A(G16), .ZN(n932) );
  XOR2_X1 U976 ( .A(n932), .B(KEYINPUT56), .Z(n903) );
  XNOR2_X1 U977 ( .A(G1966), .B(G168), .ZN(n882) );
  NAND2_X1 U978 ( .A1(n882), .A2(n881), .ZN(n883) );
  XNOR2_X1 U979 ( .A(n883), .B(KEYINPUT57), .ZN(n901) );
  XOR2_X1 U980 ( .A(G301), .B(KEYINPUT120), .Z(n884) );
  XOR2_X1 U981 ( .A(n884), .B(G1961), .Z(n887) );
  XOR2_X1 U982 ( .A(G1956), .B(n885), .Z(n886) );
  NOR2_X1 U983 ( .A1(n887), .A2(n886), .ZN(n897) );
  NAND2_X1 U984 ( .A1(G1971), .A2(G303), .ZN(n888) );
  NAND2_X1 U985 ( .A1(n889), .A2(n888), .ZN(n891) );
  XNOR2_X1 U986 ( .A(G1341), .B(n1027), .ZN(n890) );
  NOR2_X1 U987 ( .A1(n891), .A2(n890), .ZN(n892) );
  NAND2_X1 U988 ( .A1(n893), .A2(n892), .ZN(n894) );
  NOR2_X1 U989 ( .A1(n895), .A2(n894), .ZN(n896) );
  NAND2_X1 U990 ( .A1(n897), .A2(n896), .ZN(n899) );
  XOR2_X1 U991 ( .A(G1348), .B(n1028), .Z(n898) );
  NOR2_X1 U992 ( .A1(n899), .A2(n898), .ZN(n900) );
  NAND2_X1 U993 ( .A1(n901), .A2(n900), .ZN(n902) );
  NAND2_X1 U994 ( .A1(n903), .A2(n902), .ZN(n934) );
  XOR2_X1 U995 ( .A(KEYINPUT126), .B(KEYINPUT61), .Z(n930) );
  XOR2_X1 U996 ( .A(G1966), .B(G21), .Z(n905) );
  XOR2_X1 U997 ( .A(G1961), .B(G5), .Z(n904) );
  NAND2_X1 U998 ( .A1(n905), .A2(n904), .ZN(n914) );
  XNOR2_X1 U999 ( .A(KEYINPUT124), .B(KEYINPUT125), .ZN(n906) );
  XNOR2_X1 U1000 ( .A(n906), .B(KEYINPUT58), .ZN(n912) );
  XOR2_X1 U1001 ( .A(G1986), .B(G24), .Z(n910) );
  XNOR2_X1 U1002 ( .A(G1971), .B(G22), .ZN(n908) );
  XNOR2_X1 U1003 ( .A(G23), .B(G1976), .ZN(n907) );
  NOR2_X1 U1004 ( .A1(n908), .A2(n907), .ZN(n909) );
  NAND2_X1 U1005 ( .A1(n910), .A2(n909), .ZN(n911) );
  XOR2_X1 U1006 ( .A(n912), .B(n911), .Z(n913) );
  NOR2_X1 U1007 ( .A1(n914), .A2(n913), .ZN(n928) );
  XNOR2_X1 U1008 ( .A(KEYINPUT122), .B(KEYINPUT123), .ZN(n915) );
  XNOR2_X1 U1009 ( .A(n915), .B(KEYINPUT60), .ZN(n926) );
  XOR2_X1 U1010 ( .A(n916), .B(G20), .Z(n918) );
  XNOR2_X1 U1011 ( .A(G6), .B(G1981), .ZN(n917) );
  NOR2_X1 U1012 ( .A1(n918), .A2(n917), .ZN(n924) );
  XOR2_X1 U1013 ( .A(G1348), .B(KEYINPUT59), .Z(n919) );
  XNOR2_X1 U1014 ( .A(G4), .B(n919), .ZN(n922) );
  XOR2_X1 U1015 ( .A(G1341), .B(KEYINPUT121), .Z(n920) );
  XNOR2_X1 U1016 ( .A(G19), .B(n920), .ZN(n921) );
  NOR2_X1 U1017 ( .A1(n922), .A2(n921), .ZN(n923) );
  NAND2_X1 U1018 ( .A1(n924), .A2(n923), .ZN(n925) );
  XNOR2_X1 U1019 ( .A(n926), .B(n925), .ZN(n927) );
  NAND2_X1 U1020 ( .A1(n928), .A2(n927), .ZN(n929) );
  XNOR2_X1 U1021 ( .A(n930), .B(n929), .ZN(n931) );
  NAND2_X1 U1022 ( .A1(n932), .A2(n931), .ZN(n933) );
  NAND2_X1 U1023 ( .A1(n934), .A2(n933), .ZN(n960) );
  XNOR2_X1 U1024 ( .A(G27), .B(n935), .ZN(n946) );
  XOR2_X1 U1025 ( .A(G1991), .B(G25), .Z(n936) );
  NAND2_X1 U1026 ( .A1(G28), .A2(n936), .ZN(n937) );
  XNOR2_X1 U1027 ( .A(n937), .B(KEYINPUT117), .ZN(n941) );
  XNOR2_X1 U1028 ( .A(G2067), .B(G26), .ZN(n939) );
  XNOR2_X1 U1029 ( .A(G1996), .B(G32), .ZN(n938) );
  NOR2_X1 U1030 ( .A1(n939), .A2(n938), .ZN(n940) );
  NAND2_X1 U1031 ( .A1(n941), .A2(n940), .ZN(n944) );
  XNOR2_X1 U1032 ( .A(KEYINPUT118), .B(G2072), .ZN(n942) );
  XNOR2_X1 U1033 ( .A(G33), .B(n942), .ZN(n943) );
  NOR2_X1 U1034 ( .A1(n944), .A2(n943), .ZN(n945) );
  NAND2_X1 U1035 ( .A1(n946), .A2(n945), .ZN(n947) );
  XNOR2_X1 U1036 ( .A(n947), .B(KEYINPUT53), .ZN(n950) );
  XOR2_X1 U1037 ( .A(G2084), .B(G34), .Z(n948) );
  XNOR2_X1 U1038 ( .A(KEYINPUT54), .B(n948), .ZN(n949) );
  NAND2_X1 U1039 ( .A1(n950), .A2(n949), .ZN(n952) );
  XNOR2_X1 U1040 ( .A(G35), .B(G2090), .ZN(n951) );
  NOR2_X1 U1041 ( .A1(n952), .A2(n951), .ZN(n953) );
  XOR2_X1 U1042 ( .A(n954), .B(n953), .Z(n956) );
  INV_X1 U1043 ( .A(G29), .ZN(n955) );
  NAND2_X1 U1044 ( .A1(n956), .A2(n955), .ZN(n957) );
  NAND2_X1 U1045 ( .A1(n957), .A2(G11), .ZN(n958) );
  XOR2_X1 U1046 ( .A(KEYINPUT119), .B(n958), .Z(n959) );
  NOR2_X1 U1047 ( .A1(n960), .A2(n959), .ZN(n961) );
  NAND2_X1 U1048 ( .A1(n962), .A2(n961), .ZN(n963) );
  XOR2_X1 U1049 ( .A(KEYINPUT62), .B(n963), .Z(G311) );
  XNOR2_X1 U1050 ( .A(KEYINPUT127), .B(G311), .ZN(G150) );
  INV_X1 U1051 ( .A(G108), .ZN(G238) );
  INV_X1 U1052 ( .A(G96), .ZN(G221) );
  NOR2_X1 U1053 ( .A1(n965), .A2(n964), .ZN(n966) );
  XOR2_X1 U1054 ( .A(n966), .B(KEYINPUT111), .Z(G325) );
  INV_X1 U1055 ( .A(G325), .ZN(G261) );
  XOR2_X1 U1056 ( .A(G2443), .B(G2430), .Z(n968) );
  XNOR2_X1 U1057 ( .A(G1341), .B(G2451), .ZN(n967) );
  XNOR2_X1 U1058 ( .A(n968), .B(n967), .ZN(n975) );
  XOR2_X1 U1059 ( .A(G2438), .B(G2435), .Z(n970) );
  XNOR2_X1 U1060 ( .A(G1348), .B(KEYINPUT107), .ZN(n969) );
  XNOR2_X1 U1061 ( .A(n970), .B(n969), .ZN(n971) );
  XOR2_X1 U1062 ( .A(n971), .B(G2454), .Z(n973) );
  XNOR2_X1 U1063 ( .A(G2446), .B(G2427), .ZN(n972) );
  XNOR2_X1 U1064 ( .A(n973), .B(n972), .ZN(n974) );
  XNOR2_X1 U1065 ( .A(n975), .B(n974), .ZN(n976) );
  NAND2_X1 U1066 ( .A1(n976), .A2(G14), .ZN(n977) );
  XOR2_X1 U1067 ( .A(KEYINPUT108), .B(n977), .Z(G401) );
  XNOR2_X1 U1068 ( .A(n978), .B(G2096), .ZN(n980) );
  XNOR2_X1 U1069 ( .A(G2072), .B(G2090), .ZN(n979) );
  XNOR2_X1 U1070 ( .A(n980), .B(n979), .ZN(n984) );
  XOR2_X1 U1071 ( .A(G2678), .B(KEYINPUT42), .Z(n982) );
  XNOR2_X1 U1072 ( .A(G2067), .B(KEYINPUT43), .ZN(n981) );
  XNOR2_X1 U1073 ( .A(n982), .B(n981), .ZN(n983) );
  XOR2_X1 U1074 ( .A(n984), .B(n983), .Z(n986) );
  XNOR2_X1 U1075 ( .A(G2078), .B(G2084), .ZN(n985) );
  XNOR2_X1 U1076 ( .A(n986), .B(n985), .ZN(G227) );
  XNOR2_X1 U1077 ( .A(G1986), .B(G1976), .ZN(n996) );
  XOR2_X1 U1078 ( .A(G1981), .B(G1971), .Z(n988) );
  XNOR2_X1 U1079 ( .A(G1996), .B(G1961), .ZN(n987) );
  XNOR2_X1 U1080 ( .A(n988), .B(n987), .ZN(n992) );
  XOR2_X1 U1081 ( .A(KEYINPUT112), .B(G2474), .Z(n990) );
  XNOR2_X1 U1082 ( .A(G1991), .B(G1966), .ZN(n989) );
  XNOR2_X1 U1083 ( .A(n990), .B(n989), .ZN(n991) );
  XOR2_X1 U1084 ( .A(n992), .B(n991), .Z(n994) );
  XNOR2_X1 U1085 ( .A(G1956), .B(KEYINPUT41), .ZN(n993) );
  XNOR2_X1 U1086 ( .A(n994), .B(n993), .ZN(n995) );
  XNOR2_X1 U1087 ( .A(n996), .B(n995), .ZN(G229) );
  NAND2_X1 U1088 ( .A1(G130), .A2(n997), .ZN(n1000) );
  NAND2_X1 U1089 ( .A1(G118), .A2(n998), .ZN(n999) );
  NAND2_X1 U1090 ( .A1(n1000), .A2(n999), .ZN(n1008) );
  NAND2_X1 U1091 ( .A1(n1001), .A2(G142), .ZN(n1002) );
  XNOR2_X1 U1092 ( .A(n1002), .B(KEYINPUT114), .ZN(n1005) );
  NAND2_X1 U1093 ( .A1(G106), .A2(n1003), .ZN(n1004) );
  NAND2_X1 U1094 ( .A1(n1005), .A2(n1004), .ZN(n1006) );
  XOR2_X1 U1095 ( .A(KEYINPUT45), .B(n1006), .Z(n1007) );
  NOR2_X1 U1096 ( .A1(n1008), .A2(n1007), .ZN(n1009) );
  XOR2_X1 U1097 ( .A(n1010), .B(n1009), .Z(n1011) );
  XNOR2_X1 U1098 ( .A(n1012), .B(n1011), .ZN(n1016) );
  XOR2_X1 U1099 ( .A(KEYINPUT46), .B(KEYINPUT48), .Z(n1014) );
  XNOR2_X1 U1100 ( .A(G162), .B(KEYINPUT116), .ZN(n1013) );
  XNOR2_X1 U1101 ( .A(n1014), .B(n1013), .ZN(n1015) );
  XNOR2_X1 U1102 ( .A(n1016), .B(n1015), .ZN(n1021) );
  XOR2_X1 U1103 ( .A(G164), .B(n1017), .Z(n1018) );
  XNOR2_X1 U1104 ( .A(n1019), .B(n1018), .ZN(n1020) );
  XNOR2_X1 U1105 ( .A(n1021), .B(n1020), .ZN(n1024) );
  XNOR2_X1 U1106 ( .A(G160), .B(n1022), .ZN(n1023) );
  XNOR2_X1 U1107 ( .A(n1024), .B(n1023), .ZN(n1025) );
  NOR2_X1 U1108 ( .A1(G37), .A2(n1025), .ZN(G395) );
  XNOR2_X1 U1109 ( .A(n1027), .B(n1026), .ZN(n1030) );
  XOR2_X1 U1110 ( .A(G301), .B(n1028), .Z(n1029) );
  XNOR2_X1 U1111 ( .A(n1030), .B(n1029), .ZN(n1031) );
  XOR2_X1 U1112 ( .A(G286), .B(n1031), .Z(n1032) );
  NOR2_X1 U1113 ( .A1(G37), .A2(n1032), .ZN(G397) );
  OR2_X1 U1114 ( .A1(n1038), .A2(G401), .ZN(n1035) );
  NOR2_X1 U1115 ( .A1(G227), .A2(G229), .ZN(n1033) );
  XNOR2_X1 U1116 ( .A(KEYINPUT49), .B(n1033), .ZN(n1034) );
  NOR2_X1 U1117 ( .A1(n1035), .A2(n1034), .ZN(n1037) );
  NOR2_X1 U1118 ( .A1(G395), .A2(G397), .ZN(n1036) );
  NAND2_X1 U1119 ( .A1(n1037), .A2(n1036), .ZN(G225) );
  INV_X1 U1120 ( .A(G225), .ZN(G308) );
  INV_X1 U1121 ( .A(n1038), .ZN(G319) );
  INV_X1 U1122 ( .A(G69), .ZN(G235) );
endmodule

