//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 0 0 0 1 0 0 0 1 0 0 0 0 0 1 1 0 0 1 0 1 0 0 0 0 1 0 0 0 1 1 1 0 1 0 1 1 0 0 1 1 1 0 0 0 0 0 0 1 0 1 1 1 1 1 1 1 0 1 1 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:38:05 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n244, new_n245,
    new_n247, new_n248, new_n249, new_n250, new_n251, new_n252, new_n253,
    new_n254, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n822, new_n823, new_n824, new_n825, new_n826, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n901, new_n902, new_n903, new_n904, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n965, new_n966, new_n967, new_n968, new_n969,
    new_n970, new_n971, new_n972, new_n973, new_n974, new_n975, new_n976,
    new_n977, new_n978, new_n979, new_n980, new_n981, new_n982, new_n983,
    new_n984, new_n985, new_n986, new_n987, new_n988, new_n989, new_n990,
    new_n991, new_n992, new_n993, new_n994, new_n995, new_n997, new_n998,
    new_n999, new_n1000, new_n1001, new_n1002, new_n1003, new_n1004,
    new_n1005, new_n1006, new_n1007, new_n1008, new_n1009, new_n1010,
    new_n1011, new_n1012, new_n1013, new_n1014, new_n1015, new_n1016,
    new_n1017, new_n1018, new_n1019, new_n1020, new_n1022, new_n1023,
    new_n1024, new_n1025, new_n1026, new_n1027, new_n1028, new_n1029,
    new_n1030, new_n1031, new_n1032, new_n1033, new_n1034, new_n1035,
    new_n1036, new_n1037, new_n1038, new_n1039, new_n1040, new_n1041,
    new_n1042, new_n1043, new_n1044, new_n1045, new_n1046, new_n1047,
    new_n1048, new_n1049, new_n1050, new_n1051, new_n1052, new_n1053,
    new_n1054, new_n1055, new_n1056, new_n1057, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1076, new_n1077, new_n1078,
    new_n1079, new_n1080, new_n1081, new_n1082, new_n1083, new_n1084,
    new_n1085, new_n1086, new_n1087, new_n1088, new_n1089, new_n1090,
    new_n1091, new_n1092, new_n1093, new_n1094, new_n1095, new_n1096,
    new_n1097, new_n1098, new_n1099, new_n1100, new_n1101, new_n1102,
    new_n1103, new_n1104, new_n1105, new_n1106, new_n1107, new_n1108,
    new_n1109, new_n1110, new_n1111, new_n1112, new_n1113, new_n1114,
    new_n1115, new_n1116, new_n1117, new_n1118, new_n1119, new_n1120,
    new_n1121, new_n1122, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1145,
    new_n1146, new_n1147, new_n1148, new_n1149, new_n1150, new_n1151,
    new_n1152, new_n1153, new_n1154, new_n1155, new_n1156, new_n1157,
    new_n1158, new_n1159, new_n1160, new_n1161, new_n1162, new_n1163,
    new_n1164, new_n1165, new_n1166, new_n1167, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1183,
    new_n1184, new_n1185, new_n1187, new_n1188, new_n1189, new_n1190,
    new_n1191, new_n1192, new_n1193, new_n1194, new_n1195, new_n1196,
    new_n1197, new_n1198, new_n1199, new_n1200, new_n1201, new_n1202,
    new_n1203, new_n1204, new_n1205, new_n1206, new_n1207, new_n1208,
    new_n1209, new_n1210, new_n1211, new_n1212, new_n1213, new_n1214,
    new_n1215, new_n1216, new_n1217, new_n1218, new_n1219, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1231, new_n1232, new_n1233;
  INV_X1    g0000(.A(G50), .ZN(new_n201));
  INV_X1    g0001(.A(G58), .ZN(new_n202));
  INV_X1    g0002(.A(G68), .ZN(new_n203));
  NAND3_X1  g0003(.A1(new_n201), .A2(new_n202), .A3(new_n203), .ZN(new_n204));
  NOR2_X1   g0004(.A1(new_n204), .A2(G77), .ZN(G353));
  OAI21_X1  g0005(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  AOI21_X1  g0006(.A(KEYINPUT64), .B1(G1), .B2(G13), .ZN(new_n207));
  INV_X1    g0007(.A(new_n207), .ZN(new_n208));
  NAND3_X1  g0008(.A1(KEYINPUT64), .A2(G1), .A3(G13), .ZN(new_n209));
  NAND2_X1  g0009(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  INV_X1    g0010(.A(G20), .ZN(new_n211));
  NOR2_X1   g0011(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  NAND2_X1  g0012(.A1(new_n202), .A2(new_n203), .ZN(new_n213));
  NAND2_X1  g0013(.A1(new_n213), .A2(G50), .ZN(new_n214));
  INV_X1    g0014(.A(new_n214), .ZN(new_n215));
  NAND2_X1  g0015(.A1(new_n212), .A2(new_n215), .ZN(new_n216));
  INV_X1    g0016(.A(G1), .ZN(new_n217));
  NOR2_X1   g0017(.A1(new_n217), .A2(new_n211), .ZN(new_n218));
  INV_X1    g0018(.A(G13), .ZN(new_n219));
  NAND2_X1  g0019(.A1(new_n218), .A2(new_n219), .ZN(new_n220));
  INV_X1    g0020(.A(new_n220), .ZN(new_n221));
  OAI211_X1 g0021(.A(new_n221), .B(G250), .C1(G257), .C2(G264), .ZN(new_n222));
  INV_X1    g0022(.A(KEYINPUT0), .ZN(new_n223));
  OAI21_X1  g0023(.A(new_n216), .B1(new_n222), .B2(new_n223), .ZN(new_n224));
  AOI22_X1  g0024(.A1(G50), .A2(G226), .B1(G77), .B2(G244), .ZN(new_n225));
  INV_X1    g0025(.A(G116), .ZN(new_n226));
  INV_X1    g0026(.A(G270), .ZN(new_n227));
  OAI21_X1  g0027(.A(new_n225), .B1(new_n226), .B2(new_n227), .ZN(new_n228));
  AOI22_X1  g0028(.A1(G87), .A2(G250), .B1(G107), .B2(G264), .ZN(new_n229));
  NAND2_X1  g0029(.A1(G97), .A2(G257), .ZN(new_n230));
  INV_X1    g0030(.A(G238), .ZN(new_n231));
  OAI211_X1 g0031(.A(new_n229), .B(new_n230), .C1(new_n203), .C2(new_n231), .ZN(new_n232));
  AOI211_X1 g0032(.A(new_n228), .B(new_n232), .C1(G58), .C2(G232), .ZN(new_n233));
  NOR2_X1   g0033(.A1(new_n233), .A2(new_n218), .ZN(new_n234));
  XOR2_X1   g0034(.A(new_n234), .B(KEYINPUT1), .Z(new_n235));
  AOI211_X1 g0035(.A(new_n224), .B(new_n235), .C1(new_n223), .C2(new_n222), .ZN(G361));
  XOR2_X1   g0036(.A(G238), .B(G244), .Z(new_n237));
  XNOR2_X1  g0037(.A(new_n237), .B(G232), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n238), .B(KEYINPUT2), .ZN(new_n239));
  INV_X1    g0039(.A(G226), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XNOR2_X1  g0041(.A(G250), .B(G257), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n242), .B(KEYINPUT65), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n243), .B(G264), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n244), .B(new_n227), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n241), .B(new_n245), .ZN(G358));
  XNOR2_X1  g0046(.A(G50), .B(G68), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n247), .B(G58), .ZN(new_n248));
  INV_X1    g0048(.A(G77), .ZN(new_n249));
  XNOR2_X1  g0049(.A(new_n248), .B(new_n249), .ZN(new_n250));
  XOR2_X1   g0050(.A(G107), .B(G116), .Z(new_n251));
  XOR2_X1   g0051(.A(G87), .B(G97), .Z(new_n252));
  XNOR2_X1  g0052(.A(new_n251), .B(new_n252), .ZN(new_n253));
  INV_X1    g0053(.A(new_n253), .ZN(new_n254));
  XNOR2_X1  g0054(.A(new_n250), .B(new_n254), .ZN(G351));
  XNOR2_X1  g0055(.A(KEYINPUT3), .B(G33), .ZN(new_n256));
  INV_X1    g0056(.A(G1698), .ZN(new_n257));
  NAND3_X1  g0057(.A1(new_n256), .A2(G226), .A3(new_n257), .ZN(new_n258));
  NAND3_X1  g0058(.A1(new_n256), .A2(G232), .A3(G1698), .ZN(new_n259));
  NAND2_X1  g0059(.A1(G33), .A2(G97), .ZN(new_n260));
  NAND3_X1  g0060(.A1(new_n258), .A2(new_n259), .A3(new_n260), .ZN(new_n261));
  AOI21_X1  g0061(.A(new_n210), .B1(G33), .B2(G41), .ZN(new_n262));
  NAND2_X1  g0062(.A1(new_n261), .A2(new_n262), .ZN(new_n263));
  INV_X1    g0063(.A(G41), .ZN(new_n264));
  INV_X1    g0064(.A(G45), .ZN(new_n265));
  AOI21_X1  g0065(.A(G1), .B1(new_n264), .B2(new_n265), .ZN(new_n266));
  INV_X1    g0066(.A(KEYINPUT66), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n266), .A2(new_n267), .ZN(new_n268));
  INV_X1    g0068(.A(G33), .ZN(new_n269));
  OAI211_X1 g0069(.A(G1), .B(G13), .C1(new_n269), .C2(new_n264), .ZN(new_n270));
  OAI21_X1  g0070(.A(new_n217), .B1(G41), .B2(G45), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n271), .A2(KEYINPUT66), .ZN(new_n272));
  NAND3_X1  g0072(.A1(new_n268), .A2(new_n270), .A3(new_n272), .ZN(new_n273));
  INV_X1    g0073(.A(new_n273), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n274), .A2(G238), .ZN(new_n275));
  INV_X1    g0075(.A(G274), .ZN(new_n276));
  NOR2_X1   g0076(.A1(new_n271), .A2(new_n276), .ZN(new_n277));
  INV_X1    g0077(.A(new_n277), .ZN(new_n278));
  NAND3_X1  g0078(.A1(new_n263), .A2(new_n275), .A3(new_n278), .ZN(new_n279));
  NAND2_X1  g0079(.A1(new_n279), .A2(KEYINPUT13), .ZN(new_n280));
  AOI21_X1  g0080(.A(new_n277), .B1(new_n261), .B2(new_n262), .ZN(new_n281));
  INV_X1    g0081(.A(KEYINPUT13), .ZN(new_n282));
  NAND3_X1  g0082(.A1(new_n281), .A2(new_n282), .A3(new_n275), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n280), .A2(new_n283), .ZN(new_n284));
  INV_X1    g0084(.A(KEYINPUT75), .ZN(new_n285));
  NAND3_X1  g0085(.A1(new_n284), .A2(new_n285), .A3(G169), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n286), .A2(KEYINPUT14), .ZN(new_n287));
  NAND3_X1  g0087(.A1(new_n280), .A2(G179), .A3(new_n283), .ZN(new_n288));
  INV_X1    g0088(.A(KEYINPUT14), .ZN(new_n289));
  NAND4_X1  g0089(.A1(new_n284), .A2(new_n285), .A3(new_n289), .A4(G169), .ZN(new_n290));
  NAND3_X1  g0090(.A1(new_n287), .A2(new_n288), .A3(new_n290), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n203), .A2(G20), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n211), .A2(G33), .ZN(new_n293));
  NOR2_X1   g0093(.A1(G20), .A2(G33), .ZN(new_n294));
  INV_X1    g0094(.A(new_n294), .ZN(new_n295));
  OAI221_X1 g0095(.A(new_n292), .B1(new_n293), .B2(new_n249), .C1(new_n295), .C2(new_n201), .ZN(new_n296));
  NAND3_X1  g0096(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n297));
  AND3_X1   g0097(.A1(KEYINPUT64), .A2(G1), .A3(G13), .ZN(new_n298));
  OAI21_X1  g0098(.A(new_n297), .B1(new_n298), .B2(new_n207), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n299), .A2(KEYINPUT67), .ZN(new_n300));
  INV_X1    g0100(.A(KEYINPUT67), .ZN(new_n301));
  OAI211_X1 g0101(.A(new_n301), .B(new_n297), .C1(new_n298), .C2(new_n207), .ZN(new_n302));
  NAND3_X1  g0102(.A1(new_n296), .A2(new_n300), .A3(new_n302), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n303), .A2(KEYINPUT11), .ZN(new_n304));
  INV_X1    g0104(.A(KEYINPUT11), .ZN(new_n305));
  NAND4_X1  g0105(.A1(new_n296), .A2(new_n300), .A3(new_n305), .A4(new_n302), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n304), .A2(new_n306), .ZN(new_n307));
  NAND3_X1  g0107(.A1(new_n217), .A2(G13), .A3(G20), .ZN(new_n308));
  NAND4_X1  g0108(.A1(new_n210), .A2(KEYINPUT69), .A3(new_n308), .A4(new_n297), .ZN(new_n309));
  INV_X1    g0109(.A(KEYINPUT69), .ZN(new_n310));
  INV_X1    g0110(.A(new_n308), .ZN(new_n311));
  OAI21_X1  g0111(.A(new_n310), .B1(new_n299), .B2(new_n311), .ZN(new_n312));
  AOI22_X1  g0112(.A1(new_n309), .A2(new_n312), .B1(new_n217), .B2(G20), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n313), .A2(G68), .ZN(new_n314));
  AOI211_X1 g0114(.A(G68), .B(new_n308), .C1(KEYINPUT71), .C2(KEYINPUT12), .ZN(new_n315));
  NOR2_X1   g0115(.A1(KEYINPUT71), .A2(KEYINPUT12), .ZN(new_n316));
  XNOR2_X1  g0116(.A(new_n315), .B(new_n316), .ZN(new_n317));
  NAND3_X1  g0117(.A1(new_n307), .A2(new_n314), .A3(new_n317), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n318), .A2(KEYINPUT72), .ZN(new_n319));
  AOI22_X1  g0119(.A1(new_n304), .A2(new_n306), .B1(new_n313), .B2(G68), .ZN(new_n320));
  INV_X1    g0120(.A(KEYINPUT72), .ZN(new_n321));
  NAND3_X1  g0121(.A1(new_n320), .A2(new_n321), .A3(new_n317), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n319), .A2(new_n322), .ZN(new_n323));
  INV_X1    g0123(.A(new_n323), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n291), .A2(new_n324), .ZN(new_n325));
  INV_X1    g0125(.A(new_n283), .ZN(new_n326));
  AOI21_X1  g0126(.A(new_n282), .B1(new_n281), .B2(new_n275), .ZN(new_n327));
  OAI21_X1  g0127(.A(G200), .B1(new_n326), .B2(new_n327), .ZN(new_n328));
  NAND3_X1  g0128(.A1(new_n280), .A2(G190), .A3(new_n283), .ZN(new_n329));
  NOR2_X1   g0129(.A1(new_n318), .A2(KEYINPUT72), .ZN(new_n330));
  AOI21_X1  g0130(.A(new_n321), .B1(new_n320), .B2(new_n317), .ZN(new_n331));
  OAI211_X1 g0131(.A(new_n328), .B(new_n329), .C1(new_n330), .C2(new_n331), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n332), .A2(KEYINPUT73), .ZN(new_n333));
  INV_X1    g0133(.A(KEYINPUT73), .ZN(new_n334));
  NAND4_X1  g0134(.A1(new_n323), .A2(new_n334), .A3(new_n328), .A4(new_n329), .ZN(new_n335));
  AND3_X1   g0135(.A1(new_n333), .A2(KEYINPUT74), .A3(new_n335), .ZN(new_n336));
  AOI21_X1  g0136(.A(KEYINPUT74), .B1(new_n333), .B2(new_n335), .ZN(new_n337));
  OAI21_X1  g0137(.A(new_n325), .B1(new_n336), .B2(new_n337), .ZN(new_n338));
  INV_X1    g0138(.A(new_n338), .ZN(new_n339));
  NAND3_X1  g0139(.A1(new_n256), .A2(G222), .A3(new_n257), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n256), .A2(G1698), .ZN(new_n341));
  INV_X1    g0141(.A(G223), .ZN(new_n342));
  OAI221_X1 g0142(.A(new_n340), .B1(new_n249), .B2(new_n256), .C1(new_n341), .C2(new_n342), .ZN(new_n343));
  AOI21_X1  g0143(.A(new_n277), .B1(new_n343), .B2(new_n262), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n274), .A2(G226), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n344), .A2(new_n345), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n346), .A2(G200), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n347), .A2(KEYINPUT70), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n348), .A2(KEYINPUT10), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n300), .A2(new_n302), .ZN(new_n350));
  INV_X1    g0150(.A(new_n350), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n204), .A2(G20), .ZN(new_n352));
  INV_X1    g0152(.A(G150), .ZN(new_n353));
  XNOR2_X1  g0153(.A(KEYINPUT8), .B(G58), .ZN(new_n354));
  OAI221_X1 g0154(.A(new_n352), .B1(new_n353), .B2(new_n295), .C1(new_n293), .C2(new_n354), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n351), .A2(new_n355), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n311), .A2(new_n201), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n217), .A2(G20), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n358), .A2(G50), .ZN(new_n359));
  XNOR2_X1  g0159(.A(new_n359), .B(KEYINPUT68), .ZN(new_n360));
  NAND3_X1  g0160(.A1(new_n350), .A2(new_n360), .A3(new_n308), .ZN(new_n361));
  NAND3_X1  g0161(.A1(new_n356), .A2(new_n357), .A3(new_n361), .ZN(new_n362));
  INV_X1    g0162(.A(KEYINPUT9), .ZN(new_n363));
  AOI22_X1  g0163(.A1(G200), .A2(new_n346), .B1(new_n362), .B2(new_n363), .ZN(new_n364));
  NAND3_X1  g0164(.A1(new_n344), .A2(G190), .A3(new_n345), .ZN(new_n365));
  INV_X1    g0165(.A(new_n362), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n366), .A2(KEYINPUT9), .ZN(new_n367));
  NAND4_X1  g0167(.A1(new_n349), .A2(new_n364), .A3(new_n365), .A4(new_n367), .ZN(new_n368));
  NAND3_X1  g0168(.A1(new_n364), .A2(new_n365), .A3(new_n367), .ZN(new_n369));
  NAND3_X1  g0169(.A1(new_n369), .A2(KEYINPUT10), .A3(new_n348), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n368), .A2(new_n370), .ZN(new_n371));
  INV_X1    g0171(.A(G169), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n346), .A2(new_n372), .ZN(new_n373));
  INV_X1    g0173(.A(G179), .ZN(new_n374));
  NAND3_X1  g0174(.A1(new_n344), .A2(new_n374), .A3(new_n345), .ZN(new_n375));
  NAND3_X1  g0175(.A1(new_n373), .A2(new_n362), .A3(new_n375), .ZN(new_n376));
  NAND3_X1  g0176(.A1(new_n256), .A2(G232), .A3(new_n257), .ZN(new_n377));
  INV_X1    g0177(.A(G107), .ZN(new_n378));
  OAI221_X1 g0178(.A(new_n377), .B1(new_n378), .B2(new_n256), .C1(new_n341), .C2(new_n231), .ZN(new_n379));
  AOI21_X1  g0179(.A(new_n277), .B1(new_n379), .B2(new_n262), .ZN(new_n380));
  INV_X1    g0180(.A(G244), .ZN(new_n381));
  OAI21_X1  g0181(.A(new_n380), .B1(new_n381), .B2(new_n273), .ZN(new_n382));
  OR2_X1    g0182(.A1(new_n382), .A2(G179), .ZN(new_n383));
  INV_X1    g0183(.A(new_n354), .ZN(new_n384));
  AOI22_X1  g0184(.A1(new_n384), .A2(new_n294), .B1(G20), .B2(G77), .ZN(new_n385));
  XOR2_X1   g0185(.A(KEYINPUT15), .B(G87), .Z(new_n386));
  NAND3_X1  g0186(.A1(new_n386), .A2(new_n211), .A3(G33), .ZN(new_n387));
  AOI22_X1  g0187(.A1(new_n385), .A2(new_n387), .B1(new_n210), .B2(new_n297), .ZN(new_n388));
  AOI21_X1  g0188(.A(new_n388), .B1(new_n313), .B2(G77), .ZN(new_n389));
  OAI21_X1  g0189(.A(new_n389), .B1(G77), .B2(new_n308), .ZN(new_n390));
  NAND2_X1  g0190(.A1(new_n382), .A2(new_n372), .ZN(new_n391));
  NAND3_X1  g0191(.A1(new_n383), .A2(new_n390), .A3(new_n391), .ZN(new_n392));
  INV_X1    g0192(.A(new_n390), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n382), .A2(G200), .ZN(new_n394));
  INV_X1    g0194(.A(G190), .ZN(new_n395));
  OAI211_X1 g0195(.A(new_n393), .B(new_n394), .C1(new_n395), .C2(new_n382), .ZN(new_n396));
  AND4_X1   g0196(.A1(new_n371), .A2(new_n376), .A3(new_n392), .A4(new_n396), .ZN(new_n397));
  OR2_X1    g0197(.A1(KEYINPUT3), .A2(G33), .ZN(new_n398));
  NAND2_X1  g0198(.A1(KEYINPUT3), .A2(G33), .ZN(new_n399));
  NAND3_X1  g0199(.A1(new_n398), .A2(new_n211), .A3(new_n399), .ZN(new_n400));
  INV_X1    g0200(.A(KEYINPUT7), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n400), .A2(new_n401), .ZN(new_n402));
  NAND4_X1  g0202(.A1(new_n398), .A2(KEYINPUT7), .A3(new_n211), .A4(new_n399), .ZN(new_n403));
  AOI21_X1  g0203(.A(new_n203), .B1(new_n402), .B2(new_n403), .ZN(new_n404));
  INV_X1    g0204(.A(G159), .ZN(new_n405));
  NOR2_X1   g0205(.A1(new_n295), .A2(new_n405), .ZN(new_n406));
  NAND2_X1  g0206(.A1(G58), .A2(G68), .ZN(new_n407));
  AOI21_X1  g0207(.A(new_n211), .B1(new_n213), .B2(new_n407), .ZN(new_n408));
  NOR3_X1   g0208(.A1(new_n404), .A2(new_n406), .A3(new_n408), .ZN(new_n409));
  OAI21_X1  g0209(.A(KEYINPUT76), .B1(new_n409), .B2(KEYINPUT16), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n409), .A2(KEYINPUT16), .ZN(new_n411));
  AND2_X1   g0211(.A1(KEYINPUT3), .A2(G33), .ZN(new_n412));
  NOR2_X1   g0212(.A1(KEYINPUT3), .A2(G33), .ZN(new_n413));
  NOR2_X1   g0213(.A1(new_n412), .A2(new_n413), .ZN(new_n414));
  AOI21_X1  g0214(.A(KEYINPUT7), .B1(new_n414), .B2(new_n211), .ZN(new_n415));
  INV_X1    g0215(.A(new_n403), .ZN(new_n416));
  OAI21_X1  g0216(.A(G68), .B1(new_n415), .B2(new_n416), .ZN(new_n417));
  INV_X1    g0217(.A(new_n406), .ZN(new_n418));
  INV_X1    g0218(.A(new_n408), .ZN(new_n419));
  NAND3_X1  g0219(.A1(new_n417), .A2(new_n418), .A3(new_n419), .ZN(new_n420));
  INV_X1    g0220(.A(KEYINPUT76), .ZN(new_n421));
  INV_X1    g0221(.A(KEYINPUT16), .ZN(new_n422));
  NAND3_X1  g0222(.A1(new_n420), .A2(new_n421), .A3(new_n422), .ZN(new_n423));
  NAND4_X1  g0223(.A1(new_n410), .A2(new_n299), .A3(new_n411), .A4(new_n423), .ZN(new_n424));
  NAND3_X1  g0224(.A1(new_n256), .A2(G223), .A3(new_n257), .ZN(new_n425));
  INV_X1    g0225(.A(G87), .ZN(new_n426));
  OAI221_X1 g0226(.A(new_n425), .B1(new_n269), .B2(new_n426), .C1(new_n341), .C2(new_n240), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n427), .A2(new_n262), .ZN(new_n428));
  NAND4_X1  g0228(.A1(new_n268), .A2(G232), .A3(new_n272), .A4(new_n270), .ZN(new_n429));
  INV_X1    g0229(.A(KEYINPUT78), .ZN(new_n430));
  NAND3_X1  g0230(.A1(new_n429), .A2(new_n430), .A3(new_n278), .ZN(new_n431));
  INV_X1    g0231(.A(new_n431), .ZN(new_n432));
  AOI21_X1  g0232(.A(new_n430), .B1(new_n429), .B2(new_n278), .ZN(new_n433));
  OAI21_X1  g0233(.A(new_n428), .B1(new_n432), .B2(new_n433), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n434), .A2(G200), .ZN(new_n435));
  INV_X1    g0235(.A(new_n433), .ZN(new_n436));
  AOI22_X1  g0236(.A1(new_n436), .A2(new_n431), .B1(new_n262), .B2(new_n427), .ZN(new_n437));
  NAND2_X1  g0237(.A1(new_n437), .A2(G190), .ZN(new_n438));
  NOR2_X1   g0238(.A1(new_n351), .A2(new_n354), .ZN(new_n439));
  AOI22_X1  g0239(.A1(new_n439), .A2(new_n358), .B1(new_n311), .B2(new_n354), .ZN(new_n440));
  NAND4_X1  g0240(.A1(new_n424), .A2(new_n435), .A3(new_n438), .A4(new_n440), .ZN(new_n441));
  OR2_X1    g0241(.A1(new_n441), .A2(KEYINPUT17), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n441), .A2(KEYINPUT17), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n434), .A2(G169), .ZN(new_n445));
  OAI21_X1  g0245(.A(new_n445), .B1(new_n374), .B2(new_n434), .ZN(new_n446));
  NAND3_X1  g0246(.A1(new_n424), .A2(KEYINPUT77), .A3(new_n440), .ZN(new_n447));
  INV_X1    g0247(.A(new_n447), .ZN(new_n448));
  AOI21_X1  g0248(.A(KEYINPUT77), .B1(new_n424), .B2(new_n440), .ZN(new_n449));
  OAI21_X1  g0249(.A(new_n446), .B1(new_n448), .B2(new_n449), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n450), .A2(KEYINPUT18), .ZN(new_n451));
  INV_X1    g0251(.A(KEYINPUT18), .ZN(new_n452));
  OAI211_X1 g0252(.A(new_n452), .B(new_n446), .C1(new_n448), .C2(new_n449), .ZN(new_n453));
  AND2_X1   g0253(.A1(new_n451), .A2(new_n453), .ZN(new_n454));
  NAND4_X1  g0254(.A1(new_n339), .A2(new_n397), .A3(new_n444), .A4(new_n454), .ZN(new_n455));
  NAND3_X1  g0255(.A1(new_n256), .A2(G257), .A3(new_n257), .ZN(new_n456));
  NAND3_X1  g0256(.A1(new_n256), .A2(G264), .A3(G1698), .ZN(new_n457));
  INV_X1    g0257(.A(G303), .ZN(new_n458));
  OAI211_X1 g0258(.A(new_n456), .B(new_n457), .C1(new_n458), .C2(new_n256), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n459), .A2(new_n262), .ZN(new_n460));
  NOR2_X1   g0260(.A1(new_n265), .A2(G1), .ZN(new_n461));
  NAND2_X1  g0261(.A1(new_n461), .A2(G274), .ZN(new_n462));
  AND2_X1   g0262(.A1(KEYINPUT5), .A2(G41), .ZN(new_n463));
  NOR2_X1   g0263(.A1(KEYINPUT5), .A2(G41), .ZN(new_n464));
  NOR2_X1   g0264(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  OAI21_X1  g0265(.A(KEYINPUT80), .B1(new_n462), .B2(new_n465), .ZN(new_n466));
  XNOR2_X1  g0266(.A(KEYINPUT5), .B(G41), .ZN(new_n467));
  INV_X1    g0267(.A(KEYINPUT80), .ZN(new_n468));
  NAND4_X1  g0268(.A1(new_n467), .A2(new_n468), .A3(G274), .A4(new_n461), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n466), .A2(new_n469), .ZN(new_n470));
  NAND2_X1  g0270(.A1(G1), .A2(G13), .ZN(new_n471));
  AOI21_X1  g0271(.A(new_n471), .B1(G33), .B2(G41), .ZN(new_n472));
  AOI21_X1  g0272(.A(new_n472), .B1(new_n461), .B2(new_n467), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n473), .A2(G270), .ZN(new_n474));
  NAND3_X1  g0274(.A1(new_n460), .A2(new_n470), .A3(new_n474), .ZN(new_n475));
  AND2_X1   g0275(.A1(new_n475), .A2(G169), .ZN(new_n476));
  NAND2_X1  g0276(.A1(G33), .A2(G283), .ZN(new_n477));
  INV_X1    g0277(.A(G97), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n478), .A2(KEYINPUT79), .ZN(new_n479));
  INV_X1    g0279(.A(KEYINPUT79), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n480), .A2(G97), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n479), .A2(new_n481), .ZN(new_n482));
  OAI211_X1 g0282(.A(new_n211), .B(new_n477), .C1(new_n482), .C2(G33), .ZN(new_n483));
  XNOR2_X1  g0283(.A(KEYINPUT84), .B(G116), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n484), .A2(G20), .ZN(new_n485));
  NAND3_X1  g0285(.A1(new_n483), .A2(new_n299), .A3(new_n485), .ZN(new_n486));
  INV_X1    g0286(.A(KEYINPUT20), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n486), .A2(new_n487), .ZN(new_n488));
  NAND4_X1  g0288(.A1(new_n483), .A2(KEYINPUT20), .A3(new_n299), .A4(new_n485), .ZN(new_n489));
  AOI22_X1  g0289(.A1(new_n488), .A2(new_n489), .B1(new_n311), .B2(new_n484), .ZN(new_n490));
  NOR2_X1   g0290(.A1(new_n269), .A2(G1), .ZN(new_n491));
  AOI21_X1  g0291(.A(new_n491), .B1(new_n309), .B2(new_n312), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n492), .A2(G116), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n490), .A2(new_n493), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n476), .A2(new_n494), .ZN(new_n495));
  INV_X1    g0295(.A(KEYINPUT21), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  INV_X1    g0297(.A(new_n497), .ZN(new_n498));
  AND3_X1   g0298(.A1(new_n460), .A2(new_n470), .A3(new_n474), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n499), .A2(G179), .ZN(new_n500));
  NAND3_X1  g0300(.A1(new_n475), .A2(KEYINPUT21), .A3(G169), .ZN(new_n501));
  AND2_X1   g0301(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  INV_X1    g0302(.A(new_n494), .ZN(new_n503));
  OAI21_X1  g0303(.A(KEYINPUT85), .B1(new_n502), .B2(new_n503), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n500), .A2(new_n501), .ZN(new_n505));
  INV_X1    g0305(.A(KEYINPUT85), .ZN(new_n506));
  NAND3_X1  g0306(.A1(new_n505), .A2(new_n506), .A3(new_n494), .ZN(new_n507));
  AOI21_X1  g0307(.A(new_n498), .B1(new_n504), .B2(new_n507), .ZN(new_n508));
  NAND3_X1  g0308(.A1(new_n256), .A2(G257), .A3(G1698), .ZN(new_n509));
  NAND3_X1  g0309(.A1(new_n256), .A2(G250), .A3(new_n257), .ZN(new_n510));
  XNOR2_X1  g0310(.A(KEYINPUT86), .B(G294), .ZN(new_n511));
  OAI211_X1 g0311(.A(new_n509), .B(new_n510), .C1(new_n269), .C2(new_n511), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n512), .A2(new_n262), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n473), .A2(G264), .ZN(new_n514));
  NAND3_X1  g0314(.A1(new_n513), .A2(new_n470), .A3(new_n514), .ZN(new_n515));
  INV_X1    g0315(.A(new_n515), .ZN(new_n516));
  OAI21_X1  g0316(.A(KEYINPUT87), .B1(new_n516), .B2(new_n372), .ZN(new_n517));
  OR2_X1    g0317(.A1(new_n515), .A2(new_n374), .ZN(new_n518));
  INV_X1    g0318(.A(KEYINPUT87), .ZN(new_n519));
  NAND3_X1  g0319(.A1(new_n515), .A2(new_n519), .A3(G169), .ZN(new_n520));
  NAND3_X1  g0320(.A1(new_n517), .A2(new_n518), .A3(new_n520), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n521), .A2(KEYINPUT88), .ZN(new_n522));
  NAND3_X1  g0322(.A1(new_n256), .A2(KEYINPUT22), .A3(G87), .ZN(new_n523));
  OAI21_X1  g0323(.A(new_n523), .B1(new_n269), .B2(new_n484), .ZN(new_n524));
  INV_X1    g0324(.A(KEYINPUT22), .ZN(new_n525));
  NAND3_X1  g0325(.A1(new_n256), .A2(new_n211), .A3(G87), .ZN(new_n526));
  AOI22_X1  g0326(.A1(new_n524), .A2(new_n211), .B1(new_n525), .B2(new_n526), .ZN(new_n527));
  INV_X1    g0327(.A(KEYINPUT24), .ZN(new_n528));
  NOR2_X1   g0328(.A1(new_n211), .A2(G107), .ZN(new_n529));
  XNOR2_X1  g0329(.A(new_n529), .B(KEYINPUT23), .ZN(new_n530));
  AND3_X1   g0330(.A1(new_n527), .A2(new_n528), .A3(new_n530), .ZN(new_n531));
  AOI21_X1  g0331(.A(new_n528), .B1(new_n527), .B2(new_n530), .ZN(new_n532));
  OAI21_X1  g0332(.A(new_n299), .B1(new_n531), .B2(new_n532), .ZN(new_n533));
  AOI211_X1 g0333(.A(new_n311), .B(new_n491), .C1(new_n300), .C2(new_n302), .ZN(new_n534));
  NAND2_X1  g0334(.A1(new_n534), .A2(G107), .ZN(new_n535));
  NOR2_X1   g0335(.A1(new_n308), .A2(G107), .ZN(new_n536));
  XNOR2_X1  g0336(.A(new_n536), .B(KEYINPUT25), .ZN(new_n537));
  NAND3_X1  g0337(.A1(new_n533), .A2(new_n535), .A3(new_n537), .ZN(new_n538));
  INV_X1    g0338(.A(KEYINPUT88), .ZN(new_n539));
  NAND4_X1  g0339(.A1(new_n517), .A2(new_n518), .A3(new_n539), .A4(new_n520), .ZN(new_n540));
  NAND3_X1  g0340(.A1(new_n522), .A2(new_n538), .A3(new_n540), .ZN(new_n541));
  NAND3_X1  g0341(.A1(new_n256), .A2(new_n211), .A3(G68), .ZN(new_n542));
  INV_X1    g0342(.A(KEYINPUT19), .ZN(new_n543));
  OAI21_X1  g0343(.A(new_n543), .B1(new_n482), .B2(new_n293), .ZN(new_n544));
  XNOR2_X1  g0344(.A(KEYINPUT79), .B(G97), .ZN(new_n545));
  NOR3_X1   g0345(.A1(new_n545), .A2(G87), .A3(G107), .ZN(new_n546));
  NOR2_X1   g0346(.A1(new_n260), .A2(new_n543), .ZN(new_n547));
  NOR2_X1   g0347(.A1(new_n547), .A2(G20), .ZN(new_n548));
  OAI211_X1 g0348(.A(new_n542), .B(new_n544), .C1(new_n546), .C2(new_n548), .ZN(new_n549));
  INV_X1    g0349(.A(new_n386), .ZN(new_n550));
  AOI22_X1  g0350(.A1(new_n549), .A2(new_n299), .B1(new_n311), .B2(new_n550), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n534), .A2(new_n386), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  OAI211_X1 g0353(.A(G244), .B(G1698), .C1(new_n412), .C2(new_n413), .ZN(new_n554));
  OAI211_X1 g0354(.A(G238), .B(new_n257), .C1(new_n412), .C2(new_n413), .ZN(new_n555));
  OAI211_X1 g0355(.A(new_n554), .B(new_n555), .C1(new_n269), .C2(new_n484), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n262), .A2(new_n556), .ZN(new_n557));
  OAI211_X1 g0357(.A(new_n270), .B(G250), .C1(G1), .C2(new_n265), .ZN(new_n558));
  NAND3_X1  g0358(.A1(new_n557), .A2(new_n462), .A3(new_n558), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n559), .A2(new_n372), .ZN(new_n560));
  NAND4_X1  g0360(.A1(new_n557), .A2(new_n374), .A3(new_n462), .A4(new_n558), .ZN(new_n561));
  NAND3_X1  g0361(.A1(new_n553), .A2(new_n560), .A3(new_n561), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n559), .A2(G200), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n534), .A2(G87), .ZN(new_n564));
  NAND4_X1  g0364(.A1(new_n557), .A2(G190), .A3(new_n462), .A4(new_n558), .ZN(new_n565));
  NAND4_X1  g0365(.A1(new_n563), .A2(new_n551), .A3(new_n564), .A4(new_n565), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n562), .A2(new_n566), .ZN(new_n567));
  INV_X1    g0367(.A(new_n567), .ZN(new_n568));
  AND3_X1   g0368(.A1(new_n508), .A2(new_n541), .A3(new_n568), .ZN(new_n569));
  OAI211_X1 g0369(.A(G244), .B(new_n257), .C1(new_n412), .C2(new_n413), .ZN(new_n570));
  INV_X1    g0370(.A(KEYINPUT4), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n570), .A2(new_n571), .ZN(new_n572));
  NAND4_X1  g0372(.A1(new_n256), .A2(KEYINPUT4), .A3(G244), .A4(new_n257), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n572), .A2(new_n573), .ZN(new_n574));
  NAND3_X1  g0374(.A1(new_n256), .A2(G250), .A3(G1698), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n575), .A2(new_n477), .ZN(new_n576));
  OAI21_X1  g0376(.A(new_n262), .B1(new_n574), .B2(new_n576), .ZN(new_n577));
  INV_X1    g0377(.A(KEYINPUT81), .ZN(new_n578));
  AOI22_X1  g0378(.A1(new_n473), .A2(G257), .B1(new_n466), .B2(new_n469), .ZN(new_n579));
  AND3_X1   g0379(.A1(new_n577), .A2(new_n578), .A3(new_n579), .ZN(new_n580));
  AOI21_X1  g0380(.A(new_n578), .B1(new_n577), .B2(new_n579), .ZN(new_n581));
  OAI21_X1  g0381(.A(G190), .B1(new_n580), .B2(new_n581), .ZN(new_n582));
  INV_X1    g0382(.A(KEYINPUT82), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  OAI211_X1 g0384(.A(KEYINPUT82), .B(G190), .C1(new_n580), .C2(new_n581), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n584), .A2(new_n585), .ZN(new_n586));
  XOR2_X1   g0386(.A(G97), .B(G107), .Z(new_n587));
  NAND2_X1  g0387(.A1(new_n378), .A2(KEYINPUT6), .ZN(new_n588));
  OAI22_X1  g0388(.A1(new_n587), .A2(KEYINPUT6), .B1(new_n482), .B2(new_n588), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n589), .A2(G20), .ZN(new_n590));
  OAI21_X1  g0390(.A(G107), .B1(new_n415), .B2(new_n416), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n294), .A2(G77), .ZN(new_n592));
  NAND3_X1  g0392(.A1(new_n590), .A2(new_n591), .A3(new_n592), .ZN(new_n593));
  AOI22_X1  g0393(.A1(new_n593), .A2(new_n299), .B1(new_n534), .B2(G97), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n577), .A2(new_n579), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n595), .A2(G200), .ZN(new_n596));
  OAI211_X1 g0396(.A(new_n594), .B(new_n596), .C1(G97), .C2(new_n308), .ZN(new_n597));
  INV_X1    g0397(.A(new_n597), .ZN(new_n598));
  AOI21_X1  g0398(.A(KEYINPUT83), .B1(new_n586), .B2(new_n598), .ZN(new_n599));
  INV_X1    g0399(.A(KEYINPUT83), .ZN(new_n600));
  AOI211_X1 g0400(.A(new_n600), .B(new_n597), .C1(new_n584), .C2(new_n585), .ZN(new_n601));
  OAI21_X1  g0401(.A(new_n594), .B1(G97), .B2(new_n308), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n595), .A2(KEYINPUT81), .ZN(new_n603));
  NAND3_X1  g0403(.A1(new_n577), .A2(new_n578), .A3(new_n579), .ZN(new_n604));
  NAND3_X1  g0404(.A1(new_n603), .A2(new_n372), .A3(new_n604), .ZN(new_n605));
  NAND3_X1  g0405(.A1(new_n577), .A2(new_n374), .A3(new_n579), .ZN(new_n606));
  AND3_X1   g0406(.A1(new_n602), .A2(new_n605), .A3(new_n606), .ZN(new_n607));
  NOR3_X1   g0407(.A1(new_n599), .A2(new_n601), .A3(new_n607), .ZN(new_n608));
  INV_X1    g0408(.A(new_n538), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n515), .A2(G200), .ZN(new_n610));
  OR2_X1    g0410(.A1(new_n515), .A2(new_n395), .ZN(new_n611));
  NAND3_X1  g0411(.A1(new_n609), .A2(new_n610), .A3(new_n611), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n499), .A2(G190), .ZN(new_n613));
  INV_X1    g0413(.A(G200), .ZN(new_n614));
  OAI211_X1 g0414(.A(new_n503), .B(new_n613), .C1(new_n614), .C2(new_n499), .ZN(new_n615));
  NAND4_X1  g0415(.A1(new_n569), .A2(new_n608), .A3(new_n612), .A4(new_n615), .ZN(new_n616));
  NOR2_X1   g0416(.A1(new_n455), .A2(new_n616), .ZN(G372));
  NAND2_X1  g0417(.A1(new_n424), .A2(new_n440), .ZN(new_n618));
  NAND3_X1  g0418(.A1(new_n618), .A2(KEYINPUT18), .A3(new_n446), .ZN(new_n619));
  INV_X1    g0419(.A(new_n619), .ZN(new_n620));
  AOI21_X1  g0420(.A(KEYINPUT18), .B1(new_n618), .B2(new_n446), .ZN(new_n621));
  NOR2_X1   g0421(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  AND2_X1   g0422(.A1(new_n333), .A2(new_n335), .ZN(new_n623));
  OAI21_X1  g0423(.A(new_n325), .B1(new_n623), .B2(new_n392), .ZN(new_n624));
  AOI21_X1  g0424(.A(new_n622), .B1(new_n624), .B2(new_n444), .ZN(new_n625));
  INV_X1    g0425(.A(KEYINPUT90), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n371), .A2(new_n626), .ZN(new_n627));
  NAND3_X1  g0427(.A1(new_n368), .A2(new_n370), .A3(KEYINPUT90), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  OR2_X1    g0429(.A1(new_n625), .A2(new_n629), .ZN(new_n630));
  AND2_X1   g0430(.A1(new_n630), .A2(new_n376), .ZN(new_n631));
  INV_X1    g0431(.A(new_n455), .ZN(new_n632));
  INV_X1    g0432(.A(KEYINPUT26), .ZN(new_n633));
  INV_X1    g0433(.A(KEYINPUT89), .ZN(new_n634));
  AND3_X1   g0434(.A1(new_n562), .A2(new_n634), .A3(new_n566), .ZN(new_n635));
  AOI21_X1  g0435(.A(new_n634), .B1(new_n562), .B2(new_n566), .ZN(new_n636));
  OAI211_X1 g0436(.A(new_n607), .B(new_n633), .C1(new_n635), .C2(new_n636), .ZN(new_n637));
  NAND3_X1  g0437(.A1(new_n602), .A2(new_n605), .A3(new_n606), .ZN(new_n638));
  OAI21_X1  g0438(.A(KEYINPUT26), .B1(new_n638), .B2(new_n567), .ZN(new_n639));
  AND3_X1   g0439(.A1(new_n637), .A2(new_n562), .A3(new_n639), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n603), .A2(new_n604), .ZN(new_n641));
  AOI21_X1  g0441(.A(KEYINPUT82), .B1(new_n641), .B2(G190), .ZN(new_n642));
  INV_X1    g0442(.A(new_n585), .ZN(new_n643));
  OAI21_X1  g0443(.A(new_n598), .B1(new_n642), .B2(new_n643), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n644), .A2(new_n600), .ZN(new_n645));
  NAND3_X1  g0445(.A1(new_n586), .A2(KEYINPUT83), .A3(new_n598), .ZN(new_n646));
  NAND4_X1  g0446(.A1(new_n645), .A2(new_n612), .A3(new_n638), .A4(new_n646), .ZN(new_n647));
  OR2_X1    g0447(.A1(new_n635), .A2(new_n636), .ZN(new_n648));
  AND2_X1   g0448(.A1(new_n538), .A2(new_n521), .ZN(new_n649));
  OAI21_X1  g0449(.A(new_n497), .B1(new_n503), .B2(new_n502), .ZN(new_n650));
  OAI21_X1  g0450(.A(new_n648), .B1(new_n649), .B2(new_n650), .ZN(new_n651));
  OAI21_X1  g0451(.A(new_n640), .B1(new_n647), .B2(new_n651), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n632), .A2(new_n652), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n631), .A2(new_n653), .ZN(G369));
  NOR2_X1   g0454(.A1(new_n219), .A2(G20), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n655), .A2(new_n217), .ZN(new_n656));
  OR2_X1    g0456(.A1(new_n656), .A2(KEYINPUT27), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n656), .A2(KEYINPUT27), .ZN(new_n658));
  AND3_X1   g0458(.A1(new_n657), .A2(G213), .A3(new_n658), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n659), .A2(G343), .ZN(new_n660));
  XNOR2_X1  g0460(.A(new_n660), .B(KEYINPUT91), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n661), .A2(new_n494), .ZN(new_n662));
  OAI21_X1  g0462(.A(new_n615), .B1(new_n650), .B2(new_n662), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n504), .A2(new_n507), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n664), .A2(new_n497), .ZN(new_n665));
  AOI21_X1  g0465(.A(new_n663), .B1(new_n665), .B2(new_n662), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n666), .A2(G330), .ZN(new_n667));
  INV_X1    g0467(.A(new_n667), .ZN(new_n668));
  INV_X1    g0468(.A(new_n661), .ZN(new_n669));
  OAI211_X1 g0469(.A(new_n541), .B(new_n612), .C1(new_n609), .C2(new_n669), .ZN(new_n670));
  NAND4_X1  g0470(.A1(new_n522), .A2(new_n538), .A3(new_n540), .A4(new_n661), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n668), .A2(new_n672), .ZN(new_n673));
  NOR2_X1   g0473(.A1(new_n508), .A2(new_n661), .ZN(new_n674));
  AOI22_X1  g0474(.A1(new_n672), .A2(new_n674), .B1(new_n649), .B2(new_n669), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n673), .A2(new_n675), .ZN(G399));
  NOR2_X1   g0476(.A1(new_n220), .A2(G41), .ZN(new_n677));
  INV_X1    g0477(.A(new_n677), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n678), .A2(G1), .ZN(new_n679));
  NAND4_X1  g0479(.A1(new_n482), .A2(new_n426), .A3(new_n378), .A4(new_n226), .ZN(new_n680));
  OAI22_X1  g0480(.A1(new_n679), .A2(new_n680), .B1(new_n214), .B2(new_n678), .ZN(new_n681));
  XNOR2_X1  g0481(.A(new_n681), .B(KEYINPUT28), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n652), .A2(new_n669), .ZN(new_n683));
  NOR2_X1   g0483(.A1(new_n683), .A2(KEYINPUT29), .ZN(new_n684));
  NAND3_X1  g0484(.A1(new_n607), .A2(new_n568), .A3(new_n633), .ZN(new_n685));
  INV_X1    g0485(.A(new_n562), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n648), .A2(new_n607), .ZN(new_n687));
  AOI21_X1  g0487(.A(new_n686), .B1(new_n687), .B2(KEYINPUT26), .ZN(new_n688));
  NOR2_X1   g0488(.A1(new_n599), .A2(new_n601), .ZN(new_n689));
  NAND4_X1  g0489(.A1(new_n689), .A2(new_n638), .A3(new_n612), .A4(new_n648), .ZN(new_n690));
  AND2_X1   g0490(.A1(new_n508), .A2(new_n541), .ZN(new_n691));
  OAI211_X1 g0491(.A(new_n685), .B(new_n688), .C1(new_n690), .C2(new_n691), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n692), .A2(new_n669), .ZN(new_n693));
  AOI21_X1  g0493(.A(new_n684), .B1(KEYINPUT29), .B2(new_n693), .ZN(new_n694));
  NOR2_X1   g0494(.A1(new_n500), .A2(new_n559), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n513), .A2(new_n514), .ZN(new_n696));
  INV_X1    g0496(.A(KEYINPUT30), .ZN(new_n697));
  AOI21_X1  g0497(.A(new_n696), .B1(KEYINPUT93), .B2(new_n697), .ZN(new_n698));
  NAND3_X1  g0498(.A1(new_n695), .A2(new_n641), .A3(new_n698), .ZN(new_n699));
  OR3_X1    g0499(.A1(new_n699), .A2(KEYINPUT93), .A3(new_n697), .ZN(new_n700));
  NAND3_X1  g0500(.A1(new_n475), .A2(new_n374), .A3(new_n559), .ZN(new_n701));
  INV_X1    g0501(.A(KEYINPUT92), .ZN(new_n702));
  OR2_X1    g0502(.A1(new_n701), .A2(new_n702), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n701), .A2(new_n702), .ZN(new_n704));
  NAND4_X1  g0504(.A1(new_n703), .A2(new_n595), .A3(new_n515), .A4(new_n704), .ZN(new_n705));
  OAI21_X1  g0505(.A(new_n699), .B1(KEYINPUT93), .B2(new_n697), .ZN(new_n706));
  NAND3_X1  g0506(.A1(new_n700), .A2(new_n705), .A3(new_n706), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n707), .A2(new_n661), .ZN(new_n708));
  INV_X1    g0508(.A(KEYINPUT31), .ZN(new_n709));
  NAND2_X1  g0509(.A1(new_n708), .A2(new_n709), .ZN(new_n710));
  NAND3_X1  g0510(.A1(new_n707), .A2(KEYINPUT31), .A3(new_n661), .ZN(new_n711));
  OAI211_X1 g0511(.A(new_n710), .B(new_n711), .C1(new_n616), .C2(new_n661), .ZN(new_n712));
  NAND2_X1  g0512(.A1(new_n712), .A2(G330), .ZN(new_n713));
  AND2_X1   g0513(.A1(new_n694), .A2(new_n713), .ZN(new_n714));
  OAI21_X1  g0514(.A(new_n682), .B1(new_n714), .B2(G1), .ZN(G364));
  NOR2_X1   g0515(.A1(new_n666), .A2(G330), .ZN(new_n716));
  XOR2_X1   g0516(.A(new_n716), .B(KEYINPUT94), .Z(new_n717));
  AOI21_X1  g0517(.A(new_n217), .B1(new_n655), .B2(G45), .ZN(new_n718));
  INV_X1    g0518(.A(new_n718), .ZN(new_n719));
  NOR2_X1   g0519(.A1(new_n677), .A2(new_n719), .ZN(new_n720));
  INV_X1    g0520(.A(new_n720), .ZN(new_n721));
  NAND3_X1  g0521(.A1(new_n717), .A2(new_n667), .A3(new_n721), .ZN(new_n722));
  OR2_X1    g0522(.A1(new_n372), .A2(KEYINPUT97), .ZN(new_n723));
  NAND2_X1  g0523(.A1(new_n372), .A2(KEYINPUT97), .ZN(new_n724));
  NAND3_X1  g0524(.A1(new_n723), .A2(new_n724), .A3(G20), .ZN(new_n725));
  NAND3_X1  g0525(.A1(new_n725), .A2(new_n208), .A3(new_n209), .ZN(new_n726));
  XNOR2_X1  g0526(.A(new_n726), .B(KEYINPUT98), .ZN(new_n727));
  NOR2_X1   g0527(.A1(new_n211), .A2(G179), .ZN(new_n728));
  NOR2_X1   g0528(.A1(new_n614), .A2(G190), .ZN(new_n729));
  NAND2_X1  g0529(.A1(new_n728), .A2(new_n729), .ZN(new_n730));
  NOR2_X1   g0530(.A1(new_n730), .A2(new_n378), .ZN(new_n731));
  NOR2_X1   g0531(.A1(new_n211), .A2(new_n374), .ZN(new_n732));
  NOR2_X1   g0532(.A1(G190), .A2(G200), .ZN(new_n733));
  NAND2_X1  g0533(.A1(new_n732), .A2(new_n733), .ZN(new_n734));
  INV_X1    g0534(.A(new_n734), .ZN(new_n735));
  AOI21_X1  g0535(.A(new_n731), .B1(G77), .B2(new_n735), .ZN(new_n736));
  NOR2_X1   g0536(.A1(new_n395), .A2(new_n614), .ZN(new_n737));
  NAND2_X1  g0537(.A1(new_n737), .A2(new_n732), .ZN(new_n738));
  OAI21_X1  g0538(.A(new_n736), .B1(new_n201), .B2(new_n738), .ZN(new_n739));
  NAND2_X1  g0539(.A1(new_n732), .A2(new_n729), .ZN(new_n740));
  OR2_X1    g0540(.A1(new_n740), .A2(KEYINPUT99), .ZN(new_n741));
  NAND2_X1  g0541(.A1(new_n740), .A2(KEYINPUT99), .ZN(new_n742));
  NAND2_X1  g0542(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  AOI21_X1  g0543(.A(new_n739), .B1(G68), .B2(new_n743), .ZN(new_n744));
  NAND2_X1  g0544(.A1(new_n728), .A2(new_n733), .ZN(new_n745));
  INV_X1    g0545(.A(new_n745), .ZN(new_n746));
  NAND2_X1  g0546(.A1(new_n746), .A2(G159), .ZN(new_n747));
  XNOR2_X1  g0547(.A(new_n747), .B(KEYINPUT32), .ZN(new_n748));
  NAND2_X1  g0548(.A1(new_n737), .A2(new_n728), .ZN(new_n749));
  INV_X1    g0549(.A(new_n749), .ZN(new_n750));
  AOI21_X1  g0550(.A(new_n748), .B1(G87), .B2(new_n750), .ZN(new_n751));
  NAND3_X1  g0551(.A1(new_n732), .A2(G190), .A3(new_n614), .ZN(new_n752));
  INV_X1    g0552(.A(new_n752), .ZN(new_n753));
  NAND2_X1  g0553(.A1(new_n753), .A2(G58), .ZN(new_n754));
  NOR3_X1   g0554(.A1(new_n395), .A2(G179), .A3(G200), .ZN(new_n755));
  NOR2_X1   g0555(.A1(new_n755), .A2(new_n211), .ZN(new_n756));
  NOR2_X1   g0556(.A1(new_n756), .A2(new_n478), .ZN(new_n757));
  NOR2_X1   g0557(.A1(new_n757), .A2(new_n414), .ZN(new_n758));
  NAND4_X1  g0558(.A1(new_n744), .A2(new_n751), .A3(new_n754), .A4(new_n758), .ZN(new_n759));
  NOR2_X1   g0559(.A1(new_n756), .A2(new_n511), .ZN(new_n760));
  INV_X1    g0560(.A(G329), .ZN(new_n761));
  INV_X1    g0561(.A(G311), .ZN(new_n762));
  OAI221_X1 g0562(.A(new_n414), .B1(new_n745), .B2(new_n761), .C1(new_n762), .C2(new_n734), .ZN(new_n763));
  INV_X1    g0563(.A(new_n738), .ZN(new_n764));
  AOI211_X1 g0564(.A(new_n760), .B(new_n763), .C1(G326), .C2(new_n764), .ZN(new_n765));
  INV_X1    g0565(.A(G322), .ZN(new_n766));
  INV_X1    g0566(.A(G283), .ZN(new_n767));
  OAI22_X1  g0567(.A1(new_n752), .A2(new_n766), .B1(new_n730), .B2(new_n767), .ZN(new_n768));
  XNOR2_X1  g0568(.A(KEYINPUT100), .B(G317), .ZN(new_n769));
  XNOR2_X1  g0569(.A(new_n769), .B(KEYINPUT33), .ZN(new_n770));
  AOI21_X1  g0570(.A(new_n768), .B1(new_n743), .B2(new_n770), .ZN(new_n771));
  OAI211_X1 g0571(.A(new_n765), .B(new_n771), .C1(new_n458), .C2(new_n749), .ZN(new_n772));
  AOI21_X1  g0572(.A(new_n727), .B1(new_n759), .B2(new_n772), .ZN(new_n773));
  INV_X1    g0573(.A(new_n727), .ZN(new_n774));
  NAND2_X1  g0574(.A1(new_n219), .A2(new_n269), .ZN(new_n775));
  XNOR2_X1  g0575(.A(new_n775), .B(KEYINPUT96), .ZN(new_n776));
  NOR2_X1   g0576(.A1(new_n776), .A2(G20), .ZN(new_n777));
  NOR2_X1   g0577(.A1(new_n774), .A2(new_n777), .ZN(new_n778));
  NOR2_X1   g0578(.A1(new_n220), .A2(new_n256), .ZN(new_n779));
  NAND2_X1  g0579(.A1(new_n215), .A2(new_n265), .ZN(new_n780));
  OAI211_X1 g0580(.A(new_n779), .B(new_n780), .C1(new_n250), .C2(new_n265), .ZN(new_n781));
  NOR2_X1   g0581(.A1(new_n220), .A2(new_n414), .ZN(new_n782));
  XNOR2_X1  g0582(.A(new_n782), .B(KEYINPUT95), .ZN(new_n783));
  NAND2_X1  g0583(.A1(new_n783), .A2(G355), .ZN(new_n784));
  OAI211_X1 g0584(.A(new_n781), .B(new_n784), .C1(G116), .C2(new_n221), .ZN(new_n785));
  AOI21_X1  g0585(.A(new_n773), .B1(new_n778), .B2(new_n785), .ZN(new_n786));
  XNOR2_X1  g0586(.A(new_n777), .B(KEYINPUT101), .ZN(new_n787));
  INV_X1    g0587(.A(new_n787), .ZN(new_n788));
  OAI211_X1 g0588(.A(new_n720), .B(new_n786), .C1(new_n666), .C2(new_n788), .ZN(new_n789));
  NAND2_X1  g0589(.A1(new_n722), .A2(new_n789), .ZN(G396));
  OAI211_X1 g0590(.A(new_n396), .B(new_n392), .C1(new_n393), .C2(new_n669), .ZN(new_n791));
  XNOR2_X1  g0591(.A(new_n791), .B(KEYINPUT103), .ZN(new_n792));
  INV_X1    g0592(.A(new_n792), .ZN(new_n793));
  OAI21_X1  g0593(.A(new_n793), .B1(new_n392), .B2(new_n669), .ZN(new_n794));
  MUX2_X1   g0594(.A(new_n793), .B(new_n794), .S(new_n683), .Z(new_n795));
  XNOR2_X1  g0595(.A(new_n795), .B(new_n713), .ZN(new_n796));
  NAND2_X1  g0596(.A1(new_n796), .A2(new_n721), .ZN(new_n797));
  AOI22_X1  g0597(.A1(new_n753), .A2(G143), .B1(new_n735), .B2(G159), .ZN(new_n798));
  INV_X1    g0598(.A(G137), .ZN(new_n799));
  INV_X1    g0599(.A(new_n743), .ZN(new_n800));
  OAI221_X1 g0600(.A(new_n798), .B1(new_n799), .B2(new_n738), .C1(new_n800), .C2(new_n353), .ZN(new_n801));
  XNOR2_X1  g0601(.A(new_n801), .B(KEYINPUT34), .ZN(new_n802));
  NAND3_X1  g0602(.A1(new_n728), .A2(new_n729), .A3(G68), .ZN(new_n803));
  INV_X1    g0603(.A(G132), .ZN(new_n804));
  OAI221_X1 g0604(.A(new_n256), .B1(new_n745), .B2(new_n804), .C1(new_n201), .C2(new_n749), .ZN(new_n805));
  INV_X1    g0605(.A(new_n756), .ZN(new_n806));
  AOI21_X1  g0606(.A(new_n805), .B1(G58), .B2(new_n806), .ZN(new_n807));
  NAND3_X1  g0607(.A1(new_n802), .A2(new_n803), .A3(new_n807), .ZN(new_n808));
  NOR2_X1   g0608(.A1(new_n749), .A2(new_n378), .ZN(new_n809));
  OAI21_X1  g0609(.A(new_n414), .B1(new_n730), .B2(new_n426), .ZN(new_n810));
  AOI211_X1 g0610(.A(new_n810), .B(new_n757), .C1(G294), .C2(new_n753), .ZN(new_n811));
  OAI22_X1  g0611(.A1(new_n738), .A2(new_n458), .B1(new_n745), .B2(new_n762), .ZN(new_n812));
  AOI21_X1  g0612(.A(new_n812), .B1(new_n743), .B2(G283), .ZN(new_n813));
  OAI211_X1 g0613(.A(new_n811), .B(new_n813), .C1(new_n484), .C2(new_n734), .ZN(new_n814));
  OAI21_X1  g0614(.A(new_n808), .B1(new_n809), .B2(new_n814), .ZN(new_n815));
  NAND2_X1  g0615(.A1(new_n727), .A2(new_n776), .ZN(new_n816));
  XOR2_X1   g0616(.A(new_n816), .B(KEYINPUT102), .Z(new_n817));
  INV_X1    g0617(.A(new_n817), .ZN(new_n818));
  AOI22_X1  g0618(.A1(new_n815), .A2(new_n774), .B1(new_n249), .B2(new_n818), .ZN(new_n819));
  OAI211_X1 g0619(.A(new_n720), .B(new_n819), .C1(new_n794), .C2(new_n776), .ZN(new_n820));
  NAND2_X1  g0620(.A1(new_n797), .A2(new_n820), .ZN(G384));
  NAND2_X1  g0621(.A1(new_n333), .A2(new_n335), .ZN(new_n822));
  NAND2_X1  g0622(.A1(new_n324), .A2(new_n661), .ZN(new_n823));
  AND3_X1   g0623(.A1(new_n325), .A2(new_n822), .A3(new_n823), .ZN(new_n824));
  INV_X1    g0624(.A(new_n823), .ZN(new_n825));
  AOI21_X1  g0625(.A(new_n824), .B1(new_n338), .B2(new_n825), .ZN(new_n826));
  INV_X1    g0626(.A(new_n826), .ZN(new_n827));
  AND3_X1   g0627(.A1(new_n712), .A2(new_n794), .A3(new_n827), .ZN(new_n828));
  INV_X1    g0628(.A(KEYINPUT104), .ZN(new_n829));
  NAND2_X1  g0629(.A1(new_n618), .A2(new_n446), .ZN(new_n830));
  NAND2_X1  g0630(.A1(new_n830), .A2(new_n452), .ZN(new_n831));
  AOI22_X1  g0631(.A1(new_n443), .A2(new_n442), .B1(new_n831), .B2(new_n619), .ZN(new_n832));
  INV_X1    g0632(.A(new_n659), .ZN(new_n833));
  INV_X1    g0633(.A(new_n449), .ZN(new_n834));
  AOI21_X1  g0634(.A(new_n833), .B1(new_n834), .B2(new_n447), .ZN(new_n835));
  INV_X1    g0635(.A(new_n835), .ZN(new_n836));
  OAI21_X1  g0636(.A(new_n829), .B1(new_n832), .B2(new_n836), .ZN(new_n837));
  XOR2_X1   g0637(.A(new_n441), .B(KEYINPUT17), .Z(new_n838));
  OAI211_X1 g0638(.A(KEYINPUT104), .B(new_n835), .C1(new_n838), .C2(new_n622), .ZN(new_n839));
  NAND2_X1  g0639(.A1(new_n830), .A2(new_n441), .ZN(new_n840));
  OAI21_X1  g0640(.A(KEYINPUT37), .B1(new_n835), .B2(new_n840), .ZN(new_n841));
  OAI22_X1  g0641(.A1(new_n448), .A2(new_n449), .B1(new_n446), .B2(new_n659), .ZN(new_n842));
  INV_X1    g0642(.A(KEYINPUT37), .ZN(new_n843));
  AND2_X1   g0643(.A1(new_n441), .A2(new_n843), .ZN(new_n844));
  NAND2_X1  g0644(.A1(new_n842), .A2(new_n844), .ZN(new_n845));
  NAND2_X1  g0645(.A1(new_n841), .A2(new_n845), .ZN(new_n846));
  NAND3_X1  g0646(.A1(new_n837), .A2(new_n839), .A3(new_n846), .ZN(new_n847));
  INV_X1    g0647(.A(KEYINPUT38), .ZN(new_n848));
  NAND2_X1  g0648(.A1(new_n847), .A2(new_n848), .ZN(new_n849));
  INV_X1    g0649(.A(KEYINPUT105), .ZN(new_n850));
  NAND3_X1  g0650(.A1(new_n451), .A2(new_n444), .A3(new_n453), .ZN(new_n851));
  NAND2_X1  g0651(.A1(new_n420), .A2(new_n422), .ZN(new_n852));
  NAND3_X1  g0652(.A1(new_n411), .A2(new_n852), .A3(new_n351), .ZN(new_n853));
  NAND2_X1  g0653(.A1(new_n853), .A2(new_n440), .ZN(new_n854));
  NAND2_X1  g0654(.A1(new_n854), .A2(new_n659), .ZN(new_n855));
  INV_X1    g0655(.A(new_n855), .ZN(new_n856));
  NAND2_X1  g0656(.A1(new_n851), .A2(new_n856), .ZN(new_n857));
  NAND2_X1  g0657(.A1(new_n446), .A2(new_n854), .ZN(new_n858));
  NAND3_X1  g0658(.A1(new_n858), .A2(new_n441), .A3(new_n855), .ZN(new_n859));
  AOI22_X1  g0659(.A1(new_n842), .A2(new_n844), .B1(new_n859), .B2(KEYINPUT37), .ZN(new_n860));
  INV_X1    g0660(.A(new_n860), .ZN(new_n861));
  NAND3_X1  g0661(.A1(new_n857), .A2(KEYINPUT38), .A3(new_n861), .ZN(new_n862));
  AND3_X1   g0662(.A1(new_n849), .A2(new_n850), .A3(new_n862), .ZN(new_n863));
  AOI21_X1  g0663(.A(new_n850), .B1(new_n849), .B2(new_n862), .ZN(new_n864));
  OAI211_X1 g0664(.A(new_n828), .B(KEYINPUT40), .C1(new_n863), .C2(new_n864), .ZN(new_n865));
  INV_X1    g0665(.A(KEYINPUT40), .ZN(new_n866));
  NAND3_X1  g0666(.A1(new_n712), .A2(new_n794), .A3(new_n827), .ZN(new_n867));
  AOI21_X1  g0667(.A(KEYINPUT38), .B1(new_n857), .B2(new_n861), .ZN(new_n868));
  AOI211_X1 g0668(.A(new_n848), .B(new_n860), .C1(new_n851), .C2(new_n856), .ZN(new_n869));
  NOR2_X1   g0669(.A1(new_n868), .A2(new_n869), .ZN(new_n870));
  OAI21_X1  g0670(.A(new_n866), .B1(new_n867), .B2(new_n870), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n865), .A2(new_n871), .ZN(new_n872));
  AND2_X1   g0672(.A1(new_n632), .A2(new_n712), .ZN(new_n873));
  XNOR2_X1  g0673(.A(new_n872), .B(new_n873), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n874), .A2(G330), .ZN(new_n875));
  INV_X1    g0675(.A(KEYINPUT39), .ZN(new_n876));
  NAND3_X1  g0676(.A1(new_n849), .A2(new_n876), .A3(new_n862), .ZN(new_n877));
  OAI21_X1  g0677(.A(KEYINPUT39), .B1(new_n868), .B2(new_n869), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n877), .A2(new_n878), .ZN(new_n879));
  NOR2_X1   g0679(.A1(new_n325), .A2(new_n661), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n879), .A2(new_n880), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n622), .A2(new_n833), .ZN(new_n882));
  INV_X1    g0682(.A(new_n870), .ZN(new_n883));
  NAND3_X1  g0683(.A1(new_n652), .A2(new_n669), .A3(new_n792), .ZN(new_n884));
  NOR2_X1   g0684(.A1(new_n392), .A2(new_n661), .ZN(new_n885));
  INV_X1    g0685(.A(new_n885), .ZN(new_n886));
  AOI21_X1  g0686(.A(new_n826), .B1(new_n884), .B2(new_n886), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n883), .A2(new_n887), .ZN(new_n888));
  NAND3_X1  g0688(.A1(new_n881), .A2(new_n882), .A3(new_n888), .ZN(new_n889));
  OAI21_X1  g0689(.A(new_n631), .B1(new_n694), .B2(new_n455), .ZN(new_n890));
  XOR2_X1   g0690(.A(new_n889), .B(new_n890), .Z(new_n891));
  XNOR2_X1  g0691(.A(new_n875), .B(new_n891), .ZN(new_n892));
  OAI21_X1  g0692(.A(new_n892), .B1(new_n217), .B2(new_n655), .ZN(new_n893));
  AOI21_X1  g0693(.A(new_n226), .B1(new_n589), .B2(KEYINPUT35), .ZN(new_n894));
  OAI211_X1 g0694(.A(new_n894), .B(new_n212), .C1(KEYINPUT35), .C2(new_n589), .ZN(new_n895));
  XNOR2_X1  g0695(.A(new_n895), .B(KEYINPUT36), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n407), .A2(G77), .ZN(new_n897));
  OAI22_X1  g0697(.A1(new_n214), .A2(new_n897), .B1(G50), .B2(new_n203), .ZN(new_n898));
  NAND3_X1  g0698(.A1(new_n898), .A2(G1), .A3(new_n219), .ZN(new_n899));
  NAND3_X1  g0699(.A1(new_n893), .A2(new_n896), .A3(new_n899), .ZN(G367));
  NAND2_X1  g0700(.A1(new_n551), .A2(new_n564), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n661), .A2(new_n901), .ZN(new_n902));
  XNOR2_X1  g0702(.A(new_n902), .B(KEYINPUT106), .ZN(new_n903));
  AOI21_X1  g0703(.A(KEYINPUT107), .B1(new_n648), .B2(new_n903), .ZN(new_n904));
  NOR2_X1   g0704(.A1(new_n903), .A2(new_n562), .ZN(new_n905));
  MUX2_X1   g0705(.A(new_n904), .B(KEYINPUT107), .S(new_n905), .Z(new_n906));
  NAND2_X1  g0706(.A1(new_n906), .A2(new_n787), .ZN(new_n907));
  INV_X1    g0707(.A(new_n779), .ZN(new_n908));
  OAI221_X1 g0708(.A(new_n778), .B1(new_n221), .B2(new_n550), .C1(new_n245), .C2(new_n908), .ZN(new_n909));
  NOR2_X1   g0709(.A1(new_n756), .A2(new_n203), .ZN(new_n910));
  INV_X1    g0710(.A(G143), .ZN(new_n911));
  OAI221_X1 g0711(.A(new_n256), .B1(new_n749), .B2(new_n202), .C1(new_n911), .C2(new_n738), .ZN(new_n912));
  AOI211_X1 g0712(.A(new_n910), .B(new_n912), .C1(G50), .C2(new_n735), .ZN(new_n913));
  OAI22_X1  g0713(.A1(new_n730), .A2(new_n249), .B1(new_n745), .B2(new_n799), .ZN(new_n914));
  AOI21_X1  g0714(.A(new_n914), .B1(new_n743), .B2(G159), .ZN(new_n915));
  OAI211_X1 g0715(.A(new_n913), .B(new_n915), .C1(new_n353), .C2(new_n752), .ZN(new_n916));
  INV_X1    g0716(.A(new_n484), .ZN(new_n917));
  AOI21_X1  g0717(.A(KEYINPUT46), .B1(new_n750), .B2(new_n917), .ZN(new_n918));
  OAI221_X1 g0718(.A(new_n414), .B1(new_n730), .B2(new_n482), .C1(new_n762), .C2(new_n738), .ZN(new_n919));
  AOI211_X1 g0719(.A(new_n918), .B(new_n919), .C1(G107), .C2(new_n806), .ZN(new_n920));
  NAND2_X1  g0720(.A1(KEYINPUT46), .A2(G116), .ZN(new_n921));
  OAI22_X1  g0721(.A1(new_n767), .A2(new_n734), .B1(new_n749), .B2(new_n921), .ZN(new_n922));
  INV_X1    g0722(.A(new_n511), .ZN(new_n923));
  AOI21_X1  g0723(.A(new_n922), .B1(new_n743), .B2(new_n923), .ZN(new_n924));
  OAI211_X1 g0724(.A(new_n920), .B(new_n924), .C1(new_n458), .C2(new_n752), .ZN(new_n925));
  INV_X1    g0725(.A(G317), .ZN(new_n926));
  NOR2_X1   g0726(.A1(new_n745), .A2(new_n926), .ZN(new_n927));
  OAI21_X1  g0727(.A(new_n916), .B1(new_n925), .B2(new_n927), .ZN(new_n928));
  XNOR2_X1  g0728(.A(new_n928), .B(KEYINPUT47), .ZN(new_n929));
  AOI21_X1  g0729(.A(new_n721), .B1(new_n929), .B2(new_n774), .ZN(new_n930));
  NAND3_X1  g0730(.A1(new_n907), .A2(new_n909), .A3(new_n930), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n602), .A2(new_n661), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n608), .A2(new_n932), .ZN(new_n933));
  OAI21_X1  g0733(.A(new_n933), .B1(new_n638), .B2(new_n669), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n675), .A2(new_n934), .ZN(new_n935));
  XOR2_X1   g0735(.A(new_n935), .B(KEYINPUT45), .Z(new_n936));
  INV_X1    g0736(.A(KEYINPUT108), .ZN(new_n937));
  OAI211_X1 g0737(.A(new_n937), .B(KEYINPUT44), .C1(new_n675), .C2(new_n934), .ZN(new_n938));
  XOR2_X1   g0738(.A(KEYINPUT108), .B(KEYINPUT44), .Z(new_n939));
  OR3_X1    g0739(.A1(new_n675), .A2(new_n934), .A3(new_n939), .ZN(new_n940));
  NAND3_X1  g0740(.A1(new_n936), .A2(new_n938), .A3(new_n940), .ZN(new_n941));
  INV_X1    g0741(.A(new_n673), .ZN(new_n942));
  OR2_X1    g0742(.A1(new_n941), .A2(new_n942), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n941), .A2(new_n942), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n943), .A2(new_n944), .ZN(new_n945));
  XOR2_X1   g0745(.A(new_n667), .B(new_n672), .Z(new_n946));
  XNOR2_X1  g0746(.A(new_n946), .B(new_n674), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n947), .A2(new_n714), .ZN(new_n948));
  OAI21_X1  g0748(.A(new_n714), .B1(new_n945), .B2(new_n948), .ZN(new_n949));
  XNOR2_X1  g0749(.A(new_n677), .B(KEYINPUT41), .ZN(new_n950));
  AOI21_X1  g0750(.A(new_n719), .B1(new_n949), .B2(new_n950), .ZN(new_n951));
  NAND4_X1  g0751(.A1(new_n672), .A2(new_n608), .A3(new_n674), .A4(new_n932), .ZN(new_n952));
  XNOR2_X1  g0752(.A(new_n952), .B(KEYINPUT42), .ZN(new_n953));
  OR2_X1    g0753(.A1(new_n933), .A2(new_n541), .ZN(new_n954));
  AOI21_X1  g0754(.A(new_n661), .B1(new_n954), .B2(new_n638), .ZN(new_n955));
  INV_X1    g0755(.A(KEYINPUT43), .ZN(new_n956));
  OAI22_X1  g0756(.A1(new_n953), .A2(new_n955), .B1(new_n956), .B2(new_n906), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n942), .A2(new_n934), .ZN(new_n958));
  XNOR2_X1  g0758(.A(new_n957), .B(new_n958), .ZN(new_n959));
  NAND2_X1  g0759(.A1(new_n906), .A2(new_n956), .ZN(new_n960));
  XOR2_X1   g0760(.A(new_n959), .B(new_n960), .Z(new_n961));
  OAI21_X1  g0761(.A(new_n931), .B1(new_n951), .B2(new_n961), .ZN(new_n962));
  XNOR2_X1  g0762(.A(new_n962), .B(KEYINPUT109), .ZN(new_n963));
  INV_X1    g0763(.A(new_n963), .ZN(G387));
  NAND2_X1  g0764(.A1(new_n947), .A2(new_n719), .ZN(new_n965));
  XOR2_X1   g0765(.A(new_n965), .B(KEYINPUT110), .Z(new_n966));
  OR2_X1    g0766(.A1(new_n947), .A2(new_n714), .ZN(new_n967));
  NAND3_X1  g0767(.A1(new_n967), .A2(new_n677), .A3(new_n948), .ZN(new_n968));
  AOI22_X1  g0768(.A1(new_n753), .A2(G317), .B1(new_n764), .B2(G322), .ZN(new_n969));
  OAI221_X1 g0769(.A(new_n969), .B1(new_n458), .B2(new_n734), .C1(new_n800), .C2(new_n762), .ZN(new_n970));
  XNOR2_X1  g0770(.A(new_n970), .B(KEYINPUT48), .ZN(new_n971));
  OAI221_X1 g0771(.A(new_n971), .B1(new_n767), .B2(new_n756), .C1(new_n511), .C2(new_n749), .ZN(new_n972));
  XOR2_X1   g0772(.A(new_n972), .B(KEYINPUT112), .Z(new_n973));
  XNOR2_X1  g0773(.A(new_n973), .B(KEYINPUT49), .ZN(new_n974));
  AOI21_X1  g0774(.A(new_n256), .B1(new_n746), .B2(G326), .ZN(new_n975));
  OAI211_X1 g0775(.A(new_n974), .B(new_n975), .C1(new_n484), .C2(new_n730), .ZN(new_n976));
  NOR2_X1   g0776(.A1(new_n730), .A2(new_n478), .ZN(new_n977));
  OAI22_X1  g0777(.A1(new_n734), .A2(new_n203), .B1(new_n745), .B2(new_n353), .ZN(new_n978));
  AOI21_X1  g0778(.A(new_n978), .B1(new_n743), .B2(new_n384), .ZN(new_n979));
  NOR2_X1   g0779(.A1(new_n749), .A2(new_n249), .ZN(new_n980));
  AOI211_X1 g0780(.A(new_n414), .B(new_n980), .C1(G50), .C2(new_n753), .ZN(new_n981));
  AOI22_X1  g0781(.A1(new_n806), .A2(new_n386), .B1(new_n764), .B2(G159), .ZN(new_n982));
  NAND3_X1  g0782(.A1(new_n979), .A2(new_n981), .A3(new_n982), .ZN(new_n983));
  OAI21_X1  g0783(.A(new_n976), .B1(new_n977), .B2(new_n983), .ZN(new_n984));
  AOI21_X1  g0784(.A(new_n721), .B1(new_n984), .B2(new_n774), .ZN(new_n985));
  OAI21_X1  g0785(.A(new_n779), .B1(new_n241), .B2(new_n265), .ZN(new_n986));
  NOR2_X1   g0786(.A1(new_n354), .A2(G50), .ZN(new_n987));
  XNOR2_X1  g0787(.A(new_n987), .B(KEYINPUT50), .ZN(new_n988));
  OAI21_X1  g0788(.A(new_n988), .B1(new_n203), .B2(new_n249), .ZN(new_n989));
  NOR3_X1   g0789(.A1(new_n989), .A2(G45), .A3(new_n680), .ZN(new_n990));
  NOR2_X1   g0790(.A1(new_n986), .A2(new_n990), .ZN(new_n991));
  AOI22_X1  g0791(.A1(new_n783), .A2(new_n680), .B1(new_n378), .B2(new_n220), .ZN(new_n992));
  XNOR2_X1  g0792(.A(new_n992), .B(KEYINPUT111), .ZN(new_n993));
  OAI21_X1  g0793(.A(new_n778), .B1(new_n991), .B2(new_n993), .ZN(new_n994));
  OAI211_X1 g0794(.A(new_n985), .B(new_n994), .C1(new_n672), .C2(new_n788), .ZN(new_n995));
  NAND3_X1  g0795(.A1(new_n966), .A2(new_n968), .A3(new_n995), .ZN(G393));
  AOI21_X1  g0796(.A(new_n678), .B1(new_n945), .B2(new_n948), .ZN(new_n997));
  OAI21_X1  g0797(.A(new_n997), .B1(new_n945), .B2(new_n948), .ZN(new_n998));
  NAND3_X1  g0798(.A1(new_n943), .A2(new_n719), .A3(new_n944), .ZN(new_n999));
  OAI221_X1 g0799(.A(new_n778), .B1(new_n221), .B2(new_n482), .C1(new_n254), .C2(new_n908), .ZN(new_n1000));
  AOI22_X1  g0800(.A1(new_n743), .A2(G50), .B1(new_n384), .B2(new_n735), .ZN(new_n1001));
  XNOR2_X1  g0801(.A(new_n1001), .B(KEYINPUT113), .ZN(new_n1002));
  OAI22_X1  g0802(.A1(new_n752), .A2(new_n405), .B1(new_n738), .B2(new_n353), .ZN(new_n1003));
  XOR2_X1   g0803(.A(new_n1003), .B(KEYINPUT51), .Z(new_n1004));
  NOR2_X1   g0804(.A1(new_n756), .A2(new_n249), .ZN(new_n1005));
  OAI221_X1 g0805(.A(new_n256), .B1(new_n730), .B2(new_n426), .C1(new_n203), .C2(new_n749), .ZN(new_n1006));
  NOR3_X1   g0806(.A1(new_n1004), .A2(new_n1005), .A3(new_n1006), .ZN(new_n1007));
  OAI211_X1 g0807(.A(new_n1002), .B(new_n1007), .C1(new_n911), .C2(new_n745), .ZN(new_n1008));
  INV_X1    g0808(.A(G294), .ZN(new_n1009));
  OAI22_X1  g0809(.A1(new_n767), .A2(new_n749), .B1(new_n734), .B2(new_n1009), .ZN(new_n1010));
  AOI211_X1 g0810(.A(new_n731), .B(new_n1010), .C1(G322), .C2(new_n746), .ZN(new_n1011));
  OAI22_X1  g0811(.A1(new_n752), .A2(new_n762), .B1(new_n738), .B2(new_n926), .ZN(new_n1012));
  XNOR2_X1  g0812(.A(new_n1012), .B(KEYINPUT52), .ZN(new_n1013));
  NAND2_X1  g0813(.A1(new_n743), .A2(G303), .ZN(new_n1014));
  AOI21_X1  g0814(.A(new_n256), .B1(new_n806), .B2(new_n917), .ZN(new_n1015));
  NAND4_X1  g0815(.A1(new_n1011), .A2(new_n1013), .A3(new_n1014), .A4(new_n1015), .ZN(new_n1016));
  NAND2_X1  g0816(.A1(new_n1008), .A2(new_n1016), .ZN(new_n1017));
  AOI21_X1  g0817(.A(new_n721), .B1(new_n1017), .B2(new_n774), .ZN(new_n1018));
  INV_X1    g0818(.A(new_n777), .ZN(new_n1019));
  OAI211_X1 g0819(.A(new_n1000), .B(new_n1018), .C1(new_n934), .C2(new_n1019), .ZN(new_n1020));
  NAND3_X1  g0820(.A1(new_n998), .A2(new_n999), .A3(new_n1020), .ZN(G390));
  NAND3_X1  g0821(.A1(new_n632), .A2(G330), .A3(new_n712), .ZN(new_n1022));
  OAI211_X1 g0822(.A(new_n631), .B(new_n1022), .C1(new_n694), .C2(new_n455), .ZN(new_n1023));
  NAND3_X1  g0823(.A1(new_n712), .A2(new_n794), .A3(G330), .ZN(new_n1024));
  NAND2_X1  g0824(.A1(new_n1024), .A2(new_n826), .ZN(new_n1025));
  NAND4_X1  g0825(.A1(new_n712), .A2(new_n827), .A3(G330), .A4(new_n794), .ZN(new_n1026));
  NAND2_X1  g0826(.A1(new_n1025), .A2(new_n1026), .ZN(new_n1027));
  NAND2_X1  g0827(.A1(new_n884), .A2(new_n886), .ZN(new_n1028));
  NAND2_X1  g0828(.A1(new_n1027), .A2(new_n1028), .ZN(new_n1029));
  NAND3_X1  g0829(.A1(new_n692), .A2(new_n669), .A3(new_n792), .ZN(new_n1030));
  NAND4_X1  g0830(.A1(new_n1025), .A2(new_n886), .A3(new_n1030), .A4(new_n1026), .ZN(new_n1031));
  AOI21_X1  g0831(.A(new_n1023), .B1(new_n1029), .B2(new_n1031), .ZN(new_n1032));
  INV_X1    g0832(.A(new_n1032), .ZN(new_n1033));
  NAND2_X1  g0833(.A1(new_n1030), .A2(new_n886), .ZN(new_n1034));
  NAND2_X1  g0834(.A1(new_n1034), .A2(new_n827), .ZN(new_n1035));
  INV_X1    g0835(.A(new_n880), .ZN(new_n1036));
  OAI211_X1 g0836(.A(new_n1035), .B(new_n1036), .C1(new_n864), .C2(new_n863), .ZN(new_n1037));
  NAND2_X1  g0837(.A1(new_n1028), .A2(new_n827), .ZN(new_n1038));
  INV_X1    g0838(.A(KEYINPUT114), .ZN(new_n1039));
  NAND3_X1  g0839(.A1(new_n1038), .A2(new_n1039), .A3(new_n1036), .ZN(new_n1040));
  OAI21_X1  g0840(.A(KEYINPUT114), .B1(new_n887), .B2(new_n880), .ZN(new_n1041));
  NAND4_X1  g0841(.A1(new_n1040), .A2(new_n1041), .A3(new_n878), .A4(new_n877), .ZN(new_n1042));
  AOI21_X1  g0842(.A(new_n1026), .B1(new_n1037), .B2(new_n1042), .ZN(new_n1043));
  AND3_X1   g0843(.A1(new_n1037), .A2(new_n1042), .A3(new_n1026), .ZN(new_n1044));
  OAI21_X1  g0844(.A(new_n1033), .B1(new_n1043), .B2(new_n1044), .ZN(new_n1045));
  NAND2_X1  g0845(.A1(new_n1037), .A2(new_n1042), .ZN(new_n1046));
  INV_X1    g0846(.A(new_n1026), .ZN(new_n1047));
  NAND2_X1  g0847(.A1(new_n1046), .A2(new_n1047), .ZN(new_n1048));
  NAND3_X1  g0848(.A1(new_n1037), .A2(new_n1042), .A3(new_n1026), .ZN(new_n1049));
  NAND3_X1  g0849(.A1(new_n1048), .A2(new_n1049), .A3(new_n1032), .ZN(new_n1050));
  NAND3_X1  g0850(.A1(new_n1045), .A2(new_n677), .A3(new_n1050), .ZN(new_n1051));
  XOR2_X1   g0851(.A(KEYINPUT54), .B(G143), .Z(new_n1052));
  AOI22_X1  g0852(.A1(G128), .A2(new_n764), .B1(new_n735), .B2(new_n1052), .ZN(new_n1053));
  OAI221_X1 g0853(.A(new_n1053), .B1(new_n804), .B2(new_n752), .C1(new_n405), .C2(new_n756), .ZN(new_n1054));
  AOI21_X1  g0854(.A(new_n1054), .B1(G137), .B2(new_n743), .ZN(new_n1055));
  NOR2_X1   g0855(.A1(new_n749), .A2(new_n353), .ZN(new_n1056));
  XNOR2_X1  g0856(.A(new_n1056), .B(KEYINPUT53), .ZN(new_n1057));
  INV_X1    g0857(.A(G125), .ZN(new_n1058));
  OAI221_X1 g0858(.A(new_n256), .B1(new_n745), .B2(new_n1058), .C1(new_n201), .C2(new_n730), .ZN(new_n1059));
  XOR2_X1   g0859(.A(new_n1059), .B(KEYINPUT115), .Z(new_n1060));
  NAND3_X1  g0860(.A1(new_n1055), .A2(new_n1057), .A3(new_n1060), .ZN(new_n1061));
  AOI22_X1  g0861(.A1(new_n545), .A2(new_n735), .B1(new_n746), .B2(G294), .ZN(new_n1062));
  OAI221_X1 g0862(.A(new_n1062), .B1(new_n226), .B2(new_n752), .C1(new_n767), .C2(new_n738), .ZN(new_n1063));
  AOI21_X1  g0863(.A(new_n1063), .B1(G107), .B2(new_n743), .ZN(new_n1064));
  OAI21_X1  g0864(.A(new_n414), .B1(new_n749), .B2(new_n426), .ZN(new_n1065));
  XOR2_X1   g0865(.A(new_n1065), .B(KEYINPUT116), .Z(new_n1066));
  NAND3_X1  g0866(.A1(new_n1064), .A2(new_n803), .A3(new_n1066), .ZN(new_n1067));
  OAI21_X1  g0867(.A(new_n1061), .B1(new_n1067), .B2(new_n1005), .ZN(new_n1068));
  XOR2_X1   g0868(.A(new_n1068), .B(KEYINPUT117), .Z(new_n1069));
  OAI21_X1  g0869(.A(new_n720), .B1(new_n1069), .B2(new_n727), .ZN(new_n1070));
  NOR2_X1   g0870(.A1(new_n879), .A2(new_n776), .ZN(new_n1071));
  AOI211_X1 g0871(.A(new_n1070), .B(new_n1071), .C1(new_n354), .C2(new_n818), .ZN(new_n1072));
  NOR2_X1   g0872(.A1(new_n1044), .A2(new_n1043), .ZN(new_n1073));
  AOI21_X1  g0873(.A(new_n1072), .B1(new_n1073), .B2(new_n719), .ZN(new_n1074));
  NAND2_X1  g0874(.A1(new_n1051), .A2(new_n1074), .ZN(G378));
  NAND2_X1  g0875(.A1(new_n1029), .A2(new_n1031), .ZN(new_n1076));
  AOI21_X1  g0876(.A(new_n1023), .B1(new_n1073), .B2(new_n1076), .ZN(new_n1077));
  NAND3_X1  g0877(.A1(new_n865), .A2(G330), .A3(new_n871), .ZN(new_n1078));
  INV_X1    g0878(.A(KEYINPUT56), .ZN(new_n1079));
  NOR2_X1   g0879(.A1(new_n366), .A2(new_n833), .ZN(new_n1080));
  INV_X1    g0880(.A(new_n376), .ZN(new_n1081));
  OAI21_X1  g0881(.A(new_n1080), .B1(new_n629), .B2(new_n1081), .ZN(new_n1082));
  INV_X1    g0882(.A(KEYINPUT55), .ZN(new_n1083));
  INV_X1    g0883(.A(new_n1080), .ZN(new_n1084));
  NAND4_X1  g0884(.A1(new_n627), .A2(new_n376), .A3(new_n628), .A4(new_n1084), .ZN(new_n1085));
  NAND3_X1  g0885(.A1(new_n1082), .A2(new_n1083), .A3(new_n1085), .ZN(new_n1086));
  INV_X1    g0886(.A(new_n1086), .ZN(new_n1087));
  AOI21_X1  g0887(.A(new_n1083), .B1(new_n1082), .B2(new_n1085), .ZN(new_n1088));
  OAI21_X1  g0888(.A(new_n1079), .B1(new_n1087), .B2(new_n1088), .ZN(new_n1089));
  NAND2_X1  g0889(.A1(new_n1082), .A2(new_n1085), .ZN(new_n1090));
  NAND2_X1  g0890(.A1(new_n1090), .A2(KEYINPUT55), .ZN(new_n1091));
  NAND3_X1  g0891(.A1(new_n1091), .A2(KEYINPUT56), .A3(new_n1086), .ZN(new_n1092));
  NAND2_X1  g0892(.A1(new_n1089), .A2(new_n1092), .ZN(new_n1093));
  NAND2_X1  g0893(.A1(new_n1093), .A2(KEYINPUT122), .ZN(new_n1094));
  NAND2_X1  g0894(.A1(new_n1078), .A2(new_n1094), .ZN(new_n1095));
  AOI22_X1  g0895(.A1(new_n879), .A2(new_n880), .B1(new_n883), .B2(new_n887), .ZN(new_n1096));
  INV_X1    g0896(.A(KEYINPUT122), .ZN(new_n1097));
  NAND3_X1  g0897(.A1(new_n1089), .A2(new_n1092), .A3(new_n1097), .ZN(new_n1098));
  AND3_X1   g0898(.A1(new_n1096), .A2(new_n882), .A3(new_n1098), .ZN(new_n1099));
  AOI21_X1  g0899(.A(new_n1098), .B1(new_n1096), .B2(new_n882), .ZN(new_n1100));
  OAI21_X1  g0900(.A(new_n1095), .B1(new_n1099), .B2(new_n1100), .ZN(new_n1101));
  INV_X1    g0901(.A(new_n1098), .ZN(new_n1102));
  NAND2_X1  g0902(.A1(new_n889), .A2(new_n1102), .ZN(new_n1103));
  NAND3_X1  g0903(.A1(new_n1096), .A2(new_n882), .A3(new_n1098), .ZN(new_n1104));
  NAND4_X1  g0904(.A1(new_n1103), .A2(new_n1104), .A3(new_n1078), .A4(new_n1094), .ZN(new_n1105));
  NAND2_X1  g0905(.A1(new_n1101), .A2(new_n1105), .ZN(new_n1106));
  INV_X1    g0906(.A(KEYINPUT57), .ZN(new_n1107));
  NOR3_X1   g0907(.A1(new_n1077), .A2(new_n1106), .A3(new_n1107), .ZN(new_n1108));
  OAI21_X1  g0908(.A(KEYINPUT123), .B1(new_n1108), .B2(new_n678), .ZN(new_n1109));
  OAI21_X1  g0909(.A(new_n1107), .B1(new_n1077), .B2(new_n1106), .ZN(new_n1110));
  INV_X1    g0910(.A(new_n1023), .ZN(new_n1111));
  NAND2_X1  g0911(.A1(new_n1050), .A2(new_n1111), .ZN(new_n1112));
  NAND4_X1  g0912(.A1(new_n1112), .A2(KEYINPUT57), .A3(new_n1105), .A4(new_n1101), .ZN(new_n1113));
  INV_X1    g0913(.A(KEYINPUT123), .ZN(new_n1114));
  NAND3_X1  g0914(.A1(new_n1113), .A2(new_n1114), .A3(new_n677), .ZN(new_n1115));
  NAND3_X1  g0915(.A1(new_n1109), .A2(new_n1110), .A3(new_n1115), .ZN(new_n1116));
  NAND3_X1  g0916(.A1(new_n1101), .A2(new_n1105), .A3(new_n719), .ZN(new_n1117));
  OAI21_X1  g0917(.A(new_n201), .B1(new_n412), .B2(G41), .ZN(new_n1118));
  AOI22_X1  g0918(.A1(new_n753), .A2(G128), .B1(new_n750), .B2(new_n1052), .ZN(new_n1119));
  XNOR2_X1  g0919(.A(new_n1119), .B(KEYINPUT119), .ZN(new_n1120));
  OAI22_X1  g0920(.A1(new_n756), .A2(new_n353), .B1(new_n738), .B2(new_n1058), .ZN(new_n1121));
  AOI21_X1  g0921(.A(new_n1121), .B1(new_n743), .B2(G132), .ZN(new_n1122));
  OAI211_X1 g0922(.A(new_n1120), .B(new_n1122), .C1(new_n799), .C2(new_n734), .ZN(new_n1123));
  XNOR2_X1  g0923(.A(new_n1123), .B(KEYINPUT59), .ZN(new_n1124));
  AOI21_X1  g0924(.A(G41), .B1(new_n746), .B2(G124), .ZN(new_n1125));
  OAI211_X1 g0925(.A(new_n1125), .B(new_n269), .C1(new_n405), .C2(new_n730), .ZN(new_n1126));
  XNOR2_X1  g0926(.A(new_n1126), .B(KEYINPUT120), .ZN(new_n1127));
  OAI21_X1  g0927(.A(new_n1118), .B1(new_n1124), .B2(new_n1127), .ZN(new_n1128));
  OAI22_X1  g0928(.A1(new_n738), .A2(new_n226), .B1(new_n730), .B2(new_n202), .ZN(new_n1129));
  NAND2_X1  g0929(.A1(new_n414), .A2(new_n264), .ZN(new_n1130));
  NOR4_X1   g0930(.A1(new_n1129), .A2(new_n910), .A3(new_n980), .A4(new_n1130), .ZN(new_n1131));
  OAI22_X1  g0931(.A1(new_n752), .A2(new_n378), .B1(new_n745), .B2(new_n767), .ZN(new_n1132));
  AOI21_X1  g0932(.A(new_n1132), .B1(new_n743), .B2(G97), .ZN(new_n1133));
  OAI211_X1 g0933(.A(new_n1131), .B(new_n1133), .C1(new_n550), .C2(new_n734), .ZN(new_n1134));
  XNOR2_X1  g0934(.A(KEYINPUT118), .B(KEYINPUT58), .ZN(new_n1135));
  XOR2_X1   g0935(.A(new_n1134), .B(new_n1135), .Z(new_n1136));
  OAI21_X1  g0936(.A(new_n774), .B1(new_n1128), .B2(new_n1136), .ZN(new_n1137));
  INV_X1    g0937(.A(new_n1137), .ZN(new_n1138));
  OAI22_X1  g0938(.A1(new_n1138), .A2(KEYINPUT121), .B1(G50), .B2(new_n817), .ZN(new_n1139));
  AOI21_X1  g0939(.A(new_n1139), .B1(KEYINPUT121), .B2(new_n1138), .ZN(new_n1140));
  OAI211_X1 g0940(.A(new_n720), .B(new_n1140), .C1(new_n1093), .C2(new_n776), .ZN(new_n1141));
  NAND2_X1  g0941(.A1(new_n1117), .A2(new_n1141), .ZN(new_n1142));
  INV_X1    g0942(.A(new_n1142), .ZN(new_n1143));
  NAND2_X1  g0943(.A1(new_n1116), .A2(new_n1143), .ZN(G375));
  OR2_X1    g0944(.A1(new_n827), .A2(new_n776), .ZN(new_n1145));
  OAI221_X1 g0945(.A(new_n414), .B1(new_n730), .B2(new_n249), .C1(new_n1009), .C2(new_n738), .ZN(new_n1146));
  AOI21_X1  g0946(.A(new_n1146), .B1(new_n386), .B2(new_n806), .ZN(new_n1147));
  NAND2_X1  g0947(.A1(new_n753), .A2(G283), .ZN(new_n1148));
  OAI22_X1  g0948(.A1(new_n734), .A2(new_n378), .B1(new_n745), .B2(new_n458), .ZN(new_n1149));
  AOI21_X1  g0949(.A(new_n1149), .B1(new_n743), .B2(new_n917), .ZN(new_n1150));
  NAND2_X1  g0950(.A1(new_n750), .A2(G97), .ZN(new_n1151));
  NAND4_X1  g0951(.A1(new_n1147), .A2(new_n1148), .A3(new_n1150), .A4(new_n1151), .ZN(new_n1152));
  NOR2_X1   g0952(.A1(new_n738), .A2(new_n804), .ZN(new_n1153));
  OAI21_X1  g0953(.A(new_n256), .B1(new_n730), .B2(new_n202), .ZN(new_n1154));
  AOI211_X1 g0954(.A(new_n1153), .B(new_n1154), .C1(G50), .C2(new_n806), .ZN(new_n1155));
  INV_X1    g0955(.A(G128), .ZN(new_n1156));
  OAI22_X1  g0956(.A1(new_n734), .A2(new_n353), .B1(new_n745), .B2(new_n1156), .ZN(new_n1157));
  AOI21_X1  g0957(.A(new_n1157), .B1(new_n743), .B2(new_n1052), .ZN(new_n1158));
  NAND2_X1  g0958(.A1(new_n753), .A2(G137), .ZN(new_n1159));
  NAND2_X1  g0959(.A1(new_n750), .A2(G159), .ZN(new_n1160));
  NAND4_X1  g0960(.A1(new_n1155), .A2(new_n1158), .A3(new_n1159), .A4(new_n1160), .ZN(new_n1161));
  AND2_X1   g0961(.A1(new_n1152), .A2(new_n1161), .ZN(new_n1162));
  OAI221_X1 g0962(.A(new_n720), .B1(new_n727), .B2(new_n1162), .C1(new_n817), .C2(G68), .ZN(new_n1163));
  XOR2_X1   g0963(.A(new_n1163), .B(KEYINPUT124), .Z(new_n1164));
  AOI22_X1  g0964(.A1(new_n1076), .A2(new_n719), .B1(new_n1145), .B2(new_n1164), .ZN(new_n1165));
  NAND3_X1  g0965(.A1(new_n1029), .A2(new_n1023), .A3(new_n1031), .ZN(new_n1166));
  NAND2_X1  g0966(.A1(new_n1166), .A2(new_n950), .ZN(new_n1167));
  OAI21_X1  g0967(.A(new_n1165), .B1(new_n1167), .B2(new_n1032), .ZN(G381));
  INV_X1    g0968(.A(G396), .ZN(new_n1169));
  NAND4_X1  g0969(.A1(new_n966), .A2(new_n1169), .A3(new_n968), .A4(new_n995), .ZN(new_n1170));
  NOR2_X1   g0970(.A1(G390), .A2(new_n1170), .ZN(new_n1171));
  NOR2_X1   g0971(.A1(G381), .A2(G384), .ZN(new_n1172));
  NAND3_X1  g0972(.A1(new_n963), .A2(new_n1171), .A3(new_n1172), .ZN(new_n1173));
  OR2_X1    g0973(.A1(new_n1173), .A2(KEYINPUT125), .ZN(new_n1174));
  NAND2_X1  g0974(.A1(new_n1173), .A2(KEYINPUT125), .ZN(new_n1175));
  AND3_X1   g0975(.A1(new_n1113), .A2(new_n1114), .A3(new_n677), .ZN(new_n1176));
  AOI21_X1  g0976(.A(new_n1114), .B1(new_n1113), .B2(new_n677), .ZN(new_n1177));
  INV_X1    g0977(.A(new_n1110), .ZN(new_n1178));
  NOR3_X1   g0978(.A1(new_n1176), .A2(new_n1177), .A3(new_n1178), .ZN(new_n1179));
  NAND3_X1  g0979(.A1(new_n1143), .A2(new_n1074), .A3(new_n1051), .ZN(new_n1180));
  NOR2_X1   g0980(.A1(new_n1179), .A2(new_n1180), .ZN(new_n1181));
  NAND3_X1  g0981(.A1(new_n1174), .A2(new_n1175), .A3(new_n1181), .ZN(G407));
  INV_X1    g0982(.A(G213), .ZN(new_n1183));
  INV_X1    g0983(.A(G343), .ZN(new_n1184));
  AOI21_X1  g0984(.A(new_n1183), .B1(new_n1181), .B2(new_n1184), .ZN(new_n1185));
  NAND2_X1  g0985(.A1(G407), .A2(new_n1185), .ZN(G409));
  AND4_X1   g0986(.A1(new_n950), .A2(new_n1112), .A3(new_n1105), .A4(new_n1101), .ZN(new_n1187));
  OAI22_X1  g0987(.A1(new_n1180), .A2(new_n1187), .B1(new_n1183), .B2(G343), .ZN(new_n1188));
  AOI21_X1  g0988(.A(new_n1188), .B1(G375), .B2(G378), .ZN(new_n1189));
  INV_X1    g0989(.A(KEYINPUT60), .ZN(new_n1190));
  AOI21_X1  g0990(.A(new_n678), .B1(new_n1166), .B2(new_n1190), .ZN(new_n1191));
  OAI211_X1 g0991(.A(new_n1191), .B(new_n1033), .C1(new_n1190), .C2(new_n1166), .ZN(new_n1192));
  NAND2_X1  g0992(.A1(new_n1192), .A2(new_n1165), .ZN(new_n1193));
  XNOR2_X1  g0993(.A(G384), .B(KEYINPUT126), .ZN(new_n1194));
  NAND2_X1  g0994(.A1(new_n1193), .A2(new_n1194), .ZN(new_n1195));
  NAND3_X1  g0995(.A1(new_n797), .A2(KEYINPUT126), .A3(new_n820), .ZN(new_n1196));
  INV_X1    g0996(.A(new_n1196), .ZN(new_n1197));
  NAND3_X1  g0997(.A1(new_n1192), .A2(new_n1165), .A3(new_n1197), .ZN(new_n1198));
  NAND2_X1  g0998(.A1(new_n1195), .A2(new_n1198), .ZN(new_n1199));
  NAND2_X1  g0999(.A1(new_n1189), .A2(new_n1199), .ZN(new_n1200));
  NAND3_X1  g1000(.A1(new_n1184), .A2(G213), .A3(G2897), .ZN(new_n1201));
  XNOR2_X1  g1001(.A(new_n1199), .B(new_n1201), .ZN(new_n1202));
  OAI21_X1  g1002(.A(G378), .B1(new_n1179), .B2(new_n1142), .ZN(new_n1203));
  INV_X1    g1003(.A(new_n1188), .ZN(new_n1204));
  AOI21_X1  g1004(.A(new_n1202), .B1(new_n1203), .B2(new_n1204), .ZN(new_n1205));
  INV_X1    g1005(.A(KEYINPUT63), .ZN(new_n1206));
  OAI21_X1  g1006(.A(new_n1200), .B1(new_n1205), .B2(new_n1206), .ZN(new_n1207));
  NAND2_X1  g1007(.A1(G393), .A2(G396), .ZN(new_n1208));
  NAND2_X1  g1008(.A1(new_n1208), .A2(new_n1170), .ZN(new_n1209));
  NAND2_X1  g1009(.A1(new_n1209), .A2(G390), .ZN(new_n1210));
  AOI21_X1  g1010(.A(KEYINPUT109), .B1(new_n1208), .B2(new_n1170), .ZN(new_n1211));
  OAI21_X1  g1011(.A(new_n1210), .B1(G390), .B2(new_n1211), .ZN(new_n1212));
  OR2_X1    g1012(.A1(new_n951), .A2(new_n961), .ZN(new_n1213));
  NAND3_X1  g1013(.A1(new_n1212), .A2(new_n931), .A3(new_n1213), .ZN(new_n1214));
  OAI211_X1 g1014(.A(new_n1210), .B(new_n962), .C1(G390), .C2(new_n1211), .ZN(new_n1215));
  NAND2_X1  g1015(.A1(new_n1214), .A2(new_n1215), .ZN(new_n1216));
  INV_X1    g1016(.A(G378), .ZN(new_n1217));
  AOI21_X1  g1017(.A(new_n1217), .B1(new_n1116), .B2(new_n1143), .ZN(new_n1218));
  INV_X1    g1018(.A(new_n1199), .ZN(new_n1219));
  NOR3_X1   g1019(.A1(new_n1218), .A2(new_n1188), .A3(new_n1219), .ZN(new_n1220));
  AOI21_X1  g1020(.A(new_n1216), .B1(new_n1220), .B2(KEYINPUT63), .ZN(new_n1221));
  INV_X1    g1021(.A(KEYINPUT61), .ZN(new_n1222));
  NAND3_X1  g1022(.A1(new_n1207), .A2(new_n1221), .A3(new_n1222), .ZN(new_n1223));
  OAI21_X1  g1023(.A(new_n1222), .B1(new_n1189), .B2(new_n1202), .ZN(new_n1224));
  INV_X1    g1024(.A(KEYINPUT62), .ZN(new_n1225));
  AOI21_X1  g1025(.A(new_n1225), .B1(new_n1189), .B2(new_n1199), .ZN(new_n1226));
  NOR4_X1   g1026(.A1(new_n1218), .A2(KEYINPUT62), .A3(new_n1188), .A4(new_n1219), .ZN(new_n1227));
  NOR3_X1   g1027(.A1(new_n1224), .A2(new_n1226), .A3(new_n1227), .ZN(new_n1228));
  INV_X1    g1028(.A(new_n1216), .ZN(new_n1229));
  OAI21_X1  g1029(.A(new_n1223), .B1(new_n1228), .B2(new_n1229), .ZN(G405));
  OAI211_X1 g1030(.A(new_n1203), .B(new_n1199), .C1(new_n1179), .C2(new_n1180), .ZN(new_n1231));
  OAI21_X1  g1031(.A(new_n1219), .B1(new_n1181), .B2(new_n1218), .ZN(new_n1232));
  NAND2_X1  g1032(.A1(new_n1231), .A2(new_n1232), .ZN(new_n1233));
  XNOR2_X1  g1033(.A(new_n1233), .B(new_n1216), .ZN(G402));
endmodule


