//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 1 0 0 0 0 1 1 1 0 0 0 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 1 1 1 1 0 0 1 1 1 1 1 0 0 0 0 0 0 0 0 0 1 1 0 1 1 1 0 1 0 1 0 0 1 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:24:50 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n698, new_n699,
    new_n700, new_n701, new_n702, new_n703, new_n705, new_n706, new_n707,
    new_n708, new_n709, new_n710, new_n711, new_n712, new_n713, new_n714,
    new_n715, new_n717, new_n718, new_n719, new_n720, new_n721, new_n722,
    new_n723, new_n724, new_n725, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n744, new_n745,
    new_n746, new_n747, new_n748, new_n749, new_n750, new_n751, new_n752,
    new_n753, new_n754, new_n755, new_n756, new_n757, new_n758, new_n759,
    new_n760, new_n761, new_n762, new_n763, new_n764, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n781, new_n782,
    new_n784, new_n785, new_n786, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n798, new_n799,
    new_n800, new_n801, new_n802, new_n803, new_n804, new_n805, new_n806,
    new_n807, new_n808, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n820, new_n821, new_n822,
    new_n823, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n938,
    new_n939, new_n940, new_n941, new_n942, new_n943, new_n944, new_n945,
    new_n946, new_n947, new_n948, new_n949, new_n950, new_n951, new_n952,
    new_n953, new_n954, new_n955, new_n956, new_n957, new_n958, new_n959,
    new_n960, new_n961, new_n962, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n972, new_n973, new_n974, new_n975,
    new_n977, new_n978, new_n979, new_n980, new_n981, new_n982, new_n983,
    new_n985, new_n986, new_n987, new_n988, new_n989, new_n990, new_n991,
    new_n992, new_n993, new_n994, new_n995, new_n996, new_n997, new_n998,
    new_n999, new_n1000, new_n1001, new_n1003, new_n1004, new_n1005,
    new_n1006, new_n1007, new_n1008, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1017, new_n1018,
    new_n1019, new_n1020, new_n1021, new_n1022, new_n1023, new_n1024,
    new_n1025, new_n1026, new_n1027, new_n1028, new_n1029, new_n1030,
    new_n1031, new_n1032, new_n1033, new_n1034, new_n1035, new_n1036,
    new_n1037, new_n1038, new_n1039, new_n1040, new_n1041, new_n1042,
    new_n1044, new_n1045, new_n1046, new_n1047, new_n1048, new_n1049,
    new_n1050, new_n1051, new_n1052;
  INV_X1    g000(.A(G221), .ZN(new_n187));
  XOR2_X1   g001(.A(KEYINPUT9), .B(G234), .Z(new_n188));
  XNOR2_X1  g002(.A(new_n188), .B(KEYINPUT78), .ZN(new_n189));
  INV_X1    g003(.A(G902), .ZN(new_n190));
  AOI21_X1  g004(.A(new_n187), .B1(new_n189), .B2(new_n190), .ZN(new_n191));
  INV_X1    g005(.A(G137), .ZN(new_n192));
  OAI21_X1  g006(.A(KEYINPUT11), .B1(new_n192), .B2(G134), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n192), .A2(G134), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n193), .A2(new_n194), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n192), .A2(KEYINPUT64), .ZN(new_n196));
  INV_X1    g010(.A(KEYINPUT64), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n197), .A2(G137), .ZN(new_n198));
  AND2_X1   g012(.A1(KEYINPUT11), .A2(G134), .ZN(new_n199));
  NAND3_X1  g013(.A1(new_n196), .A2(new_n198), .A3(new_n199), .ZN(new_n200));
  INV_X1    g014(.A(G131), .ZN(new_n201));
  AND3_X1   g015(.A1(new_n195), .A2(new_n200), .A3(new_n201), .ZN(new_n202));
  AOI21_X1  g016(.A(new_n201), .B1(new_n195), .B2(new_n200), .ZN(new_n203));
  NOR2_X1   g017(.A1(new_n202), .A2(new_n203), .ZN(new_n204));
  INV_X1    g018(.A(new_n204), .ZN(new_n205));
  INV_X1    g019(.A(G104), .ZN(new_n206));
  AND2_X1   g020(.A1(KEYINPUT80), .A2(G107), .ZN(new_n207));
  NOR2_X1   g021(.A1(KEYINPUT80), .A2(G107), .ZN(new_n208));
  OAI21_X1  g022(.A(new_n206), .B1(new_n207), .B2(new_n208), .ZN(new_n209));
  INV_X1    g023(.A(G107), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n210), .A2(G104), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n209), .A2(new_n211), .ZN(new_n212));
  AND2_X1   g026(.A1(new_n212), .A2(G101), .ZN(new_n213));
  INV_X1    g027(.A(G128), .ZN(new_n214));
  INV_X1    g028(.A(G143), .ZN(new_n215));
  NOR2_X1   g029(.A1(new_n215), .A2(G146), .ZN(new_n216));
  INV_X1    g030(.A(G146), .ZN(new_n217));
  NOR2_X1   g031(.A1(new_n217), .A2(G143), .ZN(new_n218));
  OAI21_X1  g032(.A(new_n214), .B1(new_n216), .B2(new_n218), .ZN(new_n219));
  NOR2_X1   g033(.A1(new_n214), .A2(KEYINPUT1), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n217), .A2(G143), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n215), .A2(G146), .ZN(new_n222));
  NAND4_X1  g036(.A1(new_n220), .A2(new_n221), .A3(new_n222), .A4(KEYINPUT66), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n218), .A2(KEYINPUT1), .ZN(new_n224));
  AND3_X1   g038(.A1(new_n219), .A2(new_n223), .A3(new_n224), .ZN(new_n225));
  XNOR2_X1  g039(.A(G143), .B(G146), .ZN(new_n226));
  AOI21_X1  g040(.A(KEYINPUT66), .B1(new_n226), .B2(new_n220), .ZN(new_n227));
  INV_X1    g041(.A(new_n227), .ZN(new_n228));
  INV_X1    g042(.A(new_n208), .ZN(new_n229));
  NOR2_X1   g043(.A1(new_n206), .A2(KEYINPUT3), .ZN(new_n230));
  NAND2_X1  g044(.A1(KEYINPUT80), .A2(G107), .ZN(new_n231));
  NAND3_X1  g045(.A1(new_n229), .A2(new_n230), .A3(new_n231), .ZN(new_n232));
  NOR2_X1   g046(.A1(new_n210), .A2(G104), .ZN(new_n233));
  NOR2_X1   g047(.A1(new_n233), .A2(G101), .ZN(new_n234));
  OAI211_X1 g048(.A(KEYINPUT79), .B(KEYINPUT3), .C1(new_n206), .C2(G107), .ZN(new_n235));
  INV_X1    g049(.A(new_n235), .ZN(new_n236));
  AOI21_X1  g050(.A(KEYINPUT79), .B1(new_n211), .B2(KEYINPUT3), .ZN(new_n237));
  OAI211_X1 g051(.A(new_n232), .B(new_n234), .C1(new_n236), .C2(new_n237), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n238), .A2(KEYINPUT81), .ZN(new_n239));
  OAI21_X1  g053(.A(KEYINPUT3), .B1(new_n206), .B2(G107), .ZN(new_n240));
  INV_X1    g054(.A(KEYINPUT79), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n240), .A2(new_n241), .ZN(new_n242));
  NOR2_X1   g056(.A1(new_n207), .A2(new_n208), .ZN(new_n243));
  AOI22_X1  g057(.A1(new_n242), .A2(new_n235), .B1(new_n243), .B2(new_n230), .ZN(new_n244));
  INV_X1    g058(.A(KEYINPUT81), .ZN(new_n245));
  NAND3_X1  g059(.A1(new_n244), .A2(new_n245), .A3(new_n234), .ZN(new_n246));
  AOI221_X4 g060(.A(new_n213), .B1(new_n225), .B2(new_n228), .C1(new_n239), .C2(new_n246), .ZN(new_n247));
  NAND3_X1  g061(.A1(new_n219), .A2(new_n223), .A3(new_n224), .ZN(new_n248));
  NOR2_X1   g062(.A1(new_n248), .A2(new_n227), .ZN(new_n249));
  INV_X1    g063(.A(new_n249), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n239), .A2(new_n246), .ZN(new_n251));
  INV_X1    g065(.A(new_n213), .ZN(new_n252));
  AOI21_X1  g066(.A(new_n250), .B1(new_n251), .B2(new_n252), .ZN(new_n253));
  OAI211_X1 g067(.A(KEYINPUT12), .B(new_n205), .C1(new_n247), .C2(new_n253), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n254), .A2(KEYINPUT82), .ZN(new_n255));
  NOR2_X1   g069(.A1(new_n238), .A2(KEYINPUT81), .ZN(new_n256));
  AOI21_X1  g070(.A(new_n245), .B1(new_n244), .B2(new_n234), .ZN(new_n257));
  OAI21_X1  g071(.A(new_n252), .B1(new_n256), .B2(new_n257), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n258), .A2(new_n249), .ZN(new_n259));
  NAND3_X1  g073(.A1(new_n251), .A2(new_n250), .A3(new_n252), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n259), .A2(new_n260), .ZN(new_n261));
  INV_X1    g075(.A(KEYINPUT82), .ZN(new_n262));
  NAND4_X1  g076(.A1(new_n261), .A2(new_n262), .A3(KEYINPUT12), .A4(new_n205), .ZN(new_n263));
  OAI21_X1  g077(.A(new_n205), .B1(new_n247), .B2(new_n253), .ZN(new_n264));
  INV_X1    g078(.A(KEYINPUT12), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n264), .A2(new_n265), .ZN(new_n266));
  NAND3_X1  g080(.A1(new_n255), .A2(new_n263), .A3(new_n266), .ZN(new_n267));
  INV_X1    g081(.A(KEYINPUT84), .ZN(new_n268));
  AND2_X1   g082(.A1(new_n267), .A2(new_n268), .ZN(new_n269));
  NAND2_X1  g083(.A1(KEYINPUT0), .A2(G128), .ZN(new_n270));
  NAND2_X1  g084(.A1(new_n226), .A2(new_n270), .ZN(new_n271));
  XOR2_X1   g085(.A(KEYINPUT0), .B(G128), .Z(new_n272));
  OAI21_X1  g086(.A(new_n271), .B1(new_n272), .B2(new_n226), .ZN(new_n273));
  INV_X1    g087(.A(KEYINPUT4), .ZN(new_n274));
  OAI21_X1  g088(.A(new_n232), .B1(new_n236), .B2(new_n237), .ZN(new_n275));
  OAI21_X1  g089(.A(G101), .B1(new_n275), .B2(new_n233), .ZN(new_n276));
  AOI21_X1  g090(.A(new_n274), .B1(new_n251), .B2(new_n276), .ZN(new_n277));
  OAI21_X1  g091(.A(new_n244), .B1(G104), .B2(new_n210), .ZN(new_n278));
  AOI21_X1  g092(.A(KEYINPUT4), .B1(new_n278), .B2(G101), .ZN(new_n279));
  OAI21_X1  g093(.A(new_n273), .B1(new_n277), .B2(new_n279), .ZN(new_n280));
  AOI21_X1  g094(.A(new_n213), .B1(new_n239), .B2(new_n246), .ZN(new_n281));
  NAND3_X1  g095(.A1(new_n281), .A2(KEYINPUT10), .A3(new_n250), .ZN(new_n282));
  INV_X1    g096(.A(KEYINPUT10), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n260), .A2(new_n283), .ZN(new_n284));
  NAND4_X1  g098(.A1(new_n280), .A2(new_n204), .A3(new_n282), .A4(new_n284), .ZN(new_n285));
  XNOR2_X1  g099(.A(G110), .B(G140), .ZN(new_n286));
  INV_X1    g100(.A(G227), .ZN(new_n287));
  NOR2_X1   g101(.A1(new_n287), .A2(G953), .ZN(new_n288));
  XNOR2_X1  g102(.A(new_n286), .B(new_n288), .ZN(new_n289));
  INV_X1    g103(.A(new_n289), .ZN(new_n290));
  AND2_X1   g104(.A1(new_n285), .A2(new_n290), .ZN(new_n291));
  NAND4_X1  g105(.A1(new_n255), .A2(new_n263), .A3(new_n266), .A4(KEYINPUT84), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n291), .A2(new_n292), .ZN(new_n293));
  INV_X1    g107(.A(new_n285), .ZN(new_n294));
  OAI21_X1  g108(.A(new_n276), .B1(new_n256), .B2(new_n257), .ZN(new_n295));
  AOI21_X1  g109(.A(new_n279), .B1(new_n295), .B2(KEYINPUT4), .ZN(new_n296));
  INV_X1    g110(.A(new_n273), .ZN(new_n297));
  OAI211_X1 g111(.A(new_n282), .B(new_n284), .C1(new_n296), .C2(new_n297), .ZN(new_n298));
  INV_X1    g112(.A(KEYINPUT83), .ZN(new_n299));
  AOI21_X1  g113(.A(new_n204), .B1(new_n298), .B2(new_n299), .ZN(new_n300));
  NAND4_X1  g114(.A1(new_n280), .A2(KEYINPUT83), .A3(new_n282), .A4(new_n284), .ZN(new_n301));
  AOI21_X1  g115(.A(new_n294), .B1(new_n300), .B2(new_n301), .ZN(new_n302));
  OAI22_X1  g116(.A1(new_n269), .A2(new_n293), .B1(new_n302), .B2(new_n290), .ZN(new_n303));
  INV_X1    g117(.A(G469), .ZN(new_n304));
  NAND3_X1  g118(.A1(new_n303), .A2(new_n304), .A3(new_n190), .ZN(new_n305));
  INV_X1    g119(.A(KEYINPUT85), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n305), .A2(new_n306), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n295), .A2(KEYINPUT4), .ZN(new_n308));
  INV_X1    g122(.A(new_n279), .ZN(new_n309));
  AOI21_X1  g123(.A(new_n297), .B1(new_n308), .B2(new_n309), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n284), .A2(new_n282), .ZN(new_n311));
  OAI21_X1  g125(.A(new_n299), .B1(new_n310), .B2(new_n311), .ZN(new_n312));
  NAND3_X1  g126(.A1(new_n312), .A2(new_n205), .A3(new_n301), .ZN(new_n313));
  NAND2_X1  g127(.A1(new_n313), .A2(new_n285), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n314), .A2(new_n289), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n267), .A2(new_n268), .ZN(new_n316));
  NAND3_X1  g130(.A1(new_n316), .A2(new_n291), .A3(new_n292), .ZN(new_n317));
  AOI21_X1  g131(.A(G902), .B1(new_n315), .B2(new_n317), .ZN(new_n318));
  NAND3_X1  g132(.A1(new_n318), .A2(KEYINPUT85), .A3(new_n304), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n307), .A2(new_n319), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n267), .A2(new_n285), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n321), .A2(new_n289), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n313), .A2(new_n291), .ZN(new_n323));
  NAND2_X1  g137(.A1(new_n322), .A2(new_n323), .ZN(new_n324));
  AOI21_X1  g138(.A(new_n304), .B1(new_n324), .B2(new_n190), .ZN(new_n325));
  INV_X1    g139(.A(new_n325), .ZN(new_n326));
  AOI21_X1  g140(.A(new_n191), .B1(new_n320), .B2(new_n326), .ZN(new_n327));
  OAI21_X1  g141(.A(G210), .B1(G237), .B2(G902), .ZN(new_n328));
  INV_X1    g142(.A(new_n328), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n273), .A2(G125), .ZN(new_n330));
  OAI21_X1  g144(.A(new_n330), .B1(new_n249), .B2(G125), .ZN(new_n331));
  INV_X1    g145(.A(G224), .ZN(new_n332));
  NOR2_X1   g146(.A1(new_n332), .A2(G953), .ZN(new_n333));
  XNOR2_X1  g147(.A(new_n331), .B(new_n333), .ZN(new_n334));
  AND3_X1   g148(.A1(KEYINPUT67), .A2(KEYINPUT2), .A3(G113), .ZN(new_n335));
  AOI21_X1  g149(.A(KEYINPUT67), .B1(KEYINPUT2), .B2(G113), .ZN(new_n336));
  OAI22_X1  g150(.A1(new_n335), .A2(new_n336), .B1(KEYINPUT2), .B2(G113), .ZN(new_n337));
  XNOR2_X1  g151(.A(G116), .B(G119), .ZN(new_n338));
  XNOR2_X1  g152(.A(new_n337), .B(new_n338), .ZN(new_n339));
  INV_X1    g153(.A(new_n339), .ZN(new_n340));
  OAI21_X1  g154(.A(new_n340), .B1(new_n277), .B2(new_n279), .ZN(new_n341));
  INV_X1    g155(.A(new_n338), .ZN(new_n342));
  NOR2_X1   g156(.A1(new_n337), .A2(new_n342), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n338), .A2(KEYINPUT5), .ZN(new_n344));
  INV_X1    g158(.A(G116), .ZN(new_n345));
  NOR3_X1   g159(.A1(new_n345), .A2(KEYINPUT5), .A3(G119), .ZN(new_n346));
  INV_X1    g160(.A(G113), .ZN(new_n347));
  NOR2_X1   g161(.A1(new_n346), .A2(new_n347), .ZN(new_n348));
  AOI21_X1  g162(.A(new_n343), .B1(new_n344), .B2(new_n348), .ZN(new_n349));
  NAND3_X1  g163(.A1(new_n281), .A2(KEYINPUT86), .A3(new_n349), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n281), .A2(new_n349), .ZN(new_n351));
  INV_X1    g165(.A(KEYINPUT86), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n351), .A2(new_n352), .ZN(new_n353));
  XNOR2_X1  g167(.A(G110), .B(G122), .ZN(new_n354));
  NAND4_X1  g168(.A1(new_n341), .A2(new_n350), .A3(new_n353), .A4(new_n354), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n355), .A2(KEYINPUT6), .ZN(new_n356));
  NAND3_X1  g170(.A1(new_n341), .A2(new_n350), .A3(new_n353), .ZN(new_n357));
  XOR2_X1   g171(.A(new_n354), .B(KEYINPUT87), .Z(new_n358));
  NAND2_X1  g172(.A1(new_n357), .A2(new_n358), .ZN(new_n359));
  NAND2_X1  g173(.A1(new_n356), .A2(new_n359), .ZN(new_n360));
  NAND3_X1  g174(.A1(new_n357), .A2(KEYINPUT6), .A3(new_n358), .ZN(new_n361));
  AOI21_X1  g175(.A(new_n334), .B1(new_n360), .B2(new_n361), .ZN(new_n362));
  OAI21_X1  g176(.A(KEYINPUT7), .B1(new_n332), .B2(G953), .ZN(new_n363));
  XOR2_X1   g177(.A(new_n331), .B(new_n363), .Z(new_n364));
  XNOR2_X1  g178(.A(new_n281), .B(new_n349), .ZN(new_n365));
  XNOR2_X1  g179(.A(new_n354), .B(KEYINPUT8), .ZN(new_n366));
  AOI21_X1  g180(.A(new_n364), .B1(new_n365), .B2(new_n366), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n367), .A2(new_n355), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n368), .A2(new_n190), .ZN(new_n369));
  OAI21_X1  g183(.A(new_n329), .B1(new_n362), .B2(new_n369), .ZN(new_n370));
  INV_X1    g184(.A(KEYINPUT88), .ZN(new_n371));
  INV_X1    g185(.A(new_n334), .ZN(new_n372));
  AOI22_X1  g186(.A1(new_n355), .A2(KEYINPUT6), .B1(new_n357), .B2(new_n358), .ZN(new_n373));
  AND3_X1   g187(.A1(new_n357), .A2(KEYINPUT6), .A3(new_n358), .ZN(new_n374));
  OAI21_X1  g188(.A(new_n372), .B1(new_n373), .B2(new_n374), .ZN(new_n375));
  AOI21_X1  g189(.A(G902), .B1(new_n367), .B2(new_n355), .ZN(new_n376));
  NAND3_X1  g190(.A1(new_n375), .A2(new_n328), .A3(new_n376), .ZN(new_n377));
  NAND3_X1  g191(.A1(new_n370), .A2(new_n371), .A3(new_n377), .ZN(new_n378));
  AOI21_X1  g192(.A(new_n328), .B1(new_n375), .B2(new_n376), .ZN(new_n379));
  NAND2_X1  g193(.A1(new_n379), .A2(KEYINPUT88), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n378), .A2(new_n380), .ZN(new_n381));
  OAI21_X1  g195(.A(G214), .B1(G237), .B2(G902), .ZN(new_n382));
  INV_X1    g196(.A(new_n382), .ZN(new_n383));
  INV_X1    g197(.A(KEYINPUT20), .ZN(new_n384));
  XNOR2_X1  g198(.A(G113), .B(G122), .ZN(new_n385));
  XNOR2_X1  g199(.A(new_n385), .B(new_n206), .ZN(new_n386));
  INV_X1    g200(.A(new_n386), .ZN(new_n387));
  INV_X1    g201(.A(G140), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n388), .A2(G125), .ZN(new_n389));
  INV_X1    g203(.A(G125), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n390), .A2(G140), .ZN(new_n391));
  NAND3_X1  g205(.A1(new_n389), .A2(new_n391), .A3(KEYINPUT16), .ZN(new_n392));
  NOR2_X1   g206(.A1(new_n390), .A2(G140), .ZN(new_n393));
  INV_X1    g207(.A(KEYINPUT16), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n393), .A2(new_n394), .ZN(new_n395));
  NAND3_X1  g209(.A1(new_n392), .A2(new_n395), .A3(G146), .ZN(new_n396));
  INV_X1    g210(.A(G237), .ZN(new_n397));
  INV_X1    g211(.A(G953), .ZN(new_n398));
  NAND3_X1  g212(.A1(new_n397), .A2(new_n398), .A3(G214), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n399), .A2(new_n215), .ZN(new_n400));
  NOR2_X1   g214(.A1(G237), .A2(G953), .ZN(new_n401));
  NAND3_X1  g215(.A1(new_n401), .A2(G143), .A3(G214), .ZN(new_n402));
  NAND3_X1  g216(.A1(new_n400), .A2(new_n201), .A3(new_n402), .ZN(new_n403));
  INV_X1    g217(.A(new_n403), .ZN(new_n404));
  AOI21_X1  g218(.A(new_n201), .B1(new_n400), .B2(new_n402), .ZN(new_n405));
  OAI21_X1  g219(.A(new_n396), .B1(new_n404), .B2(new_n405), .ZN(new_n406));
  INV_X1    g220(.A(KEYINPUT89), .ZN(new_n407));
  NOR2_X1   g221(.A1(new_n388), .A2(G125), .ZN(new_n408));
  OAI21_X1  g222(.A(new_n407), .B1(new_n393), .B2(new_n408), .ZN(new_n409));
  NAND3_X1  g223(.A1(new_n389), .A2(new_n391), .A3(KEYINPUT89), .ZN(new_n410));
  NAND3_X1  g224(.A1(new_n409), .A2(KEYINPUT19), .A3(new_n410), .ZN(new_n411));
  XNOR2_X1  g225(.A(G125), .B(G140), .ZN(new_n412));
  INV_X1    g226(.A(KEYINPUT19), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n412), .A2(new_n413), .ZN(new_n414));
  NAND3_X1  g228(.A1(new_n411), .A2(new_n217), .A3(new_n414), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n415), .A2(KEYINPUT90), .ZN(new_n416));
  INV_X1    g230(.A(KEYINPUT90), .ZN(new_n417));
  NAND4_X1  g231(.A1(new_n411), .A2(new_n417), .A3(new_n217), .A4(new_n414), .ZN(new_n418));
  AOI21_X1  g232(.A(new_n406), .B1(new_n416), .B2(new_n418), .ZN(new_n419));
  NAND3_X1  g233(.A1(new_n409), .A2(G146), .A3(new_n410), .ZN(new_n420));
  NOR3_X1   g234(.A1(new_n393), .A2(new_n408), .A3(G146), .ZN(new_n421));
  INV_X1    g235(.A(new_n421), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n420), .A2(new_n422), .ZN(new_n423));
  NAND2_X1  g237(.A1(KEYINPUT18), .A2(G131), .ZN(new_n424));
  NAND3_X1  g238(.A1(new_n400), .A2(new_n402), .A3(new_n424), .ZN(new_n425));
  NAND2_X1  g239(.A1(new_n400), .A2(new_n402), .ZN(new_n426));
  NAND3_X1  g240(.A1(new_n426), .A2(KEYINPUT18), .A3(G131), .ZN(new_n427));
  NAND3_X1  g241(.A1(new_n423), .A2(new_n425), .A3(new_n427), .ZN(new_n428));
  INV_X1    g242(.A(new_n428), .ZN(new_n429));
  OAI21_X1  g243(.A(new_n387), .B1(new_n419), .B2(new_n429), .ZN(new_n430));
  INV_X1    g244(.A(new_n396), .ZN(new_n431));
  AOI21_X1  g245(.A(G146), .B1(new_n392), .B2(new_n395), .ZN(new_n432));
  NOR2_X1   g246(.A1(new_n431), .A2(new_n432), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n426), .A2(G131), .ZN(new_n434));
  INV_X1    g248(.A(KEYINPUT17), .ZN(new_n435));
  NAND3_X1  g249(.A1(new_n434), .A2(new_n435), .A3(new_n403), .ZN(new_n436));
  AND3_X1   g250(.A1(new_n405), .A2(KEYINPUT91), .A3(KEYINPUT17), .ZN(new_n437));
  AOI21_X1  g251(.A(KEYINPUT91), .B1(new_n405), .B2(KEYINPUT17), .ZN(new_n438));
  OAI211_X1 g252(.A(new_n433), .B(new_n436), .C1(new_n437), .C2(new_n438), .ZN(new_n439));
  NAND3_X1  g253(.A1(new_n439), .A2(new_n386), .A3(new_n428), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n430), .A2(new_n440), .ZN(new_n441));
  NOR2_X1   g255(.A1(G475), .A2(G902), .ZN(new_n442));
  AOI21_X1  g256(.A(new_n384), .B1(new_n441), .B2(new_n442), .ZN(new_n443));
  INV_X1    g257(.A(new_n442), .ZN(new_n444));
  AOI211_X1 g258(.A(KEYINPUT20), .B(new_n444), .C1(new_n430), .C2(new_n440), .ZN(new_n445));
  NOR2_X1   g259(.A1(new_n443), .A2(new_n445), .ZN(new_n446));
  INV_X1    g260(.A(G475), .ZN(new_n447));
  AND3_X1   g261(.A1(new_n439), .A2(new_n386), .A3(new_n428), .ZN(new_n448));
  AOI21_X1  g262(.A(new_n386), .B1(new_n439), .B2(new_n428), .ZN(new_n449));
  OR3_X1    g263(.A1(new_n448), .A2(new_n449), .A3(KEYINPUT92), .ZN(new_n450));
  AOI21_X1  g264(.A(G902), .B1(new_n449), .B2(KEYINPUT92), .ZN(new_n451));
  AOI21_X1  g265(.A(new_n447), .B1(new_n450), .B2(new_n451), .ZN(new_n452));
  NOR2_X1   g266(.A1(new_n446), .A2(new_n452), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n215), .A2(G128), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n214), .A2(G143), .ZN(new_n455));
  INV_X1    g269(.A(G134), .ZN(new_n456));
  NAND3_X1  g270(.A1(new_n454), .A2(new_n455), .A3(new_n456), .ZN(new_n457));
  XNOR2_X1  g271(.A(new_n457), .B(KEYINPUT96), .ZN(new_n458));
  INV_X1    g272(.A(G122), .ZN(new_n459));
  NOR2_X1   g273(.A1(new_n459), .A2(G116), .ZN(new_n460));
  OAI21_X1  g274(.A(KEYINPUT93), .B1(new_n345), .B2(G122), .ZN(new_n461));
  INV_X1    g275(.A(KEYINPUT93), .ZN(new_n462));
  NAND3_X1  g276(.A1(new_n462), .A2(new_n459), .A3(G116), .ZN(new_n463));
  AOI21_X1  g277(.A(new_n460), .B1(new_n461), .B2(new_n463), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n464), .A2(new_n243), .ZN(new_n465));
  INV_X1    g279(.A(new_n465), .ZN(new_n466));
  NOR2_X1   g280(.A1(new_n464), .A2(new_n243), .ZN(new_n467));
  OAI21_X1  g281(.A(new_n458), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  NAND4_X1  g282(.A1(new_n215), .A2(KEYINPUT95), .A3(KEYINPUT13), .A4(G128), .ZN(new_n469));
  NAND3_X1  g283(.A1(new_n215), .A2(KEYINPUT13), .A3(G128), .ZN(new_n470));
  INV_X1    g284(.A(new_n470), .ZN(new_n471));
  INV_X1    g285(.A(KEYINPUT95), .ZN(new_n472));
  AOI21_X1  g286(.A(new_n472), .B1(new_n214), .B2(G143), .ZN(new_n473));
  OAI21_X1  g287(.A(new_n469), .B1(new_n471), .B2(new_n473), .ZN(new_n474));
  INV_X1    g288(.A(new_n474), .ZN(new_n475));
  AOI21_X1  g289(.A(KEYINPUT13), .B1(new_n215), .B2(G128), .ZN(new_n476));
  INV_X1    g290(.A(KEYINPUT94), .ZN(new_n477));
  XNOR2_X1  g291(.A(new_n476), .B(new_n477), .ZN(new_n478));
  AOI21_X1  g292(.A(new_n456), .B1(new_n475), .B2(new_n478), .ZN(new_n479));
  INV_X1    g293(.A(KEYINPUT97), .ZN(new_n480));
  INV_X1    g294(.A(KEYINPUT14), .ZN(new_n481));
  OAI21_X1  g295(.A(new_n480), .B1(new_n460), .B2(new_n481), .ZN(new_n482));
  OAI211_X1 g296(.A(KEYINPUT97), .B(KEYINPUT14), .C1(new_n459), .C2(G116), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n482), .A2(new_n483), .ZN(new_n484));
  AOI22_X1  g298(.A1(new_n461), .A2(new_n463), .B1(new_n460), .B2(new_n481), .ZN(new_n485));
  AOI21_X1  g299(.A(new_n210), .B1(new_n484), .B2(new_n485), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n454), .A2(new_n455), .ZN(new_n487));
  NAND2_X1  g301(.A1(new_n487), .A2(G134), .ZN(new_n488));
  NAND2_X1  g302(.A1(new_n488), .A2(new_n457), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n489), .A2(new_n465), .ZN(new_n490));
  OAI22_X1  g304(.A1(new_n468), .A2(new_n479), .B1(new_n486), .B2(new_n490), .ZN(new_n491));
  INV_X1    g305(.A(G217), .ZN(new_n492));
  NOR2_X1   g306(.A1(new_n492), .A2(G953), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n189), .A2(new_n493), .ZN(new_n494));
  NAND2_X1  g308(.A1(new_n491), .A2(new_n494), .ZN(new_n495));
  XNOR2_X1  g309(.A(new_n464), .B(new_n243), .ZN(new_n496));
  XNOR2_X1  g310(.A(new_n476), .B(KEYINPUT94), .ZN(new_n497));
  OAI21_X1  g311(.A(G134), .B1(new_n497), .B2(new_n474), .ZN(new_n498));
  NAND3_X1  g312(.A1(new_n496), .A2(new_n498), .A3(new_n458), .ZN(new_n499));
  NAND2_X1  g313(.A1(new_n484), .A2(new_n485), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n500), .A2(G107), .ZN(new_n501));
  NAND3_X1  g315(.A1(new_n501), .A2(new_n489), .A3(new_n465), .ZN(new_n502));
  INV_X1    g316(.A(new_n494), .ZN(new_n503));
  NAND3_X1  g317(.A1(new_n499), .A2(new_n502), .A3(new_n503), .ZN(new_n504));
  AOI21_X1  g318(.A(G902), .B1(new_n495), .B2(new_n504), .ZN(new_n505));
  INV_X1    g319(.A(G478), .ZN(new_n506));
  NOR2_X1   g320(.A1(new_n506), .A2(KEYINPUT15), .ZN(new_n507));
  XNOR2_X1  g321(.A(new_n505), .B(new_n507), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n453), .A2(new_n508), .ZN(new_n509));
  INV_X1    g323(.A(new_n509), .ZN(new_n510));
  AND2_X1   g324(.A1(new_n398), .A2(G952), .ZN(new_n511));
  INV_X1    g325(.A(G234), .ZN(new_n512));
  OAI21_X1  g326(.A(new_n511), .B1(new_n512), .B2(new_n397), .ZN(new_n513));
  INV_X1    g327(.A(new_n513), .ZN(new_n514));
  AOI211_X1 g328(.A(new_n190), .B(new_n398), .C1(G234), .C2(G237), .ZN(new_n515));
  XNOR2_X1  g329(.A(KEYINPUT21), .B(G898), .ZN(new_n516));
  AOI21_X1  g330(.A(new_n514), .B1(new_n515), .B2(new_n516), .ZN(new_n517));
  INV_X1    g331(.A(new_n517), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n510), .A2(new_n518), .ZN(new_n519));
  NOR3_X1   g333(.A1(new_n381), .A2(new_n383), .A3(new_n519), .ZN(new_n520));
  AND2_X1   g334(.A1(new_n327), .A2(new_n520), .ZN(new_n521));
  AOI21_X1  g335(.A(new_n492), .B1(G234), .B2(new_n190), .ZN(new_n522));
  NOR2_X1   g336(.A1(new_n522), .A2(G902), .ZN(new_n523));
  INV_X1    g337(.A(new_n432), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n524), .A2(new_n396), .ZN(new_n525));
  INV_X1    g339(.A(G119), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n526), .A2(G128), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n214), .A2(G119), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  XNOR2_X1  g343(.A(KEYINPUT24), .B(G110), .ZN(new_n530));
  NOR2_X1   g344(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  INV_X1    g345(.A(KEYINPUT23), .ZN(new_n532));
  OAI21_X1  g346(.A(new_n532), .B1(new_n526), .B2(G128), .ZN(new_n533));
  NAND3_X1  g347(.A1(new_n214), .A2(KEYINPUT23), .A3(G119), .ZN(new_n534));
  NAND3_X1  g348(.A1(new_n533), .A2(new_n527), .A3(new_n534), .ZN(new_n535));
  AOI21_X1  g349(.A(new_n531), .B1(G110), .B2(new_n535), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n525), .A2(new_n536), .ZN(new_n537));
  INV_X1    g351(.A(KEYINPUT72), .ZN(new_n538));
  NOR3_X1   g352(.A1(new_n390), .A2(KEYINPUT16), .A3(G140), .ZN(new_n539));
  AOI21_X1  g353(.A(new_n539), .B1(new_n412), .B2(KEYINPUT16), .ZN(new_n540));
  AOI21_X1  g354(.A(new_n421), .B1(new_n540), .B2(G146), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n529), .A2(new_n530), .ZN(new_n542));
  INV_X1    g356(.A(G110), .ZN(new_n543));
  NAND4_X1  g357(.A1(new_n533), .A2(new_n534), .A3(new_n543), .A4(new_n527), .ZN(new_n544));
  NAND2_X1  g358(.A1(new_n542), .A2(new_n544), .ZN(new_n545));
  AOI21_X1  g359(.A(new_n538), .B1(new_n541), .B2(new_n545), .ZN(new_n546));
  AND4_X1   g360(.A1(new_n538), .A2(new_n545), .A3(new_n396), .A4(new_n422), .ZN(new_n547));
  OAI21_X1  g361(.A(new_n537), .B1(new_n546), .B2(new_n547), .ZN(new_n548));
  INV_X1    g362(.A(KEYINPUT73), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n548), .A2(new_n549), .ZN(new_n550));
  OAI211_X1 g364(.A(KEYINPUT73), .B(new_n537), .C1(new_n546), .C2(new_n547), .ZN(new_n551));
  NOR3_X1   g365(.A1(new_n187), .A2(new_n512), .A3(G953), .ZN(new_n552));
  INV_X1    g366(.A(new_n552), .ZN(new_n553));
  XOR2_X1   g367(.A(KEYINPUT22), .B(G137), .Z(new_n554));
  INV_X1    g368(.A(KEYINPUT74), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  INV_X1    g370(.A(KEYINPUT75), .ZN(new_n557));
  XNOR2_X1  g371(.A(KEYINPUT22), .B(G137), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n558), .A2(KEYINPUT74), .ZN(new_n559));
  NAND3_X1  g373(.A1(new_n556), .A2(new_n557), .A3(new_n559), .ZN(new_n560));
  INV_X1    g374(.A(new_n560), .ZN(new_n561));
  AOI21_X1  g375(.A(new_n557), .B1(new_n556), .B2(new_n559), .ZN(new_n562));
  OAI21_X1  g376(.A(new_n553), .B1(new_n561), .B2(new_n562), .ZN(new_n563));
  INV_X1    g377(.A(new_n562), .ZN(new_n564));
  NAND3_X1  g378(.A1(new_n564), .A2(new_n552), .A3(new_n560), .ZN(new_n565));
  AND2_X1   g379(.A1(new_n563), .A2(new_n565), .ZN(new_n566));
  NAND3_X1  g380(.A1(new_n550), .A2(new_n551), .A3(new_n566), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n541), .A2(new_n545), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n568), .A2(KEYINPUT72), .ZN(new_n569));
  NAND3_X1  g383(.A1(new_n541), .A2(new_n538), .A3(new_n545), .ZN(new_n570));
  AOI22_X1  g384(.A1(new_n569), .A2(new_n570), .B1(new_n525), .B2(new_n536), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n563), .A2(new_n565), .ZN(new_n572));
  AOI21_X1  g386(.A(KEYINPUT76), .B1(new_n571), .B2(new_n572), .ZN(new_n573));
  AND2_X1   g387(.A1(new_n567), .A2(new_n573), .ZN(new_n574));
  NAND4_X1  g388(.A1(new_n550), .A2(new_n566), .A3(KEYINPUT76), .A4(new_n551), .ZN(new_n575));
  INV_X1    g389(.A(new_n575), .ZN(new_n576));
  OAI21_X1  g390(.A(new_n523), .B1(new_n574), .B2(new_n576), .ZN(new_n577));
  XOR2_X1   g391(.A(new_n577), .B(KEYINPUT77), .Z(new_n578));
  OAI21_X1  g392(.A(new_n190), .B1(new_n574), .B2(new_n576), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n579), .A2(KEYINPUT25), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n567), .A2(new_n573), .ZN(new_n581));
  AOI21_X1  g395(.A(G902), .B1(new_n581), .B2(new_n575), .ZN(new_n582));
  INV_X1    g396(.A(KEYINPUT25), .ZN(new_n583));
  NAND2_X1  g397(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  XNOR2_X1  g398(.A(new_n522), .B(KEYINPUT71), .ZN(new_n585));
  NAND3_X1  g399(.A1(new_n580), .A2(new_n584), .A3(new_n585), .ZN(new_n586));
  NAND2_X1  g400(.A1(new_n578), .A2(new_n586), .ZN(new_n587));
  NAND3_X1  g401(.A1(new_n195), .A2(new_n200), .A3(new_n201), .ZN(new_n588));
  AOI21_X1  g402(.A(G134), .B1(new_n196), .B2(new_n198), .ZN(new_n589));
  INV_X1    g403(.A(KEYINPUT65), .ZN(new_n590));
  OAI21_X1  g404(.A(new_n590), .B1(new_n456), .B2(G137), .ZN(new_n591));
  NAND3_X1  g405(.A1(new_n192), .A2(KEYINPUT65), .A3(G134), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  OAI21_X1  g407(.A(G131), .B1(new_n589), .B2(new_n593), .ZN(new_n594));
  OAI211_X1 g408(.A(new_n588), .B(new_n594), .C1(new_n248), .C2(new_n227), .ZN(new_n595));
  OAI21_X1  g409(.A(new_n273), .B1(new_n202), .B2(new_n203), .ZN(new_n596));
  INV_X1    g410(.A(KEYINPUT30), .ZN(new_n597));
  AND3_X1   g411(.A1(new_n595), .A2(new_n596), .A3(new_n597), .ZN(new_n598));
  AOI21_X1  g412(.A(new_n597), .B1(new_n595), .B2(new_n596), .ZN(new_n599));
  OAI21_X1  g413(.A(new_n340), .B1(new_n598), .B2(new_n599), .ZN(new_n600));
  NAND3_X1  g414(.A1(new_n595), .A2(new_n596), .A3(new_n339), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n401), .A2(G210), .ZN(new_n602));
  XNOR2_X1  g416(.A(new_n602), .B(KEYINPUT27), .ZN(new_n603));
  XNOR2_X1  g417(.A(KEYINPUT26), .B(G101), .ZN(new_n604));
  XNOR2_X1  g418(.A(new_n603), .B(new_n604), .ZN(new_n605));
  NAND3_X1  g419(.A1(new_n600), .A2(new_n601), .A3(new_n605), .ZN(new_n606));
  INV_X1    g420(.A(KEYINPUT31), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  NAND4_X1  g422(.A1(new_n600), .A2(KEYINPUT31), .A3(new_n601), .A4(new_n605), .ZN(new_n609));
  NAND2_X1  g423(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  INV_X1    g424(.A(new_n601), .ZN(new_n611));
  AOI21_X1  g425(.A(new_n339), .B1(new_n595), .B2(new_n596), .ZN(new_n612));
  OAI21_X1  g426(.A(KEYINPUT28), .B1(new_n611), .B2(new_n612), .ZN(new_n613));
  INV_X1    g427(.A(KEYINPUT68), .ZN(new_n614));
  INV_X1    g428(.A(KEYINPUT28), .ZN(new_n615));
  AOI21_X1  g429(.A(new_n614), .B1(new_n601), .B2(new_n615), .ZN(new_n616));
  INV_X1    g430(.A(new_n616), .ZN(new_n617));
  NAND3_X1  g431(.A1(new_n601), .A2(new_n614), .A3(new_n615), .ZN(new_n618));
  NAND3_X1  g432(.A1(new_n613), .A2(new_n617), .A3(new_n618), .ZN(new_n619));
  INV_X1    g433(.A(new_n605), .ZN(new_n620));
  NAND2_X1  g434(.A1(new_n619), .A2(new_n620), .ZN(new_n621));
  NAND2_X1  g435(.A1(new_n610), .A2(new_n621), .ZN(new_n622));
  INV_X1    g436(.A(KEYINPUT32), .ZN(new_n623));
  INV_X1    g437(.A(G472), .ZN(new_n624));
  NAND4_X1  g438(.A1(new_n622), .A2(new_n623), .A3(new_n624), .A4(new_n190), .ZN(new_n625));
  AOI22_X1  g439(.A1(new_n608), .A2(new_n609), .B1(new_n619), .B2(new_n620), .ZN(new_n626));
  NAND2_X1  g440(.A1(new_n624), .A2(new_n190), .ZN(new_n627));
  OAI21_X1  g441(.A(KEYINPUT32), .B1(new_n626), .B2(new_n627), .ZN(new_n628));
  NAND2_X1  g442(.A1(new_n625), .A2(new_n628), .ZN(new_n629));
  INV_X1    g443(.A(new_n599), .ZN(new_n630));
  NAND3_X1  g444(.A1(new_n595), .A2(new_n596), .A3(new_n597), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n630), .A2(new_n631), .ZN(new_n632));
  AOI21_X1  g446(.A(new_n611), .B1(new_n632), .B2(new_n340), .ZN(new_n633));
  NOR3_X1   g447(.A1(new_n633), .A2(KEYINPUT69), .A3(new_n605), .ZN(new_n634));
  INV_X1    g448(.A(KEYINPUT29), .ZN(new_n635));
  OAI21_X1  g449(.A(new_n635), .B1(new_n619), .B2(new_n620), .ZN(new_n636));
  INV_X1    g450(.A(KEYINPUT69), .ZN(new_n637));
  NAND2_X1  g451(.A1(new_n600), .A2(new_n601), .ZN(new_n638));
  AOI21_X1  g452(.A(new_n637), .B1(new_n638), .B2(new_n620), .ZN(new_n639));
  NOR3_X1   g453(.A1(new_n634), .A2(new_n636), .A3(new_n639), .ZN(new_n640));
  INV_X1    g454(.A(new_n618), .ZN(new_n641));
  NOR2_X1   g455(.A1(new_n641), .A2(new_n616), .ZN(new_n642));
  NAND2_X1  g456(.A1(new_n595), .A2(new_n596), .ZN(new_n643));
  NAND2_X1  g457(.A1(new_n643), .A2(new_n340), .ZN(new_n644));
  INV_X1    g458(.A(KEYINPUT70), .ZN(new_n645));
  NAND3_X1  g459(.A1(new_n644), .A2(new_n645), .A3(new_n601), .ZN(new_n646));
  NAND2_X1  g460(.A1(new_n612), .A2(KEYINPUT70), .ZN(new_n647));
  NAND3_X1  g461(.A1(new_n646), .A2(KEYINPUT28), .A3(new_n647), .ZN(new_n648));
  NAND2_X1  g462(.A1(new_n642), .A2(new_n648), .ZN(new_n649));
  NAND2_X1  g463(.A1(new_n605), .A2(KEYINPUT29), .ZN(new_n650));
  OAI21_X1  g464(.A(new_n190), .B1(new_n649), .B2(new_n650), .ZN(new_n651));
  OAI21_X1  g465(.A(G472), .B1(new_n640), .B2(new_n651), .ZN(new_n652));
  AOI21_X1  g466(.A(new_n587), .B1(new_n629), .B2(new_n652), .ZN(new_n653));
  NAND2_X1  g467(.A1(new_n521), .A2(new_n653), .ZN(new_n654));
  XNOR2_X1  g468(.A(new_n654), .B(G101), .ZN(G3));
  NOR2_X1   g469(.A1(new_n305), .A2(new_n306), .ZN(new_n656));
  AOI21_X1  g470(.A(KEYINPUT85), .B1(new_n318), .B2(new_n304), .ZN(new_n657));
  OAI21_X1  g471(.A(new_n326), .B1(new_n656), .B2(new_n657), .ZN(new_n658));
  INV_X1    g472(.A(new_n191), .ZN(new_n659));
  NAND2_X1  g473(.A1(new_n622), .A2(new_n190), .ZN(new_n660));
  NAND2_X1  g474(.A1(new_n660), .A2(G472), .ZN(new_n661));
  OAI21_X1  g475(.A(new_n661), .B1(new_n626), .B2(new_n627), .ZN(new_n662));
  NOR2_X1   g476(.A1(new_n587), .A2(new_n662), .ZN(new_n663));
  NAND3_X1  g477(.A1(new_n658), .A2(new_n659), .A3(new_n663), .ZN(new_n664));
  INV_X1    g478(.A(KEYINPUT98), .ZN(new_n665));
  NAND2_X1  g479(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  NAND3_X1  g480(.A1(new_n327), .A2(KEYINPUT98), .A3(new_n663), .ZN(new_n667));
  AND2_X1   g481(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  AOI21_X1  g482(.A(new_n383), .B1(new_n370), .B2(new_n377), .ZN(new_n669));
  NAND2_X1  g483(.A1(new_n669), .A2(new_n518), .ZN(new_n670));
  AND3_X1   g484(.A1(new_n499), .A2(new_n502), .A3(new_n503), .ZN(new_n671));
  AOI21_X1  g485(.A(new_n503), .B1(new_n499), .B2(new_n502), .ZN(new_n672));
  INV_X1    g486(.A(KEYINPUT33), .ZN(new_n673));
  INV_X1    g487(.A(KEYINPUT99), .ZN(new_n674));
  AOI21_X1  g488(.A(new_n673), .B1(new_n494), .B2(new_n674), .ZN(new_n675));
  INV_X1    g489(.A(new_n675), .ZN(new_n676));
  NOR3_X1   g490(.A1(new_n671), .A2(new_n672), .A3(new_n676), .ZN(new_n677));
  AOI21_X1  g491(.A(new_n675), .B1(new_n495), .B2(new_n504), .ZN(new_n678));
  OAI21_X1  g492(.A(G478), .B1(new_n677), .B2(new_n678), .ZN(new_n679));
  NOR2_X1   g493(.A1(new_n506), .A2(new_n190), .ZN(new_n680));
  AOI21_X1  g494(.A(new_n680), .B1(new_n505), .B2(new_n506), .ZN(new_n681));
  NAND2_X1  g495(.A1(new_n679), .A2(new_n681), .ZN(new_n682));
  NAND2_X1  g496(.A1(new_n441), .A2(new_n442), .ZN(new_n683));
  NAND2_X1  g497(.A1(new_n683), .A2(KEYINPUT20), .ZN(new_n684));
  NAND3_X1  g498(.A1(new_n441), .A2(new_n384), .A3(new_n442), .ZN(new_n685));
  NAND2_X1  g499(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  NOR3_X1   g500(.A1(new_n448), .A2(new_n449), .A3(KEYINPUT92), .ZN(new_n687));
  NAND2_X1  g501(.A1(new_n439), .A2(new_n428), .ZN(new_n688));
  NAND3_X1  g502(.A1(new_n688), .A2(KEYINPUT92), .A3(new_n387), .ZN(new_n689));
  NAND2_X1  g503(.A1(new_n689), .A2(new_n190), .ZN(new_n690));
  OAI21_X1  g504(.A(G475), .B1(new_n687), .B2(new_n690), .ZN(new_n691));
  AOI21_X1  g505(.A(new_n682), .B1(new_n686), .B2(new_n691), .ZN(new_n692));
  INV_X1    g506(.A(new_n692), .ZN(new_n693));
  NOR2_X1   g507(.A1(new_n670), .A2(new_n693), .ZN(new_n694));
  NAND2_X1  g508(.A1(new_n668), .A2(new_n694), .ZN(new_n695));
  XOR2_X1   g509(.A(KEYINPUT34), .B(G104), .Z(new_n696));
  XNOR2_X1  g510(.A(new_n695), .B(new_n696), .ZN(G6));
  INV_X1    g511(.A(new_n508), .ZN(new_n698));
  NAND2_X1  g512(.A1(new_n453), .A2(new_n698), .ZN(new_n699));
  NOR2_X1   g513(.A1(new_n670), .A2(new_n699), .ZN(new_n700));
  NAND2_X1  g514(.A1(new_n668), .A2(new_n700), .ZN(new_n701));
  XNOR2_X1  g515(.A(new_n701), .B(KEYINPUT100), .ZN(new_n702));
  XOR2_X1   g516(.A(KEYINPUT35), .B(G107), .Z(new_n703));
  XNOR2_X1  g517(.A(new_n702), .B(new_n703), .ZN(G9));
  NAND2_X1  g518(.A1(new_n550), .A2(new_n551), .ZN(new_n705));
  NOR2_X1   g519(.A1(new_n566), .A2(KEYINPUT36), .ZN(new_n706));
  XOR2_X1   g520(.A(new_n705), .B(new_n706), .Z(new_n707));
  NAND2_X1  g521(.A1(new_n707), .A2(new_n523), .ZN(new_n708));
  OAI21_X1  g522(.A(new_n585), .B1(new_n582), .B2(new_n583), .ZN(new_n709));
  AOI211_X1 g523(.A(KEYINPUT25), .B(G902), .C1(new_n581), .C2(new_n575), .ZN(new_n710));
  OAI21_X1  g524(.A(new_n708), .B1(new_n709), .B2(new_n710), .ZN(new_n711));
  INV_X1    g525(.A(new_n711), .ZN(new_n712));
  NOR2_X1   g526(.A1(new_n662), .A2(new_n712), .ZN(new_n713));
  NAND2_X1  g527(.A1(new_n521), .A2(new_n713), .ZN(new_n714));
  XOR2_X1   g528(.A(KEYINPUT37), .B(G110), .Z(new_n715));
  XNOR2_X1  g529(.A(new_n714), .B(new_n715), .ZN(G12));
  NAND2_X1  g530(.A1(new_n629), .A2(new_n652), .ZN(new_n717));
  NAND2_X1  g531(.A1(new_n717), .A2(new_n711), .ZN(new_n718));
  NOR3_X1   g532(.A1(new_n362), .A2(new_n329), .A3(new_n369), .ZN(new_n719));
  OAI21_X1  g533(.A(new_n382), .B1(new_n719), .B2(new_n379), .ZN(new_n720));
  INV_X1    g534(.A(new_n515), .ZN(new_n721));
  OAI21_X1  g535(.A(new_n513), .B1(new_n721), .B2(G900), .ZN(new_n722));
  NAND3_X1  g536(.A1(new_n453), .A2(new_n698), .A3(new_n722), .ZN(new_n723));
  NOR3_X1   g537(.A1(new_n718), .A2(new_n720), .A3(new_n723), .ZN(new_n724));
  NAND2_X1  g538(.A1(new_n327), .A2(new_n724), .ZN(new_n725));
  XNOR2_X1  g539(.A(new_n725), .B(G128), .ZN(G30));
  XOR2_X1   g540(.A(new_n381), .B(KEYINPUT38), .Z(new_n727));
  NOR3_X1   g541(.A1(new_n453), .A2(new_n508), .A3(new_n383), .ZN(new_n728));
  NAND2_X1  g542(.A1(new_n712), .A2(new_n728), .ZN(new_n729));
  NAND2_X1  g543(.A1(new_n729), .A2(KEYINPUT102), .ZN(new_n730));
  OR2_X1    g544(.A1(new_n729), .A2(KEYINPUT102), .ZN(new_n731));
  NOR2_X1   g545(.A1(new_n633), .A2(new_n620), .ZN(new_n732));
  AOI21_X1  g546(.A(new_n605), .B1(new_n646), .B2(new_n647), .ZN(new_n733));
  NOR3_X1   g547(.A1(new_n732), .A2(G902), .A3(new_n733), .ZN(new_n734));
  OAI21_X1  g548(.A(new_n629), .B1(new_n624), .B2(new_n734), .ZN(new_n735));
  XNOR2_X1  g549(.A(new_n735), .B(KEYINPUT101), .ZN(new_n736));
  AND4_X1   g550(.A1(new_n727), .A2(new_n730), .A3(new_n731), .A4(new_n736), .ZN(new_n737));
  XNOR2_X1  g551(.A(new_n722), .B(KEYINPUT39), .ZN(new_n738));
  NAND2_X1  g552(.A1(new_n327), .A2(new_n738), .ZN(new_n739));
  OR2_X1    g553(.A1(new_n739), .A2(KEYINPUT40), .ZN(new_n740));
  NAND2_X1  g554(.A1(new_n739), .A2(KEYINPUT40), .ZN(new_n741));
  NAND3_X1  g555(.A1(new_n737), .A2(new_n740), .A3(new_n741), .ZN(new_n742));
  XNOR2_X1  g556(.A(new_n742), .B(G143), .ZN(G45));
  AOI22_X1  g557(.A1(new_n629), .A2(new_n652), .B1(new_n586), .B2(new_n708), .ZN(new_n744));
  INV_X1    g558(.A(new_n680), .ZN(new_n745));
  OAI21_X1  g559(.A(new_n190), .B1(new_n671), .B2(new_n672), .ZN(new_n746));
  OAI21_X1  g560(.A(new_n745), .B1(new_n746), .B2(G478), .ZN(new_n747));
  OAI21_X1  g561(.A(new_n676), .B1(new_n671), .B2(new_n672), .ZN(new_n748));
  NAND3_X1  g562(.A1(new_n495), .A2(new_n504), .A3(new_n675), .ZN(new_n749));
  AOI21_X1  g563(.A(new_n506), .B1(new_n748), .B2(new_n749), .ZN(new_n750));
  NOR2_X1   g564(.A1(new_n747), .A2(new_n750), .ZN(new_n751));
  OAI211_X1 g565(.A(new_n751), .B(new_n722), .C1(new_n446), .C2(new_n452), .ZN(new_n752));
  NAND2_X1  g566(.A1(new_n752), .A2(KEYINPUT103), .ZN(new_n753));
  OAI21_X1  g567(.A(new_n691), .B1(new_n443), .B2(new_n445), .ZN(new_n754));
  INV_X1    g568(.A(KEYINPUT103), .ZN(new_n755));
  NAND4_X1  g569(.A1(new_n754), .A2(new_n755), .A3(new_n751), .A4(new_n722), .ZN(new_n756));
  AND2_X1   g570(.A1(new_n753), .A2(new_n756), .ZN(new_n757));
  NAND3_X1  g571(.A1(new_n744), .A2(new_n757), .A3(new_n669), .ZN(new_n758));
  INV_X1    g572(.A(new_n758), .ZN(new_n759));
  NAND3_X1  g573(.A1(new_n759), .A2(new_n658), .A3(new_n659), .ZN(new_n760));
  INV_X1    g574(.A(KEYINPUT104), .ZN(new_n761));
  NAND2_X1  g575(.A1(new_n760), .A2(new_n761), .ZN(new_n762));
  NAND3_X1  g576(.A1(new_n327), .A2(KEYINPUT104), .A3(new_n759), .ZN(new_n763));
  NAND2_X1  g577(.A1(new_n762), .A2(new_n763), .ZN(new_n764));
  XNOR2_X1  g578(.A(new_n764), .B(G146), .ZN(G48));
  INV_X1    g579(.A(KEYINPUT106), .ZN(new_n766));
  NAND2_X1  g580(.A1(new_n303), .A2(new_n190), .ZN(new_n767));
  AOI21_X1  g581(.A(new_n191), .B1(new_n767), .B2(G469), .ZN(new_n768));
  OAI211_X1 g582(.A(KEYINPUT105), .B(new_n768), .C1(new_n656), .C2(new_n657), .ZN(new_n769));
  INV_X1    g583(.A(new_n769), .ZN(new_n770));
  AOI21_X1  g584(.A(KEYINPUT105), .B1(new_n320), .B2(new_n768), .ZN(new_n771));
  OAI21_X1  g585(.A(new_n766), .B1(new_n770), .B2(new_n771), .ZN(new_n772));
  OAI21_X1  g586(.A(new_n768), .B1(new_n656), .B2(new_n657), .ZN(new_n773));
  INV_X1    g587(.A(KEYINPUT105), .ZN(new_n774));
  NAND2_X1  g588(.A1(new_n773), .A2(new_n774), .ZN(new_n775));
  NAND3_X1  g589(.A1(new_n775), .A2(KEYINPUT106), .A3(new_n769), .ZN(new_n776));
  NAND4_X1  g590(.A1(new_n772), .A2(new_n776), .A3(new_n653), .A4(new_n694), .ZN(new_n777));
  XOR2_X1   g591(.A(KEYINPUT41), .B(G113), .Z(new_n778));
  XNOR2_X1  g592(.A(new_n778), .B(KEYINPUT107), .ZN(new_n779));
  XNOR2_X1  g593(.A(new_n777), .B(new_n779), .ZN(G15));
  AND2_X1   g594(.A1(new_n700), .A2(new_n653), .ZN(new_n781));
  NAND3_X1  g595(.A1(new_n772), .A2(new_n776), .A3(new_n781), .ZN(new_n782));
  XNOR2_X1  g596(.A(new_n782), .B(G116), .ZN(G18));
  NOR2_X1   g597(.A1(new_n770), .A2(new_n771), .ZN(new_n784));
  NOR3_X1   g598(.A1(new_n718), .A2(new_n720), .A3(new_n519), .ZN(new_n785));
  NAND2_X1  g599(.A1(new_n784), .A2(new_n785), .ZN(new_n786));
  XNOR2_X1  g600(.A(new_n786), .B(G119), .ZN(G21));
  INV_X1    g601(.A(new_n587), .ZN(new_n788));
  NAND2_X1  g602(.A1(new_n649), .A2(new_n620), .ZN(new_n789));
  AOI21_X1  g603(.A(new_n627), .B1(new_n789), .B2(new_n610), .ZN(new_n790));
  AOI21_X1  g604(.A(new_n790), .B1(new_n660), .B2(G472), .ZN(new_n791));
  NAND2_X1  g605(.A1(new_n788), .A2(new_n791), .ZN(new_n792));
  NAND2_X1  g606(.A1(new_n370), .A2(new_n377), .ZN(new_n793));
  NAND2_X1  g607(.A1(new_n793), .A2(new_n728), .ZN(new_n794));
  NOR3_X1   g608(.A1(new_n792), .A2(new_n517), .A3(new_n794), .ZN(new_n795));
  NAND3_X1  g609(.A1(new_n772), .A2(new_n776), .A3(new_n795), .ZN(new_n796));
  XNOR2_X1  g610(.A(new_n796), .B(G122), .ZN(G24));
  INV_X1    g611(.A(KEYINPUT109), .ZN(new_n798));
  AOI21_X1  g612(.A(new_n755), .B1(new_n692), .B2(new_n722), .ZN(new_n799));
  INV_X1    g613(.A(new_n756), .ZN(new_n800));
  OAI21_X1  g614(.A(new_n798), .B1(new_n799), .B2(new_n800), .ZN(new_n801));
  NAND3_X1  g615(.A1(new_n753), .A2(KEYINPUT109), .A3(new_n756), .ZN(new_n802));
  INV_X1    g616(.A(KEYINPUT108), .ZN(new_n803));
  AND3_X1   g617(.A1(new_n791), .A2(new_n711), .A3(new_n803), .ZN(new_n804));
  AOI21_X1  g618(.A(new_n803), .B1(new_n791), .B2(new_n711), .ZN(new_n805));
  OAI211_X1 g619(.A(new_n801), .B(new_n802), .C1(new_n804), .C2(new_n805), .ZN(new_n806));
  INV_X1    g620(.A(new_n806), .ZN(new_n807));
  NAND4_X1  g621(.A1(new_n775), .A2(new_n807), .A3(new_n669), .A4(new_n769), .ZN(new_n808));
  XNOR2_X1  g622(.A(new_n808), .B(G125), .ZN(G27));
  AOI21_X1  g623(.A(new_n383), .B1(new_n378), .B2(new_n380), .ZN(new_n810));
  AND3_X1   g624(.A1(new_n658), .A2(new_n659), .A3(new_n810), .ZN(new_n811));
  NAND2_X1  g625(.A1(new_n801), .A2(new_n802), .ZN(new_n812));
  INV_X1    g626(.A(new_n812), .ZN(new_n813));
  NAND4_X1  g627(.A1(new_n811), .A2(KEYINPUT42), .A3(new_n653), .A4(new_n813), .ZN(new_n814));
  INV_X1    g628(.A(KEYINPUT42), .ZN(new_n815));
  NAND4_X1  g629(.A1(new_n658), .A2(new_n653), .A3(new_n659), .A4(new_n810), .ZN(new_n816));
  OAI21_X1  g630(.A(new_n815), .B1(new_n816), .B2(new_n812), .ZN(new_n817));
  NAND2_X1  g631(.A1(new_n814), .A2(new_n817), .ZN(new_n818));
  XNOR2_X1  g632(.A(new_n818), .B(G131), .ZN(G33));
  INV_X1    g633(.A(new_n816), .ZN(new_n820));
  INV_X1    g634(.A(new_n723), .ZN(new_n821));
  NAND2_X1  g635(.A1(new_n820), .A2(new_n821), .ZN(new_n822));
  XOR2_X1   g636(.A(KEYINPUT110), .B(G134), .Z(new_n823));
  XNOR2_X1  g637(.A(new_n822), .B(new_n823), .ZN(G36));
  NAND2_X1  g638(.A1(new_n453), .A2(new_n751), .ZN(new_n825));
  XOR2_X1   g639(.A(new_n825), .B(KEYINPUT43), .Z(new_n826));
  NAND3_X1  g640(.A1(new_n826), .A2(new_n662), .A3(new_n711), .ZN(new_n827));
  XNOR2_X1  g641(.A(new_n827), .B(KEYINPUT44), .ZN(new_n828));
  NAND2_X1  g642(.A1(new_n828), .A2(new_n810), .ZN(new_n829));
  INV_X1    g643(.A(KEYINPUT45), .ZN(new_n830));
  AOI21_X1  g644(.A(new_n304), .B1(new_n324), .B2(new_n830), .ZN(new_n831));
  OAI21_X1  g645(.A(new_n831), .B1(new_n830), .B2(new_n324), .ZN(new_n832));
  NAND2_X1  g646(.A1(G469), .A2(G902), .ZN(new_n833));
  NAND2_X1  g647(.A1(new_n832), .A2(new_n833), .ZN(new_n834));
  INV_X1    g648(.A(KEYINPUT46), .ZN(new_n835));
  NAND2_X1  g649(.A1(new_n834), .A2(new_n835), .ZN(new_n836));
  NAND3_X1  g650(.A1(new_n832), .A2(KEYINPUT46), .A3(new_n833), .ZN(new_n837));
  NAND3_X1  g651(.A1(new_n836), .A2(new_n320), .A3(new_n837), .ZN(new_n838));
  NAND3_X1  g652(.A1(new_n838), .A2(new_n659), .A3(new_n738), .ZN(new_n839));
  NAND2_X1  g653(.A1(new_n839), .A2(KEYINPUT111), .ZN(new_n840));
  INV_X1    g654(.A(KEYINPUT111), .ZN(new_n841));
  NAND4_X1  g655(.A1(new_n838), .A2(new_n841), .A3(new_n659), .A4(new_n738), .ZN(new_n842));
  AOI21_X1  g656(.A(new_n829), .B1(new_n840), .B2(new_n842), .ZN(new_n843));
  XNOR2_X1  g657(.A(new_n843), .B(new_n192), .ZN(G39));
  NOR2_X1   g658(.A1(new_n788), .A2(new_n717), .ZN(new_n845));
  NAND3_X1  g659(.A1(new_n845), .A2(new_n757), .A3(new_n810), .ZN(new_n846));
  NAND2_X1  g660(.A1(new_n838), .A2(new_n659), .ZN(new_n847));
  INV_X1    g661(.A(KEYINPUT47), .ZN(new_n848));
  NAND2_X1  g662(.A1(new_n847), .A2(new_n848), .ZN(new_n849));
  NAND3_X1  g663(.A1(new_n838), .A2(KEYINPUT47), .A3(new_n659), .ZN(new_n850));
  AOI21_X1  g664(.A(new_n846), .B1(new_n849), .B2(new_n850), .ZN(new_n851));
  XNOR2_X1  g665(.A(new_n851), .B(new_n388), .ZN(G42));
  OR4_X1    g666(.A1(new_n587), .A2(new_n191), .A3(new_n383), .A4(new_n825), .ZN(new_n853));
  OAI21_X1  g667(.A(new_n320), .B1(new_n304), .B2(new_n318), .ZN(new_n854));
  AOI21_X1  g668(.A(new_n853), .B1(new_n854), .B2(KEYINPUT49), .ZN(new_n855));
  XOR2_X1   g669(.A(new_n855), .B(KEYINPUT112), .Z(new_n856));
  NOR2_X1   g670(.A1(new_n727), .A2(new_n736), .ZN(new_n857));
  OAI211_X1 g671(.A(new_n856), .B(new_n857), .C1(KEYINPUT49), .C2(new_n854), .ZN(new_n858));
  XNOR2_X1  g672(.A(new_n858), .B(KEYINPUT113), .ZN(new_n859));
  NAND2_X1  g673(.A1(new_n826), .A2(new_n514), .ZN(new_n860));
  OAI21_X1  g674(.A(new_n383), .B1(KEYINPUT116), .B2(KEYINPUT50), .ZN(new_n861));
  NOR4_X1   g675(.A1(new_n727), .A2(new_n792), .A3(new_n860), .A4(new_n861), .ZN(new_n862));
  NAND2_X1  g676(.A1(new_n862), .A2(new_n784), .ZN(new_n863));
  NAND2_X1  g677(.A1(KEYINPUT116), .A2(KEYINPUT50), .ZN(new_n864));
  XNOR2_X1  g678(.A(new_n863), .B(new_n864), .ZN(new_n865));
  OAI211_X1 g679(.A(new_n849), .B(new_n850), .C1(new_n659), .C2(new_n854), .ZN(new_n866));
  NOR2_X1   g680(.A1(new_n860), .A2(new_n792), .ZN(new_n867));
  NAND3_X1  g681(.A1(new_n866), .A2(new_n810), .A3(new_n867), .ZN(new_n868));
  AND2_X1   g682(.A1(new_n784), .A2(new_n810), .ZN(new_n869));
  INV_X1    g683(.A(new_n860), .ZN(new_n870));
  OAI211_X1 g684(.A(new_n869), .B(new_n870), .C1(new_n804), .C2(new_n805), .ZN(new_n871));
  NOR3_X1   g685(.A1(new_n736), .A2(new_n587), .A3(new_n513), .ZN(new_n872));
  NAND4_X1  g686(.A1(new_n869), .A2(new_n453), .A3(new_n682), .A4(new_n872), .ZN(new_n873));
  NAND4_X1  g687(.A1(new_n865), .A2(new_n868), .A3(new_n871), .A4(new_n873), .ZN(new_n874));
  INV_X1    g688(.A(KEYINPUT51), .ZN(new_n875));
  NOR2_X1   g689(.A1(new_n874), .A2(new_n875), .ZN(new_n876));
  NAND3_X1  g690(.A1(new_n869), .A2(new_n653), .A3(new_n870), .ZN(new_n877));
  AND2_X1   g691(.A1(new_n877), .A2(KEYINPUT48), .ZN(new_n878));
  NOR2_X1   g692(.A1(new_n877), .A2(KEYINPUT48), .ZN(new_n879));
  NOR2_X1   g693(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  NAND3_X1  g694(.A1(new_n869), .A2(new_n692), .A3(new_n872), .ZN(new_n881));
  NAND3_X1  g695(.A1(new_n784), .A2(new_n669), .A3(new_n867), .ZN(new_n882));
  NAND3_X1  g696(.A1(new_n881), .A2(new_n511), .A3(new_n882), .ZN(new_n883));
  NOR3_X1   g697(.A1(new_n876), .A2(new_n880), .A3(new_n883), .ZN(new_n884));
  INV_X1    g698(.A(KEYINPUT117), .ZN(new_n885));
  NAND3_X1  g699(.A1(new_n874), .A2(new_n885), .A3(new_n875), .ZN(new_n886));
  INV_X1    g700(.A(new_n886), .ZN(new_n887));
  AOI21_X1  g701(.A(new_n885), .B1(new_n874), .B2(new_n875), .ZN(new_n888));
  OAI21_X1  g702(.A(new_n884), .B1(new_n887), .B2(new_n888), .ZN(new_n889));
  INV_X1    g703(.A(KEYINPUT115), .ZN(new_n890));
  OAI211_X1 g704(.A(new_n772), .B(new_n776), .C1(new_n781), .C2(new_n795), .ZN(new_n891));
  AND3_X1   g705(.A1(new_n891), .A2(new_n777), .A3(new_n786), .ZN(new_n892));
  NAND3_X1  g706(.A1(new_n744), .A2(new_n510), .A3(new_n722), .ZN(new_n893));
  NAND2_X1  g707(.A1(new_n806), .A2(new_n893), .ZN(new_n894));
  AOI22_X1  g708(.A1(new_n820), .A2(new_n821), .B1(new_n811), .B2(new_n894), .ZN(new_n895));
  NAND2_X1  g709(.A1(new_n693), .A2(new_n699), .ZN(new_n896));
  NAND2_X1  g710(.A1(new_n896), .A2(new_n518), .ZN(new_n897));
  NOR3_X1   g711(.A1(new_n381), .A2(new_n383), .A3(new_n897), .ZN(new_n898));
  NAND3_X1  g712(.A1(new_n666), .A2(new_n667), .A3(new_n898), .ZN(new_n899));
  OAI21_X1  g713(.A(new_n521), .B1(new_n653), .B2(new_n713), .ZN(new_n900));
  AND3_X1   g714(.A1(new_n895), .A2(new_n899), .A3(new_n900), .ZN(new_n901));
  NAND4_X1  g715(.A1(new_n892), .A2(new_n901), .A3(KEYINPUT53), .A4(new_n818), .ZN(new_n902));
  AOI21_X1  g716(.A(KEYINPUT104), .B1(new_n327), .B2(new_n759), .ZN(new_n903));
  AOI21_X1  g717(.A(new_n325), .B1(new_n307), .B2(new_n319), .ZN(new_n904));
  NOR4_X1   g718(.A1(new_n904), .A2(new_n758), .A3(new_n761), .A4(new_n191), .ZN(new_n905));
  OAI211_X1 g719(.A(new_n808), .B(new_n725), .C1(new_n903), .C2(new_n905), .ZN(new_n906));
  INV_X1    g720(.A(new_n327), .ZN(new_n907));
  NAND3_X1  g721(.A1(new_n735), .A2(new_n712), .A3(new_n722), .ZN(new_n908));
  NOR3_X1   g722(.A1(new_n907), .A2(new_n794), .A3(new_n908), .ZN(new_n909));
  OAI21_X1  g723(.A(KEYINPUT52), .B1(new_n906), .B2(new_n909), .ZN(new_n910));
  AOI22_X1  g724(.A1(new_n762), .A2(new_n763), .B1(new_n327), .B2(new_n724), .ZN(new_n911));
  INV_X1    g725(.A(KEYINPUT52), .ZN(new_n912));
  OR3_X1    g726(.A1(new_n907), .A2(new_n794), .A3(new_n908), .ZN(new_n913));
  NAND4_X1  g727(.A1(new_n911), .A2(new_n912), .A3(new_n808), .A4(new_n913), .ZN(new_n914));
  NAND2_X1  g728(.A1(new_n910), .A2(new_n914), .ZN(new_n915));
  OAI21_X1  g729(.A(new_n890), .B1(new_n902), .B2(new_n915), .ZN(new_n916));
  AND2_X1   g730(.A1(new_n910), .A2(new_n914), .ZN(new_n917));
  NAND4_X1  g731(.A1(new_n818), .A2(new_n891), .A3(new_n777), .A4(new_n786), .ZN(new_n918));
  NAND4_X1  g732(.A1(new_n895), .A2(new_n900), .A3(new_n899), .A4(KEYINPUT53), .ZN(new_n919));
  NOR2_X1   g733(.A1(new_n918), .A2(new_n919), .ZN(new_n920));
  NAND3_X1  g734(.A1(new_n917), .A2(new_n920), .A3(KEYINPUT115), .ZN(new_n921));
  INV_X1    g735(.A(KEYINPUT53), .ZN(new_n922));
  INV_X1    g736(.A(new_n918), .ZN(new_n923));
  NAND4_X1  g737(.A1(new_n923), .A2(new_n910), .A3(new_n914), .A4(new_n901), .ZN(new_n924));
  AOI22_X1  g738(.A1(new_n916), .A2(new_n921), .B1(new_n922), .B2(new_n924), .ZN(new_n925));
  INV_X1    g739(.A(KEYINPUT54), .ZN(new_n926));
  NAND2_X1  g740(.A1(new_n925), .A2(new_n926), .ZN(new_n927));
  NAND2_X1  g741(.A1(new_n924), .A2(new_n922), .ZN(new_n928));
  NAND2_X1  g742(.A1(new_n917), .A2(new_n920), .ZN(new_n929));
  NAND2_X1  g743(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  NAND2_X1  g744(.A1(new_n930), .A2(KEYINPUT54), .ZN(new_n931));
  NAND3_X1  g745(.A1(new_n927), .A2(KEYINPUT114), .A3(new_n931), .ZN(new_n932));
  INV_X1    g746(.A(KEYINPUT114), .ZN(new_n933));
  NAND3_X1  g747(.A1(new_n930), .A2(new_n933), .A3(KEYINPUT54), .ZN(new_n934));
  AOI21_X1  g748(.A(new_n889), .B1(new_n932), .B2(new_n934), .ZN(new_n935));
  NOR2_X1   g749(.A1(G952), .A2(G953), .ZN(new_n936));
  OAI21_X1  g750(.A(new_n859), .B1(new_n935), .B2(new_n936), .ZN(G75));
  NOR3_X1   g751(.A1(new_n373), .A2(new_n374), .A3(new_n372), .ZN(new_n938));
  NOR2_X1   g752(.A1(new_n938), .A2(new_n362), .ZN(new_n939));
  XOR2_X1   g753(.A(new_n939), .B(KEYINPUT55), .Z(new_n940));
  INV_X1    g754(.A(new_n940), .ZN(new_n941));
  NOR4_X1   g755(.A1(new_n915), .A2(new_n890), .A3(new_n918), .A4(new_n919), .ZN(new_n942));
  AOI21_X1  g756(.A(KEYINPUT115), .B1(new_n917), .B2(new_n920), .ZN(new_n943));
  OAI21_X1  g757(.A(new_n928), .B1(new_n942), .B2(new_n943), .ZN(new_n944));
  NAND2_X1  g758(.A1(G210), .A2(G902), .ZN(new_n945));
  INV_X1    g759(.A(new_n945), .ZN(new_n946));
  NAND2_X1  g760(.A1(new_n944), .A2(new_n946), .ZN(new_n947));
  INV_X1    g761(.A(KEYINPUT118), .ZN(new_n948));
  AOI21_X1  g762(.A(KEYINPUT56), .B1(new_n947), .B2(new_n948), .ZN(new_n949));
  NAND3_X1  g763(.A1(new_n944), .A2(KEYINPUT118), .A3(new_n946), .ZN(new_n950));
  AOI21_X1  g764(.A(new_n941), .B1(new_n949), .B2(new_n950), .ZN(new_n951));
  NOR2_X1   g765(.A1(new_n398), .A2(G952), .ZN(new_n952));
  NOR2_X1   g766(.A1(new_n940), .A2(KEYINPUT56), .ZN(new_n953));
  AOI21_X1  g767(.A(new_n952), .B1(new_n947), .B2(new_n953), .ZN(new_n954));
  INV_X1    g768(.A(new_n954), .ZN(new_n955));
  OAI21_X1  g769(.A(KEYINPUT119), .B1(new_n951), .B2(new_n955), .ZN(new_n956));
  OAI21_X1  g770(.A(new_n948), .B1(new_n925), .B2(new_n945), .ZN(new_n957));
  INV_X1    g771(.A(KEYINPUT56), .ZN(new_n958));
  NAND3_X1  g772(.A1(new_n957), .A2(new_n950), .A3(new_n958), .ZN(new_n959));
  NAND2_X1  g773(.A1(new_n959), .A2(new_n940), .ZN(new_n960));
  INV_X1    g774(.A(KEYINPUT119), .ZN(new_n961));
  NAND3_X1  g775(.A1(new_n960), .A2(new_n961), .A3(new_n954), .ZN(new_n962));
  NAND2_X1  g776(.A1(new_n956), .A2(new_n962), .ZN(G51));
  NAND2_X1  g777(.A1(new_n944), .A2(KEYINPUT54), .ZN(new_n964));
  NAND3_X1  g778(.A1(new_n927), .A2(new_n964), .A3(KEYINPUT120), .ZN(new_n965));
  OR3_X1    g779(.A1(new_n925), .A2(KEYINPUT120), .A3(new_n926), .ZN(new_n966));
  XOR2_X1   g780(.A(new_n833), .B(KEYINPUT57), .Z(new_n967));
  NAND3_X1  g781(.A1(new_n965), .A2(new_n966), .A3(new_n967), .ZN(new_n968));
  NAND2_X1  g782(.A1(new_n968), .A2(new_n303), .ZN(new_n969));
  OR3_X1    g783(.A1(new_n925), .A2(new_n190), .A3(new_n832), .ZN(new_n970));
  AOI21_X1  g784(.A(new_n952), .B1(new_n969), .B2(new_n970), .ZN(G54));
  NAND4_X1  g785(.A1(new_n944), .A2(KEYINPUT58), .A3(G475), .A4(G902), .ZN(new_n972));
  INV_X1    g786(.A(new_n441), .ZN(new_n973));
  AND2_X1   g787(.A1(new_n972), .A2(new_n973), .ZN(new_n974));
  NOR2_X1   g788(.A1(new_n972), .A2(new_n973), .ZN(new_n975));
  NOR3_X1   g789(.A1(new_n974), .A2(new_n975), .A3(new_n952), .ZN(G60));
  XOR2_X1   g790(.A(new_n680), .B(KEYINPUT59), .Z(new_n977));
  NAND3_X1  g791(.A1(new_n932), .A2(new_n934), .A3(new_n977), .ZN(new_n978));
  NOR2_X1   g792(.A1(new_n677), .A2(new_n678), .ZN(new_n979));
  INV_X1    g793(.A(new_n979), .ZN(new_n980));
  NAND2_X1  g794(.A1(new_n978), .A2(new_n980), .ZN(new_n981));
  INV_X1    g795(.A(new_n952), .ZN(new_n982));
  NAND4_X1  g796(.A1(new_n965), .A2(new_n966), .A3(new_n979), .A4(new_n977), .ZN(new_n983));
  AND3_X1   g797(.A1(new_n981), .A2(new_n982), .A3(new_n983), .ZN(G63));
  NOR2_X1   g798(.A1(new_n574), .A2(new_n576), .ZN(new_n985));
  NAND2_X1  g799(.A1(G217), .A2(G902), .ZN(new_n986));
  XNOR2_X1  g800(.A(new_n986), .B(KEYINPUT60), .ZN(new_n987));
  OAI21_X1  g801(.A(new_n985), .B1(new_n925), .B2(new_n987), .ZN(new_n988));
  INV_X1    g802(.A(new_n987), .ZN(new_n989));
  NAND3_X1  g803(.A1(new_n944), .A2(new_n707), .A3(new_n989), .ZN(new_n990));
  NAND4_X1  g804(.A1(new_n988), .A2(KEYINPUT61), .A3(new_n990), .A4(new_n982), .ZN(new_n991));
  NAND2_X1  g805(.A1(new_n991), .A2(KEYINPUT122), .ZN(new_n992));
  NAND2_X1  g806(.A1(new_n944), .A2(new_n989), .ZN(new_n993));
  AOI21_X1  g807(.A(new_n952), .B1(new_n993), .B2(new_n985), .ZN(new_n994));
  INV_X1    g808(.A(KEYINPUT122), .ZN(new_n995));
  NAND4_X1  g809(.A1(new_n994), .A2(new_n995), .A3(KEYINPUT61), .A4(new_n990), .ZN(new_n996));
  NAND2_X1  g810(.A1(new_n992), .A2(new_n996), .ZN(new_n997));
  NAND3_X1  g811(.A1(new_n988), .A2(new_n982), .A3(new_n990), .ZN(new_n998));
  INV_X1    g812(.A(KEYINPUT61), .ZN(new_n999));
  AOI21_X1  g813(.A(KEYINPUT121), .B1(new_n998), .B2(new_n999), .ZN(new_n1000));
  AND3_X1   g814(.A1(new_n998), .A2(KEYINPUT121), .A3(new_n999), .ZN(new_n1001));
  OAI21_X1  g815(.A(new_n997), .B1(new_n1000), .B2(new_n1001), .ZN(G66));
  NAND3_X1  g816(.A1(new_n892), .A2(new_n899), .A3(new_n900), .ZN(new_n1003));
  NAND2_X1  g817(.A1(new_n1003), .A2(new_n398), .ZN(new_n1004));
  OAI21_X1  g818(.A(G953), .B1(new_n516), .B2(new_n332), .ZN(new_n1005));
  XOR2_X1   g819(.A(new_n1005), .B(KEYINPUT123), .Z(new_n1006));
  NAND2_X1  g820(.A1(new_n1004), .A2(new_n1006), .ZN(new_n1007));
  OAI211_X1 g821(.A(new_n360), .B(new_n361), .C1(G898), .C2(new_n398), .ZN(new_n1008));
  XNOR2_X1  g822(.A(new_n1007), .B(new_n1008), .ZN(G69));
  INV_X1    g823(.A(KEYINPUT125), .ZN(new_n1010));
  INV_X1    g824(.A(new_n906), .ZN(new_n1011));
  NAND2_X1  g825(.A1(new_n742), .A2(new_n1011), .ZN(new_n1012));
  NAND2_X1  g826(.A1(new_n1012), .A2(KEYINPUT62), .ZN(new_n1013));
  NOR2_X1   g827(.A1(new_n843), .A2(new_n851), .ZN(new_n1014));
  INV_X1    g828(.A(KEYINPUT62), .ZN(new_n1015));
  NAND3_X1  g829(.A1(new_n742), .A2(new_n1011), .A3(new_n1015), .ZN(new_n1016));
  INV_X1    g830(.A(new_n739), .ZN(new_n1017));
  NAND4_X1  g831(.A1(new_n1017), .A2(new_n653), .A3(new_n810), .A4(new_n896), .ZN(new_n1018));
  NAND4_X1  g832(.A1(new_n1013), .A2(new_n1014), .A3(new_n1016), .A4(new_n1018), .ZN(new_n1019));
  NAND2_X1  g833(.A1(new_n1019), .A2(new_n398), .ZN(new_n1020));
  NAND2_X1  g834(.A1(new_n411), .A2(new_n414), .ZN(new_n1021));
  XOR2_X1   g835(.A(new_n632), .B(new_n1021), .Z(new_n1022));
  XOR2_X1   g836(.A(new_n1022), .B(KEYINPUT124), .Z(new_n1023));
  INV_X1    g837(.A(new_n1023), .ZN(new_n1024));
  AOI21_X1  g838(.A(new_n1010), .B1(new_n1020), .B2(new_n1024), .ZN(new_n1025));
  AOI211_X1 g839(.A(KEYINPUT125), .B(new_n1023), .C1(new_n1019), .C2(new_n398), .ZN(new_n1026));
  NOR2_X1   g840(.A1(new_n398), .A2(G900), .ZN(new_n1027));
  NAND2_X1  g841(.A1(new_n818), .A2(new_n822), .ZN(new_n1028));
  INV_X1    g842(.A(KEYINPUT127), .ZN(new_n1029));
  XNOR2_X1  g843(.A(new_n1028), .B(new_n1029), .ZN(new_n1030));
  NAND2_X1  g844(.A1(new_n840), .A2(new_n842), .ZN(new_n1031));
  NAND4_X1  g845(.A1(new_n1031), .A2(new_n653), .A3(new_n793), .A4(new_n728), .ZN(new_n1032));
  NAND4_X1  g846(.A1(new_n1030), .A2(new_n1011), .A3(new_n1014), .A4(new_n1032), .ZN(new_n1033));
  AOI21_X1  g847(.A(new_n1027), .B1(new_n1033), .B2(new_n398), .ZN(new_n1034));
  INV_X1    g848(.A(new_n1022), .ZN(new_n1035));
  OAI22_X1  g849(.A1(new_n1025), .A2(new_n1026), .B1(new_n1034), .B2(new_n1035), .ZN(new_n1036));
  NAND2_X1  g850(.A1(new_n1036), .A2(KEYINPUT126), .ZN(new_n1037));
  INV_X1    g851(.A(KEYINPUT126), .ZN(new_n1038));
  OAI221_X1 g852(.A(new_n1038), .B1(new_n1034), .B2(new_n1035), .C1(new_n1025), .C2(new_n1026), .ZN(new_n1039));
  AOI21_X1  g853(.A(new_n1027), .B1(new_n287), .B2(G953), .ZN(new_n1040));
  AND3_X1   g854(.A1(new_n1037), .A2(new_n1039), .A3(new_n1040), .ZN(new_n1041));
  AOI21_X1  g855(.A(new_n1040), .B1(new_n1037), .B2(new_n1039), .ZN(new_n1042));
  NOR2_X1   g856(.A1(new_n1041), .A2(new_n1042), .ZN(G72));
  NAND2_X1  g857(.A1(G472), .A2(G902), .ZN(new_n1044));
  XOR2_X1   g858(.A(new_n1044), .B(KEYINPUT63), .Z(new_n1045));
  OAI21_X1  g859(.A(new_n1045), .B1(new_n1033), .B2(new_n1003), .ZN(new_n1046));
  NAND3_X1  g860(.A1(new_n1046), .A2(new_n620), .A3(new_n633), .ZN(new_n1047));
  INV_X1    g861(.A(new_n606), .ZN(new_n1048));
  OR2_X1    g862(.A1(new_n634), .A2(new_n639), .ZN(new_n1049));
  OAI211_X1 g863(.A(new_n930), .B(new_n1045), .C1(new_n1048), .C2(new_n1049), .ZN(new_n1050));
  NAND2_X1  g864(.A1(new_n1047), .A2(new_n1050), .ZN(new_n1051));
  OAI21_X1  g865(.A(new_n1045), .B1(new_n1019), .B2(new_n1003), .ZN(new_n1052));
  AOI211_X1 g866(.A(new_n952), .B(new_n1051), .C1(new_n732), .C2(new_n1052), .ZN(G57));
endmodule


