

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
         n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598,
         n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609,
         n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620,
         n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631,
         n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642,
         n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653,
         n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664,
         n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675,
         n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686,
         n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697,
         n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708,
         n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719,
         n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, n730,
         n731, n732, n733, n734, n735, n736, n737, n738, n739, n740, n741,
         n742, n743, n744, n745, n746, n747, n748, n749, n750, n751, n752,
         n753, n754, n755, n756, n757, n758, n759, n760, n761, n762, n763,
         n764, n765, n766, n767, n768, n769, n770, n771, n772, n773, n774,
         n775, n776, n777, n778, n779, n780, n781, n782, n783, n784, n785,
         n786, n787, n788, n789, n790, n791, n792, n793, n794, n795, n796,
         n797, n798, n799, n800, n801, n802, n803, n804, n805, n806, n807,
         n808, n809, n810, n811, n812, n813, n814, n815, n816, n817, n818,
         n819, n820, n821, n822, n823, n824, n825, n826, n827, n828, n829,
         n830, n831, n832, n833, n834, n835, n836, n837, n838, n839, n840,
         n841, n842, n843, n844, n845, n846, n847, n848, n849, n850, n851,
         n852, n853, n854, n855, n856, n857, n858, n859, n860, n861, n862,
         n863, n864, n865, n866, n867, n868, n869, n870, n871, n872, n873,
         n874, n875, n876, n877, n878, n879, n880, n881, n882, n883, n884,
         n885, n886, n887, n888, n889, n890, n891, n892, n893, n894, n895,
         n896, n897, n898, n899, n900, n901, n902, n903, n904, n905, n906,
         n907, n908, n909, n910, n911, n912, n913, n914, n915, n916, n917,
         n918, n919, n920, n921, n922, n923, n924, n925, n926, n927, n928,
         n929, n930, n931, n932, n933, n934, n935, n936, n937, n938, n939,
         n940, n941, n942, n943, n944, n945, n946, n947, n948, n949, n950,
         n951, n952, n953, n954, n955, n956, n957, n958, n959, n960, n961,
         n962, n963, n964, n965, n966, n967, n968, n969, n970, n971, n972,
         n973, n974, n975, n976, n977, n978, n979, n980, n981, n982, n983,
         n984, n985, n986, n987, n988, n989, n990, n991, n992, n993, n994,
         n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
         n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
         n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
         n1025;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  INV_X1 U552 ( .A(n727), .ZN(n708) );
  NOR2_X1 U553 ( .A1(G2105), .A2(G2104), .ZN(n523) );
  BUF_X2 U554 ( .A(n874), .Z(n518) );
  XOR2_X1 U555 ( .A(KEYINPUT17), .B(n523), .Z(n874) );
  AND2_X1 U556 ( .A1(G40), .A2(n682), .ZN(n753) );
  XNOR2_X1 U557 ( .A(n699), .B(KEYINPUT97), .ZN(n702) );
  AND2_X1 U558 ( .A1(n687), .A2(n686), .ZN(n693) );
  INV_X1 U559 ( .A(KEYINPUT100), .ZN(n696) );
  XOR2_X1 U560 ( .A(n698), .B(KEYINPUT27), .Z(n519) );
  OR2_X1 U561 ( .A1(n708), .A2(n990), .ZN(n520) );
  XOR2_X1 U562 ( .A(n703), .B(KEYINPUT28), .Z(n521) );
  NOR2_X1 U563 ( .A1(n745), .A2(n795), .ZN(n522) );
  XNOR2_X1 U564 ( .A(n717), .B(KEYINPUT103), .ZN(n718) );
  XNOR2_X1 U565 ( .A(n719), .B(n718), .ZN(n720) );
  NOR2_X1 U566 ( .A1(G651), .A2(n651), .ZN(n646) );
  XNOR2_X1 U567 ( .A(n535), .B(n534), .ZN(n682) );
  BUF_X1 U568 ( .A(n682), .Z(G160) );
  NAND2_X1 U569 ( .A1(G137), .A2(n518), .ZN(n525) );
  INV_X1 U570 ( .A(G2104), .ZN(n530) );
  AND2_X1 U571 ( .A1(G2105), .A2(G2104), .ZN(n869) );
  NAND2_X1 U572 ( .A1(G113), .A2(n869), .ZN(n524) );
  NAND2_X1 U573 ( .A1(n525), .A2(n524), .ZN(n526) );
  XNOR2_X1 U574 ( .A(n526), .B(KEYINPUT68), .ZN(n529) );
  NOR2_X2 U575 ( .A1(G2105), .A2(n530), .ZN(n873) );
  NAND2_X1 U576 ( .A1(G101), .A2(n873), .ZN(n527) );
  XNOR2_X1 U577 ( .A(KEYINPUT23), .B(n527), .ZN(n528) );
  NOR2_X1 U578 ( .A1(n529), .A2(n528), .ZN(n533) );
  NAND2_X1 U579 ( .A1(n530), .A2(G2105), .ZN(n531) );
  XNOR2_X1 U580 ( .A(n531), .B(KEYINPUT67), .ZN(n870) );
  NAND2_X1 U581 ( .A1(n870), .A2(G125), .ZN(n532) );
  NAND2_X1 U582 ( .A1(n533), .A2(n532), .ZN(n535) );
  INV_X1 U583 ( .A(KEYINPUT66), .ZN(n534) );
  NOR2_X1 U584 ( .A1(G651), .A2(G543), .ZN(n638) );
  NAND2_X1 U585 ( .A1(G85), .A2(n638), .ZN(n537) );
  XOR2_X1 U586 ( .A(KEYINPUT0), .B(G543), .Z(n651) );
  INV_X1 U587 ( .A(G651), .ZN(n538) );
  NOR2_X1 U588 ( .A1(n651), .A2(n538), .ZN(n636) );
  NAND2_X1 U589 ( .A1(G72), .A2(n636), .ZN(n536) );
  NAND2_X1 U590 ( .A1(n537), .A2(n536), .ZN(n543) );
  NOR2_X1 U591 ( .A1(G543), .A2(n538), .ZN(n539) );
  XOR2_X1 U592 ( .A(KEYINPUT1), .B(n539), .Z(n650) );
  NAND2_X1 U593 ( .A1(G60), .A2(n650), .ZN(n541) );
  NAND2_X1 U594 ( .A1(G47), .A2(n646), .ZN(n540) );
  NAND2_X1 U595 ( .A1(n541), .A2(n540), .ZN(n542) );
  OR2_X1 U596 ( .A1(n543), .A2(n542), .ZN(G290) );
  AND2_X1 U597 ( .A1(G452), .A2(G94), .ZN(G173) );
  NAND2_X1 U598 ( .A1(G123), .A2(n870), .ZN(n544) );
  XNOR2_X1 U599 ( .A(n544), .B(KEYINPUT18), .ZN(n551) );
  NAND2_X1 U600 ( .A1(G111), .A2(n869), .ZN(n546) );
  NAND2_X1 U601 ( .A1(G99), .A2(n873), .ZN(n545) );
  NAND2_X1 U602 ( .A1(n546), .A2(n545), .ZN(n549) );
  NAND2_X1 U603 ( .A1(n518), .A2(G135), .ZN(n547) );
  XOR2_X1 U604 ( .A(KEYINPUT80), .B(n547), .Z(n548) );
  NOR2_X1 U605 ( .A1(n549), .A2(n548), .ZN(n550) );
  NAND2_X1 U606 ( .A1(n551), .A2(n550), .ZN(n913) );
  XNOR2_X1 U607 ( .A(G2096), .B(n913), .ZN(n552) );
  OR2_X1 U608 ( .A1(G2100), .A2(n552), .ZN(G156) );
  INV_X1 U609 ( .A(G57), .ZN(G237) );
  INV_X1 U610 ( .A(G69), .ZN(G235) );
  INV_X1 U611 ( .A(G108), .ZN(G238) );
  INV_X1 U612 ( .A(G120), .ZN(G236) );
  INV_X1 U613 ( .A(G82), .ZN(G220) );
  NAND2_X1 U614 ( .A1(G64), .A2(n650), .ZN(n554) );
  NAND2_X1 U615 ( .A1(G52), .A2(n646), .ZN(n553) );
  NAND2_X1 U616 ( .A1(n554), .A2(n553), .ZN(n560) );
  NAND2_X1 U617 ( .A1(G90), .A2(n638), .ZN(n556) );
  NAND2_X1 U618 ( .A1(G77), .A2(n636), .ZN(n555) );
  NAND2_X1 U619 ( .A1(n556), .A2(n555), .ZN(n557) );
  XNOR2_X1 U620 ( .A(KEYINPUT69), .B(n557), .ZN(n558) );
  XNOR2_X1 U621 ( .A(KEYINPUT9), .B(n558), .ZN(n559) );
  NOR2_X1 U622 ( .A1(n560), .A2(n559), .ZN(G171) );
  INV_X1 U623 ( .A(G171), .ZN(G301) );
  NAND2_X1 U624 ( .A1(G88), .A2(n638), .ZN(n562) );
  NAND2_X1 U625 ( .A1(G75), .A2(n636), .ZN(n561) );
  NAND2_X1 U626 ( .A1(n562), .A2(n561), .ZN(n563) );
  XOR2_X1 U627 ( .A(KEYINPUT82), .B(n563), .Z(n567) );
  NAND2_X1 U628 ( .A1(G62), .A2(n650), .ZN(n565) );
  NAND2_X1 U629 ( .A1(G50), .A2(n646), .ZN(n564) );
  AND2_X1 U630 ( .A1(n565), .A2(n564), .ZN(n566) );
  NAND2_X1 U631 ( .A1(n567), .A2(n566), .ZN(G303) );
  NAND2_X1 U632 ( .A1(G114), .A2(n869), .ZN(n569) );
  NAND2_X1 U633 ( .A1(G102), .A2(n873), .ZN(n568) );
  NAND2_X1 U634 ( .A1(n569), .A2(n568), .ZN(n574) );
  NAND2_X1 U635 ( .A1(G138), .A2(n518), .ZN(n570) );
  XNOR2_X1 U636 ( .A(n570), .B(KEYINPUT88), .ZN(n572) );
  NAND2_X1 U637 ( .A1(n870), .A2(G126), .ZN(n571) );
  NAND2_X1 U638 ( .A1(n572), .A2(n571), .ZN(n573) );
  NOR2_X1 U639 ( .A1(n574), .A2(n573), .ZN(G164) );
  NAND2_X1 U640 ( .A1(n636), .A2(G76), .ZN(n575) );
  XNOR2_X1 U641 ( .A(KEYINPUT76), .B(n575), .ZN(n579) );
  XOR2_X1 U642 ( .A(KEYINPUT75), .B(KEYINPUT4), .Z(n577) );
  NAND2_X1 U643 ( .A1(G89), .A2(n638), .ZN(n576) );
  XNOR2_X1 U644 ( .A(n577), .B(n576), .ZN(n578) );
  NAND2_X1 U645 ( .A1(n579), .A2(n578), .ZN(n580) );
  XNOR2_X1 U646 ( .A(n580), .B(KEYINPUT5), .ZN(n586) );
  NAND2_X1 U647 ( .A1(n646), .A2(G51), .ZN(n581) );
  XOR2_X1 U648 ( .A(KEYINPUT77), .B(n581), .Z(n583) );
  NAND2_X1 U649 ( .A1(n650), .A2(G63), .ZN(n582) );
  NAND2_X1 U650 ( .A1(n583), .A2(n582), .ZN(n584) );
  XOR2_X1 U651 ( .A(KEYINPUT6), .B(n584), .Z(n585) );
  NAND2_X1 U652 ( .A1(n586), .A2(n585), .ZN(n587) );
  XNOR2_X1 U653 ( .A(n587), .B(KEYINPUT7), .ZN(G168) );
  XOR2_X1 U654 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U655 ( .A1(G7), .A2(G661), .ZN(n588) );
  XNOR2_X1 U656 ( .A(n588), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U657 ( .A(G223), .ZN(n818) );
  NAND2_X1 U658 ( .A1(n818), .A2(G567), .ZN(n589) );
  XOR2_X1 U659 ( .A(KEYINPUT11), .B(n589), .Z(G234) );
  XOR2_X1 U660 ( .A(KEYINPUT72), .B(KEYINPUT14), .Z(n591) );
  NAND2_X1 U661 ( .A1(G56), .A2(n650), .ZN(n590) );
  XNOR2_X1 U662 ( .A(n591), .B(n590), .ZN(n598) );
  XNOR2_X1 U663 ( .A(KEYINPUT73), .B(KEYINPUT13), .ZN(n596) );
  NAND2_X1 U664 ( .A1(n638), .A2(G81), .ZN(n592) );
  XNOR2_X1 U665 ( .A(n592), .B(KEYINPUT12), .ZN(n594) );
  NAND2_X1 U666 ( .A1(G68), .A2(n636), .ZN(n593) );
  NAND2_X1 U667 ( .A1(n594), .A2(n593), .ZN(n595) );
  XNOR2_X1 U668 ( .A(n596), .B(n595), .ZN(n597) );
  NOR2_X1 U669 ( .A1(n598), .A2(n597), .ZN(n600) );
  NAND2_X1 U670 ( .A1(n646), .A2(G43), .ZN(n599) );
  NAND2_X1 U671 ( .A1(n600), .A2(n599), .ZN(n973) );
  INV_X1 U672 ( .A(G860), .ZN(n620) );
  OR2_X1 U673 ( .A1(n973), .A2(n620), .ZN(G153) );
  INV_X1 U674 ( .A(G868), .ZN(n662) );
  NOR2_X1 U675 ( .A1(G301), .A2(n662), .ZN(n610) );
  NAND2_X1 U676 ( .A1(G66), .A2(n650), .ZN(n602) );
  NAND2_X1 U677 ( .A1(G92), .A2(n638), .ZN(n601) );
  NAND2_X1 U678 ( .A1(n602), .A2(n601), .ZN(n606) );
  NAND2_X1 U679 ( .A1(G79), .A2(n636), .ZN(n604) );
  NAND2_X1 U680 ( .A1(G54), .A2(n646), .ZN(n603) );
  NAND2_X1 U681 ( .A1(n604), .A2(n603), .ZN(n605) );
  NOR2_X1 U682 ( .A1(n606), .A2(n605), .ZN(n607) );
  XOR2_X1 U683 ( .A(KEYINPUT15), .B(n607), .Z(n608) );
  XNOR2_X1 U684 ( .A(KEYINPUT74), .B(n608), .ZN(n956) );
  AND2_X1 U685 ( .A1(n956), .A2(n662), .ZN(n609) );
  NOR2_X1 U686 ( .A1(n610), .A2(n609), .ZN(G284) );
  NAND2_X1 U687 ( .A1(G65), .A2(n650), .ZN(n612) );
  NAND2_X1 U688 ( .A1(G91), .A2(n638), .ZN(n611) );
  NAND2_X1 U689 ( .A1(n612), .A2(n611), .ZN(n615) );
  NAND2_X1 U690 ( .A1(n636), .A2(G78), .ZN(n613) );
  XOR2_X1 U691 ( .A(KEYINPUT70), .B(n613), .Z(n614) );
  NOR2_X1 U692 ( .A1(n615), .A2(n614), .ZN(n617) );
  NAND2_X1 U693 ( .A1(n646), .A2(G53), .ZN(n616) );
  NAND2_X1 U694 ( .A1(n617), .A2(n616), .ZN(G299) );
  NOR2_X1 U695 ( .A1(G286), .A2(n662), .ZN(n619) );
  NOR2_X1 U696 ( .A1(G868), .A2(G299), .ZN(n618) );
  NOR2_X1 U697 ( .A1(n619), .A2(n618), .ZN(G297) );
  NAND2_X1 U698 ( .A1(n620), .A2(G559), .ZN(n621) );
  NAND2_X1 U699 ( .A1(n621), .A2(n956), .ZN(n622) );
  XNOR2_X1 U700 ( .A(n622), .B(KEYINPUT16), .ZN(n623) );
  XNOR2_X1 U701 ( .A(KEYINPUT78), .B(n623), .ZN(G148) );
  NAND2_X1 U702 ( .A1(G868), .A2(n956), .ZN(n624) );
  XOR2_X1 U703 ( .A(KEYINPUT79), .B(n624), .Z(n625) );
  NOR2_X1 U704 ( .A1(G559), .A2(n625), .ZN(n627) );
  NOR2_X1 U705 ( .A1(G868), .A2(n973), .ZN(n626) );
  NOR2_X1 U706 ( .A1(n627), .A2(n626), .ZN(G282) );
  NAND2_X1 U707 ( .A1(n956), .A2(G559), .ZN(n628) );
  XNOR2_X1 U708 ( .A(n973), .B(n628), .ZN(n660) );
  NOR2_X1 U709 ( .A1(n660), .A2(G860), .ZN(n635) );
  NAND2_X1 U710 ( .A1(G67), .A2(n650), .ZN(n630) );
  NAND2_X1 U711 ( .A1(G55), .A2(n646), .ZN(n629) );
  NAND2_X1 U712 ( .A1(n630), .A2(n629), .ZN(n634) );
  NAND2_X1 U713 ( .A1(G93), .A2(n638), .ZN(n632) );
  NAND2_X1 U714 ( .A1(G80), .A2(n636), .ZN(n631) );
  NAND2_X1 U715 ( .A1(n632), .A2(n631), .ZN(n633) );
  NOR2_X1 U716 ( .A1(n634), .A2(n633), .ZN(n654) );
  XNOR2_X1 U717 ( .A(n635), .B(n654), .ZN(G145) );
  INV_X1 U718 ( .A(G303), .ZN(G166) );
  NAND2_X1 U719 ( .A1(G73), .A2(n636), .ZN(n637) );
  XOR2_X1 U720 ( .A(KEYINPUT2), .B(n637), .Z(n643) );
  NAND2_X1 U721 ( .A1(G61), .A2(n650), .ZN(n640) );
  NAND2_X1 U722 ( .A1(G86), .A2(n638), .ZN(n639) );
  NAND2_X1 U723 ( .A1(n640), .A2(n639), .ZN(n641) );
  XOR2_X1 U724 ( .A(KEYINPUT81), .B(n641), .Z(n642) );
  NOR2_X1 U725 ( .A1(n643), .A2(n642), .ZN(n645) );
  NAND2_X1 U726 ( .A1(n646), .A2(G48), .ZN(n644) );
  NAND2_X1 U727 ( .A1(n645), .A2(n644), .ZN(G305) );
  NAND2_X1 U728 ( .A1(G49), .A2(n646), .ZN(n648) );
  NAND2_X1 U729 ( .A1(G74), .A2(G651), .ZN(n647) );
  NAND2_X1 U730 ( .A1(n648), .A2(n647), .ZN(n649) );
  NOR2_X1 U731 ( .A1(n650), .A2(n649), .ZN(n653) );
  NAND2_X1 U732 ( .A1(n651), .A2(G87), .ZN(n652) );
  NAND2_X1 U733 ( .A1(n653), .A2(n652), .ZN(G288) );
  NOR2_X1 U734 ( .A1(G868), .A2(n654), .ZN(n664) );
  XNOR2_X1 U735 ( .A(n654), .B(G305), .ZN(n655) );
  XNOR2_X1 U736 ( .A(n655), .B(G288), .ZN(n656) );
  XNOR2_X1 U737 ( .A(KEYINPUT19), .B(n656), .ZN(n658) );
  INV_X1 U738 ( .A(G299), .ZN(n959) );
  XNOR2_X1 U739 ( .A(G290), .B(n959), .ZN(n657) );
  XNOR2_X1 U740 ( .A(n658), .B(n657), .ZN(n659) );
  XNOR2_X1 U741 ( .A(G166), .B(n659), .ZN(n897) );
  XOR2_X1 U742 ( .A(n660), .B(n897), .Z(n661) );
  NOR2_X1 U743 ( .A1(n662), .A2(n661), .ZN(n663) );
  NOR2_X1 U744 ( .A1(n664), .A2(n663), .ZN(n665) );
  XNOR2_X1 U745 ( .A(n665), .B(KEYINPUT83), .ZN(G295) );
  NAND2_X1 U746 ( .A1(G2078), .A2(G2084), .ZN(n666) );
  XOR2_X1 U747 ( .A(KEYINPUT20), .B(n666), .Z(n667) );
  NAND2_X1 U748 ( .A1(G2090), .A2(n667), .ZN(n668) );
  XNOR2_X1 U749 ( .A(KEYINPUT21), .B(n668), .ZN(n669) );
  NAND2_X1 U750 ( .A1(n669), .A2(G2072), .ZN(n670) );
  XNOR2_X1 U751 ( .A(KEYINPUT84), .B(n670), .ZN(G158) );
  XNOR2_X1 U752 ( .A(KEYINPUT71), .B(G132), .ZN(G219) );
  XNOR2_X1 U753 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U754 ( .A1(G220), .A2(G219), .ZN(n672) );
  XNOR2_X1 U755 ( .A(KEYINPUT22), .B(KEYINPUT85), .ZN(n671) );
  XNOR2_X1 U756 ( .A(n672), .B(n671), .ZN(n673) );
  NOR2_X1 U757 ( .A1(n673), .A2(G218), .ZN(n674) );
  NAND2_X1 U758 ( .A1(G96), .A2(n674), .ZN(n822) );
  NAND2_X1 U759 ( .A1(G2106), .A2(n822), .ZN(n680) );
  NOR2_X1 U760 ( .A1(G236), .A2(G238), .ZN(n676) );
  NOR2_X1 U761 ( .A1(G235), .A2(G237), .ZN(n675) );
  NAND2_X1 U762 ( .A1(n676), .A2(n675), .ZN(n677) );
  XNOR2_X1 U763 ( .A(KEYINPUT86), .B(n677), .ZN(n823) );
  NAND2_X1 U764 ( .A1(n823), .A2(G567), .ZN(n678) );
  XOR2_X1 U765 ( .A(KEYINPUT87), .B(n678), .Z(n679) );
  NAND2_X1 U766 ( .A1(n680), .A2(n679), .ZN(n908) );
  NAND2_X1 U767 ( .A1(G483), .A2(G661), .ZN(n681) );
  NOR2_X1 U768 ( .A1(n908), .A2(n681), .ZN(n821) );
  NAND2_X1 U769 ( .A1(n821), .A2(G36), .ZN(G176) );
  NOR2_X1 U770 ( .A1(G164), .A2(G1384), .ZN(n755) );
  NAND2_X2 U771 ( .A1(n753), .A2(n755), .ZN(n727) );
  XOR2_X1 U772 ( .A(G1996), .B(KEYINPUT98), .Z(n940) );
  NOR2_X1 U773 ( .A1(n727), .A2(n940), .ZN(n684) );
  XNOR2_X1 U774 ( .A(KEYINPUT65), .B(KEYINPUT26), .ZN(n683) );
  XNOR2_X1 U775 ( .A(n684), .B(n683), .ZN(n687) );
  AND2_X1 U776 ( .A1(n727), .A2(G1341), .ZN(n685) );
  NOR2_X1 U777 ( .A1(n685), .A2(n973), .ZN(n686) );
  NAND2_X1 U778 ( .A1(n693), .A2(n956), .ZN(n691) );
  NOR2_X1 U779 ( .A1(n708), .A2(G1348), .ZN(n689) );
  NOR2_X1 U780 ( .A1(G2067), .A2(n727), .ZN(n688) );
  NOR2_X1 U781 ( .A1(n689), .A2(n688), .ZN(n690) );
  NAND2_X1 U782 ( .A1(n691), .A2(n690), .ZN(n692) );
  XNOR2_X1 U783 ( .A(n692), .B(KEYINPUT99), .ZN(n695) );
  NOR2_X1 U784 ( .A1(n956), .A2(n693), .ZN(n694) );
  NOR2_X1 U785 ( .A1(n695), .A2(n694), .ZN(n697) );
  XNOR2_X1 U786 ( .A(n697), .B(n696), .ZN(n701) );
  NAND2_X1 U787 ( .A1(n708), .A2(G2072), .ZN(n698) );
  XOR2_X1 U788 ( .A(G1956), .B(KEYINPUT96), .Z(n990) );
  NAND2_X1 U789 ( .A1(n519), .A2(n520), .ZN(n699) );
  NAND2_X1 U790 ( .A1(n702), .A2(n959), .ZN(n700) );
  NAND2_X1 U791 ( .A1(n701), .A2(n700), .ZN(n704) );
  NOR2_X1 U792 ( .A1(n702), .A2(n959), .ZN(n703) );
  NAND2_X1 U793 ( .A1(n704), .A2(n521), .ZN(n706) );
  XNOR2_X1 U794 ( .A(KEYINPUT29), .B(KEYINPUT101), .ZN(n705) );
  XNOR2_X1 U795 ( .A(n706), .B(n705), .ZN(n713) );
  XNOR2_X1 U796 ( .A(G1961), .B(KEYINPUT93), .ZN(n1000) );
  NAND2_X1 U797 ( .A1(n727), .A2(n1000), .ZN(n707) );
  XNOR2_X1 U798 ( .A(n707), .B(KEYINPUT94), .ZN(n710) );
  XNOR2_X1 U799 ( .A(KEYINPUT25), .B(G2078), .ZN(n941) );
  NAND2_X1 U800 ( .A1(n708), .A2(n941), .ZN(n709) );
  NAND2_X1 U801 ( .A1(n710), .A2(n709), .ZN(n721) );
  AND2_X1 U802 ( .A1(n721), .A2(G171), .ZN(n711) );
  XNOR2_X1 U803 ( .A(KEYINPUT95), .B(n711), .ZN(n712) );
  NAND2_X1 U804 ( .A1(n713), .A2(n712), .ZN(n726) );
  NAND2_X1 U805 ( .A1(G8), .A2(n727), .ZN(n795) );
  NOR2_X1 U806 ( .A1(G1966), .A2(n795), .ZN(n737) );
  NOR2_X1 U807 ( .A1(n727), .A2(G2084), .ZN(n714) );
  XNOR2_X1 U808 ( .A(n714), .B(KEYINPUT92), .ZN(n736) );
  NOR2_X1 U809 ( .A1(n737), .A2(n736), .ZN(n715) );
  XNOR2_X1 U810 ( .A(n715), .B(KEYINPUT102), .ZN(n716) );
  NAND2_X1 U811 ( .A1(n716), .A2(G8), .ZN(n719) );
  INV_X1 U812 ( .A(KEYINPUT30), .ZN(n717) );
  NOR2_X1 U813 ( .A1(G168), .A2(n720), .ZN(n723) );
  NOR2_X1 U814 ( .A1(G171), .A2(n721), .ZN(n722) );
  NOR2_X1 U815 ( .A1(n723), .A2(n722), .ZN(n724) );
  XOR2_X1 U816 ( .A(KEYINPUT31), .B(n724), .Z(n725) );
  NAND2_X1 U817 ( .A1(n726), .A2(n725), .ZN(n738) );
  NAND2_X1 U818 ( .A1(n738), .A2(G286), .ZN(n734) );
  INV_X1 U819 ( .A(G8), .ZN(n732) );
  NOR2_X1 U820 ( .A1(G1971), .A2(n795), .ZN(n729) );
  NOR2_X1 U821 ( .A1(G2090), .A2(n727), .ZN(n728) );
  NOR2_X1 U822 ( .A1(n729), .A2(n728), .ZN(n730) );
  NAND2_X1 U823 ( .A1(G303), .A2(n730), .ZN(n731) );
  OR2_X1 U824 ( .A1(n732), .A2(n731), .ZN(n733) );
  AND2_X1 U825 ( .A1(n734), .A2(n733), .ZN(n735) );
  XNOR2_X1 U826 ( .A(n735), .B(KEYINPUT32), .ZN(n743) );
  NAND2_X1 U827 ( .A1(n736), .A2(G8), .ZN(n741) );
  INV_X1 U828 ( .A(n738), .ZN(n739) );
  NOR2_X1 U829 ( .A1(n737), .A2(n739), .ZN(n740) );
  NAND2_X1 U830 ( .A1(n741), .A2(n740), .ZN(n742) );
  NAND2_X1 U831 ( .A1(n743), .A2(n742), .ZN(n790) );
  NOR2_X1 U832 ( .A1(G1976), .A2(G288), .ZN(n749) );
  NOR2_X1 U833 ( .A1(G1971), .A2(G303), .ZN(n744) );
  NOR2_X1 U834 ( .A1(n749), .A2(n744), .ZN(n962) );
  NAND2_X1 U835 ( .A1(n790), .A2(n962), .ZN(n746) );
  NAND2_X1 U836 ( .A1(G1976), .A2(G288), .ZN(n961) );
  INV_X1 U837 ( .A(n961), .ZN(n745) );
  AND2_X1 U838 ( .A1(n746), .A2(n522), .ZN(n747) );
  XNOR2_X1 U839 ( .A(n747), .B(KEYINPUT64), .ZN(n748) );
  NOR2_X1 U840 ( .A1(KEYINPUT33), .A2(n748), .ZN(n752) );
  NAND2_X1 U841 ( .A1(n749), .A2(KEYINPUT33), .ZN(n750) );
  NOR2_X1 U842 ( .A1(n750), .A2(n795), .ZN(n751) );
  NOR2_X1 U843 ( .A1(n752), .A2(n751), .ZN(n787) );
  XOR2_X1 U844 ( .A(G1981), .B(G305), .Z(n969) );
  INV_X1 U845 ( .A(n753), .ZN(n754) );
  NOR2_X1 U846 ( .A1(n755), .A2(n754), .ZN(n813) );
  XNOR2_X1 U847 ( .A(G2067), .B(KEYINPUT37), .ZN(n811) );
  NAND2_X1 U848 ( .A1(n518), .A2(G140), .ZN(n756) );
  XOR2_X1 U849 ( .A(KEYINPUT89), .B(n756), .Z(n758) );
  NAND2_X1 U850 ( .A1(n873), .A2(G104), .ZN(n757) );
  NAND2_X1 U851 ( .A1(n758), .A2(n757), .ZN(n759) );
  XNOR2_X1 U852 ( .A(KEYINPUT34), .B(n759), .ZN(n764) );
  NAND2_X1 U853 ( .A1(G116), .A2(n869), .ZN(n761) );
  NAND2_X1 U854 ( .A1(G128), .A2(n870), .ZN(n760) );
  NAND2_X1 U855 ( .A1(n761), .A2(n760), .ZN(n762) );
  XOR2_X1 U856 ( .A(KEYINPUT35), .B(n762), .Z(n763) );
  NOR2_X1 U857 ( .A1(n764), .A2(n763), .ZN(n765) );
  XNOR2_X1 U858 ( .A(KEYINPUT36), .B(n765), .ZN(n894) );
  NOR2_X1 U859 ( .A1(n811), .A2(n894), .ZN(n928) );
  NAND2_X1 U860 ( .A1(n813), .A2(n928), .ZN(n809) );
  NAND2_X1 U861 ( .A1(G95), .A2(n873), .ZN(n767) );
  NAND2_X1 U862 ( .A1(G131), .A2(n518), .ZN(n766) );
  NAND2_X1 U863 ( .A1(n767), .A2(n766), .ZN(n771) );
  NAND2_X1 U864 ( .A1(G107), .A2(n869), .ZN(n769) );
  NAND2_X1 U865 ( .A1(G119), .A2(n870), .ZN(n768) );
  NAND2_X1 U866 ( .A1(n769), .A2(n768), .ZN(n770) );
  NOR2_X1 U867 ( .A1(n771), .A2(n770), .ZN(n885) );
  INV_X1 U868 ( .A(G1991), .ZN(n936) );
  NOR2_X1 U869 ( .A1(n885), .A2(n936), .ZN(n782) );
  NAND2_X1 U870 ( .A1(G141), .A2(n518), .ZN(n772) );
  XNOR2_X1 U871 ( .A(n772), .B(KEYINPUT90), .ZN(n779) );
  NAND2_X1 U872 ( .A1(G117), .A2(n869), .ZN(n774) );
  NAND2_X1 U873 ( .A1(G129), .A2(n870), .ZN(n773) );
  NAND2_X1 U874 ( .A1(n774), .A2(n773), .ZN(n777) );
  NAND2_X1 U875 ( .A1(n873), .A2(G105), .ZN(n775) );
  XOR2_X1 U876 ( .A(KEYINPUT38), .B(n775), .Z(n776) );
  NOR2_X1 U877 ( .A1(n777), .A2(n776), .ZN(n778) );
  NAND2_X1 U878 ( .A1(n779), .A2(n778), .ZN(n780) );
  XOR2_X1 U879 ( .A(KEYINPUT91), .B(n780), .Z(n889) );
  AND2_X1 U880 ( .A1(G1996), .A2(n889), .ZN(n781) );
  NOR2_X1 U881 ( .A1(n782), .A2(n781), .ZN(n918) );
  INV_X1 U882 ( .A(n813), .ZN(n783) );
  NOR2_X1 U883 ( .A1(n918), .A2(n783), .ZN(n806) );
  INV_X1 U884 ( .A(n806), .ZN(n784) );
  NAND2_X1 U885 ( .A1(n809), .A2(n784), .ZN(n799) );
  INV_X1 U886 ( .A(n799), .ZN(n785) );
  AND2_X1 U887 ( .A1(n969), .A2(n785), .ZN(n786) );
  NAND2_X1 U888 ( .A1(n787), .A2(n786), .ZN(n801) );
  NOR2_X1 U889 ( .A1(G2090), .A2(G303), .ZN(n788) );
  XNOR2_X1 U890 ( .A(n788), .B(KEYINPUT104), .ZN(n789) );
  NAND2_X1 U891 ( .A1(n789), .A2(G8), .ZN(n791) );
  NAND2_X1 U892 ( .A1(n791), .A2(n790), .ZN(n792) );
  AND2_X1 U893 ( .A1(n792), .A2(n795), .ZN(n797) );
  NOR2_X1 U894 ( .A1(G1981), .A2(G305), .ZN(n793) );
  XOR2_X1 U895 ( .A(n793), .B(KEYINPUT24), .Z(n794) );
  NOR2_X1 U896 ( .A1(n795), .A2(n794), .ZN(n796) );
  NOR2_X1 U897 ( .A1(n797), .A2(n796), .ZN(n798) );
  OR2_X1 U898 ( .A1(n799), .A2(n798), .ZN(n800) );
  NAND2_X1 U899 ( .A1(n801), .A2(n800), .ZN(n803) );
  XNOR2_X1 U900 ( .A(G1986), .B(G290), .ZN(n958) );
  NAND2_X1 U901 ( .A1(n958), .A2(n813), .ZN(n802) );
  NAND2_X1 U902 ( .A1(n803), .A2(n802), .ZN(n816) );
  NOR2_X1 U903 ( .A1(G1996), .A2(n889), .ZN(n920) );
  AND2_X1 U904 ( .A1(n936), .A2(n885), .ZN(n916) );
  NOR2_X1 U905 ( .A1(G1986), .A2(G290), .ZN(n804) );
  NOR2_X1 U906 ( .A1(n916), .A2(n804), .ZN(n805) );
  NOR2_X1 U907 ( .A1(n806), .A2(n805), .ZN(n807) );
  NOR2_X1 U908 ( .A1(n920), .A2(n807), .ZN(n808) );
  XNOR2_X1 U909 ( .A(KEYINPUT39), .B(n808), .ZN(n810) );
  NAND2_X1 U910 ( .A1(n810), .A2(n809), .ZN(n812) );
  NAND2_X1 U911 ( .A1(n811), .A2(n894), .ZN(n925) );
  NAND2_X1 U912 ( .A1(n812), .A2(n925), .ZN(n814) );
  NAND2_X1 U913 ( .A1(n814), .A2(n813), .ZN(n815) );
  NAND2_X1 U914 ( .A1(n816), .A2(n815), .ZN(n817) );
  XNOR2_X1 U915 ( .A(KEYINPUT40), .B(n817), .ZN(G329) );
  NAND2_X1 U916 ( .A1(G2106), .A2(n818), .ZN(G217) );
  AND2_X1 U917 ( .A1(G15), .A2(G2), .ZN(n819) );
  NAND2_X1 U918 ( .A1(G661), .A2(n819), .ZN(G259) );
  NAND2_X1 U919 ( .A1(G3), .A2(G1), .ZN(n820) );
  NAND2_X1 U920 ( .A1(n821), .A2(n820), .ZN(G188) );
  INV_X1 U922 ( .A(G96), .ZN(G221) );
  NOR2_X1 U923 ( .A1(n823), .A2(n822), .ZN(G325) );
  INV_X1 U924 ( .A(G325), .ZN(G261) );
  XOR2_X1 U925 ( .A(G2454), .B(G2435), .Z(n825) );
  XNOR2_X1 U926 ( .A(G2438), .B(G2427), .ZN(n824) );
  XNOR2_X1 U927 ( .A(n825), .B(n824), .ZN(n832) );
  XOR2_X1 U928 ( .A(KEYINPUT105), .B(G2446), .Z(n827) );
  XNOR2_X1 U929 ( .A(G2443), .B(G2430), .ZN(n826) );
  XNOR2_X1 U930 ( .A(n827), .B(n826), .ZN(n828) );
  XOR2_X1 U931 ( .A(n828), .B(G2451), .Z(n830) );
  XNOR2_X1 U932 ( .A(G1341), .B(G1348), .ZN(n829) );
  XNOR2_X1 U933 ( .A(n830), .B(n829), .ZN(n831) );
  XNOR2_X1 U934 ( .A(n832), .B(n831), .ZN(n833) );
  NAND2_X1 U935 ( .A1(n833), .A2(G14), .ZN(n834) );
  XOR2_X1 U936 ( .A(KEYINPUT106), .B(n834), .Z(G401) );
  XOR2_X1 U937 ( .A(G2100), .B(G2096), .Z(n836) );
  XNOR2_X1 U938 ( .A(KEYINPUT42), .B(G2678), .ZN(n835) );
  XNOR2_X1 U939 ( .A(n836), .B(n835), .ZN(n840) );
  XOR2_X1 U940 ( .A(KEYINPUT43), .B(G2090), .Z(n838) );
  XNOR2_X1 U941 ( .A(G2067), .B(G2072), .ZN(n837) );
  XNOR2_X1 U942 ( .A(n838), .B(n837), .ZN(n839) );
  XOR2_X1 U943 ( .A(n840), .B(n839), .Z(n842) );
  XNOR2_X1 U944 ( .A(G2078), .B(G2084), .ZN(n841) );
  XNOR2_X1 U945 ( .A(n842), .B(n841), .ZN(G227) );
  XOR2_X1 U946 ( .A(G1976), .B(G1971), .Z(n844) );
  XNOR2_X1 U947 ( .A(G1986), .B(G1961), .ZN(n843) );
  XNOR2_X1 U948 ( .A(n844), .B(n843), .ZN(n848) );
  XOR2_X1 U949 ( .A(G1981), .B(G1966), .Z(n846) );
  XNOR2_X1 U950 ( .A(G1996), .B(G1991), .ZN(n845) );
  XNOR2_X1 U951 ( .A(n846), .B(n845), .ZN(n847) );
  XOR2_X1 U952 ( .A(n848), .B(n847), .Z(n850) );
  XNOR2_X1 U953 ( .A(KEYINPUT41), .B(KEYINPUT107), .ZN(n849) );
  XNOR2_X1 U954 ( .A(n850), .B(n849), .ZN(n852) );
  XOR2_X1 U955 ( .A(G1956), .B(G2474), .Z(n851) );
  XNOR2_X1 U956 ( .A(n852), .B(n851), .ZN(G229) );
  NAND2_X1 U957 ( .A1(n873), .A2(G100), .ZN(n853) );
  XNOR2_X1 U958 ( .A(n853), .B(KEYINPUT108), .ZN(n855) );
  NAND2_X1 U959 ( .A1(G112), .A2(n869), .ZN(n854) );
  NAND2_X1 U960 ( .A1(n855), .A2(n854), .ZN(n856) );
  XNOR2_X1 U961 ( .A(n856), .B(KEYINPUT109), .ZN(n858) );
  NAND2_X1 U962 ( .A1(G136), .A2(n518), .ZN(n857) );
  NAND2_X1 U963 ( .A1(n858), .A2(n857), .ZN(n861) );
  NAND2_X1 U964 ( .A1(n870), .A2(G124), .ZN(n859) );
  XOR2_X1 U965 ( .A(KEYINPUT44), .B(n859), .Z(n860) );
  NOR2_X1 U966 ( .A1(n861), .A2(n860), .ZN(G162) );
  NAND2_X1 U967 ( .A1(G103), .A2(n873), .ZN(n863) );
  NAND2_X1 U968 ( .A1(G139), .A2(n518), .ZN(n862) );
  NAND2_X1 U969 ( .A1(n863), .A2(n862), .ZN(n868) );
  NAND2_X1 U970 ( .A1(G115), .A2(n869), .ZN(n865) );
  NAND2_X1 U971 ( .A1(G127), .A2(n870), .ZN(n864) );
  NAND2_X1 U972 ( .A1(n865), .A2(n864), .ZN(n866) );
  XOR2_X1 U973 ( .A(KEYINPUT47), .B(n866), .Z(n867) );
  NOR2_X1 U974 ( .A1(n868), .A2(n867), .ZN(n909) );
  XNOR2_X1 U975 ( .A(n909), .B(G162), .ZN(n893) );
  NAND2_X1 U976 ( .A1(G118), .A2(n869), .ZN(n872) );
  NAND2_X1 U977 ( .A1(G130), .A2(n870), .ZN(n871) );
  NAND2_X1 U978 ( .A1(n872), .A2(n871), .ZN(n880) );
  NAND2_X1 U979 ( .A1(G106), .A2(n873), .ZN(n876) );
  NAND2_X1 U980 ( .A1(G142), .A2(n518), .ZN(n875) );
  NAND2_X1 U981 ( .A1(n876), .A2(n875), .ZN(n877) );
  XOR2_X1 U982 ( .A(KEYINPUT110), .B(n877), .Z(n878) );
  XNOR2_X1 U983 ( .A(KEYINPUT45), .B(n878), .ZN(n879) );
  NOR2_X1 U984 ( .A1(n880), .A2(n879), .ZN(n884) );
  XOR2_X1 U985 ( .A(KEYINPUT111), .B(KEYINPUT112), .Z(n882) );
  XNOR2_X1 U986 ( .A(KEYINPUT48), .B(KEYINPUT46), .ZN(n881) );
  XNOR2_X1 U987 ( .A(n882), .B(n881), .ZN(n883) );
  XNOR2_X1 U988 ( .A(n884), .B(n883), .ZN(n887) );
  XNOR2_X1 U989 ( .A(G160), .B(n885), .ZN(n886) );
  XNOR2_X1 U990 ( .A(n887), .B(n886), .ZN(n888) );
  XNOR2_X1 U991 ( .A(n913), .B(n888), .ZN(n891) );
  XOR2_X1 U992 ( .A(G164), .B(n889), .Z(n890) );
  XNOR2_X1 U993 ( .A(n891), .B(n890), .ZN(n892) );
  XNOR2_X1 U994 ( .A(n893), .B(n892), .ZN(n895) );
  XOR2_X1 U995 ( .A(n895), .B(n894), .Z(n896) );
  NOR2_X1 U996 ( .A1(G37), .A2(n896), .ZN(G395) );
  XNOR2_X1 U997 ( .A(G286), .B(n973), .ZN(n900) );
  XNOR2_X1 U998 ( .A(n956), .B(G301), .ZN(n898) );
  XNOR2_X1 U999 ( .A(n898), .B(n897), .ZN(n899) );
  XNOR2_X1 U1000 ( .A(n900), .B(n899), .ZN(n901) );
  NOR2_X1 U1001 ( .A1(G37), .A2(n901), .ZN(G397) );
  OR2_X1 U1002 ( .A1(n908), .A2(G401), .ZN(n905) );
  NOR2_X1 U1003 ( .A1(G227), .A2(G229), .ZN(n902) );
  XOR2_X1 U1004 ( .A(KEYINPUT113), .B(n902), .Z(n903) );
  XNOR2_X1 U1005 ( .A(n903), .B(KEYINPUT49), .ZN(n904) );
  NOR2_X1 U1006 ( .A1(n905), .A2(n904), .ZN(n907) );
  NOR2_X1 U1007 ( .A1(G395), .A2(G397), .ZN(n906) );
  NAND2_X1 U1008 ( .A1(n907), .A2(n906), .ZN(G225) );
  INV_X1 U1009 ( .A(G225), .ZN(G308) );
  INV_X1 U1010 ( .A(n908), .ZN(G319) );
  XOR2_X1 U1011 ( .A(G2072), .B(n909), .Z(n911) );
  XOR2_X1 U1012 ( .A(G164), .B(G2078), .Z(n910) );
  NOR2_X1 U1013 ( .A1(n911), .A2(n910), .ZN(n912) );
  XOR2_X1 U1014 ( .A(KEYINPUT50), .B(n912), .Z(n931) );
  XNOR2_X1 U1015 ( .A(G160), .B(G2084), .ZN(n914) );
  NAND2_X1 U1016 ( .A1(n914), .A2(n913), .ZN(n915) );
  NOR2_X1 U1017 ( .A1(n916), .A2(n915), .ZN(n917) );
  NAND2_X1 U1018 ( .A1(n918), .A2(n917), .ZN(n924) );
  XOR2_X1 U1019 ( .A(G2090), .B(G162), .Z(n919) );
  NOR2_X1 U1020 ( .A1(n920), .A2(n919), .ZN(n921) );
  XOR2_X1 U1021 ( .A(KEYINPUT114), .B(n921), .Z(n922) );
  XOR2_X1 U1022 ( .A(KEYINPUT51), .B(n922), .Z(n923) );
  NOR2_X1 U1023 ( .A1(n924), .A2(n923), .ZN(n926) );
  NAND2_X1 U1024 ( .A1(n926), .A2(n925), .ZN(n927) );
  NOR2_X1 U1025 ( .A1(n928), .A2(n927), .ZN(n929) );
  XNOR2_X1 U1026 ( .A(KEYINPUT115), .B(n929), .ZN(n930) );
  NOR2_X1 U1027 ( .A1(n931), .A2(n930), .ZN(n932) );
  XNOR2_X1 U1028 ( .A(KEYINPUT52), .B(n932), .ZN(n934) );
  INV_X1 U1029 ( .A(KEYINPUT55), .ZN(n933) );
  NAND2_X1 U1030 ( .A1(n934), .A2(n933), .ZN(n935) );
  NAND2_X1 U1031 ( .A1(n935), .A2(G29), .ZN(n1024) );
  XOR2_X1 U1032 ( .A(G2090), .B(G35), .Z(n951) );
  XNOR2_X1 U1033 ( .A(G25), .B(n936), .ZN(n937) );
  NAND2_X1 U1034 ( .A1(n937), .A2(G28), .ZN(n947) );
  XNOR2_X1 U1035 ( .A(G2067), .B(G26), .ZN(n939) );
  XNOR2_X1 U1036 ( .A(G33), .B(G2072), .ZN(n938) );
  NOR2_X1 U1037 ( .A1(n939), .A2(n938), .ZN(n945) );
  XOR2_X1 U1038 ( .A(n940), .B(G32), .Z(n943) );
  XOR2_X1 U1039 ( .A(n941), .B(G27), .Z(n942) );
  NOR2_X1 U1040 ( .A1(n943), .A2(n942), .ZN(n944) );
  NAND2_X1 U1041 ( .A1(n945), .A2(n944), .ZN(n946) );
  NOR2_X1 U1042 ( .A1(n947), .A2(n946), .ZN(n948) );
  XOR2_X1 U1043 ( .A(KEYINPUT53), .B(n948), .Z(n949) );
  XNOR2_X1 U1044 ( .A(n949), .B(KEYINPUT116), .ZN(n950) );
  NAND2_X1 U1045 ( .A1(n951), .A2(n950), .ZN(n954) );
  XNOR2_X1 U1046 ( .A(KEYINPUT54), .B(G2084), .ZN(n952) );
  XNOR2_X1 U1047 ( .A(G34), .B(n952), .ZN(n953) );
  NOR2_X1 U1048 ( .A1(n954), .A2(n953), .ZN(n1016) );
  NAND2_X1 U1049 ( .A1(KEYINPUT55), .A2(n1016), .ZN(n955) );
  NAND2_X1 U1050 ( .A1(G11), .A2(n955), .ZN(n1022) );
  XNOR2_X1 U1051 ( .A(G16), .B(KEYINPUT56), .ZN(n983) );
  XOR2_X1 U1052 ( .A(G1348), .B(n956), .Z(n957) );
  NOR2_X1 U1053 ( .A1(n958), .A2(n957), .ZN(n981) );
  NAND2_X1 U1054 ( .A1(G303), .A2(G1971), .ZN(n966) );
  XNOR2_X1 U1055 ( .A(n959), .B(G1956), .ZN(n960) );
  XNOR2_X1 U1056 ( .A(n960), .B(KEYINPUT119), .ZN(n964) );
  NAND2_X1 U1057 ( .A1(n962), .A2(n961), .ZN(n963) );
  NOR2_X1 U1058 ( .A1(n964), .A2(n963), .ZN(n965) );
  NAND2_X1 U1059 ( .A1(n966), .A2(n965), .ZN(n967) );
  XNOR2_X1 U1060 ( .A(n967), .B(KEYINPUT120), .ZN(n979) );
  XOR2_X1 U1061 ( .A(G1966), .B(G168), .Z(n968) );
  XNOR2_X1 U1062 ( .A(KEYINPUT117), .B(n968), .ZN(n970) );
  NAND2_X1 U1063 ( .A1(n970), .A2(n969), .ZN(n972) );
  XNOR2_X1 U1064 ( .A(KEYINPUT118), .B(KEYINPUT57), .ZN(n971) );
  XNOR2_X1 U1065 ( .A(n972), .B(n971), .ZN(n977) );
  XNOR2_X1 U1066 ( .A(n973), .B(G1341), .ZN(n975) );
  XNOR2_X1 U1067 ( .A(G301), .B(G1961), .ZN(n974) );
  NOR2_X1 U1068 ( .A1(n975), .A2(n974), .ZN(n976) );
  NAND2_X1 U1069 ( .A1(n977), .A2(n976), .ZN(n978) );
  NOR2_X1 U1070 ( .A1(n979), .A2(n978), .ZN(n980) );
  NAND2_X1 U1071 ( .A1(n981), .A2(n980), .ZN(n982) );
  NAND2_X1 U1072 ( .A1(n983), .A2(n982), .ZN(n1014) );
  INV_X1 U1073 ( .A(G16), .ZN(n1012) );
  XOR2_X1 U1074 ( .A(G1966), .B(G21), .Z(n997) );
  XNOR2_X1 U1075 ( .A(KEYINPUT124), .B(KEYINPUT60), .ZN(n995) );
  XNOR2_X1 U1076 ( .A(KEYINPUT59), .B(G1348), .ZN(n984) );
  XNOR2_X1 U1077 ( .A(n984), .B(G4), .ZN(n989) );
  XOR2_X1 U1078 ( .A(G1981), .B(KEYINPUT123), .Z(n985) );
  XNOR2_X1 U1079 ( .A(G6), .B(n985), .ZN(n987) );
  XNOR2_X1 U1080 ( .A(G19), .B(G1341), .ZN(n986) );
  NOR2_X1 U1081 ( .A1(n987), .A2(n986), .ZN(n988) );
  NAND2_X1 U1082 ( .A1(n989), .A2(n988), .ZN(n993) );
  XOR2_X1 U1083 ( .A(G20), .B(n990), .Z(n991) );
  XNOR2_X1 U1084 ( .A(KEYINPUT122), .B(n991), .ZN(n992) );
  NOR2_X1 U1085 ( .A1(n993), .A2(n992), .ZN(n994) );
  XNOR2_X1 U1086 ( .A(n995), .B(n994), .ZN(n996) );
  NAND2_X1 U1087 ( .A1(n997), .A2(n996), .ZN(n998) );
  XNOR2_X1 U1088 ( .A(KEYINPUT125), .B(n998), .ZN(n1002) );
  XOR2_X1 U1089 ( .A(KEYINPUT121), .B(G5), .Z(n999) );
  XNOR2_X1 U1090 ( .A(n1000), .B(n999), .ZN(n1001) );
  NAND2_X1 U1091 ( .A1(n1002), .A2(n1001), .ZN(n1009) );
  XNOR2_X1 U1092 ( .A(G1971), .B(G22), .ZN(n1004) );
  XNOR2_X1 U1093 ( .A(G23), .B(G1976), .ZN(n1003) );
  NOR2_X1 U1094 ( .A1(n1004), .A2(n1003), .ZN(n1006) );
  XOR2_X1 U1095 ( .A(G1986), .B(G24), .Z(n1005) );
  NAND2_X1 U1096 ( .A1(n1006), .A2(n1005), .ZN(n1007) );
  XNOR2_X1 U1097 ( .A(KEYINPUT58), .B(n1007), .ZN(n1008) );
  NOR2_X1 U1098 ( .A1(n1009), .A2(n1008), .ZN(n1010) );
  XNOR2_X1 U1099 ( .A(KEYINPUT61), .B(n1010), .ZN(n1011) );
  NAND2_X1 U1100 ( .A1(n1012), .A2(n1011), .ZN(n1013) );
  NAND2_X1 U1101 ( .A1(n1014), .A2(n1013), .ZN(n1015) );
  XOR2_X1 U1102 ( .A(KEYINPUT126), .B(n1015), .Z(n1020) );
  INV_X1 U1103 ( .A(n1016), .ZN(n1018) );
  NOR2_X1 U1104 ( .A1(G29), .A2(KEYINPUT55), .ZN(n1017) );
  NAND2_X1 U1105 ( .A1(n1018), .A2(n1017), .ZN(n1019) );
  NAND2_X1 U1106 ( .A1(n1020), .A2(n1019), .ZN(n1021) );
  NOR2_X1 U1107 ( .A1(n1022), .A2(n1021), .ZN(n1023) );
  NAND2_X1 U1108 ( .A1(n1024), .A2(n1023), .ZN(n1025) );
  XOR2_X1 U1109 ( .A(KEYINPUT62), .B(n1025), .Z(G311) );
  INV_X1 U1110 ( .A(G311), .ZN(G150) );
endmodule

