//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 1 0 0 0 1 0 0 0 0 0 1 0 0 1 0 0 1 1 1 0 1 0 1 1 1 0 0 0 1 1 1 0 1 0 0 0 0 1 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 0 1 0 0 1 0 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:17:14 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n675, new_n676, new_n677, new_n678, new_n680,
    new_n681, new_n682, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n706, new_n707, new_n708, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n733, new_n734, new_n736,
    new_n737, new_n738, new_n740, new_n742, new_n743, new_n744, new_n745,
    new_n746, new_n747, new_n748, new_n749, new_n750, new_n751, new_n752,
    new_n753, new_n754, new_n755, new_n756, new_n757, new_n758, new_n759,
    new_n760, new_n761, new_n762, new_n763, new_n764, new_n765, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n785, new_n786, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n879, new_n880, new_n882, new_n883, new_n884,
    new_n885, new_n886, new_n887, new_n888, new_n889, new_n891, new_n892,
    new_n893, new_n894, new_n895, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n929, new_n930,
    new_n931, new_n933, new_n934, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n944, new_n945, new_n946, new_n948,
    new_n949, new_n950, new_n951, new_n952, new_n953, new_n954, new_n955,
    new_n956, new_n957, new_n958, new_n960, new_n961, new_n962, new_n963,
    new_n964, new_n965, new_n966, new_n967, new_n969, new_n970, new_n971,
    new_n972, new_n973, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n981, new_n982, new_n983, new_n984, new_n985, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993;
  INV_X1    g000(.A(KEYINPUT91), .ZN(new_n202));
  XOR2_X1   g001(.A(G43gat), .B(G50gat), .Z(new_n203));
  INV_X1    g002(.A(KEYINPUT15), .ZN(new_n204));
  INV_X1    g003(.A(G29gat), .ZN(new_n205));
  INV_X1    g004(.A(G36gat), .ZN(new_n206));
  OAI21_X1  g005(.A(KEYINPUT14), .B1(new_n205), .B2(new_n206), .ZN(new_n207));
  NAND2_X1  g006(.A1(new_n205), .A2(new_n206), .ZN(new_n208));
  AND2_X1   g007(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  AND3_X1   g008(.A1(new_n205), .A2(new_n206), .A3(KEYINPUT14), .ZN(new_n210));
  OAI21_X1  g009(.A(new_n204), .B1(new_n209), .B2(new_n210), .ZN(new_n211));
  AOI21_X1  g010(.A(new_n210), .B1(new_n208), .B2(new_n207), .ZN(new_n212));
  NAND2_X1  g011(.A1(new_n212), .A2(KEYINPUT15), .ZN(new_n213));
  AOI21_X1  g012(.A(new_n203), .B1(new_n211), .B2(new_n213), .ZN(new_n214));
  AND2_X1   g013(.A1(new_n213), .A2(new_n203), .ZN(new_n215));
  NOR2_X1   g014(.A1(new_n214), .A2(new_n215), .ZN(new_n216));
  INV_X1    g015(.A(KEYINPUT88), .ZN(new_n217));
  NAND2_X1  g016(.A1(new_n216), .A2(new_n217), .ZN(new_n218));
  OAI21_X1  g017(.A(KEYINPUT88), .B1(new_n214), .B2(new_n215), .ZN(new_n219));
  NAND2_X1  g018(.A1(new_n218), .A2(new_n219), .ZN(new_n220));
  XOR2_X1   g019(.A(G15gat), .B(G22gat), .Z(new_n221));
  INV_X1    g020(.A(G1gat), .ZN(new_n222));
  NAND2_X1  g021(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  INV_X1    g022(.A(KEYINPUT89), .ZN(new_n224));
  NAND2_X1  g023(.A1(new_n223), .A2(new_n224), .ZN(new_n225));
  XNOR2_X1  g024(.A(G15gat), .B(G22gat), .ZN(new_n226));
  INV_X1    g025(.A(KEYINPUT16), .ZN(new_n227));
  OAI21_X1  g026(.A(new_n226), .B1(new_n227), .B2(G1gat), .ZN(new_n228));
  NAND2_X1  g027(.A1(new_n223), .A2(new_n228), .ZN(new_n229));
  NAND3_X1  g028(.A1(new_n225), .A2(new_n229), .A3(G8gat), .ZN(new_n230));
  INV_X1    g029(.A(G8gat), .ZN(new_n231));
  OAI211_X1 g030(.A(new_n223), .B(new_n228), .C1(new_n224), .C2(new_n231), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n230), .A2(new_n232), .ZN(new_n233));
  INV_X1    g032(.A(KEYINPUT90), .ZN(new_n234));
  XNOR2_X1  g033(.A(new_n233), .B(new_n234), .ZN(new_n235));
  OAI21_X1  g034(.A(new_n202), .B1(new_n220), .B2(new_n235), .ZN(new_n236));
  XNOR2_X1  g035(.A(new_n233), .B(KEYINPUT90), .ZN(new_n237));
  NAND4_X1  g036(.A1(new_n237), .A2(KEYINPUT91), .A3(new_n219), .A4(new_n218), .ZN(new_n238));
  NAND2_X1  g037(.A1(new_n236), .A2(new_n238), .ZN(new_n239));
  NAND2_X1  g038(.A1(G229gat), .A2(G233gat), .ZN(new_n240));
  INV_X1    g039(.A(new_n233), .ZN(new_n241));
  OAI21_X1  g040(.A(KEYINPUT17), .B1(new_n214), .B2(new_n215), .ZN(new_n242));
  OAI211_X1 g041(.A(new_n241), .B(new_n242), .C1(new_n220), .C2(KEYINPUT17), .ZN(new_n243));
  NAND3_X1  g042(.A1(new_n239), .A2(new_n240), .A3(new_n243), .ZN(new_n244));
  INV_X1    g043(.A(KEYINPUT18), .ZN(new_n245));
  NAND2_X1  g044(.A1(new_n244), .A2(new_n245), .ZN(new_n246));
  NAND2_X1  g045(.A1(new_n220), .A2(new_n235), .ZN(new_n247));
  NAND2_X1  g046(.A1(new_n239), .A2(new_n247), .ZN(new_n248));
  XNOR2_X1  g047(.A(new_n240), .B(KEYINPUT13), .ZN(new_n249));
  INV_X1    g048(.A(new_n249), .ZN(new_n250));
  NAND2_X1  g049(.A1(new_n248), .A2(new_n250), .ZN(new_n251));
  NAND4_X1  g050(.A1(new_n239), .A2(KEYINPUT18), .A3(new_n240), .A4(new_n243), .ZN(new_n252));
  NAND3_X1  g051(.A1(new_n246), .A2(new_n251), .A3(new_n252), .ZN(new_n253));
  XNOR2_X1  g052(.A(G113gat), .B(G141gat), .ZN(new_n254));
  XNOR2_X1  g053(.A(new_n254), .B(G197gat), .ZN(new_n255));
  XNOR2_X1  g054(.A(new_n255), .B(KEYINPUT11), .ZN(new_n256));
  INV_X1    g055(.A(G169gat), .ZN(new_n257));
  XNOR2_X1  g056(.A(new_n256), .B(new_n257), .ZN(new_n258));
  XNOR2_X1  g057(.A(new_n258), .B(KEYINPUT12), .ZN(new_n259));
  INV_X1    g058(.A(new_n259), .ZN(new_n260));
  NAND2_X1  g059(.A1(new_n253), .A2(new_n260), .ZN(new_n261));
  NAND4_X1  g060(.A1(new_n246), .A2(new_n251), .A3(new_n259), .A4(new_n252), .ZN(new_n262));
  NAND2_X1  g061(.A1(new_n261), .A2(new_n262), .ZN(new_n263));
  INV_X1    g062(.A(new_n263), .ZN(new_n264));
  NAND2_X1  g063(.A1(G230gat), .A2(G233gat), .ZN(new_n265));
  INV_X1    g064(.A(KEYINPUT92), .ZN(new_n266));
  NAND2_X1  g065(.A1(new_n266), .A2(G57gat), .ZN(new_n267));
  XNOR2_X1  g066(.A(new_n267), .B(G64gat), .ZN(new_n268));
  XNOR2_X1  g067(.A(G71gat), .B(G78gat), .ZN(new_n269));
  AND2_X1   g068(.A1(G71gat), .A2(G78gat), .ZN(new_n270));
  OAI211_X1 g069(.A(new_n268), .B(new_n269), .C1(KEYINPUT9), .C2(new_n270), .ZN(new_n271));
  OR2_X1    g070(.A1(G57gat), .A2(G64gat), .ZN(new_n272));
  NAND2_X1  g071(.A1(G57gat), .A2(G64gat), .ZN(new_n273));
  AND3_X1   g072(.A1(new_n272), .A2(KEYINPUT9), .A3(new_n273), .ZN(new_n274));
  OR2_X1    g073(.A1(new_n274), .A2(new_n269), .ZN(new_n275));
  NAND2_X1  g074(.A1(new_n271), .A2(new_n275), .ZN(new_n276));
  NAND2_X1  g075(.A1(G85gat), .A2(G92gat), .ZN(new_n277));
  XNOR2_X1  g076(.A(new_n277), .B(KEYINPUT7), .ZN(new_n278));
  NAND2_X1  g077(.A1(G99gat), .A2(G106gat), .ZN(new_n279));
  INV_X1    g078(.A(G85gat), .ZN(new_n280));
  INV_X1    g079(.A(G92gat), .ZN(new_n281));
  AOI22_X1  g080(.A1(KEYINPUT8), .A2(new_n279), .B1(new_n280), .B2(new_n281), .ZN(new_n282));
  NAND2_X1  g081(.A1(new_n278), .A2(new_n282), .ZN(new_n283));
  INV_X1    g082(.A(new_n283), .ZN(new_n284));
  NOR2_X1   g083(.A1(new_n284), .A2(KEYINPUT95), .ZN(new_n285));
  NOR2_X1   g084(.A1(new_n276), .A2(new_n285), .ZN(new_n286));
  XOR2_X1   g085(.A(G99gat), .B(G106gat), .Z(new_n287));
  XNOR2_X1  g086(.A(new_n283), .B(new_n287), .ZN(new_n288));
  NAND2_X1  g087(.A1(new_n286), .A2(new_n288), .ZN(new_n289));
  NOR2_X1   g088(.A1(new_n284), .A2(new_n287), .ZN(new_n290));
  AND2_X1   g089(.A1(new_n284), .A2(new_n287), .ZN(new_n291));
  OAI22_X1  g090(.A1(new_n290), .A2(new_n291), .B1(new_n276), .B2(new_n285), .ZN(new_n292));
  AOI21_X1  g091(.A(KEYINPUT10), .B1(new_n289), .B2(new_n292), .ZN(new_n293));
  INV_X1    g092(.A(new_n288), .ZN(new_n294));
  INV_X1    g093(.A(new_n276), .ZN(new_n295));
  NAND3_X1  g094(.A1(new_n294), .A2(KEYINPUT10), .A3(new_n295), .ZN(new_n296));
  INV_X1    g095(.A(new_n296), .ZN(new_n297));
  OAI21_X1  g096(.A(new_n265), .B1(new_n293), .B2(new_n297), .ZN(new_n298));
  NAND2_X1  g097(.A1(new_n298), .A2(KEYINPUT97), .ZN(new_n299));
  INV_X1    g098(.A(new_n265), .ZN(new_n300));
  NAND3_X1  g099(.A1(new_n289), .A2(new_n300), .A3(new_n292), .ZN(new_n301));
  INV_X1    g100(.A(KEYINPUT97), .ZN(new_n302));
  OAI211_X1 g101(.A(new_n302), .B(new_n265), .C1(new_n293), .C2(new_n297), .ZN(new_n303));
  NAND3_X1  g102(.A1(new_n299), .A2(new_n301), .A3(new_n303), .ZN(new_n304));
  XNOR2_X1  g103(.A(G120gat), .B(G148gat), .ZN(new_n305));
  INV_X1    g104(.A(G176gat), .ZN(new_n306));
  XNOR2_X1  g105(.A(new_n305), .B(new_n306), .ZN(new_n307));
  XOR2_X1   g106(.A(new_n307), .B(G204gat), .Z(new_n308));
  NAND2_X1  g107(.A1(new_n304), .A2(new_n308), .ZN(new_n309));
  INV_X1    g108(.A(KEYINPUT96), .ZN(new_n310));
  NAND2_X1  g109(.A1(new_n289), .A2(new_n292), .ZN(new_n311));
  INV_X1    g110(.A(KEYINPUT10), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n311), .A2(new_n312), .ZN(new_n313));
  AOI21_X1  g112(.A(new_n310), .B1(new_n313), .B2(new_n296), .ZN(new_n314));
  NOR3_X1   g113(.A1(new_n293), .A2(KEYINPUT96), .A3(new_n297), .ZN(new_n315));
  OAI21_X1  g114(.A(new_n265), .B1(new_n314), .B2(new_n315), .ZN(new_n316));
  INV_X1    g115(.A(new_n308), .ZN(new_n317));
  NAND3_X1  g116(.A1(new_n316), .A2(new_n301), .A3(new_n317), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n309), .A2(new_n318), .ZN(new_n319));
  NAND2_X1  g118(.A1(new_n319), .A2(KEYINPUT98), .ZN(new_n320));
  INV_X1    g119(.A(KEYINPUT98), .ZN(new_n321));
  NAND3_X1  g120(.A1(new_n309), .A2(new_n318), .A3(new_n321), .ZN(new_n322));
  NAND2_X1  g121(.A1(new_n320), .A2(new_n322), .ZN(new_n323));
  NOR2_X1   g122(.A1(new_n264), .A2(new_n323), .ZN(new_n324));
  INV_X1    g123(.A(KEYINPUT72), .ZN(new_n325));
  NAND2_X1  g124(.A1(G226gat), .A2(G233gat), .ZN(new_n326));
  INV_X1    g125(.A(new_n326), .ZN(new_n327));
  INV_X1    g126(.A(KEYINPUT26), .ZN(new_n328));
  NAND3_X1  g127(.A1(new_n328), .A2(new_n257), .A3(new_n306), .ZN(new_n329));
  NAND2_X1  g128(.A1(G169gat), .A2(G176gat), .ZN(new_n330));
  OAI21_X1  g129(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n331));
  NAND3_X1  g130(.A1(new_n329), .A2(new_n330), .A3(new_n331), .ZN(new_n332));
  INV_X1    g131(.A(KEYINPUT28), .ZN(new_n333));
  INV_X1    g132(.A(G190gat), .ZN(new_n334));
  AND2_X1   g133(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n335));
  NOR2_X1   g134(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n336));
  OAI211_X1 g135(.A(new_n333), .B(new_n334), .C1(new_n335), .C2(new_n336), .ZN(new_n337));
  NAND2_X1  g136(.A1(G183gat), .A2(G190gat), .ZN(new_n338));
  AND3_X1   g137(.A1(new_n332), .A2(new_n337), .A3(new_n338), .ZN(new_n339));
  OR2_X1    g138(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n340));
  INV_X1    g139(.A(KEYINPUT66), .ZN(new_n341));
  NAND2_X1  g140(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n342));
  NAND3_X1  g141(.A1(new_n340), .A2(new_n341), .A3(new_n342), .ZN(new_n343));
  OAI21_X1  g142(.A(KEYINPUT66), .B1(new_n335), .B2(new_n336), .ZN(new_n344));
  AOI21_X1  g143(.A(G190gat), .B1(new_n343), .B2(new_n344), .ZN(new_n345));
  OAI21_X1  g144(.A(new_n339), .B1(new_n333), .B2(new_n345), .ZN(new_n346));
  INV_X1    g145(.A(KEYINPUT24), .ZN(new_n347));
  NAND3_X1  g146(.A1(new_n347), .A2(G183gat), .A3(G190gat), .ZN(new_n348));
  NAND2_X1  g147(.A1(new_n338), .A2(KEYINPUT24), .ZN(new_n349));
  NOR2_X1   g148(.A1(G183gat), .A2(G190gat), .ZN(new_n350));
  OAI21_X1  g149(.A(new_n348), .B1(new_n349), .B2(new_n350), .ZN(new_n351));
  INV_X1    g150(.A(new_n351), .ZN(new_n352));
  INV_X1    g151(.A(KEYINPUT23), .ZN(new_n353));
  OAI21_X1  g152(.A(new_n353), .B1(G169gat), .B2(G176gat), .ZN(new_n354));
  AOI21_X1  g153(.A(KEYINPUT25), .B1(G169gat), .B2(G176gat), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n354), .A2(new_n355), .ZN(new_n356));
  INV_X1    g155(.A(KEYINPUT64), .ZN(new_n357));
  AND4_X1   g156(.A1(new_n357), .A2(new_n257), .A3(new_n306), .A4(KEYINPUT23), .ZN(new_n358));
  NOR2_X1   g157(.A1(G169gat), .A2(G176gat), .ZN(new_n359));
  AOI21_X1  g158(.A(new_n357), .B1(new_n359), .B2(KEYINPUT23), .ZN(new_n360));
  NOR3_X1   g159(.A1(new_n356), .A2(new_n358), .A3(new_n360), .ZN(new_n361));
  INV_X1    g160(.A(KEYINPUT65), .ZN(new_n362));
  INV_X1    g161(.A(KEYINPUT25), .ZN(new_n363));
  NOR2_X1   g162(.A1(new_n362), .A2(new_n363), .ZN(new_n364));
  OAI21_X1  g163(.A(new_n352), .B1(new_n361), .B2(new_n364), .ZN(new_n365));
  INV_X1    g164(.A(new_n350), .ZN(new_n366));
  NAND3_X1  g165(.A1(new_n366), .A2(KEYINPUT24), .A3(new_n338), .ZN(new_n367));
  AOI21_X1  g166(.A(KEYINPUT65), .B1(new_n367), .B2(new_n348), .ZN(new_n368));
  NAND3_X1  g167(.A1(new_n257), .A2(new_n306), .A3(KEYINPUT23), .ZN(new_n369));
  NAND3_X1  g168(.A1(new_n369), .A2(new_n354), .A3(new_n330), .ZN(new_n370));
  OAI21_X1  g169(.A(KEYINPUT25), .B1(new_n368), .B2(new_n370), .ZN(new_n371));
  NAND3_X1  g170(.A1(new_n346), .A2(new_n365), .A3(new_n371), .ZN(new_n372));
  INV_X1    g171(.A(KEYINPUT29), .ZN(new_n373));
  AOI21_X1  g172(.A(new_n327), .B1(new_n372), .B2(new_n373), .ZN(new_n374));
  AND2_X1   g173(.A1(new_n354), .A2(new_n355), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n369), .A2(KEYINPUT64), .ZN(new_n376));
  NAND3_X1  g175(.A1(new_n359), .A2(new_n357), .A3(KEYINPUT23), .ZN(new_n377));
  NAND3_X1  g176(.A1(new_n375), .A2(new_n376), .A3(new_n377), .ZN(new_n378));
  INV_X1    g177(.A(new_n364), .ZN(new_n379));
  AOI21_X1  g178(.A(new_n351), .B1(new_n378), .B2(new_n379), .ZN(new_n380));
  NAND2_X1  g179(.A1(new_n351), .A2(new_n362), .ZN(new_n381));
  INV_X1    g180(.A(new_n370), .ZN(new_n382));
  AOI21_X1  g181(.A(new_n363), .B1(new_n381), .B2(new_n382), .ZN(new_n383));
  NOR2_X1   g182(.A1(new_n380), .A2(new_n383), .ZN(new_n384));
  AOI21_X1  g183(.A(new_n326), .B1(new_n384), .B2(new_n346), .ZN(new_n385));
  OAI21_X1  g184(.A(new_n325), .B1(new_n374), .B2(new_n385), .ZN(new_n386));
  XNOR2_X1  g185(.A(G197gat), .B(G204gat), .ZN(new_n387));
  INV_X1    g186(.A(KEYINPUT22), .ZN(new_n388));
  INV_X1    g187(.A(G211gat), .ZN(new_n389));
  INV_X1    g188(.A(G218gat), .ZN(new_n390));
  OAI21_X1  g189(.A(new_n388), .B1(new_n389), .B2(new_n390), .ZN(new_n391));
  NAND2_X1  g190(.A1(new_n387), .A2(new_n391), .ZN(new_n392));
  XNOR2_X1  g191(.A(G211gat), .B(G218gat), .ZN(new_n393));
  INV_X1    g192(.A(new_n393), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n392), .A2(new_n394), .ZN(new_n395));
  NAND3_X1  g194(.A1(new_n393), .A2(new_n387), .A3(new_n391), .ZN(new_n396));
  NAND2_X1  g195(.A1(new_n395), .A2(new_n396), .ZN(new_n397));
  AOI21_X1  g196(.A(KEYINPUT29), .B1(new_n384), .B2(new_n346), .ZN(new_n398));
  OAI21_X1  g197(.A(KEYINPUT72), .B1(new_n398), .B2(new_n327), .ZN(new_n399));
  NAND3_X1  g198(.A1(new_n386), .A2(new_n397), .A3(new_n399), .ZN(new_n400));
  INV_X1    g199(.A(new_n397), .ZN(new_n401));
  OAI21_X1  g200(.A(new_n401), .B1(new_n374), .B2(new_n385), .ZN(new_n402));
  NAND2_X1  g201(.A1(new_n402), .A2(KEYINPUT71), .ZN(new_n403));
  INV_X1    g202(.A(KEYINPUT71), .ZN(new_n404));
  OAI211_X1 g203(.A(new_n404), .B(new_n401), .C1(new_n374), .C2(new_n385), .ZN(new_n405));
  XNOR2_X1  g204(.A(G8gat), .B(G36gat), .ZN(new_n406));
  XNOR2_X1  g205(.A(new_n406), .B(KEYINPUT73), .ZN(new_n407));
  XOR2_X1   g206(.A(new_n407), .B(G64gat), .Z(new_n408));
  XNOR2_X1  g207(.A(new_n408), .B(new_n281), .ZN(new_n409));
  NAND4_X1  g208(.A1(new_n400), .A2(new_n403), .A3(new_n405), .A4(new_n409), .ZN(new_n410));
  INV_X1    g209(.A(new_n410), .ZN(new_n411));
  NAND2_X1  g210(.A1(G225gat), .A2(G233gat), .ZN(new_n412));
  AND2_X1   g211(.A1(G155gat), .A2(G162gat), .ZN(new_n413));
  INV_X1    g212(.A(KEYINPUT2), .ZN(new_n414));
  NOR2_X1   g213(.A1(G155gat), .A2(G162gat), .ZN(new_n415));
  AOI21_X1  g214(.A(new_n413), .B1(new_n414), .B2(new_n415), .ZN(new_n416));
  INV_X1    g215(.A(KEYINPUT76), .ZN(new_n417));
  NOR2_X1   g216(.A1(new_n417), .A2(G148gat), .ZN(new_n418));
  INV_X1    g217(.A(G148gat), .ZN(new_n419));
  NOR2_X1   g218(.A1(new_n419), .A2(KEYINPUT76), .ZN(new_n420));
  OAI21_X1  g219(.A(G141gat), .B1(new_n418), .B2(new_n420), .ZN(new_n421));
  INV_X1    g220(.A(G141gat), .ZN(new_n422));
  NAND2_X1  g221(.A1(new_n422), .A2(G148gat), .ZN(new_n423));
  AOI21_X1  g222(.A(new_n416), .B1(new_n421), .B2(new_n423), .ZN(new_n424));
  XNOR2_X1  g223(.A(G155gat), .B(G162gat), .ZN(new_n425));
  NAND2_X1  g224(.A1(new_n419), .A2(G141gat), .ZN(new_n426));
  NAND2_X1  g225(.A1(new_n423), .A2(new_n426), .ZN(new_n427));
  XNOR2_X1  g226(.A(KEYINPUT75), .B(KEYINPUT2), .ZN(new_n428));
  AOI21_X1  g227(.A(new_n425), .B1(new_n427), .B2(new_n428), .ZN(new_n429));
  OAI21_X1  g228(.A(KEYINPUT3), .B1(new_n424), .B2(new_n429), .ZN(new_n430));
  NOR2_X1   g229(.A1(new_n413), .A2(new_n415), .ZN(new_n431));
  AND2_X1   g230(.A1(KEYINPUT75), .A2(KEYINPUT2), .ZN(new_n432));
  NOR2_X1   g231(.A1(KEYINPUT75), .A2(KEYINPUT2), .ZN(new_n433));
  NOR2_X1   g232(.A1(new_n432), .A2(new_n433), .ZN(new_n434));
  XNOR2_X1  g233(.A(G141gat), .B(G148gat), .ZN(new_n435));
  OAI21_X1  g234(.A(new_n431), .B1(new_n434), .B2(new_n435), .ZN(new_n436));
  INV_X1    g235(.A(KEYINPUT3), .ZN(new_n437));
  INV_X1    g236(.A(new_n423), .ZN(new_n438));
  NAND2_X1  g237(.A1(new_n419), .A2(KEYINPUT76), .ZN(new_n439));
  NAND2_X1  g238(.A1(new_n417), .A2(G148gat), .ZN(new_n440));
  NAND2_X1  g239(.A1(new_n439), .A2(new_n440), .ZN(new_n441));
  AOI21_X1  g240(.A(new_n438), .B1(new_n441), .B2(G141gat), .ZN(new_n442));
  OAI211_X1 g241(.A(new_n436), .B(new_n437), .C1(new_n442), .C2(new_n416), .ZN(new_n443));
  INV_X1    g242(.A(G113gat), .ZN(new_n444));
  INV_X1    g243(.A(G120gat), .ZN(new_n445));
  AOI21_X1  g244(.A(KEYINPUT1), .B1(new_n444), .B2(new_n445), .ZN(new_n446));
  NAND2_X1  g245(.A1(G113gat), .A2(G120gat), .ZN(new_n447));
  NAND2_X1  g246(.A1(new_n446), .A2(new_n447), .ZN(new_n448));
  OR2_X1    g247(.A1(G127gat), .A2(G134gat), .ZN(new_n449));
  OR2_X1    g248(.A1(KEYINPUT67), .A2(G127gat), .ZN(new_n450));
  NAND2_X1  g249(.A1(KEYINPUT67), .A2(G127gat), .ZN(new_n451));
  NAND3_X1  g250(.A1(new_n450), .A2(G134gat), .A3(new_n451), .ZN(new_n452));
  NAND3_X1  g251(.A1(new_n448), .A2(new_n449), .A3(new_n452), .ZN(new_n453));
  XNOR2_X1  g252(.A(G127gat), .B(G134gat), .ZN(new_n454));
  XNOR2_X1  g253(.A(KEYINPUT68), .B(G113gat), .ZN(new_n455));
  OAI211_X1 g254(.A(new_n446), .B(new_n454), .C1(new_n455), .C2(new_n445), .ZN(new_n456));
  NAND2_X1  g255(.A1(new_n453), .A2(new_n456), .ZN(new_n457));
  NAND3_X1  g256(.A1(new_n430), .A2(new_n443), .A3(new_n457), .ZN(new_n458));
  INV_X1    g257(.A(KEYINPUT4), .ZN(new_n459));
  AND2_X1   g258(.A1(new_n453), .A2(new_n456), .ZN(new_n460));
  XNOR2_X1  g259(.A(KEYINPUT76), .B(G148gat), .ZN(new_n461));
  OAI21_X1  g260(.A(new_n423), .B1(new_n461), .B2(new_n422), .ZN(new_n462));
  INV_X1    g261(.A(new_n416), .ZN(new_n463));
  NAND2_X1  g262(.A1(new_n427), .A2(new_n428), .ZN(new_n464));
  AOI22_X1  g263(.A1(new_n462), .A2(new_n463), .B1(new_n464), .B2(new_n431), .ZN(new_n465));
  AOI21_X1  g264(.A(new_n459), .B1(new_n460), .B2(new_n465), .ZN(new_n466));
  OAI21_X1  g265(.A(new_n436), .B1(new_n442), .B2(new_n416), .ZN(new_n467));
  NOR3_X1   g266(.A1(new_n467), .A2(new_n457), .A3(KEYINPUT4), .ZN(new_n468));
  OAI211_X1 g267(.A(new_n412), .B(new_n458), .C1(new_n466), .C2(new_n468), .ZN(new_n469));
  XNOR2_X1  g268(.A(new_n467), .B(new_n457), .ZN(new_n470));
  INV_X1    g269(.A(new_n412), .ZN(new_n471));
  NAND2_X1  g270(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  NAND2_X1  g271(.A1(new_n469), .A2(new_n472), .ZN(new_n473));
  NAND2_X1  g272(.A1(new_n473), .A2(KEYINPUT5), .ZN(new_n474));
  XNOR2_X1  g273(.A(G1gat), .B(G29gat), .ZN(new_n475));
  XNOR2_X1  g274(.A(new_n475), .B(KEYINPUT0), .ZN(new_n476));
  XNOR2_X1  g275(.A(new_n476), .B(G57gat), .ZN(new_n477));
  XNOR2_X1  g276(.A(new_n477), .B(new_n280), .ZN(new_n478));
  INV_X1    g277(.A(new_n478), .ZN(new_n479));
  INV_X1    g278(.A(KEYINPUT5), .ZN(new_n480));
  NAND2_X1  g279(.A1(new_n469), .A2(new_n480), .ZN(new_n481));
  NAND3_X1  g280(.A1(new_n474), .A2(new_n479), .A3(new_n481), .ZN(new_n482));
  AOI21_X1  g281(.A(new_n479), .B1(new_n474), .B2(new_n481), .ZN(new_n483));
  OAI21_X1  g282(.A(new_n482), .B1(new_n483), .B2(KEYINPUT6), .ZN(new_n484));
  AOI21_X1  g283(.A(new_n480), .B1(new_n469), .B2(new_n472), .ZN(new_n485));
  AND2_X1   g284(.A1(new_n443), .A2(new_n457), .ZN(new_n486));
  NAND3_X1  g285(.A1(new_n460), .A2(new_n465), .A3(new_n459), .ZN(new_n487));
  OAI21_X1  g286(.A(KEYINPUT4), .B1(new_n467), .B2(new_n457), .ZN(new_n488));
  AOI22_X1  g287(.A1(new_n430), .A2(new_n486), .B1(new_n487), .B2(new_n488), .ZN(new_n489));
  AOI21_X1  g288(.A(KEYINPUT5), .B1(new_n489), .B2(new_n412), .ZN(new_n490));
  NOR3_X1   g289(.A1(new_n485), .A2(new_n490), .A3(new_n478), .ZN(new_n491));
  INV_X1    g290(.A(KEYINPUT6), .ZN(new_n492));
  NAND2_X1  g291(.A1(new_n491), .A2(new_n492), .ZN(new_n493));
  AOI21_X1  g292(.A(new_n411), .B1(new_n484), .B2(new_n493), .ZN(new_n494));
  INV_X1    g293(.A(KEYINPUT37), .ZN(new_n495));
  NAND4_X1  g294(.A1(new_n400), .A2(new_n403), .A3(new_n495), .A4(new_n405), .ZN(new_n496));
  INV_X1    g295(.A(KEYINPUT84), .ZN(new_n497));
  XNOR2_X1  g296(.A(new_n496), .B(new_n497), .ZN(new_n498));
  NOR2_X1   g297(.A1(new_n409), .A2(KEYINPUT38), .ZN(new_n499));
  NAND3_X1  g298(.A1(new_n386), .A2(new_n401), .A3(new_n399), .ZN(new_n500));
  NAND2_X1  g299(.A1(new_n372), .A2(new_n327), .ZN(new_n501));
  OAI21_X1  g300(.A(new_n501), .B1(new_n398), .B2(new_n327), .ZN(new_n502));
  AOI21_X1  g301(.A(new_n495), .B1(new_n502), .B2(new_n397), .ZN(new_n503));
  INV_X1    g302(.A(KEYINPUT83), .ZN(new_n504));
  AND3_X1   g303(.A1(new_n500), .A2(new_n503), .A3(new_n504), .ZN(new_n505));
  AOI21_X1  g304(.A(new_n504), .B1(new_n500), .B2(new_n503), .ZN(new_n506));
  OAI21_X1  g305(.A(new_n499), .B1(new_n505), .B2(new_n506), .ZN(new_n507));
  OAI21_X1  g306(.A(new_n494), .B1(new_n498), .B2(new_n507), .ZN(new_n508));
  INV_X1    g307(.A(KEYINPUT85), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  XNOR2_X1  g309(.A(new_n496), .B(KEYINPUT84), .ZN(new_n511));
  INV_X1    g310(.A(new_n409), .ZN(new_n512));
  NAND3_X1  g311(.A1(new_n400), .A2(new_n403), .A3(new_n405), .ZN(new_n513));
  NAND2_X1  g312(.A1(new_n513), .A2(KEYINPUT37), .ZN(new_n514));
  NAND3_X1  g313(.A1(new_n511), .A2(new_n512), .A3(new_n514), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n515), .A2(KEYINPUT38), .ZN(new_n516));
  OAI211_X1 g315(.A(KEYINPUT85), .B(new_n494), .C1(new_n498), .C2(new_n507), .ZN(new_n517));
  NAND3_X1  g316(.A1(new_n510), .A2(new_n516), .A3(new_n517), .ZN(new_n518));
  AOI21_X1  g317(.A(KEYINPUT29), .B1(new_n395), .B2(new_n396), .ZN(new_n519));
  OAI21_X1  g318(.A(new_n467), .B1(new_n519), .B2(KEYINPUT3), .ZN(new_n520));
  AOI21_X1  g319(.A(KEYINPUT29), .B1(new_n465), .B2(new_n437), .ZN(new_n521));
  OAI21_X1  g320(.A(new_n520), .B1(new_n521), .B2(new_n397), .ZN(new_n522));
  NAND2_X1  g321(.A1(G228gat), .A2(G233gat), .ZN(new_n523));
  XNOR2_X1  g322(.A(new_n523), .B(G22gat), .ZN(new_n524));
  INV_X1    g323(.A(new_n524), .ZN(new_n525));
  NAND2_X1  g324(.A1(new_n522), .A2(new_n525), .ZN(new_n526));
  OAI211_X1 g325(.A(new_n520), .B(new_n524), .C1(new_n521), .C2(new_n397), .ZN(new_n527));
  NAND3_X1  g326(.A1(new_n526), .A2(new_n527), .A3(KEYINPUT79), .ZN(new_n528));
  XNOR2_X1  g327(.A(G78gat), .B(G106gat), .ZN(new_n529));
  INV_X1    g328(.A(G50gat), .ZN(new_n530));
  XNOR2_X1  g329(.A(new_n529), .B(new_n530), .ZN(new_n531));
  XNOR2_X1  g330(.A(KEYINPUT78), .B(KEYINPUT31), .ZN(new_n532));
  XNOR2_X1  g331(.A(new_n531), .B(new_n532), .ZN(new_n533));
  XNOR2_X1  g332(.A(new_n528), .B(new_n533), .ZN(new_n534));
  INV_X1    g333(.A(new_n534), .ZN(new_n535));
  INV_X1    g334(.A(KEYINPUT39), .ZN(new_n536));
  OR2_X1    g335(.A1(new_n470), .A2(new_n471), .ZN(new_n537));
  AOI21_X1  g336(.A(new_n536), .B1(new_n537), .B2(KEYINPUT81), .ZN(new_n538));
  OAI221_X1 g337(.A(new_n538), .B1(KEYINPUT81), .B2(new_n537), .C1(new_n412), .C2(new_n489), .ZN(new_n539));
  XOR2_X1   g338(.A(KEYINPUT80), .B(KEYINPUT39), .Z(new_n540));
  OR3_X1    g339(.A1(new_n489), .A2(new_n412), .A3(new_n540), .ZN(new_n541));
  NAND3_X1  g340(.A1(new_n539), .A2(new_n478), .A3(new_n541), .ZN(new_n542));
  INV_X1    g341(.A(KEYINPUT40), .ZN(new_n543));
  NAND3_X1  g342(.A1(new_n542), .A2(KEYINPUT82), .A3(new_n543), .ZN(new_n544));
  NAND2_X1  g343(.A1(new_n543), .A2(KEYINPUT82), .ZN(new_n545));
  NAND4_X1  g344(.A1(new_n539), .A2(new_n478), .A3(new_n545), .A4(new_n541), .ZN(new_n546));
  AND3_X1   g345(.A1(new_n544), .A2(new_n482), .A3(new_n546), .ZN(new_n547));
  NAND2_X1  g346(.A1(new_n513), .A2(new_n512), .ZN(new_n548));
  INV_X1    g347(.A(KEYINPUT74), .ZN(new_n549));
  NAND2_X1  g348(.A1(new_n548), .A2(new_n549), .ZN(new_n550));
  NAND3_X1  g349(.A1(new_n513), .A2(KEYINPUT74), .A3(new_n512), .ZN(new_n551));
  NAND2_X1  g350(.A1(new_n410), .A2(KEYINPUT30), .ZN(new_n552));
  AOI21_X1  g351(.A(new_n404), .B1(new_n502), .B2(new_n401), .ZN(new_n553));
  INV_X1    g352(.A(new_n405), .ZN(new_n554));
  NOR2_X1   g353(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  INV_X1    g354(.A(KEYINPUT30), .ZN(new_n556));
  NAND4_X1  g355(.A1(new_n555), .A2(new_n556), .A3(new_n400), .A4(new_n409), .ZN(new_n557));
  AOI22_X1  g356(.A1(new_n550), .A2(new_n551), .B1(new_n552), .B2(new_n557), .ZN(new_n558));
  INV_X1    g357(.A(new_n558), .ZN(new_n559));
  AOI21_X1  g358(.A(new_n535), .B1(new_n547), .B2(new_n559), .ZN(new_n560));
  NAND2_X1  g359(.A1(new_n518), .A2(new_n560), .ZN(new_n561));
  INV_X1    g360(.A(new_n493), .ZN(new_n562));
  OAI21_X1  g361(.A(new_n478), .B1(new_n485), .B2(new_n490), .ZN(new_n563));
  NAND2_X1  g362(.A1(new_n563), .A2(new_n492), .ZN(new_n564));
  AOI21_X1  g363(.A(new_n491), .B1(new_n564), .B2(KEYINPUT77), .ZN(new_n565));
  INV_X1    g364(.A(KEYINPUT77), .ZN(new_n566));
  NAND3_X1  g365(.A1(new_n563), .A2(new_n566), .A3(new_n492), .ZN(new_n567));
  AOI21_X1  g366(.A(new_n562), .B1(new_n565), .B2(new_n567), .ZN(new_n568));
  AOI21_X1  g367(.A(new_n534), .B1(new_n558), .B2(new_n568), .ZN(new_n569));
  NOR2_X1   g368(.A1(new_n358), .A2(new_n360), .ZN(new_n570));
  AOI21_X1  g369(.A(new_n364), .B1(new_n570), .B2(new_n375), .ZN(new_n571));
  AOI21_X1  g370(.A(new_n370), .B1(new_n351), .B2(new_n362), .ZN(new_n572));
  OAI22_X1  g371(.A1(new_n571), .A2(new_n351), .B1(new_n363), .B2(new_n572), .ZN(new_n573));
  NAND3_X1  g372(.A1(new_n332), .A2(new_n337), .A3(new_n338), .ZN(new_n574));
  INV_X1    g373(.A(new_n345), .ZN(new_n575));
  AOI21_X1  g374(.A(new_n574), .B1(new_n575), .B2(KEYINPUT28), .ZN(new_n576));
  OAI21_X1  g375(.A(new_n460), .B1(new_n573), .B2(new_n576), .ZN(new_n577));
  NAND2_X1  g376(.A1(G227gat), .A2(G233gat), .ZN(new_n578));
  INV_X1    g377(.A(new_n578), .ZN(new_n579));
  NAND4_X1  g378(.A1(new_n346), .A2(new_n365), .A3(new_n371), .A4(new_n457), .ZN(new_n580));
  NAND3_X1  g379(.A1(new_n577), .A2(new_n579), .A3(new_n580), .ZN(new_n581));
  XNOR2_X1  g380(.A(G15gat), .B(G43gat), .ZN(new_n582));
  XNOR2_X1  g381(.A(new_n582), .B(G71gat), .ZN(new_n583));
  INV_X1    g382(.A(G99gat), .ZN(new_n584));
  XNOR2_X1  g383(.A(new_n583), .B(new_n584), .ZN(new_n585));
  NAND2_X1  g384(.A1(new_n585), .A2(KEYINPUT33), .ZN(new_n586));
  NAND3_X1  g385(.A1(new_n581), .A2(KEYINPUT32), .A3(new_n586), .ZN(new_n587));
  INV_X1    g386(.A(KEYINPUT69), .ZN(new_n588));
  NAND2_X1  g387(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  NAND4_X1  g388(.A1(new_n581), .A2(KEYINPUT69), .A3(KEYINPUT32), .A4(new_n586), .ZN(new_n590));
  NAND2_X1  g389(.A1(new_n589), .A2(new_n590), .ZN(new_n591));
  INV_X1    g390(.A(KEYINPUT33), .ZN(new_n592));
  OAI21_X1  g391(.A(new_n581), .B1(KEYINPUT32), .B2(new_n592), .ZN(new_n593));
  NAND2_X1  g392(.A1(new_n593), .A2(new_n585), .ZN(new_n594));
  NAND2_X1  g393(.A1(new_n591), .A2(new_n594), .ZN(new_n595));
  AOI21_X1  g394(.A(new_n579), .B1(new_n577), .B2(new_n580), .ZN(new_n596));
  XNOR2_X1  g395(.A(new_n596), .B(KEYINPUT34), .ZN(new_n597));
  INV_X1    g396(.A(new_n597), .ZN(new_n598));
  NAND2_X1  g397(.A1(new_n595), .A2(new_n598), .ZN(new_n599));
  NAND3_X1  g398(.A1(new_n591), .A2(new_n597), .A3(new_n594), .ZN(new_n600));
  NAND3_X1  g399(.A1(new_n599), .A2(KEYINPUT36), .A3(new_n600), .ZN(new_n601));
  NAND3_X1  g400(.A1(new_n599), .A2(KEYINPUT70), .A3(new_n600), .ZN(new_n602));
  INV_X1    g401(.A(KEYINPUT36), .ZN(new_n603));
  AOI21_X1  g402(.A(new_n597), .B1(new_n591), .B2(new_n594), .ZN(new_n604));
  INV_X1    g403(.A(KEYINPUT70), .ZN(new_n605));
  NAND2_X1  g404(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  NAND3_X1  g405(.A1(new_n602), .A2(new_n603), .A3(new_n606), .ZN(new_n607));
  AOI21_X1  g406(.A(new_n569), .B1(new_n601), .B2(new_n607), .ZN(new_n608));
  NAND2_X1  g407(.A1(new_n561), .A2(new_n608), .ZN(new_n609));
  AND3_X1   g408(.A1(new_n591), .A2(new_n597), .A3(new_n594), .ZN(new_n610));
  NOR3_X1   g409(.A1(new_n610), .A2(new_n604), .A3(new_n535), .ZN(new_n611));
  NAND3_X1  g410(.A1(new_n558), .A2(new_n611), .A3(new_n568), .ZN(new_n612));
  NAND2_X1  g411(.A1(new_n612), .A2(KEYINPUT35), .ZN(new_n613));
  NAND2_X1  g412(.A1(new_n613), .A2(KEYINPUT87), .ZN(new_n614));
  INV_X1    g413(.A(KEYINPUT87), .ZN(new_n615));
  NAND3_X1  g414(.A1(new_n612), .A2(new_n615), .A3(KEYINPUT35), .ZN(new_n616));
  INV_X1    g415(.A(KEYINPUT86), .ZN(new_n617));
  NAND2_X1  g416(.A1(new_n602), .A2(new_n606), .ZN(new_n618));
  INV_X1    g417(.A(new_n618), .ZN(new_n619));
  INV_X1    g418(.A(KEYINPUT35), .ZN(new_n620));
  NAND4_X1  g419(.A1(new_n484), .A2(new_n620), .A3(new_n493), .A4(new_n534), .ZN(new_n621));
  INV_X1    g420(.A(new_n621), .ZN(new_n622));
  NAND2_X1  g421(.A1(new_n558), .A2(new_n622), .ZN(new_n623));
  OAI21_X1  g422(.A(new_n617), .B1(new_n619), .B2(new_n623), .ZN(new_n624));
  AND3_X1   g423(.A1(new_n513), .A2(KEYINPUT74), .A3(new_n512), .ZN(new_n625));
  AOI21_X1  g424(.A(KEYINPUT74), .B1(new_n513), .B2(new_n512), .ZN(new_n626));
  NOR2_X1   g425(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  XNOR2_X1  g426(.A(new_n410), .B(new_n556), .ZN(new_n628));
  NOR3_X1   g427(.A1(new_n627), .A2(new_n628), .A3(new_n621), .ZN(new_n629));
  NAND3_X1  g428(.A1(new_n629), .A2(KEYINPUT86), .A3(new_n618), .ZN(new_n630));
  NAND4_X1  g429(.A1(new_n614), .A2(new_n616), .A3(new_n624), .A4(new_n630), .ZN(new_n631));
  NAND2_X1  g430(.A1(new_n609), .A2(new_n631), .ZN(new_n632));
  INV_X1    g431(.A(KEYINPUT21), .ZN(new_n633));
  OAI21_X1  g432(.A(new_n235), .B1(new_n633), .B2(new_n276), .ZN(new_n634));
  NAND2_X1  g433(.A1(new_n276), .A2(new_n633), .ZN(new_n635));
  XOR2_X1   g434(.A(new_n635), .B(G127gat), .Z(new_n636));
  XNOR2_X1  g435(.A(new_n634), .B(new_n636), .ZN(new_n637));
  XNOR2_X1  g436(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n638));
  XNOR2_X1  g437(.A(G155gat), .B(G183gat), .ZN(new_n639));
  XNOR2_X1  g438(.A(new_n638), .B(new_n639), .ZN(new_n640));
  XNOR2_X1  g439(.A(new_n637), .B(new_n640), .ZN(new_n641));
  NAND2_X1  g440(.A1(G231gat), .A2(G233gat), .ZN(new_n642));
  XNOR2_X1  g441(.A(new_n642), .B(new_n389), .ZN(new_n643));
  INV_X1    g442(.A(new_n643), .ZN(new_n644));
  XNOR2_X1  g443(.A(new_n641), .B(new_n644), .ZN(new_n645));
  AOI21_X1  g444(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n646));
  XNOR2_X1  g445(.A(new_n646), .B(G134gat), .ZN(new_n647));
  XNOR2_X1  g446(.A(new_n647), .B(G162gat), .ZN(new_n648));
  OAI211_X1 g447(.A(new_n288), .B(new_n242), .C1(new_n220), .C2(KEYINPUT17), .ZN(new_n649));
  NAND3_X1  g448(.A1(new_n218), .A2(new_n294), .A3(new_n219), .ZN(new_n650));
  NAND3_X1  g449(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n651));
  NAND3_X1  g450(.A1(new_n649), .A2(new_n650), .A3(new_n651), .ZN(new_n652));
  XNOR2_X1  g451(.A(G190gat), .B(G218gat), .ZN(new_n653));
  NAND2_X1  g452(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  INV_X1    g453(.A(KEYINPUT94), .ZN(new_n655));
  AOI21_X1  g454(.A(new_n648), .B1(new_n654), .B2(new_n655), .ZN(new_n656));
  INV_X1    g455(.A(KEYINPUT93), .ZN(new_n657));
  NAND2_X1  g456(.A1(new_n654), .A2(new_n657), .ZN(new_n658));
  NAND2_X1  g457(.A1(new_n656), .A2(new_n658), .ZN(new_n659));
  NOR2_X1   g458(.A1(new_n652), .A2(new_n653), .ZN(new_n660));
  OAI211_X1 g459(.A(new_n654), .B(new_n657), .C1(new_n655), .C2(new_n648), .ZN(new_n661));
  AND3_X1   g460(.A1(new_n659), .A2(new_n660), .A3(new_n661), .ZN(new_n662));
  AOI21_X1  g461(.A(new_n660), .B1(new_n659), .B2(new_n661), .ZN(new_n663));
  NOR2_X1   g462(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  AND4_X1   g463(.A1(new_n324), .A2(new_n632), .A3(new_n645), .A4(new_n664), .ZN(new_n665));
  INV_X1    g464(.A(new_n568), .ZN(new_n666));
  NAND2_X1  g465(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  XNOR2_X1  g466(.A(new_n667), .B(G1gat), .ZN(G1324gat));
  NAND2_X1  g467(.A1(KEYINPUT16), .A2(G8gat), .ZN(new_n669));
  NAND3_X1  g468(.A1(new_n665), .A2(new_n559), .A3(new_n669), .ZN(new_n670));
  AOI21_X1  g469(.A(new_n670), .B1(new_n227), .B2(new_n231), .ZN(new_n671));
  AOI21_X1  g470(.A(new_n231), .B1(new_n665), .B2(new_n559), .ZN(new_n672));
  OAI21_X1  g471(.A(KEYINPUT42), .B1(new_n671), .B2(new_n672), .ZN(new_n673));
  OAI21_X1  g472(.A(new_n673), .B1(KEYINPUT42), .B2(new_n671), .ZN(G1325gat));
  AOI21_X1  g473(.A(G15gat), .B1(new_n665), .B2(new_n618), .ZN(new_n675));
  NAND2_X1  g474(.A1(new_n607), .A2(new_n601), .ZN(new_n676));
  INV_X1    g475(.A(new_n676), .ZN(new_n677));
  AND2_X1   g476(.A1(new_n677), .A2(G15gat), .ZN(new_n678));
  AOI21_X1  g477(.A(new_n675), .B1(new_n665), .B2(new_n678), .ZN(G1326gat));
  NAND2_X1  g478(.A1(new_n665), .A2(new_n535), .ZN(new_n680));
  XOR2_X1   g479(.A(new_n680), .B(KEYINPUT99), .Z(new_n681));
  XNOR2_X1  g480(.A(new_n681), .B(KEYINPUT43), .ZN(new_n682));
  XNOR2_X1  g481(.A(new_n682), .B(G22gat), .ZN(G1327gat));
  AND3_X1   g482(.A1(new_n612), .A2(new_n615), .A3(KEYINPUT35), .ZN(new_n684));
  AOI21_X1  g483(.A(new_n615), .B1(new_n612), .B2(KEYINPUT35), .ZN(new_n685));
  NOR2_X1   g484(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  AND4_X1   g485(.A1(KEYINPUT86), .A2(new_n618), .A3(new_n558), .A4(new_n622), .ZN(new_n687));
  AOI21_X1  g486(.A(KEYINPUT86), .B1(new_n629), .B2(new_n618), .ZN(new_n688));
  NOR2_X1   g487(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  AOI22_X1  g488(.A1(new_n686), .A2(new_n689), .B1(new_n561), .B2(new_n608), .ZN(new_n690));
  OAI21_X1  g489(.A(KEYINPUT44), .B1(new_n690), .B2(new_n664), .ZN(new_n691));
  INV_X1    g490(.A(KEYINPUT44), .ZN(new_n692));
  INV_X1    g491(.A(new_n664), .ZN(new_n693));
  NAND3_X1  g492(.A1(new_n632), .A2(new_n692), .A3(new_n693), .ZN(new_n694));
  NAND2_X1  g493(.A1(new_n691), .A2(new_n694), .ZN(new_n695));
  INV_X1    g494(.A(new_n695), .ZN(new_n696));
  INV_X1    g495(.A(new_n645), .ZN(new_n697));
  NAND2_X1  g496(.A1(new_n324), .A2(new_n697), .ZN(new_n698));
  NOR2_X1   g497(.A1(new_n696), .A2(new_n698), .ZN(new_n699));
  INV_X1    g498(.A(new_n699), .ZN(new_n700));
  OAI21_X1  g499(.A(G29gat), .B1(new_n700), .B2(new_n568), .ZN(new_n701));
  NOR3_X1   g500(.A1(new_n690), .A2(new_n664), .A3(new_n698), .ZN(new_n702));
  NAND3_X1  g501(.A1(new_n702), .A2(new_n205), .A3(new_n666), .ZN(new_n703));
  XNOR2_X1  g502(.A(new_n703), .B(KEYINPUT45), .ZN(new_n704));
  NAND2_X1  g503(.A1(new_n701), .A2(new_n704), .ZN(G1328gat));
  OAI21_X1  g504(.A(G36gat), .B1(new_n700), .B2(new_n558), .ZN(new_n706));
  NAND3_X1  g505(.A1(new_n702), .A2(new_n206), .A3(new_n559), .ZN(new_n707));
  XOR2_X1   g506(.A(new_n707), .B(KEYINPUT46), .Z(new_n708));
  NAND2_X1  g507(.A1(new_n706), .A2(new_n708), .ZN(G1329gat));
  OR3_X1    g508(.A1(new_n700), .A2(KEYINPUT100), .A3(new_n676), .ZN(new_n710));
  OAI21_X1  g509(.A(KEYINPUT100), .B1(new_n700), .B2(new_n676), .ZN(new_n711));
  NAND3_X1  g510(.A1(new_n710), .A2(G43gat), .A3(new_n711), .ZN(new_n712));
  INV_X1    g511(.A(G43gat), .ZN(new_n713));
  NAND3_X1  g512(.A1(new_n702), .A2(new_n713), .A3(new_n618), .ZN(new_n714));
  NAND3_X1  g513(.A1(new_n712), .A2(KEYINPUT47), .A3(new_n714), .ZN(new_n715));
  OAI21_X1  g514(.A(G43gat), .B1(new_n700), .B2(new_n676), .ZN(new_n716));
  AND2_X1   g515(.A1(new_n716), .A2(new_n714), .ZN(new_n717));
  OAI21_X1  g516(.A(new_n715), .B1(KEYINPUT47), .B2(new_n717), .ZN(G1330gat));
  INV_X1    g517(.A(KEYINPUT48), .ZN(new_n719));
  NAND2_X1  g518(.A1(new_n699), .A2(new_n535), .ZN(new_n720));
  NAND2_X1  g519(.A1(new_n720), .A2(G50gat), .ZN(new_n721));
  AOI21_X1  g520(.A(new_n719), .B1(new_n721), .B2(KEYINPUT102), .ZN(new_n722));
  NAND2_X1  g521(.A1(new_n535), .A2(new_n530), .ZN(new_n723));
  XNOR2_X1  g522(.A(new_n723), .B(KEYINPUT101), .ZN(new_n724));
  AOI22_X1  g523(.A1(new_n720), .A2(G50gat), .B1(new_n702), .B2(new_n724), .ZN(new_n725));
  XNOR2_X1  g524(.A(new_n722), .B(new_n725), .ZN(G1331gat));
  NAND3_X1  g525(.A1(new_n664), .A2(new_n264), .A3(new_n645), .ZN(new_n727));
  NOR2_X1   g526(.A1(new_n690), .A2(new_n727), .ZN(new_n728));
  NAND2_X1  g527(.A1(new_n728), .A2(new_n323), .ZN(new_n729));
  NOR2_X1   g528(.A1(new_n729), .A2(new_n568), .ZN(new_n730));
  XOR2_X1   g529(.A(KEYINPUT103), .B(G57gat), .Z(new_n731));
  XNOR2_X1  g530(.A(new_n730), .B(new_n731), .ZN(G1332gat));
  AOI211_X1 g531(.A(new_n558), .B(new_n729), .C1(KEYINPUT49), .C2(G64gat), .ZN(new_n733));
  NOR2_X1   g532(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n734));
  XNOR2_X1  g533(.A(new_n733), .B(new_n734), .ZN(G1333gat));
  OAI21_X1  g534(.A(G71gat), .B1(new_n729), .B2(new_n676), .ZN(new_n736));
  OR2_X1    g535(.A1(new_n619), .A2(G71gat), .ZN(new_n737));
  OAI21_X1  g536(.A(new_n736), .B1(new_n729), .B2(new_n737), .ZN(new_n738));
  XOR2_X1   g537(.A(new_n738), .B(KEYINPUT50), .Z(G1334gat));
  NOR2_X1   g538(.A1(new_n729), .A2(new_n534), .ZN(new_n740));
  XOR2_X1   g539(.A(new_n740), .B(G78gat), .Z(G1335gat));
  NOR2_X1   g540(.A1(new_n645), .A2(new_n263), .ZN(new_n742));
  NAND2_X1  g541(.A1(new_n742), .A2(new_n323), .ZN(new_n743));
  NAND2_X1  g542(.A1(new_n743), .A2(KEYINPUT104), .ZN(new_n744));
  INV_X1    g543(.A(KEYINPUT104), .ZN(new_n745));
  NAND3_X1  g544(.A1(new_n742), .A2(new_n745), .A3(new_n323), .ZN(new_n746));
  NAND2_X1  g545(.A1(new_n744), .A2(new_n746), .ZN(new_n747));
  INV_X1    g546(.A(new_n747), .ZN(new_n748));
  AOI21_X1  g547(.A(KEYINPUT105), .B1(new_n695), .B2(new_n748), .ZN(new_n749));
  INV_X1    g548(.A(KEYINPUT105), .ZN(new_n750));
  AOI211_X1 g549(.A(new_n750), .B(new_n747), .C1(new_n691), .C2(new_n694), .ZN(new_n751));
  NOR2_X1   g550(.A1(new_n749), .A2(new_n751), .ZN(new_n752));
  OAI21_X1  g551(.A(G85gat), .B1(new_n752), .B2(new_n568), .ZN(new_n753));
  NOR2_X1   g552(.A1(new_n690), .A2(new_n664), .ZN(new_n754));
  NAND2_X1  g553(.A1(new_n754), .A2(new_n742), .ZN(new_n755));
  INV_X1    g554(.A(KEYINPUT51), .ZN(new_n756));
  NAND2_X1  g555(.A1(new_n755), .A2(new_n756), .ZN(new_n757));
  INV_X1    g556(.A(KEYINPUT106), .ZN(new_n758));
  NAND3_X1  g557(.A1(new_n754), .A2(KEYINPUT51), .A3(new_n742), .ZN(new_n759));
  NAND3_X1  g558(.A1(new_n757), .A2(new_n758), .A3(new_n759), .ZN(new_n760));
  NAND3_X1  g559(.A1(new_n755), .A2(KEYINPUT106), .A3(new_n756), .ZN(new_n761));
  NAND2_X1  g560(.A1(new_n760), .A2(new_n761), .ZN(new_n762));
  INV_X1    g561(.A(new_n762), .ZN(new_n763));
  NAND3_X1  g562(.A1(new_n763), .A2(new_n280), .A3(new_n666), .ZN(new_n764));
  AND2_X1   g563(.A1(new_n320), .A2(new_n322), .ZN(new_n765));
  OAI21_X1  g564(.A(new_n753), .B1(new_n764), .B2(new_n765), .ZN(G1336gat));
  NOR3_X1   g565(.A1(new_n765), .A2(G92gat), .A3(new_n558), .ZN(new_n767));
  NAND2_X1  g566(.A1(new_n763), .A2(new_n767), .ZN(new_n768));
  INV_X1    g567(.A(KEYINPUT52), .ZN(new_n769));
  INV_X1    g568(.A(KEYINPUT108), .ZN(new_n770));
  AOI21_X1  g569(.A(new_n692), .B1(new_n632), .B2(new_n693), .ZN(new_n771));
  AOI211_X1 g570(.A(KEYINPUT44), .B(new_n664), .C1(new_n609), .C2(new_n631), .ZN(new_n772));
  OAI21_X1  g571(.A(new_n748), .B1(new_n771), .B2(new_n772), .ZN(new_n773));
  OAI21_X1  g572(.A(new_n770), .B1(new_n773), .B2(new_n558), .ZN(new_n774));
  NAND4_X1  g573(.A1(new_n695), .A2(KEYINPUT108), .A3(new_n559), .A4(new_n748), .ZN(new_n775));
  NAND3_X1  g574(.A1(new_n774), .A2(G92gat), .A3(new_n775), .ZN(new_n776));
  NAND3_X1  g575(.A1(new_n768), .A2(new_n769), .A3(new_n776), .ZN(new_n777));
  INV_X1    g576(.A(KEYINPUT107), .ZN(new_n778));
  NAND3_X1  g577(.A1(new_n757), .A2(new_n778), .A3(new_n759), .ZN(new_n779));
  NAND3_X1  g578(.A1(new_n755), .A2(KEYINPUT107), .A3(new_n756), .ZN(new_n780));
  AND2_X1   g579(.A1(new_n779), .A2(new_n780), .ZN(new_n781));
  OAI21_X1  g580(.A(new_n559), .B1(new_n749), .B2(new_n751), .ZN(new_n782));
  AOI22_X1  g581(.A1(new_n781), .A2(new_n767), .B1(new_n782), .B2(G92gat), .ZN(new_n783));
  OAI21_X1  g582(.A(new_n777), .B1(new_n769), .B2(new_n783), .ZN(G1337gat));
  OAI21_X1  g583(.A(G99gat), .B1(new_n752), .B2(new_n676), .ZN(new_n785));
  NAND3_X1  g584(.A1(new_n323), .A2(new_n584), .A3(new_n618), .ZN(new_n786));
  OAI21_X1  g585(.A(new_n785), .B1(new_n762), .B2(new_n786), .ZN(G1338gat));
  OAI21_X1  g586(.A(G106gat), .B1(new_n773), .B2(new_n534), .ZN(new_n788));
  INV_X1    g587(.A(KEYINPUT53), .ZN(new_n789));
  INV_X1    g588(.A(G106gat), .ZN(new_n790));
  NAND3_X1  g589(.A1(new_n323), .A2(new_n790), .A3(new_n535), .ZN(new_n791));
  OAI211_X1 g590(.A(new_n788), .B(new_n789), .C1(new_n762), .C2(new_n791), .ZN(new_n792));
  INV_X1    g591(.A(KEYINPUT109), .ZN(new_n793));
  NAND2_X1  g592(.A1(new_n773), .A2(new_n750), .ZN(new_n794));
  NAND3_X1  g593(.A1(new_n695), .A2(KEYINPUT105), .A3(new_n748), .ZN(new_n795));
  AOI21_X1  g594(.A(new_n534), .B1(new_n794), .B2(new_n795), .ZN(new_n796));
  OAI21_X1  g595(.A(new_n793), .B1(new_n796), .B2(new_n790), .ZN(new_n797));
  INV_X1    g596(.A(new_n791), .ZN(new_n798));
  NAND3_X1  g597(.A1(new_n779), .A2(new_n780), .A3(new_n798), .ZN(new_n799));
  OAI21_X1  g598(.A(new_n535), .B1(new_n749), .B2(new_n751), .ZN(new_n800));
  NAND3_X1  g599(.A1(new_n800), .A2(KEYINPUT109), .A3(G106gat), .ZN(new_n801));
  NAND3_X1  g600(.A1(new_n797), .A2(new_n799), .A3(new_n801), .ZN(new_n802));
  AND3_X1   g601(.A1(new_n802), .A2(KEYINPUT110), .A3(KEYINPUT53), .ZN(new_n803));
  AOI21_X1  g602(.A(KEYINPUT110), .B1(new_n802), .B2(KEYINPUT53), .ZN(new_n804));
  OAI21_X1  g603(.A(new_n792), .B1(new_n803), .B2(new_n804), .ZN(G1339gat));
  INV_X1    g604(.A(KEYINPUT117), .ZN(new_n806));
  NOR2_X1   g605(.A1(new_n727), .A2(new_n323), .ZN(new_n807));
  XNOR2_X1  g606(.A(new_n807), .B(KEYINPUT111), .ZN(new_n808));
  AND3_X1   g607(.A1(new_n239), .A2(new_n247), .A3(new_n249), .ZN(new_n809));
  AOI21_X1  g608(.A(new_n240), .B1(new_n239), .B2(new_n243), .ZN(new_n810));
  OAI21_X1  g609(.A(new_n258), .B1(new_n809), .B2(new_n810), .ZN(new_n811));
  NAND2_X1  g610(.A1(new_n811), .A2(KEYINPUT114), .ZN(new_n812));
  INV_X1    g611(.A(KEYINPUT114), .ZN(new_n813));
  OAI211_X1 g612(.A(new_n813), .B(new_n258), .C1(new_n809), .C2(new_n810), .ZN(new_n814));
  NAND2_X1  g613(.A1(new_n812), .A2(new_n814), .ZN(new_n815));
  NAND2_X1  g614(.A1(new_n815), .A2(new_n262), .ZN(new_n816));
  OAI21_X1  g615(.A(KEYINPUT115), .B1(new_n816), .B2(new_n765), .ZN(new_n817));
  INV_X1    g616(.A(KEYINPUT55), .ZN(new_n818));
  INV_X1    g617(.A(KEYINPUT112), .ZN(new_n819));
  INV_X1    g618(.A(KEYINPUT54), .ZN(new_n820));
  NAND3_X1  g619(.A1(new_n313), .A2(new_n310), .A3(new_n296), .ZN(new_n821));
  OAI21_X1  g620(.A(KEYINPUT96), .B1(new_n293), .B2(new_n297), .ZN(new_n822));
  NAND2_X1  g621(.A1(new_n821), .A2(new_n822), .ZN(new_n823));
  AOI21_X1  g622(.A(new_n820), .B1(new_n823), .B2(new_n265), .ZN(new_n824));
  NOR3_X1   g623(.A1(new_n293), .A2(new_n265), .A3(new_n297), .ZN(new_n825));
  INV_X1    g624(.A(new_n825), .ZN(new_n826));
  AOI21_X1  g625(.A(new_n819), .B1(new_n824), .B2(new_n826), .ZN(new_n827));
  AOI21_X1  g626(.A(new_n300), .B1(new_n821), .B2(new_n822), .ZN(new_n828));
  NOR4_X1   g627(.A1(new_n828), .A2(KEYINPUT112), .A3(new_n825), .A4(new_n820), .ZN(new_n829));
  NOR2_X1   g628(.A1(new_n827), .A2(new_n829), .ZN(new_n830));
  NAND2_X1  g629(.A1(new_n299), .A2(new_n303), .ZN(new_n831));
  NAND2_X1  g630(.A1(new_n831), .A2(new_n820), .ZN(new_n832));
  INV_X1    g631(.A(KEYINPUT113), .ZN(new_n833));
  NAND3_X1  g632(.A1(new_n832), .A2(new_n833), .A3(new_n308), .ZN(new_n834));
  AOI21_X1  g633(.A(KEYINPUT54), .B1(new_n299), .B2(new_n303), .ZN(new_n835));
  OAI21_X1  g634(.A(KEYINPUT113), .B1(new_n835), .B2(new_n317), .ZN(new_n836));
  NAND2_X1  g635(.A1(new_n834), .A2(new_n836), .ZN(new_n837));
  OAI21_X1  g636(.A(new_n818), .B1(new_n830), .B2(new_n837), .ZN(new_n838));
  NAND3_X1  g637(.A1(new_n316), .A2(KEYINPUT54), .A3(new_n826), .ZN(new_n839));
  NAND2_X1  g638(.A1(new_n839), .A2(KEYINPUT112), .ZN(new_n840));
  NAND3_X1  g639(.A1(new_n824), .A2(new_n819), .A3(new_n826), .ZN(new_n841));
  NAND2_X1  g640(.A1(new_n840), .A2(new_n841), .ZN(new_n842));
  NAND4_X1  g641(.A1(new_n842), .A2(KEYINPUT55), .A3(new_n834), .A4(new_n836), .ZN(new_n843));
  NAND4_X1  g642(.A1(new_n838), .A2(new_n843), .A3(new_n318), .A4(new_n263), .ZN(new_n844));
  INV_X1    g643(.A(KEYINPUT115), .ZN(new_n845));
  NAND4_X1  g644(.A1(new_n323), .A2(new_n815), .A3(new_n845), .A4(new_n262), .ZN(new_n846));
  NAND3_X1  g645(.A1(new_n817), .A2(new_n844), .A3(new_n846), .ZN(new_n847));
  OAI21_X1  g646(.A(new_n838), .B1(new_n662), .B2(new_n663), .ZN(new_n848));
  NAND2_X1  g647(.A1(new_n843), .A2(new_n318), .ZN(new_n849));
  NOR2_X1   g648(.A1(new_n848), .A2(new_n849), .ZN(new_n850));
  INV_X1    g649(.A(new_n816), .ZN(new_n851));
  AOI22_X1  g650(.A1(new_n847), .A2(new_n664), .B1(new_n850), .B2(new_n851), .ZN(new_n852));
  INV_X1    g651(.A(KEYINPUT116), .ZN(new_n853));
  AOI21_X1  g652(.A(new_n645), .B1(new_n852), .B2(new_n853), .ZN(new_n854));
  NAND2_X1  g653(.A1(new_n847), .A2(new_n664), .ZN(new_n855));
  NAND2_X1  g654(.A1(new_n850), .A2(new_n851), .ZN(new_n856));
  NAND2_X1  g655(.A1(new_n855), .A2(new_n856), .ZN(new_n857));
  NAND2_X1  g656(.A1(new_n857), .A2(KEYINPUT116), .ZN(new_n858));
  AOI21_X1  g657(.A(new_n808), .B1(new_n854), .B2(new_n858), .ZN(new_n859));
  OAI21_X1  g658(.A(new_n806), .B1(new_n859), .B2(new_n535), .ZN(new_n860));
  INV_X1    g659(.A(KEYINPUT111), .ZN(new_n861));
  XNOR2_X1  g660(.A(new_n807), .B(new_n861), .ZN(new_n862));
  NAND3_X1  g661(.A1(new_n855), .A2(new_n853), .A3(new_n856), .ZN(new_n863));
  NAND2_X1  g662(.A1(new_n863), .A2(new_n697), .ZN(new_n864));
  NOR2_X1   g663(.A1(new_n852), .A2(new_n853), .ZN(new_n865));
  OAI21_X1  g664(.A(new_n862), .B1(new_n864), .B2(new_n865), .ZN(new_n866));
  NAND3_X1  g665(.A1(new_n866), .A2(KEYINPUT117), .A3(new_n534), .ZN(new_n867));
  NAND2_X1  g666(.A1(new_n860), .A2(new_n867), .ZN(new_n868));
  NOR2_X1   g667(.A1(new_n559), .A2(new_n568), .ZN(new_n869));
  NAND3_X1  g668(.A1(new_n868), .A2(new_n618), .A3(new_n869), .ZN(new_n870));
  OAI21_X1  g669(.A(G113gat), .B1(new_n870), .B2(new_n264), .ZN(new_n871));
  INV_X1    g670(.A(new_n611), .ZN(new_n872));
  NOR2_X1   g671(.A1(new_n859), .A2(new_n872), .ZN(new_n873));
  AND2_X1   g672(.A1(new_n873), .A2(new_n869), .ZN(new_n874));
  NAND2_X1  g673(.A1(new_n263), .A2(new_n455), .ZN(new_n875));
  XNOR2_X1  g674(.A(new_n875), .B(KEYINPUT118), .ZN(new_n876));
  NAND2_X1  g675(.A1(new_n874), .A2(new_n876), .ZN(new_n877));
  NAND2_X1  g676(.A1(new_n871), .A2(new_n877), .ZN(G1340gat));
  OAI21_X1  g677(.A(G120gat), .B1(new_n870), .B2(new_n765), .ZN(new_n879));
  NAND3_X1  g678(.A1(new_n874), .A2(new_n445), .A3(new_n323), .ZN(new_n880));
  NAND2_X1  g679(.A1(new_n879), .A2(new_n880), .ZN(G1341gat));
  NAND2_X1  g680(.A1(new_n450), .A2(new_n451), .ZN(new_n882));
  AND4_X1   g681(.A1(new_n882), .A2(new_n873), .A3(new_n645), .A4(new_n869), .ZN(new_n883));
  NAND4_X1  g682(.A1(new_n868), .A2(new_n645), .A3(new_n618), .A4(new_n869), .ZN(new_n884));
  INV_X1    g683(.A(new_n882), .ZN(new_n885));
  AOI21_X1  g684(.A(new_n883), .B1(new_n884), .B2(new_n885), .ZN(new_n886));
  INV_X1    g685(.A(KEYINPUT119), .ZN(new_n887));
  NOR2_X1   g686(.A1(new_n886), .A2(new_n887), .ZN(new_n888));
  AOI211_X1 g687(.A(KEYINPUT119), .B(new_n883), .C1(new_n884), .C2(new_n885), .ZN(new_n889));
  NOR2_X1   g688(.A1(new_n888), .A2(new_n889), .ZN(G1342gat));
  INV_X1    g689(.A(G134gat), .ZN(new_n891));
  NAND3_X1  g690(.A1(new_n874), .A2(new_n891), .A3(new_n693), .ZN(new_n892));
  OR2_X1    g691(.A1(new_n892), .A2(KEYINPUT56), .ZN(new_n893));
  OAI21_X1  g692(.A(G134gat), .B1(new_n870), .B2(new_n664), .ZN(new_n894));
  NAND2_X1  g693(.A1(new_n892), .A2(KEYINPUT56), .ZN(new_n895));
  NAND3_X1  g694(.A1(new_n893), .A2(new_n894), .A3(new_n895), .ZN(G1343gat));
  NOR2_X1   g695(.A1(new_n859), .A2(new_n534), .ZN(new_n897));
  INV_X1    g696(.A(KEYINPUT57), .ZN(new_n898));
  NAND2_X1  g697(.A1(new_n897), .A2(new_n898), .ZN(new_n899));
  AND2_X1   g698(.A1(new_n869), .A2(new_n676), .ZN(new_n900));
  XNOR2_X1  g699(.A(new_n900), .B(KEYINPUT120), .ZN(new_n901));
  INV_X1    g700(.A(new_n901), .ZN(new_n902));
  OR3_X1    g701(.A1(new_n816), .A2(new_n765), .A3(KEYINPUT121), .ZN(new_n903));
  OAI21_X1  g702(.A(KEYINPUT121), .B1(new_n816), .B2(new_n765), .ZN(new_n904));
  NAND3_X1  g703(.A1(new_n903), .A2(new_n844), .A3(new_n904), .ZN(new_n905));
  NAND2_X1  g704(.A1(new_n905), .A2(new_n664), .ZN(new_n906));
  AOI21_X1  g705(.A(new_n645), .B1(new_n906), .B2(new_n856), .ZN(new_n907));
  OAI21_X1  g706(.A(new_n535), .B1(new_n907), .B2(new_n808), .ZN(new_n908));
  AOI21_X1  g707(.A(new_n902), .B1(new_n908), .B2(KEYINPUT57), .ZN(new_n909));
  NAND2_X1  g708(.A1(new_n899), .A2(new_n909), .ZN(new_n910));
  OAI21_X1  g709(.A(G141gat), .B1(new_n910), .B2(new_n264), .ZN(new_n911));
  AND2_X1   g710(.A1(new_n897), .A2(new_n900), .ZN(new_n912));
  NAND3_X1  g711(.A1(new_n912), .A2(new_n422), .A3(new_n263), .ZN(new_n913));
  NAND2_X1  g712(.A1(new_n911), .A2(new_n913), .ZN(new_n914));
  NAND2_X1  g713(.A1(new_n914), .A2(KEYINPUT58), .ZN(new_n915));
  INV_X1    g714(.A(KEYINPUT58), .ZN(new_n916));
  NAND3_X1  g715(.A1(new_n911), .A2(new_n916), .A3(new_n913), .ZN(new_n917));
  NAND2_X1  g716(.A1(new_n915), .A2(new_n917), .ZN(G1344gat));
  NAND3_X1  g717(.A1(new_n912), .A2(new_n441), .A3(new_n323), .ZN(new_n919));
  INV_X1    g718(.A(new_n910), .ZN(new_n920));
  AOI211_X1 g719(.A(KEYINPUT59), .B(new_n441), .C1(new_n920), .C2(new_n323), .ZN(new_n921));
  INV_X1    g720(.A(KEYINPUT59), .ZN(new_n922));
  OAI21_X1  g721(.A(KEYINPUT57), .B1(new_n859), .B2(new_n534), .ZN(new_n923));
  OAI211_X1 g722(.A(new_n898), .B(new_n535), .C1(new_n907), .C2(new_n807), .ZN(new_n924));
  AND2_X1   g723(.A1(new_n923), .A2(new_n924), .ZN(new_n925));
  NAND3_X1  g724(.A1(new_n925), .A2(new_n323), .A3(new_n901), .ZN(new_n926));
  AOI21_X1  g725(.A(new_n922), .B1(new_n926), .B2(G148gat), .ZN(new_n927));
  OAI21_X1  g726(.A(new_n919), .B1(new_n921), .B2(new_n927), .ZN(G1345gat));
  OAI21_X1  g727(.A(G155gat), .B1(new_n910), .B2(new_n697), .ZN(new_n929));
  INV_X1    g728(.A(G155gat), .ZN(new_n930));
  NAND3_X1  g729(.A1(new_n912), .A2(new_n930), .A3(new_n645), .ZN(new_n931));
  NAND2_X1  g730(.A1(new_n929), .A2(new_n931), .ZN(G1346gat));
  AOI21_X1  g731(.A(G162gat), .B1(new_n912), .B2(new_n693), .ZN(new_n933));
  AND2_X1   g732(.A1(new_n693), .A2(G162gat), .ZN(new_n934));
  AOI21_X1  g733(.A(new_n933), .B1(new_n920), .B2(new_n934), .ZN(G1347gat));
  NOR2_X1   g734(.A1(new_n666), .A2(new_n558), .ZN(new_n936));
  INV_X1    g735(.A(new_n936), .ZN(new_n937));
  NOR3_X1   g736(.A1(new_n859), .A2(new_n872), .A3(new_n937), .ZN(new_n938));
  NAND3_X1  g737(.A1(new_n938), .A2(new_n257), .A3(new_n263), .ZN(new_n939));
  NAND4_X1  g738(.A1(new_n868), .A2(new_n263), .A3(new_n618), .A4(new_n936), .ZN(new_n940));
  AND3_X1   g739(.A1(new_n940), .A2(KEYINPUT122), .A3(G169gat), .ZN(new_n941));
  AOI21_X1  g740(.A(KEYINPUT122), .B1(new_n940), .B2(G169gat), .ZN(new_n942));
  OAI21_X1  g741(.A(new_n939), .B1(new_n941), .B2(new_n942), .ZN(G1348gat));
  AOI21_X1  g742(.A(G176gat), .B1(new_n938), .B2(new_n323), .ZN(new_n944));
  AOI211_X1 g743(.A(new_n619), .B(new_n937), .C1(new_n860), .C2(new_n867), .ZN(new_n945));
  NOR2_X1   g744(.A1(new_n765), .A2(new_n306), .ZN(new_n946));
  AOI21_X1  g745(.A(new_n944), .B1(new_n945), .B2(new_n946), .ZN(G1349gat));
  INV_X1    g746(.A(G183gat), .ZN(new_n948));
  AOI21_X1  g747(.A(new_n948), .B1(new_n945), .B2(new_n645), .ZN(new_n949));
  INV_X1    g748(.A(new_n344), .ZN(new_n950));
  INV_X1    g749(.A(new_n343), .ZN(new_n951));
  OAI211_X1 g750(.A(new_n938), .B(new_n645), .C1(new_n950), .C2(new_n951), .ZN(new_n952));
  NAND2_X1  g751(.A1(new_n952), .A2(KEYINPUT123), .ZN(new_n953));
  OAI21_X1  g752(.A(KEYINPUT60), .B1(new_n949), .B2(new_n953), .ZN(new_n954));
  NAND3_X1  g753(.A1(new_n868), .A2(new_n618), .A3(new_n936), .ZN(new_n955));
  OAI21_X1  g754(.A(G183gat), .B1(new_n955), .B2(new_n697), .ZN(new_n956));
  INV_X1    g755(.A(KEYINPUT60), .ZN(new_n957));
  NAND4_X1  g756(.A1(new_n956), .A2(KEYINPUT123), .A3(new_n957), .A4(new_n952), .ZN(new_n958));
  NAND2_X1  g757(.A1(new_n954), .A2(new_n958), .ZN(G1350gat));
  NAND4_X1  g758(.A1(new_n868), .A2(new_n693), .A3(new_n618), .A4(new_n936), .ZN(new_n960));
  NAND2_X1  g759(.A1(KEYINPUT124), .A2(KEYINPUT61), .ZN(new_n961));
  NAND3_X1  g760(.A1(new_n960), .A2(G190gat), .A3(new_n961), .ZN(new_n962));
  NOR2_X1   g761(.A1(KEYINPUT124), .A2(KEYINPUT61), .ZN(new_n963));
  NAND2_X1  g762(.A1(new_n962), .A2(new_n963), .ZN(new_n964));
  NAND3_X1  g763(.A1(new_n938), .A2(new_n334), .A3(new_n693), .ZN(new_n965));
  INV_X1    g764(.A(new_n963), .ZN(new_n966));
  NAND4_X1  g765(.A1(new_n960), .A2(G190gat), .A3(new_n961), .A4(new_n966), .ZN(new_n967));
  NAND3_X1  g766(.A1(new_n964), .A2(new_n965), .A3(new_n967), .ZN(G1351gat));
  NOR2_X1   g767(.A1(new_n677), .A2(new_n937), .ZN(new_n969));
  NAND3_X1  g768(.A1(new_n923), .A2(new_n924), .A3(new_n969), .ZN(new_n970));
  OAI21_X1  g769(.A(G197gat), .B1(new_n970), .B2(new_n264), .ZN(new_n971));
  NAND2_X1  g770(.A1(new_n897), .A2(new_n969), .ZN(new_n972));
  OR2_X1    g771(.A1(new_n264), .A2(G197gat), .ZN(new_n973));
  OAI21_X1  g772(.A(new_n971), .B1(new_n972), .B2(new_n973), .ZN(G1352gat));
  XNOR2_X1  g773(.A(KEYINPUT125), .B(G204gat), .ZN(new_n975));
  NOR3_X1   g774(.A1(new_n972), .A2(new_n765), .A3(new_n975), .ZN(new_n976));
  XNOR2_X1  g775(.A(new_n976), .B(KEYINPUT62), .ZN(new_n977));
  NAND3_X1  g776(.A1(new_n925), .A2(new_n323), .A3(new_n969), .ZN(new_n978));
  NAND2_X1  g777(.A1(new_n978), .A2(new_n975), .ZN(new_n979));
  NAND2_X1  g778(.A1(new_n977), .A2(new_n979), .ZN(G1353gat));
  OAI21_X1  g779(.A(G211gat), .B1(new_n970), .B2(new_n697), .ZN(new_n981));
  INV_X1    g780(.A(KEYINPUT63), .ZN(new_n982));
  AND2_X1   g781(.A1(new_n981), .A2(new_n982), .ZN(new_n983));
  NOR2_X1   g782(.A1(new_n981), .A2(new_n982), .ZN(new_n984));
  NAND2_X1  g783(.A1(new_n645), .A2(new_n389), .ZN(new_n985));
  OAI22_X1  g784(.A1(new_n983), .A2(new_n984), .B1(new_n972), .B2(new_n985), .ZN(G1354gat));
  OR2_X1    g785(.A1(new_n970), .A2(KEYINPUT126), .ZN(new_n987));
  NAND3_X1  g786(.A1(new_n693), .A2(KEYINPUT127), .A3(G218gat), .ZN(new_n988));
  NAND2_X1  g787(.A1(new_n970), .A2(KEYINPUT126), .ZN(new_n989));
  INV_X1    g788(.A(KEYINPUT127), .ZN(new_n990));
  OAI21_X1  g789(.A(new_n990), .B1(new_n664), .B2(new_n390), .ZN(new_n991));
  NAND4_X1  g790(.A1(new_n987), .A2(new_n988), .A3(new_n989), .A4(new_n991), .ZN(new_n992));
  OAI21_X1  g791(.A(new_n390), .B1(new_n972), .B2(new_n664), .ZN(new_n993));
  AND2_X1   g792(.A1(new_n992), .A2(new_n993), .ZN(G1355gat));
endmodule


