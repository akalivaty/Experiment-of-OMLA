//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 0 0 1 0 0 1 0 0 0 0 0 1 0 1 1 1 1 1 0 1 0 1 0 0 0 0 1 1 1 0 1 0 1 0 1 0 1 0 0 1 1 1 0 0 0 1 0 1 1 0 0 0 0 0 1 1 1 0 1 0 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:40:44 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n204, new_n205, new_n206, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n245, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1239, new_n1240, new_n1242, new_n1243,
    new_n1244, new_n1245, new_n1246, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1301, new_n1302, new_n1303, new_n1304, new_n1305,
    new_n1306, new_n1307, new_n1308, new_n1309, new_n1310, new_n1311,
    new_n1312, new_n1313;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(new_n201), .ZN(new_n202));
  NOR3_X1   g0002(.A1(new_n202), .A2(G50), .A3(G77), .ZN(G353));
  INV_X1    g0003(.A(G97), .ZN(new_n204));
  INV_X1    g0004(.A(G107), .ZN(new_n205));
  NAND2_X1  g0005(.A1(new_n204), .A2(new_n205), .ZN(new_n206));
  NAND2_X1  g0006(.A1(new_n206), .A2(G87), .ZN(G355));
  INV_X1    g0007(.A(KEYINPUT64), .ZN(new_n208));
  NAND2_X1  g0008(.A1(G1), .A2(G20), .ZN(new_n209));
  OAI21_X1  g0009(.A(new_n208), .B1(new_n209), .B2(G13), .ZN(new_n210));
  INV_X1    g0010(.A(G13), .ZN(new_n211));
  NAND4_X1  g0011(.A1(new_n211), .A2(KEYINPUT64), .A3(G1), .A4(G20), .ZN(new_n212));
  NAND2_X1  g0012(.A1(new_n210), .A2(new_n212), .ZN(new_n213));
  OAI211_X1 g0013(.A(new_n213), .B(G250), .C1(G257), .C2(G264), .ZN(new_n214));
  XOR2_X1   g0014(.A(new_n214), .B(KEYINPUT0), .Z(new_n215));
  XNOR2_X1  g0015(.A(KEYINPUT65), .B(G238), .ZN(new_n216));
  INV_X1    g0016(.A(G68), .ZN(new_n217));
  NOR2_X1   g0017(.A1(new_n216), .A2(new_n217), .ZN(new_n218));
  AOI22_X1  g0018(.A1(G87), .A2(G250), .B1(G116), .B2(G270), .ZN(new_n219));
  AOI22_X1  g0019(.A1(G58), .A2(G232), .B1(G77), .B2(G244), .ZN(new_n220));
  AOI22_X1  g0020(.A1(G50), .A2(G226), .B1(G97), .B2(G257), .ZN(new_n221));
  NAND2_X1  g0021(.A1(G107), .A2(G264), .ZN(new_n222));
  NAND4_X1  g0022(.A1(new_n219), .A2(new_n220), .A3(new_n221), .A4(new_n222), .ZN(new_n223));
  OAI21_X1  g0023(.A(new_n209), .B1(new_n218), .B2(new_n223), .ZN(new_n224));
  XNOR2_X1  g0024(.A(new_n224), .B(KEYINPUT1), .ZN(new_n225));
  NAND2_X1  g0025(.A1(new_n202), .A2(G50), .ZN(new_n226));
  INV_X1    g0026(.A(G20), .ZN(new_n227));
  NAND2_X1  g0027(.A1(G1), .A2(G13), .ZN(new_n228));
  NOR3_X1   g0028(.A1(new_n226), .A2(new_n227), .A3(new_n228), .ZN(new_n229));
  NOR3_X1   g0029(.A1(new_n215), .A2(new_n225), .A3(new_n229), .ZN(G361));
  XNOR2_X1  g0030(.A(G238), .B(G244), .ZN(new_n231));
  INV_X1    g0031(.A(G232), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n231), .B(new_n232), .ZN(new_n233));
  XOR2_X1   g0033(.A(KEYINPUT2), .B(G226), .Z(new_n234));
  XNOR2_X1  g0034(.A(new_n233), .B(new_n234), .ZN(new_n235));
  XOR2_X1   g0035(.A(G264), .B(G270), .Z(new_n236));
  XNOR2_X1  g0036(.A(G250), .B(G257), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n235), .B(new_n238), .ZN(G358));
  XNOR2_X1  g0039(.A(G87), .B(G97), .ZN(new_n240));
  XNOR2_X1  g0040(.A(G107), .B(G116), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XNOR2_X1  g0042(.A(G50), .B(G68), .ZN(new_n243));
  XNOR2_X1  g0043(.A(G58), .B(G77), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n242), .B(new_n245), .ZN(G351));
  NAND3_X1  g0046(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n247));
  NAND2_X1  g0047(.A1(new_n247), .A2(new_n228), .ZN(new_n248));
  INV_X1    g0048(.A(new_n248), .ZN(new_n249));
  INV_X1    g0049(.A(G50), .ZN(new_n250));
  AOI21_X1  g0050(.A(new_n227), .B1(new_n201), .B2(new_n250), .ZN(new_n251));
  INV_X1    g0051(.A(KEYINPUT68), .ZN(new_n252));
  XNOR2_X1  g0052(.A(new_n251), .B(new_n252), .ZN(new_n253));
  XNOR2_X1  g0053(.A(KEYINPUT8), .B(G58), .ZN(new_n254));
  INV_X1    g0054(.A(new_n254), .ZN(new_n255));
  INV_X1    g0055(.A(G33), .ZN(new_n256));
  NOR2_X1   g0056(.A1(new_n256), .A2(G20), .ZN(new_n257));
  NOR2_X1   g0057(.A1(G20), .A2(G33), .ZN(new_n258));
  AOI22_X1  g0058(.A1(new_n255), .A2(new_n257), .B1(G150), .B2(new_n258), .ZN(new_n259));
  AOI21_X1  g0059(.A(new_n249), .B1(new_n253), .B2(new_n259), .ZN(new_n260));
  INV_X1    g0060(.A(G1), .ZN(new_n261));
  NAND3_X1  g0061(.A1(new_n261), .A2(G13), .A3(G20), .ZN(new_n262));
  INV_X1    g0062(.A(new_n262), .ZN(new_n263));
  NOR2_X1   g0063(.A1(new_n263), .A2(new_n248), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n261), .A2(G20), .ZN(new_n265));
  NAND3_X1  g0065(.A1(new_n264), .A2(G50), .A3(new_n265), .ZN(new_n266));
  OAI21_X1  g0066(.A(new_n266), .B1(G50), .B2(new_n262), .ZN(new_n267));
  NOR2_X1   g0067(.A1(new_n260), .A2(new_n267), .ZN(new_n268));
  AOI21_X1  g0068(.A(new_n228), .B1(G33), .B2(G41), .ZN(new_n269));
  INV_X1    g0069(.A(G274), .ZN(new_n270));
  OAI21_X1  g0070(.A(new_n261), .B1(G41), .B2(G45), .ZN(new_n271));
  NOR3_X1   g0071(.A1(new_n269), .A2(new_n270), .A3(new_n271), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n271), .A2(KEYINPUT66), .ZN(new_n273));
  NAND2_X1  g0073(.A1(G33), .A2(G41), .ZN(new_n274));
  NAND3_X1  g0074(.A1(new_n274), .A2(G1), .A3(G13), .ZN(new_n275));
  INV_X1    g0075(.A(KEYINPUT66), .ZN(new_n276));
  OAI211_X1 g0076(.A(new_n276), .B(new_n261), .C1(G41), .C2(G45), .ZN(new_n277));
  AND3_X1   g0077(.A1(new_n273), .A2(new_n275), .A3(new_n277), .ZN(new_n278));
  AOI21_X1  g0078(.A(new_n272), .B1(new_n278), .B2(G226), .ZN(new_n279));
  INV_X1    g0079(.A(KEYINPUT3), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n280), .A2(new_n256), .ZN(new_n281));
  NAND2_X1  g0081(.A1(KEYINPUT3), .A2(G33), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n281), .A2(new_n282), .ZN(new_n283));
  INV_X1    g0083(.A(G1698), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n283), .A2(new_n284), .ZN(new_n285));
  INV_X1    g0085(.A(G222), .ZN(new_n286));
  INV_X1    g0086(.A(G77), .ZN(new_n287));
  OAI22_X1  g0087(.A1(new_n285), .A2(new_n286), .B1(new_n287), .B2(new_n283), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n283), .A2(G1698), .ZN(new_n289));
  XNOR2_X1  g0089(.A(new_n289), .B(KEYINPUT67), .ZN(new_n290));
  AOI21_X1  g0090(.A(new_n288), .B1(new_n290), .B2(G223), .ZN(new_n291));
  OAI21_X1  g0091(.A(new_n279), .B1(new_n291), .B2(new_n275), .ZN(new_n292));
  NOR2_X1   g0092(.A1(new_n292), .A2(G179), .ZN(new_n293));
  INV_X1    g0093(.A(G169), .ZN(new_n294));
  AOI211_X1 g0094(.A(new_n268), .B(new_n293), .C1(new_n294), .C2(new_n292), .ZN(new_n295));
  INV_X1    g0095(.A(new_n268), .ZN(new_n296));
  AND2_X1   g0096(.A1(new_n296), .A2(KEYINPUT9), .ZN(new_n297));
  NOR2_X1   g0097(.A1(new_n296), .A2(KEYINPUT9), .ZN(new_n298));
  NOR2_X1   g0098(.A1(new_n297), .A2(new_n298), .ZN(new_n299));
  INV_X1    g0099(.A(G190), .ZN(new_n300));
  NOR2_X1   g0100(.A1(new_n292), .A2(new_n300), .ZN(new_n301));
  NOR2_X1   g0101(.A1(new_n299), .A2(new_n301), .ZN(new_n302));
  INV_X1    g0102(.A(KEYINPUT10), .ZN(new_n303));
  INV_X1    g0103(.A(KEYINPUT70), .ZN(new_n304));
  AOI21_X1  g0104(.A(new_n304), .B1(new_n292), .B2(G200), .ZN(new_n305));
  INV_X1    g0105(.A(new_n305), .ZN(new_n306));
  NAND3_X1  g0106(.A1(new_n292), .A2(new_n304), .A3(G200), .ZN(new_n307));
  NAND4_X1  g0107(.A1(new_n302), .A2(new_n303), .A3(new_n306), .A4(new_n307), .ZN(new_n308));
  OAI221_X1 g0108(.A(new_n307), .B1(new_n300), .B2(new_n292), .C1(new_n297), .C2(new_n298), .ZN(new_n309));
  OAI21_X1  g0109(.A(KEYINPUT10), .B1(new_n309), .B2(new_n305), .ZN(new_n310));
  AOI21_X1  g0110(.A(new_n295), .B1(new_n308), .B2(new_n310), .ZN(new_n311));
  AOI22_X1  g0111(.A1(new_n258), .A2(G50), .B1(G20), .B2(new_n217), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n227), .A2(G33), .ZN(new_n313));
  OAI21_X1  g0113(.A(new_n312), .B1(new_n287), .B2(new_n313), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n314), .A2(new_n248), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n315), .A2(KEYINPUT11), .ZN(new_n316));
  INV_X1    g0116(.A(KEYINPUT11), .ZN(new_n317));
  NAND3_X1  g0117(.A1(new_n314), .A2(new_n317), .A3(new_n248), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n316), .A2(new_n318), .ZN(new_n319));
  NAND3_X1  g0119(.A1(new_n264), .A2(G68), .A3(new_n265), .ZN(new_n320));
  OAI22_X1  g0120(.A1(new_n262), .A2(G68), .B1(KEYINPUT71), .B2(KEYINPUT12), .ZN(new_n321));
  NAND2_X1  g0121(.A1(KEYINPUT71), .A2(KEYINPUT12), .ZN(new_n322));
  XNOR2_X1  g0122(.A(new_n321), .B(new_n322), .ZN(new_n323));
  NAND3_X1  g0123(.A1(new_n319), .A2(new_n320), .A3(new_n323), .ZN(new_n324));
  NAND2_X1  g0124(.A1(G33), .A2(G97), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n232), .A2(G1698), .ZN(new_n326));
  OAI21_X1  g0126(.A(new_n326), .B1(G226), .B2(G1698), .ZN(new_n327));
  AND2_X1   g0127(.A1(KEYINPUT3), .A2(G33), .ZN(new_n328));
  NOR2_X1   g0128(.A1(KEYINPUT3), .A2(G33), .ZN(new_n329));
  NOR2_X1   g0129(.A1(new_n328), .A2(new_n329), .ZN(new_n330));
  OAI21_X1  g0130(.A(new_n325), .B1(new_n327), .B2(new_n330), .ZN(new_n331));
  AOI21_X1  g0131(.A(new_n272), .B1(new_n331), .B2(new_n269), .ZN(new_n332));
  INV_X1    g0132(.A(KEYINPUT13), .ZN(new_n333));
  NAND4_X1  g0133(.A1(new_n273), .A2(G238), .A3(new_n275), .A4(new_n277), .ZN(new_n334));
  NAND3_X1  g0134(.A1(new_n332), .A2(new_n333), .A3(new_n334), .ZN(new_n335));
  INV_X1    g0135(.A(new_n228), .ZN(new_n336));
  AOI21_X1  g0136(.A(new_n270), .B1(new_n336), .B2(new_n274), .ZN(new_n337));
  INV_X1    g0137(.A(new_n271), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n337), .A2(new_n338), .ZN(new_n339));
  NOR2_X1   g0139(.A1(G226), .A2(G1698), .ZN(new_n340));
  AOI21_X1  g0140(.A(new_n340), .B1(new_n232), .B2(G1698), .ZN(new_n341));
  AOI22_X1  g0141(.A1(new_n341), .A2(new_n283), .B1(G33), .B2(G97), .ZN(new_n342));
  OAI211_X1 g0142(.A(new_n339), .B(new_n334), .C1(new_n342), .C2(new_n275), .ZN(new_n343));
  NAND2_X1  g0143(.A1(new_n343), .A2(KEYINPUT13), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n335), .A2(new_n344), .ZN(new_n345));
  INV_X1    g0145(.A(KEYINPUT14), .ZN(new_n346));
  NAND3_X1  g0146(.A1(new_n345), .A2(new_n346), .A3(G169), .ZN(new_n347));
  NAND3_X1  g0147(.A1(new_n335), .A2(new_n344), .A3(G179), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n347), .A2(new_n348), .ZN(new_n349));
  AOI21_X1  g0149(.A(new_n346), .B1(new_n345), .B2(G169), .ZN(new_n350));
  OAI21_X1  g0150(.A(new_n324), .B1(new_n349), .B2(new_n350), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n345), .A2(G200), .ZN(new_n352));
  INV_X1    g0152(.A(new_n324), .ZN(new_n353));
  NAND3_X1  g0153(.A1(new_n335), .A2(new_n344), .A3(G190), .ZN(new_n354));
  NAND3_X1  g0154(.A1(new_n352), .A2(new_n353), .A3(new_n354), .ZN(new_n355));
  AND2_X1   g0155(.A1(new_n351), .A2(new_n355), .ZN(new_n356));
  INV_X1    g0156(.A(KEYINPUT18), .ZN(new_n357));
  INV_X1    g0157(.A(KEYINPUT16), .ZN(new_n358));
  NAND3_X1  g0158(.A1(new_n281), .A2(new_n227), .A3(new_n282), .ZN(new_n359));
  INV_X1    g0159(.A(KEYINPUT7), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n359), .A2(new_n360), .ZN(new_n361));
  NAND4_X1  g0161(.A1(new_n281), .A2(KEYINPUT7), .A3(new_n227), .A4(new_n282), .ZN(new_n362));
  AOI21_X1  g0162(.A(new_n217), .B1(new_n361), .B2(new_n362), .ZN(new_n363));
  INV_X1    g0163(.A(G58), .ZN(new_n364));
  NOR2_X1   g0164(.A1(new_n364), .A2(new_n217), .ZN(new_n365));
  OAI21_X1  g0165(.A(G20), .B1(new_n365), .B2(new_n201), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n258), .A2(G159), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n366), .A2(new_n367), .ZN(new_n368));
  OAI21_X1  g0168(.A(new_n358), .B1(new_n363), .B2(new_n368), .ZN(new_n369));
  AOI21_X1  g0169(.A(KEYINPUT7), .B1(new_n330), .B2(new_n227), .ZN(new_n370));
  INV_X1    g0170(.A(new_n362), .ZN(new_n371));
  OAI21_X1  g0171(.A(G68), .B1(new_n370), .B2(new_n371), .ZN(new_n372));
  INV_X1    g0172(.A(new_n368), .ZN(new_n373));
  NAND3_X1  g0173(.A1(new_n372), .A2(KEYINPUT16), .A3(new_n373), .ZN(new_n374));
  NAND3_X1  g0174(.A1(new_n369), .A2(new_n374), .A3(new_n248), .ZN(new_n375));
  AOI21_X1  g0175(.A(new_n254), .B1(new_n261), .B2(G20), .ZN(new_n376));
  AOI22_X1  g0176(.A1(new_n376), .A2(new_n264), .B1(new_n254), .B2(new_n263), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n375), .A2(new_n377), .ZN(new_n378));
  NOR2_X1   g0178(.A1(G223), .A2(G1698), .ZN(new_n379));
  INV_X1    g0179(.A(G226), .ZN(new_n380));
  AOI21_X1  g0180(.A(new_n379), .B1(new_n380), .B2(G1698), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n381), .A2(new_n283), .ZN(new_n382));
  NAND2_X1  g0182(.A1(G33), .A2(G87), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n382), .A2(new_n383), .ZN(new_n384));
  NAND2_X1  g0184(.A1(new_n384), .A2(new_n269), .ZN(new_n385));
  NAND4_X1  g0185(.A1(new_n273), .A2(G232), .A3(new_n275), .A4(new_n277), .ZN(new_n386));
  NAND4_X1  g0186(.A1(new_n385), .A2(G179), .A3(new_n339), .A4(new_n386), .ZN(new_n387));
  AOI22_X1  g0187(.A1(new_n381), .A2(new_n283), .B1(G33), .B2(G87), .ZN(new_n388));
  OAI211_X1 g0188(.A(new_n339), .B(new_n386), .C1(new_n388), .C2(new_n275), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n389), .A2(G169), .ZN(new_n390));
  NAND2_X1  g0190(.A1(new_n387), .A2(new_n390), .ZN(new_n391));
  AOI21_X1  g0191(.A(new_n357), .B1(new_n378), .B2(new_n391), .ZN(new_n392));
  INV_X1    g0192(.A(new_n392), .ZN(new_n393));
  NAND3_X1  g0193(.A1(new_n378), .A2(new_n357), .A3(new_n391), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n393), .A2(new_n394), .ZN(new_n395));
  NAND4_X1  g0195(.A1(new_n385), .A2(G190), .A3(new_n339), .A4(new_n386), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n389), .A2(G200), .ZN(new_n397));
  NAND4_X1  g0197(.A1(new_n375), .A2(new_n377), .A3(new_n396), .A4(new_n397), .ZN(new_n398));
  INV_X1    g0198(.A(KEYINPUT17), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n398), .A2(new_n399), .ZN(new_n400));
  AND2_X1   g0200(.A1(new_n396), .A2(new_n397), .ZN(new_n401));
  NAND4_X1  g0201(.A1(new_n401), .A2(KEYINPUT17), .A3(new_n375), .A4(new_n377), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n400), .A2(new_n402), .ZN(new_n403));
  NOR2_X1   g0203(.A1(new_n395), .A2(new_n403), .ZN(new_n404));
  INV_X1    g0204(.A(KEYINPUT69), .ZN(new_n405));
  INV_X1    g0205(.A(new_n258), .ZN(new_n406));
  AOI21_X1  g0206(.A(new_n254), .B1(new_n405), .B2(new_n406), .ZN(new_n407));
  OAI21_X1  g0207(.A(new_n407), .B1(new_n405), .B2(new_n406), .ZN(new_n408));
  XNOR2_X1  g0208(.A(KEYINPUT15), .B(G87), .ZN(new_n409));
  INV_X1    g0209(.A(new_n409), .ZN(new_n410));
  AOI22_X1  g0210(.A1(new_n410), .A2(new_n257), .B1(G20), .B2(G77), .ZN(new_n411));
  AOI21_X1  g0211(.A(new_n249), .B1(new_n408), .B2(new_n411), .ZN(new_n412));
  NAND3_X1  g0212(.A1(new_n264), .A2(G77), .A3(new_n265), .ZN(new_n413));
  OAI21_X1  g0213(.A(new_n413), .B1(G77), .B2(new_n262), .ZN(new_n414));
  NOR2_X1   g0214(.A1(new_n412), .A2(new_n414), .ZN(new_n415));
  OAI22_X1  g0215(.A1(new_n285), .A2(new_n232), .B1(new_n205), .B2(new_n283), .ZN(new_n416));
  INV_X1    g0216(.A(new_n216), .ZN(new_n417));
  AOI21_X1  g0217(.A(new_n416), .B1(new_n290), .B2(new_n417), .ZN(new_n418));
  OR2_X1    g0218(.A1(new_n418), .A2(new_n275), .ZN(new_n419));
  AOI21_X1  g0219(.A(new_n272), .B1(new_n278), .B2(G244), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n419), .A2(new_n420), .ZN(new_n421));
  AOI21_X1  g0221(.A(new_n415), .B1(new_n421), .B2(new_n294), .ZN(new_n422));
  INV_X1    g0222(.A(G179), .ZN(new_n423));
  NAND3_X1  g0223(.A1(new_n419), .A2(new_n423), .A3(new_n420), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n422), .A2(new_n424), .ZN(new_n425));
  INV_X1    g0225(.A(new_n425), .ZN(new_n426));
  INV_X1    g0226(.A(G200), .ZN(new_n427));
  AOI21_X1  g0227(.A(new_n427), .B1(new_n419), .B2(new_n420), .ZN(new_n428));
  OAI211_X1 g0228(.A(G190), .B(new_n420), .C1(new_n418), .C2(new_n275), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n429), .A2(new_n415), .ZN(new_n430));
  NOR2_X1   g0230(.A1(new_n428), .A2(new_n430), .ZN(new_n431));
  NOR2_X1   g0231(.A1(new_n426), .A2(new_n431), .ZN(new_n432));
  AND4_X1   g0232(.A1(new_n311), .A2(new_n356), .A3(new_n404), .A4(new_n432), .ZN(new_n433));
  INV_X1    g0233(.A(new_n433), .ZN(new_n434));
  INV_X1    g0234(.A(KEYINPUT81), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n261), .A2(G33), .ZN(new_n436));
  AND3_X1   g0236(.A1(new_n249), .A2(new_n262), .A3(new_n436), .ZN(new_n437));
  INV_X1    g0237(.A(KEYINPUT25), .ZN(new_n438));
  NOR3_X1   g0238(.A1(new_n262), .A2(new_n438), .A3(G107), .ZN(new_n439));
  INV_X1    g0239(.A(new_n439), .ZN(new_n440));
  OAI21_X1  g0240(.A(new_n438), .B1(new_n262), .B2(G107), .ZN(new_n441));
  AOI22_X1  g0241(.A1(new_n437), .A2(G107), .B1(new_n440), .B2(new_n441), .ZN(new_n442));
  INV_X1    g0242(.A(new_n442), .ZN(new_n443));
  INV_X1    g0243(.A(KEYINPUT24), .ZN(new_n444));
  OAI21_X1  g0244(.A(KEYINPUT23), .B1(new_n227), .B2(G107), .ZN(new_n445));
  INV_X1    g0245(.A(KEYINPUT23), .ZN(new_n446));
  NAND3_X1  g0246(.A1(new_n446), .A2(new_n205), .A3(G20), .ZN(new_n447));
  INV_X1    g0247(.A(G116), .ZN(new_n448));
  OAI211_X1 g0248(.A(new_n445), .B(new_n447), .C1(new_n448), .C2(new_n313), .ZN(new_n449));
  INV_X1    g0249(.A(KEYINPUT80), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n449), .A2(new_n450), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n257), .A2(G116), .ZN(new_n452));
  NAND4_X1  g0252(.A1(new_n452), .A2(KEYINPUT80), .A3(new_n447), .A4(new_n445), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n451), .A2(new_n453), .ZN(new_n454));
  OAI211_X1 g0254(.A(new_n227), .B(G87), .C1(new_n328), .C2(new_n329), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n455), .A2(KEYINPUT22), .ZN(new_n456));
  INV_X1    g0256(.A(KEYINPUT22), .ZN(new_n457));
  NAND4_X1  g0257(.A1(new_n283), .A2(new_n457), .A3(new_n227), .A4(G87), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n456), .A2(new_n458), .ZN(new_n459));
  AOI21_X1  g0259(.A(new_n444), .B1(new_n454), .B2(new_n459), .ZN(new_n460));
  INV_X1    g0260(.A(new_n460), .ZN(new_n461));
  NAND3_X1  g0261(.A1(new_n454), .A2(new_n444), .A3(new_n459), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  AOI21_X1  g0263(.A(new_n443), .B1(new_n463), .B2(new_n248), .ZN(new_n464));
  OAI211_X1 g0264(.A(G257), .B(G1698), .C1(new_n328), .C2(new_n329), .ZN(new_n465));
  OAI211_X1 g0265(.A(G250), .B(new_n284), .C1(new_n328), .C2(new_n329), .ZN(new_n466));
  INV_X1    g0266(.A(G294), .ZN(new_n467));
  OAI211_X1 g0267(.A(new_n465), .B(new_n466), .C1(new_n256), .C2(new_n467), .ZN(new_n468));
  NAND2_X1  g0268(.A1(new_n261), .A2(G45), .ZN(new_n469));
  INV_X1    g0269(.A(KEYINPUT5), .ZN(new_n470));
  NOR2_X1   g0270(.A1(new_n470), .A2(G41), .ZN(new_n471));
  INV_X1    g0271(.A(KEYINPUT75), .ZN(new_n472));
  AOI21_X1  g0272(.A(new_n469), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  INV_X1    g0273(.A(G41), .ZN(new_n474));
  OAI21_X1  g0274(.A(new_n472), .B1(new_n474), .B2(KEYINPUT5), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n474), .A2(KEYINPUT5), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n475), .A2(new_n476), .ZN(new_n477));
  AOI21_X1  g0277(.A(new_n269), .B1(new_n473), .B2(new_n477), .ZN(new_n478));
  AOI22_X1  g0278(.A1(new_n269), .A2(new_n468), .B1(new_n478), .B2(G264), .ZN(new_n479));
  NAND3_X1  g0279(.A1(new_n473), .A2(new_n337), .A3(new_n477), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n479), .A2(new_n480), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n481), .A2(new_n294), .ZN(new_n482));
  OAI21_X1  g0282(.A(new_n482), .B1(G179), .B2(new_n481), .ZN(new_n483));
  OAI21_X1  g0283(.A(new_n435), .B1(new_n464), .B2(new_n483), .ZN(new_n484));
  AOI22_X1  g0284(.A1(new_n247), .A2(new_n228), .B1(G20), .B2(new_n448), .ZN(new_n485));
  NAND2_X1  g0285(.A1(G33), .A2(G283), .ZN(new_n486));
  OAI211_X1 g0286(.A(new_n486), .B(new_n227), .C1(G33), .C2(new_n204), .ZN(new_n487));
  NAND3_X1  g0287(.A1(new_n485), .A2(KEYINPUT20), .A3(new_n487), .ZN(new_n488));
  INV_X1    g0288(.A(KEYINPUT77), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  AOI21_X1  g0290(.A(KEYINPUT20), .B1(new_n485), .B2(new_n487), .ZN(new_n491));
  INV_X1    g0291(.A(new_n491), .ZN(new_n492));
  NAND4_X1  g0292(.A1(new_n485), .A2(KEYINPUT77), .A3(new_n487), .A4(KEYINPUT20), .ZN(new_n493));
  NAND3_X1  g0293(.A1(new_n490), .A2(new_n492), .A3(new_n493), .ZN(new_n494));
  NAND3_X1  g0294(.A1(new_n249), .A2(new_n262), .A3(new_n436), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n495), .A2(G116), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n262), .A2(new_n448), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n494), .A2(new_n498), .ZN(new_n499));
  OAI211_X1 g0299(.A(G264), .B(G1698), .C1(new_n328), .C2(new_n329), .ZN(new_n500));
  OAI211_X1 g0300(.A(G257), .B(new_n284), .C1(new_n328), .C2(new_n329), .ZN(new_n501));
  INV_X1    g0301(.A(G303), .ZN(new_n502));
  OAI211_X1 g0302(.A(new_n500), .B(new_n501), .C1(new_n502), .C2(new_n283), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n503), .A2(new_n269), .ZN(new_n504));
  AOI21_X1  g0304(.A(KEYINPUT75), .B1(new_n470), .B2(G41), .ZN(new_n505));
  NOR2_X1   g0305(.A1(new_n505), .A2(new_n471), .ZN(new_n506));
  INV_X1    g0306(.A(G45), .ZN(new_n507));
  NOR2_X1   g0307(.A1(new_n507), .A2(G1), .ZN(new_n508));
  OAI21_X1  g0308(.A(new_n508), .B1(new_n476), .B2(KEYINPUT75), .ZN(new_n509));
  OAI211_X1 g0309(.A(G270), .B(new_n275), .C1(new_n506), .C2(new_n509), .ZN(new_n510));
  NAND3_X1  g0310(.A1(new_n504), .A2(new_n480), .A3(new_n510), .ZN(new_n511));
  NAND4_X1  g0311(.A1(new_n499), .A2(new_n511), .A3(KEYINPUT21), .A4(G169), .ZN(new_n512));
  INV_X1    g0312(.A(KEYINPUT78), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  AND2_X1   g0314(.A1(new_n510), .A2(new_n480), .ZN(new_n515));
  AOI21_X1  g0315(.A(new_n294), .B1(new_n515), .B2(new_n504), .ZN(new_n516));
  NAND4_X1  g0316(.A1(new_n516), .A2(KEYINPUT78), .A3(KEYINPUT21), .A4(new_n499), .ZN(new_n517));
  NOR2_X1   g0317(.A1(new_n511), .A2(new_n423), .ZN(new_n518));
  AOI22_X1  g0318(.A1(new_n514), .A2(new_n517), .B1(new_n499), .B2(new_n518), .ZN(new_n519));
  AOI21_X1  g0319(.A(G169), .B1(new_n479), .B2(new_n480), .ZN(new_n520));
  INV_X1    g0320(.A(new_n481), .ZN(new_n521));
  AOI21_X1  g0321(.A(new_n520), .B1(new_n521), .B2(new_n423), .ZN(new_n522));
  AND3_X1   g0322(.A1(new_n454), .A2(new_n444), .A3(new_n459), .ZN(new_n523));
  OAI21_X1  g0323(.A(new_n248), .B1(new_n523), .B2(new_n460), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n524), .A2(new_n442), .ZN(new_n525));
  NAND3_X1  g0325(.A1(new_n522), .A2(new_n525), .A3(KEYINPUT81), .ZN(new_n526));
  INV_X1    g0326(.A(KEYINPUT79), .ZN(new_n527));
  AND2_X1   g0327(.A1(new_n503), .A2(new_n269), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n510), .A2(new_n480), .ZN(new_n529));
  OAI21_X1  g0329(.A(G169), .B1(new_n528), .B2(new_n529), .ZN(new_n530));
  AOI21_X1  g0330(.A(new_n491), .B1(new_n489), .B2(new_n488), .ZN(new_n531));
  AOI22_X1  g0331(.A1(new_n531), .A2(new_n493), .B1(new_n496), .B2(new_n497), .ZN(new_n532));
  OAI21_X1  g0332(.A(new_n527), .B1(new_n530), .B2(new_n532), .ZN(new_n533));
  INV_X1    g0333(.A(KEYINPUT21), .ZN(new_n534));
  NAND4_X1  g0334(.A1(new_n499), .A2(new_n511), .A3(KEYINPUT79), .A4(G169), .ZN(new_n535));
  NAND3_X1  g0335(.A1(new_n533), .A2(new_n534), .A3(new_n535), .ZN(new_n536));
  NAND4_X1  g0336(.A1(new_n484), .A2(new_n519), .A3(new_n526), .A4(new_n536), .ZN(new_n537));
  NOR2_X1   g0337(.A1(new_n262), .A2(G97), .ZN(new_n538));
  AOI21_X1  g0338(.A(new_n538), .B1(new_n437), .B2(G97), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n258), .A2(G77), .ZN(new_n540));
  INV_X1    g0340(.A(KEYINPUT6), .ZN(new_n541));
  NAND2_X1  g0341(.A1(new_n541), .A2(KEYINPUT72), .ZN(new_n542));
  INV_X1    g0342(.A(KEYINPUT72), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n543), .A2(KEYINPUT6), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n542), .A2(new_n544), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n205), .A2(G97), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n545), .A2(new_n546), .ZN(new_n547));
  NAND2_X1  g0347(.A1(G97), .A2(G107), .ZN(new_n548));
  NAND4_X1  g0348(.A1(new_n206), .A2(new_n542), .A3(new_n544), .A4(new_n548), .ZN(new_n549));
  NAND3_X1  g0349(.A1(new_n547), .A2(G20), .A3(new_n549), .ZN(new_n550));
  AOI21_X1  g0350(.A(new_n205), .B1(new_n361), .B2(new_n362), .ZN(new_n551));
  INV_X1    g0351(.A(KEYINPUT73), .ZN(new_n552));
  OAI211_X1 g0352(.A(new_n540), .B(new_n550), .C1(new_n551), .C2(new_n552), .ZN(new_n553));
  OAI21_X1  g0353(.A(G107), .B1(new_n370), .B2(new_n371), .ZN(new_n554));
  NOR2_X1   g0354(.A1(new_n554), .A2(KEYINPUT73), .ZN(new_n555));
  OAI211_X1 g0355(.A(KEYINPUT74), .B(new_n248), .C1(new_n553), .C2(new_n555), .ZN(new_n556));
  INV_X1    g0356(.A(new_n556), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n554), .A2(KEYINPUT73), .ZN(new_n558));
  AND2_X1   g0358(.A1(new_n550), .A2(new_n540), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n551), .A2(new_n552), .ZN(new_n560));
  NAND3_X1  g0360(.A1(new_n558), .A2(new_n559), .A3(new_n560), .ZN(new_n561));
  AOI21_X1  g0361(.A(KEYINPUT74), .B1(new_n561), .B2(new_n248), .ZN(new_n562));
  OAI21_X1  g0362(.A(new_n539), .B1(new_n557), .B2(new_n562), .ZN(new_n563));
  NAND3_X1  g0363(.A1(new_n283), .A2(G250), .A3(G1698), .ZN(new_n564));
  NAND3_X1  g0364(.A1(new_n283), .A2(G244), .A3(new_n284), .ZN(new_n565));
  INV_X1    g0365(.A(KEYINPUT4), .ZN(new_n566));
  OAI211_X1 g0366(.A(new_n486), .B(new_n564), .C1(new_n565), .C2(new_n566), .ZN(new_n567));
  NOR2_X1   g0367(.A1(new_n330), .A2(G1698), .ZN(new_n568));
  AOI21_X1  g0368(.A(KEYINPUT4), .B1(new_n568), .B2(G244), .ZN(new_n569));
  OAI21_X1  g0369(.A(new_n269), .B1(new_n567), .B2(new_n569), .ZN(new_n570));
  NOR2_X1   g0370(.A1(new_n506), .A2(new_n509), .ZN(new_n571));
  AOI22_X1  g0371(.A1(new_n478), .A2(G257), .B1(new_n571), .B2(new_n337), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n570), .A2(new_n572), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n573), .A2(G169), .ZN(new_n574));
  OAI21_X1  g0374(.A(new_n574), .B1(new_n423), .B2(new_n573), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n563), .A2(new_n575), .ZN(new_n576));
  OAI211_X1 g0376(.A(G244), .B(G1698), .C1(new_n328), .C2(new_n329), .ZN(new_n577));
  OAI211_X1 g0377(.A(G238), .B(new_n284), .C1(new_n328), .C2(new_n329), .ZN(new_n578));
  OAI211_X1 g0378(.A(new_n577), .B(new_n578), .C1(new_n256), .C2(new_n448), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n579), .A2(new_n269), .ZN(new_n580));
  INV_X1    g0380(.A(KEYINPUT76), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n508), .A2(new_n581), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n469), .A2(KEYINPUT76), .ZN(new_n583));
  NAND4_X1  g0383(.A1(new_n582), .A2(new_n583), .A3(G250), .A4(new_n275), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n337), .A2(new_n508), .ZN(new_n585));
  AND2_X1   g0385(.A1(new_n584), .A2(new_n585), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n580), .A2(new_n586), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n587), .A2(G200), .ZN(new_n588));
  INV_X1    g0388(.A(KEYINPUT19), .ZN(new_n589));
  OAI21_X1  g0389(.A(new_n227), .B1(new_n325), .B2(new_n589), .ZN(new_n590));
  OAI21_X1  g0390(.A(new_n590), .B1(G87), .B2(new_n206), .ZN(new_n591));
  OAI211_X1 g0391(.A(new_n227), .B(G68), .C1(new_n328), .C2(new_n329), .ZN(new_n592));
  OAI21_X1  g0392(.A(new_n589), .B1(new_n313), .B2(new_n204), .ZN(new_n593));
  NAND3_X1  g0393(.A1(new_n591), .A2(new_n592), .A3(new_n593), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n594), .A2(new_n248), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n409), .A2(new_n263), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n437), .A2(G87), .ZN(new_n597));
  AND3_X1   g0397(.A1(new_n595), .A2(new_n596), .A3(new_n597), .ZN(new_n598));
  NAND3_X1  g0398(.A1(new_n580), .A2(new_n586), .A3(G190), .ZN(new_n599));
  NAND3_X1  g0399(.A1(new_n588), .A2(new_n598), .A3(new_n599), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n437), .A2(new_n410), .ZN(new_n601));
  NAND3_X1  g0401(.A1(new_n595), .A2(new_n601), .A3(new_n596), .ZN(new_n602));
  NAND3_X1  g0402(.A1(new_n580), .A2(new_n586), .A3(new_n423), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n584), .A2(new_n585), .ZN(new_n604));
  AOI21_X1  g0404(.A(new_n604), .B1(new_n269), .B2(new_n579), .ZN(new_n605));
  OAI211_X1 g0405(.A(new_n602), .B(new_n603), .C1(new_n605), .C2(G169), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n600), .A2(new_n606), .ZN(new_n607));
  AOI21_X1  g0407(.A(new_n427), .B1(new_n479), .B2(new_n480), .ZN(new_n608));
  AOI21_X1  g0408(.A(new_n608), .B1(new_n521), .B2(G190), .ZN(new_n609));
  AOI21_X1  g0409(.A(new_n607), .B1(new_n464), .B2(new_n609), .ZN(new_n610));
  AND3_X1   g0410(.A1(new_n570), .A2(G190), .A3(new_n572), .ZN(new_n611));
  AOI21_X1  g0411(.A(new_n427), .B1(new_n570), .B2(new_n572), .ZN(new_n612));
  NOR2_X1   g0412(.A1(new_n611), .A2(new_n612), .ZN(new_n613));
  OAI211_X1 g0413(.A(new_n613), .B(new_n539), .C1(new_n562), .C2(new_n557), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n511), .A2(G200), .ZN(new_n615));
  OAI211_X1 g0415(.A(new_n615), .B(new_n532), .C1(new_n300), .C2(new_n511), .ZN(new_n616));
  NAND4_X1  g0416(.A1(new_n576), .A2(new_n610), .A3(new_n614), .A4(new_n616), .ZN(new_n617));
  NOR3_X1   g0417(.A1(new_n434), .A2(new_n537), .A3(new_n617), .ZN(G372));
  AOI221_X4 g0418(.A(KEYINPUT18), .B1(new_n387), .B2(new_n390), .C1(new_n375), .C2(new_n377), .ZN(new_n619));
  NOR2_X1   g0419(.A1(new_n619), .A2(new_n392), .ZN(new_n620));
  INV_X1    g0420(.A(new_n351), .ZN(new_n621));
  AOI21_X1  g0421(.A(new_n621), .B1(new_n426), .B2(new_n355), .ZN(new_n622));
  OAI21_X1  g0422(.A(new_n620), .B1(new_n622), .B2(new_n403), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n308), .A2(new_n310), .ZN(new_n624));
  AOI21_X1  g0424(.A(new_n295), .B1(new_n623), .B2(new_n624), .ZN(new_n625));
  AND2_X1   g0425(.A1(new_n600), .A2(new_n606), .ZN(new_n626));
  XNOR2_X1  g0426(.A(KEYINPUT84), .B(KEYINPUT26), .ZN(new_n627));
  INV_X1    g0427(.A(new_n627), .ZN(new_n628));
  NAND4_X1  g0428(.A1(new_n563), .A2(new_n575), .A3(new_n626), .A4(new_n628), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n629), .A2(KEYINPUT83), .ZN(new_n630));
  NAND3_X1  g0430(.A1(new_n563), .A2(new_n575), .A3(new_n626), .ZN(new_n631));
  INV_X1    g0431(.A(KEYINPUT26), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n631), .A2(new_n632), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n630), .A2(new_n633), .ZN(new_n634));
  NAND3_X1  g0434(.A1(new_n631), .A2(KEYINPUT83), .A3(new_n632), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  INV_X1    g0436(.A(new_n606), .ZN(new_n637));
  AND3_X1   g0437(.A1(new_n576), .A2(new_n614), .A3(new_n610), .ZN(new_n638));
  INV_X1    g0438(.A(KEYINPUT82), .ZN(new_n639));
  AND3_X1   g0439(.A1(new_n522), .A2(new_n525), .A3(new_n639), .ZN(new_n640));
  AOI21_X1  g0440(.A(new_n639), .B1(new_n522), .B2(new_n525), .ZN(new_n641));
  OAI211_X1 g0441(.A(new_n536), .B(new_n519), .C1(new_n640), .C2(new_n641), .ZN(new_n642));
  AOI21_X1  g0442(.A(new_n637), .B1(new_n638), .B2(new_n642), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n636), .A2(new_n643), .ZN(new_n644));
  INV_X1    g0444(.A(new_n644), .ZN(new_n645));
  OAI21_X1  g0445(.A(new_n625), .B1(new_n434), .B2(new_n645), .ZN(new_n646));
  XNOR2_X1  g0446(.A(new_n646), .B(KEYINPUT85), .ZN(G369));
  NAND3_X1  g0447(.A1(new_n261), .A2(new_n227), .A3(G13), .ZN(new_n648));
  OR2_X1    g0448(.A1(new_n648), .A2(KEYINPUT27), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n648), .A2(KEYINPUT27), .ZN(new_n650));
  AND3_X1   g0450(.A1(new_n649), .A2(G213), .A3(new_n650), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n651), .A2(G343), .ZN(new_n652));
  XNOR2_X1  g0452(.A(new_n652), .B(KEYINPUT86), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n525), .A2(new_n653), .ZN(new_n654));
  XNOR2_X1  g0454(.A(new_n654), .B(KEYINPUT87), .ZN(new_n655));
  AND2_X1   g0455(.A1(new_n484), .A2(new_n526), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n464), .A2(new_n609), .ZN(new_n657));
  AND3_X1   g0457(.A1(new_n655), .A2(new_n656), .A3(new_n657), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n522), .A2(new_n525), .ZN(new_n659));
  INV_X1    g0459(.A(new_n659), .ZN(new_n660));
  AOI21_X1  g0460(.A(new_n658), .B1(new_n660), .B2(new_n653), .ZN(new_n661));
  INV_X1    g0461(.A(new_n661), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n514), .A2(new_n517), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n518), .A2(new_n499), .ZN(new_n664));
  NAND3_X1  g0464(.A1(new_n663), .A2(new_n536), .A3(new_n664), .ZN(new_n665));
  INV_X1    g0465(.A(new_n653), .ZN(new_n666));
  NOR2_X1   g0466(.A1(new_n666), .A2(new_n532), .ZN(new_n667));
  XNOR2_X1  g0467(.A(new_n665), .B(new_n667), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n668), .A2(new_n616), .ZN(new_n669));
  INV_X1    g0469(.A(G330), .ZN(new_n670));
  NOR2_X1   g0470(.A1(new_n669), .A2(new_n670), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n662), .A2(new_n671), .ZN(new_n672));
  INV_X1    g0472(.A(new_n641), .ZN(new_n673));
  NAND3_X1  g0473(.A1(new_n522), .A2(new_n525), .A3(new_n639), .ZN(new_n674));
  NAND3_X1  g0474(.A1(new_n673), .A2(new_n674), .A3(new_n666), .ZN(new_n675));
  NAND3_X1  g0475(.A1(new_n655), .A2(new_n656), .A3(new_n657), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n665), .A2(new_n666), .ZN(new_n677));
  OAI21_X1  g0477(.A(new_n675), .B1(new_n676), .B2(new_n677), .ZN(new_n678));
  INV_X1    g0478(.A(new_n678), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n672), .A2(new_n679), .ZN(G399));
  INV_X1    g0480(.A(new_n213), .ZN(new_n681));
  NOR2_X1   g0481(.A1(new_n681), .A2(G41), .ZN(new_n682));
  INV_X1    g0482(.A(G87), .ZN(new_n683));
  NAND4_X1  g0483(.A1(new_n683), .A2(new_n204), .A3(new_n205), .A4(new_n448), .ZN(new_n684));
  NOR3_X1   g0484(.A1(new_n682), .A2(new_n261), .A3(new_n684), .ZN(new_n685));
  INV_X1    g0485(.A(new_n226), .ZN(new_n686));
  AOI21_X1  g0486(.A(new_n685), .B1(new_n686), .B2(new_n682), .ZN(new_n687));
  XOR2_X1   g0487(.A(new_n687), .B(KEYINPUT28), .Z(new_n688));
  AND2_X1   g0488(.A1(new_n638), .A2(new_n537), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n631), .A2(new_n628), .ZN(new_n690));
  OAI211_X1 g0490(.A(new_n690), .B(new_n606), .C1(KEYINPUT26), .C2(new_n631), .ZN(new_n691));
  OAI211_X1 g0491(.A(KEYINPUT29), .B(new_n666), .C1(new_n689), .C2(new_n691), .ZN(new_n692));
  AOI21_X1  g0492(.A(new_n653), .B1(new_n636), .B2(new_n643), .ZN(new_n693));
  OAI21_X1  g0493(.A(new_n692), .B1(new_n693), .B2(KEYINPUT29), .ZN(new_n694));
  INV_X1    g0494(.A(KEYINPUT30), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n468), .A2(new_n269), .ZN(new_n696));
  NAND2_X1  g0496(.A1(new_n478), .A2(G264), .ZN(new_n697));
  AND4_X1   g0497(.A1(new_n696), .A2(new_n580), .A3(new_n586), .A4(new_n697), .ZN(new_n698));
  NAND4_X1  g0498(.A1(new_n518), .A2(new_n698), .A3(new_n570), .A4(new_n572), .ZN(new_n699));
  AND2_X1   g0499(.A1(new_n573), .A2(new_n481), .ZN(new_n700));
  AND3_X1   g0500(.A1(new_n511), .A2(new_n423), .A3(new_n587), .ZN(new_n701));
  AOI22_X1  g0501(.A1(new_n695), .A2(new_n699), .B1(new_n700), .B2(new_n701), .ZN(new_n702));
  OR2_X1    g0502(.A1(new_n699), .A2(new_n695), .ZN(new_n703));
  AOI21_X1  g0503(.A(new_n666), .B1(new_n702), .B2(new_n703), .ZN(new_n704));
  OAI21_X1  g0504(.A(KEYINPUT88), .B1(new_n704), .B2(KEYINPUT31), .ZN(new_n705));
  NAND2_X1  g0505(.A1(new_n699), .A2(new_n695), .ZN(new_n706));
  NAND2_X1  g0506(.A1(new_n700), .A2(new_n701), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  NOR2_X1   g0508(.A1(new_n699), .A2(new_n695), .ZN(new_n709));
  OAI21_X1  g0509(.A(new_n653), .B1(new_n708), .B2(new_n709), .ZN(new_n710));
  INV_X1    g0510(.A(KEYINPUT88), .ZN(new_n711));
  INV_X1    g0511(.A(KEYINPUT31), .ZN(new_n712));
  NAND3_X1  g0512(.A1(new_n710), .A2(new_n711), .A3(new_n712), .ZN(new_n713));
  NAND2_X1  g0513(.A1(new_n704), .A2(KEYINPUT31), .ZN(new_n714));
  NAND3_X1  g0514(.A1(new_n705), .A2(new_n713), .A3(new_n714), .ZN(new_n715));
  NOR3_X1   g0515(.A1(new_n617), .A2(new_n537), .A3(new_n653), .ZN(new_n716));
  OAI21_X1  g0516(.A(G330), .B1(new_n715), .B2(new_n716), .ZN(new_n717));
  NAND2_X1  g0517(.A1(new_n694), .A2(new_n717), .ZN(new_n718));
  INV_X1    g0518(.A(new_n718), .ZN(new_n719));
  OAI21_X1  g0519(.A(new_n688), .B1(new_n719), .B2(G1), .ZN(G364));
  NAND2_X1  g0520(.A1(new_n669), .A2(new_n670), .ZN(new_n721));
  XNOR2_X1  g0521(.A(new_n721), .B(KEYINPUT89), .ZN(new_n722));
  INV_X1    g0522(.A(new_n682), .ZN(new_n723));
  NOR2_X1   g0523(.A1(new_n211), .A2(G20), .ZN(new_n724));
  AOI21_X1  g0524(.A(new_n261), .B1(new_n724), .B2(G45), .ZN(new_n725));
  AOI211_X1 g0525(.A(new_n671), .B(new_n722), .C1(new_n723), .C2(new_n725), .ZN(new_n726));
  INV_X1    g0526(.A(new_n725), .ZN(new_n727));
  NOR2_X1   g0527(.A1(new_n682), .A2(new_n727), .ZN(new_n728));
  INV_X1    g0528(.A(new_n728), .ZN(new_n729));
  AOI21_X1  g0529(.A(new_n228), .B1(G20), .B2(new_n294), .ZN(new_n730));
  INV_X1    g0530(.A(new_n730), .ZN(new_n731));
  NOR2_X1   g0531(.A1(new_n227), .A2(new_n423), .ZN(new_n732));
  NOR2_X1   g0532(.A1(G190), .A2(G200), .ZN(new_n733));
  NAND2_X1  g0533(.A1(new_n732), .A2(new_n733), .ZN(new_n734));
  INV_X1    g0534(.A(G311), .ZN(new_n735));
  NAND3_X1  g0535(.A1(new_n732), .A2(new_n300), .A3(G200), .ZN(new_n736));
  XOR2_X1   g0536(.A(KEYINPUT33), .B(G317), .Z(new_n737));
  OAI221_X1 g0537(.A(new_n330), .B1(new_n734), .B2(new_n735), .C1(new_n736), .C2(new_n737), .ZN(new_n738));
  NAND2_X1  g0538(.A1(new_n732), .A2(G190), .ZN(new_n739));
  NOR2_X1   g0539(.A1(new_n739), .A2(G200), .ZN(new_n740));
  NOR2_X1   g0540(.A1(new_n227), .A2(G179), .ZN(new_n741));
  NAND3_X1  g0541(.A1(new_n741), .A2(G190), .A3(G200), .ZN(new_n742));
  INV_X1    g0542(.A(new_n742), .ZN(new_n743));
  AOI22_X1  g0543(.A1(new_n740), .A2(G322), .B1(new_n743), .B2(G303), .ZN(new_n744));
  NOR2_X1   g0544(.A1(new_n739), .A2(new_n427), .ZN(new_n745));
  NAND3_X1  g0545(.A1(new_n741), .A2(new_n300), .A3(G200), .ZN(new_n746));
  INV_X1    g0546(.A(new_n746), .ZN(new_n747));
  AOI22_X1  g0547(.A1(new_n745), .A2(G326), .B1(new_n747), .B2(G283), .ZN(new_n748));
  NAND2_X1  g0548(.A1(new_n744), .A2(new_n748), .ZN(new_n749));
  OR3_X1    g0549(.A1(KEYINPUT91), .A2(G179), .A3(G200), .ZN(new_n750));
  OAI21_X1  g0550(.A(KEYINPUT91), .B1(G179), .B2(G200), .ZN(new_n751));
  NAND2_X1  g0551(.A1(new_n750), .A2(new_n751), .ZN(new_n752));
  NOR2_X1   g0552(.A1(new_n227), .A2(G190), .ZN(new_n753));
  AND2_X1   g0553(.A1(new_n752), .A2(new_n753), .ZN(new_n754));
  AOI211_X1 g0554(.A(new_n738), .B(new_n749), .C1(G329), .C2(new_n754), .ZN(new_n755));
  AOI21_X1  g0555(.A(new_n300), .B1(new_n750), .B2(new_n751), .ZN(new_n756));
  NOR2_X1   g0556(.A1(new_n756), .A2(new_n227), .ZN(new_n757));
  OAI21_X1  g0557(.A(new_n755), .B1(new_n467), .B2(new_n757), .ZN(new_n758));
  INV_X1    g0558(.A(new_n740), .ZN(new_n759));
  OAI22_X1  g0559(.A1(new_n759), .A2(new_n364), .B1(new_n742), .B2(new_n683), .ZN(new_n760));
  INV_X1    g0560(.A(new_n745), .ZN(new_n761));
  NOR2_X1   g0561(.A1(new_n761), .A2(new_n250), .ZN(new_n762));
  OAI221_X1 g0562(.A(new_n283), .B1(new_n734), .B2(new_n287), .C1(new_n217), .C2(new_n736), .ZN(new_n763));
  NOR2_X1   g0563(.A1(new_n746), .A2(new_n205), .ZN(new_n764));
  NOR4_X1   g0564(.A1(new_n760), .A2(new_n762), .A3(new_n763), .A4(new_n764), .ZN(new_n765));
  INV_X1    g0565(.A(new_n754), .ZN(new_n766));
  INV_X1    g0566(.A(G159), .ZN(new_n767));
  OR3_X1    g0567(.A1(new_n766), .A2(KEYINPUT32), .A3(new_n767), .ZN(new_n768));
  INV_X1    g0568(.A(new_n757), .ZN(new_n769));
  NAND2_X1  g0569(.A1(new_n769), .A2(G97), .ZN(new_n770));
  OAI21_X1  g0570(.A(KEYINPUT32), .B1(new_n766), .B2(new_n767), .ZN(new_n771));
  NAND4_X1  g0571(.A1(new_n765), .A2(new_n768), .A3(new_n770), .A4(new_n771), .ZN(new_n772));
  AOI21_X1  g0572(.A(new_n731), .B1(new_n758), .B2(new_n772), .ZN(new_n773));
  NOR2_X1   g0573(.A1(G13), .A2(G33), .ZN(new_n774));
  INV_X1    g0574(.A(new_n774), .ZN(new_n775));
  NOR2_X1   g0575(.A1(new_n775), .A2(G20), .ZN(new_n776));
  NOR2_X1   g0576(.A1(new_n776), .A2(new_n730), .ZN(new_n777));
  XOR2_X1   g0577(.A(new_n777), .B(KEYINPUT90), .Z(new_n778));
  NOR2_X1   g0578(.A1(new_n681), .A2(new_n330), .ZN(new_n779));
  AOI22_X1  g0579(.A1(new_n779), .A2(G355), .B1(new_n448), .B2(new_n681), .ZN(new_n780));
  AND2_X1   g0580(.A1(new_n245), .A2(G45), .ZN(new_n781));
  NOR2_X1   g0581(.A1(new_n681), .A2(new_n283), .ZN(new_n782));
  OAI21_X1  g0582(.A(new_n782), .B1(G45), .B2(new_n226), .ZN(new_n783));
  OAI21_X1  g0583(.A(new_n780), .B1(new_n781), .B2(new_n783), .ZN(new_n784));
  AOI211_X1 g0584(.A(new_n729), .B(new_n773), .C1(new_n778), .C2(new_n784), .ZN(new_n785));
  XOR2_X1   g0585(.A(new_n785), .B(KEYINPUT92), .Z(new_n786));
  AOI21_X1  g0586(.A(new_n786), .B1(new_n669), .B2(new_n776), .ZN(new_n787));
  NOR2_X1   g0587(.A1(new_n726), .A2(new_n787), .ZN(new_n788));
  INV_X1    g0588(.A(new_n788), .ZN(G396));
  OAI211_X1 g0589(.A(new_n425), .B(new_n666), .C1(new_n428), .C2(new_n430), .ZN(new_n790));
  INV_X1    g0590(.A(new_n790), .ZN(new_n791));
  AOI22_X1  g0591(.A1(KEYINPUT83), .A2(new_n629), .B1(new_n631), .B2(new_n632), .ZN(new_n792));
  AND3_X1   g0592(.A1(new_n631), .A2(KEYINPUT83), .A3(new_n632), .ZN(new_n793));
  NOR2_X1   g0593(.A1(new_n792), .A2(new_n793), .ZN(new_n794));
  AOI21_X1  g0594(.A(new_n665), .B1(new_n673), .B2(new_n674), .ZN(new_n795));
  NAND3_X1  g0595(.A1(new_n576), .A2(new_n610), .A3(new_n614), .ZN(new_n796));
  OAI21_X1  g0596(.A(new_n606), .B1(new_n795), .B2(new_n796), .ZN(new_n797));
  OAI21_X1  g0597(.A(new_n791), .B1(new_n794), .B2(new_n797), .ZN(new_n798));
  INV_X1    g0598(.A(new_n415), .ZN(new_n799));
  NOR2_X1   g0599(.A1(new_n418), .A2(new_n275), .ZN(new_n800));
  INV_X1    g0600(.A(new_n420), .ZN(new_n801));
  OAI21_X1  g0601(.A(new_n294), .B1(new_n800), .B2(new_n801), .ZN(new_n802));
  AND4_X1   g0602(.A1(new_n424), .A2(new_n799), .A3(new_n802), .A4(new_n666), .ZN(new_n803));
  OAI22_X1  g0603(.A1(new_n428), .A2(new_n430), .B1(new_n415), .B2(new_n666), .ZN(new_n804));
  AOI21_X1  g0604(.A(new_n803), .B1(new_n425), .B2(new_n804), .ZN(new_n805));
  OAI21_X1  g0605(.A(new_n798), .B1(new_n693), .B2(new_n805), .ZN(new_n806));
  AOI21_X1  g0606(.A(new_n728), .B1(new_n806), .B2(new_n717), .ZN(new_n807));
  OAI21_X1  g0607(.A(new_n807), .B1(new_n717), .B2(new_n806), .ZN(new_n808));
  NOR2_X1   g0608(.A1(new_n730), .A2(new_n774), .ZN(new_n809));
  AOI21_X1  g0609(.A(new_n729), .B1(new_n287), .B2(new_n809), .ZN(new_n810));
  INV_X1    g0610(.A(new_n736), .ZN(new_n811));
  INV_X1    g0611(.A(new_n734), .ZN(new_n812));
  AOI22_X1  g0612(.A1(new_n811), .A2(G150), .B1(new_n812), .B2(G159), .ZN(new_n813));
  INV_X1    g0613(.A(G143), .ZN(new_n814));
  INV_X1    g0614(.A(G137), .ZN(new_n815));
  OAI221_X1 g0615(.A(new_n813), .B1(new_n759), .B2(new_n814), .C1(new_n815), .C2(new_n761), .ZN(new_n816));
  XNOR2_X1  g0616(.A(new_n816), .B(KEYINPUT34), .ZN(new_n817));
  OAI221_X1 g0617(.A(new_n283), .B1(new_n742), .B2(new_n250), .C1(new_n217), .C2(new_n746), .ZN(new_n818));
  NOR2_X1   g0618(.A1(new_n757), .A2(new_n364), .ZN(new_n819));
  AOI211_X1 g0619(.A(new_n818), .B(new_n819), .C1(G132), .C2(new_n754), .ZN(new_n820));
  NOR2_X1   g0620(.A1(new_n766), .A2(new_n735), .ZN(new_n821));
  OAI22_X1  g0621(.A1(new_n759), .A2(new_n467), .B1(new_n742), .B2(new_n205), .ZN(new_n822));
  OAI22_X1  g0622(.A1(new_n761), .A2(new_n502), .B1(new_n746), .B2(new_n683), .ZN(new_n823));
  INV_X1    g0623(.A(G283), .ZN(new_n824));
  OAI221_X1 g0624(.A(new_n330), .B1(new_n734), .B2(new_n448), .C1(new_n824), .C2(new_n736), .ZN(new_n825));
  NOR4_X1   g0625(.A1(new_n821), .A2(new_n822), .A3(new_n823), .A4(new_n825), .ZN(new_n826));
  AOI22_X1  g0626(.A1(new_n817), .A2(new_n820), .B1(new_n770), .B2(new_n826), .ZN(new_n827));
  OAI221_X1 g0627(.A(new_n810), .B1(new_n731), .B2(new_n827), .C1(new_n805), .C2(new_n775), .ZN(new_n828));
  AND2_X1   g0628(.A1(new_n808), .A2(new_n828), .ZN(new_n829));
  INV_X1    g0629(.A(new_n829), .ZN(G384));
  NOR3_X1   g0630(.A1(new_n228), .A2(new_n227), .A3(new_n448), .ZN(new_n831));
  NAND2_X1  g0631(.A1(new_n547), .A2(new_n549), .ZN(new_n832));
  INV_X1    g0632(.A(KEYINPUT35), .ZN(new_n833));
  OAI21_X1  g0633(.A(new_n831), .B1(new_n832), .B2(new_n833), .ZN(new_n834));
  AOI21_X1  g0634(.A(new_n834), .B1(new_n833), .B2(new_n832), .ZN(new_n835));
  XNOR2_X1  g0635(.A(KEYINPUT93), .B(KEYINPUT36), .ZN(new_n836));
  XNOR2_X1  g0636(.A(new_n835), .B(new_n836), .ZN(new_n837));
  OR3_X1    g0637(.A1(new_n226), .A2(new_n287), .A3(new_n365), .ZN(new_n838));
  NAND2_X1  g0638(.A1(new_n250), .A2(G68), .ZN(new_n839));
  AOI211_X1 g0639(.A(new_n261), .B(G13), .C1(new_n838), .C2(new_n839), .ZN(new_n840));
  NOR2_X1   g0640(.A1(new_n837), .A2(new_n840), .ZN(new_n841));
  OAI211_X1 g0641(.A(new_n433), .B(new_n692), .C1(KEYINPUT29), .C2(new_n693), .ZN(new_n842));
  NAND2_X1  g0642(.A1(new_n842), .A2(new_n625), .ZN(new_n843));
  XNOR2_X1  g0643(.A(new_n843), .B(KEYINPUT99), .ZN(new_n844));
  INV_X1    g0644(.A(new_n377), .ZN(new_n845));
  AND2_X1   g0645(.A1(new_n374), .A2(new_n248), .ZN(new_n846));
  OAI21_X1  g0646(.A(KEYINPUT95), .B1(new_n363), .B2(new_n368), .ZN(new_n847));
  INV_X1    g0647(.A(KEYINPUT95), .ZN(new_n848));
  NAND3_X1  g0648(.A1(new_n372), .A2(new_n848), .A3(new_n373), .ZN(new_n849));
  NAND3_X1  g0649(.A1(new_n847), .A2(new_n849), .A3(new_n358), .ZN(new_n850));
  AOI21_X1  g0650(.A(new_n845), .B1(new_n846), .B2(new_n850), .ZN(new_n851));
  INV_X1    g0651(.A(new_n651), .ZN(new_n852));
  NOR2_X1   g0652(.A1(new_n851), .A2(new_n852), .ZN(new_n853));
  OAI21_X1  g0653(.A(new_n853), .B1(new_n395), .B2(new_n403), .ZN(new_n854));
  INV_X1    g0654(.A(new_n391), .ZN(new_n855));
  OAI21_X1  g0655(.A(new_n398), .B1(new_n851), .B2(new_n855), .ZN(new_n856));
  OAI21_X1  g0656(.A(KEYINPUT37), .B1(new_n856), .B2(new_n853), .ZN(new_n857));
  NAND2_X1  g0657(.A1(new_n378), .A2(new_n391), .ZN(new_n858));
  NAND2_X1  g0658(.A1(new_n378), .A2(new_n651), .ZN(new_n859));
  INV_X1    g0659(.A(KEYINPUT37), .ZN(new_n860));
  NAND4_X1  g0660(.A1(new_n858), .A2(new_n859), .A3(new_n860), .A4(new_n398), .ZN(new_n861));
  NAND2_X1  g0661(.A1(new_n857), .A2(new_n861), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n854), .A2(new_n862), .ZN(new_n863));
  INV_X1    g0663(.A(KEYINPUT38), .ZN(new_n864));
  NAND2_X1  g0664(.A1(new_n863), .A2(new_n864), .ZN(new_n865));
  NAND3_X1  g0665(.A1(new_n854), .A2(new_n862), .A3(KEYINPUT38), .ZN(new_n866));
  NAND2_X1  g0666(.A1(new_n865), .A2(new_n866), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n345), .A2(G169), .ZN(new_n868));
  NAND2_X1  g0668(.A1(new_n868), .A2(KEYINPUT14), .ZN(new_n869));
  NAND4_X1  g0669(.A1(new_n355), .A2(new_n869), .A3(new_n348), .A4(new_n347), .ZN(new_n870));
  INV_X1    g0670(.A(KEYINPUT94), .ZN(new_n871));
  NOR2_X1   g0671(.A1(new_n666), .A2(new_n353), .ZN(new_n872));
  NAND3_X1  g0672(.A1(new_n870), .A2(new_n871), .A3(new_n872), .ZN(new_n873));
  INV_X1    g0673(.A(new_n873), .ZN(new_n874));
  INV_X1    g0674(.A(new_n872), .ZN(new_n875));
  NAND3_X1  g0675(.A1(new_n351), .A2(new_n355), .A3(new_n875), .ZN(new_n876));
  AOI21_X1  g0676(.A(new_n871), .B1(new_n870), .B2(new_n872), .ZN(new_n877));
  AOI21_X1  g0677(.A(new_n874), .B1(new_n876), .B2(new_n877), .ZN(new_n878));
  AOI21_X1  g0678(.A(new_n790), .B1(new_n636), .B2(new_n643), .ZN(new_n879));
  OAI211_X1 g0679(.A(new_n867), .B(new_n878), .C1(new_n879), .C2(new_n803), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n395), .A2(new_n852), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n880), .A2(new_n881), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n882), .A2(KEYINPUT96), .ZN(new_n883));
  INV_X1    g0683(.A(KEYINPUT96), .ZN(new_n884));
  NAND3_X1  g0684(.A1(new_n880), .A2(new_n884), .A3(new_n881), .ZN(new_n885));
  INV_X1    g0685(.A(KEYINPUT39), .ZN(new_n886));
  INV_X1    g0686(.A(new_n859), .ZN(new_n887));
  INV_X1    g0687(.A(KEYINPUT98), .ZN(new_n888));
  NAND3_X1  g0688(.A1(new_n400), .A2(new_n888), .A3(new_n402), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n620), .A2(new_n889), .ZN(new_n890));
  AOI21_X1  g0690(.A(new_n888), .B1(new_n400), .B2(new_n402), .ZN(new_n891));
  OAI21_X1  g0691(.A(new_n887), .B1(new_n890), .B2(new_n891), .ZN(new_n892));
  NAND3_X1  g0692(.A1(new_n858), .A2(new_n859), .A3(new_n398), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n893), .A2(KEYINPUT37), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n894), .A2(new_n861), .ZN(new_n895));
  AOI21_X1  g0695(.A(KEYINPUT38), .B1(new_n892), .B2(new_n895), .ZN(new_n896));
  AND3_X1   g0696(.A1(new_n854), .A2(new_n862), .A3(KEYINPUT38), .ZN(new_n897));
  OAI21_X1  g0697(.A(new_n886), .B1(new_n896), .B2(new_n897), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n621), .A2(new_n666), .ZN(new_n899));
  XNOR2_X1  g0699(.A(new_n899), .B(KEYINPUT97), .ZN(new_n900));
  NAND3_X1  g0700(.A1(new_n865), .A2(KEYINPUT39), .A3(new_n866), .ZN(new_n901));
  AND3_X1   g0701(.A1(new_n898), .A2(new_n900), .A3(new_n901), .ZN(new_n902));
  INV_X1    g0702(.A(new_n902), .ZN(new_n903));
  NAND3_X1  g0703(.A1(new_n883), .A2(new_n885), .A3(new_n903), .ZN(new_n904));
  XOR2_X1   g0704(.A(new_n844), .B(new_n904), .Z(new_n905));
  INV_X1    g0705(.A(KEYINPUT40), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n877), .A2(new_n876), .ZN(new_n907));
  NAND3_X1  g0707(.A1(new_n907), .A2(new_n805), .A3(new_n873), .ZN(new_n908));
  OR3_X1    g0708(.A1(new_n617), .A2(new_n537), .A3(new_n653), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n710), .A2(new_n712), .ZN(new_n910));
  AND2_X1   g0710(.A1(new_n910), .A2(new_n714), .ZN(new_n911));
  AOI21_X1  g0711(.A(new_n908), .B1(new_n909), .B2(new_n911), .ZN(new_n912));
  INV_X1    g0712(.A(new_n891), .ZN(new_n913));
  NAND3_X1  g0713(.A1(new_n913), .A2(new_n620), .A3(new_n889), .ZN(new_n914));
  AOI22_X1  g0714(.A1(new_n914), .A2(new_n887), .B1(new_n861), .B2(new_n894), .ZN(new_n915));
  OAI21_X1  g0715(.A(new_n866), .B1(new_n915), .B2(KEYINPUT38), .ZN(new_n916));
  AOI21_X1  g0716(.A(new_n906), .B1(new_n912), .B2(new_n916), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n910), .A2(new_n714), .ZN(new_n918));
  OAI211_X1 g0718(.A(new_n878), .B(new_n805), .C1(new_n918), .C2(new_n716), .ZN(new_n919));
  AOI21_X1  g0719(.A(KEYINPUT38), .B1(new_n854), .B2(new_n862), .ZN(new_n920));
  OAI21_X1  g0720(.A(new_n906), .B1(new_n897), .B2(new_n920), .ZN(new_n921));
  NOR2_X1   g0721(.A1(new_n919), .A2(new_n921), .ZN(new_n922));
  NOR2_X1   g0722(.A1(new_n917), .A2(new_n922), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n911), .A2(new_n909), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n433), .A2(new_n924), .ZN(new_n925));
  OR2_X1    g0725(.A1(new_n923), .A2(new_n925), .ZN(new_n926));
  NAND2_X1  g0726(.A1(new_n923), .A2(new_n925), .ZN(new_n927));
  NAND3_X1  g0727(.A1(new_n926), .A2(G330), .A3(new_n927), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n905), .A2(new_n928), .ZN(new_n929));
  OAI21_X1  g0729(.A(new_n929), .B1(new_n261), .B2(new_n724), .ZN(new_n930));
  NOR2_X1   g0730(.A1(new_n905), .A2(new_n928), .ZN(new_n931));
  OAI21_X1  g0731(.A(new_n841), .B1(new_n930), .B2(new_n931), .ZN(G367));
  NAND2_X1  g0732(.A1(new_n563), .A2(new_n653), .ZN(new_n933));
  NAND3_X1  g0733(.A1(new_n576), .A2(new_n933), .A3(new_n614), .ZN(new_n934));
  NAND3_X1  g0734(.A1(new_n563), .A2(new_n575), .A3(new_n653), .ZN(new_n935));
  AND2_X1   g0735(.A1(new_n935), .A2(KEYINPUT100), .ZN(new_n936));
  NOR2_X1   g0736(.A1(new_n935), .A2(KEYINPUT100), .ZN(new_n937));
  OAI21_X1  g0737(.A(new_n934), .B1(new_n936), .B2(new_n937), .ZN(new_n938));
  INV_X1    g0738(.A(KEYINPUT101), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n938), .A2(new_n939), .ZN(new_n940));
  OAI211_X1 g0740(.A(new_n934), .B(KEYINPUT101), .C1(new_n936), .C2(new_n937), .ZN(new_n941));
  NAND2_X1  g0741(.A1(new_n940), .A2(new_n941), .ZN(new_n942));
  INV_X1    g0742(.A(new_n677), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n658), .A2(new_n943), .ZN(new_n944));
  INV_X1    g0744(.A(new_n944), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n942), .A2(new_n945), .ZN(new_n946));
  INV_X1    g0746(.A(KEYINPUT42), .ZN(new_n947));
  XNOR2_X1  g0747(.A(new_n946), .B(new_n947), .ZN(new_n948));
  INV_X1    g0748(.A(new_n942), .ZN(new_n949));
  OAI21_X1  g0749(.A(new_n576), .B1(new_n949), .B2(new_n656), .ZN(new_n950));
  NAND2_X1  g0750(.A1(new_n950), .A2(new_n666), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n948), .A2(new_n951), .ZN(new_n952));
  OR2_X1    g0752(.A1(new_n666), .A2(new_n598), .ZN(new_n953));
  XNOR2_X1  g0753(.A(new_n953), .B(new_n607), .ZN(new_n954));
  INV_X1    g0754(.A(KEYINPUT43), .ZN(new_n955));
  NAND2_X1  g0755(.A1(new_n954), .A2(new_n955), .ZN(new_n956));
  INV_X1    g0756(.A(new_n954), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n957), .A2(KEYINPUT43), .ZN(new_n958));
  NAND3_X1  g0758(.A1(new_n952), .A2(new_n956), .A3(new_n958), .ZN(new_n959));
  NAND4_X1  g0759(.A1(new_n948), .A2(new_n955), .A3(new_n951), .A4(new_n954), .ZN(new_n960));
  NAND2_X1  g0760(.A1(new_n959), .A2(new_n960), .ZN(new_n961));
  OAI21_X1  g0761(.A(new_n961), .B1(new_n672), .B2(new_n949), .ZN(new_n962));
  INV_X1    g0762(.A(new_n672), .ZN(new_n963));
  NAND4_X1  g0763(.A1(new_n959), .A2(new_n963), .A3(new_n942), .A4(new_n960), .ZN(new_n964));
  XOR2_X1   g0764(.A(new_n682), .B(KEYINPUT41), .Z(new_n965));
  NAND3_X1  g0765(.A1(new_n940), .A2(new_n678), .A3(new_n941), .ZN(new_n966));
  XOR2_X1   g0766(.A(KEYINPUT102), .B(KEYINPUT44), .Z(new_n967));
  XNOR2_X1  g0767(.A(new_n966), .B(new_n967), .ZN(new_n968));
  INV_X1    g0768(.A(new_n968), .ZN(new_n969));
  NAND3_X1  g0769(.A1(new_n942), .A2(new_n679), .A3(KEYINPUT45), .ZN(new_n970));
  INV_X1    g0770(.A(new_n970), .ZN(new_n971));
  AOI21_X1  g0771(.A(KEYINPUT45), .B1(new_n942), .B2(new_n679), .ZN(new_n972));
  NOR2_X1   g0772(.A1(new_n971), .A2(new_n972), .ZN(new_n973));
  OAI21_X1  g0773(.A(new_n963), .B1(new_n969), .B2(new_n973), .ZN(new_n974));
  OAI211_X1 g0774(.A(new_n968), .B(new_n672), .C1(new_n971), .C2(new_n972), .ZN(new_n975));
  OAI21_X1  g0775(.A(new_n944), .B1(new_n662), .B2(new_n943), .ZN(new_n976));
  XNOR2_X1  g0776(.A(new_n976), .B(new_n671), .ZN(new_n977));
  NAND4_X1  g0777(.A1(new_n974), .A2(new_n975), .A3(new_n719), .A4(new_n977), .ZN(new_n978));
  AOI21_X1  g0778(.A(new_n965), .B1(new_n978), .B2(new_n719), .ZN(new_n979));
  OAI211_X1 g0779(.A(new_n962), .B(new_n964), .C1(new_n979), .C2(new_n727), .ZN(new_n980));
  NOR3_X1   g0780(.A1(new_n238), .A2(new_n681), .A3(new_n283), .ZN(new_n981));
  OAI21_X1  g0781(.A(new_n777), .B1(new_n213), .B2(new_n409), .ZN(new_n982));
  OAI21_X1  g0782(.A(new_n728), .B1(new_n981), .B2(new_n982), .ZN(new_n983));
  INV_X1    g0783(.A(G150), .ZN(new_n984));
  OAI22_X1  g0784(.A1(new_n759), .A2(new_n984), .B1(new_n746), .B2(new_n287), .ZN(new_n985));
  OAI22_X1  g0785(.A1(new_n761), .A2(new_n814), .B1(new_n742), .B2(new_n364), .ZN(new_n986));
  NOR2_X1   g0786(.A1(new_n985), .A2(new_n986), .ZN(new_n987));
  NAND2_X1  g0787(.A1(new_n769), .A2(G68), .ZN(new_n988));
  NAND2_X1  g0788(.A1(new_n754), .A2(G137), .ZN(new_n989));
  OAI21_X1  g0789(.A(new_n283), .B1(new_n736), .B2(new_n767), .ZN(new_n990));
  AOI21_X1  g0790(.A(new_n990), .B1(G50), .B2(new_n812), .ZN(new_n991));
  NAND4_X1  g0791(.A1(new_n987), .A2(new_n988), .A3(new_n989), .A4(new_n991), .ZN(new_n992));
  OAI221_X1 g0792(.A(new_n330), .B1(new_n734), .B2(new_n824), .C1(new_n467), .C2(new_n736), .ZN(new_n993));
  AOI21_X1  g0793(.A(new_n993), .B1(G317), .B2(new_n754), .ZN(new_n994));
  INV_X1    g0794(.A(KEYINPUT46), .ZN(new_n995));
  OAI21_X1  g0795(.A(new_n995), .B1(new_n742), .B2(new_n448), .ZN(new_n996));
  NAND3_X1  g0796(.A1(new_n743), .A2(KEYINPUT46), .A3(G116), .ZN(new_n997));
  NAND3_X1  g0797(.A1(new_n994), .A2(new_n996), .A3(new_n997), .ZN(new_n998));
  AOI22_X1  g0798(.A1(new_n740), .A2(G303), .B1(new_n747), .B2(G97), .ZN(new_n999));
  OAI221_X1 g0799(.A(new_n999), .B1(new_n735), .B2(new_n761), .C1(new_n205), .C2(new_n757), .ZN(new_n1000));
  OAI21_X1  g0800(.A(new_n992), .B1(new_n998), .B2(new_n1000), .ZN(new_n1001));
  XOR2_X1   g0801(.A(KEYINPUT103), .B(KEYINPUT47), .Z(new_n1002));
  XNOR2_X1  g0802(.A(new_n1001), .B(new_n1002), .ZN(new_n1003));
  AOI21_X1  g0803(.A(new_n983), .B1(new_n1003), .B2(new_n730), .ZN(new_n1004));
  INV_X1    g0804(.A(new_n776), .ZN(new_n1005));
  OAI21_X1  g0805(.A(new_n1004), .B1(new_n957), .B2(new_n1005), .ZN(new_n1006));
  NAND2_X1  g0806(.A1(new_n980), .A2(new_n1006), .ZN(G387));
  NAND2_X1  g0807(.A1(new_n977), .A2(new_n727), .ZN(new_n1008));
  AOI22_X1  g0808(.A1(new_n769), .A2(G283), .B1(G294), .B2(new_n743), .ZN(new_n1009));
  AOI22_X1  g0809(.A1(new_n811), .A2(G311), .B1(new_n812), .B2(G303), .ZN(new_n1010));
  NAND2_X1  g0810(.A1(new_n740), .A2(G317), .ZN(new_n1011));
  NAND2_X1  g0811(.A1(new_n745), .A2(G322), .ZN(new_n1012));
  NAND3_X1  g0812(.A1(new_n1010), .A2(new_n1011), .A3(new_n1012), .ZN(new_n1013));
  INV_X1    g0813(.A(KEYINPUT48), .ZN(new_n1014));
  OAI21_X1  g0814(.A(new_n1009), .B1(new_n1013), .B2(new_n1014), .ZN(new_n1015));
  XOR2_X1   g0815(.A(new_n1015), .B(KEYINPUT105), .Z(new_n1016));
  NAND2_X1  g0816(.A1(new_n1013), .A2(new_n1014), .ZN(new_n1017));
  NAND2_X1  g0817(.A1(new_n1016), .A2(new_n1017), .ZN(new_n1018));
  XOR2_X1   g0818(.A(new_n1018), .B(KEYINPUT106), .Z(new_n1019));
  OR2_X1    g0819(.A1(new_n1019), .A2(KEYINPUT49), .ZN(new_n1020));
  NAND2_X1  g0820(.A1(new_n1019), .A2(KEYINPUT49), .ZN(new_n1021));
  OAI21_X1  g0821(.A(new_n330), .B1(new_n746), .B2(new_n448), .ZN(new_n1022));
  AOI21_X1  g0822(.A(new_n1022), .B1(new_n754), .B2(G326), .ZN(new_n1023));
  NAND3_X1  g0823(.A1(new_n1020), .A2(new_n1021), .A3(new_n1023), .ZN(new_n1024));
  OAI221_X1 g0824(.A(new_n283), .B1(new_n742), .B2(new_n287), .C1(new_n204), .C2(new_n746), .ZN(new_n1025));
  AOI21_X1  g0825(.A(new_n1025), .B1(G150), .B2(new_n754), .ZN(new_n1026));
  XOR2_X1   g0826(.A(new_n1026), .B(KEYINPUT104), .Z(new_n1027));
  NAND2_X1  g0827(.A1(new_n769), .A2(new_n410), .ZN(new_n1028));
  AOI22_X1  g0828(.A1(new_n811), .A2(new_n255), .B1(new_n812), .B2(G68), .ZN(new_n1029));
  OAI21_X1  g0829(.A(new_n1029), .B1(new_n767), .B2(new_n761), .ZN(new_n1030));
  AOI21_X1  g0830(.A(new_n1030), .B1(G50), .B2(new_n740), .ZN(new_n1031));
  NAND3_X1  g0831(.A1(new_n1027), .A2(new_n1028), .A3(new_n1031), .ZN(new_n1032));
  AOI21_X1  g0832(.A(new_n731), .B1(new_n1024), .B2(new_n1032), .ZN(new_n1033));
  OR2_X1    g0833(.A1(new_n235), .A2(new_n507), .ZN(new_n1034));
  AOI22_X1  g0834(.A1(new_n1034), .A2(new_n782), .B1(new_n684), .B2(new_n779), .ZN(new_n1035));
  INV_X1    g0835(.A(KEYINPUT50), .ZN(new_n1036));
  AOI21_X1  g0836(.A(new_n1036), .B1(new_n255), .B2(new_n250), .ZN(new_n1037));
  NOR3_X1   g0837(.A1(new_n254), .A2(KEYINPUT50), .A3(G50), .ZN(new_n1038));
  OAI21_X1  g0838(.A(new_n507), .B1(new_n217), .B2(new_n287), .ZN(new_n1039));
  NOR4_X1   g0839(.A1(new_n1037), .A2(new_n1038), .A3(new_n684), .A4(new_n1039), .ZN(new_n1040));
  OAI22_X1  g0840(.A1(new_n1035), .A2(new_n1040), .B1(G107), .B2(new_n213), .ZN(new_n1041));
  AOI21_X1  g0841(.A(new_n729), .B1(new_n1041), .B2(new_n778), .ZN(new_n1042));
  OAI21_X1  g0842(.A(new_n1042), .B1(new_n662), .B2(new_n1005), .ZN(new_n1043));
  NAND2_X1  g0843(.A1(new_n977), .A2(new_n719), .ZN(new_n1044));
  NAND2_X1  g0844(.A1(new_n1044), .A2(new_n682), .ZN(new_n1045));
  NOR2_X1   g0845(.A1(new_n977), .A2(new_n719), .ZN(new_n1046));
  OAI221_X1 g0846(.A(new_n1008), .B1(new_n1033), .B2(new_n1043), .C1(new_n1045), .C2(new_n1046), .ZN(G393));
  INV_X1    g0847(.A(KEYINPUT107), .ZN(new_n1048));
  NAND2_X1  g0848(.A1(new_n974), .A2(new_n1048), .ZN(new_n1049));
  INV_X1    g0849(.A(new_n1049), .ZN(new_n1050));
  AOI21_X1  g0850(.A(new_n1048), .B1(new_n974), .B2(new_n975), .ZN(new_n1051));
  OAI21_X1  g0851(.A(new_n1044), .B1(new_n1050), .B2(new_n1051), .ZN(new_n1052));
  AND2_X1   g0852(.A1(new_n978), .A2(new_n682), .ZN(new_n1053));
  NAND2_X1  g0853(.A1(new_n949), .A2(new_n776), .ZN(new_n1054));
  OAI21_X1  g0854(.A(new_n777), .B1(new_n204), .B2(new_n213), .ZN(new_n1055));
  AOI21_X1  g0855(.A(new_n1055), .B1(new_n242), .B2(new_n782), .ZN(new_n1056));
  XOR2_X1   g0856(.A(new_n1056), .B(KEYINPUT109), .Z(new_n1057));
  AOI22_X1  g0857(.A1(new_n740), .A2(G159), .B1(new_n745), .B2(G150), .ZN(new_n1058));
  XOR2_X1   g0858(.A(new_n1058), .B(KEYINPUT51), .Z(new_n1059));
  NAND2_X1  g0859(.A1(new_n769), .A2(G77), .ZN(new_n1060));
  OAI22_X1  g0860(.A1(new_n217), .A2(new_n742), .B1(new_n746), .B2(new_n683), .ZN(new_n1061));
  OAI221_X1 g0861(.A(new_n283), .B1(new_n734), .B2(new_n254), .C1(new_n250), .C2(new_n736), .ZN(new_n1062));
  AOI211_X1 g0862(.A(new_n1061), .B(new_n1062), .C1(G143), .C2(new_n754), .ZN(new_n1063));
  NAND3_X1  g0863(.A1(new_n1059), .A2(new_n1060), .A3(new_n1063), .ZN(new_n1064));
  XOR2_X1   g0864(.A(new_n1064), .B(KEYINPUT110), .Z(new_n1065));
  AOI22_X1  g0865(.A1(new_n811), .A2(G303), .B1(new_n812), .B2(G294), .ZN(new_n1066));
  OAI21_X1  g0866(.A(new_n1066), .B1(new_n448), .B2(new_n757), .ZN(new_n1067));
  XOR2_X1   g0867(.A(new_n1067), .B(KEYINPUT111), .Z(new_n1068));
  AOI22_X1  g0868(.A1(new_n740), .A2(G311), .B1(new_n745), .B2(G317), .ZN(new_n1069));
  XOR2_X1   g0869(.A(new_n1069), .B(KEYINPUT52), .Z(new_n1070));
  OAI221_X1 g0870(.A(new_n330), .B1(new_n742), .B2(new_n824), .C1(new_n205), .C2(new_n746), .ZN(new_n1071));
  AOI21_X1  g0871(.A(new_n1071), .B1(G322), .B2(new_n754), .ZN(new_n1072));
  NAND3_X1  g0872(.A1(new_n1068), .A2(new_n1070), .A3(new_n1072), .ZN(new_n1073));
  NAND2_X1  g0873(.A1(new_n1073), .A2(KEYINPUT112), .ZN(new_n1074));
  OR2_X1    g0874(.A1(new_n1073), .A2(KEYINPUT112), .ZN(new_n1075));
  NAND3_X1  g0875(.A1(new_n1065), .A2(new_n1074), .A3(new_n1075), .ZN(new_n1076));
  AOI211_X1 g0876(.A(new_n729), .B(new_n1057), .C1(new_n1076), .C2(new_n730), .ZN(new_n1077));
  AOI22_X1  g0877(.A1(new_n1052), .A2(new_n1053), .B1(new_n1054), .B2(new_n1077), .ZN(new_n1078));
  INV_X1    g0878(.A(new_n1051), .ZN(new_n1079));
  NAND3_X1  g0879(.A1(new_n1079), .A2(KEYINPUT108), .A3(new_n1049), .ZN(new_n1080));
  INV_X1    g0880(.A(KEYINPUT108), .ZN(new_n1081));
  OAI21_X1  g0881(.A(new_n1081), .B1(new_n1050), .B2(new_n1051), .ZN(new_n1082));
  NAND3_X1  g0882(.A1(new_n1080), .A2(new_n1082), .A3(new_n727), .ZN(new_n1083));
  NAND2_X1  g0883(.A1(new_n1078), .A2(new_n1083), .ZN(G390));
  INV_X1    g0884(.A(KEYINPUT113), .ZN(new_n1085));
  NAND2_X1  g0885(.A1(new_n907), .A2(new_n873), .ZN(new_n1086));
  INV_X1    g0886(.A(new_n803), .ZN(new_n1087));
  AOI21_X1  g0887(.A(new_n1086), .B1(new_n798), .B2(new_n1087), .ZN(new_n1088));
  OAI21_X1  g0888(.A(new_n1085), .B1(new_n1088), .B2(new_n900), .ZN(new_n1089));
  NAND2_X1  g0889(.A1(new_n898), .A2(new_n901), .ZN(new_n1090));
  INV_X1    g0890(.A(new_n900), .ZN(new_n1091));
  AOI21_X1  g0891(.A(new_n803), .B1(new_n644), .B2(new_n791), .ZN(new_n1092));
  OAI211_X1 g0892(.A(KEYINPUT113), .B(new_n1091), .C1(new_n1092), .C2(new_n1086), .ZN(new_n1093));
  NAND3_X1  g0893(.A1(new_n1089), .A2(new_n1090), .A3(new_n1093), .ZN(new_n1094));
  NAND2_X1  g0894(.A1(new_n916), .A2(new_n1091), .ZN(new_n1095));
  NAND2_X1  g0895(.A1(new_n425), .A2(new_n804), .ZN(new_n1096));
  OAI211_X1 g0896(.A(new_n666), .B(new_n1096), .C1(new_n689), .C2(new_n691), .ZN(new_n1097));
  NAND2_X1  g0897(.A1(new_n1097), .A2(new_n1087), .ZN(new_n1098));
  AOI21_X1  g0898(.A(new_n1095), .B1(new_n878), .B2(new_n1098), .ZN(new_n1099));
  INV_X1    g0899(.A(new_n1099), .ZN(new_n1100));
  OAI211_X1 g0900(.A(G330), .B(new_n805), .C1(new_n715), .C2(new_n716), .ZN(new_n1101));
  OR2_X1    g0901(.A1(new_n1101), .A2(new_n1086), .ZN(new_n1102));
  NAND3_X1  g0902(.A1(new_n1094), .A2(new_n1100), .A3(new_n1102), .ZN(new_n1103));
  NAND3_X1  g0903(.A1(new_n433), .A2(G330), .A3(new_n924), .ZN(new_n1104));
  NAND3_X1  g0904(.A1(new_n842), .A2(new_n625), .A3(new_n1104), .ZN(new_n1105));
  NAND3_X1  g0905(.A1(new_n924), .A2(G330), .A3(new_n805), .ZN(new_n1106));
  NAND2_X1  g0906(.A1(new_n1106), .A2(new_n1086), .ZN(new_n1107));
  NAND4_X1  g0907(.A1(new_n1102), .A2(new_n1107), .A3(new_n1087), .A4(new_n1097), .ZN(new_n1108));
  AND2_X1   g0908(.A1(new_n1101), .A2(new_n1086), .ZN(new_n1109));
  INV_X1    g0909(.A(new_n908), .ZN(new_n1110));
  NAND3_X1  g0910(.A1(new_n924), .A2(new_n1110), .A3(G330), .ZN(new_n1111));
  INV_X1    g0911(.A(new_n1111), .ZN(new_n1112));
  OAI22_X1  g0912(.A1(new_n1109), .A2(new_n1112), .B1(new_n879), .B2(new_n803), .ZN(new_n1113));
  AOI21_X1  g0913(.A(new_n1105), .B1(new_n1108), .B2(new_n1113), .ZN(new_n1114));
  INV_X1    g0914(.A(new_n1090), .ZN(new_n1115));
  OAI21_X1  g0915(.A(new_n1091), .B1(new_n1092), .B2(new_n1086), .ZN(new_n1116));
  AOI21_X1  g0916(.A(new_n1115), .B1(new_n1116), .B2(new_n1085), .ZN(new_n1117));
  AOI21_X1  g0917(.A(new_n1099), .B1(new_n1117), .B2(new_n1093), .ZN(new_n1118));
  OAI211_X1 g0918(.A(new_n1103), .B(new_n1114), .C1(new_n1118), .C2(new_n1111), .ZN(new_n1119));
  NAND2_X1  g0919(.A1(new_n1119), .A2(KEYINPUT114), .ZN(new_n1120));
  NAND2_X1  g0920(.A1(new_n1094), .A2(new_n1100), .ZN(new_n1121));
  NAND2_X1  g0921(.A1(new_n1121), .A2(new_n1112), .ZN(new_n1122));
  INV_X1    g0922(.A(KEYINPUT114), .ZN(new_n1123));
  NAND4_X1  g0923(.A1(new_n1122), .A2(new_n1123), .A3(new_n1103), .A4(new_n1114), .ZN(new_n1124));
  NAND2_X1  g0924(.A1(new_n1120), .A2(new_n1124), .ZN(new_n1125));
  NAND2_X1  g0925(.A1(new_n1122), .A2(new_n1103), .ZN(new_n1126));
  INV_X1    g0926(.A(new_n1114), .ZN(new_n1127));
  AOI21_X1  g0927(.A(new_n723), .B1(new_n1126), .B2(new_n1127), .ZN(new_n1128));
  NAND2_X1  g0928(.A1(new_n1125), .A2(new_n1128), .ZN(new_n1129));
  OAI22_X1  g0929(.A1(new_n448), .A2(new_n759), .B1(new_n761), .B2(new_n824), .ZN(new_n1130));
  OAI22_X1  g0930(.A1(new_n217), .A2(new_n746), .B1(new_n742), .B2(new_n683), .ZN(new_n1131));
  NOR2_X1   g0931(.A1(new_n1130), .A2(new_n1131), .ZN(new_n1132));
  NAND2_X1  g0932(.A1(new_n754), .A2(G294), .ZN(new_n1133));
  OAI21_X1  g0933(.A(new_n330), .B1(new_n736), .B2(new_n205), .ZN(new_n1134));
  AOI21_X1  g0934(.A(new_n1134), .B1(G97), .B2(new_n812), .ZN(new_n1135));
  NAND4_X1  g0935(.A1(new_n1132), .A2(new_n1060), .A3(new_n1133), .A4(new_n1135), .ZN(new_n1136));
  OAI21_X1  g0936(.A(new_n283), .B1(new_n736), .B2(new_n815), .ZN(new_n1137));
  AOI21_X1  g0937(.A(new_n1137), .B1(G128), .B2(new_n745), .ZN(new_n1138));
  AOI22_X1  g0938(.A1(new_n740), .A2(G132), .B1(new_n747), .B2(G50), .ZN(new_n1139));
  XNOR2_X1  g0939(.A(KEYINPUT54), .B(G143), .ZN(new_n1140));
  XNOR2_X1  g0940(.A(new_n1140), .B(KEYINPUT115), .ZN(new_n1141));
  NAND2_X1  g0941(.A1(new_n1141), .A2(new_n812), .ZN(new_n1142));
  NAND2_X1  g0942(.A1(new_n754), .A2(G125), .ZN(new_n1143));
  NAND4_X1  g0943(.A1(new_n1138), .A2(new_n1139), .A3(new_n1142), .A4(new_n1143), .ZN(new_n1144));
  NOR2_X1   g0944(.A1(new_n742), .A2(new_n984), .ZN(new_n1145));
  XNOR2_X1  g0945(.A(new_n1145), .B(KEYINPUT53), .ZN(new_n1146));
  OAI21_X1  g0946(.A(new_n1146), .B1(new_n767), .B2(new_n757), .ZN(new_n1147));
  OAI21_X1  g0947(.A(new_n1136), .B1(new_n1144), .B2(new_n1147), .ZN(new_n1148));
  NAND2_X1  g0948(.A1(new_n1148), .A2(new_n730), .ZN(new_n1149));
  INV_X1    g0949(.A(new_n809), .ZN(new_n1150));
  OAI211_X1 g0950(.A(new_n1149), .B(new_n728), .C1(new_n255), .C2(new_n1150), .ZN(new_n1151));
  AOI21_X1  g0951(.A(new_n1151), .B1(new_n1090), .B2(new_n774), .ZN(new_n1152));
  XNOR2_X1  g0952(.A(new_n1152), .B(KEYINPUT116), .ZN(new_n1153));
  NAND3_X1  g0953(.A1(new_n1122), .A2(new_n727), .A3(new_n1103), .ZN(new_n1154));
  NAND3_X1  g0954(.A1(new_n1129), .A2(new_n1153), .A3(new_n1154), .ZN(G378));
  NOR2_X1   g0955(.A1(new_n268), .A2(new_n852), .ZN(new_n1156));
  XNOR2_X1  g0956(.A(new_n1156), .B(KEYINPUT55), .ZN(new_n1157));
  XNOR2_X1  g0957(.A(new_n311), .B(new_n1157), .ZN(new_n1158));
  XOR2_X1   g0958(.A(KEYINPUT118), .B(KEYINPUT56), .Z(new_n1159));
  XOR2_X1   g0959(.A(new_n1158), .B(new_n1159), .Z(new_n1160));
  INV_X1    g0960(.A(new_n1160), .ZN(new_n1161));
  OAI21_X1  g0961(.A(G330), .B1(new_n917), .B2(new_n922), .ZN(new_n1162));
  AND4_X1   g0962(.A1(new_n885), .A2(new_n883), .A3(new_n903), .A4(new_n1162), .ZN(new_n1163));
  AOI21_X1  g0963(.A(new_n902), .B1(new_n882), .B2(KEYINPUT96), .ZN(new_n1164));
  AOI21_X1  g0964(.A(new_n1162), .B1(new_n1164), .B2(new_n885), .ZN(new_n1165));
  OAI21_X1  g0965(.A(new_n1161), .B1(new_n1163), .B2(new_n1165), .ZN(new_n1166));
  INV_X1    g0966(.A(new_n1162), .ZN(new_n1167));
  NAND2_X1  g0967(.A1(new_n904), .A2(new_n1167), .ZN(new_n1168));
  NAND3_X1  g0968(.A1(new_n1164), .A2(new_n885), .A3(new_n1162), .ZN(new_n1169));
  NAND3_X1  g0969(.A1(new_n1168), .A2(new_n1169), .A3(new_n1160), .ZN(new_n1170));
  AND3_X1   g0970(.A1(new_n1166), .A2(KEYINPUT120), .A3(new_n1170), .ZN(new_n1171));
  AOI21_X1  g0971(.A(KEYINPUT120), .B1(new_n1166), .B2(new_n1170), .ZN(new_n1172));
  NOR2_X1   g0972(.A1(new_n1171), .A2(new_n1172), .ZN(new_n1173));
  INV_X1    g0973(.A(new_n1105), .ZN(new_n1174));
  NAND2_X1  g0974(.A1(new_n1125), .A2(new_n1174), .ZN(new_n1175));
  AOI21_X1  g0975(.A(KEYINPUT57), .B1(new_n1173), .B2(new_n1175), .ZN(new_n1176));
  AOI21_X1  g0976(.A(new_n1105), .B1(new_n1120), .B2(new_n1124), .ZN(new_n1177));
  NAND2_X1  g0977(.A1(new_n1166), .A2(new_n1170), .ZN(new_n1178));
  NAND2_X1  g0978(.A1(new_n1178), .A2(KEYINPUT57), .ZN(new_n1179));
  OAI21_X1  g0979(.A(new_n682), .B1(new_n1177), .B2(new_n1179), .ZN(new_n1180));
  OR2_X1    g0980(.A1(new_n1176), .A2(new_n1180), .ZN(new_n1181));
  OAI21_X1  g0981(.A(new_n728), .B1(G50), .B2(new_n1150), .ZN(new_n1182));
  NAND2_X1  g0982(.A1(new_n330), .A2(new_n474), .ZN(new_n1183));
  OAI211_X1 g0983(.A(new_n1183), .B(new_n250), .C1(G33), .C2(G41), .ZN(new_n1184));
  NOR2_X1   g0984(.A1(new_n746), .A2(new_n364), .ZN(new_n1185));
  OAI22_X1  g0985(.A1(new_n761), .A2(new_n448), .B1(new_n742), .B2(new_n287), .ZN(new_n1186));
  AOI211_X1 g0986(.A(new_n1185), .B(new_n1186), .C1(G107), .C2(new_n740), .ZN(new_n1187));
  NAND2_X1  g0987(.A1(new_n754), .A2(G283), .ZN(new_n1188));
  NOR2_X1   g0988(.A1(new_n734), .A2(new_n409), .ZN(new_n1189));
  AOI211_X1 g0989(.A(new_n1183), .B(new_n1189), .C1(G97), .C2(new_n811), .ZN(new_n1190));
  NAND4_X1  g0990(.A1(new_n1187), .A2(new_n988), .A3(new_n1188), .A4(new_n1190), .ZN(new_n1191));
  INV_X1    g0991(.A(KEYINPUT58), .ZN(new_n1192));
  OAI21_X1  g0992(.A(new_n1184), .B1(new_n1191), .B2(new_n1192), .ZN(new_n1193));
  AOI21_X1  g0993(.A(new_n1193), .B1(new_n1192), .B2(new_n1191), .ZN(new_n1194));
  AOI22_X1  g0994(.A1(new_n811), .A2(G132), .B1(new_n812), .B2(G137), .ZN(new_n1195));
  INV_X1    g0995(.A(G128), .ZN(new_n1196));
  OAI21_X1  g0996(.A(new_n1195), .B1(new_n1196), .B2(new_n759), .ZN(new_n1197));
  AOI21_X1  g0997(.A(new_n1197), .B1(G125), .B2(new_n745), .ZN(new_n1198));
  NAND2_X1  g0998(.A1(new_n1141), .A2(new_n743), .ZN(new_n1199));
  OAI211_X1 g0999(.A(new_n1198), .B(new_n1199), .C1(new_n984), .C2(new_n757), .ZN(new_n1200));
  XNOR2_X1  g1000(.A(new_n1200), .B(KEYINPUT117), .ZN(new_n1201));
  INV_X1    g1001(.A(new_n1201), .ZN(new_n1202));
  NOR2_X1   g1002(.A1(new_n1202), .A2(KEYINPUT59), .ZN(new_n1203));
  OAI211_X1 g1003(.A(new_n256), .B(new_n474), .C1(new_n746), .C2(new_n767), .ZN(new_n1204));
  AOI21_X1  g1004(.A(new_n1204), .B1(new_n754), .B2(G124), .ZN(new_n1205));
  INV_X1    g1005(.A(KEYINPUT59), .ZN(new_n1206));
  OAI21_X1  g1006(.A(new_n1205), .B1(new_n1201), .B2(new_n1206), .ZN(new_n1207));
  OAI21_X1  g1007(.A(new_n1194), .B1(new_n1203), .B2(new_n1207), .ZN(new_n1208));
  AOI21_X1  g1008(.A(new_n1182), .B1(new_n1208), .B2(new_n730), .ZN(new_n1209));
  OAI21_X1  g1009(.A(new_n1209), .B1(new_n1161), .B2(new_n775), .ZN(new_n1210));
  XNOR2_X1  g1010(.A(new_n1210), .B(KEYINPUT119), .ZN(new_n1211));
  AOI21_X1  g1011(.A(new_n1211), .B1(new_n1173), .B2(new_n727), .ZN(new_n1212));
  NAND2_X1  g1012(.A1(new_n1181), .A2(new_n1212), .ZN(G375));
  NAND2_X1  g1013(.A1(new_n1086), .A2(new_n774), .ZN(new_n1214));
  XNOR2_X1  g1014(.A(new_n1214), .B(KEYINPUT121), .ZN(new_n1215));
  OAI21_X1  g1015(.A(new_n728), .B1(G68), .B2(new_n1150), .ZN(new_n1216));
  XOR2_X1   g1016(.A(new_n1216), .B(KEYINPUT122), .Z(new_n1217));
  AOI211_X1 g1017(.A(new_n330), .B(new_n1185), .C1(G150), .C2(new_n812), .ZN(new_n1218));
  NAND2_X1  g1018(.A1(new_n1141), .A2(new_n811), .ZN(new_n1219));
  AOI22_X1  g1019(.A1(new_n740), .A2(G137), .B1(new_n745), .B2(G132), .ZN(new_n1220));
  NAND3_X1  g1020(.A1(new_n1218), .A2(new_n1219), .A3(new_n1220), .ZN(new_n1221));
  AOI21_X1  g1021(.A(new_n1221), .B1(G50), .B2(new_n769), .ZN(new_n1222));
  AOI22_X1  g1022(.A1(new_n754), .A2(G128), .B1(G159), .B2(new_n743), .ZN(new_n1223));
  XOR2_X1   g1023(.A(new_n1223), .B(KEYINPUT123), .Z(new_n1224));
  NOR2_X1   g1024(.A1(new_n766), .A2(new_n502), .ZN(new_n1225));
  OAI22_X1  g1025(.A1(new_n824), .A2(new_n759), .B1(new_n761), .B2(new_n467), .ZN(new_n1226));
  OAI22_X1  g1026(.A1(new_n287), .A2(new_n746), .B1(new_n742), .B2(new_n204), .ZN(new_n1227));
  OAI221_X1 g1027(.A(new_n330), .B1(new_n734), .B2(new_n205), .C1(new_n448), .C2(new_n736), .ZN(new_n1228));
  NOR4_X1   g1028(.A1(new_n1225), .A2(new_n1226), .A3(new_n1227), .A4(new_n1228), .ZN(new_n1229));
  AOI22_X1  g1029(.A1(new_n1222), .A2(new_n1224), .B1(new_n1028), .B2(new_n1229), .ZN(new_n1230));
  OAI211_X1 g1030(.A(new_n1215), .B(new_n1217), .C1(new_n731), .C2(new_n1230), .ZN(new_n1231));
  AND2_X1   g1031(.A1(new_n1108), .A2(new_n1113), .ZN(new_n1232));
  OAI21_X1  g1032(.A(new_n1231), .B1(new_n1232), .B2(new_n725), .ZN(new_n1233));
  INV_X1    g1033(.A(KEYINPUT124), .ZN(new_n1234));
  XNOR2_X1  g1034(.A(new_n1233), .B(new_n1234), .ZN(new_n1235));
  AND2_X1   g1035(.A1(new_n1232), .A2(new_n1105), .ZN(new_n1236));
  OR2_X1    g1036(.A1(new_n1114), .A2(new_n965), .ZN(new_n1237));
  OAI21_X1  g1037(.A(new_n1235), .B1(new_n1236), .B2(new_n1237), .ZN(G381));
  OR2_X1    g1038(.A1(G393), .A2(G396), .ZN(new_n1239));
  OR4_X1    g1039(.A1(G384), .A2(G387), .A3(new_n1239), .A4(G381), .ZN(new_n1240));
  OR4_X1    g1040(.A1(G390), .A2(G375), .A3(new_n1240), .A4(G378), .ZN(G407));
  AND3_X1   g1041(.A1(new_n1129), .A2(new_n1153), .A3(new_n1154), .ZN(new_n1242));
  INV_X1    g1042(.A(G343), .ZN(new_n1243));
  NAND2_X1  g1043(.A1(new_n1243), .A2(G213), .ZN(new_n1244));
  XNOR2_X1  g1044(.A(new_n1244), .B(KEYINPUT125), .ZN(new_n1245));
  NAND2_X1  g1045(.A1(new_n1242), .A2(new_n1245), .ZN(new_n1246));
  OAI211_X1 g1046(.A(G407), .B(G213), .C1(G375), .C2(new_n1246), .ZN(G409));
  NAND3_X1  g1047(.A1(G390), .A2(new_n1006), .A3(new_n980), .ZN(new_n1248));
  XNOR2_X1  g1048(.A(G393), .B(new_n788), .ZN(new_n1249));
  INV_X1    g1049(.A(new_n1249), .ZN(new_n1250));
  AND2_X1   g1050(.A1(new_n1248), .A2(new_n1250), .ZN(new_n1251));
  INV_X1    g1051(.A(KEYINPUT126), .ZN(new_n1252));
  AOI22_X1  g1052(.A1(G390), .A2(new_n1252), .B1(new_n1006), .B2(new_n980), .ZN(new_n1253));
  NAND3_X1  g1053(.A1(new_n1078), .A2(new_n1083), .A3(KEYINPUT126), .ZN(new_n1254));
  NAND3_X1  g1054(.A1(new_n1253), .A2(KEYINPUT127), .A3(new_n1254), .ZN(new_n1255));
  INV_X1    g1055(.A(new_n1255), .ZN(new_n1256));
  AOI21_X1  g1056(.A(KEYINPUT127), .B1(new_n1253), .B2(new_n1254), .ZN(new_n1257));
  OAI21_X1  g1057(.A(new_n1251), .B1(new_n1256), .B2(new_n1257), .ZN(new_n1258));
  NAND3_X1  g1058(.A1(G387), .A2(new_n1083), .A3(new_n1078), .ZN(new_n1259));
  AOI21_X1  g1059(.A(new_n1250), .B1(new_n1248), .B2(new_n1259), .ZN(new_n1260));
  INV_X1    g1060(.A(new_n1260), .ZN(new_n1261));
  NAND2_X1  g1061(.A1(new_n1258), .A2(new_n1261), .ZN(new_n1262));
  INV_X1    g1062(.A(KEYINPUT63), .ZN(new_n1263));
  OAI211_X1 g1063(.A(G378), .B(new_n1212), .C1(new_n1176), .C2(new_n1180), .ZN(new_n1264));
  NOR4_X1   g1064(.A1(new_n1177), .A2(new_n1171), .A3(new_n1172), .A4(new_n965), .ZN(new_n1265));
  AOI21_X1  g1065(.A(new_n725), .B1(new_n1166), .B2(new_n1170), .ZN(new_n1266));
  OR2_X1    g1066(.A1(new_n1211), .A2(new_n1266), .ZN(new_n1267));
  OAI21_X1  g1067(.A(new_n1242), .B1(new_n1265), .B2(new_n1267), .ZN(new_n1268));
  NAND2_X1  g1068(.A1(new_n1264), .A2(new_n1268), .ZN(new_n1269));
  INV_X1    g1069(.A(new_n1245), .ZN(new_n1270));
  NAND2_X1  g1070(.A1(new_n1269), .A2(new_n1270), .ZN(new_n1271));
  NAND3_X1  g1071(.A1(new_n1232), .A2(KEYINPUT60), .A3(new_n1105), .ZN(new_n1272));
  AND2_X1   g1072(.A1(new_n1272), .A2(new_n682), .ZN(new_n1273));
  AND2_X1   g1073(.A1(new_n1127), .A2(KEYINPUT60), .ZN(new_n1274));
  OAI21_X1  g1074(.A(new_n1273), .B1(new_n1236), .B2(new_n1274), .ZN(new_n1275));
  NAND2_X1  g1075(.A1(new_n1275), .A2(new_n1235), .ZN(new_n1276));
  NAND2_X1  g1076(.A1(new_n1276), .A2(new_n829), .ZN(new_n1277));
  INV_X1    g1077(.A(new_n1277), .ZN(new_n1278));
  NOR2_X1   g1078(.A1(new_n1276), .A2(new_n829), .ZN(new_n1279));
  NOR2_X1   g1079(.A1(new_n1278), .A2(new_n1279), .ZN(new_n1280));
  INV_X1    g1080(.A(new_n1280), .ZN(new_n1281));
  OAI21_X1  g1081(.A(new_n1263), .B1(new_n1271), .B2(new_n1281), .ZN(new_n1282));
  NAND2_X1  g1082(.A1(new_n1245), .A2(G2897), .ZN(new_n1283));
  INV_X1    g1083(.A(new_n1283), .ZN(new_n1284));
  OAI21_X1  g1084(.A(new_n1284), .B1(new_n1278), .B2(new_n1279), .ZN(new_n1285));
  INV_X1    g1085(.A(new_n1279), .ZN(new_n1286));
  NAND3_X1  g1086(.A1(new_n1286), .A2(new_n1277), .A3(new_n1283), .ZN(new_n1287));
  AND2_X1   g1087(.A1(new_n1285), .A2(new_n1287), .ZN(new_n1288));
  AOI21_X1  g1088(.A(KEYINPUT61), .B1(new_n1271), .B2(new_n1288), .ZN(new_n1289));
  AOI21_X1  g1089(.A(new_n1245), .B1(new_n1264), .B2(new_n1268), .ZN(new_n1290));
  NAND3_X1  g1090(.A1(new_n1290), .A2(KEYINPUT63), .A3(new_n1280), .ZN(new_n1291));
  NAND4_X1  g1091(.A1(new_n1262), .A2(new_n1282), .A3(new_n1289), .A4(new_n1291), .ZN(new_n1292));
  INV_X1    g1092(.A(KEYINPUT62), .ZN(new_n1293));
  AND3_X1   g1093(.A1(new_n1290), .A2(new_n1293), .A3(new_n1280), .ZN(new_n1294));
  INV_X1    g1094(.A(KEYINPUT61), .ZN(new_n1295));
  NAND2_X1  g1095(.A1(new_n1285), .A2(new_n1287), .ZN(new_n1296));
  OAI21_X1  g1096(.A(new_n1295), .B1(new_n1290), .B2(new_n1296), .ZN(new_n1297));
  AOI21_X1  g1097(.A(new_n1293), .B1(new_n1290), .B2(new_n1280), .ZN(new_n1298));
  NOR3_X1   g1098(.A1(new_n1294), .A2(new_n1297), .A3(new_n1298), .ZN(new_n1299));
  OAI21_X1  g1099(.A(new_n1292), .B1(new_n1299), .B2(new_n1262), .ZN(G405));
  NAND2_X1  g1100(.A1(G390), .A2(new_n1252), .ZN(new_n1301));
  NAND3_X1  g1101(.A1(new_n1301), .A2(G387), .A3(new_n1254), .ZN(new_n1302));
  INV_X1    g1102(.A(KEYINPUT127), .ZN(new_n1303));
  NAND2_X1  g1103(.A1(new_n1302), .A2(new_n1303), .ZN(new_n1304));
  NAND2_X1  g1104(.A1(new_n1304), .A2(new_n1255), .ZN(new_n1305));
  AOI21_X1  g1105(.A(new_n1260), .B1(new_n1305), .B2(new_n1251), .ZN(new_n1306));
  NAND2_X1  g1106(.A1(G375), .A2(new_n1242), .ZN(new_n1307));
  NAND3_X1  g1107(.A1(new_n1307), .A2(new_n1281), .A3(new_n1264), .ZN(new_n1308));
  AOI21_X1  g1108(.A(G378), .B1(new_n1181), .B2(new_n1212), .ZN(new_n1309));
  INV_X1    g1109(.A(new_n1264), .ZN(new_n1310));
  OAI21_X1  g1110(.A(new_n1280), .B1(new_n1309), .B2(new_n1310), .ZN(new_n1311));
  AND3_X1   g1111(.A1(new_n1306), .A2(new_n1308), .A3(new_n1311), .ZN(new_n1312));
  AOI21_X1  g1112(.A(new_n1306), .B1(new_n1311), .B2(new_n1308), .ZN(new_n1313));
  NOR2_X1   g1113(.A1(new_n1312), .A2(new_n1313), .ZN(G402));
endmodule


