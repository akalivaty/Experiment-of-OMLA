//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 0 0 1 0 1 0 1 1 0 1 0 1 0 1 1 1 1 0 1 0 1 1 0 0 0 0 1 0 1 0 0 0 1 1 0 1 0 1 0 1 1 1 1 1 1 0 0 0 0 1 0 1 0 1 0 1 1 1 0 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:17:18 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n713, new_n714,
    new_n716, new_n717, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n733, new_n734, new_n735, new_n736, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n762,
    new_n763, new_n764, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n775, new_n776, new_n777, new_n778,
    new_n779, new_n781, new_n783, new_n784, new_n785, new_n786, new_n787,
    new_n788, new_n789, new_n790, new_n791, new_n792, new_n793, new_n794,
    new_n795, new_n796, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n812, new_n813, new_n814, new_n815, new_n816, new_n817,
    new_n818, new_n819, new_n820, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n866, new_n867, new_n869, new_n870,
    new_n871, new_n873, new_n874, new_n875, new_n876, new_n877, new_n878,
    new_n879, new_n880, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n930,
    new_n931, new_n932, new_n933, new_n935, new_n936, new_n937, new_n938,
    new_n939, new_n940, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n953, new_n954,
    new_n955, new_n957, new_n958, new_n959, new_n961, new_n962, new_n963,
    new_n964, new_n965, new_n966, new_n967, new_n968, new_n970, new_n971,
    new_n972, new_n973, new_n974, new_n975, new_n976, new_n977, new_n978,
    new_n979, new_n980, new_n981, new_n982, new_n983, new_n984, new_n985,
    new_n986, new_n987, new_n988, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010;
  XOR2_X1   g000(.A(G183gat), .B(G211gat), .Z(new_n202));
  INV_X1    g001(.A(KEYINPUT9), .ZN(new_n203));
  INV_X1    g002(.A(G71gat), .ZN(new_n204));
  INV_X1    g003(.A(G78gat), .ZN(new_n205));
  OAI21_X1  g004(.A(new_n203), .B1(new_n204), .B2(new_n205), .ZN(new_n206));
  INV_X1    g005(.A(KEYINPUT92), .ZN(new_n207));
  NAND2_X1  g006(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  XOR2_X1   g007(.A(G57gat), .B(G64gat), .Z(new_n209));
  OAI211_X1 g008(.A(KEYINPUT92), .B(new_n203), .C1(new_n204), .C2(new_n205), .ZN(new_n210));
  NAND3_X1  g009(.A1(new_n208), .A2(new_n209), .A3(new_n210), .ZN(new_n211));
  XOR2_X1   g010(.A(G71gat), .B(G78gat), .Z(new_n212));
  NOR2_X1   g011(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  INV_X1    g012(.A(KEYINPUT94), .ZN(new_n214));
  XNOR2_X1  g013(.A(new_n213), .B(new_n214), .ZN(new_n215));
  NAND2_X1  g014(.A1(new_n211), .A2(new_n212), .ZN(new_n216));
  INV_X1    g015(.A(KEYINPUT93), .ZN(new_n217));
  XNOR2_X1  g016(.A(new_n216), .B(new_n217), .ZN(new_n218));
  AOI21_X1  g017(.A(KEYINPUT21), .B1(new_n215), .B2(new_n218), .ZN(new_n219));
  AND2_X1   g018(.A1(G231gat), .A2(G233gat), .ZN(new_n220));
  XNOR2_X1  g019(.A(new_n219), .B(new_n220), .ZN(new_n221));
  XOR2_X1   g020(.A(G127gat), .B(G155gat), .Z(new_n222));
  XNOR2_X1  g021(.A(new_n222), .B(KEYINPUT20), .ZN(new_n223));
  INV_X1    g022(.A(new_n223), .ZN(new_n224));
  NAND2_X1  g023(.A1(new_n221), .A2(new_n224), .ZN(new_n225));
  INV_X1    g024(.A(new_n225), .ZN(new_n226));
  NOR2_X1   g025(.A1(new_n221), .A2(new_n224), .ZN(new_n227));
  OAI21_X1  g026(.A(new_n202), .B1(new_n226), .B2(new_n227), .ZN(new_n228));
  INV_X1    g027(.A(new_n227), .ZN(new_n229));
  INV_X1    g028(.A(new_n202), .ZN(new_n230));
  NAND3_X1  g029(.A1(new_n229), .A2(new_n225), .A3(new_n230), .ZN(new_n231));
  NAND3_X1  g030(.A1(new_n215), .A2(KEYINPUT21), .A3(new_n218), .ZN(new_n232));
  XNOR2_X1  g031(.A(G15gat), .B(G22gat), .ZN(new_n233));
  OR2_X1    g032(.A1(new_n233), .A2(G1gat), .ZN(new_n234));
  NAND2_X1  g033(.A1(new_n234), .A2(KEYINPUT88), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n235), .A2(G8gat), .ZN(new_n236));
  INV_X1    g035(.A(KEYINPUT87), .ZN(new_n237));
  INV_X1    g036(.A(KEYINPUT16), .ZN(new_n238));
  NOR3_X1   g037(.A1(new_n237), .A2(new_n238), .A3(G1gat), .ZN(new_n239));
  OAI21_X1  g038(.A(new_n237), .B1(new_n238), .B2(G1gat), .ZN(new_n240));
  NAND2_X1  g039(.A1(new_n233), .A2(new_n240), .ZN(new_n241));
  OAI21_X1  g040(.A(new_n234), .B1(new_n239), .B2(new_n241), .ZN(new_n242));
  XNOR2_X1  g041(.A(new_n236), .B(new_n242), .ZN(new_n243));
  NAND2_X1  g042(.A1(new_n232), .A2(new_n243), .ZN(new_n244));
  XOR2_X1   g043(.A(KEYINPUT95), .B(KEYINPUT19), .Z(new_n245));
  XNOR2_X1  g044(.A(new_n244), .B(new_n245), .ZN(new_n246));
  AND3_X1   g045(.A1(new_n228), .A2(new_n231), .A3(new_n246), .ZN(new_n247));
  AOI21_X1  g046(.A(new_n246), .B1(new_n228), .B2(new_n231), .ZN(new_n248));
  NOR2_X1   g047(.A1(new_n247), .A2(new_n248), .ZN(new_n249));
  NAND2_X1  g048(.A1(G232gat), .A2(G233gat), .ZN(new_n250));
  XOR2_X1   g049(.A(new_n250), .B(KEYINPUT96), .Z(new_n251));
  INV_X1    g050(.A(KEYINPUT41), .ZN(new_n252));
  NAND2_X1  g051(.A1(new_n251), .A2(new_n252), .ZN(new_n253));
  XNOR2_X1  g052(.A(new_n253), .B(KEYINPUT97), .ZN(new_n254));
  XOR2_X1   g053(.A(G134gat), .B(G162gat), .Z(new_n255));
  XNOR2_X1  g054(.A(new_n254), .B(new_n255), .ZN(new_n256));
  INV_X1    g055(.A(new_n256), .ZN(new_n257));
  INV_X1    g056(.A(KEYINPUT15), .ZN(new_n258));
  INV_X1    g057(.A(G50gat), .ZN(new_n259));
  NAND2_X1  g058(.A1(new_n259), .A2(G43gat), .ZN(new_n260));
  INV_X1    g059(.A(KEYINPUT84), .ZN(new_n261));
  XNOR2_X1  g060(.A(new_n260), .B(new_n261), .ZN(new_n262));
  XNOR2_X1  g061(.A(KEYINPUT85), .B(G50gat), .ZN(new_n263));
  NOR2_X1   g062(.A1(new_n263), .A2(G43gat), .ZN(new_n264));
  OAI211_X1 g063(.A(KEYINPUT86), .B(new_n258), .C1(new_n262), .C2(new_n264), .ZN(new_n265));
  INV_X1    g064(.A(G43gat), .ZN(new_n266));
  NAND2_X1  g065(.A1(new_n266), .A2(G50gat), .ZN(new_n267));
  NAND3_X1  g066(.A1(new_n267), .A2(new_n260), .A3(KEYINPUT15), .ZN(new_n268));
  NAND2_X1  g067(.A1(new_n265), .A2(new_n268), .ZN(new_n269));
  XNOR2_X1  g068(.A(KEYINPUT14), .B(G29gat), .ZN(new_n270));
  INV_X1    g069(.A(G36gat), .ZN(new_n271));
  NAND2_X1  g070(.A1(new_n270), .A2(new_n271), .ZN(new_n272));
  INV_X1    g071(.A(G29gat), .ZN(new_n273));
  NAND2_X1  g072(.A1(new_n273), .A2(KEYINPUT14), .ZN(new_n274));
  OAI21_X1  g073(.A(new_n272), .B1(new_n271), .B2(new_n274), .ZN(new_n275));
  AND2_X1   g074(.A1(new_n269), .A2(new_n275), .ZN(new_n276));
  INV_X1    g075(.A(new_n268), .ZN(new_n277));
  OAI21_X1  g076(.A(new_n258), .B1(new_n262), .B2(new_n264), .ZN(new_n278));
  INV_X1    g077(.A(KEYINPUT86), .ZN(new_n279));
  NAND2_X1  g078(.A1(new_n278), .A2(new_n279), .ZN(new_n280));
  AOI21_X1  g079(.A(new_n277), .B1(new_n280), .B2(new_n275), .ZN(new_n281));
  OAI21_X1  g080(.A(KEYINPUT17), .B1(new_n276), .B2(new_n281), .ZN(new_n282));
  INV_X1    g081(.A(KEYINPUT17), .ZN(new_n283));
  NAND2_X1  g082(.A1(new_n269), .A2(new_n275), .ZN(new_n284));
  AND2_X1   g083(.A1(new_n280), .A2(new_n275), .ZN(new_n285));
  OAI211_X1 g084(.A(new_n283), .B(new_n284), .C1(new_n285), .C2(new_n277), .ZN(new_n286));
  INV_X1    g085(.A(G85gat), .ZN(new_n287));
  INV_X1    g086(.A(G92gat), .ZN(new_n288));
  OAI21_X1  g087(.A(KEYINPUT98), .B1(new_n287), .B2(new_n288), .ZN(new_n289));
  INV_X1    g088(.A(KEYINPUT98), .ZN(new_n290));
  NAND3_X1  g089(.A1(new_n290), .A2(G85gat), .A3(G92gat), .ZN(new_n291));
  NAND3_X1  g090(.A1(new_n289), .A2(KEYINPUT7), .A3(new_n291), .ZN(new_n292));
  NAND2_X1  g091(.A1(G99gat), .A2(G106gat), .ZN(new_n293));
  AOI22_X1  g092(.A1(KEYINPUT8), .A2(new_n293), .B1(new_n287), .B2(new_n288), .ZN(new_n294));
  OAI211_X1 g093(.A(new_n292), .B(new_n294), .C1(KEYINPUT7), .C2(new_n289), .ZN(new_n295));
  XNOR2_X1  g094(.A(G99gat), .B(G106gat), .ZN(new_n296));
  XNOR2_X1  g095(.A(new_n295), .B(new_n296), .ZN(new_n297));
  INV_X1    g096(.A(new_n297), .ZN(new_n298));
  NAND3_X1  g097(.A1(new_n282), .A2(new_n286), .A3(new_n298), .ZN(new_n299));
  NOR2_X1   g098(.A1(new_n251), .A2(new_n252), .ZN(new_n300));
  NOR2_X1   g099(.A1(new_n276), .A2(new_n281), .ZN(new_n301));
  AOI21_X1  g100(.A(new_n300), .B1(new_n301), .B2(new_n297), .ZN(new_n302));
  XOR2_X1   g101(.A(G190gat), .B(G218gat), .Z(new_n303));
  INV_X1    g102(.A(new_n303), .ZN(new_n304));
  NAND3_X1  g103(.A1(new_n299), .A2(new_n302), .A3(new_n304), .ZN(new_n305));
  INV_X1    g104(.A(new_n305), .ZN(new_n306));
  AOI21_X1  g105(.A(new_n304), .B1(new_n299), .B2(new_n302), .ZN(new_n307));
  OAI21_X1  g106(.A(new_n257), .B1(new_n306), .B2(new_n307), .ZN(new_n308));
  INV_X1    g107(.A(new_n307), .ZN(new_n309));
  NAND3_X1  g108(.A1(new_n309), .A2(new_n256), .A3(new_n305), .ZN(new_n310));
  NAND2_X1  g109(.A1(new_n308), .A2(new_n310), .ZN(new_n311));
  INV_X1    g110(.A(new_n311), .ZN(new_n312));
  XNOR2_X1  g111(.A(G120gat), .B(G148gat), .ZN(new_n313));
  XNOR2_X1  g112(.A(G176gat), .B(G204gat), .ZN(new_n314));
  XOR2_X1   g113(.A(new_n313), .B(new_n314), .Z(new_n315));
  INV_X1    g114(.A(new_n315), .ZN(new_n316));
  NAND2_X1  g115(.A1(G230gat), .A2(G233gat), .ZN(new_n317));
  INV_X1    g116(.A(new_n317), .ZN(new_n318));
  NAND3_X1  g117(.A1(new_n215), .A2(new_n218), .A3(new_n297), .ZN(new_n319));
  INV_X1    g118(.A(KEYINPUT10), .ZN(new_n320));
  OR2_X1    g119(.A1(new_n319), .A2(new_n320), .ZN(new_n321));
  XNOR2_X1  g120(.A(new_n213), .B(KEYINPUT94), .ZN(new_n322));
  XNOR2_X1  g121(.A(new_n216), .B(KEYINPUT93), .ZN(new_n323));
  OAI21_X1  g122(.A(new_n298), .B1(new_n322), .B2(new_n323), .ZN(new_n324));
  NAND3_X1  g123(.A1(new_n324), .A2(new_n320), .A3(new_n319), .ZN(new_n325));
  AOI21_X1  g124(.A(new_n318), .B1(new_n321), .B2(new_n325), .ZN(new_n326));
  AOI21_X1  g125(.A(new_n317), .B1(new_n324), .B2(new_n319), .ZN(new_n327));
  OAI21_X1  g126(.A(new_n316), .B1(new_n326), .B2(new_n327), .ZN(new_n328));
  NAND2_X1  g127(.A1(new_n321), .A2(new_n325), .ZN(new_n329));
  NAND2_X1  g128(.A1(new_n329), .A2(new_n317), .ZN(new_n330));
  NAND2_X1  g129(.A1(new_n330), .A2(new_n315), .ZN(new_n331));
  XNOR2_X1  g130(.A(new_n327), .B(KEYINPUT99), .ZN(new_n332));
  OAI21_X1  g131(.A(new_n328), .B1(new_n331), .B2(new_n332), .ZN(new_n333));
  INV_X1    g132(.A(new_n333), .ZN(new_n334));
  NAND3_X1  g133(.A1(new_n249), .A2(new_n312), .A3(new_n334), .ZN(new_n335));
  NAND3_X1  g134(.A1(new_n282), .A2(new_n286), .A3(new_n243), .ZN(new_n336));
  INV_X1    g135(.A(new_n243), .ZN(new_n337));
  NAND2_X1  g136(.A1(new_n301), .A2(new_n337), .ZN(new_n338));
  NAND2_X1  g137(.A1(G229gat), .A2(G233gat), .ZN(new_n339));
  NAND4_X1  g138(.A1(new_n336), .A2(new_n338), .A3(KEYINPUT18), .A4(new_n339), .ZN(new_n340));
  XOR2_X1   g139(.A(new_n339), .B(KEYINPUT13), .Z(new_n341));
  NOR2_X1   g140(.A1(new_n301), .A2(new_n337), .ZN(new_n342));
  NOR3_X1   g141(.A1(new_n243), .A2(new_n276), .A3(new_n281), .ZN(new_n343));
  OAI21_X1  g142(.A(new_n341), .B1(new_n342), .B2(new_n343), .ZN(new_n344));
  XNOR2_X1  g143(.A(G113gat), .B(G141gat), .ZN(new_n345));
  XNOR2_X1  g144(.A(new_n345), .B(G197gat), .ZN(new_n346));
  XOR2_X1   g145(.A(KEYINPUT11), .B(G169gat), .Z(new_n347));
  XNOR2_X1  g146(.A(new_n346), .B(new_n347), .ZN(new_n348));
  XNOR2_X1  g147(.A(new_n348), .B(KEYINPUT12), .ZN(new_n349));
  AND3_X1   g148(.A1(new_n340), .A2(new_n344), .A3(new_n349), .ZN(new_n350));
  NAND3_X1  g149(.A1(new_n336), .A2(new_n338), .A3(new_n339), .ZN(new_n351));
  XNOR2_X1  g150(.A(KEYINPUT89), .B(KEYINPUT18), .ZN(new_n352));
  NAND2_X1  g151(.A1(new_n351), .A2(new_n352), .ZN(new_n353));
  NAND2_X1  g152(.A1(new_n353), .A2(KEYINPUT90), .ZN(new_n354));
  INV_X1    g153(.A(KEYINPUT90), .ZN(new_n355));
  NAND3_X1  g154(.A1(new_n351), .A2(new_n355), .A3(new_n352), .ZN(new_n356));
  NAND3_X1  g155(.A1(new_n350), .A2(new_n354), .A3(new_n356), .ZN(new_n357));
  NAND3_X1  g156(.A1(new_n353), .A2(new_n344), .A3(new_n340), .ZN(new_n358));
  XNOR2_X1  g157(.A(new_n349), .B(KEYINPUT83), .ZN(new_n359));
  NAND2_X1  g158(.A1(new_n358), .A2(new_n359), .ZN(new_n360));
  AND2_X1   g159(.A1(new_n357), .A2(new_n360), .ZN(new_n361));
  INV_X1    g160(.A(new_n361), .ZN(new_n362));
  XOR2_X1   g161(.A(G1gat), .B(G29gat), .Z(new_n363));
  XNOR2_X1  g162(.A(KEYINPUT76), .B(KEYINPUT0), .ZN(new_n364));
  XNOR2_X1  g163(.A(new_n363), .B(new_n364), .ZN(new_n365));
  XNOR2_X1  g164(.A(G57gat), .B(G85gat), .ZN(new_n366));
  XNOR2_X1  g165(.A(new_n365), .B(new_n366), .ZN(new_n367));
  INV_X1    g166(.A(new_n367), .ZN(new_n368));
  NAND2_X1  g167(.A1(G225gat), .A2(G233gat), .ZN(new_n369));
  XNOR2_X1  g168(.A(G127gat), .B(G134gat), .ZN(new_n370));
  INV_X1    g169(.A(new_n370), .ZN(new_n371));
  INV_X1    g170(.A(G120gat), .ZN(new_n372));
  NAND2_X1  g171(.A1(new_n372), .A2(G113gat), .ZN(new_n373));
  INV_X1    g172(.A(G113gat), .ZN(new_n374));
  NAND2_X1  g173(.A1(new_n374), .A2(G120gat), .ZN(new_n375));
  AOI21_X1  g174(.A(KEYINPUT1), .B1(new_n373), .B2(new_n375), .ZN(new_n376));
  NAND3_X1  g175(.A1(new_n371), .A2(new_n376), .A3(KEYINPUT65), .ZN(new_n377));
  OAI21_X1  g176(.A(new_n370), .B1(new_n376), .B2(KEYINPUT65), .ZN(new_n378));
  INV_X1    g177(.A(KEYINPUT65), .ZN(new_n379));
  AOI211_X1 g178(.A(new_n379), .B(KEYINPUT1), .C1(new_n373), .C2(new_n375), .ZN(new_n380));
  OAI21_X1  g179(.A(new_n377), .B1(new_n378), .B2(new_n380), .ZN(new_n381));
  INV_X1    g180(.A(G141gat), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n382), .A2(G148gat), .ZN(new_n383));
  INV_X1    g182(.A(G148gat), .ZN(new_n384));
  NAND2_X1  g183(.A1(new_n384), .A2(G141gat), .ZN(new_n385));
  NAND2_X1  g184(.A1(G155gat), .A2(G162gat), .ZN(new_n386));
  AOI22_X1  g185(.A1(new_n383), .A2(new_n385), .B1(KEYINPUT2), .B2(new_n386), .ZN(new_n387));
  INV_X1    g186(.A(new_n386), .ZN(new_n388));
  NOR2_X1   g187(.A1(G155gat), .A2(G162gat), .ZN(new_n389));
  OAI21_X1  g188(.A(KEYINPUT73), .B1(new_n388), .B2(new_n389), .ZN(new_n390));
  OR2_X1    g189(.A1(G155gat), .A2(G162gat), .ZN(new_n391));
  INV_X1    g190(.A(KEYINPUT73), .ZN(new_n392));
  NAND3_X1  g191(.A1(new_n391), .A2(new_n392), .A3(new_n386), .ZN(new_n393));
  NAND3_X1  g192(.A1(new_n387), .A2(new_n390), .A3(new_n393), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n391), .A2(new_n386), .ZN(new_n395));
  XNOR2_X1  g194(.A(G141gat), .B(G148gat), .ZN(new_n396));
  INV_X1    g195(.A(KEYINPUT2), .ZN(new_n397));
  AOI21_X1  g196(.A(new_n397), .B1(G155gat), .B2(G162gat), .ZN(new_n398));
  OAI211_X1 g197(.A(new_n395), .B(KEYINPUT73), .C1(new_n396), .C2(new_n398), .ZN(new_n399));
  NAND2_X1  g198(.A1(new_n394), .A2(new_n399), .ZN(new_n400));
  NAND2_X1  g199(.A1(new_n381), .A2(new_n400), .ZN(new_n401));
  NAND2_X1  g200(.A1(new_n401), .A2(KEYINPUT4), .ZN(new_n402));
  INV_X1    g201(.A(KEYINPUT4), .ZN(new_n403));
  NAND3_X1  g202(.A1(new_n381), .A2(new_n403), .A3(new_n400), .ZN(new_n404));
  INV_X1    g203(.A(KEYINPUT74), .ZN(new_n405));
  NAND2_X1  g204(.A1(new_n400), .A2(new_n405), .ZN(new_n406));
  NAND3_X1  g205(.A1(new_n394), .A2(KEYINPUT74), .A3(new_n399), .ZN(new_n407));
  NAND3_X1  g206(.A1(new_n406), .A2(KEYINPUT3), .A3(new_n407), .ZN(new_n408));
  XNOR2_X1  g207(.A(KEYINPUT75), .B(KEYINPUT3), .ZN(new_n409));
  AOI21_X1  g208(.A(new_n409), .B1(new_n394), .B2(new_n399), .ZN(new_n410));
  NOR2_X1   g209(.A1(new_n381), .A2(new_n410), .ZN(new_n411));
  AOI22_X1  g210(.A1(new_n402), .A2(new_n404), .B1(new_n408), .B2(new_n411), .ZN(new_n412));
  INV_X1    g211(.A(new_n369), .ZN(new_n413));
  INV_X1    g212(.A(new_n407), .ZN(new_n414));
  AOI21_X1  g213(.A(KEYINPUT74), .B1(new_n394), .B2(new_n399), .ZN(new_n415));
  NOR3_X1   g214(.A1(new_n414), .A2(new_n381), .A3(new_n415), .ZN(new_n416));
  INV_X1    g215(.A(new_n401), .ZN(new_n417));
  OAI21_X1  g216(.A(new_n413), .B1(new_n416), .B2(new_n417), .ZN(new_n418));
  AOI22_X1  g217(.A1(new_n369), .A2(new_n412), .B1(new_n418), .B2(KEYINPUT5), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n402), .A2(new_n404), .ZN(new_n420));
  NAND2_X1  g219(.A1(new_n408), .A2(new_n411), .ZN(new_n421));
  AND4_X1   g220(.A1(KEYINPUT5), .A2(new_n420), .A3(new_n421), .A4(new_n369), .ZN(new_n422));
  OAI21_X1  g221(.A(new_n368), .B1(new_n419), .B2(new_n422), .ZN(new_n423));
  INV_X1    g222(.A(KEYINPUT6), .ZN(new_n424));
  NAND3_X1  g223(.A1(new_n412), .A2(KEYINPUT5), .A3(new_n369), .ZN(new_n425));
  AND3_X1   g224(.A1(new_n420), .A2(new_n421), .A3(new_n369), .ZN(new_n426));
  INV_X1    g225(.A(KEYINPUT5), .ZN(new_n427));
  NAND2_X1  g226(.A1(new_n406), .A2(new_n407), .ZN(new_n428));
  OAI21_X1  g227(.A(new_n401), .B1(new_n428), .B2(new_n381), .ZN(new_n429));
  AOI21_X1  g228(.A(new_n427), .B1(new_n429), .B2(new_n413), .ZN(new_n430));
  OAI211_X1 g229(.A(new_n425), .B(new_n367), .C1(new_n426), .C2(new_n430), .ZN(new_n431));
  NAND3_X1  g230(.A1(new_n423), .A2(new_n424), .A3(new_n431), .ZN(new_n432));
  NOR2_X1   g231(.A1(new_n419), .A2(new_n422), .ZN(new_n433));
  NAND3_X1  g232(.A1(new_n433), .A2(KEYINPUT6), .A3(new_n367), .ZN(new_n434));
  AND2_X1   g233(.A1(G211gat), .A2(G218gat), .ZN(new_n435));
  OR2_X1    g234(.A1(new_n435), .A2(KEYINPUT22), .ZN(new_n436));
  AND2_X1   g235(.A1(KEYINPUT67), .A2(G197gat), .ZN(new_n437));
  NOR2_X1   g236(.A1(KEYINPUT67), .A2(G197gat), .ZN(new_n438));
  INV_X1    g237(.A(G204gat), .ZN(new_n439));
  NOR3_X1   g238(.A1(new_n437), .A2(new_n438), .A3(new_n439), .ZN(new_n440));
  INV_X1    g239(.A(KEYINPUT67), .ZN(new_n441));
  INV_X1    g240(.A(G197gat), .ZN(new_n442));
  NAND2_X1  g241(.A1(new_n441), .A2(new_n442), .ZN(new_n443));
  NAND2_X1  g242(.A1(KEYINPUT67), .A2(G197gat), .ZN(new_n444));
  AOI21_X1  g243(.A(G204gat), .B1(new_n443), .B2(new_n444), .ZN(new_n445));
  OAI21_X1  g244(.A(new_n436), .B1(new_n440), .B2(new_n445), .ZN(new_n446));
  NOR2_X1   g245(.A1(G211gat), .A2(G218gat), .ZN(new_n447));
  NOR2_X1   g246(.A1(new_n435), .A2(new_n447), .ZN(new_n448));
  NAND2_X1  g247(.A1(new_n446), .A2(new_n448), .ZN(new_n449));
  OAI21_X1  g248(.A(new_n439), .B1(new_n437), .B2(new_n438), .ZN(new_n450));
  NAND3_X1  g249(.A1(new_n443), .A2(G204gat), .A3(new_n444), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n450), .A2(new_n451), .ZN(new_n452));
  INV_X1    g251(.A(new_n448), .ZN(new_n453));
  NAND3_X1  g252(.A1(new_n452), .A2(new_n453), .A3(new_n436), .ZN(new_n454));
  NAND2_X1  g253(.A1(new_n449), .A2(new_n454), .ZN(new_n455));
  NAND2_X1  g254(.A1(G169gat), .A2(G176gat), .ZN(new_n456));
  INV_X1    g255(.A(KEYINPUT64), .ZN(new_n457));
  NAND2_X1  g256(.A1(new_n456), .A2(new_n457), .ZN(new_n458));
  NAND3_X1  g257(.A1(KEYINPUT64), .A2(G169gat), .A3(G176gat), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  NOR3_X1   g259(.A1(KEYINPUT26), .A2(G169gat), .A3(G176gat), .ZN(new_n461));
  INV_X1    g260(.A(new_n461), .ZN(new_n462));
  OAI21_X1  g261(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n463));
  NAND3_X1  g262(.A1(new_n460), .A2(new_n462), .A3(new_n463), .ZN(new_n464));
  INV_X1    g263(.A(G183gat), .ZN(new_n465));
  INV_X1    g264(.A(G190gat), .ZN(new_n466));
  NOR2_X1   g265(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  INV_X1    g266(.A(new_n467), .ZN(new_n468));
  XNOR2_X1  g267(.A(KEYINPUT27), .B(G183gat), .ZN(new_n469));
  AOI21_X1  g268(.A(KEYINPUT28), .B1(new_n469), .B2(new_n466), .ZN(new_n470));
  NAND2_X1  g269(.A1(new_n465), .A2(KEYINPUT27), .ZN(new_n471));
  INV_X1    g270(.A(KEYINPUT27), .ZN(new_n472));
  NAND2_X1  g271(.A1(new_n472), .A2(G183gat), .ZN(new_n473));
  AND4_X1   g272(.A1(KEYINPUT28), .A2(new_n471), .A3(new_n473), .A4(new_n466), .ZN(new_n474));
  OAI211_X1 g273(.A(new_n464), .B(new_n468), .C1(new_n470), .C2(new_n474), .ZN(new_n475));
  OAI21_X1  g274(.A(G190gat), .B1(KEYINPUT24), .B2(G183gat), .ZN(new_n476));
  AND2_X1   g275(.A1(KEYINPUT24), .A2(G183gat), .ZN(new_n477));
  NOR2_X1   g276(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  INV_X1    g277(.A(KEYINPUT24), .ZN(new_n479));
  NOR3_X1   g278(.A1(new_n479), .A2(new_n465), .A3(G190gat), .ZN(new_n480));
  NOR2_X1   g279(.A1(new_n478), .A2(new_n480), .ZN(new_n481));
  OAI21_X1  g280(.A(KEYINPUT23), .B1(G169gat), .B2(G176gat), .ZN(new_n482));
  INV_X1    g281(.A(KEYINPUT23), .ZN(new_n483));
  INV_X1    g282(.A(G169gat), .ZN(new_n484));
  INV_X1    g283(.A(G176gat), .ZN(new_n485));
  NAND3_X1  g284(.A1(new_n483), .A2(new_n484), .A3(new_n485), .ZN(new_n486));
  AOI22_X1  g285(.A1(new_n482), .A2(new_n486), .B1(new_n458), .B2(new_n459), .ZN(new_n487));
  AND3_X1   g286(.A1(new_n481), .A2(new_n487), .A3(KEYINPUT25), .ZN(new_n488));
  AOI21_X1  g287(.A(KEYINPUT25), .B1(new_n481), .B2(new_n487), .ZN(new_n489));
  OAI21_X1  g288(.A(new_n475), .B1(new_n488), .B2(new_n489), .ZN(new_n490));
  NAND2_X1  g289(.A1(G226gat), .A2(G233gat), .ZN(new_n491));
  INV_X1    g290(.A(new_n491), .ZN(new_n492));
  NAND2_X1  g291(.A1(new_n490), .A2(new_n492), .ZN(new_n493));
  NAND2_X1  g292(.A1(new_n493), .A2(KEYINPUT69), .ZN(new_n494));
  INV_X1    g293(.A(KEYINPUT25), .ZN(new_n495));
  NAND2_X1  g294(.A1(new_n479), .A2(new_n465), .ZN(new_n496));
  NAND2_X1  g295(.A1(KEYINPUT24), .A2(G183gat), .ZN(new_n497));
  NAND3_X1  g296(.A1(new_n496), .A2(G190gat), .A3(new_n497), .ZN(new_n498));
  NAND2_X1  g297(.A1(new_n476), .A2(new_n477), .ZN(new_n499));
  NAND2_X1  g298(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  INV_X1    g299(.A(new_n482), .ZN(new_n501));
  NOR3_X1   g300(.A1(KEYINPUT23), .A2(G169gat), .A3(G176gat), .ZN(new_n502));
  AND3_X1   g301(.A1(KEYINPUT64), .A2(G169gat), .A3(G176gat), .ZN(new_n503));
  AOI21_X1  g302(.A(KEYINPUT64), .B1(G169gat), .B2(G176gat), .ZN(new_n504));
  OAI22_X1  g303(.A1(new_n501), .A2(new_n502), .B1(new_n503), .B2(new_n504), .ZN(new_n505));
  OAI21_X1  g304(.A(new_n495), .B1(new_n500), .B2(new_n505), .ZN(new_n506));
  NAND3_X1  g305(.A1(new_n481), .A2(new_n487), .A3(KEYINPUT25), .ZN(new_n507));
  NAND2_X1  g306(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  AOI21_X1  g307(.A(new_n491), .B1(new_n508), .B2(new_n475), .ZN(new_n509));
  INV_X1    g308(.A(KEYINPUT29), .ZN(new_n510));
  NAND2_X1  g309(.A1(new_n490), .A2(new_n510), .ZN(new_n511));
  AOI21_X1  g310(.A(new_n509), .B1(new_n511), .B2(new_n491), .ZN(new_n512));
  OAI211_X1 g311(.A(new_n455), .B(new_n494), .C1(new_n512), .C2(KEYINPUT69), .ZN(new_n513));
  INV_X1    g312(.A(KEYINPUT68), .ZN(new_n514));
  OAI21_X1  g313(.A(new_n514), .B1(new_n512), .B2(new_n455), .ZN(new_n515));
  NAND3_X1  g314(.A1(new_n471), .A2(new_n473), .A3(new_n466), .ZN(new_n516));
  INV_X1    g315(.A(KEYINPUT28), .ZN(new_n517));
  NAND2_X1  g316(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  NAND3_X1  g317(.A1(new_n469), .A2(KEYINPUT28), .A3(new_n466), .ZN(new_n519));
  NAND2_X1  g318(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  INV_X1    g319(.A(new_n463), .ZN(new_n521));
  NOR2_X1   g320(.A1(new_n521), .A2(new_n461), .ZN(new_n522));
  AOI21_X1  g321(.A(new_n467), .B1(new_n522), .B2(new_n460), .ZN(new_n523));
  AOI22_X1  g322(.A1(new_n506), .A2(new_n507), .B1(new_n520), .B2(new_n523), .ZN(new_n524));
  OAI21_X1  g323(.A(new_n491), .B1(new_n524), .B2(KEYINPUT29), .ZN(new_n525));
  NAND2_X1  g324(.A1(new_n525), .A2(new_n493), .ZN(new_n526));
  INV_X1    g325(.A(new_n455), .ZN(new_n527));
  NAND3_X1  g326(.A1(new_n526), .A2(KEYINPUT68), .A3(new_n527), .ZN(new_n528));
  XOR2_X1   g327(.A(G8gat), .B(G36gat), .Z(new_n529));
  XNOR2_X1  g328(.A(new_n529), .B(KEYINPUT70), .ZN(new_n530));
  XNOR2_X1  g329(.A(G64gat), .B(G92gat), .ZN(new_n531));
  XNOR2_X1  g330(.A(new_n530), .B(new_n531), .ZN(new_n532));
  NAND4_X1  g331(.A1(new_n513), .A2(new_n515), .A3(new_n528), .A4(new_n532), .ZN(new_n533));
  AND3_X1   g332(.A1(new_n432), .A2(new_n434), .A3(new_n533), .ZN(new_n534));
  INV_X1    g333(.A(KEYINPUT37), .ZN(new_n535));
  NAND4_X1  g334(.A1(new_n513), .A2(new_n515), .A3(new_n535), .A4(new_n528), .ZN(new_n536));
  INV_X1    g335(.A(new_n532), .ZN(new_n537));
  NAND2_X1  g336(.A1(new_n536), .A2(new_n537), .ZN(new_n538));
  AOI21_X1  g337(.A(KEYINPUT68), .B1(new_n526), .B2(new_n527), .ZN(new_n539));
  AOI211_X1 g338(.A(new_n514), .B(new_n455), .C1(new_n525), .C2(new_n493), .ZN(new_n540));
  NOR2_X1   g339(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  AOI21_X1  g340(.A(new_n535), .B1(new_n541), .B2(new_n513), .ZN(new_n542));
  OAI21_X1  g341(.A(KEYINPUT38), .B1(new_n538), .B2(new_n542), .ZN(new_n543));
  INV_X1    g342(.A(KEYINPUT38), .ZN(new_n544));
  XNOR2_X1  g343(.A(new_n532), .B(KEYINPUT71), .ZN(new_n545));
  AND3_X1   g344(.A1(new_n536), .A2(new_n544), .A3(new_n545), .ZN(new_n546));
  NOR2_X1   g345(.A1(new_n526), .A2(new_n527), .ZN(new_n547));
  AOI21_X1  g346(.A(KEYINPUT69), .B1(new_n525), .B2(new_n493), .ZN(new_n548));
  AND2_X1   g347(.A1(new_n493), .A2(KEYINPUT69), .ZN(new_n549));
  OAI21_X1  g348(.A(new_n527), .B1(new_n548), .B2(new_n549), .ZN(new_n550));
  INV_X1    g349(.A(KEYINPUT80), .ZN(new_n551));
  AOI21_X1  g350(.A(new_n547), .B1(new_n550), .B2(new_n551), .ZN(new_n552));
  OAI211_X1 g351(.A(KEYINPUT80), .B(new_n527), .C1(new_n548), .C2(new_n549), .ZN(new_n553));
  AOI21_X1  g352(.A(new_n535), .B1(new_n552), .B2(new_n553), .ZN(new_n554));
  OAI21_X1  g353(.A(new_n546), .B1(new_n554), .B2(KEYINPUT81), .ZN(new_n555));
  INV_X1    g354(.A(KEYINPUT81), .ZN(new_n556));
  AOI211_X1 g355(.A(new_n556), .B(new_n535), .C1(new_n552), .C2(new_n553), .ZN(new_n557));
  OAI211_X1 g356(.A(new_n534), .B(new_n543), .C1(new_n555), .C2(new_n557), .ZN(new_n558));
  XNOR2_X1  g357(.A(G78gat), .B(G106gat), .ZN(new_n559));
  XNOR2_X1  g358(.A(new_n559), .B(G22gat), .ZN(new_n560));
  INV_X1    g359(.A(new_n560), .ZN(new_n561));
  XNOR2_X1  g360(.A(KEYINPUT31), .B(G50gat), .ZN(new_n562));
  INV_X1    g361(.A(new_n562), .ZN(new_n563));
  OAI21_X1  g362(.A(new_n527), .B1(KEYINPUT29), .B2(new_n410), .ZN(new_n564));
  INV_X1    g363(.A(G228gat), .ZN(new_n565));
  INV_X1    g364(.A(G233gat), .ZN(new_n566));
  NOR2_X1   g365(.A1(new_n565), .A2(new_n566), .ZN(new_n567));
  INV_X1    g366(.A(new_n567), .ZN(new_n568));
  NAND2_X1  g367(.A1(new_n564), .A2(new_n568), .ZN(new_n569));
  INV_X1    g368(.A(new_n569), .ZN(new_n570));
  NAND3_X1  g369(.A1(new_n449), .A2(KEYINPUT77), .A3(new_n454), .ZN(new_n571));
  AOI21_X1  g370(.A(new_n453), .B1(new_n452), .B2(new_n436), .ZN(new_n572));
  INV_X1    g371(.A(KEYINPUT77), .ZN(new_n573));
  AOI21_X1  g372(.A(KEYINPUT29), .B1(new_n572), .B2(new_n573), .ZN(new_n574));
  INV_X1    g373(.A(KEYINPUT78), .ZN(new_n575));
  AND3_X1   g374(.A1(new_n571), .A2(new_n574), .A3(new_n575), .ZN(new_n576));
  AOI21_X1  g375(.A(new_n575), .B1(new_n571), .B2(new_n574), .ZN(new_n577));
  NOR3_X1   g376(.A1(new_n576), .A2(new_n577), .A3(new_n409), .ZN(new_n578));
  OAI21_X1  g377(.A(new_n570), .B1(new_n578), .B2(new_n400), .ZN(new_n579));
  NAND2_X1  g378(.A1(new_n455), .A2(new_n510), .ZN(new_n580));
  INV_X1    g379(.A(KEYINPUT3), .ZN(new_n581));
  AOI21_X1  g380(.A(new_n428), .B1(new_n580), .B2(new_n581), .ZN(new_n582));
  NOR2_X1   g381(.A1(new_n410), .A2(KEYINPUT29), .ZN(new_n583));
  NOR2_X1   g382(.A1(new_n583), .A2(new_n455), .ZN(new_n584));
  OAI21_X1  g383(.A(new_n567), .B1(new_n582), .B2(new_n584), .ZN(new_n585));
  AOI21_X1  g384(.A(new_n563), .B1(new_n579), .B2(new_n585), .ZN(new_n586));
  AND3_X1   g385(.A1(new_n452), .A2(new_n453), .A3(new_n436), .ZN(new_n587));
  NOR3_X1   g386(.A1(new_n587), .A2(new_n572), .A3(new_n573), .ZN(new_n588));
  NAND3_X1  g387(.A1(new_n446), .A2(new_n573), .A3(new_n448), .ZN(new_n589));
  NAND2_X1  g388(.A1(new_n589), .A2(new_n510), .ZN(new_n590));
  OAI21_X1  g389(.A(KEYINPUT78), .B1(new_n588), .B2(new_n590), .ZN(new_n591));
  INV_X1    g390(.A(new_n409), .ZN(new_n592));
  NAND3_X1  g391(.A1(new_n571), .A2(new_n574), .A3(new_n575), .ZN(new_n593));
  NAND3_X1  g392(.A1(new_n591), .A2(new_n592), .A3(new_n593), .ZN(new_n594));
  INV_X1    g393(.A(new_n400), .ZN(new_n595));
  AOI21_X1  g394(.A(new_n569), .B1(new_n594), .B2(new_n595), .ZN(new_n596));
  NAND2_X1  g395(.A1(new_n580), .A2(new_n581), .ZN(new_n597));
  INV_X1    g396(.A(new_n428), .ZN(new_n598));
  NAND2_X1  g397(.A1(new_n597), .A2(new_n598), .ZN(new_n599));
  AOI21_X1  g398(.A(new_n568), .B1(new_n599), .B2(new_n564), .ZN(new_n600));
  NOR3_X1   g399(.A1(new_n596), .A2(new_n600), .A3(new_n562), .ZN(new_n601));
  OAI21_X1  g400(.A(new_n561), .B1(new_n586), .B2(new_n601), .ZN(new_n602));
  OAI21_X1  g401(.A(new_n562), .B1(new_n596), .B2(new_n600), .ZN(new_n603));
  NOR2_X1   g402(.A1(new_n577), .A2(new_n409), .ZN(new_n604));
  AOI21_X1  g403(.A(new_n400), .B1(new_n604), .B2(new_n593), .ZN(new_n605));
  OAI211_X1 g404(.A(new_n585), .B(new_n563), .C1(new_n605), .C2(new_n569), .ZN(new_n606));
  NAND3_X1  g405(.A1(new_n603), .A2(new_n606), .A3(new_n560), .ZN(new_n607));
  NAND2_X1  g406(.A1(new_n602), .A2(new_n607), .ZN(new_n608));
  NAND2_X1  g407(.A1(new_n533), .A2(KEYINPUT30), .ZN(new_n609));
  INV_X1    g408(.A(KEYINPUT30), .ZN(new_n610));
  NAND4_X1  g409(.A1(new_n541), .A2(new_n610), .A3(new_n513), .A4(new_n532), .ZN(new_n611));
  NAND2_X1  g410(.A1(new_n609), .A2(new_n611), .ZN(new_n612));
  INV_X1    g411(.A(KEYINPUT72), .ZN(new_n613));
  NAND3_X1  g412(.A1(new_n513), .A2(new_n515), .A3(new_n528), .ZN(new_n614));
  AOI21_X1  g413(.A(new_n613), .B1(new_n614), .B2(new_n545), .ZN(new_n615));
  AND3_X1   g414(.A1(new_n614), .A2(new_n613), .A3(new_n545), .ZN(new_n616));
  OAI21_X1  g415(.A(new_n612), .B1(new_n615), .B2(new_n616), .ZN(new_n617));
  NAND2_X1  g416(.A1(new_n420), .A2(new_n421), .ZN(new_n618));
  NAND2_X1  g417(.A1(new_n618), .A2(new_n413), .ZN(new_n619));
  INV_X1    g418(.A(KEYINPUT39), .ZN(new_n620));
  NOR2_X1   g419(.A1(new_n416), .A2(new_n417), .ZN(new_n621));
  AOI21_X1  g420(.A(new_n620), .B1(new_n621), .B2(new_n369), .ZN(new_n622));
  AOI21_X1  g421(.A(new_n367), .B1(new_n619), .B2(new_n622), .ZN(new_n623));
  XOR2_X1   g422(.A(KEYINPUT79), .B(KEYINPUT39), .Z(new_n624));
  NAND3_X1  g423(.A1(new_n618), .A2(new_n413), .A3(new_n624), .ZN(new_n625));
  NAND3_X1  g424(.A1(new_n623), .A2(KEYINPUT40), .A3(new_n625), .ZN(new_n626));
  NAND2_X1  g425(.A1(new_n626), .A2(new_n431), .ZN(new_n627));
  AOI21_X1  g426(.A(KEYINPUT40), .B1(new_n623), .B2(new_n625), .ZN(new_n628));
  NOR2_X1   g427(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  AOI21_X1  g428(.A(new_n608), .B1(new_n617), .B2(new_n629), .ZN(new_n630));
  NAND2_X1  g429(.A1(new_n558), .A2(new_n630), .ZN(new_n631));
  NAND2_X1  g430(.A1(new_n614), .A2(new_n545), .ZN(new_n632));
  NAND2_X1  g431(.A1(new_n632), .A2(KEYINPUT72), .ZN(new_n633));
  NAND3_X1  g432(.A1(new_n614), .A2(new_n613), .A3(new_n545), .ZN(new_n634));
  NAND2_X1  g433(.A1(new_n633), .A2(new_n634), .ZN(new_n635));
  NAND2_X1  g434(.A1(new_n432), .A2(new_n434), .ZN(new_n636));
  NAND3_X1  g435(.A1(new_n635), .A2(new_n636), .A3(new_n612), .ZN(new_n637));
  NAND2_X1  g436(.A1(new_n637), .A2(new_n608), .ZN(new_n638));
  INV_X1    g437(.A(KEYINPUT66), .ZN(new_n639));
  INV_X1    g438(.A(KEYINPUT36), .ZN(new_n640));
  NAND2_X1  g439(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  NAND2_X1  g440(.A1(KEYINPUT66), .A2(KEYINPUT36), .ZN(new_n642));
  INV_X1    g441(.A(new_n381), .ZN(new_n643));
  NAND2_X1  g442(.A1(new_n490), .A2(new_n643), .ZN(new_n644));
  NAND2_X1  g443(.A1(G227gat), .A2(G233gat), .ZN(new_n645));
  NAND3_X1  g444(.A1(new_n508), .A2(new_n381), .A3(new_n475), .ZN(new_n646));
  NAND3_X1  g445(.A1(new_n644), .A2(new_n645), .A3(new_n646), .ZN(new_n647));
  NAND2_X1  g446(.A1(new_n647), .A2(KEYINPUT34), .ZN(new_n648));
  INV_X1    g447(.A(KEYINPUT34), .ZN(new_n649));
  NAND4_X1  g448(.A1(new_n644), .A2(new_n649), .A3(new_n645), .A4(new_n646), .ZN(new_n650));
  NAND2_X1  g449(.A1(new_n648), .A2(new_n650), .ZN(new_n651));
  XOR2_X1   g450(.A(G15gat), .B(G43gat), .Z(new_n652));
  XNOR2_X1  g451(.A(G71gat), .B(G99gat), .ZN(new_n653));
  XNOR2_X1  g452(.A(new_n652), .B(new_n653), .ZN(new_n654));
  INV_X1    g453(.A(new_n654), .ZN(new_n655));
  INV_X1    g454(.A(new_n645), .ZN(new_n656));
  AND3_X1   g455(.A1(new_n508), .A2(new_n381), .A3(new_n475), .ZN(new_n657));
  AOI21_X1  g456(.A(new_n381), .B1(new_n508), .B2(new_n475), .ZN(new_n658));
  OAI21_X1  g457(.A(new_n656), .B1(new_n657), .B2(new_n658), .ZN(new_n659));
  INV_X1    g458(.A(KEYINPUT33), .ZN(new_n660));
  AOI21_X1  g459(.A(new_n655), .B1(new_n659), .B2(new_n660), .ZN(new_n661));
  NAND2_X1  g460(.A1(new_n651), .A2(new_n661), .ZN(new_n662));
  AOI21_X1  g461(.A(new_n645), .B1(new_n644), .B2(new_n646), .ZN(new_n663));
  OAI21_X1  g462(.A(new_n654), .B1(new_n663), .B2(KEYINPUT33), .ZN(new_n664));
  NAND3_X1  g463(.A1(new_n664), .A2(new_n648), .A3(new_n650), .ZN(new_n665));
  NAND2_X1  g464(.A1(new_n659), .A2(KEYINPUT32), .ZN(new_n666));
  INV_X1    g465(.A(new_n666), .ZN(new_n667));
  NAND3_X1  g466(.A1(new_n662), .A2(new_n665), .A3(new_n667), .ZN(new_n668));
  INV_X1    g467(.A(new_n668), .ZN(new_n669));
  AOI21_X1  g468(.A(new_n667), .B1(new_n662), .B2(new_n665), .ZN(new_n670));
  OAI211_X1 g469(.A(new_n641), .B(new_n642), .C1(new_n669), .C2(new_n670), .ZN(new_n671));
  AOI21_X1  g470(.A(new_n664), .B1(new_n648), .B2(new_n650), .ZN(new_n672));
  NOR2_X1   g471(.A1(new_n651), .A2(new_n661), .ZN(new_n673));
  OAI21_X1  g472(.A(new_n666), .B1(new_n672), .B2(new_n673), .ZN(new_n674));
  NAND4_X1  g473(.A1(new_n674), .A2(new_n639), .A3(new_n640), .A4(new_n668), .ZN(new_n675));
  AND2_X1   g474(.A1(new_n671), .A2(new_n675), .ZN(new_n676));
  NAND3_X1  g475(.A1(new_n631), .A2(new_n638), .A3(new_n676), .ZN(new_n677));
  INV_X1    g476(.A(KEYINPUT82), .ZN(new_n678));
  NAND2_X1  g477(.A1(new_n674), .A2(new_n668), .ZN(new_n679));
  AND3_X1   g478(.A1(new_n603), .A2(new_n606), .A3(new_n560), .ZN(new_n680));
  AOI21_X1  g479(.A(new_n560), .B1(new_n603), .B2(new_n606), .ZN(new_n681));
  NOR3_X1   g480(.A1(new_n679), .A2(new_n680), .A3(new_n681), .ZN(new_n682));
  INV_X1    g481(.A(KEYINPUT35), .ZN(new_n683));
  AOI22_X1  g482(.A1(new_n633), .A2(new_n634), .B1(new_n609), .B2(new_n611), .ZN(new_n684));
  NAND4_X1  g483(.A1(new_n682), .A2(new_n683), .A3(new_n636), .A4(new_n684), .ZN(new_n685));
  NAND4_X1  g484(.A1(new_n602), .A2(new_n607), .A3(new_n668), .A4(new_n674), .ZN(new_n686));
  OAI21_X1  g485(.A(KEYINPUT35), .B1(new_n637), .B2(new_n686), .ZN(new_n687));
  NAND2_X1  g486(.A1(new_n685), .A2(new_n687), .ZN(new_n688));
  AND3_X1   g487(.A1(new_n677), .A2(new_n678), .A3(new_n688), .ZN(new_n689));
  AOI21_X1  g488(.A(new_n678), .B1(new_n677), .B2(new_n688), .ZN(new_n690));
  OAI21_X1  g489(.A(new_n362), .B1(new_n689), .B2(new_n690), .ZN(new_n691));
  NAND2_X1  g490(.A1(new_n691), .A2(KEYINPUT91), .ZN(new_n692));
  AND2_X1   g491(.A1(new_n558), .A2(new_n630), .ZN(new_n693));
  NAND2_X1  g492(.A1(new_n638), .A2(new_n676), .ZN(new_n694));
  OAI21_X1  g493(.A(new_n688), .B1(new_n693), .B2(new_n694), .ZN(new_n695));
  NAND2_X1  g494(.A1(new_n695), .A2(KEYINPUT82), .ZN(new_n696));
  NAND3_X1  g495(.A1(new_n677), .A2(new_n678), .A3(new_n688), .ZN(new_n697));
  NAND2_X1  g496(.A1(new_n696), .A2(new_n697), .ZN(new_n698));
  INV_X1    g497(.A(KEYINPUT91), .ZN(new_n699));
  NAND3_X1  g498(.A1(new_n698), .A2(new_n699), .A3(new_n362), .ZN(new_n700));
  AOI21_X1  g499(.A(new_n335), .B1(new_n692), .B2(new_n700), .ZN(new_n701));
  INV_X1    g500(.A(new_n636), .ZN(new_n702));
  NAND2_X1  g501(.A1(new_n701), .A2(new_n702), .ZN(new_n703));
  XNOR2_X1  g502(.A(new_n703), .B(G1gat), .ZN(G1324gat));
  XOR2_X1   g503(.A(KEYINPUT16), .B(G8gat), .Z(new_n705));
  NAND3_X1  g504(.A1(new_n701), .A2(new_n617), .A3(new_n705), .ZN(new_n706));
  INV_X1    g505(.A(KEYINPUT42), .ZN(new_n707));
  OR2_X1    g506(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  INV_X1    g507(.A(new_n701), .ZN(new_n709));
  OAI21_X1  g508(.A(G8gat), .B1(new_n709), .B2(new_n684), .ZN(new_n710));
  NAND2_X1  g509(.A1(new_n706), .A2(new_n707), .ZN(new_n711));
  NAND3_X1  g510(.A1(new_n708), .A2(new_n710), .A3(new_n711), .ZN(G1325gat));
  OR3_X1    g511(.A1(new_n709), .A2(G15gat), .A3(new_n679), .ZN(new_n713));
  OAI21_X1  g512(.A(G15gat), .B1(new_n709), .B2(new_n676), .ZN(new_n714));
  NAND2_X1  g513(.A1(new_n713), .A2(new_n714), .ZN(G1326gat));
  NAND2_X1  g514(.A1(new_n701), .A2(new_n608), .ZN(new_n716));
  XNOR2_X1  g515(.A(KEYINPUT43), .B(G22gat), .ZN(new_n717));
  XNOR2_X1  g516(.A(new_n716), .B(new_n717), .ZN(G1327gat));
  INV_X1    g517(.A(new_n249), .ZN(new_n719));
  NAND3_X1  g518(.A1(new_n719), .A2(new_n311), .A3(new_n334), .ZN(new_n720));
  AOI21_X1  g519(.A(new_n720), .B1(new_n692), .B2(new_n700), .ZN(new_n721));
  NAND3_X1  g520(.A1(new_n721), .A2(new_n273), .A3(new_n702), .ZN(new_n722));
  XNOR2_X1  g521(.A(new_n722), .B(KEYINPUT45), .ZN(new_n723));
  NAND3_X1  g522(.A1(new_n698), .A2(KEYINPUT44), .A3(new_n311), .ZN(new_n724));
  INV_X1    g523(.A(KEYINPUT44), .ZN(new_n725));
  INV_X1    g524(.A(new_n695), .ZN(new_n726));
  OAI21_X1  g525(.A(new_n725), .B1(new_n726), .B2(new_n312), .ZN(new_n727));
  AND2_X1   g526(.A1(new_n724), .A2(new_n727), .ZN(new_n728));
  NOR3_X1   g527(.A1(new_n249), .A2(new_n361), .A3(new_n333), .ZN(new_n729));
  NAND2_X1  g528(.A1(new_n728), .A2(new_n729), .ZN(new_n730));
  OAI21_X1  g529(.A(G29gat), .B1(new_n730), .B2(new_n636), .ZN(new_n731));
  NAND2_X1  g530(.A1(new_n723), .A2(new_n731), .ZN(G1328gat));
  NAND3_X1  g531(.A1(new_n721), .A2(new_n271), .A3(new_n617), .ZN(new_n733));
  OR2_X1    g532(.A1(new_n733), .A2(KEYINPUT46), .ZN(new_n734));
  OAI21_X1  g533(.A(G36gat), .B1(new_n730), .B2(new_n684), .ZN(new_n735));
  NAND2_X1  g534(.A1(new_n733), .A2(KEYINPUT46), .ZN(new_n736));
  NAND3_X1  g535(.A1(new_n734), .A2(new_n735), .A3(new_n736), .ZN(G1329gat));
  INV_X1    g536(.A(new_n720), .ZN(new_n738));
  AOI21_X1  g537(.A(new_n699), .B1(new_n698), .B2(new_n362), .ZN(new_n739));
  AOI211_X1 g538(.A(KEYINPUT91), .B(new_n361), .C1(new_n696), .C2(new_n697), .ZN(new_n740));
  OAI21_X1  g539(.A(new_n738), .B1(new_n739), .B2(new_n740), .ZN(new_n741));
  OAI21_X1  g540(.A(new_n266), .B1(new_n741), .B2(new_n679), .ZN(new_n742));
  NOR2_X1   g541(.A1(new_n676), .A2(new_n266), .ZN(new_n743));
  INV_X1    g542(.A(new_n743), .ZN(new_n744));
  OAI21_X1  g543(.A(new_n742), .B1(new_n730), .B2(new_n744), .ZN(new_n745));
  XNOR2_X1  g544(.A(new_n745), .B(KEYINPUT47), .ZN(G1330gat));
  INV_X1    g545(.A(new_n263), .ZN(new_n747));
  INV_X1    g546(.A(new_n608), .ZN(new_n748));
  INV_X1    g547(.A(KEYINPUT100), .ZN(new_n749));
  AOI21_X1  g548(.A(new_n748), .B1(new_n741), .B2(new_n749), .ZN(new_n750));
  NAND2_X1  g549(.A1(new_n721), .A2(KEYINPUT100), .ZN(new_n751));
  AOI21_X1  g550(.A(new_n747), .B1(new_n750), .B2(new_n751), .ZN(new_n752));
  NAND4_X1  g551(.A1(new_n728), .A2(new_n608), .A3(new_n747), .A4(new_n729), .ZN(new_n753));
  INV_X1    g552(.A(new_n753), .ZN(new_n754));
  OAI21_X1  g553(.A(KEYINPUT48), .B1(new_n752), .B2(new_n754), .ZN(new_n755));
  OAI21_X1  g554(.A(new_n608), .B1(new_n721), .B2(KEYINPUT100), .ZN(new_n756));
  NOR2_X1   g555(.A1(new_n741), .A2(new_n749), .ZN(new_n757));
  OAI21_X1  g556(.A(new_n263), .B1(new_n756), .B2(new_n757), .ZN(new_n758));
  INV_X1    g557(.A(KEYINPUT48), .ZN(new_n759));
  NAND3_X1  g558(.A1(new_n758), .A2(new_n753), .A3(new_n759), .ZN(new_n760));
  NAND2_X1  g559(.A1(new_n755), .A2(new_n760), .ZN(G1331gat));
  NAND4_X1  g560(.A1(new_n249), .A2(new_n361), .A3(new_n312), .A4(new_n333), .ZN(new_n762));
  NOR2_X1   g561(.A1(new_n726), .A2(new_n762), .ZN(new_n763));
  NAND2_X1  g562(.A1(new_n763), .A2(new_n702), .ZN(new_n764));
  XNOR2_X1  g563(.A(new_n764), .B(G57gat), .ZN(G1332gat));
  OR2_X1    g564(.A1(new_n617), .A2(KEYINPUT101), .ZN(new_n766));
  NAND2_X1  g565(.A1(new_n617), .A2(KEYINPUT101), .ZN(new_n767));
  NAND2_X1  g566(.A1(new_n766), .A2(new_n767), .ZN(new_n768));
  INV_X1    g567(.A(new_n768), .ZN(new_n769));
  AOI21_X1  g568(.A(new_n769), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n770));
  NAND2_X1  g569(.A1(new_n763), .A2(new_n770), .ZN(new_n771));
  XNOR2_X1  g570(.A(new_n771), .B(KEYINPUT102), .ZN(new_n772));
  NOR2_X1   g571(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n773));
  XNOR2_X1  g572(.A(new_n772), .B(new_n773), .ZN(G1333gat));
  INV_X1    g573(.A(new_n763), .ZN(new_n775));
  OAI21_X1  g574(.A(G71gat), .B1(new_n775), .B2(new_n676), .ZN(new_n776));
  INV_X1    g575(.A(new_n679), .ZN(new_n777));
  NAND3_X1  g576(.A1(new_n763), .A2(new_n204), .A3(new_n777), .ZN(new_n778));
  NAND2_X1  g577(.A1(new_n776), .A2(new_n778), .ZN(new_n779));
  XOR2_X1   g578(.A(new_n779), .B(KEYINPUT50), .Z(G1334gat));
  NAND2_X1  g579(.A1(new_n763), .A2(new_n608), .ZN(new_n781));
  XNOR2_X1  g580(.A(new_n781), .B(G78gat), .ZN(G1335gat));
  INV_X1    g581(.A(KEYINPUT103), .ZN(new_n783));
  NOR2_X1   g582(.A1(new_n726), .A2(new_n312), .ZN(new_n784));
  NOR2_X1   g583(.A1(new_n249), .A2(new_n362), .ZN(new_n785));
  NAND2_X1  g584(.A1(new_n784), .A2(new_n785), .ZN(new_n786));
  INV_X1    g585(.A(KEYINPUT51), .ZN(new_n787));
  OAI21_X1  g586(.A(new_n783), .B1(new_n786), .B2(new_n787), .ZN(new_n788));
  NAND4_X1  g587(.A1(new_n784), .A2(KEYINPUT103), .A3(KEYINPUT51), .A4(new_n785), .ZN(new_n789));
  AOI21_X1  g588(.A(KEYINPUT51), .B1(new_n784), .B2(new_n785), .ZN(new_n790));
  INV_X1    g589(.A(new_n790), .ZN(new_n791));
  NAND3_X1  g590(.A1(new_n788), .A2(new_n789), .A3(new_n791), .ZN(new_n792));
  NAND4_X1  g591(.A1(new_n792), .A2(new_n287), .A3(new_n702), .A4(new_n333), .ZN(new_n793));
  NOR3_X1   g592(.A1(new_n249), .A2(new_n362), .A3(new_n334), .ZN(new_n794));
  NAND3_X1  g593(.A1(new_n728), .A2(new_n702), .A3(new_n794), .ZN(new_n795));
  NAND2_X1  g594(.A1(new_n795), .A2(G85gat), .ZN(new_n796));
  NAND2_X1  g595(.A1(new_n793), .A2(new_n796), .ZN(G1336gat));
  NAND3_X1  g596(.A1(new_n768), .A2(new_n288), .A3(new_n333), .ZN(new_n798));
  XOR2_X1   g597(.A(new_n798), .B(KEYINPUT104), .Z(new_n799));
  INV_X1    g598(.A(new_n799), .ZN(new_n800));
  NAND2_X1  g599(.A1(new_n792), .A2(new_n800), .ZN(new_n801));
  INV_X1    g600(.A(KEYINPUT105), .ZN(new_n802));
  NAND4_X1  g601(.A1(new_n724), .A2(new_n727), .A3(new_n768), .A4(new_n794), .ZN(new_n803));
  AOI21_X1  g602(.A(KEYINPUT52), .B1(new_n803), .B2(G92gat), .ZN(new_n804));
  AND3_X1   g603(.A1(new_n801), .A2(new_n802), .A3(new_n804), .ZN(new_n805));
  AOI21_X1  g604(.A(new_n802), .B1(new_n801), .B2(new_n804), .ZN(new_n806));
  XNOR2_X1  g605(.A(new_n786), .B(new_n787), .ZN(new_n807));
  NAND3_X1  g606(.A1(new_n728), .A2(new_n617), .A3(new_n794), .ZN(new_n808));
  AOI22_X1  g607(.A1(new_n807), .A2(new_n800), .B1(G92gat), .B2(new_n808), .ZN(new_n809));
  INV_X1    g608(.A(KEYINPUT52), .ZN(new_n810));
  OAI22_X1  g609(.A1(new_n805), .A2(new_n806), .B1(new_n809), .B2(new_n810), .ZN(G1337gat));
  INV_X1    g610(.A(new_n676), .ZN(new_n812));
  NAND3_X1  g611(.A1(new_n728), .A2(new_n812), .A3(new_n794), .ZN(new_n813));
  NAND2_X1  g612(.A1(new_n813), .A2(G99gat), .ZN(new_n814));
  NOR3_X1   g613(.A1(new_n334), .A2(G99gat), .A3(new_n679), .ZN(new_n815));
  NAND2_X1  g614(.A1(new_n792), .A2(new_n815), .ZN(new_n816));
  NAND2_X1  g615(.A1(new_n814), .A2(new_n816), .ZN(new_n817));
  NAND2_X1  g616(.A1(new_n817), .A2(KEYINPUT106), .ZN(new_n818));
  INV_X1    g617(.A(KEYINPUT106), .ZN(new_n819));
  NAND3_X1  g618(.A1(new_n814), .A2(new_n819), .A3(new_n816), .ZN(new_n820));
  NAND2_X1  g619(.A1(new_n818), .A2(new_n820), .ZN(G1338gat));
  NAND3_X1  g620(.A1(new_n728), .A2(new_n608), .A3(new_n794), .ZN(new_n822));
  NAND2_X1  g621(.A1(new_n822), .A2(G106gat), .ZN(new_n823));
  INV_X1    g622(.A(KEYINPUT53), .ZN(new_n824));
  NAND2_X1  g623(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  NOR3_X1   g624(.A1(new_n748), .A2(new_n334), .A3(G106gat), .ZN(new_n826));
  XNOR2_X1  g625(.A(new_n826), .B(KEYINPUT107), .ZN(new_n827));
  AND2_X1   g626(.A1(new_n792), .A2(new_n827), .ZN(new_n828));
  AOI22_X1  g627(.A1(new_n822), .A2(G106gat), .B1(new_n807), .B2(new_n827), .ZN(new_n829));
  OAI22_X1  g628(.A1(new_n825), .A2(new_n828), .B1(new_n829), .B2(new_n824), .ZN(G1339gat));
  NAND4_X1  g629(.A1(new_n249), .A2(new_n361), .A3(new_n312), .A4(new_n334), .ZN(new_n831));
  INV_X1    g630(.A(KEYINPUT55), .ZN(new_n832));
  NAND3_X1  g631(.A1(new_n321), .A2(new_n325), .A3(new_n318), .ZN(new_n833));
  INV_X1    g632(.A(new_n833), .ZN(new_n834));
  INV_X1    g633(.A(KEYINPUT54), .ZN(new_n835));
  NOR3_X1   g634(.A1(new_n834), .A2(new_n326), .A3(new_n835), .ZN(new_n836));
  OAI21_X1  g635(.A(new_n316), .B1(new_n330), .B2(KEYINPUT54), .ZN(new_n837));
  OAI21_X1  g636(.A(new_n832), .B1(new_n836), .B2(new_n837), .ZN(new_n838));
  OR2_X1    g637(.A1(new_n331), .A2(new_n332), .ZN(new_n839));
  NAND3_X1  g638(.A1(new_n330), .A2(KEYINPUT54), .A3(new_n833), .ZN(new_n840));
  AOI21_X1  g639(.A(new_n315), .B1(new_n326), .B2(new_n835), .ZN(new_n841));
  NAND3_X1  g640(.A1(new_n840), .A2(KEYINPUT55), .A3(new_n841), .ZN(new_n842));
  NAND3_X1  g641(.A1(new_n838), .A2(new_n839), .A3(new_n842), .ZN(new_n843));
  AOI21_X1  g642(.A(new_n339), .B1(new_n336), .B2(new_n338), .ZN(new_n844));
  NOR3_X1   g643(.A1(new_n342), .A2(new_n343), .A3(new_n341), .ZN(new_n845));
  OAI21_X1  g644(.A(new_n348), .B1(new_n844), .B2(new_n845), .ZN(new_n846));
  NAND3_X1  g645(.A1(new_n357), .A2(new_n311), .A3(new_n846), .ZN(new_n847));
  NOR2_X1   g646(.A1(new_n843), .A2(new_n847), .ZN(new_n848));
  NAND3_X1  g647(.A1(new_n357), .A2(new_n333), .A3(new_n846), .ZN(new_n849));
  OAI21_X1  g648(.A(new_n849), .B1(new_n843), .B2(new_n361), .ZN(new_n850));
  AOI21_X1  g649(.A(new_n848), .B1(new_n850), .B2(new_n312), .ZN(new_n851));
  OAI21_X1  g650(.A(new_n831), .B1(new_n851), .B2(new_n249), .ZN(new_n852));
  AND2_X1   g651(.A1(new_n852), .A2(new_n748), .ZN(new_n853));
  NOR2_X1   g652(.A1(new_n679), .A2(new_n636), .ZN(new_n854));
  NAND2_X1  g653(.A1(new_n853), .A2(new_n854), .ZN(new_n855));
  INV_X1    g654(.A(KEYINPUT108), .ZN(new_n856));
  NAND2_X1  g655(.A1(new_n855), .A2(new_n856), .ZN(new_n857));
  NAND3_X1  g656(.A1(new_n853), .A2(KEYINPUT108), .A3(new_n854), .ZN(new_n858));
  AOI21_X1  g657(.A(new_n768), .B1(new_n857), .B2(new_n858), .ZN(new_n859));
  AND2_X1   g658(.A1(new_n859), .A2(KEYINPUT109), .ZN(new_n860));
  NOR2_X1   g659(.A1(new_n859), .A2(KEYINPUT109), .ZN(new_n861));
  OAI211_X1 g660(.A(new_n374), .B(new_n362), .C1(new_n860), .C2(new_n861), .ZN(new_n862));
  NAND3_X1  g661(.A1(new_n853), .A2(new_n769), .A3(new_n854), .ZN(new_n863));
  OAI21_X1  g662(.A(G113gat), .B1(new_n863), .B2(new_n361), .ZN(new_n864));
  NAND2_X1  g663(.A1(new_n862), .A2(new_n864), .ZN(G1340gat));
  OAI211_X1 g664(.A(new_n372), .B(new_n333), .C1(new_n860), .C2(new_n861), .ZN(new_n866));
  OAI21_X1  g665(.A(G120gat), .B1(new_n863), .B2(new_n334), .ZN(new_n867));
  NAND2_X1  g666(.A1(new_n866), .A2(new_n867), .ZN(G1341gat));
  INV_X1    g667(.A(G127gat), .ZN(new_n869));
  NAND3_X1  g668(.A1(new_n859), .A2(new_n869), .A3(new_n249), .ZN(new_n870));
  OAI21_X1  g669(.A(G127gat), .B1(new_n863), .B2(new_n719), .ZN(new_n871));
  NAND2_X1  g670(.A1(new_n870), .A2(new_n871), .ZN(G1342gat));
  NAND2_X1  g671(.A1(new_n857), .A2(new_n858), .ZN(new_n873));
  NAND2_X1  g672(.A1(new_n684), .A2(new_n311), .ZN(new_n874));
  XNOR2_X1  g673(.A(new_n874), .B(KEYINPUT110), .ZN(new_n875));
  NOR2_X1   g674(.A1(new_n875), .A2(G134gat), .ZN(new_n876));
  NAND2_X1  g675(.A1(new_n873), .A2(new_n876), .ZN(new_n877));
  OR2_X1    g676(.A1(new_n877), .A2(KEYINPUT56), .ZN(new_n878));
  OAI21_X1  g677(.A(G134gat), .B1(new_n863), .B2(new_n312), .ZN(new_n879));
  NAND2_X1  g678(.A1(new_n877), .A2(KEYINPUT56), .ZN(new_n880));
  NAND3_X1  g679(.A1(new_n878), .A2(new_n879), .A3(new_n880), .ZN(G1343gat));
  NAND2_X1  g680(.A1(new_n676), .A2(new_n702), .ZN(new_n882));
  NOR2_X1   g681(.A1(new_n768), .A2(new_n882), .ZN(new_n883));
  INV_X1    g682(.A(KEYINPUT113), .ZN(new_n884));
  NAND4_X1  g683(.A1(new_n357), .A2(new_n333), .A3(new_n884), .A4(new_n846), .ZN(new_n885));
  OAI21_X1  g684(.A(new_n885), .B1(new_n843), .B2(new_n361), .ZN(new_n886));
  NAND2_X1  g685(.A1(new_n849), .A2(KEYINPUT113), .ZN(new_n887));
  INV_X1    g686(.A(new_n887), .ZN(new_n888));
  OAI21_X1  g687(.A(new_n312), .B1(new_n886), .B2(new_n888), .ZN(new_n889));
  INV_X1    g688(.A(new_n848), .ZN(new_n890));
  AOI21_X1  g689(.A(new_n249), .B1(new_n889), .B2(new_n890), .ZN(new_n891));
  INV_X1    g690(.A(new_n831), .ZN(new_n892));
  OAI211_X1 g691(.A(KEYINPUT57), .B(new_n608), .C1(new_n891), .C2(new_n892), .ZN(new_n893));
  XNOR2_X1  g692(.A(KEYINPUT111), .B(KEYINPUT57), .ZN(new_n894));
  INV_X1    g693(.A(new_n894), .ZN(new_n895));
  AOI21_X1  g694(.A(new_n895), .B1(new_n852), .B2(new_n608), .ZN(new_n896));
  INV_X1    g695(.A(KEYINPUT112), .ZN(new_n897));
  OAI21_X1  g696(.A(new_n893), .B1(new_n896), .B2(new_n897), .ZN(new_n898));
  AOI211_X1 g697(.A(KEYINPUT112), .B(new_n895), .C1(new_n852), .C2(new_n608), .ZN(new_n899));
  OAI211_X1 g698(.A(new_n362), .B(new_n883), .C1(new_n898), .C2(new_n899), .ZN(new_n900));
  NAND2_X1  g699(.A1(new_n900), .A2(G141gat), .ZN(new_n901));
  NAND2_X1  g700(.A1(new_n901), .A2(KEYINPUT114), .ZN(new_n902));
  NAND2_X1  g701(.A1(new_n852), .A2(new_n608), .ZN(new_n903));
  NOR3_X1   g702(.A1(new_n903), .A2(new_n768), .A3(new_n882), .ZN(new_n904));
  NAND3_X1  g703(.A1(new_n904), .A2(new_n382), .A3(new_n362), .ZN(new_n905));
  NAND2_X1  g704(.A1(new_n901), .A2(new_n905), .ZN(new_n906));
  NAND3_X1  g705(.A1(new_n902), .A2(new_n906), .A3(KEYINPUT58), .ZN(new_n907));
  INV_X1    g706(.A(KEYINPUT58), .ZN(new_n908));
  OAI211_X1 g707(.A(new_n901), .B(new_n905), .C1(KEYINPUT114), .C2(new_n908), .ZN(new_n909));
  NAND2_X1  g708(.A1(new_n907), .A2(new_n909), .ZN(G1344gat));
  OAI211_X1 g709(.A(new_n333), .B(new_n883), .C1(new_n898), .C2(new_n899), .ZN(new_n911));
  NOR2_X1   g710(.A1(new_n384), .A2(KEYINPUT59), .ZN(new_n912));
  OAI211_X1 g711(.A(new_n887), .B(new_n885), .C1(new_n361), .C2(new_n843), .ZN(new_n913));
  AOI21_X1  g712(.A(new_n848), .B1(new_n913), .B2(new_n312), .ZN(new_n914));
  OAI21_X1  g713(.A(new_n831), .B1(new_n914), .B2(new_n249), .ZN(new_n915));
  AOI21_X1  g714(.A(KEYINPUT57), .B1(new_n915), .B2(new_n608), .ZN(new_n916));
  AND3_X1   g715(.A1(new_n852), .A2(new_n608), .A3(new_n895), .ZN(new_n917));
  OAI211_X1 g716(.A(new_n333), .B(new_n883), .C1(new_n916), .C2(new_n917), .ZN(new_n918));
  NAND2_X1  g717(.A1(new_n918), .A2(G148gat), .ZN(new_n919));
  AOI22_X1  g718(.A1(new_n911), .A2(new_n912), .B1(new_n919), .B2(KEYINPUT59), .ZN(new_n920));
  NAND3_X1  g719(.A1(new_n904), .A2(new_n384), .A3(new_n333), .ZN(new_n921));
  INV_X1    g720(.A(new_n921), .ZN(new_n922));
  OAI21_X1  g721(.A(KEYINPUT115), .B1(new_n920), .B2(new_n922), .ZN(new_n923));
  INV_X1    g722(.A(KEYINPUT115), .ZN(new_n924));
  AND2_X1   g723(.A1(new_n911), .A2(new_n912), .ZN(new_n925));
  INV_X1    g724(.A(KEYINPUT59), .ZN(new_n926));
  AOI21_X1  g725(.A(new_n926), .B1(new_n918), .B2(G148gat), .ZN(new_n927));
  OAI211_X1 g726(.A(new_n924), .B(new_n921), .C1(new_n925), .C2(new_n927), .ZN(new_n928));
  NAND2_X1  g727(.A1(new_n923), .A2(new_n928), .ZN(G1345gat));
  OAI21_X1  g728(.A(new_n883), .B1(new_n898), .B2(new_n899), .ZN(new_n930));
  OAI21_X1  g729(.A(G155gat), .B1(new_n930), .B2(new_n719), .ZN(new_n931));
  INV_X1    g730(.A(G155gat), .ZN(new_n932));
  NAND3_X1  g731(.A1(new_n904), .A2(new_n932), .A3(new_n249), .ZN(new_n933));
  NAND2_X1  g732(.A1(new_n931), .A2(new_n933), .ZN(G1346gat));
  OAI21_X1  g733(.A(G162gat), .B1(new_n930), .B2(new_n312), .ZN(new_n935));
  OR4_X1    g734(.A1(G162gat), .A2(new_n903), .A3(new_n875), .A4(new_n882), .ZN(new_n936));
  NAND2_X1  g735(.A1(new_n935), .A2(new_n936), .ZN(new_n937));
  INV_X1    g736(.A(KEYINPUT116), .ZN(new_n938));
  NAND2_X1  g737(.A1(new_n937), .A2(new_n938), .ZN(new_n939));
  NAND3_X1  g738(.A1(new_n935), .A2(KEYINPUT116), .A3(new_n936), .ZN(new_n940));
  NAND2_X1  g739(.A1(new_n939), .A2(new_n940), .ZN(G1347gat));
  NOR2_X1   g740(.A1(new_n684), .A2(new_n702), .ZN(new_n942));
  XNOR2_X1  g741(.A(new_n942), .B(KEYINPUT117), .ZN(new_n943));
  AND2_X1   g742(.A1(new_n943), .A2(new_n777), .ZN(new_n944));
  NAND2_X1  g743(.A1(new_n853), .A2(new_n944), .ZN(new_n945));
  NOR3_X1   g744(.A1(new_n945), .A2(new_n484), .A3(new_n361), .ZN(new_n946));
  AND2_X1   g745(.A1(new_n852), .A2(new_n636), .ZN(new_n947));
  NOR2_X1   g746(.A1(new_n769), .A2(new_n686), .ZN(new_n948));
  NAND2_X1  g747(.A1(new_n947), .A2(new_n948), .ZN(new_n949));
  INV_X1    g748(.A(new_n949), .ZN(new_n950));
  NAND2_X1  g749(.A1(new_n950), .A2(new_n362), .ZN(new_n951));
  AOI21_X1  g750(.A(new_n946), .B1(new_n484), .B2(new_n951), .ZN(G1348gat));
  OAI21_X1  g751(.A(new_n485), .B1(new_n949), .B2(new_n334), .ZN(new_n953));
  XNOR2_X1  g752(.A(new_n953), .B(KEYINPUT118), .ZN(new_n954));
  NOR3_X1   g753(.A1(new_n945), .A2(new_n485), .A3(new_n334), .ZN(new_n955));
  NOR2_X1   g754(.A1(new_n954), .A2(new_n955), .ZN(G1349gat));
  NAND3_X1  g755(.A1(new_n950), .A2(new_n469), .A3(new_n249), .ZN(new_n957));
  OAI21_X1  g756(.A(G183gat), .B1(new_n945), .B2(new_n719), .ZN(new_n958));
  NAND3_X1  g757(.A1(new_n957), .A2(KEYINPUT119), .A3(new_n958), .ZN(new_n959));
  XNOR2_X1  g758(.A(new_n959), .B(KEYINPUT60), .ZN(G1350gat));
  NOR3_X1   g759(.A1(new_n949), .A2(G190gat), .A3(new_n312), .ZN(new_n961));
  NAND3_X1  g760(.A1(new_n853), .A2(new_n311), .A3(new_n944), .ZN(new_n962));
  AND2_X1   g761(.A1(new_n962), .A2(G190gat), .ZN(new_n963));
  NOR2_X1   g762(.A1(new_n963), .A2(KEYINPUT120), .ZN(new_n964));
  INV_X1    g763(.A(KEYINPUT61), .ZN(new_n965));
  AOI21_X1  g764(.A(new_n961), .B1(new_n964), .B2(new_n965), .ZN(new_n966));
  AND2_X1   g765(.A1(new_n963), .A2(KEYINPUT120), .ZN(new_n967));
  OAI21_X1  g766(.A(KEYINPUT61), .B1(new_n963), .B2(KEYINPUT120), .ZN(new_n968));
  OAI21_X1  g767(.A(new_n966), .B1(new_n967), .B2(new_n968), .ZN(G1351gat));
  INV_X1    g768(.A(KEYINPUT124), .ZN(new_n970));
  NAND2_X1  g769(.A1(new_n943), .A2(new_n676), .ZN(new_n971));
  INV_X1    g770(.A(KEYINPUT122), .ZN(new_n972));
  XNOR2_X1  g771(.A(new_n971), .B(new_n972), .ZN(new_n973));
  INV_X1    g772(.A(KEYINPUT123), .ZN(new_n974));
  XNOR2_X1  g773(.A(new_n973), .B(new_n974), .ZN(new_n975));
  NOR2_X1   g774(.A1(new_n975), .A2(new_n361), .ZN(new_n976));
  NOR2_X1   g775(.A1(new_n916), .A2(new_n917), .ZN(new_n977));
  INV_X1    g776(.A(new_n977), .ZN(new_n978));
  AOI21_X1  g777(.A(new_n442), .B1(new_n976), .B2(new_n978), .ZN(new_n979));
  NOR3_X1   g778(.A1(new_n769), .A2(new_n748), .A3(new_n812), .ZN(new_n980));
  NAND4_X1  g779(.A1(new_n947), .A2(new_n442), .A3(new_n362), .A4(new_n980), .ZN(new_n981));
  XNOR2_X1  g780(.A(new_n981), .B(KEYINPUT121), .ZN(new_n982));
  INV_X1    g781(.A(new_n982), .ZN(new_n983));
  OAI21_X1  g782(.A(new_n970), .B1(new_n979), .B2(new_n983), .ZN(new_n984));
  XNOR2_X1  g783(.A(new_n973), .B(KEYINPUT123), .ZN(new_n985));
  NAND2_X1  g784(.A1(new_n985), .A2(new_n362), .ZN(new_n986));
  OAI21_X1  g785(.A(G197gat), .B1(new_n986), .B2(new_n977), .ZN(new_n987));
  NAND3_X1  g786(.A1(new_n987), .A2(KEYINPUT124), .A3(new_n982), .ZN(new_n988));
  NAND2_X1  g787(.A1(new_n984), .A2(new_n988), .ZN(G1352gat));
  NAND2_X1  g788(.A1(new_n947), .A2(new_n980), .ZN(new_n990));
  NOR3_X1   g789(.A1(new_n990), .A2(G204gat), .A3(new_n334), .ZN(new_n991));
  XNOR2_X1  g790(.A(KEYINPUT125), .B(KEYINPUT62), .ZN(new_n992));
  XNOR2_X1  g791(.A(new_n991), .B(new_n992), .ZN(new_n993));
  NAND3_X1  g792(.A1(new_n985), .A2(new_n978), .A3(new_n333), .ZN(new_n994));
  NAND2_X1  g793(.A1(new_n994), .A2(G204gat), .ZN(new_n995));
  NAND2_X1  g794(.A1(new_n993), .A2(new_n995), .ZN(G1353gat));
  OR3_X1    g795(.A1(new_n990), .A2(G211gat), .A3(new_n719), .ZN(new_n997));
  OAI211_X1 g796(.A(new_n249), .B(new_n973), .C1(new_n916), .C2(new_n917), .ZN(new_n998));
  AND3_X1   g797(.A1(new_n998), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n999));
  AOI21_X1  g798(.A(KEYINPUT63), .B1(new_n998), .B2(G211gat), .ZN(new_n1000));
  OAI21_X1  g799(.A(new_n997), .B1(new_n999), .B2(new_n1000), .ZN(new_n1001));
  INV_X1    g800(.A(KEYINPUT126), .ZN(new_n1002));
  NAND2_X1  g801(.A1(new_n1001), .A2(new_n1002), .ZN(new_n1003));
  OAI211_X1 g802(.A(KEYINPUT126), .B(new_n997), .C1(new_n999), .C2(new_n1000), .ZN(new_n1004));
  NAND2_X1  g803(.A1(new_n1003), .A2(new_n1004), .ZN(G1354gat));
  INV_X1    g804(.A(G218gat), .ZN(new_n1006));
  NOR2_X1   g805(.A1(new_n312), .A2(new_n1006), .ZN(new_n1007));
  NAND3_X1  g806(.A1(new_n985), .A2(new_n978), .A3(new_n1007), .ZN(new_n1008));
  OAI21_X1  g807(.A(new_n1006), .B1(new_n990), .B2(new_n312), .ZN(new_n1009));
  NAND2_X1  g808(.A1(new_n1008), .A2(new_n1009), .ZN(new_n1010));
  XNOR2_X1  g809(.A(new_n1010), .B(KEYINPUT127), .ZN(G1355gat));
endmodule


