//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 1 0 1 1 1 0 0 0 1 1 1 1 1 1 1 1 0 1 1 0 0 1 0 0 1 0 0 0 0 1 1 0 0 0 1 0 1 0 1 0 0 0 1 1 1 1 0 1 0 1 1 1 1 0 1 0 1 1 1 0 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:38:09 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n241, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n692, new_n693, new_n694, new_n695, new_n696,
    new_n697, new_n698, new_n699, new_n700, new_n701, new_n702, new_n703,
    new_n704, new_n705, new_n706, new_n707, new_n708, new_n709, new_n710,
    new_n711, new_n712, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n772, new_n773, new_n774, new_n775,
    new_n776, new_n777, new_n778, new_n779, new_n780, new_n781, new_n782,
    new_n783, new_n784, new_n785, new_n786, new_n787, new_n788, new_n789,
    new_n790, new_n791, new_n792, new_n793, new_n794, new_n795, new_n796,
    new_n797, new_n798, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n906, new_n907, new_n908, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1087,
    new_n1088, new_n1089, new_n1090, new_n1091, new_n1092, new_n1093,
    new_n1094, new_n1095, new_n1096, new_n1097, new_n1098, new_n1099,
    new_n1100, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1108, new_n1109, new_n1110, new_n1111, new_n1112,
    new_n1113, new_n1114, new_n1115, new_n1116, new_n1117, new_n1118,
    new_n1119, new_n1120, new_n1121, new_n1122, new_n1123, new_n1124,
    new_n1125, new_n1126, new_n1127, new_n1128, new_n1129, new_n1130,
    new_n1131, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1186, new_n1187, new_n1188, new_n1189, new_n1190, new_n1191,
    new_n1192, new_n1193, new_n1194, new_n1195, new_n1196, new_n1197,
    new_n1198, new_n1199, new_n1200, new_n1201, new_n1202, new_n1203,
    new_n1204, new_n1205, new_n1206, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1251, new_n1252,
    new_n1253, new_n1254, new_n1255, new_n1256, new_n1257, new_n1258,
    new_n1259, new_n1260, new_n1261, new_n1263, new_n1264, new_n1265,
    new_n1266, new_n1267, new_n1268, new_n1269, new_n1270, new_n1271,
    new_n1272, new_n1273, new_n1274, new_n1275, new_n1276, new_n1277,
    new_n1278, new_n1279, new_n1280, new_n1281, new_n1282, new_n1283,
    new_n1285, new_n1286, new_n1287, new_n1288, new_n1289, new_n1290,
    new_n1291, new_n1292, new_n1293, new_n1294, new_n1296, new_n1297,
    new_n1298, new_n1299, new_n1300, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1346,
    new_n1347, new_n1348, new_n1349, new_n1350, new_n1351, new_n1352,
    new_n1353, new_n1354, new_n1355, new_n1356, new_n1357, new_n1358,
    new_n1359, new_n1360, new_n1361, new_n1362, new_n1363, new_n1364,
    new_n1365, new_n1366, new_n1367, new_n1368, new_n1369, new_n1370,
    new_n1371, new_n1372, new_n1373, new_n1374, new_n1376, new_n1377,
    new_n1378, new_n1379, new_n1380;
  INV_X1    g0000(.A(G50), .ZN(new_n201));
  INV_X1    g0001(.A(G58), .ZN(new_n202));
  INV_X1    g0002(.A(G68), .ZN(new_n203));
  NAND3_X1  g0003(.A1(new_n201), .A2(new_n202), .A3(new_n203), .ZN(new_n204));
  NOR2_X1   g0004(.A1(new_n204), .A2(G77), .ZN(G353));
  OAI21_X1  g0005(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0006(.A1(G1), .A2(G20), .ZN(new_n207));
  AOI22_X1  g0007(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n208));
  INV_X1    g0008(.A(G232), .ZN(new_n209));
  INV_X1    g0009(.A(G97), .ZN(new_n210));
  INV_X1    g0010(.A(G257), .ZN(new_n211));
  OAI221_X1 g0011(.A(new_n208), .B1(new_n202), .B2(new_n209), .C1(new_n210), .C2(new_n211), .ZN(new_n212));
  AOI22_X1  g0012(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n213));
  AOI22_X1  g0013(.A1(G68), .A2(G238), .B1(G87), .B2(G250), .ZN(new_n214));
  NAND2_X1  g0014(.A1(new_n213), .A2(new_n214), .ZN(new_n215));
  OAI21_X1  g0015(.A(new_n207), .B1(new_n212), .B2(new_n215), .ZN(new_n216));
  XNOR2_X1  g0016(.A(new_n216), .B(KEYINPUT1), .ZN(new_n217));
  NOR2_X1   g0017(.A1(new_n207), .A2(G13), .ZN(new_n218));
  INV_X1    g0018(.A(new_n218), .ZN(new_n219));
  OAI21_X1  g0019(.A(G250), .B1(G257), .B2(G264), .ZN(new_n220));
  NOR2_X1   g0020(.A1(new_n219), .A2(new_n220), .ZN(new_n221));
  XNOR2_X1  g0021(.A(KEYINPUT64), .B(KEYINPUT0), .ZN(new_n222));
  NAND2_X1  g0022(.A1(G1), .A2(G13), .ZN(new_n223));
  INV_X1    g0023(.A(G20), .ZN(new_n224));
  NOR2_X1   g0024(.A1(new_n223), .A2(new_n224), .ZN(new_n225));
  NAND2_X1  g0025(.A1(new_n202), .A2(new_n203), .ZN(new_n226));
  NAND2_X1  g0026(.A1(new_n226), .A2(G50), .ZN(new_n227));
  INV_X1    g0027(.A(new_n227), .ZN(new_n228));
  AOI22_X1  g0028(.A1(new_n221), .A2(new_n222), .B1(new_n225), .B2(new_n228), .ZN(new_n229));
  OAI21_X1  g0029(.A(new_n229), .B1(new_n221), .B2(new_n222), .ZN(new_n230));
  NOR2_X1   g0030(.A1(new_n217), .A2(new_n230), .ZN(G361));
  XOR2_X1   g0031(.A(G238), .B(G244), .Z(new_n232));
  XNOR2_X1  g0032(.A(KEYINPUT65), .B(KEYINPUT2), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n232), .B(new_n233), .ZN(new_n234));
  XNOR2_X1  g0034(.A(G226), .B(G232), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XNOR2_X1  g0036(.A(G250), .B(G257), .ZN(new_n237));
  XNOR2_X1  g0037(.A(G264), .B(G270), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n236), .B(new_n239), .ZN(G358));
  XNOR2_X1  g0040(.A(G68), .B(G77), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n241), .B(G58), .ZN(new_n242));
  XNOR2_X1  g0042(.A(KEYINPUT66), .B(G50), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XOR2_X1   g0044(.A(G87), .B(G97), .Z(new_n245));
  XOR2_X1   g0045(.A(G107), .B(G116), .Z(new_n246));
  XNOR2_X1  g0046(.A(new_n245), .B(new_n246), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n244), .B(new_n247), .ZN(G351));
  NAND4_X1  g0048(.A1(KEYINPUT69), .A2(G1), .A3(G20), .A4(G33), .ZN(new_n249));
  NAND2_X1  g0049(.A1(new_n249), .A2(new_n223), .ZN(new_n250));
  INV_X1    g0050(.A(new_n250), .ZN(new_n251));
  NAND3_X1  g0051(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n252));
  INV_X1    g0052(.A(KEYINPUT69), .ZN(new_n253));
  NAND2_X1  g0053(.A1(new_n252), .A2(new_n253), .ZN(new_n254));
  NAND2_X1  g0054(.A1(new_n251), .A2(new_n254), .ZN(new_n255));
  INV_X1    g0055(.A(G77), .ZN(new_n256));
  INV_X1    g0056(.A(KEYINPUT70), .ZN(new_n257));
  INV_X1    g0057(.A(G33), .ZN(new_n258));
  OAI21_X1  g0058(.A(new_n257), .B1(new_n258), .B2(G20), .ZN(new_n259));
  NAND3_X1  g0059(.A1(new_n224), .A2(KEYINPUT70), .A3(G33), .ZN(new_n260));
  AOI21_X1  g0060(.A(new_n256), .B1(new_n259), .B2(new_n260), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n224), .A2(new_n258), .ZN(new_n262));
  OAI22_X1  g0062(.A1(new_n262), .A2(new_n201), .B1(new_n224), .B2(G68), .ZN(new_n263));
  OAI21_X1  g0063(.A(new_n255), .B1(new_n261), .B2(new_n263), .ZN(new_n264));
  INV_X1    g0064(.A(KEYINPUT11), .ZN(new_n265));
  OR2_X1    g0065(.A1(new_n264), .A2(new_n265), .ZN(new_n266));
  NAND2_X1  g0066(.A1(new_n264), .A2(new_n265), .ZN(new_n267));
  INV_X1    g0067(.A(G13), .ZN(new_n268));
  NOR3_X1   g0068(.A1(new_n268), .A2(new_n224), .A3(G1), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n269), .A2(new_n203), .ZN(new_n270));
  XNOR2_X1  g0070(.A(new_n270), .B(KEYINPUT12), .ZN(new_n271));
  INV_X1    g0071(.A(new_n269), .ZN(new_n272));
  NAND3_X1  g0072(.A1(new_n251), .A2(new_n272), .A3(new_n254), .ZN(new_n273));
  NOR2_X1   g0073(.A1(new_n224), .A2(G1), .ZN(new_n274));
  OR3_X1    g0074(.A1(new_n273), .A2(new_n203), .A3(new_n274), .ZN(new_n275));
  NAND4_X1  g0075(.A1(new_n266), .A2(new_n267), .A3(new_n271), .A4(new_n275), .ZN(new_n276));
  NAND2_X1  g0076(.A1(G33), .A2(G41), .ZN(new_n277));
  NAND3_X1  g0077(.A1(new_n277), .A2(G1), .A3(G13), .ZN(new_n278));
  INV_X1    g0078(.A(new_n278), .ZN(new_n279));
  NOR2_X1   g0079(.A1(G41), .A2(G45), .ZN(new_n280));
  NOR2_X1   g0080(.A1(new_n280), .A2(G1), .ZN(new_n281));
  NOR2_X1   g0081(.A1(new_n279), .A2(new_n281), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n282), .A2(G238), .ZN(new_n283));
  OAI21_X1  g0083(.A(KEYINPUT67), .B1(new_n280), .B2(G1), .ZN(new_n284));
  INV_X1    g0084(.A(KEYINPUT67), .ZN(new_n285));
  INV_X1    g0085(.A(G1), .ZN(new_n286));
  OAI211_X1 g0086(.A(new_n285), .B(new_n286), .C1(G41), .C2(G45), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n284), .A2(new_n287), .ZN(new_n288));
  INV_X1    g0088(.A(KEYINPUT68), .ZN(new_n289));
  INV_X1    g0089(.A(G274), .ZN(new_n290));
  INV_X1    g0090(.A(new_n223), .ZN(new_n291));
  AOI21_X1  g0091(.A(new_n290), .B1(new_n291), .B2(new_n277), .ZN(new_n292));
  AND3_X1   g0092(.A1(new_n288), .A2(new_n289), .A3(new_n292), .ZN(new_n293));
  AOI21_X1  g0093(.A(new_n289), .B1(new_n288), .B2(new_n292), .ZN(new_n294));
  OAI21_X1  g0094(.A(new_n283), .B1(new_n293), .B2(new_n294), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n295), .A2(KEYINPUT75), .ZN(new_n296));
  INV_X1    g0096(.A(KEYINPUT13), .ZN(new_n297));
  INV_X1    g0097(.A(KEYINPUT75), .ZN(new_n298));
  OAI211_X1 g0098(.A(new_n298), .B(new_n283), .C1(new_n293), .C2(new_n294), .ZN(new_n299));
  INV_X1    g0099(.A(KEYINPUT74), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n209), .A2(G1698), .ZN(new_n301));
  AND2_X1   g0101(.A1(KEYINPUT3), .A2(G33), .ZN(new_n302));
  NOR2_X1   g0102(.A1(KEYINPUT3), .A2(G33), .ZN(new_n303));
  OAI221_X1 g0103(.A(new_n301), .B1(G226), .B2(G1698), .C1(new_n302), .C2(new_n303), .ZN(new_n304));
  INV_X1    g0104(.A(new_n304), .ZN(new_n305));
  NOR2_X1   g0105(.A1(new_n258), .A2(new_n210), .ZN(new_n306));
  OAI211_X1 g0106(.A(new_n300), .B(new_n279), .C1(new_n305), .C2(new_n306), .ZN(new_n307));
  NOR2_X1   g0107(.A1(G226), .A2(G1698), .ZN(new_n308));
  AOI21_X1  g0108(.A(new_n308), .B1(new_n209), .B2(G1698), .ZN(new_n309));
  XNOR2_X1  g0109(.A(KEYINPUT3), .B(G33), .ZN(new_n310));
  AOI21_X1  g0110(.A(new_n306), .B1(new_n309), .B2(new_n310), .ZN(new_n311));
  OAI21_X1  g0111(.A(KEYINPUT74), .B1(new_n311), .B2(new_n278), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n307), .A2(new_n312), .ZN(new_n313));
  NAND4_X1  g0113(.A1(new_n296), .A2(new_n297), .A3(new_n299), .A4(new_n313), .ZN(new_n314));
  INV_X1    g0114(.A(KEYINPUT76), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n314), .A2(new_n315), .ZN(new_n316));
  AND2_X1   g0116(.A1(new_n313), .A2(new_n299), .ZN(new_n317));
  NAND4_X1  g0117(.A1(new_n317), .A2(KEYINPUT76), .A3(new_n297), .A4(new_n296), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n313), .A2(new_n299), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n288), .A2(new_n292), .ZN(new_n320));
  NAND2_X1  g0120(.A1(new_n320), .A2(KEYINPUT68), .ZN(new_n321));
  NAND3_X1  g0121(.A1(new_n288), .A2(new_n289), .A3(new_n292), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n321), .A2(new_n322), .ZN(new_n323));
  AOI21_X1  g0123(.A(new_n298), .B1(new_n323), .B2(new_n283), .ZN(new_n324));
  OAI21_X1  g0124(.A(KEYINPUT13), .B1(new_n319), .B2(new_n324), .ZN(new_n325));
  NAND3_X1  g0125(.A1(new_n316), .A2(new_n318), .A3(new_n325), .ZN(new_n326));
  AOI21_X1  g0126(.A(new_n276), .B1(new_n326), .B2(G200), .ZN(new_n327));
  INV_X1    g0127(.A(KEYINPUT77), .ZN(new_n328));
  OAI21_X1  g0128(.A(new_n328), .B1(new_n319), .B2(new_n324), .ZN(new_n329));
  NAND4_X1  g0129(.A1(new_n296), .A2(KEYINPUT77), .A3(new_n299), .A4(new_n313), .ZN(new_n330));
  NAND3_X1  g0130(.A1(new_n329), .A2(KEYINPUT13), .A3(new_n330), .ZN(new_n331));
  AND2_X1   g0131(.A1(new_n314), .A2(G190), .ZN(new_n332));
  INV_X1    g0132(.A(KEYINPUT78), .ZN(new_n333));
  AND3_X1   g0133(.A1(new_n331), .A2(new_n332), .A3(new_n333), .ZN(new_n334));
  AOI21_X1  g0134(.A(new_n333), .B1(new_n331), .B2(new_n332), .ZN(new_n335));
  OAI21_X1  g0135(.A(new_n327), .B1(new_n334), .B2(new_n335), .ZN(new_n336));
  INV_X1    g0136(.A(KEYINPUT14), .ZN(new_n337));
  AND3_X1   g0137(.A1(new_n326), .A2(new_n337), .A3(G169), .ZN(new_n338));
  AOI21_X1  g0138(.A(new_n337), .B1(new_n326), .B2(G169), .ZN(new_n339));
  NAND3_X1  g0139(.A1(new_n331), .A2(G179), .A3(new_n314), .ZN(new_n340));
  INV_X1    g0140(.A(new_n340), .ZN(new_n341));
  NOR3_X1   g0141(.A1(new_n338), .A2(new_n339), .A3(new_n341), .ZN(new_n342));
  INV_X1    g0142(.A(new_n276), .ZN(new_n343));
  OAI21_X1  g0143(.A(new_n336), .B1(new_n342), .B2(new_n343), .ZN(new_n344));
  AOI22_X1  g0144(.A1(new_n321), .A2(new_n322), .B1(G232), .B2(new_n282), .ZN(new_n345));
  INV_X1    g0145(.A(KEYINPUT82), .ZN(new_n346));
  OR2_X1    g0146(.A1(G223), .A2(G1698), .ZN(new_n347));
  INV_X1    g0147(.A(G226), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n348), .A2(G1698), .ZN(new_n349));
  OAI211_X1 g0149(.A(new_n347), .B(new_n349), .C1(new_n302), .C2(new_n303), .ZN(new_n350));
  NAND2_X1  g0150(.A1(G33), .A2(G87), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n350), .A2(new_n351), .ZN(new_n352));
  AOI21_X1  g0152(.A(new_n346), .B1(new_n352), .B2(new_n279), .ZN(new_n353));
  AOI211_X1 g0153(.A(KEYINPUT82), .B(new_n278), .C1(new_n350), .C2(new_n351), .ZN(new_n354));
  NOR2_X1   g0154(.A1(new_n353), .A2(new_n354), .ZN(new_n355));
  INV_X1    g0155(.A(G179), .ZN(new_n356));
  NAND3_X1  g0156(.A1(new_n345), .A2(new_n355), .A3(new_n356), .ZN(new_n357));
  INV_X1    g0157(.A(KEYINPUT83), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n357), .A2(new_n358), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n282), .A2(G232), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n352), .A2(new_n279), .ZN(new_n361));
  OAI211_X1 g0161(.A(new_n360), .B(new_n361), .C1(new_n293), .C2(new_n294), .ZN(new_n362));
  INV_X1    g0162(.A(G169), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n362), .A2(new_n363), .ZN(new_n364));
  NAND4_X1  g0164(.A1(new_n345), .A2(new_n355), .A3(KEYINPUT83), .A4(new_n356), .ZN(new_n365));
  AND3_X1   g0165(.A1(new_n359), .A2(new_n364), .A3(new_n365), .ZN(new_n366));
  INV_X1    g0166(.A(new_n273), .ZN(new_n367));
  XOR2_X1   g0167(.A(KEYINPUT8), .B(G58), .Z(new_n368));
  INV_X1    g0168(.A(new_n368), .ZN(new_n369));
  NOR2_X1   g0169(.A1(new_n369), .A2(new_n274), .ZN(new_n370));
  AOI22_X1  g0170(.A1(new_n367), .A2(new_n370), .B1(new_n269), .B2(new_n369), .ZN(new_n371));
  INV_X1    g0171(.A(KEYINPUT81), .ZN(new_n372));
  NOR2_X1   g0172(.A1(new_n302), .A2(new_n303), .ZN(new_n373));
  AOI21_X1  g0173(.A(KEYINPUT7), .B1(new_n373), .B2(new_n224), .ZN(new_n374));
  INV_X1    g0174(.A(KEYINPUT7), .ZN(new_n375));
  NOR4_X1   g0175(.A1(new_n302), .A2(new_n303), .A3(new_n375), .A4(G20), .ZN(new_n376));
  OAI21_X1  g0176(.A(G68), .B1(new_n374), .B2(new_n376), .ZN(new_n377));
  NAND2_X1  g0177(.A1(G58), .A2(G68), .ZN(new_n378));
  INV_X1    g0178(.A(KEYINPUT79), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n378), .A2(new_n379), .ZN(new_n380));
  NAND3_X1  g0180(.A1(KEYINPUT79), .A2(G58), .A3(G68), .ZN(new_n381));
  NAND3_X1  g0181(.A1(new_n380), .A2(new_n226), .A3(new_n381), .ZN(new_n382));
  INV_X1    g0182(.A(G159), .ZN(new_n383));
  OAI21_X1  g0183(.A(KEYINPUT80), .B1(new_n262), .B2(new_n383), .ZN(new_n384));
  NOR2_X1   g0184(.A1(G20), .A2(G33), .ZN(new_n385));
  INV_X1    g0185(.A(KEYINPUT80), .ZN(new_n386));
  NAND3_X1  g0186(.A1(new_n385), .A2(new_n386), .A3(G159), .ZN(new_n387));
  AOI22_X1  g0187(.A1(new_n382), .A2(G20), .B1(new_n384), .B2(new_n387), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n377), .A2(new_n388), .ZN(new_n389));
  INV_X1    g0189(.A(KEYINPUT16), .ZN(new_n390));
  AOI22_X1  g0190(.A1(new_n389), .A2(new_n390), .B1(new_n254), .B2(new_n251), .ZN(new_n391));
  NAND3_X1  g0191(.A1(new_n377), .A2(KEYINPUT16), .A3(new_n388), .ZN(new_n392));
  AOI21_X1  g0192(.A(new_n372), .B1(new_n391), .B2(new_n392), .ZN(new_n393));
  OAI21_X1  g0193(.A(new_n375), .B1(new_n310), .B2(G20), .ZN(new_n394));
  NAND3_X1  g0194(.A1(new_n373), .A2(KEYINPUT7), .A3(new_n224), .ZN(new_n395));
  AOI21_X1  g0195(.A(new_n203), .B1(new_n394), .B2(new_n395), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n382), .A2(G20), .ZN(new_n397));
  NAND2_X1  g0197(.A1(new_n384), .A2(new_n387), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n397), .A2(new_n398), .ZN(new_n399));
  OAI21_X1  g0199(.A(new_n390), .B1(new_n396), .B2(new_n399), .ZN(new_n400));
  AND4_X1   g0200(.A1(new_n372), .A2(new_n400), .A3(new_n392), .A4(new_n255), .ZN(new_n401));
  OAI21_X1  g0201(.A(new_n371), .B1(new_n393), .B2(new_n401), .ZN(new_n402));
  INV_X1    g0202(.A(KEYINPUT18), .ZN(new_n403));
  NAND3_X1  g0203(.A1(new_n366), .A2(new_n402), .A3(new_n403), .ZN(new_n404));
  INV_X1    g0204(.A(new_n371), .ZN(new_n405));
  NAND3_X1  g0205(.A1(new_n391), .A2(new_n372), .A3(new_n392), .ZN(new_n406));
  NAND3_X1  g0206(.A1(new_n400), .A2(new_n392), .A3(new_n255), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n407), .A2(KEYINPUT81), .ZN(new_n408));
  AOI21_X1  g0208(.A(new_n405), .B1(new_n406), .B2(new_n408), .ZN(new_n409));
  NAND3_X1  g0209(.A1(new_n359), .A2(new_n364), .A3(new_n365), .ZN(new_n410));
  OAI21_X1  g0210(.A(KEYINPUT18), .B1(new_n409), .B2(new_n410), .ZN(new_n411));
  INV_X1    g0211(.A(G190), .ZN(new_n412));
  NAND3_X1  g0212(.A1(new_n345), .A2(new_n355), .A3(new_n412), .ZN(new_n413));
  INV_X1    g0213(.A(G200), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n362), .A2(new_n414), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n413), .A2(new_n415), .ZN(new_n416));
  OAI211_X1 g0216(.A(new_n416), .B(new_n371), .C1(new_n393), .C2(new_n401), .ZN(new_n417));
  INV_X1    g0217(.A(KEYINPUT17), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n417), .A2(new_n418), .ZN(new_n419));
  NAND3_X1  g0219(.A1(new_n409), .A2(KEYINPUT17), .A3(new_n416), .ZN(new_n420));
  NAND4_X1  g0220(.A1(new_n404), .A2(new_n411), .A3(new_n419), .A4(new_n420), .ZN(new_n421));
  NOR3_X1   g0221(.A1(new_n273), .A2(new_n201), .A3(new_n274), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n259), .A2(new_n260), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n368), .A2(new_n423), .ZN(new_n424));
  AOI22_X1  g0224(.A1(new_n204), .A2(G20), .B1(G150), .B2(new_n385), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n424), .A2(new_n425), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n426), .A2(new_n255), .ZN(new_n427));
  AOI21_X1  g0227(.A(new_n422), .B1(KEYINPUT71), .B2(new_n427), .ZN(new_n428));
  OR2_X1    g0228(.A1(new_n427), .A2(KEYINPUT71), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n269), .A2(new_n201), .ZN(new_n430));
  NAND3_X1  g0230(.A1(new_n428), .A2(new_n429), .A3(new_n430), .ZN(new_n431));
  INV_X1    g0231(.A(KEYINPUT9), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n431), .A2(new_n432), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n282), .A2(G226), .ZN(new_n434));
  INV_X1    g0234(.A(G1698), .ZN(new_n435));
  OR2_X1    g0235(.A1(KEYINPUT3), .A2(G33), .ZN(new_n436));
  NAND2_X1  g0236(.A1(KEYINPUT3), .A2(G33), .ZN(new_n437));
  AOI21_X1  g0237(.A(new_n435), .B1(new_n436), .B2(new_n437), .ZN(new_n438));
  AOI22_X1  g0238(.A1(new_n438), .A2(G223), .B1(new_n373), .B2(G77), .ZN(new_n439));
  NAND3_X1  g0239(.A1(new_n310), .A2(G222), .A3(new_n435), .ZN(new_n440));
  AND2_X1   g0240(.A1(new_n439), .A2(new_n440), .ZN(new_n441));
  OAI211_X1 g0241(.A(new_n323), .B(new_n434), .C1(new_n441), .C2(new_n278), .ZN(new_n442));
  OR2_X1    g0242(.A1(new_n442), .A2(new_n412), .ZN(new_n443));
  NAND4_X1  g0243(.A1(new_n428), .A2(new_n429), .A3(KEYINPUT9), .A4(new_n430), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n442), .A2(G200), .ZN(new_n445));
  NAND4_X1  g0245(.A1(new_n433), .A2(new_n443), .A3(new_n444), .A4(new_n445), .ZN(new_n446));
  XNOR2_X1  g0246(.A(new_n446), .B(KEYINPUT10), .ZN(new_n447));
  NAND2_X1  g0247(.A1(new_n442), .A2(new_n363), .ZN(new_n448));
  OAI211_X1 g0248(.A(new_n431), .B(new_n448), .C1(G179), .C2(new_n442), .ZN(new_n449));
  XOR2_X1   g0249(.A(new_n449), .B(KEYINPUT72), .Z(new_n450));
  NAND2_X1  g0250(.A1(new_n282), .A2(G244), .ZN(new_n451));
  AOI22_X1  g0251(.A1(new_n438), .A2(G238), .B1(new_n373), .B2(G107), .ZN(new_n452));
  NAND3_X1  g0252(.A1(new_n310), .A2(G232), .A3(new_n435), .ZN(new_n453));
  AND2_X1   g0253(.A1(new_n452), .A2(new_n453), .ZN(new_n454));
  OAI211_X1 g0254(.A(new_n323), .B(new_n451), .C1(new_n454), .C2(new_n278), .ZN(new_n455));
  OR2_X1    g0255(.A1(new_n455), .A2(G179), .ZN(new_n456));
  XNOR2_X1  g0256(.A(KEYINPUT15), .B(G87), .ZN(new_n457));
  INV_X1    g0257(.A(new_n457), .ZN(new_n458));
  AOI22_X1  g0258(.A1(new_n458), .A2(new_n423), .B1(G20), .B2(G77), .ZN(new_n459));
  AND2_X1   g0259(.A1(new_n385), .A2(KEYINPUT73), .ZN(new_n460));
  OAI21_X1  g0260(.A(new_n368), .B1(KEYINPUT73), .B2(new_n385), .ZN(new_n461));
  OAI21_X1  g0261(.A(new_n459), .B1(new_n460), .B2(new_n461), .ZN(new_n462));
  AND2_X1   g0262(.A1(new_n462), .A2(new_n255), .ZN(new_n463));
  NOR3_X1   g0263(.A1(new_n273), .A2(new_n256), .A3(new_n274), .ZN(new_n464));
  NOR2_X1   g0264(.A1(new_n272), .A2(G77), .ZN(new_n465));
  OR3_X1    g0265(.A1(new_n463), .A2(new_n464), .A3(new_n465), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n455), .A2(new_n363), .ZN(new_n467));
  NAND3_X1  g0267(.A1(new_n456), .A2(new_n466), .A3(new_n467), .ZN(new_n468));
  NOR3_X1   g0268(.A1(new_n463), .A2(new_n464), .A3(new_n465), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n455), .A2(G200), .ZN(new_n470));
  OAI211_X1 g0270(.A(new_n469), .B(new_n470), .C1(new_n412), .C2(new_n455), .ZN(new_n471));
  AND2_X1   g0271(.A1(new_n468), .A2(new_n471), .ZN(new_n472));
  NAND3_X1  g0272(.A1(new_n447), .A2(new_n450), .A3(new_n472), .ZN(new_n473));
  NOR3_X1   g0273(.A1(new_n344), .A2(new_n421), .A3(new_n473), .ZN(new_n474));
  INV_X1    g0274(.A(new_n474), .ZN(new_n475));
  OAI211_X1 g0275(.A(G257), .B(G1698), .C1(new_n302), .C2(new_n303), .ZN(new_n476));
  OAI211_X1 g0276(.A(G250), .B(new_n435), .C1(new_n302), .C2(new_n303), .ZN(new_n477));
  NAND2_X1  g0277(.A1(G33), .A2(G294), .ZN(new_n478));
  NAND3_X1  g0278(.A1(new_n476), .A2(new_n477), .A3(new_n478), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n479), .A2(KEYINPUT94), .ZN(new_n480));
  INV_X1    g0280(.A(KEYINPUT94), .ZN(new_n481));
  NAND4_X1  g0281(.A1(new_n476), .A2(new_n477), .A3(new_n481), .A4(new_n478), .ZN(new_n482));
  NAND3_X1  g0282(.A1(new_n480), .A2(new_n279), .A3(new_n482), .ZN(new_n483));
  INV_X1    g0283(.A(G45), .ZN(new_n484));
  NOR2_X1   g0284(.A1(new_n484), .A2(G1), .ZN(new_n485));
  NOR2_X1   g0285(.A1(KEYINPUT5), .A2(G41), .ZN(new_n486));
  AND2_X1   g0286(.A1(KEYINPUT5), .A2(G41), .ZN(new_n487));
  OAI211_X1 g0287(.A(new_n292), .B(new_n485), .C1(new_n486), .C2(new_n487), .ZN(new_n488));
  OAI21_X1  g0288(.A(new_n485), .B1(new_n487), .B2(new_n486), .ZN(new_n489));
  AND3_X1   g0289(.A1(new_n489), .A2(G264), .A3(new_n278), .ZN(new_n490));
  INV_X1    g0290(.A(new_n490), .ZN(new_n491));
  NAND4_X1  g0291(.A1(new_n483), .A2(new_n412), .A3(new_n488), .A4(new_n491), .ZN(new_n492));
  NOR3_X1   g0292(.A1(new_n489), .A2(new_n279), .A3(new_n290), .ZN(new_n493));
  AOI21_X1  g0293(.A(new_n278), .B1(new_n479), .B2(KEYINPUT94), .ZN(new_n494));
  AOI211_X1 g0294(.A(new_n493), .B(new_n490), .C1(new_n494), .C2(new_n482), .ZN(new_n495));
  OAI21_X1  g0295(.A(new_n492), .B1(new_n495), .B2(G200), .ZN(new_n496));
  INV_X1    g0296(.A(G107), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n269), .A2(new_n497), .ZN(new_n498));
  XOR2_X1   g0298(.A(new_n498), .B(KEYINPUT25), .Z(new_n499));
  NAND2_X1  g0299(.A1(new_n286), .A2(G33), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n367), .A2(new_n500), .ZN(new_n501));
  OAI21_X1  g0301(.A(new_n499), .B1(new_n501), .B2(new_n497), .ZN(new_n502));
  OAI211_X1 g0302(.A(new_n224), .B(G87), .C1(new_n302), .C2(new_n303), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n503), .A2(KEYINPUT22), .ZN(new_n504));
  INV_X1    g0304(.A(KEYINPUT22), .ZN(new_n505));
  NAND4_X1  g0305(.A1(new_n310), .A2(new_n505), .A3(new_n224), .A4(G87), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n504), .A2(new_n506), .ZN(new_n507));
  INV_X1    g0307(.A(G116), .ZN(new_n508));
  NOR3_X1   g0308(.A1(new_n258), .A2(new_n508), .A3(G20), .ZN(new_n509));
  INV_X1    g0309(.A(KEYINPUT93), .ZN(new_n510));
  OAI21_X1  g0310(.A(new_n510), .B1(new_n224), .B2(G107), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n511), .A2(KEYINPUT23), .ZN(new_n512));
  INV_X1    g0312(.A(KEYINPUT23), .ZN(new_n513));
  OAI211_X1 g0313(.A(new_n510), .B(new_n513), .C1(new_n224), .C2(G107), .ZN(new_n514));
  AOI21_X1  g0314(.A(new_n509), .B1(new_n512), .B2(new_n514), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n507), .A2(new_n515), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n516), .A2(KEYINPUT24), .ZN(new_n517));
  INV_X1    g0317(.A(KEYINPUT24), .ZN(new_n518));
  NAND3_X1  g0318(.A1(new_n507), .A2(new_n518), .A3(new_n515), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n517), .A2(new_n519), .ZN(new_n520));
  AOI21_X1  g0320(.A(new_n502), .B1(new_n520), .B2(new_n255), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n496), .A2(new_n521), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n522), .A2(KEYINPUT95), .ZN(new_n523));
  INV_X1    g0323(.A(KEYINPUT95), .ZN(new_n524));
  NAND3_X1  g0324(.A1(new_n496), .A2(new_n521), .A3(new_n524), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n523), .A2(new_n525), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n489), .A2(new_n278), .ZN(new_n527));
  OAI21_X1  g0327(.A(new_n488), .B1(new_n211), .B2(new_n527), .ZN(new_n528));
  INV_X1    g0328(.A(new_n528), .ZN(new_n529));
  OAI211_X1 g0329(.A(G244), .B(new_n435), .C1(new_n302), .C2(new_n303), .ZN(new_n530));
  INV_X1    g0330(.A(KEYINPUT4), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n530), .A2(new_n531), .ZN(new_n532));
  INV_X1    g0332(.A(KEYINPUT84), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  OR2_X1    g0334(.A1(new_n530), .A2(new_n531), .ZN(new_n535));
  NAND3_X1  g0335(.A1(new_n530), .A2(KEYINPUT84), .A3(new_n531), .ZN(new_n536));
  OAI211_X1 g0336(.A(G250), .B(G1698), .C1(new_n302), .C2(new_n303), .ZN(new_n537));
  NAND2_X1  g0337(.A1(G33), .A2(G283), .ZN(new_n538));
  AND2_X1   g0338(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  NAND4_X1  g0339(.A1(new_n534), .A2(new_n535), .A3(new_n536), .A4(new_n539), .ZN(new_n540));
  AND3_X1   g0340(.A1(new_n540), .A2(KEYINPUT85), .A3(new_n279), .ZN(new_n541));
  AOI21_X1  g0341(.A(KEYINPUT85), .B1(new_n540), .B2(new_n279), .ZN(new_n542));
  OAI211_X1 g0342(.A(new_n356), .B(new_n529), .C1(new_n541), .C2(new_n542), .ZN(new_n543));
  INV_X1    g0343(.A(new_n536), .ZN(new_n544));
  OAI211_X1 g0344(.A(new_n538), .B(new_n537), .C1(new_n530), .C2(new_n531), .ZN(new_n545));
  AOI21_X1  g0345(.A(KEYINPUT84), .B1(new_n530), .B2(new_n531), .ZN(new_n546));
  NOR3_X1   g0346(.A1(new_n544), .A2(new_n545), .A3(new_n546), .ZN(new_n547));
  OAI21_X1  g0347(.A(new_n529), .B1(new_n547), .B2(new_n278), .ZN(new_n548));
  NOR2_X1   g0348(.A1(new_n272), .A2(G97), .ZN(new_n549));
  OAI21_X1  g0349(.A(G107), .B1(new_n374), .B2(new_n376), .ZN(new_n550));
  INV_X1    g0350(.A(KEYINPUT6), .ZN(new_n551));
  AND2_X1   g0351(.A1(G97), .A2(G107), .ZN(new_n552));
  NOR2_X1   g0352(.A1(G97), .A2(G107), .ZN(new_n553));
  OAI21_X1  g0353(.A(new_n551), .B1(new_n552), .B2(new_n553), .ZN(new_n554));
  NAND3_X1  g0354(.A1(new_n497), .A2(KEYINPUT6), .A3(G97), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  AOI22_X1  g0356(.A1(new_n556), .A2(G20), .B1(G77), .B2(new_n385), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n550), .A2(new_n557), .ZN(new_n558));
  AOI21_X1  g0358(.A(new_n549), .B1(new_n558), .B2(new_n255), .ZN(new_n559));
  NAND3_X1  g0359(.A1(new_n367), .A2(G97), .A3(new_n500), .ZN(new_n560));
  AOI22_X1  g0360(.A1(new_n548), .A2(new_n363), .B1(new_n559), .B2(new_n560), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n543), .A2(new_n561), .ZN(new_n562));
  XNOR2_X1  g0362(.A(G97), .B(G107), .ZN(new_n563));
  NOR2_X1   g0363(.A1(new_n551), .A2(new_n210), .ZN(new_n564));
  AOI22_X1  g0364(.A1(new_n563), .A2(new_n551), .B1(new_n497), .B2(new_n564), .ZN(new_n565));
  OAI22_X1  g0365(.A1(new_n565), .A2(new_n224), .B1(new_n256), .B2(new_n262), .ZN(new_n566));
  AOI21_X1  g0366(.A(new_n497), .B1(new_n394), .B2(new_n395), .ZN(new_n567));
  OAI21_X1  g0367(.A(new_n255), .B1(new_n566), .B2(new_n567), .ZN(new_n568));
  INV_X1    g0368(.A(new_n549), .ZN(new_n569));
  NAND3_X1  g0369(.A1(new_n568), .A2(new_n560), .A3(new_n569), .ZN(new_n570));
  AOI21_X1  g0370(.A(new_n528), .B1(new_n540), .B2(new_n279), .ZN(new_n571));
  AOI21_X1  g0371(.A(new_n570), .B1(G190), .B2(new_n571), .ZN(new_n572));
  INV_X1    g0372(.A(KEYINPUT85), .ZN(new_n573));
  OAI21_X1  g0373(.A(new_n573), .B1(new_n547), .B2(new_n278), .ZN(new_n574));
  NAND3_X1  g0374(.A1(new_n540), .A2(KEYINPUT85), .A3(new_n279), .ZN(new_n575));
  AOI21_X1  g0375(.A(new_n528), .B1(new_n574), .B2(new_n575), .ZN(new_n576));
  OAI211_X1 g0376(.A(new_n572), .B(KEYINPUT86), .C1(new_n576), .C2(new_n414), .ZN(new_n577));
  INV_X1    g0377(.A(new_n577), .ZN(new_n578));
  OAI21_X1  g0378(.A(new_n529), .B1(new_n541), .B2(new_n542), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n579), .A2(G200), .ZN(new_n580));
  AOI21_X1  g0380(.A(KEYINPUT86), .B1(new_n580), .B2(new_n572), .ZN(new_n581));
  OAI211_X1 g0381(.A(new_n526), .B(new_n562), .C1(new_n578), .C2(new_n581), .ZN(new_n582));
  NAND3_X1  g0382(.A1(new_n489), .A2(G270), .A3(new_n278), .ZN(new_n583));
  INV_X1    g0383(.A(KEYINPUT89), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  NAND4_X1  g0385(.A1(new_n489), .A2(KEYINPUT89), .A3(G270), .A4(new_n278), .ZN(new_n586));
  AOI21_X1  g0386(.A(new_n493), .B1(new_n585), .B2(new_n586), .ZN(new_n587));
  OAI211_X1 g0387(.A(G264), .B(G1698), .C1(new_n302), .C2(new_n303), .ZN(new_n588));
  INV_X1    g0388(.A(KEYINPUT90), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n588), .A2(new_n589), .ZN(new_n590));
  NAND4_X1  g0390(.A1(new_n310), .A2(KEYINPUT90), .A3(G264), .A4(G1698), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n373), .A2(G303), .ZN(new_n592));
  NAND3_X1  g0392(.A1(new_n310), .A2(G257), .A3(new_n435), .ZN(new_n593));
  NAND4_X1  g0393(.A1(new_n590), .A2(new_n591), .A3(new_n592), .A4(new_n593), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n594), .A2(new_n279), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n587), .A2(new_n595), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n596), .A2(KEYINPUT91), .ZN(new_n597));
  INV_X1    g0397(.A(KEYINPUT91), .ZN(new_n598));
  NAND3_X1  g0398(.A1(new_n587), .A2(new_n595), .A3(new_n598), .ZN(new_n599));
  NAND4_X1  g0399(.A1(new_n597), .A2(KEYINPUT21), .A3(G169), .A4(new_n599), .ZN(new_n600));
  NAND3_X1  g0400(.A1(new_n587), .A2(new_n595), .A3(G179), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  NOR2_X1   g0402(.A1(new_n272), .A2(G116), .ZN(new_n603));
  AOI21_X1  g0403(.A(new_n273), .B1(new_n286), .B2(G33), .ZN(new_n604));
  AOI21_X1  g0404(.A(new_n603), .B1(new_n604), .B2(G116), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n508), .A2(G20), .ZN(new_n606));
  AND2_X1   g0406(.A1(new_n252), .A2(new_n253), .ZN(new_n607));
  OAI21_X1  g0407(.A(new_n606), .B1(new_n607), .B2(new_n250), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n608), .A2(KEYINPUT92), .ZN(new_n609));
  INV_X1    g0409(.A(KEYINPUT92), .ZN(new_n610));
  OAI211_X1 g0410(.A(new_n610), .B(new_n606), .C1(new_n607), .C2(new_n250), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n609), .A2(new_n611), .ZN(new_n612));
  OAI211_X1 g0412(.A(new_n538), .B(new_n224), .C1(G33), .C2(new_n210), .ZN(new_n613));
  AOI21_X1  g0413(.A(KEYINPUT20), .B1(new_n612), .B2(new_n613), .ZN(new_n614));
  INV_X1    g0414(.A(KEYINPUT20), .ZN(new_n615));
  INV_X1    g0415(.A(new_n613), .ZN(new_n616));
  AOI211_X1 g0416(.A(new_n615), .B(new_n616), .C1(new_n609), .C2(new_n611), .ZN(new_n617));
  OAI21_X1  g0417(.A(new_n605), .B1(new_n614), .B2(new_n617), .ZN(new_n618));
  NAND4_X1  g0418(.A1(new_n618), .A2(G169), .A3(new_n597), .A4(new_n599), .ZN(new_n619));
  INV_X1    g0419(.A(KEYINPUT21), .ZN(new_n620));
  AOI22_X1  g0420(.A1(new_n602), .A2(new_n618), .B1(new_n619), .B2(new_n620), .ZN(new_n621));
  OAI211_X1 g0421(.A(new_n224), .B(G68), .C1(new_n302), .C2(new_n303), .ZN(new_n622));
  AOI21_X1  g0422(.A(new_n210), .B1(new_n259), .B2(new_n260), .ZN(new_n623));
  OAI21_X1  g0423(.A(new_n622), .B1(new_n623), .B2(KEYINPUT19), .ZN(new_n624));
  NAND3_X1  g0424(.A1(KEYINPUT19), .A2(G33), .A3(G97), .ZN(new_n625));
  AND3_X1   g0425(.A1(new_n625), .A2(KEYINPUT87), .A3(new_n224), .ZN(new_n626));
  AOI21_X1  g0426(.A(KEYINPUT87), .B1(new_n625), .B2(new_n224), .ZN(new_n627));
  NOR3_X1   g0427(.A1(G87), .A2(G97), .A3(G107), .ZN(new_n628));
  NOR3_X1   g0428(.A1(new_n626), .A2(new_n627), .A3(new_n628), .ZN(new_n629));
  OAI21_X1  g0429(.A(new_n255), .B1(new_n624), .B2(new_n629), .ZN(new_n630));
  INV_X1    g0430(.A(KEYINPUT88), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n457), .A2(new_n269), .ZN(new_n632));
  AND3_X1   g0432(.A1(new_n630), .A2(new_n631), .A3(new_n632), .ZN(new_n633));
  AOI21_X1  g0433(.A(new_n631), .B1(new_n630), .B2(new_n632), .ZN(new_n634));
  OAI22_X1  g0434(.A1(new_n633), .A2(new_n634), .B1(new_n457), .B2(new_n501), .ZN(new_n635));
  OAI211_X1 g0435(.A(new_n278), .B(G250), .C1(G1), .C2(new_n484), .ZN(new_n636));
  NAND3_X1  g0436(.A1(new_n278), .A2(G274), .A3(new_n485), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  NAND3_X1  g0438(.A1(new_n310), .A2(G244), .A3(G1698), .ZN(new_n639));
  NAND3_X1  g0439(.A1(new_n310), .A2(G238), .A3(new_n435), .ZN(new_n640));
  NAND2_X1  g0440(.A1(G33), .A2(G116), .ZN(new_n641));
  NAND3_X1  g0441(.A1(new_n639), .A2(new_n640), .A3(new_n641), .ZN(new_n642));
  AOI21_X1  g0442(.A(new_n638), .B1(new_n642), .B2(new_n279), .ZN(new_n643));
  NOR2_X1   g0443(.A1(new_n643), .A2(G169), .ZN(new_n644));
  AOI21_X1  g0444(.A(new_n644), .B1(new_n356), .B2(new_n643), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n635), .A2(new_n645), .ZN(new_n646));
  AND3_X1   g0446(.A1(new_n507), .A2(new_n518), .A3(new_n515), .ZN(new_n647));
  AOI21_X1  g0447(.A(new_n518), .B1(new_n507), .B2(new_n515), .ZN(new_n648));
  OAI21_X1  g0448(.A(new_n255), .B1(new_n647), .B2(new_n648), .ZN(new_n649));
  XNOR2_X1  g0449(.A(new_n498), .B(KEYINPUT25), .ZN(new_n650));
  AOI21_X1  g0450(.A(new_n650), .B1(new_n604), .B2(G107), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n649), .A2(new_n651), .ZN(new_n652));
  NAND4_X1  g0452(.A1(new_n483), .A2(new_n356), .A3(new_n488), .A4(new_n491), .ZN(new_n653));
  NAND3_X1  g0453(.A1(new_n483), .A2(new_n488), .A3(new_n491), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n654), .A2(new_n363), .ZN(new_n655));
  NAND3_X1  g0455(.A1(new_n652), .A2(new_n653), .A3(new_n655), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n630), .A2(new_n632), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n657), .A2(KEYINPUT88), .ZN(new_n658));
  NAND3_X1  g0458(.A1(new_n630), .A2(new_n631), .A3(new_n632), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  INV_X1    g0460(.A(G87), .ZN(new_n661));
  NOR2_X1   g0461(.A1(new_n501), .A2(new_n661), .ZN(new_n662));
  INV_X1    g0462(.A(new_n662), .ZN(new_n663));
  AOI211_X1 g0463(.A(new_n412), .B(new_n638), .C1(new_n642), .C2(new_n279), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n642), .A2(new_n279), .ZN(new_n665));
  INV_X1    g0465(.A(new_n638), .ZN(new_n666));
  AOI21_X1  g0466(.A(new_n414), .B1(new_n665), .B2(new_n666), .ZN(new_n667));
  NOR2_X1   g0467(.A1(new_n664), .A2(new_n667), .ZN(new_n668));
  NAND3_X1  g0468(.A1(new_n660), .A2(new_n663), .A3(new_n668), .ZN(new_n669));
  AND3_X1   g0469(.A1(new_n646), .A2(new_n656), .A3(new_n669), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n597), .A2(new_n599), .ZN(new_n671));
  AOI21_X1  g0471(.A(new_n618), .B1(new_n671), .B2(G190), .ZN(new_n672));
  OAI21_X1  g0472(.A(new_n672), .B1(new_n414), .B2(new_n671), .ZN(new_n673));
  NAND3_X1  g0473(.A1(new_n621), .A2(new_n670), .A3(new_n673), .ZN(new_n674));
  NOR3_X1   g0474(.A1(new_n475), .A2(new_n582), .A3(new_n674), .ZN(G372));
  AND2_X1   g0475(.A1(new_n543), .A2(new_n561), .ZN(new_n676));
  NAND3_X1  g0476(.A1(new_n676), .A2(new_n669), .A3(new_n646), .ZN(new_n677));
  INV_X1    g0477(.A(KEYINPUT26), .ZN(new_n678));
  NOR2_X1   g0478(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  AOI21_X1  g0479(.A(KEYINPUT96), .B1(new_n660), .B2(new_n663), .ZN(new_n680));
  INV_X1    g0480(.A(KEYINPUT96), .ZN(new_n681));
  AOI211_X1 g0481(.A(new_n681), .B(new_n662), .C1(new_n658), .C2(new_n659), .ZN(new_n682));
  OAI21_X1  g0482(.A(new_n668), .B1(new_n680), .B2(new_n682), .ZN(new_n683));
  INV_X1    g0483(.A(KEYINPUT97), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n562), .A2(new_n684), .ZN(new_n685));
  NAND3_X1  g0485(.A1(new_n543), .A2(new_n561), .A3(KEYINPUT97), .ZN(new_n686));
  NAND4_X1  g0486(.A1(new_n683), .A2(new_n685), .A3(new_n646), .A4(new_n686), .ZN(new_n687));
  AOI21_X1  g0487(.A(new_n679), .B1(new_n678), .B2(new_n687), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n602), .A2(new_n618), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n619), .A2(new_n620), .ZN(new_n690));
  NAND3_X1  g0490(.A1(new_n689), .A2(new_n690), .A3(new_n656), .ZN(new_n691));
  INV_X1    g0491(.A(new_n646), .ZN(new_n692));
  OAI21_X1  g0492(.A(new_n663), .B1(new_n633), .B2(new_n634), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n693), .A2(new_n681), .ZN(new_n694));
  NAND3_X1  g0494(.A1(new_n660), .A2(KEYINPUT96), .A3(new_n663), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n694), .A2(new_n695), .ZN(new_n696));
  AOI21_X1  g0496(.A(new_n692), .B1(new_n696), .B2(new_n668), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n691), .A2(new_n697), .ZN(new_n698));
  OAI21_X1  g0498(.A(new_n646), .B1(new_n582), .B2(new_n698), .ZN(new_n699));
  OAI21_X1  g0499(.A(new_n474), .B1(new_n688), .B2(new_n699), .ZN(new_n700));
  INV_X1    g0500(.A(new_n450), .ZN(new_n701));
  AND2_X1   g0501(.A1(new_n404), .A2(new_n411), .ZN(new_n702));
  NAND2_X1  g0502(.A1(new_n326), .A2(G169), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n703), .A2(KEYINPUT14), .ZN(new_n704));
  NAND3_X1  g0504(.A1(new_n326), .A2(new_n337), .A3(G169), .ZN(new_n705));
  NAND3_X1  g0505(.A1(new_n704), .A2(new_n705), .A3(new_n340), .ZN(new_n706));
  INV_X1    g0506(.A(new_n468), .ZN(new_n707));
  AOI22_X1  g0507(.A1(new_n706), .A2(new_n276), .B1(new_n336), .B2(new_n707), .ZN(new_n708));
  AND2_X1   g0508(.A1(new_n419), .A2(new_n420), .ZN(new_n709));
  INV_X1    g0509(.A(new_n709), .ZN(new_n710));
  OAI21_X1  g0510(.A(new_n702), .B1(new_n708), .B2(new_n710), .ZN(new_n711));
  AOI21_X1  g0511(.A(new_n701), .B1(new_n711), .B2(new_n447), .ZN(new_n712));
  NAND2_X1  g0512(.A1(new_n700), .A2(new_n712), .ZN(G369));
  NAND3_X1  g0513(.A1(new_n286), .A2(new_n224), .A3(G13), .ZN(new_n714));
  OR2_X1    g0514(.A1(new_n714), .A2(KEYINPUT27), .ZN(new_n715));
  NAND2_X1  g0515(.A1(new_n714), .A2(KEYINPUT27), .ZN(new_n716));
  NAND3_X1  g0516(.A1(new_n715), .A2(G213), .A3(new_n716), .ZN(new_n717));
  XNOR2_X1  g0517(.A(new_n717), .B(KEYINPUT98), .ZN(new_n718));
  INV_X1    g0518(.A(new_n718), .ZN(new_n719));
  INV_X1    g0519(.A(G343), .ZN(new_n720));
  NOR2_X1   g0520(.A1(new_n719), .A2(new_n720), .ZN(new_n721));
  NAND2_X1  g0521(.A1(new_n721), .A2(new_n618), .ZN(new_n722));
  NAND3_X1  g0522(.A1(new_n621), .A2(new_n673), .A3(new_n722), .ZN(new_n723));
  OAI21_X1  g0523(.A(new_n723), .B1(new_n621), .B2(new_n722), .ZN(new_n724));
  NAND2_X1  g0524(.A1(new_n724), .A2(G330), .ZN(new_n725));
  INV_X1    g0525(.A(new_n526), .ZN(new_n726));
  INV_X1    g0526(.A(new_n721), .ZN(new_n727));
  NOR2_X1   g0527(.A1(new_n727), .A2(new_n521), .ZN(new_n728));
  OAI21_X1  g0528(.A(new_n656), .B1(new_n726), .B2(new_n728), .ZN(new_n729));
  NOR2_X1   g0529(.A1(new_n656), .A2(new_n721), .ZN(new_n730));
  INV_X1    g0530(.A(new_n730), .ZN(new_n731));
  NAND2_X1  g0531(.A1(new_n729), .A2(new_n731), .ZN(new_n732));
  NOR2_X1   g0532(.A1(new_n725), .A2(new_n732), .ZN(new_n733));
  INV_X1    g0533(.A(new_n733), .ZN(new_n734));
  OR2_X1    g0534(.A1(new_n621), .A2(new_n721), .ZN(new_n735));
  OAI21_X1  g0535(.A(new_n731), .B1(new_n732), .B2(new_n735), .ZN(new_n736));
  INV_X1    g0536(.A(new_n736), .ZN(new_n737));
  NAND2_X1  g0537(.A1(new_n734), .A2(new_n737), .ZN(G399));
  NOR2_X1   g0538(.A1(new_n219), .A2(G41), .ZN(new_n739));
  INV_X1    g0539(.A(new_n739), .ZN(new_n740));
  NAND2_X1  g0540(.A1(new_n628), .A2(new_n508), .ZN(new_n741));
  INV_X1    g0541(.A(new_n741), .ZN(new_n742));
  NAND3_X1  g0542(.A1(new_n740), .A2(G1), .A3(new_n742), .ZN(new_n743));
  OAI21_X1  g0543(.A(new_n743), .B1(new_n227), .B2(new_n740), .ZN(new_n744));
  XNOR2_X1  g0544(.A(new_n744), .B(KEYINPUT28), .ZN(new_n745));
  AND3_X1   g0545(.A1(new_n691), .A2(new_n697), .A3(new_n526), .ZN(new_n746));
  OAI21_X1  g0546(.A(new_n562), .B1(new_n578), .B2(new_n581), .ZN(new_n747));
  INV_X1    g0547(.A(KEYINPUT103), .ZN(new_n748));
  NAND2_X1  g0548(.A1(new_n747), .A2(new_n748), .ZN(new_n749));
  INV_X1    g0549(.A(KEYINPUT86), .ZN(new_n750));
  NAND2_X1  g0550(.A1(new_n574), .A2(new_n575), .ZN(new_n751));
  AOI21_X1  g0551(.A(new_n414), .B1(new_n751), .B2(new_n529), .ZN(new_n752));
  OAI211_X1 g0552(.A(new_n560), .B(new_n559), .C1(new_n548), .C2(new_n412), .ZN(new_n753));
  OAI21_X1  g0553(.A(new_n750), .B1(new_n752), .B2(new_n753), .ZN(new_n754));
  AOI21_X1  g0554(.A(new_n676), .B1(new_n754), .B2(new_n577), .ZN(new_n755));
  NAND2_X1  g0555(.A1(new_n755), .A2(KEYINPUT103), .ZN(new_n756));
  NAND3_X1  g0556(.A1(new_n746), .A2(new_n749), .A3(new_n756), .ZN(new_n757));
  AND3_X1   g0557(.A1(new_n543), .A2(new_n561), .A3(KEYINPUT97), .ZN(new_n758));
  AOI21_X1  g0558(.A(KEYINPUT97), .B1(new_n543), .B2(new_n561), .ZN(new_n759));
  NOR2_X1   g0559(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  AOI21_X1  g0560(.A(new_n678), .B1(new_n697), .B2(new_n760), .ZN(new_n761));
  OAI21_X1  g0561(.A(new_n646), .B1(new_n677), .B2(KEYINPUT26), .ZN(new_n762));
  OAI21_X1  g0562(.A(KEYINPUT102), .B1(new_n761), .B2(new_n762), .ZN(new_n763));
  NAND2_X1  g0563(.A1(new_n687), .A2(KEYINPUT26), .ZN(new_n764));
  AND4_X1   g0564(.A1(new_n543), .A2(new_n646), .A3(new_n669), .A4(new_n561), .ZN(new_n765));
  AOI21_X1  g0565(.A(new_n692), .B1(new_n765), .B2(new_n678), .ZN(new_n766));
  INV_X1    g0566(.A(KEYINPUT102), .ZN(new_n767));
  NAND3_X1  g0567(.A1(new_n764), .A2(new_n766), .A3(new_n767), .ZN(new_n768));
  NAND3_X1  g0568(.A1(new_n757), .A2(new_n763), .A3(new_n768), .ZN(new_n769));
  NAND3_X1  g0569(.A1(new_n769), .A2(KEYINPUT29), .A3(new_n727), .ZN(new_n770));
  OAI21_X1  g0570(.A(new_n727), .B1(new_n699), .B2(new_n688), .ZN(new_n771));
  XNOR2_X1  g0571(.A(KEYINPUT101), .B(KEYINPUT29), .ZN(new_n772));
  NAND2_X1  g0572(.A1(new_n771), .A2(new_n772), .ZN(new_n773));
  NAND3_X1  g0573(.A1(new_n483), .A2(new_n643), .A3(new_n491), .ZN(new_n774));
  NOR3_X1   g0574(.A1(new_n548), .A2(new_n774), .A3(new_n601), .ZN(new_n775));
  OAI21_X1  g0575(.A(KEYINPUT30), .B1(new_n775), .B2(KEYINPUT99), .ZN(new_n776));
  INV_X1    g0576(.A(KEYINPUT99), .ZN(new_n777));
  INV_X1    g0577(.A(KEYINPUT30), .ZN(new_n778));
  NAND4_X1  g0578(.A1(new_n571), .A2(G179), .A3(new_n595), .A4(new_n587), .ZN(new_n779));
  OAI211_X1 g0579(.A(new_n777), .B(new_n778), .C1(new_n779), .C2(new_n774), .ZN(new_n780));
  NOR3_X1   g0580(.A1(new_n495), .A2(G179), .A3(new_n643), .ZN(new_n781));
  INV_X1    g0581(.A(new_n599), .ZN(new_n782));
  AOI21_X1  g0582(.A(new_n598), .B1(new_n587), .B2(new_n595), .ZN(new_n783));
  NOR2_X1   g0583(.A1(new_n782), .A2(new_n783), .ZN(new_n784));
  NAND3_X1  g0584(.A1(new_n781), .A2(new_n784), .A3(new_n579), .ZN(new_n785));
  NAND3_X1  g0585(.A1(new_n776), .A2(new_n780), .A3(new_n785), .ZN(new_n786));
  AND3_X1   g0586(.A1(new_n786), .A2(KEYINPUT31), .A3(new_n721), .ZN(new_n787));
  AOI21_X1  g0587(.A(KEYINPUT31), .B1(new_n786), .B2(new_n721), .ZN(new_n788));
  OAI21_X1  g0588(.A(KEYINPUT100), .B1(new_n787), .B2(new_n788), .ZN(new_n789));
  AND3_X1   g0589(.A1(new_n621), .A2(new_n673), .A3(new_n670), .ZN(new_n790));
  NAND4_X1  g0590(.A1(new_n790), .A2(new_n526), .A3(new_n755), .A4(new_n727), .ZN(new_n791));
  NAND2_X1  g0591(.A1(new_n786), .A2(new_n721), .ZN(new_n792));
  INV_X1    g0592(.A(KEYINPUT31), .ZN(new_n793));
  NAND2_X1  g0593(.A1(new_n792), .A2(new_n793), .ZN(new_n794));
  INV_X1    g0594(.A(KEYINPUT100), .ZN(new_n795));
  NAND2_X1  g0595(.A1(new_n794), .A2(new_n795), .ZN(new_n796));
  NAND3_X1  g0596(.A1(new_n789), .A2(new_n791), .A3(new_n796), .ZN(new_n797));
  AOI22_X1  g0597(.A1(new_n770), .A2(new_n773), .B1(G330), .B2(new_n797), .ZN(new_n798));
  OAI21_X1  g0598(.A(new_n745), .B1(new_n798), .B2(G1), .ZN(G364));
  NOR2_X1   g0599(.A1(new_n268), .A2(G20), .ZN(new_n800));
  AOI21_X1  g0600(.A(new_n286), .B1(new_n800), .B2(G45), .ZN(new_n801));
  INV_X1    g0601(.A(new_n801), .ZN(new_n802));
  NOR2_X1   g0602(.A1(new_n739), .A2(new_n802), .ZN(new_n803));
  NAND2_X1  g0603(.A1(new_n310), .A2(new_n218), .ZN(new_n804));
  INV_X1    g0604(.A(G355), .ZN(new_n805));
  OAI22_X1  g0605(.A1(new_n804), .A2(new_n805), .B1(G116), .B2(new_n218), .ZN(new_n806));
  NAND2_X1  g0606(.A1(new_n244), .A2(G45), .ZN(new_n807));
  NOR2_X1   g0607(.A1(new_n219), .A2(new_n310), .ZN(new_n808));
  INV_X1    g0608(.A(new_n808), .ZN(new_n809));
  AOI21_X1  g0609(.A(new_n809), .B1(new_n484), .B2(new_n228), .ZN(new_n810));
  AOI21_X1  g0610(.A(new_n806), .B1(new_n807), .B2(new_n810), .ZN(new_n811));
  NOR2_X1   g0611(.A1(G13), .A2(G33), .ZN(new_n812));
  INV_X1    g0612(.A(new_n812), .ZN(new_n813));
  NOR2_X1   g0613(.A1(new_n813), .A2(G20), .ZN(new_n814));
  AOI21_X1  g0614(.A(new_n223), .B1(G20), .B2(new_n363), .ZN(new_n815));
  NOR2_X1   g0615(.A1(new_n814), .A2(new_n815), .ZN(new_n816));
  INV_X1    g0616(.A(new_n816), .ZN(new_n817));
  OAI21_X1  g0617(.A(new_n803), .B1(new_n811), .B2(new_n817), .ZN(new_n818));
  INV_X1    g0618(.A(G303), .ZN(new_n819));
  NOR2_X1   g0619(.A1(new_n224), .A2(new_n412), .ZN(new_n820));
  NOR2_X1   g0620(.A1(new_n414), .A2(G179), .ZN(new_n821));
  NAND2_X1  g0621(.A1(new_n820), .A2(new_n821), .ZN(new_n822));
  NOR2_X1   g0622(.A1(new_n356), .A2(G200), .ZN(new_n823));
  NAND2_X1  g0623(.A1(new_n820), .A2(new_n823), .ZN(new_n824));
  INV_X1    g0624(.A(G322), .ZN(new_n825));
  OAI22_X1  g0625(.A1(new_n819), .A2(new_n822), .B1(new_n824), .B2(new_n825), .ZN(new_n826));
  NOR2_X1   g0626(.A1(new_n224), .A2(G190), .ZN(new_n827));
  NAND2_X1  g0627(.A1(new_n827), .A2(new_n821), .ZN(new_n828));
  INV_X1    g0628(.A(new_n828), .ZN(new_n829));
  AOI21_X1  g0629(.A(new_n826), .B1(G283), .B2(new_n829), .ZN(new_n830));
  NAND2_X1  g0630(.A1(new_n823), .A2(new_n827), .ZN(new_n831));
  INV_X1    g0631(.A(G311), .ZN(new_n832));
  OAI21_X1  g0632(.A(new_n373), .B1(new_n831), .B2(new_n832), .ZN(new_n833));
  NAND3_X1  g0633(.A1(G20), .A2(G179), .A3(G200), .ZN(new_n834));
  NOR2_X1   g0634(.A1(new_n834), .A2(G190), .ZN(new_n835));
  XNOR2_X1  g0635(.A(KEYINPUT33), .B(G317), .ZN(new_n836));
  AOI21_X1  g0636(.A(new_n833), .B1(new_n835), .B2(new_n836), .ZN(new_n837));
  NOR2_X1   g0637(.A1(G179), .A2(G200), .ZN(new_n838));
  NAND2_X1  g0638(.A1(new_n827), .A2(new_n838), .ZN(new_n839));
  XNOR2_X1  g0639(.A(new_n839), .B(KEYINPUT106), .ZN(new_n840));
  NAND2_X1  g0640(.A1(new_n840), .A2(G329), .ZN(new_n841));
  AOI21_X1  g0641(.A(new_n224), .B1(new_n838), .B2(G190), .ZN(new_n842));
  INV_X1    g0642(.A(new_n842), .ZN(new_n843));
  NOR2_X1   g0643(.A1(new_n834), .A2(new_n412), .ZN(new_n844));
  AOI22_X1  g0644(.A1(new_n843), .A2(G294), .B1(G326), .B2(new_n844), .ZN(new_n845));
  NAND4_X1  g0645(.A1(new_n830), .A2(new_n837), .A3(new_n841), .A4(new_n845), .ZN(new_n846));
  OAI22_X1  g0646(.A1(new_n824), .A2(new_n202), .B1(new_n831), .B2(new_n256), .ZN(new_n847));
  AOI22_X1  g0647(.A1(new_n847), .A2(KEYINPUT104), .B1(G50), .B2(new_n844), .ZN(new_n848));
  OAI21_X1  g0648(.A(new_n848), .B1(KEYINPUT104), .B2(new_n847), .ZN(new_n849));
  XOR2_X1   g0649(.A(new_n849), .B(KEYINPUT105), .Z(new_n850));
  NOR2_X1   g0650(.A1(new_n828), .A2(new_n497), .ZN(new_n851));
  INV_X1    g0651(.A(new_n822), .ZN(new_n852));
  AOI211_X1 g0652(.A(new_n373), .B(new_n851), .C1(G87), .C2(new_n852), .ZN(new_n853));
  NOR2_X1   g0653(.A1(new_n842), .A2(new_n210), .ZN(new_n854));
  AOI21_X1  g0654(.A(new_n854), .B1(new_n835), .B2(G68), .ZN(new_n855));
  NOR2_X1   g0655(.A1(new_n839), .A2(new_n383), .ZN(new_n856));
  XNOR2_X1  g0656(.A(new_n856), .B(KEYINPUT32), .ZN(new_n857));
  NAND3_X1  g0657(.A1(new_n853), .A2(new_n855), .A3(new_n857), .ZN(new_n858));
  OAI21_X1  g0658(.A(new_n846), .B1(new_n850), .B2(new_n858), .ZN(new_n859));
  AOI21_X1  g0659(.A(new_n818), .B1(new_n859), .B2(new_n815), .ZN(new_n860));
  INV_X1    g0660(.A(new_n814), .ZN(new_n861));
  OAI21_X1  g0661(.A(new_n860), .B1(new_n724), .B2(new_n861), .ZN(new_n862));
  INV_X1    g0662(.A(new_n803), .ZN(new_n863));
  NAND2_X1  g0663(.A1(new_n725), .A2(new_n863), .ZN(new_n864));
  NOR2_X1   g0664(.A1(new_n724), .A2(G330), .ZN(new_n865));
  OAI21_X1  g0665(.A(new_n862), .B1(new_n864), .B2(new_n865), .ZN(G396));
  NOR2_X1   g0666(.A1(new_n815), .A2(new_n812), .ZN(new_n867));
  AOI21_X1  g0667(.A(new_n863), .B1(new_n256), .B2(new_n867), .ZN(new_n868));
  INV_X1    g0668(.A(new_n815), .ZN(new_n869));
  NOR2_X1   g0669(.A1(new_n828), .A2(new_n661), .ZN(new_n870));
  INV_X1    g0670(.A(new_n831), .ZN(new_n871));
  AOI21_X1  g0671(.A(new_n870), .B1(G116), .B2(new_n871), .ZN(new_n872));
  INV_X1    g0672(.A(G294), .ZN(new_n873));
  INV_X1    g0673(.A(new_n840), .ZN(new_n874));
  OAI221_X1 g0674(.A(new_n872), .B1(new_n873), .B2(new_n824), .C1(new_n874), .C2(new_n832), .ZN(new_n875));
  OAI21_X1  g0675(.A(new_n373), .B1(new_n822), .B2(new_n497), .ZN(new_n876));
  INV_X1    g0676(.A(new_n835), .ZN(new_n877));
  INV_X1    g0677(.A(G283), .ZN(new_n878));
  INV_X1    g0678(.A(new_n844), .ZN(new_n879));
  OAI22_X1  g0679(.A1(new_n877), .A2(new_n878), .B1(new_n879), .B2(new_n819), .ZN(new_n880));
  NOR4_X1   g0680(.A1(new_n875), .A2(new_n854), .A3(new_n876), .A4(new_n880), .ZN(new_n881));
  AOI21_X1  g0681(.A(new_n373), .B1(new_n829), .B2(G68), .ZN(new_n882));
  OAI221_X1 g0682(.A(new_n882), .B1(new_n201), .B2(new_n822), .C1(new_n202), .C2(new_n842), .ZN(new_n883));
  INV_X1    g0683(.A(new_n824), .ZN(new_n884));
  AOI22_X1  g0684(.A1(G143), .A2(new_n884), .B1(new_n871), .B2(G159), .ZN(new_n885));
  INV_X1    g0685(.A(G137), .ZN(new_n886));
  INV_X1    g0686(.A(G150), .ZN(new_n887));
  OAI221_X1 g0687(.A(new_n885), .B1(new_n879), .B2(new_n886), .C1(new_n887), .C2(new_n877), .ZN(new_n888));
  INV_X1    g0688(.A(KEYINPUT34), .ZN(new_n889));
  NOR2_X1   g0689(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  AOI211_X1 g0690(.A(new_n883), .B(new_n890), .C1(G132), .C2(new_n840), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n888), .A2(new_n889), .ZN(new_n892));
  AOI21_X1  g0692(.A(new_n881), .B1(new_n891), .B2(new_n892), .ZN(new_n893));
  OAI21_X1  g0693(.A(new_n472), .B1(new_n469), .B2(new_n727), .ZN(new_n894));
  NAND4_X1  g0694(.A1(new_n456), .A2(new_n466), .A3(new_n467), .A4(new_n721), .ZN(new_n895));
  INV_X1    g0695(.A(KEYINPUT107), .ZN(new_n896));
  XNOR2_X1  g0696(.A(new_n895), .B(new_n896), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n894), .A2(new_n897), .ZN(new_n898));
  OAI221_X1 g0698(.A(new_n868), .B1(new_n869), .B2(new_n893), .C1(new_n898), .C2(new_n813), .ZN(new_n899));
  INV_X1    g0699(.A(new_n898), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n771), .A2(new_n900), .ZN(new_n901));
  AOI21_X1  g0701(.A(new_n721), .B1(new_n894), .B2(new_n897), .ZN(new_n902));
  OAI21_X1  g0702(.A(new_n902), .B1(new_n699), .B2(new_n688), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n901), .A2(new_n903), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n797), .A2(G330), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n906), .A2(new_n863), .ZN(new_n907));
  NOR2_X1   g0707(.A1(new_n904), .A2(new_n905), .ZN(new_n908));
  OAI21_X1  g0708(.A(new_n899), .B1(new_n907), .B2(new_n908), .ZN(G384));
  NOR2_X1   g0709(.A1(new_n800), .A2(new_n286), .ZN(new_n910));
  INV_X1    g0710(.A(new_n336), .ZN(new_n911));
  OAI211_X1 g0711(.A(new_n276), .B(new_n721), .C1(new_n911), .C2(new_n706), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n721), .A2(new_n276), .ZN(new_n913));
  OAI211_X1 g0713(.A(new_n336), .B(new_n913), .C1(new_n342), .C2(new_n343), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n912), .A2(new_n914), .ZN(new_n915));
  NOR2_X1   g0715(.A1(new_n787), .A2(new_n788), .ZN(new_n916));
  AOI21_X1  g0716(.A(new_n900), .B1(new_n791), .B2(new_n916), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n407), .A2(new_n371), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n918), .A2(new_n718), .ZN(new_n919));
  INV_X1    g0719(.A(new_n919), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n421), .A2(new_n920), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n366), .A2(new_n402), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n402), .A2(new_n718), .ZN(new_n923));
  INV_X1    g0723(.A(KEYINPUT37), .ZN(new_n924));
  NAND4_X1  g0724(.A1(new_n922), .A2(new_n923), .A3(new_n924), .A4(new_n417), .ZN(new_n925));
  NAND4_X1  g0725(.A1(new_n359), .A2(new_n918), .A3(new_n364), .A4(new_n365), .ZN(new_n926));
  NAND3_X1  g0726(.A1(new_n417), .A2(new_n926), .A3(new_n919), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n927), .A2(KEYINPUT37), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n925), .A2(new_n928), .ZN(new_n929));
  NAND4_X1  g0729(.A1(new_n921), .A2(KEYINPUT110), .A3(new_n929), .A4(KEYINPUT38), .ZN(new_n930));
  AOI22_X1  g0730(.A1(new_n421), .A2(new_n920), .B1(new_n925), .B2(new_n928), .ZN(new_n931));
  OAI21_X1  g0731(.A(new_n930), .B1(KEYINPUT38), .B2(new_n931), .ZN(new_n932));
  AOI21_X1  g0732(.A(KEYINPUT110), .B1(new_n931), .B2(KEYINPUT38), .ZN(new_n933));
  OAI211_X1 g0733(.A(new_n915), .B(new_n917), .C1(new_n932), .C2(new_n933), .ZN(new_n934));
  INV_X1    g0734(.A(KEYINPUT40), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n934), .A2(new_n935), .ZN(new_n936));
  INV_X1    g0736(.A(KEYINPUT38), .ZN(new_n937));
  OAI21_X1  g0737(.A(new_n417), .B1(new_n409), .B2(new_n410), .ZN(new_n938));
  NOR2_X1   g0738(.A1(new_n409), .A2(new_n719), .ZN(new_n939));
  NOR2_X1   g0739(.A1(new_n938), .A2(new_n939), .ZN(new_n940));
  INV_X1    g0740(.A(KEYINPUT111), .ZN(new_n941));
  AOI21_X1  g0741(.A(new_n924), .B1(new_n923), .B2(new_n941), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n940), .A2(new_n942), .ZN(new_n943));
  AOI21_X1  g0743(.A(KEYINPUT111), .B1(new_n402), .B2(new_n718), .ZN(new_n944));
  OAI22_X1  g0744(.A1(new_n938), .A2(new_n939), .B1(new_n944), .B2(new_n924), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n943), .A2(new_n945), .ZN(new_n946));
  AOI21_X1  g0746(.A(new_n923), .B1(new_n702), .B2(new_n709), .ZN(new_n947));
  OAI21_X1  g0747(.A(new_n937), .B1(new_n946), .B2(new_n947), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n931), .A2(KEYINPUT38), .ZN(new_n949));
  NAND2_X1  g0749(.A1(new_n948), .A2(new_n949), .ZN(new_n950));
  NAND4_X1  g0750(.A1(new_n950), .A2(new_n915), .A3(KEYINPUT40), .A4(new_n917), .ZN(new_n951));
  AND2_X1   g0751(.A1(new_n936), .A2(new_n951), .ZN(new_n952));
  NOR3_X1   g0752(.A1(new_n582), .A2(new_n674), .A3(new_n721), .ZN(new_n953));
  NAND3_X1  g0753(.A1(new_n786), .A2(KEYINPUT31), .A3(new_n721), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n794), .A2(new_n954), .ZN(new_n955));
  NOR2_X1   g0755(.A1(new_n953), .A2(new_n955), .ZN(new_n956));
  NOR2_X1   g0756(.A1(new_n475), .A2(new_n956), .ZN(new_n957));
  NOR2_X1   g0757(.A1(new_n952), .A2(new_n957), .ZN(new_n958));
  INV_X1    g0758(.A(G330), .ZN(new_n959));
  NOR2_X1   g0759(.A1(new_n958), .A2(new_n959), .ZN(new_n960));
  AOI22_X1  g0760(.A1(new_n960), .A2(KEYINPUT112), .B1(new_n952), .B2(new_n957), .ZN(new_n961));
  OAI21_X1  g0761(.A(new_n961), .B1(KEYINPUT112), .B2(new_n960), .ZN(new_n962));
  OAI21_X1  g0762(.A(KEYINPUT39), .B1(new_n932), .B2(new_n933), .ZN(new_n963));
  INV_X1    g0763(.A(KEYINPUT39), .ZN(new_n964));
  NAND3_X1  g0764(.A1(new_n948), .A2(new_n964), .A3(new_n949), .ZN(new_n965));
  NAND2_X1  g0765(.A1(new_n963), .A2(new_n965), .ZN(new_n966));
  NAND3_X1  g0766(.A1(new_n706), .A2(new_n276), .A3(new_n727), .ZN(new_n967));
  INV_X1    g0767(.A(new_n967), .ZN(new_n968));
  NAND2_X1  g0768(.A1(new_n966), .A2(new_n968), .ZN(new_n969));
  AOI21_X1  g0769(.A(KEYINPUT38), .B1(new_n921), .B2(new_n929), .ZN(new_n970));
  AND3_X1   g0770(.A1(new_n921), .A2(KEYINPUT38), .A3(new_n929), .ZN(new_n971));
  AOI21_X1  g0771(.A(new_n970), .B1(new_n971), .B2(KEYINPUT110), .ZN(new_n972));
  INV_X1    g0772(.A(new_n933), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n972), .A2(new_n973), .ZN(new_n974));
  INV_X1    g0774(.A(KEYINPUT109), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n707), .A2(new_n727), .ZN(new_n976));
  XNOR2_X1  g0776(.A(new_n976), .B(KEYINPUT108), .ZN(new_n977));
  AND3_X1   g0777(.A1(new_n903), .A2(new_n975), .A3(new_n977), .ZN(new_n978));
  AOI21_X1  g0778(.A(new_n975), .B1(new_n903), .B2(new_n977), .ZN(new_n979));
  OAI211_X1 g0779(.A(new_n974), .B(new_n915), .C1(new_n978), .C2(new_n979), .ZN(new_n980));
  INV_X1    g0780(.A(new_n702), .ZN(new_n981));
  NAND2_X1  g0781(.A1(new_n981), .A2(new_n719), .ZN(new_n982));
  NAND3_X1  g0782(.A1(new_n969), .A2(new_n980), .A3(new_n982), .ZN(new_n983));
  NAND3_X1  g0783(.A1(new_n770), .A2(new_n474), .A3(new_n773), .ZN(new_n984));
  NAND2_X1  g0784(.A1(new_n984), .A2(new_n712), .ZN(new_n985));
  XNOR2_X1  g0785(.A(new_n983), .B(new_n985), .ZN(new_n986));
  AOI21_X1  g0786(.A(new_n910), .B1(new_n962), .B2(new_n986), .ZN(new_n987));
  OAI21_X1  g0787(.A(new_n987), .B1(new_n986), .B2(new_n962), .ZN(new_n988));
  OR2_X1    g0788(.A1(new_n556), .A2(KEYINPUT35), .ZN(new_n989));
  NAND2_X1  g0789(.A1(new_n556), .A2(KEYINPUT35), .ZN(new_n990));
  NAND4_X1  g0790(.A1(new_n989), .A2(new_n990), .A3(G116), .A4(new_n225), .ZN(new_n991));
  XNOR2_X1  g0791(.A(new_n991), .B(KEYINPUT36), .ZN(new_n992));
  NAND4_X1  g0792(.A1(new_n228), .A2(G77), .A3(new_n380), .A4(new_n381), .ZN(new_n993));
  OAI21_X1  g0793(.A(new_n993), .B1(G50), .B2(new_n203), .ZN(new_n994));
  NAND3_X1  g0794(.A1(new_n994), .A2(G1), .A3(new_n268), .ZN(new_n995));
  NAND3_X1  g0795(.A1(new_n988), .A2(new_n992), .A3(new_n995), .ZN(G367));
  INV_X1    g0796(.A(new_n839), .ZN(new_n997));
  AOI22_X1  g0797(.A1(new_n871), .A2(G50), .B1(new_n997), .B2(G137), .ZN(new_n998));
  OAI221_X1 g0798(.A(new_n998), .B1(new_n256), .B2(new_n828), .C1(new_n887), .C2(new_n824), .ZN(new_n999));
  NOR2_X1   g0799(.A1(new_n842), .A2(new_n203), .ZN(new_n1000));
  INV_X1    g0800(.A(G143), .ZN(new_n1001));
  OAI22_X1  g0801(.A1(new_n877), .A2(new_n383), .B1(new_n879), .B2(new_n1001), .ZN(new_n1002));
  OAI21_X1  g0802(.A(new_n310), .B1(new_n822), .B2(new_n202), .ZN(new_n1003));
  NOR4_X1   g0803(.A1(new_n999), .A2(new_n1000), .A3(new_n1002), .A4(new_n1003), .ZN(new_n1004));
  NOR2_X1   g0804(.A1(new_n822), .A2(new_n508), .ZN(new_n1005));
  AOI22_X1  g0805(.A1(new_n1005), .A2(KEYINPUT46), .B1(G294), .B2(new_n835), .ZN(new_n1006));
  OAI221_X1 g0806(.A(new_n1006), .B1(new_n497), .B2(new_n842), .C1(new_n832), .C2(new_n879), .ZN(new_n1007));
  AOI22_X1  g0807(.A1(G303), .A2(new_n884), .B1(new_n829), .B2(G97), .ZN(new_n1008));
  INV_X1    g0808(.A(G317), .ZN(new_n1009));
  OAI21_X1  g0809(.A(new_n1008), .B1(new_n1009), .B2(new_n839), .ZN(new_n1010));
  OAI221_X1 g0810(.A(new_n373), .B1(new_n878), .B2(new_n831), .C1(new_n1005), .C2(KEYINPUT46), .ZN(new_n1011));
  NOR3_X1   g0811(.A1(new_n1007), .A2(new_n1010), .A3(new_n1011), .ZN(new_n1012));
  NOR2_X1   g0812(.A1(new_n1004), .A2(new_n1012), .ZN(new_n1013));
  XOR2_X1   g0813(.A(new_n1013), .B(KEYINPUT47), .Z(new_n1014));
  NAND2_X1  g0814(.A1(new_n1014), .A2(new_n815), .ZN(new_n1015));
  AOI21_X1  g0815(.A(new_n817), .B1(new_n219), .B2(new_n458), .ZN(new_n1016));
  NAND2_X1  g0816(.A1(new_n239), .A2(new_n808), .ZN(new_n1017));
  AOI21_X1  g0817(.A(new_n863), .B1(new_n1016), .B2(new_n1017), .ZN(new_n1018));
  NAND3_X1  g0818(.A1(new_n694), .A2(new_n695), .A3(new_n721), .ZN(new_n1019));
  NAND2_X1  g0819(.A1(new_n697), .A2(new_n1019), .ZN(new_n1020));
  OR2_X1    g0820(.A1(new_n1019), .A2(new_n646), .ZN(new_n1021));
  NAND2_X1  g0821(.A1(new_n1020), .A2(new_n1021), .ZN(new_n1022));
  OAI211_X1 g0822(.A(new_n1015), .B(new_n1018), .C1(new_n1022), .C2(new_n861), .ZN(new_n1023));
  NAND2_X1  g0823(.A1(new_n721), .A2(new_n570), .ZN(new_n1024));
  NAND3_X1  g0824(.A1(new_n749), .A2(new_n756), .A3(new_n1024), .ZN(new_n1025));
  NAND2_X1  g0825(.A1(new_n676), .A2(new_n721), .ZN(new_n1026));
  AND2_X1   g0826(.A1(new_n1025), .A2(new_n1026), .ZN(new_n1027));
  NAND2_X1  g0827(.A1(new_n1027), .A2(new_n736), .ZN(new_n1028));
  INV_X1    g0828(.A(KEYINPUT44), .ZN(new_n1029));
  XNOR2_X1  g0829(.A(new_n1028), .B(new_n1029), .ZN(new_n1030));
  INV_X1    g0830(.A(new_n1027), .ZN(new_n1031));
  NAND3_X1  g0831(.A1(new_n1031), .A2(KEYINPUT45), .A3(new_n737), .ZN(new_n1032));
  INV_X1    g0832(.A(KEYINPUT45), .ZN(new_n1033));
  OAI21_X1  g0833(.A(new_n1033), .B1(new_n1027), .B2(new_n736), .ZN(new_n1034));
  NAND2_X1  g0834(.A1(new_n1032), .A2(new_n1034), .ZN(new_n1035));
  NAND2_X1  g0835(.A1(new_n1030), .A2(new_n1035), .ZN(new_n1036));
  NAND2_X1  g0836(.A1(new_n1036), .A2(new_n733), .ZN(new_n1037));
  XOR2_X1   g0837(.A(new_n732), .B(new_n735), .Z(new_n1038));
  XNOR2_X1  g0838(.A(new_n1038), .B(new_n725), .ZN(new_n1039));
  AND2_X1   g0839(.A1(new_n1039), .A2(new_n798), .ZN(new_n1040));
  NAND3_X1  g0840(.A1(new_n1030), .A2(new_n734), .A3(new_n1035), .ZN(new_n1041));
  NAND3_X1  g0841(.A1(new_n1037), .A2(new_n1040), .A3(new_n1041), .ZN(new_n1042));
  NAND2_X1  g0842(.A1(new_n1042), .A2(new_n798), .ZN(new_n1043));
  XOR2_X1   g0843(.A(new_n739), .B(KEYINPUT41), .Z(new_n1044));
  INV_X1    g0844(.A(new_n1044), .ZN(new_n1045));
  NAND2_X1  g0845(.A1(new_n1043), .A2(new_n1045), .ZN(new_n1046));
  NAND2_X1  g0846(.A1(new_n1046), .A2(KEYINPUT113), .ZN(new_n1047));
  INV_X1    g0847(.A(KEYINPUT113), .ZN(new_n1048));
  NAND3_X1  g0848(.A1(new_n1043), .A2(new_n1048), .A3(new_n1045), .ZN(new_n1049));
  AOI21_X1  g0849(.A(new_n802), .B1(new_n1047), .B2(new_n1049), .ZN(new_n1050));
  OR3_X1    g0850(.A1(new_n1027), .A2(new_n732), .A3(new_n735), .ZN(new_n1051));
  NOR2_X1   g0851(.A1(new_n1051), .A2(KEYINPUT42), .ZN(new_n1052));
  INV_X1    g0852(.A(new_n1052), .ZN(new_n1053));
  OR2_X1    g0853(.A1(new_n1025), .A2(new_n656), .ZN(new_n1054));
  AOI21_X1  g0854(.A(new_n721), .B1(new_n1054), .B2(new_n562), .ZN(new_n1055));
  AOI21_X1  g0855(.A(new_n1055), .B1(new_n1051), .B2(KEYINPUT42), .ZN(new_n1056));
  AOI22_X1  g0856(.A1(new_n1053), .A2(new_n1056), .B1(KEYINPUT43), .B2(new_n1022), .ZN(new_n1057));
  NOR2_X1   g0857(.A1(new_n1022), .A2(KEYINPUT43), .ZN(new_n1058));
  INV_X1    g0858(.A(new_n1058), .ZN(new_n1059));
  OR2_X1    g0859(.A1(new_n1057), .A2(new_n1059), .ZN(new_n1060));
  NAND2_X1  g0860(.A1(new_n1057), .A2(new_n1059), .ZN(new_n1061));
  NAND2_X1  g0861(.A1(new_n1060), .A2(new_n1061), .ZN(new_n1062));
  NOR2_X1   g0862(.A1(new_n734), .A2(new_n1027), .ZN(new_n1063));
  INV_X1    g0863(.A(new_n1063), .ZN(new_n1064));
  NAND2_X1  g0864(.A1(new_n1062), .A2(new_n1064), .ZN(new_n1065));
  NAND3_X1  g0865(.A1(new_n1060), .A2(new_n1063), .A3(new_n1061), .ZN(new_n1066));
  NAND2_X1  g0866(.A1(new_n1065), .A2(new_n1066), .ZN(new_n1067));
  OAI21_X1  g0867(.A(new_n1023), .B1(new_n1050), .B2(new_n1067), .ZN(G387));
  OAI22_X1  g0868(.A1(new_n742), .A2(new_n804), .B1(G107), .B2(new_n218), .ZN(new_n1069));
  XOR2_X1   g0869(.A(new_n1069), .B(KEYINPUT114), .Z(new_n1070));
  NAND2_X1  g0870(.A1(new_n236), .A2(G45), .ZN(new_n1071));
  NAND2_X1  g0871(.A1(new_n368), .A2(new_n201), .ZN(new_n1072));
  XOR2_X1   g0872(.A(new_n1072), .B(KEYINPUT50), .Z(new_n1073));
  AOI211_X1 g0873(.A(G45), .B(new_n741), .C1(G68), .C2(G77), .ZN(new_n1074));
  AOI21_X1  g0874(.A(new_n809), .B1(new_n1073), .B2(new_n1074), .ZN(new_n1075));
  AOI21_X1  g0875(.A(new_n1070), .B1(new_n1071), .B2(new_n1075), .ZN(new_n1076));
  OAI21_X1  g0876(.A(new_n803), .B1(new_n1076), .B2(new_n817), .ZN(new_n1077));
  XOR2_X1   g0877(.A(new_n1077), .B(KEYINPUT115), .Z(new_n1078));
  OAI221_X1 g0878(.A(new_n310), .B1(new_n210), .B2(new_n828), .C1(new_n369), .C2(new_n877), .ZN(new_n1079));
  OAI22_X1  g0879(.A1(new_n879), .A2(new_n383), .B1(new_n842), .B2(new_n457), .ZN(new_n1080));
  OAI22_X1  g0880(.A1(new_n831), .A2(new_n203), .B1(new_n839), .B2(new_n887), .ZN(new_n1081));
  OAI22_X1  g0881(.A1(new_n201), .A2(new_n824), .B1(new_n822), .B2(new_n256), .ZN(new_n1082));
  NOR4_X1   g0882(.A1(new_n1079), .A2(new_n1080), .A3(new_n1081), .A4(new_n1082), .ZN(new_n1083));
  OAI22_X1  g0883(.A1(new_n822), .A2(new_n873), .B1(new_n842), .B2(new_n878), .ZN(new_n1084));
  AOI22_X1  g0884(.A1(G317), .A2(new_n884), .B1(new_n871), .B2(G303), .ZN(new_n1085));
  OAI221_X1 g0885(.A(new_n1085), .B1(new_n879), .B2(new_n825), .C1(new_n832), .C2(new_n877), .ZN(new_n1086));
  INV_X1    g0886(.A(KEYINPUT48), .ZN(new_n1087));
  AOI21_X1  g0887(.A(new_n1084), .B1(new_n1086), .B2(new_n1087), .ZN(new_n1088));
  OAI21_X1  g0888(.A(new_n1088), .B1(new_n1087), .B2(new_n1086), .ZN(new_n1089));
  XOR2_X1   g0889(.A(new_n1089), .B(KEYINPUT49), .Z(new_n1090));
  OR2_X1    g0890(.A1(new_n1090), .A2(KEYINPUT116), .ZN(new_n1091));
  AOI21_X1  g0891(.A(new_n310), .B1(new_n997), .B2(G326), .ZN(new_n1092));
  OAI21_X1  g0892(.A(new_n1092), .B1(new_n508), .B2(new_n828), .ZN(new_n1093));
  AOI21_X1  g0893(.A(new_n1093), .B1(new_n1090), .B2(KEYINPUT116), .ZN(new_n1094));
  AOI21_X1  g0894(.A(new_n1083), .B1(new_n1091), .B2(new_n1094), .ZN(new_n1095));
  OAI21_X1  g0895(.A(new_n1078), .B1(new_n1095), .B2(new_n869), .ZN(new_n1096));
  AOI21_X1  g0896(.A(new_n1096), .B1(new_n732), .B2(new_n814), .ZN(new_n1097));
  AOI21_X1  g0897(.A(new_n1097), .B1(new_n1039), .B2(new_n802), .ZN(new_n1098));
  OR2_X1    g0898(.A1(new_n1040), .A2(new_n740), .ZN(new_n1099));
  NOR2_X1   g0899(.A1(new_n1039), .A2(new_n798), .ZN(new_n1100));
  OAI21_X1  g0900(.A(new_n1098), .B1(new_n1099), .B2(new_n1100), .ZN(G393));
  NAND3_X1  g0901(.A1(new_n1037), .A2(new_n802), .A3(new_n1041), .ZN(new_n1102));
  AOI21_X1  g0902(.A(new_n817), .B1(G97), .B2(new_n219), .ZN(new_n1103));
  NAND2_X1  g0903(.A1(new_n247), .A2(new_n808), .ZN(new_n1104));
  AOI21_X1  g0904(.A(new_n863), .B1(new_n1103), .B2(new_n1104), .ZN(new_n1105));
  AOI211_X1 g0905(.A(new_n310), .B(new_n851), .C1(G303), .C2(new_n835), .ZN(new_n1106));
  OAI22_X1  g0906(.A1(new_n831), .A2(new_n873), .B1(new_n839), .B2(new_n825), .ZN(new_n1107));
  AOI21_X1  g0907(.A(new_n1107), .B1(G283), .B2(new_n852), .ZN(new_n1108));
  OAI211_X1 g0908(.A(new_n1106), .B(new_n1108), .C1(new_n508), .C2(new_n842), .ZN(new_n1109));
  AOI22_X1  g0909(.A1(new_n884), .A2(G311), .B1(G317), .B2(new_n844), .ZN(new_n1110));
  XNOR2_X1  g0910(.A(new_n1110), .B(KEYINPUT52), .ZN(new_n1111));
  NOR2_X1   g0911(.A1(new_n1109), .A2(new_n1111), .ZN(new_n1112));
  OR2_X1    g0912(.A1(new_n1112), .A2(KEYINPUT118), .ZN(new_n1113));
  NAND2_X1  g0913(.A1(new_n1112), .A2(KEYINPUT118), .ZN(new_n1114));
  AOI22_X1  g0914(.A1(new_n871), .A2(new_n368), .B1(G50), .B2(new_n835), .ZN(new_n1115));
  INV_X1    g0915(.A(new_n1115), .ZN(new_n1116));
  OR2_X1    g0916(.A1(new_n1116), .A2(KEYINPUT117), .ZN(new_n1117));
  OAI22_X1  g0917(.A1(new_n879), .A2(new_n887), .B1(new_n824), .B2(new_n383), .ZN(new_n1118));
  XNOR2_X1  g0918(.A(new_n1118), .B(KEYINPUT51), .ZN(new_n1119));
  NAND2_X1  g0919(.A1(new_n1116), .A2(KEYINPUT117), .ZN(new_n1120));
  OAI22_X1  g0920(.A1(new_n822), .A2(new_n203), .B1(new_n839), .B2(new_n1001), .ZN(new_n1121));
  NOR2_X1   g0921(.A1(new_n842), .A2(new_n256), .ZN(new_n1122));
  NOR4_X1   g0922(.A1(new_n1121), .A2(new_n870), .A3(new_n1122), .A4(new_n373), .ZN(new_n1123));
  NAND4_X1  g0923(.A1(new_n1117), .A2(new_n1119), .A3(new_n1120), .A4(new_n1123), .ZN(new_n1124));
  AND3_X1   g0924(.A1(new_n1113), .A2(new_n1114), .A3(new_n1124), .ZN(new_n1125));
  OAI221_X1 g0925(.A(new_n1105), .B1(new_n869), .B2(new_n1125), .C1(new_n1031), .C2(new_n861), .ZN(new_n1126));
  NAND2_X1  g0926(.A1(new_n1102), .A2(new_n1126), .ZN(new_n1127));
  AND2_X1   g0927(.A1(new_n1037), .A2(new_n1041), .ZN(new_n1128));
  OR2_X1    g0928(.A1(new_n1128), .A2(new_n1040), .ZN(new_n1129));
  AND2_X1   g0929(.A1(new_n1042), .A2(new_n739), .ZN(new_n1130));
  AOI21_X1  g0930(.A(new_n1127), .B1(new_n1129), .B2(new_n1130), .ZN(new_n1131));
  INV_X1    g0931(.A(new_n1131), .ZN(G390));
  NAND3_X1  g0932(.A1(new_n915), .A2(G330), .A3(new_n917), .ZN(new_n1133));
  INV_X1    g0933(.A(new_n1133), .ZN(new_n1134));
  OAI21_X1  g0934(.A(new_n915), .B1(new_n978), .B2(new_n979), .ZN(new_n1135));
  AOI21_X1  g0935(.A(new_n966), .B1(new_n1135), .B2(new_n967), .ZN(new_n1136));
  NAND2_X1  g0936(.A1(new_n950), .A2(new_n967), .ZN(new_n1137));
  NAND3_X1  g0937(.A1(new_n769), .A2(new_n727), .A3(new_n898), .ZN(new_n1138));
  NAND2_X1  g0938(.A1(new_n1138), .A2(new_n977), .ZN(new_n1139));
  AOI21_X1  g0939(.A(new_n1137), .B1(new_n1139), .B2(new_n915), .ZN(new_n1140));
  OAI21_X1  g0940(.A(new_n1134), .B1(new_n1136), .B2(new_n1140), .ZN(new_n1141));
  INV_X1    g0941(.A(new_n966), .ZN(new_n1142));
  AND2_X1   g0942(.A1(new_n912), .A2(new_n914), .ZN(new_n1143));
  NAND2_X1  g0943(.A1(new_n898), .A2(new_n727), .ZN(new_n1144));
  NAND2_X1  g0944(.A1(new_n754), .A2(new_n577), .ZN(new_n1145));
  AND3_X1   g0945(.A1(new_n1145), .A2(new_n526), .A3(new_n562), .ZN(new_n1146));
  AND2_X1   g0946(.A1(new_n691), .A2(new_n697), .ZN(new_n1147));
  AOI21_X1  g0947(.A(new_n692), .B1(new_n1146), .B2(new_n1147), .ZN(new_n1148));
  NAND2_X1  g0948(.A1(new_n687), .A2(new_n678), .ZN(new_n1149));
  OAI21_X1  g0949(.A(new_n1149), .B1(new_n678), .B2(new_n677), .ZN(new_n1150));
  AOI21_X1  g0950(.A(new_n1144), .B1(new_n1148), .B2(new_n1150), .ZN(new_n1151));
  INV_X1    g0951(.A(new_n977), .ZN(new_n1152));
  OAI21_X1  g0952(.A(KEYINPUT109), .B1(new_n1151), .B2(new_n1152), .ZN(new_n1153));
  NAND3_X1  g0953(.A1(new_n903), .A2(new_n975), .A3(new_n977), .ZN(new_n1154));
  AOI21_X1  g0954(.A(new_n1143), .B1(new_n1153), .B2(new_n1154), .ZN(new_n1155));
  OAI21_X1  g0955(.A(new_n1142), .B1(new_n1155), .B2(new_n968), .ZN(new_n1156));
  NAND4_X1  g0956(.A1(new_n915), .A2(G330), .A3(new_n797), .A4(new_n898), .ZN(new_n1157));
  INV_X1    g0957(.A(new_n1140), .ZN(new_n1158));
  NAND3_X1  g0958(.A1(new_n1156), .A2(new_n1157), .A3(new_n1158), .ZN(new_n1159));
  NAND2_X1  g0959(.A1(new_n1141), .A2(new_n1159), .ZN(new_n1160));
  OAI211_X1 g0960(.A(new_n474), .B(G330), .C1(new_n953), .C2(new_n955), .ZN(new_n1161));
  NAND3_X1  g0961(.A1(new_n984), .A2(new_n712), .A3(new_n1161), .ZN(new_n1162));
  INV_X1    g0962(.A(new_n1162), .ZN(new_n1163));
  OAI21_X1  g0963(.A(new_n898), .B1(new_n953), .B2(new_n955), .ZN(new_n1164));
  OAI21_X1  g0964(.A(new_n1143), .B1(new_n959), .B2(new_n1164), .ZN(new_n1165));
  NAND4_X1  g0965(.A1(new_n1165), .A2(new_n1157), .A3(new_n977), .A4(new_n1138), .ZN(new_n1166));
  INV_X1    g0966(.A(new_n1166), .ZN(new_n1167));
  NAND3_X1  g0967(.A1(new_n797), .A2(G330), .A3(new_n898), .ZN(new_n1168));
  NAND2_X1  g0968(.A1(new_n1168), .A2(new_n1143), .ZN(new_n1169));
  AOI22_X1  g0969(.A1(new_n1133), .A2(new_n1169), .B1(new_n1153), .B2(new_n1154), .ZN(new_n1170));
  OAI21_X1  g0970(.A(new_n1163), .B1(new_n1167), .B2(new_n1170), .ZN(new_n1171));
  NAND2_X1  g0971(.A1(new_n1160), .A2(new_n1171), .ZN(new_n1172));
  NAND2_X1  g0972(.A1(new_n1169), .A2(new_n1133), .ZN(new_n1173));
  NAND2_X1  g0973(.A1(new_n1153), .A2(new_n1154), .ZN(new_n1174));
  NAND2_X1  g0974(.A1(new_n1173), .A2(new_n1174), .ZN(new_n1175));
  AOI21_X1  g0975(.A(new_n1162), .B1(new_n1175), .B2(new_n1166), .ZN(new_n1176));
  NAND3_X1  g0976(.A1(new_n1141), .A2(new_n1159), .A3(new_n1176), .ZN(new_n1177));
  NAND3_X1  g0977(.A1(new_n1172), .A2(new_n739), .A3(new_n1177), .ZN(new_n1178));
  NAND3_X1  g0978(.A1(new_n1141), .A2(new_n1159), .A3(new_n802), .ZN(new_n1179));
  AOI21_X1  g0979(.A(new_n863), .B1(new_n369), .B2(new_n867), .ZN(new_n1180));
  AOI211_X1 g0980(.A(new_n310), .B(new_n1122), .C1(G87), .C2(new_n852), .ZN(new_n1181));
  AOI22_X1  g0981(.A1(G107), .A2(new_n835), .B1(new_n844), .B2(G283), .ZN(new_n1182));
  OAI22_X1  g0982(.A1(new_n203), .A2(new_n828), .B1(new_n831), .B2(new_n210), .ZN(new_n1183));
  AOI21_X1  g0983(.A(new_n1183), .B1(G116), .B2(new_n884), .ZN(new_n1184));
  NAND2_X1  g0984(.A1(new_n840), .A2(G294), .ZN(new_n1185));
  NAND4_X1  g0985(.A1(new_n1181), .A2(new_n1182), .A3(new_n1184), .A4(new_n1185), .ZN(new_n1186));
  INV_X1    g0986(.A(G125), .ZN(new_n1187));
  OAI221_X1 g0987(.A(new_n310), .B1(new_n201), .B2(new_n828), .C1(new_n874), .C2(new_n1187), .ZN(new_n1188));
  XOR2_X1   g0988(.A(new_n1188), .B(KEYINPUT119), .Z(new_n1189));
  NOR2_X1   g0989(.A1(new_n822), .A2(new_n887), .ZN(new_n1190));
  INV_X1    g0990(.A(KEYINPUT53), .ZN(new_n1191));
  NAND2_X1  g0991(.A1(new_n1190), .A2(new_n1191), .ZN(new_n1192));
  INV_X1    g0992(.A(G132), .ZN(new_n1193));
  XNOR2_X1  g0993(.A(KEYINPUT54), .B(G143), .ZN(new_n1194));
  OAI221_X1 g0994(.A(new_n1192), .B1(new_n1193), .B2(new_n824), .C1(new_n831), .C2(new_n1194), .ZN(new_n1195));
  AOI22_X1  g0995(.A1(new_n843), .A2(G159), .B1(G137), .B2(new_n835), .ZN(new_n1196));
  INV_X1    g0996(.A(G128), .ZN(new_n1197));
  OAI221_X1 g0997(.A(new_n1196), .B1(new_n1191), .B2(new_n1190), .C1(new_n1197), .C2(new_n879), .ZN(new_n1198));
  OR2_X1    g0998(.A1(new_n1195), .A2(new_n1198), .ZN(new_n1199));
  OAI21_X1  g0999(.A(new_n1186), .B1(new_n1189), .B2(new_n1199), .ZN(new_n1200));
  INV_X1    g1000(.A(KEYINPUT120), .ZN(new_n1201));
  NOR2_X1   g1001(.A1(new_n1200), .A2(new_n1201), .ZN(new_n1202));
  NAND2_X1  g1002(.A1(new_n1200), .A2(new_n1201), .ZN(new_n1203));
  NAND2_X1  g1003(.A1(new_n1203), .A2(new_n815), .ZN(new_n1204));
  OAI221_X1 g1004(.A(new_n1180), .B1(new_n1202), .B2(new_n1204), .C1(new_n966), .C2(new_n813), .ZN(new_n1205));
  AND2_X1   g1005(.A1(new_n1179), .A2(new_n1205), .ZN(new_n1206));
  NAND2_X1  g1006(.A1(new_n1178), .A2(new_n1206), .ZN(G378));
  NAND2_X1  g1007(.A1(new_n447), .A2(new_n449), .ZN(new_n1208));
  NAND2_X1  g1008(.A1(new_n431), .A2(new_n718), .ZN(new_n1209));
  XNOR2_X1  g1009(.A(new_n1208), .B(new_n1209), .ZN(new_n1210));
  XNOR2_X1  g1010(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1211));
  XNOR2_X1  g1011(.A(new_n1210), .B(new_n1211), .ZN(new_n1212));
  INV_X1    g1012(.A(new_n1212), .ZN(new_n1213));
  NAND2_X1  g1013(.A1(new_n1213), .A2(new_n812), .ZN(new_n1214));
  OAI22_X1  g1014(.A1(new_n877), .A2(new_n210), .B1(new_n879), .B2(new_n508), .ZN(new_n1215));
  NOR2_X1   g1015(.A1(new_n822), .A2(new_n256), .ZN(new_n1216));
  OR2_X1    g1016(.A1(new_n310), .A2(G41), .ZN(new_n1217));
  NOR4_X1   g1017(.A1(new_n1215), .A2(new_n1216), .A3(new_n1217), .A4(new_n1000), .ZN(new_n1218));
  NOR2_X1   g1018(.A1(new_n831), .A2(new_n457), .ZN(new_n1219));
  NOR2_X1   g1019(.A1(new_n828), .A2(new_n202), .ZN(new_n1220));
  AOI211_X1 g1020(.A(new_n1219), .B(new_n1220), .C1(G107), .C2(new_n884), .ZN(new_n1221));
  OAI211_X1 g1021(.A(new_n1218), .B(new_n1221), .C1(new_n878), .C2(new_n874), .ZN(new_n1222));
  INV_X1    g1022(.A(KEYINPUT58), .ZN(new_n1223));
  NOR2_X1   g1023(.A1(G33), .A2(G41), .ZN(new_n1224));
  NOR2_X1   g1024(.A1(new_n1224), .A2(G50), .ZN(new_n1225));
  AOI22_X1  g1025(.A1(new_n1222), .A2(new_n1223), .B1(new_n1217), .B2(new_n1225), .ZN(new_n1226));
  AOI22_X1  g1026(.A1(new_n871), .A2(G137), .B1(G132), .B2(new_n835), .ZN(new_n1227));
  XNOR2_X1  g1027(.A(new_n1227), .B(KEYINPUT121), .ZN(new_n1228));
  NOR2_X1   g1028(.A1(new_n879), .A2(new_n1187), .ZN(new_n1229));
  NOR2_X1   g1029(.A1(new_n842), .A2(new_n887), .ZN(new_n1230));
  OAI22_X1  g1030(.A1(new_n1197), .A2(new_n824), .B1(new_n822), .B2(new_n1194), .ZN(new_n1231));
  NOR4_X1   g1031(.A1(new_n1228), .A2(new_n1229), .A3(new_n1230), .A4(new_n1231), .ZN(new_n1232));
  INV_X1    g1032(.A(new_n1232), .ZN(new_n1233));
  NOR2_X1   g1033(.A1(new_n1233), .A2(KEYINPUT59), .ZN(new_n1234));
  OAI21_X1  g1034(.A(new_n1224), .B1(new_n828), .B2(new_n383), .ZN(new_n1235));
  AOI21_X1  g1035(.A(new_n1235), .B1(G124), .B2(new_n997), .ZN(new_n1236));
  INV_X1    g1036(.A(KEYINPUT59), .ZN(new_n1237));
  OAI21_X1  g1037(.A(new_n1236), .B1(new_n1232), .B2(new_n1237), .ZN(new_n1238));
  OAI221_X1 g1038(.A(new_n1226), .B1(new_n1223), .B2(new_n1222), .C1(new_n1234), .C2(new_n1238), .ZN(new_n1239));
  AND2_X1   g1039(.A1(new_n1239), .A2(new_n815), .ZN(new_n1240));
  AOI211_X1 g1040(.A(new_n863), .B(new_n1240), .C1(new_n201), .C2(new_n867), .ZN(new_n1241));
  NAND2_X1  g1041(.A1(new_n1214), .A2(new_n1241), .ZN(new_n1242));
  XOR2_X1   g1042(.A(new_n1242), .B(KEYINPUT122), .Z(new_n1243));
  AOI21_X1  g1043(.A(new_n1164), .B1(new_n914), .B2(new_n912), .ZN(new_n1244));
  AOI21_X1  g1044(.A(new_n935), .B1(new_n948), .B2(new_n949), .ZN(new_n1245));
  AOI21_X1  g1045(.A(new_n959), .B1(new_n1244), .B2(new_n1245), .ZN(new_n1246));
  AND3_X1   g1046(.A1(new_n1246), .A2(new_n936), .A3(new_n1212), .ZN(new_n1247));
  AOI21_X1  g1047(.A(new_n1212), .B1(new_n1246), .B2(new_n936), .ZN(new_n1248));
  OAI21_X1  g1048(.A(new_n983), .B1(new_n1247), .B2(new_n1248), .ZN(new_n1249));
  AOI21_X1  g1049(.A(KEYINPUT40), .B1(new_n974), .B2(new_n1244), .ZN(new_n1250));
  NAND2_X1  g1050(.A1(new_n951), .A2(G330), .ZN(new_n1251));
  OAI21_X1  g1051(.A(new_n1213), .B1(new_n1250), .B2(new_n1251), .ZN(new_n1252));
  AOI22_X1  g1052(.A1(new_n966), .A2(new_n968), .B1(new_n981), .B2(new_n719), .ZN(new_n1253));
  NAND3_X1  g1053(.A1(new_n1246), .A2(new_n936), .A3(new_n1212), .ZN(new_n1254));
  NAND4_X1  g1054(.A1(new_n1252), .A2(new_n980), .A3(new_n1253), .A4(new_n1254), .ZN(new_n1255));
  NAND2_X1  g1055(.A1(new_n1249), .A2(new_n1255), .ZN(new_n1256));
  AOI21_X1  g1056(.A(new_n1243), .B1(new_n802), .B2(new_n1256), .ZN(new_n1257));
  AOI22_X1  g1057(.A1(new_n1177), .A2(new_n1163), .B1(new_n1255), .B2(new_n1249), .ZN(new_n1258));
  OAI21_X1  g1058(.A(new_n739), .B1(new_n1258), .B2(KEYINPUT57), .ZN(new_n1259));
  NAND2_X1  g1059(.A1(new_n1177), .A2(new_n1163), .ZN(new_n1260));
  AND3_X1   g1060(.A1(new_n1260), .A2(KEYINPUT57), .A3(new_n1256), .ZN(new_n1261));
  OAI21_X1  g1061(.A(new_n1257), .B1(new_n1259), .B2(new_n1261), .ZN(G375));
  AOI21_X1  g1062(.A(new_n801), .B1(new_n1175), .B2(new_n1166), .ZN(new_n1263));
  NAND2_X1  g1063(.A1(new_n1143), .A2(new_n812), .ZN(new_n1264));
  OAI22_X1  g1064(.A1(new_n822), .A2(new_n383), .B1(new_n831), .B2(new_n887), .ZN(new_n1265));
  AOI21_X1  g1065(.A(new_n1265), .B1(G137), .B2(new_n884), .ZN(new_n1266));
  NAND2_X1  g1066(.A1(new_n840), .A2(G128), .ZN(new_n1267));
  NOR2_X1   g1067(.A1(new_n877), .A2(new_n1194), .ZN(new_n1268));
  NOR3_X1   g1068(.A1(new_n1268), .A2(new_n1220), .A3(new_n373), .ZN(new_n1269));
  AOI22_X1  g1069(.A1(new_n843), .A2(G50), .B1(G132), .B2(new_n844), .ZN(new_n1270));
  NAND4_X1  g1070(.A1(new_n1266), .A2(new_n1267), .A3(new_n1269), .A4(new_n1270), .ZN(new_n1271));
  OAI22_X1  g1071(.A1(new_n824), .A2(new_n878), .B1(new_n831), .B2(new_n497), .ZN(new_n1272));
  AOI21_X1  g1072(.A(new_n1272), .B1(G97), .B2(new_n852), .ZN(new_n1273));
  NAND2_X1  g1073(.A1(new_n840), .A2(G303), .ZN(new_n1274));
  AOI22_X1  g1074(.A1(G116), .A2(new_n835), .B1(new_n844), .B2(G294), .ZN(new_n1275));
  OAI21_X1  g1075(.A(new_n373), .B1(new_n828), .B2(new_n256), .ZN(new_n1276));
  AOI21_X1  g1076(.A(new_n1276), .B1(new_n458), .B2(new_n843), .ZN(new_n1277));
  NAND4_X1  g1077(.A1(new_n1273), .A2(new_n1274), .A3(new_n1275), .A4(new_n1277), .ZN(new_n1278));
  AOI21_X1  g1078(.A(new_n869), .B1(new_n1271), .B2(new_n1278), .ZN(new_n1279));
  AOI211_X1 g1079(.A(new_n863), .B(new_n1279), .C1(new_n203), .C2(new_n867), .ZN(new_n1280));
  AOI21_X1  g1080(.A(new_n1263), .B1(new_n1264), .B2(new_n1280), .ZN(new_n1281));
  NAND3_X1  g1081(.A1(new_n1175), .A2(new_n1162), .A3(new_n1166), .ZN(new_n1282));
  NAND3_X1  g1082(.A1(new_n1171), .A2(new_n1045), .A3(new_n1282), .ZN(new_n1283));
  NAND2_X1  g1083(.A1(new_n1281), .A2(new_n1283), .ZN(G381));
  INV_X1    g1084(.A(G384), .ZN(new_n1285));
  NAND2_X1  g1085(.A1(new_n1131), .A2(new_n1285), .ZN(new_n1286));
  NOR4_X1   g1086(.A1(new_n1286), .A2(G396), .A3(G393), .A4(G381), .ZN(new_n1287));
  AND2_X1   g1087(.A1(new_n1065), .A2(new_n1066), .ZN(new_n1288));
  AOI21_X1  g1088(.A(new_n1048), .B1(new_n1043), .B2(new_n1045), .ZN(new_n1289));
  AOI211_X1 g1089(.A(KEYINPUT113), .B(new_n1044), .C1(new_n1042), .C2(new_n798), .ZN(new_n1290));
  OAI21_X1  g1090(.A(new_n801), .B1(new_n1289), .B2(new_n1290), .ZN(new_n1291));
  NAND2_X1  g1091(.A1(new_n1288), .A2(new_n1291), .ZN(new_n1292));
  INV_X1    g1092(.A(G378), .ZN(new_n1293));
  NAND4_X1  g1093(.A1(new_n1287), .A2(new_n1292), .A3(new_n1023), .A4(new_n1293), .ZN(new_n1294));
  OR2_X1    g1094(.A1(new_n1294), .A2(G375), .ZN(G407));
  OAI21_X1  g1095(.A(G213), .B1(new_n1294), .B2(G375), .ZN(new_n1296));
  NAND2_X1  g1096(.A1(new_n720), .A2(G213), .ZN(new_n1297));
  NOR3_X1   g1097(.A1(G375), .A2(G378), .A3(new_n1297), .ZN(new_n1298));
  OR3_X1    g1098(.A1(new_n1296), .A2(KEYINPUT123), .A3(new_n1298), .ZN(new_n1299));
  OAI21_X1  g1099(.A(KEYINPUT123), .B1(new_n1296), .B2(new_n1298), .ZN(new_n1300));
  NAND2_X1  g1100(.A1(new_n1299), .A2(new_n1300), .ZN(G409));
  AOI221_X4 g1101(.A(new_n1044), .B1(new_n1255), .B2(new_n1249), .C1(new_n1177), .C2(new_n1163), .ZN(new_n1302));
  INV_X1    g1102(.A(new_n1242), .ZN(new_n1303));
  INV_X1    g1103(.A(KEYINPUT124), .ZN(new_n1304));
  AOI21_X1  g1104(.A(new_n801), .B1(new_n1256), .B2(new_n1304), .ZN(new_n1305));
  NAND3_X1  g1105(.A1(new_n1249), .A2(new_n1255), .A3(KEYINPUT124), .ZN(new_n1306));
  AOI21_X1  g1106(.A(new_n1303), .B1(new_n1305), .B2(new_n1306), .ZN(new_n1307));
  AOI21_X1  g1107(.A(new_n1302), .B1(new_n1307), .B2(KEYINPUT125), .ZN(new_n1308));
  NAND2_X1  g1108(.A1(new_n1256), .A2(new_n1304), .ZN(new_n1309));
  NAND3_X1  g1109(.A1(new_n1309), .A2(new_n802), .A3(new_n1306), .ZN(new_n1310));
  NAND2_X1  g1110(.A1(new_n1310), .A2(new_n1242), .ZN(new_n1311));
  INV_X1    g1111(.A(KEYINPUT125), .ZN(new_n1312));
  NAND2_X1  g1112(.A1(new_n1311), .A2(new_n1312), .ZN(new_n1313));
  AOI21_X1  g1113(.A(G378), .B1(new_n1308), .B2(new_n1313), .ZN(new_n1314));
  OAI211_X1 g1114(.A(G378), .B(new_n1257), .C1(new_n1259), .C2(new_n1261), .ZN(new_n1315));
  INV_X1    g1115(.A(new_n1315), .ZN(new_n1316));
  OAI21_X1  g1116(.A(new_n1297), .B1(new_n1314), .B2(new_n1316), .ZN(new_n1317));
  NAND3_X1  g1117(.A1(new_n720), .A2(G213), .A3(G2897), .ZN(new_n1318));
  INV_X1    g1118(.A(KEYINPUT60), .ZN(new_n1319));
  NAND2_X1  g1119(.A1(new_n1282), .A2(new_n1319), .ZN(new_n1320));
  NAND4_X1  g1120(.A1(new_n1175), .A2(new_n1162), .A3(new_n1166), .A4(KEYINPUT60), .ZN(new_n1321));
  NAND4_X1  g1121(.A1(new_n1320), .A2(new_n739), .A3(new_n1171), .A4(new_n1321), .ZN(new_n1322));
  AND3_X1   g1122(.A1(new_n1322), .A2(G384), .A3(new_n1281), .ZN(new_n1323));
  AOI21_X1  g1123(.A(G384), .B1(new_n1322), .B2(new_n1281), .ZN(new_n1324));
  NOR3_X1   g1124(.A1(new_n1323), .A2(new_n1324), .A3(KEYINPUT126), .ZN(new_n1325));
  INV_X1    g1125(.A(KEYINPUT126), .ZN(new_n1326));
  NAND2_X1  g1126(.A1(new_n1322), .A2(new_n1281), .ZN(new_n1327));
  NAND2_X1  g1127(.A1(new_n1327), .A2(new_n1285), .ZN(new_n1328));
  NAND3_X1  g1128(.A1(new_n1322), .A2(G384), .A3(new_n1281), .ZN(new_n1329));
  AOI21_X1  g1129(.A(new_n1326), .B1(new_n1328), .B2(new_n1329), .ZN(new_n1330));
  OAI21_X1  g1130(.A(new_n1318), .B1(new_n1325), .B2(new_n1330), .ZN(new_n1331));
  NAND3_X1  g1131(.A1(new_n1328), .A2(new_n1326), .A3(new_n1329), .ZN(new_n1332));
  INV_X1    g1132(.A(new_n1318), .ZN(new_n1333));
  NAND2_X1  g1133(.A1(new_n1332), .A2(new_n1333), .ZN(new_n1334));
  NAND3_X1  g1134(.A1(new_n1331), .A2(KEYINPUT127), .A3(new_n1334), .ZN(new_n1335));
  INV_X1    g1135(.A(KEYINPUT127), .ZN(new_n1336));
  OAI21_X1  g1136(.A(KEYINPUT126), .B1(new_n1323), .B2(new_n1324), .ZN(new_n1337));
  AOI21_X1  g1137(.A(new_n1333), .B1(new_n1337), .B2(new_n1332), .ZN(new_n1338));
  NOR2_X1   g1138(.A1(new_n1323), .A2(new_n1324), .ZN(new_n1339));
  AOI21_X1  g1139(.A(new_n1318), .B1(new_n1339), .B2(new_n1326), .ZN(new_n1340));
  OAI21_X1  g1140(.A(new_n1336), .B1(new_n1338), .B2(new_n1340), .ZN(new_n1341));
  NAND3_X1  g1141(.A1(new_n1317), .A2(new_n1335), .A3(new_n1341), .ZN(new_n1342));
  OAI211_X1 g1142(.A(new_n1297), .B(new_n1339), .C1(new_n1314), .C2(new_n1316), .ZN(new_n1343));
  NAND2_X1  g1143(.A1(new_n1343), .A2(KEYINPUT62), .ZN(new_n1344));
  INV_X1    g1144(.A(KEYINPUT61), .ZN(new_n1345));
  NAND3_X1  g1145(.A1(new_n1310), .A2(KEYINPUT125), .A3(new_n1242), .ZN(new_n1346));
  INV_X1    g1146(.A(new_n1302), .ZN(new_n1347));
  NAND2_X1  g1147(.A1(new_n1346), .A2(new_n1347), .ZN(new_n1348));
  NOR2_X1   g1148(.A1(new_n1307), .A2(KEYINPUT125), .ZN(new_n1349));
  OAI21_X1  g1149(.A(new_n1293), .B1(new_n1348), .B2(new_n1349), .ZN(new_n1350));
  NAND2_X1  g1150(.A1(new_n1350), .A2(new_n1315), .ZN(new_n1351));
  INV_X1    g1151(.A(KEYINPUT62), .ZN(new_n1352));
  NAND4_X1  g1152(.A1(new_n1351), .A2(new_n1352), .A3(new_n1297), .A4(new_n1339), .ZN(new_n1353));
  NAND4_X1  g1153(.A1(new_n1342), .A2(new_n1344), .A3(new_n1345), .A4(new_n1353), .ZN(new_n1354));
  XOR2_X1   g1154(.A(G393), .B(G396), .Z(new_n1355));
  INV_X1    g1155(.A(new_n1355), .ZN(new_n1356));
  AOI21_X1  g1156(.A(G390), .B1(new_n1292), .B2(new_n1023), .ZN(new_n1357));
  INV_X1    g1157(.A(new_n1023), .ZN(new_n1358));
  AOI211_X1 g1158(.A(new_n1358), .B(new_n1131), .C1(new_n1288), .C2(new_n1291), .ZN(new_n1359));
  OAI21_X1  g1159(.A(new_n1356), .B1(new_n1357), .B2(new_n1359), .ZN(new_n1360));
  NAND2_X1  g1160(.A1(G387), .A2(new_n1131), .ZN(new_n1361));
  NAND3_X1  g1161(.A1(new_n1292), .A2(new_n1023), .A3(G390), .ZN(new_n1362));
  NAND3_X1  g1162(.A1(new_n1361), .A2(new_n1355), .A3(new_n1362), .ZN(new_n1363));
  NAND2_X1  g1163(.A1(new_n1360), .A2(new_n1363), .ZN(new_n1364));
  NAND2_X1  g1164(.A1(new_n1354), .A2(new_n1364), .ZN(new_n1365));
  AOI21_X1  g1165(.A(KEYINPUT127), .B1(new_n1331), .B2(new_n1334), .ZN(new_n1366));
  NOR3_X1   g1166(.A1(new_n1338), .A2(new_n1340), .A3(new_n1336), .ZN(new_n1367));
  NOR2_X1   g1167(.A1(new_n1366), .A2(new_n1367), .ZN(new_n1368));
  AOI21_X1  g1168(.A(KEYINPUT61), .B1(new_n1368), .B2(new_n1317), .ZN(new_n1369));
  AND2_X1   g1169(.A1(new_n1360), .A2(new_n1363), .ZN(new_n1370));
  INV_X1    g1170(.A(KEYINPUT63), .ZN(new_n1371));
  OR2_X1    g1171(.A1(new_n1343), .A2(new_n1371), .ZN(new_n1372));
  NAND2_X1  g1172(.A1(new_n1343), .A2(new_n1371), .ZN(new_n1373));
  NAND4_X1  g1173(.A1(new_n1369), .A2(new_n1370), .A3(new_n1372), .A4(new_n1373), .ZN(new_n1374));
  NAND2_X1  g1174(.A1(new_n1365), .A2(new_n1374), .ZN(G405));
  AND2_X1   g1175(.A1(G375), .A2(new_n1293), .ZN(new_n1376));
  OAI21_X1  g1176(.A(new_n1339), .B1(new_n1376), .B2(new_n1316), .ZN(new_n1377));
  NAND2_X1  g1177(.A1(G375), .A2(new_n1293), .ZN(new_n1378));
  OAI211_X1 g1178(.A(new_n1378), .B(new_n1315), .C1(new_n1324), .C2(new_n1323), .ZN(new_n1379));
  NAND2_X1  g1179(.A1(new_n1377), .A2(new_n1379), .ZN(new_n1380));
  XNOR2_X1  g1180(.A(new_n1364), .B(new_n1380), .ZN(G402));
endmodule


