//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 0 0 0 0 0 1 1 1 0 0 0 0 0 1 1 0 0 1 1 0 1 0 1 1 0 1 1 1 0 1 0 1 1 0 1 0 1 1 1 0 1 1 1 0 1 0 1 1 0 0 0 1 1 0 1 0 0 0 1 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:38:32 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n205, new_n207, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n244, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n251, new_n252, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n692, new_n693, new_n694, new_n695, new_n696,
    new_n697, new_n698, new_n699, new_n700, new_n701, new_n702, new_n703,
    new_n704, new_n705, new_n706, new_n707, new_n708, new_n709, new_n710,
    new_n711, new_n712, new_n713, new_n714, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n772, new_n773, new_n774, new_n775,
    new_n776, new_n777, new_n778, new_n779, new_n780, new_n781, new_n782,
    new_n783, new_n784, new_n785, new_n786, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1087,
    new_n1088, new_n1089, new_n1090, new_n1091, new_n1092, new_n1093,
    new_n1094, new_n1095, new_n1096, new_n1097, new_n1098, new_n1099,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1108, new_n1109, new_n1110, new_n1111, new_n1112,
    new_n1113, new_n1114, new_n1115, new_n1116, new_n1117, new_n1118,
    new_n1119, new_n1120, new_n1121, new_n1122, new_n1123, new_n1124,
    new_n1125, new_n1126, new_n1127, new_n1128, new_n1129, new_n1130,
    new_n1131, new_n1132, new_n1133, new_n1134, new_n1135, new_n1136,
    new_n1137, new_n1138, new_n1139, new_n1140, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1186, new_n1187, new_n1188, new_n1189, new_n1190, new_n1191,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1251, new_n1252,
    new_n1253, new_n1255, new_n1256, new_n1257, new_n1258, new_n1259,
    new_n1260, new_n1261, new_n1262, new_n1263, new_n1264, new_n1265,
    new_n1266, new_n1267, new_n1268, new_n1269, new_n1270, new_n1271,
    new_n1272, new_n1273, new_n1274, new_n1275, new_n1277, new_n1278,
    new_n1279, new_n1281, new_n1282, new_n1283, new_n1284, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1344, new_n1345, new_n1346;
  INV_X1    g0000(.A(G58), .ZN(new_n201));
  INV_X1    g0001(.A(G68), .ZN(new_n202));
  NAND3_X1  g0002(.A1(new_n201), .A2(new_n202), .A3(KEYINPUT64), .ZN(new_n203));
  INV_X1    g0003(.A(KEYINPUT64), .ZN(new_n204));
  OAI21_X1  g0004(.A(new_n204), .B1(G58), .B2(G68), .ZN(new_n205));
  AOI211_X1 g0005(.A(G50), .B(G77), .C1(new_n203), .C2(new_n205), .ZN(G353));
  OAI21_X1  g0006(.A(G87), .B1(G97), .B2(G107), .ZN(new_n207));
  XOR2_X1   g0007(.A(new_n207), .B(KEYINPUT65), .Z(G355));
  NAND2_X1  g0008(.A1(G1), .A2(G20), .ZN(new_n209));
  OR3_X1    g0009(.A1(new_n209), .A2(KEYINPUT66), .A3(G13), .ZN(new_n210));
  OAI21_X1  g0010(.A(KEYINPUT66), .B1(new_n209), .B2(G13), .ZN(new_n211));
  NAND2_X1  g0011(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  INV_X1    g0012(.A(new_n212), .ZN(new_n213));
  OAI21_X1  g0013(.A(G250), .B1(G257), .B2(G264), .ZN(new_n214));
  NOR2_X1   g0014(.A1(new_n213), .A2(new_n214), .ZN(new_n215));
  NAND2_X1  g0015(.A1(G1), .A2(G13), .ZN(new_n216));
  INV_X1    g0016(.A(G20), .ZN(new_n217));
  NOR2_X1   g0017(.A1(new_n216), .A2(new_n217), .ZN(new_n218));
  NAND2_X1  g0018(.A1(new_n203), .A2(new_n205), .ZN(new_n219));
  INV_X1    g0019(.A(G50), .ZN(new_n220));
  NOR2_X1   g0020(.A1(new_n219), .A2(new_n220), .ZN(new_n221));
  AOI22_X1  g0021(.A1(new_n215), .A2(KEYINPUT0), .B1(new_n218), .B2(new_n221), .ZN(new_n222));
  AOI22_X1  g0022(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n223));
  INV_X1    g0023(.A(G238), .ZN(new_n224));
  INV_X1    g0024(.A(G77), .ZN(new_n225));
  INV_X1    g0025(.A(G244), .ZN(new_n226));
  OAI221_X1 g0026(.A(new_n223), .B1(new_n202), .B2(new_n224), .C1(new_n225), .C2(new_n226), .ZN(new_n227));
  XOR2_X1   g0027(.A(new_n227), .B(KEYINPUT67), .Z(new_n228));
  AOI22_X1  g0028(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n229));
  XOR2_X1   g0029(.A(new_n229), .B(KEYINPUT68), .Z(new_n230));
  AOI22_X1  g0030(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n231));
  NAND2_X1  g0031(.A1(new_n230), .A2(new_n231), .ZN(new_n232));
  OAI21_X1  g0032(.A(new_n209), .B1(new_n228), .B2(new_n232), .ZN(new_n233));
  OAI221_X1 g0033(.A(new_n222), .B1(KEYINPUT0), .B2(new_n215), .C1(new_n233), .C2(KEYINPUT1), .ZN(new_n234));
  AOI21_X1  g0034(.A(new_n234), .B1(KEYINPUT1), .B2(new_n233), .ZN(new_n235));
  XOR2_X1   g0035(.A(new_n235), .B(KEYINPUT69), .Z(G361));
  XNOR2_X1  g0036(.A(G238), .B(G244), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n237), .B(G232), .ZN(new_n238));
  XNOR2_X1  g0038(.A(KEYINPUT2), .B(G226), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XNOR2_X1  g0040(.A(G250), .B(G257), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n241), .B(KEYINPUT70), .ZN(new_n242));
  XNOR2_X1  g0042(.A(G264), .B(G270), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n240), .B(new_n244), .ZN(G358));
  XNOR2_X1  g0045(.A(G87), .B(G97), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n246), .B(KEYINPUT71), .ZN(new_n247));
  XNOR2_X1  g0047(.A(G107), .B(G116), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n247), .B(new_n248), .ZN(new_n249));
  XNOR2_X1  g0049(.A(G50), .B(G68), .ZN(new_n250));
  XNOR2_X1  g0050(.A(G58), .B(G77), .ZN(new_n251));
  XNOR2_X1  g0051(.A(new_n250), .B(new_n251), .ZN(new_n252));
  XNOR2_X1  g0052(.A(new_n249), .B(new_n252), .ZN(G351));
  INV_X1    g0053(.A(G1), .ZN(new_n254));
  OAI21_X1  g0054(.A(new_n254), .B1(G41), .B2(G45), .ZN(new_n255));
  INV_X1    g0055(.A(KEYINPUT72), .ZN(new_n256));
  NAND2_X1  g0056(.A1(new_n255), .A2(new_n256), .ZN(new_n257));
  OAI211_X1 g0057(.A(new_n254), .B(KEYINPUT72), .C1(G41), .C2(G45), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n257), .A2(new_n258), .ZN(new_n259));
  INV_X1    g0059(.A(G274), .ZN(new_n260));
  AND2_X1   g0060(.A1(G1), .A2(G13), .ZN(new_n261));
  NAND2_X1  g0061(.A1(G33), .A2(G41), .ZN(new_n262));
  AOI21_X1  g0062(.A(new_n260), .B1(new_n261), .B2(new_n262), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n259), .A2(new_n263), .ZN(new_n264));
  NOR2_X1   g0064(.A1(G226), .A2(G1698), .ZN(new_n265));
  INV_X1    g0065(.A(G232), .ZN(new_n266));
  AOI21_X1  g0066(.A(new_n265), .B1(new_n266), .B2(G1698), .ZN(new_n267));
  XNOR2_X1  g0067(.A(KEYINPUT3), .B(G33), .ZN(new_n268));
  AOI22_X1  g0068(.A1(new_n267), .A2(new_n268), .B1(G33), .B2(G97), .ZN(new_n269));
  NAND3_X1  g0069(.A1(new_n262), .A2(G1), .A3(G13), .ZN(new_n270));
  OAI21_X1  g0070(.A(new_n264), .B1(new_n269), .B2(new_n270), .ZN(new_n271));
  AOI21_X1  g0071(.A(KEYINPUT73), .B1(new_n270), .B2(new_n255), .ZN(new_n272));
  INV_X1    g0072(.A(new_n272), .ZN(new_n273));
  NAND3_X1  g0073(.A1(new_n270), .A2(KEYINPUT73), .A3(new_n255), .ZN(new_n274));
  AOI21_X1  g0074(.A(new_n224), .B1(new_n273), .B2(new_n274), .ZN(new_n275));
  NOR3_X1   g0075(.A1(new_n271), .A2(new_n275), .A3(KEYINPUT13), .ZN(new_n276));
  INV_X1    g0076(.A(KEYINPUT13), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n266), .A2(G1698), .ZN(new_n278));
  OAI21_X1  g0078(.A(new_n278), .B1(G226), .B2(G1698), .ZN(new_n279));
  AND2_X1   g0079(.A1(KEYINPUT3), .A2(G33), .ZN(new_n280));
  NOR2_X1   g0080(.A1(KEYINPUT3), .A2(G33), .ZN(new_n281));
  NOR2_X1   g0081(.A1(new_n280), .A2(new_n281), .ZN(new_n282));
  INV_X1    g0082(.A(G33), .ZN(new_n283));
  INV_X1    g0083(.A(G97), .ZN(new_n284));
  OAI22_X1  g0084(.A1(new_n279), .A2(new_n282), .B1(new_n283), .B2(new_n284), .ZN(new_n285));
  AOI21_X1  g0085(.A(new_n216), .B1(G33), .B2(G41), .ZN(new_n286));
  AOI22_X1  g0086(.A1(new_n285), .A2(new_n286), .B1(new_n259), .B2(new_n263), .ZN(new_n287));
  INV_X1    g0087(.A(new_n274), .ZN(new_n288));
  OAI21_X1  g0088(.A(G238), .B1(new_n288), .B2(new_n272), .ZN(new_n289));
  AOI21_X1  g0089(.A(new_n277), .B1(new_n287), .B2(new_n289), .ZN(new_n290));
  NOR2_X1   g0090(.A1(new_n276), .A2(new_n290), .ZN(new_n291));
  NAND3_X1  g0091(.A1(new_n291), .A2(KEYINPUT74), .A3(G190), .ZN(new_n292));
  INV_X1    g0092(.A(KEYINPUT74), .ZN(new_n293));
  OAI21_X1  g0093(.A(KEYINPUT13), .B1(new_n271), .B2(new_n275), .ZN(new_n294));
  NAND3_X1  g0094(.A1(new_n287), .A2(new_n289), .A3(new_n277), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n294), .A2(new_n295), .ZN(new_n296));
  INV_X1    g0096(.A(G190), .ZN(new_n297));
  OAI21_X1  g0097(.A(new_n293), .B1(new_n296), .B2(new_n297), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n292), .A2(new_n298), .ZN(new_n299));
  NAND3_X1  g0099(.A1(new_n254), .A2(G13), .A3(G20), .ZN(new_n300));
  INV_X1    g0100(.A(new_n300), .ZN(new_n301));
  NAND3_X1  g0101(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n302), .A2(new_n216), .ZN(new_n303));
  NOR2_X1   g0103(.A1(new_n301), .A2(new_n303), .ZN(new_n304));
  AOI21_X1  g0104(.A(new_n202), .B1(new_n254), .B2(G20), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n304), .A2(new_n305), .ZN(new_n306));
  INV_X1    g0106(.A(KEYINPUT75), .ZN(new_n307));
  XNOR2_X1  g0107(.A(new_n306), .B(new_n307), .ZN(new_n308));
  NOR2_X1   g0108(.A1(G20), .A2(G33), .ZN(new_n309));
  AOI22_X1  g0109(.A1(new_n309), .A2(G50), .B1(G20), .B2(new_n202), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n217), .A2(G33), .ZN(new_n311));
  OAI21_X1  g0111(.A(new_n310), .B1(new_n225), .B2(new_n311), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n312), .A2(new_n303), .ZN(new_n313));
  INV_X1    g0113(.A(KEYINPUT11), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n313), .A2(new_n314), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n301), .A2(new_n202), .ZN(new_n316));
  XNOR2_X1  g0116(.A(new_n316), .B(KEYINPUT12), .ZN(new_n317));
  NAND3_X1  g0117(.A1(new_n312), .A2(KEYINPUT11), .A3(new_n303), .ZN(new_n318));
  NAND4_X1  g0118(.A1(new_n308), .A2(new_n315), .A3(new_n317), .A4(new_n318), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n319), .A2(KEYINPUT76), .ZN(new_n320));
  AND2_X1   g0120(.A1(new_n317), .A2(new_n318), .ZN(new_n321));
  INV_X1    g0121(.A(KEYINPUT76), .ZN(new_n322));
  NAND4_X1  g0122(.A1(new_n321), .A2(new_n322), .A3(new_n308), .A4(new_n315), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n320), .A2(new_n323), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n296), .A2(G200), .ZN(new_n325));
  NAND3_X1  g0125(.A1(new_n299), .A2(new_n324), .A3(new_n325), .ZN(new_n326));
  INV_X1    g0126(.A(G169), .ZN(new_n327));
  AOI21_X1  g0127(.A(new_n327), .B1(new_n294), .B2(new_n295), .ZN(new_n328));
  INV_X1    g0128(.A(KEYINPUT14), .ZN(new_n329));
  INV_X1    g0129(.A(G179), .ZN(new_n330));
  OAI22_X1  g0130(.A1(new_n328), .A2(new_n329), .B1(new_n296), .B2(new_n330), .ZN(new_n331));
  INV_X1    g0131(.A(KEYINPUT77), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n296), .A2(G169), .ZN(new_n333));
  OAI21_X1  g0133(.A(new_n332), .B1(new_n333), .B2(KEYINPUT14), .ZN(new_n334));
  NAND3_X1  g0134(.A1(new_n328), .A2(KEYINPUT77), .A3(new_n329), .ZN(new_n335));
  AOI21_X1  g0135(.A(new_n331), .B1(new_n334), .B2(new_n335), .ZN(new_n336));
  OAI21_X1  g0136(.A(new_n326), .B1(new_n336), .B2(new_n324), .ZN(new_n337));
  NAND2_X1  g0137(.A1(G20), .A2(G77), .ZN(new_n338));
  XNOR2_X1  g0138(.A(KEYINPUT8), .B(G58), .ZN(new_n339));
  INV_X1    g0139(.A(new_n309), .ZN(new_n340));
  XNOR2_X1  g0140(.A(KEYINPUT15), .B(G87), .ZN(new_n341));
  OAI221_X1 g0141(.A(new_n338), .B1(new_n339), .B2(new_n340), .C1(new_n311), .C2(new_n341), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n342), .A2(new_n303), .ZN(new_n343));
  AOI21_X1  g0143(.A(new_n225), .B1(new_n254), .B2(G20), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n304), .A2(new_n344), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n301), .A2(new_n225), .ZN(new_n346));
  AND2_X1   g0146(.A1(new_n345), .A2(new_n346), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n343), .A2(new_n347), .ZN(new_n348));
  INV_X1    g0148(.A(G1698), .ZN(new_n349));
  NAND3_X1  g0149(.A1(new_n268), .A2(G232), .A3(new_n349), .ZN(new_n350));
  NAND3_X1  g0150(.A1(new_n268), .A2(G238), .A3(G1698), .ZN(new_n351));
  INV_X1    g0151(.A(G107), .ZN(new_n352));
  OAI211_X1 g0152(.A(new_n350), .B(new_n351), .C1(new_n352), .C2(new_n268), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n353), .A2(new_n286), .ZN(new_n354));
  OAI21_X1  g0154(.A(G244), .B1(new_n288), .B2(new_n272), .ZN(new_n355));
  NAND3_X1  g0155(.A1(new_n354), .A2(new_n264), .A3(new_n355), .ZN(new_n356));
  AOI21_X1  g0156(.A(new_n348), .B1(new_n356), .B2(G200), .ZN(new_n357));
  OAI21_X1  g0157(.A(new_n357), .B1(new_n297), .B2(new_n356), .ZN(new_n358));
  AOI22_X1  g0158(.A1(new_n356), .A2(new_n327), .B1(new_n343), .B2(new_n347), .ZN(new_n359));
  NAND4_X1  g0159(.A1(new_n354), .A2(new_n330), .A3(new_n264), .A4(new_n355), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n359), .A2(new_n360), .ZN(new_n361));
  AND2_X1   g0161(.A1(new_n358), .A2(new_n361), .ZN(new_n362));
  NAND3_X1  g0162(.A1(new_n268), .A2(G222), .A3(new_n349), .ZN(new_n363));
  NAND3_X1  g0163(.A1(new_n268), .A2(G223), .A3(G1698), .ZN(new_n364));
  OAI211_X1 g0164(.A(new_n363), .B(new_n364), .C1(new_n225), .C2(new_n268), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n365), .A2(new_n286), .ZN(new_n366));
  OAI21_X1  g0166(.A(G226), .B1(new_n288), .B2(new_n272), .ZN(new_n367));
  NAND3_X1  g0167(.A1(new_n366), .A2(new_n264), .A3(new_n367), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n368), .A2(new_n327), .ZN(new_n369));
  AOI21_X1  g0169(.A(new_n217), .B1(new_n219), .B2(new_n220), .ZN(new_n370));
  INV_X1    g0170(.A(G150), .ZN(new_n371));
  OAI22_X1  g0171(.A1(new_n339), .A2(new_n311), .B1(new_n371), .B2(new_n340), .ZN(new_n372));
  OAI21_X1  g0172(.A(new_n303), .B1(new_n370), .B2(new_n372), .ZN(new_n373));
  AOI21_X1  g0173(.A(new_n220), .B1(new_n254), .B2(G20), .ZN(new_n374));
  AOI22_X1  g0174(.A1(new_n304), .A2(new_n374), .B1(new_n220), .B2(new_n301), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n373), .A2(new_n375), .ZN(new_n376));
  OAI211_X1 g0176(.A(new_n369), .B(new_n376), .C1(G179), .C2(new_n368), .ZN(new_n377));
  INV_X1    g0177(.A(KEYINPUT10), .ZN(new_n378));
  INV_X1    g0178(.A(KEYINPUT9), .ZN(new_n379));
  NOR2_X1   g0179(.A1(new_n376), .A2(new_n379), .ZN(new_n380));
  INV_X1    g0180(.A(new_n368), .ZN(new_n381));
  AOI21_X1  g0181(.A(new_n380), .B1(new_n381), .B2(G190), .ZN(new_n382));
  AOI22_X1  g0182(.A1(new_n368), .A2(G200), .B1(new_n379), .B2(new_n376), .ZN(new_n383));
  AOI21_X1  g0183(.A(new_n378), .B1(new_n382), .B2(new_n383), .ZN(new_n384));
  NAND2_X1  g0184(.A1(new_n376), .A2(new_n379), .ZN(new_n385));
  INV_X1    g0185(.A(G200), .ZN(new_n386));
  OAI21_X1  g0186(.A(new_n385), .B1(new_n381), .B2(new_n386), .ZN(new_n387));
  OAI22_X1  g0187(.A1(new_n368), .A2(new_n297), .B1(new_n379), .B2(new_n376), .ZN(new_n388));
  NOR3_X1   g0188(.A1(new_n387), .A2(new_n388), .A3(KEYINPUT10), .ZN(new_n389));
  OAI211_X1 g0189(.A(new_n362), .B(new_n377), .C1(new_n384), .C2(new_n389), .ZN(new_n390));
  INV_X1    g0190(.A(KEYINPUT17), .ZN(new_n391));
  AOI21_X1  g0191(.A(new_n339), .B1(new_n254), .B2(G20), .ZN(new_n392));
  AOI22_X1  g0192(.A1(new_n392), .A2(new_n304), .B1(new_n301), .B2(new_n339), .ZN(new_n393));
  NAND2_X1  g0193(.A1(G58), .A2(G68), .ZN(new_n394));
  NAND3_X1  g0194(.A1(new_n203), .A2(new_n205), .A3(new_n394), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n395), .A2(G20), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n309), .A2(G159), .ZN(new_n397));
  NAND2_X1  g0197(.A1(new_n396), .A2(new_n397), .ZN(new_n398));
  AOI21_X1  g0198(.A(KEYINPUT7), .B1(new_n282), .B2(new_n217), .ZN(new_n399));
  INV_X1    g0199(.A(KEYINPUT3), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n400), .A2(new_n283), .ZN(new_n401));
  NAND2_X1  g0201(.A1(KEYINPUT3), .A2(G33), .ZN(new_n402));
  NAND4_X1  g0202(.A1(new_n401), .A2(KEYINPUT7), .A3(new_n217), .A4(new_n402), .ZN(new_n403));
  INV_X1    g0203(.A(new_n403), .ZN(new_n404));
  OAI21_X1  g0204(.A(G68), .B1(new_n399), .B2(new_n404), .ZN(new_n405));
  INV_X1    g0205(.A(KEYINPUT79), .ZN(new_n406));
  AOI21_X1  g0206(.A(new_n398), .B1(new_n405), .B2(new_n406), .ZN(new_n407));
  NAND3_X1  g0207(.A1(new_n401), .A2(new_n217), .A3(new_n402), .ZN(new_n408));
  INV_X1    g0208(.A(KEYINPUT7), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n408), .A2(new_n409), .ZN(new_n410));
  AOI211_X1 g0210(.A(new_n406), .B(new_n202), .C1(new_n410), .C2(new_n403), .ZN(new_n411));
  INV_X1    g0211(.A(new_n411), .ZN(new_n412));
  AOI21_X1  g0212(.A(KEYINPUT16), .B1(new_n407), .B2(new_n412), .ZN(new_n413));
  AOI22_X1  g0213(.A1(new_n395), .A2(G20), .B1(G159), .B2(new_n309), .ZN(new_n414));
  INV_X1    g0214(.A(KEYINPUT78), .ZN(new_n415));
  AND3_X1   g0215(.A1(new_n410), .A2(new_n415), .A3(new_n403), .ZN(new_n416));
  NOR2_X1   g0216(.A1(new_n415), .A2(KEYINPUT7), .ZN(new_n417));
  NAND3_X1  g0217(.A1(new_n408), .A2(new_n409), .A3(new_n417), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n418), .A2(G68), .ZN(new_n419));
  OAI211_X1 g0219(.A(KEYINPUT16), .B(new_n414), .C1(new_n416), .C2(new_n419), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n420), .A2(new_n303), .ZN(new_n421));
  OAI21_X1  g0221(.A(new_n393), .B1(new_n413), .B2(new_n421), .ZN(new_n422));
  OAI211_X1 g0222(.A(G223), .B(new_n349), .C1(new_n280), .C2(new_n281), .ZN(new_n423));
  OAI211_X1 g0223(.A(G226), .B(G1698), .C1(new_n280), .C2(new_n281), .ZN(new_n424));
  AND3_X1   g0224(.A1(KEYINPUT80), .A2(G33), .A3(G87), .ZN(new_n425));
  AOI21_X1  g0225(.A(KEYINPUT80), .B1(G33), .B2(G87), .ZN(new_n426));
  NOR2_X1   g0226(.A1(new_n425), .A2(new_n426), .ZN(new_n427));
  NAND3_X1  g0227(.A1(new_n423), .A2(new_n424), .A3(new_n427), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n428), .A2(new_n286), .ZN(new_n429));
  INV_X1    g0229(.A(G41), .ZN(new_n430));
  INV_X1    g0230(.A(G45), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n430), .A2(new_n431), .ZN(new_n432));
  AOI22_X1  g0232(.A1(new_n254), .A2(new_n432), .B1(new_n261), .B2(new_n262), .ZN(new_n433));
  AOI22_X1  g0233(.A1(new_n259), .A2(new_n263), .B1(new_n433), .B2(G232), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n429), .A2(new_n434), .ZN(new_n435));
  NOR2_X1   g0235(.A1(new_n435), .A2(G190), .ZN(new_n436));
  INV_X1    g0236(.A(KEYINPUT81), .ZN(new_n437));
  NAND2_X1  g0237(.A1(new_n435), .A2(new_n437), .ZN(new_n438));
  NAND3_X1  g0238(.A1(new_n429), .A2(new_n434), .A3(KEYINPUT81), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n438), .A2(new_n439), .ZN(new_n440));
  AOI21_X1  g0240(.A(new_n436), .B1(new_n440), .B2(new_n386), .ZN(new_n441));
  OAI21_X1  g0241(.A(new_n391), .B1(new_n422), .B2(new_n441), .ZN(new_n442));
  INV_X1    g0242(.A(new_n393), .ZN(new_n443));
  INV_X1    g0243(.A(new_n303), .ZN(new_n444));
  AOI21_X1  g0244(.A(new_n202), .B1(new_n399), .B2(new_n417), .ZN(new_n445));
  NAND3_X1  g0245(.A1(new_n410), .A2(new_n415), .A3(new_n403), .ZN(new_n446));
  AOI21_X1  g0246(.A(new_n398), .B1(new_n445), .B2(new_n446), .ZN(new_n447));
  AOI21_X1  g0247(.A(new_n444), .B1(new_n447), .B2(KEYINPUT16), .ZN(new_n448));
  INV_X1    g0248(.A(KEYINPUT16), .ZN(new_n449));
  AOI21_X1  g0249(.A(new_n202), .B1(new_n410), .B2(new_n403), .ZN(new_n450));
  OAI21_X1  g0250(.A(new_n414), .B1(new_n450), .B2(KEYINPUT79), .ZN(new_n451));
  OAI21_X1  g0251(.A(new_n449), .B1(new_n451), .B2(new_n411), .ZN(new_n452));
  AOI21_X1  g0252(.A(new_n443), .B1(new_n448), .B2(new_n452), .ZN(new_n453));
  AND3_X1   g0253(.A1(new_n429), .A2(new_n434), .A3(KEYINPUT81), .ZN(new_n454));
  AOI21_X1  g0254(.A(KEYINPUT81), .B1(new_n429), .B2(new_n434), .ZN(new_n455));
  OAI21_X1  g0255(.A(new_n327), .B1(new_n454), .B2(new_n455), .ZN(new_n456));
  NOR2_X1   g0256(.A1(new_n435), .A2(G179), .ZN(new_n457));
  INV_X1    g0257(.A(new_n457), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n456), .A2(new_n458), .ZN(new_n459));
  OAI21_X1  g0259(.A(KEYINPUT18), .B1(new_n453), .B2(new_n459), .ZN(new_n460));
  AOI21_X1  g0260(.A(new_n457), .B1(new_n440), .B2(new_n327), .ZN(new_n461));
  INV_X1    g0261(.A(KEYINPUT18), .ZN(new_n462));
  NAND3_X1  g0262(.A1(new_n422), .A2(new_n461), .A3(new_n462), .ZN(new_n463));
  OAI21_X1  g0263(.A(new_n386), .B1(new_n454), .B2(new_n455), .ZN(new_n464));
  INV_X1    g0264(.A(new_n436), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  NAND3_X1  g0266(.A1(new_n453), .A2(new_n466), .A3(KEYINPUT17), .ZN(new_n467));
  NAND4_X1  g0267(.A1(new_n442), .A2(new_n460), .A3(new_n463), .A4(new_n467), .ZN(new_n468));
  NOR3_X1   g0268(.A1(new_n337), .A2(new_n390), .A3(new_n468), .ZN(new_n469));
  INV_X1    g0269(.A(G116), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n301), .A2(new_n470), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n254), .A2(G33), .ZN(new_n472));
  NAND4_X1  g0272(.A1(new_n300), .A2(new_n472), .A3(new_n216), .A4(new_n302), .ZN(new_n473));
  OAI21_X1  g0273(.A(new_n471), .B1(new_n473), .B2(new_n470), .ZN(new_n474));
  INV_X1    g0274(.A(new_n474), .ZN(new_n475));
  NAND2_X1  g0275(.A1(G33), .A2(G283), .ZN(new_n476));
  AND2_X1   g0276(.A1(KEYINPUT83), .A2(G97), .ZN(new_n477));
  NOR2_X1   g0277(.A1(KEYINPUT83), .A2(G97), .ZN(new_n478));
  NOR2_X1   g0278(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  OAI211_X1 g0279(.A(new_n217), .B(new_n476), .C1(new_n479), .C2(G33), .ZN(new_n480));
  AOI22_X1  g0280(.A1(new_n302), .A2(new_n216), .B1(G20), .B2(new_n470), .ZN(new_n481));
  AOI21_X1  g0281(.A(KEYINPUT20), .B1(new_n480), .B2(new_n481), .ZN(new_n482));
  INV_X1    g0282(.A(KEYINPUT83), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n483), .A2(new_n284), .ZN(new_n484));
  NAND2_X1  g0284(.A1(KEYINPUT83), .A2(G97), .ZN(new_n485));
  AOI21_X1  g0285(.A(G33), .B1(new_n484), .B2(new_n485), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n476), .A2(new_n217), .ZN(new_n487));
  OAI211_X1 g0287(.A(KEYINPUT20), .B(new_n481), .C1(new_n486), .C2(new_n487), .ZN(new_n488));
  INV_X1    g0288(.A(new_n488), .ZN(new_n489));
  OAI21_X1  g0289(.A(new_n475), .B1(new_n482), .B2(new_n489), .ZN(new_n490));
  NOR2_X1   g0290(.A1(new_n431), .A2(G1), .ZN(new_n491));
  AND2_X1   g0291(.A1(KEYINPUT5), .A2(G41), .ZN(new_n492));
  NOR2_X1   g0292(.A1(KEYINPUT5), .A2(G41), .ZN(new_n493));
  OAI21_X1  g0293(.A(new_n491), .B1(new_n492), .B2(new_n493), .ZN(new_n494));
  NAND3_X1  g0294(.A1(new_n494), .A2(G270), .A3(new_n270), .ZN(new_n495));
  XNOR2_X1  g0295(.A(KEYINPUT5), .B(G41), .ZN(new_n496));
  NAND3_X1  g0296(.A1(new_n263), .A2(new_n491), .A3(new_n496), .ZN(new_n497));
  AND2_X1   g0297(.A1(new_n495), .A2(new_n497), .ZN(new_n498));
  OAI211_X1 g0298(.A(G264), .B(G1698), .C1(new_n280), .C2(new_n281), .ZN(new_n499));
  OAI211_X1 g0299(.A(G257), .B(new_n349), .C1(new_n280), .C2(new_n281), .ZN(new_n500));
  NAND3_X1  g0300(.A1(new_n401), .A2(G303), .A3(new_n402), .ZN(new_n501));
  NAND3_X1  g0301(.A1(new_n499), .A2(new_n500), .A3(new_n501), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n502), .A2(new_n286), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n498), .A2(new_n503), .ZN(new_n504));
  AOI21_X1  g0304(.A(new_n490), .B1(G200), .B2(new_n504), .ZN(new_n505));
  OAI21_X1  g0305(.A(new_n505), .B1(new_n297), .B2(new_n504), .ZN(new_n506));
  AOI21_X1  g0306(.A(new_n327), .B1(new_n498), .B2(new_n503), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n507), .A2(KEYINPUT21), .ZN(new_n508));
  NAND3_X1  g0308(.A1(new_n498), .A2(G179), .A3(new_n503), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n510), .A2(new_n490), .ZN(new_n511));
  INV_X1    g0311(.A(KEYINPUT88), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n507), .A2(new_n490), .ZN(new_n513));
  INV_X1    g0313(.A(KEYINPUT21), .ZN(new_n514));
  AOI21_X1  g0314(.A(new_n512), .B1(new_n513), .B2(new_n514), .ZN(new_n515));
  AOI211_X1 g0315(.A(KEYINPUT88), .B(KEYINPUT21), .C1(new_n507), .C2(new_n490), .ZN(new_n516));
  OAI211_X1 g0316(.A(new_n506), .B(new_n511), .C1(new_n515), .C2(new_n516), .ZN(new_n517));
  INV_X1    g0317(.A(new_n517), .ZN(new_n518));
  OAI211_X1 g0318(.A(new_n217), .B(G87), .C1(new_n280), .C2(new_n281), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n519), .A2(KEYINPUT22), .ZN(new_n520));
  INV_X1    g0320(.A(KEYINPUT22), .ZN(new_n521));
  NAND4_X1  g0321(.A1(new_n268), .A2(new_n521), .A3(new_n217), .A4(G87), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n520), .A2(new_n522), .ZN(new_n523));
  NOR3_X1   g0323(.A1(new_n283), .A2(new_n470), .A3(G20), .ZN(new_n524));
  INV_X1    g0324(.A(KEYINPUT23), .ZN(new_n525));
  OAI21_X1  g0325(.A(new_n525), .B1(new_n217), .B2(G107), .ZN(new_n526));
  NAND3_X1  g0326(.A1(new_n352), .A2(KEYINPUT23), .A3(G20), .ZN(new_n527));
  AOI21_X1  g0327(.A(new_n524), .B1(new_n526), .B2(new_n527), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n523), .A2(new_n528), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n529), .A2(KEYINPUT24), .ZN(new_n530));
  INV_X1    g0330(.A(KEYINPUT24), .ZN(new_n531));
  NAND3_X1  g0331(.A1(new_n523), .A2(new_n531), .A3(new_n528), .ZN(new_n532));
  AOI21_X1  g0332(.A(new_n444), .B1(new_n530), .B2(new_n532), .ZN(new_n533));
  XOR2_X1   g0333(.A(KEYINPUT89), .B(KEYINPUT25), .Z(new_n534));
  NOR2_X1   g0334(.A1(new_n300), .A2(G107), .ZN(new_n535));
  XNOR2_X1  g0335(.A(new_n534), .B(new_n535), .ZN(new_n536));
  NOR2_X1   g0336(.A1(new_n473), .A2(new_n352), .ZN(new_n537));
  NOR2_X1   g0337(.A1(new_n536), .A2(new_n537), .ZN(new_n538));
  INV_X1    g0338(.A(new_n538), .ZN(new_n539));
  OAI21_X1  g0339(.A(KEYINPUT90), .B1(new_n533), .B2(new_n539), .ZN(new_n540));
  INV_X1    g0340(.A(new_n532), .ZN(new_n541));
  AOI21_X1  g0341(.A(new_n531), .B1(new_n523), .B2(new_n528), .ZN(new_n542));
  OAI21_X1  g0342(.A(new_n303), .B1(new_n541), .B2(new_n542), .ZN(new_n543));
  INV_X1    g0343(.A(KEYINPUT90), .ZN(new_n544));
  NAND3_X1  g0344(.A1(new_n543), .A2(new_n544), .A3(new_n538), .ZN(new_n545));
  OAI211_X1 g0345(.A(G257), .B(G1698), .C1(new_n280), .C2(new_n281), .ZN(new_n546));
  OAI211_X1 g0346(.A(G250), .B(new_n349), .C1(new_n280), .C2(new_n281), .ZN(new_n547));
  INV_X1    g0347(.A(G294), .ZN(new_n548));
  OAI211_X1 g0348(.A(new_n546), .B(new_n547), .C1(new_n283), .C2(new_n548), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n549), .A2(new_n286), .ZN(new_n550));
  AOI21_X1  g0350(.A(new_n286), .B1(new_n491), .B2(new_n496), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n551), .A2(G264), .ZN(new_n552));
  NAND3_X1  g0352(.A1(new_n550), .A2(new_n497), .A3(new_n552), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n553), .A2(G169), .ZN(new_n554));
  AOI22_X1  g0354(.A1(new_n549), .A2(new_n286), .B1(new_n551), .B2(G264), .ZN(new_n555));
  NAND3_X1  g0355(.A1(new_n555), .A2(G179), .A3(new_n497), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n554), .A2(new_n556), .ZN(new_n557));
  NAND3_X1  g0357(.A1(new_n540), .A2(new_n545), .A3(new_n557), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n553), .A2(G200), .ZN(new_n559));
  NAND3_X1  g0359(.A1(new_n555), .A2(G190), .A3(new_n497), .ZN(new_n560));
  NAND4_X1  g0360(.A1(new_n543), .A2(new_n538), .A3(new_n559), .A4(new_n560), .ZN(new_n561));
  AND2_X1   g0361(.A1(new_n558), .A2(new_n561), .ZN(new_n562));
  OAI211_X1 g0362(.A(G244), .B(new_n349), .C1(new_n280), .C2(new_n281), .ZN(new_n563));
  INV_X1    g0363(.A(KEYINPUT4), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n563), .A2(new_n564), .ZN(new_n565));
  INV_X1    g0365(.A(new_n476), .ZN(new_n566));
  NAND2_X1  g0366(.A1(G250), .A2(G1698), .ZN(new_n567));
  NAND2_X1  g0367(.A1(KEYINPUT4), .A2(G244), .ZN(new_n568));
  OAI21_X1  g0368(.A(new_n567), .B1(new_n568), .B2(G1698), .ZN(new_n569));
  AOI21_X1  g0369(.A(new_n566), .B1(new_n268), .B2(new_n569), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n565), .A2(new_n570), .ZN(new_n571));
  INV_X1    g0371(.A(KEYINPUT85), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n571), .A2(new_n572), .ZN(new_n573));
  NAND3_X1  g0373(.A1(new_n565), .A2(new_n570), .A3(KEYINPUT85), .ZN(new_n574));
  AOI21_X1  g0374(.A(new_n270), .B1(new_n573), .B2(new_n574), .ZN(new_n575));
  INV_X1    g0375(.A(KEYINPUT86), .ZN(new_n576));
  AOI21_X1  g0376(.A(new_n576), .B1(new_n551), .B2(G257), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n494), .A2(new_n270), .ZN(new_n578));
  INV_X1    g0378(.A(G257), .ZN(new_n579));
  NOR3_X1   g0379(.A1(new_n578), .A2(KEYINPUT86), .A3(new_n579), .ZN(new_n580));
  OAI21_X1  g0380(.A(new_n497), .B1(new_n577), .B2(new_n580), .ZN(new_n581));
  OAI21_X1  g0381(.A(new_n386), .B1(new_n575), .B2(new_n581), .ZN(new_n582));
  AND3_X1   g0382(.A1(new_n565), .A2(new_n570), .A3(KEYINPUT85), .ZN(new_n583));
  AOI21_X1  g0383(.A(KEYINPUT85), .B1(new_n565), .B2(new_n570), .ZN(new_n584));
  OAI21_X1  g0384(.A(new_n286), .B1(new_n583), .B2(new_n584), .ZN(new_n585));
  INV_X1    g0385(.A(new_n497), .ZN(new_n586));
  NAND3_X1  g0386(.A1(new_n551), .A2(new_n576), .A3(G257), .ZN(new_n587));
  OAI21_X1  g0387(.A(KEYINPUT86), .B1(new_n578), .B2(new_n579), .ZN(new_n588));
  AOI21_X1  g0388(.A(new_n586), .B1(new_n587), .B2(new_n588), .ZN(new_n589));
  NAND3_X1  g0389(.A1(new_n585), .A2(new_n297), .A3(new_n589), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n582), .A2(new_n590), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n301), .A2(new_n284), .ZN(new_n592));
  OAI21_X1  g0392(.A(new_n592), .B1(new_n473), .B2(new_n284), .ZN(new_n593));
  AOI21_X1  g0393(.A(new_n352), .B1(new_n410), .B2(new_n403), .ZN(new_n594));
  NAND3_X1  g0394(.A1(new_n484), .A2(KEYINPUT6), .A3(new_n485), .ZN(new_n595));
  INV_X1    g0395(.A(KEYINPUT6), .ZN(new_n596));
  NAND3_X1  g0396(.A1(new_n596), .A2(new_n352), .A3(G97), .ZN(new_n597));
  OAI21_X1  g0397(.A(G107), .B1(new_n284), .B2(KEYINPUT6), .ZN(new_n598));
  NAND4_X1  g0398(.A1(new_n595), .A2(G20), .A3(new_n597), .A4(new_n598), .ZN(new_n599));
  NOR4_X1   g0399(.A1(new_n225), .A2(KEYINPUT82), .A3(G20), .A4(G33), .ZN(new_n600));
  INV_X1    g0400(.A(KEYINPUT82), .ZN(new_n601));
  AOI21_X1  g0401(.A(new_n601), .B1(new_n309), .B2(G77), .ZN(new_n602));
  NOR2_X1   g0402(.A1(new_n600), .A2(new_n602), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n599), .A2(new_n603), .ZN(new_n604));
  OAI21_X1  g0404(.A(new_n303), .B1(new_n594), .B2(new_n604), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n605), .A2(KEYINPUT84), .ZN(new_n606));
  INV_X1    g0406(.A(KEYINPUT84), .ZN(new_n607));
  OAI211_X1 g0407(.A(new_n607), .B(new_n303), .C1(new_n594), .C2(new_n604), .ZN(new_n608));
  AOI21_X1  g0408(.A(new_n593), .B1(new_n606), .B2(new_n608), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n591), .A2(new_n609), .ZN(new_n610));
  INV_X1    g0410(.A(new_n593), .ZN(new_n611));
  OAI21_X1  g0411(.A(G107), .B1(new_n399), .B2(new_n404), .ZN(new_n612));
  NAND3_X1  g0412(.A1(new_n612), .A2(new_n599), .A3(new_n603), .ZN(new_n613));
  AOI21_X1  g0413(.A(new_n607), .B1(new_n613), .B2(new_n303), .ZN(new_n614));
  INV_X1    g0414(.A(new_n608), .ZN(new_n615));
  OAI21_X1  g0415(.A(new_n611), .B1(new_n614), .B2(new_n615), .ZN(new_n616));
  AOI21_X1  g0416(.A(G169), .B1(new_n585), .B2(new_n589), .ZN(new_n617));
  INV_X1    g0417(.A(new_n617), .ZN(new_n618));
  NAND3_X1  g0418(.A1(new_n585), .A2(new_n330), .A3(new_n589), .ZN(new_n619));
  NAND3_X1  g0419(.A1(new_n616), .A2(new_n618), .A3(new_n619), .ZN(new_n620));
  INV_X1    g0420(.A(new_n341), .ZN(new_n621));
  NOR2_X1   g0421(.A1(new_n621), .A2(new_n300), .ZN(new_n622));
  INV_X1    g0422(.A(KEYINPUT19), .ZN(new_n623));
  OAI21_X1  g0423(.A(new_n623), .B1(new_n479), .B2(new_n311), .ZN(new_n624));
  NOR2_X1   g0424(.A1(G87), .A2(G107), .ZN(new_n625));
  NAND3_X1  g0425(.A1(new_n484), .A2(new_n485), .A3(new_n625), .ZN(new_n626));
  NAND3_X1  g0426(.A1(KEYINPUT19), .A2(G33), .A3(G97), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n627), .A2(new_n217), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n626), .A2(new_n628), .ZN(new_n629));
  NAND3_X1  g0429(.A1(new_n268), .A2(new_n217), .A3(G68), .ZN(new_n630));
  NAND3_X1  g0430(.A1(new_n624), .A2(new_n629), .A3(new_n630), .ZN(new_n631));
  AOI21_X1  g0431(.A(new_n622), .B1(new_n631), .B2(new_n303), .ZN(new_n632));
  OR2_X1    g0432(.A1(new_n473), .A2(new_n341), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n254), .A2(G45), .ZN(new_n635));
  NAND3_X1  g0435(.A1(new_n270), .A2(G250), .A3(new_n635), .ZN(new_n636));
  NOR2_X1   g0436(.A1(G238), .A2(G1698), .ZN(new_n637));
  AOI21_X1  g0437(.A(new_n637), .B1(new_n226), .B2(G1698), .ZN(new_n638));
  AOI22_X1  g0438(.A1(new_n638), .A2(new_n268), .B1(G33), .B2(G116), .ZN(new_n639));
  OAI21_X1  g0439(.A(new_n636), .B1(new_n639), .B2(new_n270), .ZN(new_n640));
  AOI21_X1  g0440(.A(KEYINPUT87), .B1(new_n263), .B2(new_n491), .ZN(new_n641));
  AND4_X1   g0441(.A1(KEYINPUT87), .A2(new_n270), .A3(G274), .A4(new_n491), .ZN(new_n642));
  NOR2_X1   g0442(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  OAI21_X1  g0443(.A(new_n327), .B1(new_n640), .B2(new_n643), .ZN(new_n644));
  INV_X1    g0444(.A(new_n636), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n226), .A2(G1698), .ZN(new_n646));
  OAI21_X1  g0446(.A(new_n646), .B1(G238), .B2(G1698), .ZN(new_n647));
  OAI22_X1  g0447(.A1(new_n647), .A2(new_n282), .B1(new_n283), .B2(new_n470), .ZN(new_n648));
  AOI21_X1  g0448(.A(new_n645), .B1(new_n648), .B2(new_n286), .ZN(new_n649));
  INV_X1    g0449(.A(KEYINPUT87), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n270), .A2(G274), .ZN(new_n651));
  OAI21_X1  g0451(.A(new_n650), .B1(new_n651), .B2(new_n635), .ZN(new_n652));
  NAND3_X1  g0452(.A1(new_n263), .A2(KEYINPUT87), .A3(new_n491), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  NAND3_X1  g0454(.A1(new_n649), .A2(new_n330), .A3(new_n654), .ZN(new_n655));
  NAND3_X1  g0455(.A1(new_n634), .A2(new_n644), .A3(new_n655), .ZN(new_n656));
  INV_X1    g0456(.A(G87), .ZN(new_n657));
  NOR2_X1   g0457(.A1(new_n473), .A2(new_n657), .ZN(new_n658));
  AOI211_X1 g0458(.A(new_n622), .B(new_n658), .C1(new_n631), .C2(new_n303), .ZN(new_n659));
  OAI21_X1  g0459(.A(G200), .B1(new_n640), .B2(new_n643), .ZN(new_n660));
  NAND3_X1  g0460(.A1(new_n649), .A2(G190), .A3(new_n654), .ZN(new_n661));
  NAND3_X1  g0461(.A1(new_n659), .A2(new_n660), .A3(new_n661), .ZN(new_n662));
  AND2_X1   g0462(.A1(new_n656), .A2(new_n662), .ZN(new_n663));
  AND3_X1   g0463(.A1(new_n610), .A2(new_n620), .A3(new_n663), .ZN(new_n664));
  AND4_X1   g0464(.A1(new_n469), .A2(new_n518), .A3(new_n562), .A4(new_n664), .ZN(G372));
  NAND2_X1  g0465(.A1(new_n460), .A2(new_n463), .ZN(new_n666));
  INV_X1    g0466(.A(KEYINPUT93), .ZN(new_n667));
  NAND3_X1  g0467(.A1(new_n359), .A2(new_n667), .A3(new_n360), .ZN(new_n668));
  INV_X1    g0468(.A(new_n668), .ZN(new_n669));
  AOI21_X1  g0469(.A(new_n667), .B1(new_n359), .B2(new_n360), .ZN(new_n670));
  NOR2_X1   g0470(.A1(new_n669), .A2(new_n670), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n326), .A2(new_n671), .ZN(new_n672));
  AOI22_X1  g0472(.A1(new_n333), .A2(KEYINPUT14), .B1(new_n291), .B2(G179), .ZN(new_n673));
  AND3_X1   g0473(.A1(new_n328), .A2(KEYINPUT77), .A3(new_n329), .ZN(new_n674));
  AOI21_X1  g0474(.A(KEYINPUT77), .B1(new_n328), .B2(new_n329), .ZN(new_n675));
  OAI21_X1  g0475(.A(new_n673), .B1(new_n674), .B2(new_n675), .ZN(new_n676));
  INV_X1    g0476(.A(new_n324), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n672), .A2(new_n678), .ZN(new_n679));
  AND2_X1   g0479(.A1(new_n442), .A2(new_n467), .ZN(new_n680));
  AOI21_X1  g0480(.A(new_n666), .B1(new_n679), .B2(new_n680), .ZN(new_n681));
  NOR2_X1   g0481(.A1(new_n389), .A2(new_n384), .ZN(new_n682));
  OAI21_X1  g0482(.A(new_n377), .B1(new_n681), .B2(new_n682), .ZN(new_n683));
  INV_X1    g0483(.A(new_n683), .ZN(new_n684));
  OR3_X1    g0484(.A1(new_n337), .A2(new_n390), .A3(new_n468), .ZN(new_n685));
  INV_X1    g0485(.A(KEYINPUT26), .ZN(new_n686));
  INV_X1    g0486(.A(KEYINPUT91), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n649), .A2(new_n654), .ZN(new_n688));
  AOI21_X1  g0488(.A(new_n687), .B1(new_n688), .B2(new_n327), .ZN(new_n689));
  AOI211_X1 g0489(.A(KEYINPUT91), .B(G169), .C1(new_n649), .C2(new_n654), .ZN(new_n690));
  NOR2_X1   g0490(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  NOR2_X1   g0491(.A1(new_n640), .A2(new_n643), .ZN(new_n692));
  AOI22_X1  g0492(.A1(new_n692), .A2(new_n330), .B1(new_n632), .B2(new_n633), .ZN(new_n693));
  INV_X1    g0493(.A(new_n693), .ZN(new_n694));
  OAI21_X1  g0494(.A(new_n662), .B1(new_n691), .B2(new_n694), .ZN(new_n695));
  OAI21_X1  g0495(.A(new_n686), .B1(new_n695), .B2(new_n620), .ZN(new_n696));
  AND3_X1   g0496(.A1(new_n585), .A2(new_n330), .A3(new_n589), .ZN(new_n697));
  NOR2_X1   g0497(.A1(new_n609), .A2(new_n697), .ZN(new_n698));
  NAND4_X1  g0498(.A1(new_n698), .A2(new_n663), .A3(KEYINPUT26), .A4(new_n618), .ZN(new_n699));
  NAND3_X1  g0499(.A1(new_n696), .A2(KEYINPUT92), .A3(new_n699), .ZN(new_n700));
  NAND2_X1  g0500(.A1(new_n644), .A2(KEYINPUT91), .ZN(new_n701));
  NAND3_X1  g0501(.A1(new_n688), .A2(new_n687), .A3(new_n327), .ZN(new_n702));
  NAND2_X1  g0502(.A1(new_n701), .A2(new_n702), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n703), .A2(new_n693), .ZN(new_n704));
  AOI22_X1  g0504(.A1(new_n698), .A2(new_n618), .B1(new_n609), .B2(new_n591), .ZN(new_n705));
  AND3_X1   g0505(.A1(new_n704), .A2(new_n561), .A3(new_n662), .ZN(new_n706));
  OAI21_X1  g0506(.A(new_n557), .B1(new_n533), .B2(new_n539), .ZN(new_n707));
  OAI211_X1 g0507(.A(new_n707), .B(new_n511), .C1(new_n515), .C2(new_n516), .ZN(new_n708));
  NAND3_X1  g0508(.A1(new_n705), .A2(new_n706), .A3(new_n708), .ZN(new_n709));
  NOR3_X1   g0509(.A1(new_n609), .A2(new_n697), .A3(new_n617), .ZN(new_n710));
  INV_X1    g0510(.A(KEYINPUT92), .ZN(new_n711));
  NAND4_X1  g0511(.A1(new_n710), .A2(new_n711), .A3(KEYINPUT26), .A4(new_n663), .ZN(new_n712));
  NAND4_X1  g0512(.A1(new_n700), .A2(new_n704), .A3(new_n709), .A4(new_n712), .ZN(new_n713));
  INV_X1    g0513(.A(new_n713), .ZN(new_n714));
  OAI21_X1  g0514(.A(new_n684), .B1(new_n685), .B2(new_n714), .ZN(G369));
  INV_X1    g0515(.A(KEYINPUT20), .ZN(new_n716));
  NOR2_X1   g0516(.A1(new_n486), .A2(new_n487), .ZN(new_n717));
  INV_X1    g0517(.A(new_n481), .ZN(new_n718));
  OAI21_X1  g0518(.A(new_n716), .B1(new_n717), .B2(new_n718), .ZN(new_n719));
  AOI21_X1  g0519(.A(new_n474), .B1(new_n719), .B2(new_n488), .ZN(new_n720));
  AOI21_X1  g0520(.A(new_n720), .B1(new_n508), .B2(new_n509), .ZN(new_n721));
  AND2_X1   g0521(.A1(new_n502), .A2(new_n286), .ZN(new_n722));
  NAND2_X1  g0522(.A1(new_n495), .A2(new_n497), .ZN(new_n723));
  OAI21_X1  g0523(.A(G169), .B1(new_n722), .B2(new_n723), .ZN(new_n724));
  OAI21_X1  g0524(.A(new_n514), .B1(new_n724), .B2(new_n720), .ZN(new_n725));
  NAND2_X1  g0525(.A1(new_n725), .A2(KEYINPUT88), .ZN(new_n726));
  NAND3_X1  g0526(.A1(new_n513), .A2(new_n512), .A3(new_n514), .ZN(new_n727));
  AOI21_X1  g0527(.A(new_n721), .B1(new_n726), .B2(new_n727), .ZN(new_n728));
  INV_X1    g0528(.A(new_n728), .ZN(new_n729));
  NAND3_X1  g0529(.A1(new_n254), .A2(new_n217), .A3(G13), .ZN(new_n730));
  OR2_X1    g0530(.A1(new_n730), .A2(KEYINPUT27), .ZN(new_n731));
  NAND2_X1  g0531(.A1(new_n730), .A2(KEYINPUT27), .ZN(new_n732));
  NAND3_X1  g0532(.A1(new_n731), .A2(G213), .A3(new_n732), .ZN(new_n733));
  INV_X1    g0533(.A(G343), .ZN(new_n734));
  NOR2_X1   g0534(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  INV_X1    g0535(.A(new_n735), .ZN(new_n736));
  NOR2_X1   g0536(.A1(new_n720), .A2(new_n736), .ZN(new_n737));
  NAND2_X1  g0537(.A1(new_n729), .A2(new_n737), .ZN(new_n738));
  OAI21_X1  g0538(.A(new_n738), .B1(new_n517), .B2(new_n737), .ZN(new_n739));
  AND2_X1   g0539(.A1(new_n739), .A2(G330), .ZN(new_n740));
  NAND3_X1  g0540(.A1(new_n540), .A2(new_n545), .A3(new_n735), .ZN(new_n741));
  NAND2_X1  g0541(.A1(new_n562), .A2(new_n741), .ZN(new_n742));
  OAI21_X1  g0542(.A(new_n742), .B1(new_n558), .B2(new_n736), .ZN(new_n743));
  NAND2_X1  g0543(.A1(new_n740), .A2(new_n743), .ZN(new_n744));
  NOR2_X1   g0544(.A1(new_n728), .A2(new_n735), .ZN(new_n745));
  AND2_X1   g0545(.A1(new_n562), .A2(new_n745), .ZN(new_n746));
  INV_X1    g0546(.A(new_n707), .ZN(new_n747));
  AOI21_X1  g0547(.A(new_n746), .B1(new_n747), .B2(new_n736), .ZN(new_n748));
  NAND2_X1  g0548(.A1(new_n744), .A2(new_n748), .ZN(G399));
  NOR2_X1   g0549(.A1(new_n213), .A2(G41), .ZN(new_n750));
  NAND3_X1  g0550(.A1(new_n479), .A2(new_n470), .A3(new_n625), .ZN(new_n751));
  NOR3_X1   g0551(.A1(new_n750), .A2(new_n254), .A3(new_n751), .ZN(new_n752));
  AOI21_X1  g0552(.A(new_n752), .B1(new_n221), .B2(new_n750), .ZN(new_n753));
  XOR2_X1   g0553(.A(new_n753), .B(KEYINPUT28), .Z(new_n754));
  NAND2_X1  g0554(.A1(new_n728), .A2(new_n558), .ZN(new_n755));
  NAND3_X1  g0555(.A1(new_n755), .A2(new_n705), .A3(new_n706), .ZN(new_n756));
  NAND2_X1  g0556(.A1(new_n656), .A2(new_n662), .ZN(new_n757));
  OAI21_X1  g0557(.A(new_n686), .B1(new_n620), .B2(new_n757), .ZN(new_n758));
  AND2_X1   g0558(.A1(new_n660), .A2(new_n661), .ZN(new_n759));
  AOI22_X1  g0559(.A1(new_n703), .A2(new_n693), .B1(new_n759), .B2(new_n659), .ZN(new_n760));
  NAND3_X1  g0560(.A1(new_n710), .A2(new_n760), .A3(KEYINPUT26), .ZN(new_n761));
  NAND2_X1  g0561(.A1(new_n758), .A2(new_n761), .ZN(new_n762));
  NAND3_X1  g0562(.A1(new_n756), .A2(new_n762), .A3(new_n704), .ZN(new_n763));
  INV_X1    g0563(.A(KEYINPUT94), .ZN(new_n764));
  AND3_X1   g0564(.A1(new_n763), .A2(new_n764), .A3(new_n736), .ZN(new_n765));
  AOI21_X1  g0565(.A(new_n764), .B1(new_n763), .B2(new_n736), .ZN(new_n766));
  OAI21_X1  g0566(.A(KEYINPUT29), .B1(new_n765), .B2(new_n766), .ZN(new_n767));
  AOI21_X1  g0567(.A(KEYINPUT29), .B1(new_n713), .B2(new_n736), .ZN(new_n768));
  INV_X1    g0568(.A(new_n768), .ZN(new_n769));
  INV_X1    g0569(.A(KEYINPUT30), .ZN(new_n770));
  AOI21_X1  g0570(.A(new_n723), .B1(new_n286), .B2(new_n502), .ZN(new_n771));
  NAND4_X1  g0571(.A1(new_n692), .A2(new_n771), .A3(G179), .A4(new_n555), .ZN(new_n772));
  NAND2_X1  g0572(.A1(new_n585), .A2(new_n589), .ZN(new_n773));
  OAI21_X1  g0573(.A(new_n770), .B1(new_n772), .B2(new_n773), .ZN(new_n774));
  NAND4_X1  g0574(.A1(new_n649), .A2(new_n550), .A3(new_n552), .A4(new_n654), .ZN(new_n775));
  NOR2_X1   g0575(.A1(new_n775), .A2(new_n509), .ZN(new_n776));
  NAND4_X1  g0576(.A1(new_n776), .A2(KEYINPUT30), .A3(new_n585), .A4(new_n589), .ZN(new_n777));
  NOR2_X1   g0577(.A1(new_n692), .A2(G179), .ZN(new_n778));
  NAND4_X1  g0578(.A1(new_n778), .A2(new_n773), .A3(new_n504), .A4(new_n553), .ZN(new_n779));
  NAND3_X1  g0579(.A1(new_n774), .A2(new_n777), .A3(new_n779), .ZN(new_n780));
  AND3_X1   g0580(.A1(new_n780), .A2(KEYINPUT31), .A3(new_n735), .ZN(new_n781));
  AOI21_X1  g0581(.A(KEYINPUT31), .B1(new_n780), .B2(new_n735), .ZN(new_n782));
  NOR2_X1   g0582(.A1(new_n781), .A2(new_n782), .ZN(new_n783));
  NAND4_X1  g0583(.A1(new_n664), .A2(new_n562), .A3(new_n518), .A4(new_n736), .ZN(new_n784));
  NAND2_X1  g0584(.A1(new_n783), .A2(new_n784), .ZN(new_n785));
  AOI22_X1  g0585(.A1(new_n767), .A2(new_n769), .B1(G330), .B2(new_n785), .ZN(new_n786));
  OAI21_X1  g0586(.A(new_n754), .B1(new_n786), .B2(G1), .ZN(G364));
  AND2_X1   g0587(.A1(new_n217), .A2(G13), .ZN(new_n788));
  AOI21_X1  g0588(.A(new_n254), .B1(new_n788), .B2(G45), .ZN(new_n789));
  INV_X1    g0589(.A(new_n789), .ZN(new_n790));
  NOR2_X1   g0590(.A1(new_n750), .A2(new_n790), .ZN(new_n791));
  NOR2_X1   g0591(.A1(new_n740), .A2(new_n791), .ZN(new_n792));
  OAI21_X1  g0592(.A(new_n792), .B1(G330), .B2(new_n739), .ZN(new_n793));
  NAND3_X1  g0593(.A1(G355), .A2(new_n212), .A3(new_n268), .ZN(new_n794));
  OAI21_X1  g0594(.A(new_n794), .B1(G116), .B2(new_n212), .ZN(new_n795));
  NOR2_X1   g0595(.A1(new_n213), .A2(new_n268), .ZN(new_n796));
  INV_X1    g0596(.A(new_n796), .ZN(new_n797));
  AOI21_X1  g0597(.A(new_n797), .B1(new_n431), .B2(new_n221), .ZN(new_n798));
  NAND2_X1  g0598(.A1(new_n252), .A2(G45), .ZN(new_n799));
  AOI21_X1  g0599(.A(new_n795), .B1(new_n798), .B2(new_n799), .ZN(new_n800));
  NOR2_X1   g0600(.A1(G13), .A2(G33), .ZN(new_n801));
  INV_X1    g0601(.A(new_n801), .ZN(new_n802));
  NOR2_X1   g0602(.A1(new_n802), .A2(G20), .ZN(new_n803));
  AOI21_X1  g0603(.A(new_n216), .B1(G20), .B2(new_n327), .ZN(new_n804));
  NOR2_X1   g0604(.A1(new_n803), .A2(new_n804), .ZN(new_n805));
  INV_X1    g0605(.A(new_n805), .ZN(new_n806));
  OAI21_X1  g0606(.A(new_n791), .B1(new_n800), .B2(new_n806), .ZN(new_n807));
  NOR2_X1   g0607(.A1(new_n297), .A2(G200), .ZN(new_n808));
  NAND2_X1  g0608(.A1(new_n808), .A2(new_n330), .ZN(new_n809));
  NAND2_X1  g0609(.A1(new_n809), .A2(G20), .ZN(new_n810));
  INV_X1    g0610(.A(new_n810), .ZN(new_n811));
  NOR2_X1   g0611(.A1(new_n217), .A2(G179), .ZN(new_n812));
  NAND3_X1  g0612(.A1(new_n812), .A2(G190), .A3(G200), .ZN(new_n813));
  INV_X1    g0613(.A(G303), .ZN(new_n814));
  OAI22_X1  g0614(.A1(new_n811), .A2(new_n548), .B1(new_n813), .B2(new_n814), .ZN(new_n815));
  NOR2_X1   g0615(.A1(new_n217), .A2(new_n330), .ZN(new_n816));
  NAND2_X1  g0616(.A1(new_n816), .A2(G200), .ZN(new_n817));
  NOR2_X1   g0617(.A1(new_n817), .A2(G190), .ZN(new_n818));
  INV_X1    g0618(.A(new_n818), .ZN(new_n819));
  XOR2_X1   g0619(.A(KEYINPUT33), .B(G317), .Z(new_n820));
  NOR2_X1   g0620(.A1(new_n819), .A2(new_n820), .ZN(new_n821));
  NOR2_X1   g0621(.A1(new_n817), .A2(new_n297), .ZN(new_n822));
  AOI211_X1 g0622(.A(new_n815), .B(new_n821), .C1(G326), .C2(new_n822), .ZN(new_n823));
  NOR2_X1   g0623(.A1(G190), .A2(G200), .ZN(new_n824));
  NAND2_X1  g0624(.A1(new_n812), .A2(new_n824), .ZN(new_n825));
  INV_X1    g0625(.A(new_n825), .ZN(new_n826));
  AOI21_X1  g0626(.A(new_n268), .B1(new_n826), .B2(G329), .ZN(new_n827));
  INV_X1    g0627(.A(G283), .ZN(new_n828));
  NAND3_X1  g0628(.A1(new_n812), .A2(new_n297), .A3(G200), .ZN(new_n829));
  OAI21_X1  g0629(.A(new_n827), .B1(new_n828), .B2(new_n829), .ZN(new_n830));
  XOR2_X1   g0630(.A(new_n816), .B(KEYINPUT95), .Z(new_n831));
  INV_X1    g0631(.A(new_n831), .ZN(new_n832));
  NAND2_X1  g0632(.A1(new_n832), .A2(new_n808), .ZN(new_n833));
  INV_X1    g0633(.A(new_n833), .ZN(new_n834));
  AOI21_X1  g0634(.A(new_n830), .B1(new_n834), .B2(G322), .ZN(new_n835));
  INV_X1    g0635(.A(G311), .ZN(new_n836));
  NAND2_X1  g0636(.A1(new_n832), .A2(new_n824), .ZN(new_n837));
  OAI211_X1 g0637(.A(new_n823), .B(new_n835), .C1(new_n836), .C2(new_n837), .ZN(new_n838));
  INV_X1    g0638(.A(new_n822), .ZN(new_n839));
  OAI22_X1  g0639(.A1(new_n839), .A2(new_n220), .B1(new_n811), .B2(new_n284), .ZN(new_n840));
  AOI211_X1 g0640(.A(new_n282), .B(new_n840), .C1(G68), .C2(new_n818), .ZN(new_n841));
  OAI221_X1 g0641(.A(new_n841), .B1(new_n201), .B2(new_n833), .C1(new_n225), .C2(new_n837), .ZN(new_n842));
  INV_X1    g0642(.A(G159), .ZN(new_n843));
  NOR2_X1   g0643(.A1(new_n825), .A2(new_n843), .ZN(new_n844));
  XNOR2_X1  g0644(.A(new_n844), .B(KEYINPUT32), .ZN(new_n845));
  OAI221_X1 g0645(.A(new_n845), .B1(new_n657), .B2(new_n813), .C1(new_n352), .C2(new_n829), .ZN(new_n846));
  OAI21_X1  g0646(.A(new_n838), .B1(new_n842), .B2(new_n846), .ZN(new_n847));
  OR2_X1    g0647(.A1(new_n847), .A2(KEYINPUT96), .ZN(new_n848));
  INV_X1    g0648(.A(new_n804), .ZN(new_n849));
  AOI21_X1  g0649(.A(new_n849), .B1(new_n847), .B2(KEYINPUT96), .ZN(new_n850));
  AOI21_X1  g0650(.A(new_n807), .B1(new_n848), .B2(new_n850), .ZN(new_n851));
  INV_X1    g0651(.A(new_n803), .ZN(new_n852));
  OAI21_X1  g0652(.A(new_n851), .B1(new_n739), .B2(new_n852), .ZN(new_n853));
  NAND2_X1  g0653(.A1(new_n793), .A2(new_n853), .ZN(new_n854));
  XNOR2_X1  g0654(.A(new_n854), .B(KEYINPUT97), .ZN(G396));
  NAND2_X1  g0655(.A1(new_n713), .A2(new_n736), .ZN(new_n856));
  INV_X1    g0656(.A(KEYINPUT101), .ZN(new_n857));
  NAND2_X1  g0657(.A1(new_n348), .A2(new_n735), .ZN(new_n858));
  NOR3_X1   g0658(.A1(new_n669), .A2(new_n670), .A3(new_n858), .ZN(new_n859));
  NAND3_X1  g0659(.A1(new_n358), .A2(new_n361), .A3(new_n858), .ZN(new_n860));
  INV_X1    g0660(.A(new_n860), .ZN(new_n861));
  OAI21_X1  g0661(.A(new_n857), .B1(new_n859), .B2(new_n861), .ZN(new_n862));
  INV_X1    g0662(.A(new_n670), .ZN(new_n863));
  NAND2_X1  g0663(.A1(new_n863), .A2(new_n668), .ZN(new_n864));
  OAI211_X1 g0664(.A(KEYINPUT101), .B(new_n860), .C1(new_n864), .C2(new_n858), .ZN(new_n865));
  NAND2_X1  g0665(.A1(new_n862), .A2(new_n865), .ZN(new_n866));
  INV_X1    g0666(.A(new_n866), .ZN(new_n867));
  AND2_X1   g0667(.A1(new_n362), .A2(new_n736), .ZN(new_n868));
  AOI22_X1  g0668(.A1(new_n856), .A2(new_n867), .B1(new_n713), .B2(new_n868), .ZN(new_n869));
  INV_X1    g0669(.A(new_n869), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n785), .A2(G330), .ZN(new_n871));
  NOR2_X1   g0671(.A1(new_n870), .A2(new_n871), .ZN(new_n872));
  INV_X1    g0672(.A(new_n872), .ZN(new_n873));
  AOI21_X1  g0673(.A(new_n791), .B1(new_n870), .B2(new_n871), .ZN(new_n874));
  NOR2_X1   g0674(.A1(new_n859), .A2(new_n861), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n875), .A2(new_n801), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n849), .A2(new_n802), .ZN(new_n877));
  OAI21_X1  g0677(.A(new_n791), .B1(G77), .B2(new_n877), .ZN(new_n878));
  XNOR2_X1  g0678(.A(new_n878), .B(KEYINPUT98), .ZN(new_n879));
  AOI22_X1  g0679(.A1(new_n818), .A2(G150), .B1(new_n822), .B2(G137), .ZN(new_n880));
  INV_X1    g0680(.A(G143), .ZN(new_n881));
  OAI221_X1 g0681(.A(new_n880), .B1(new_n837), .B2(new_n843), .C1(new_n881), .C2(new_n833), .ZN(new_n882));
  INV_X1    g0682(.A(KEYINPUT34), .ZN(new_n883));
  AND2_X1   g0683(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  AOI21_X1  g0684(.A(new_n282), .B1(new_n826), .B2(G132), .ZN(new_n885));
  OAI21_X1  g0685(.A(new_n885), .B1(new_n202), .B2(new_n829), .ZN(new_n886));
  OAI22_X1  g0686(.A1(new_n811), .A2(new_n201), .B1(new_n813), .B2(new_n220), .ZN(new_n887));
  NOR3_X1   g0687(.A1(new_n884), .A2(new_n886), .A3(new_n887), .ZN(new_n888));
  OAI21_X1  g0688(.A(new_n888), .B1(new_n883), .B2(new_n882), .ZN(new_n889));
  AOI22_X1  g0689(.A1(new_n818), .A2(G283), .B1(new_n822), .B2(G303), .ZN(new_n890));
  OAI21_X1  g0690(.A(new_n890), .B1(new_n837), .B2(new_n470), .ZN(new_n891));
  XOR2_X1   g0691(.A(new_n891), .B(KEYINPUT99), .Z(new_n892));
  OAI22_X1  g0692(.A1(new_n833), .A2(new_n548), .B1(new_n284), .B2(new_n811), .ZN(new_n893));
  XOR2_X1   g0693(.A(new_n893), .B(KEYINPUT100), .Z(new_n894));
  NOR2_X1   g0694(.A1(new_n829), .A2(new_n657), .ZN(new_n895));
  OAI21_X1  g0695(.A(new_n282), .B1(new_n825), .B2(new_n836), .ZN(new_n896));
  INV_X1    g0696(.A(new_n813), .ZN(new_n897));
  AOI211_X1 g0697(.A(new_n895), .B(new_n896), .C1(G107), .C2(new_n897), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n894), .A2(new_n898), .ZN(new_n899));
  OAI21_X1  g0699(.A(new_n889), .B1(new_n892), .B2(new_n899), .ZN(new_n900));
  AOI21_X1  g0700(.A(new_n879), .B1(new_n900), .B2(new_n804), .ZN(new_n901));
  AOI22_X1  g0701(.A1(new_n873), .A2(new_n874), .B1(new_n876), .B2(new_n901), .ZN(new_n902));
  INV_X1    g0702(.A(new_n902), .ZN(G384));
  NAND3_X1  g0703(.A1(new_n595), .A2(new_n597), .A3(new_n598), .ZN(new_n904));
  INV_X1    g0704(.A(KEYINPUT35), .ZN(new_n905));
  OAI211_X1 g0705(.A(G116), .B(new_n218), .C1(new_n904), .C2(new_n905), .ZN(new_n906));
  AOI21_X1  g0706(.A(new_n906), .B1(new_n905), .B2(new_n904), .ZN(new_n907));
  XNOR2_X1  g0707(.A(new_n907), .B(KEYINPUT36), .ZN(new_n908));
  NAND3_X1  g0708(.A1(new_n221), .A2(G77), .A3(new_n394), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n220), .A2(G68), .ZN(new_n910));
  AOI211_X1 g0710(.A(new_n254), .B(G13), .C1(new_n909), .C2(new_n910), .ZN(new_n911));
  NOR2_X1   g0711(.A1(new_n908), .A2(new_n911), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n445), .A2(new_n446), .ZN(new_n913));
  AOI21_X1  g0713(.A(KEYINPUT16), .B1(new_n913), .B2(new_n414), .ZN(new_n914));
  OAI21_X1  g0714(.A(new_n393), .B1(new_n421), .B2(new_n914), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n461), .A2(new_n915), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n453), .A2(new_n466), .ZN(new_n917));
  INV_X1    g0717(.A(new_n733), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n915), .A2(new_n918), .ZN(new_n919));
  NAND3_X1  g0719(.A1(new_n916), .A2(new_n917), .A3(new_n919), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n920), .A2(KEYINPUT37), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n422), .A2(new_n461), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n422), .A2(new_n918), .ZN(new_n923));
  INV_X1    g0723(.A(KEYINPUT37), .ZN(new_n924));
  NAND4_X1  g0724(.A1(new_n922), .A2(new_n923), .A3(new_n917), .A4(new_n924), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n921), .A2(new_n925), .ZN(new_n926));
  INV_X1    g0726(.A(new_n919), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n468), .A2(new_n927), .ZN(new_n928));
  AND3_X1   g0728(.A1(new_n926), .A2(new_n928), .A3(KEYINPUT38), .ZN(new_n929));
  AOI21_X1  g0729(.A(KEYINPUT38), .B1(new_n926), .B2(new_n928), .ZN(new_n930));
  NOR2_X1   g0730(.A1(new_n929), .A2(new_n930), .ZN(new_n931));
  NOR2_X1   g0731(.A1(new_n361), .A2(new_n735), .ZN(new_n932));
  AOI21_X1  g0732(.A(new_n932), .B1(new_n713), .B2(new_n868), .ZN(new_n933));
  NAND3_X1  g0733(.A1(new_n320), .A2(new_n323), .A3(new_n735), .ZN(new_n934));
  XNOR2_X1  g0734(.A(new_n934), .B(KEYINPUT102), .ZN(new_n935));
  NAND3_X1  g0735(.A1(new_n678), .A2(new_n326), .A3(new_n935), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n336), .A2(new_n326), .ZN(new_n937));
  NAND3_X1  g0737(.A1(new_n937), .A2(new_n677), .A3(new_n735), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n936), .A2(new_n938), .ZN(new_n939));
  INV_X1    g0739(.A(new_n939), .ZN(new_n940));
  NOR3_X1   g0740(.A1(new_n931), .A2(new_n933), .A3(new_n940), .ZN(new_n941));
  NAND2_X1  g0741(.A1(new_n666), .A2(new_n733), .ZN(new_n942));
  INV_X1    g0742(.A(new_n942), .ZN(new_n943));
  OAI21_X1  g0743(.A(KEYINPUT103), .B1(new_n941), .B2(new_n943), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n926), .A2(new_n928), .ZN(new_n945));
  INV_X1    g0745(.A(KEYINPUT38), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n945), .A2(new_n946), .ZN(new_n947));
  NAND3_X1  g0747(.A1(new_n926), .A2(new_n928), .A3(KEYINPUT38), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n947), .A2(new_n948), .ZN(new_n949));
  NAND4_X1  g0749(.A1(new_n610), .A2(new_n760), .A3(new_n620), .A4(new_n561), .ZN(new_n950));
  INV_X1    g0750(.A(new_n708), .ZN(new_n951));
  OAI211_X1 g0751(.A(new_n704), .B(new_n712), .C1(new_n950), .C2(new_n951), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n699), .A2(KEYINPUT92), .ZN(new_n953));
  AOI21_X1  g0753(.A(KEYINPUT26), .B1(new_n710), .B2(new_n760), .ZN(new_n954));
  NOR2_X1   g0754(.A1(new_n953), .A2(new_n954), .ZN(new_n955));
  OAI21_X1  g0755(.A(new_n868), .B1(new_n952), .B2(new_n955), .ZN(new_n956));
  INV_X1    g0756(.A(new_n932), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n956), .A2(new_n957), .ZN(new_n958));
  NAND3_X1  g0758(.A1(new_n949), .A2(new_n958), .A3(new_n939), .ZN(new_n959));
  INV_X1    g0759(.A(KEYINPUT103), .ZN(new_n960));
  NAND3_X1  g0760(.A1(new_n959), .A2(new_n960), .A3(new_n942), .ZN(new_n961));
  INV_X1    g0761(.A(KEYINPUT39), .ZN(new_n962));
  NAND3_X1  g0762(.A1(new_n922), .A2(new_n923), .A3(new_n917), .ZN(new_n963));
  NAND2_X1  g0763(.A1(new_n963), .A2(KEYINPUT37), .ZN(new_n964));
  NAND2_X1  g0764(.A1(new_n964), .A2(new_n925), .ZN(new_n965));
  INV_X1    g0765(.A(new_n923), .ZN(new_n966));
  NAND2_X1  g0766(.A1(new_n468), .A2(new_n966), .ZN(new_n967));
  AOI21_X1  g0767(.A(KEYINPUT38), .B1(new_n965), .B2(new_n967), .ZN(new_n968));
  OAI21_X1  g0768(.A(new_n962), .B1(new_n929), .B2(new_n968), .ZN(new_n969));
  NAND3_X1  g0769(.A1(new_n947), .A2(KEYINPUT39), .A3(new_n948), .ZN(new_n970));
  AND2_X1   g0770(.A1(new_n969), .A2(new_n970), .ZN(new_n971));
  NOR2_X1   g0771(.A1(new_n678), .A2(new_n735), .ZN(new_n972));
  NAND2_X1  g0772(.A1(new_n971), .A2(new_n972), .ZN(new_n973));
  NAND3_X1  g0773(.A1(new_n944), .A2(new_n961), .A3(new_n973), .ZN(new_n974));
  INV_X1    g0774(.A(KEYINPUT29), .ZN(new_n975));
  AOI21_X1  g0775(.A(new_n685), .B1(new_n856), .B2(new_n975), .ZN(new_n976));
  AOI21_X1  g0776(.A(new_n683), .B1(new_n767), .B2(new_n976), .ZN(new_n977));
  XOR2_X1   g0777(.A(new_n974), .B(new_n977), .Z(new_n978));
  INV_X1    g0778(.A(G330), .ZN(new_n979));
  AOI21_X1  g0779(.A(new_n875), .B1(new_n783), .B2(new_n784), .ZN(new_n980));
  OAI211_X1 g0780(.A(new_n939), .B(new_n980), .C1(new_n929), .C2(new_n968), .ZN(new_n981));
  NAND2_X1  g0781(.A1(new_n981), .A2(KEYINPUT40), .ZN(new_n982));
  INV_X1    g0782(.A(KEYINPUT40), .ZN(new_n983));
  NAND4_X1  g0783(.A1(new_n949), .A2(new_n983), .A3(new_n939), .A4(new_n980), .ZN(new_n984));
  NAND2_X1  g0784(.A1(new_n982), .A2(new_n984), .ZN(new_n985));
  AND2_X1   g0785(.A1(new_n469), .A2(new_n785), .ZN(new_n986));
  AOI21_X1  g0786(.A(new_n979), .B1(new_n985), .B2(new_n986), .ZN(new_n987));
  OAI21_X1  g0787(.A(new_n987), .B1(new_n986), .B2(new_n985), .ZN(new_n988));
  NAND2_X1  g0788(.A1(new_n978), .A2(new_n988), .ZN(new_n989));
  OAI21_X1  g0789(.A(new_n989), .B1(new_n254), .B2(new_n788), .ZN(new_n990));
  NOR2_X1   g0790(.A1(new_n978), .A2(new_n988), .ZN(new_n991));
  OAI21_X1  g0791(.A(new_n912), .B1(new_n990), .B2(new_n991), .ZN(G367));
  OAI21_X1  g0792(.A(new_n705), .B1(new_n609), .B2(new_n736), .ZN(new_n993));
  XNOR2_X1  g0793(.A(new_n993), .B(KEYINPUT104), .ZN(new_n994));
  OAI21_X1  g0794(.A(new_n994), .B1(new_n620), .B2(new_n736), .ZN(new_n995));
  NAND2_X1  g0795(.A1(new_n995), .A2(new_n746), .ZN(new_n996));
  OR2_X1    g0796(.A1(new_n996), .A2(KEYINPUT42), .ZN(new_n997));
  OAI21_X1  g0797(.A(new_n620), .B1(new_n994), .B2(new_n558), .ZN(new_n998));
  NAND2_X1  g0798(.A1(new_n998), .A2(new_n736), .ZN(new_n999));
  NAND2_X1  g0799(.A1(new_n996), .A2(KEYINPUT42), .ZN(new_n1000));
  NAND3_X1  g0800(.A1(new_n997), .A2(new_n999), .A3(new_n1000), .ZN(new_n1001));
  INV_X1    g0801(.A(KEYINPUT105), .ZN(new_n1002));
  XNOR2_X1  g0802(.A(new_n1001), .B(new_n1002), .ZN(new_n1003));
  NOR2_X1   g0803(.A1(new_n659), .A2(new_n736), .ZN(new_n1004));
  NAND3_X1  g0804(.A1(new_n703), .A2(new_n693), .A3(new_n1004), .ZN(new_n1005));
  OAI21_X1  g0805(.A(new_n1005), .B1(new_n695), .B2(new_n1004), .ZN(new_n1006));
  XNOR2_X1  g0806(.A(new_n1006), .B(KEYINPUT43), .ZN(new_n1007));
  AND2_X1   g0807(.A1(new_n1003), .A2(new_n1007), .ZN(new_n1008));
  NOR2_X1   g0808(.A1(new_n1006), .A2(KEYINPUT43), .ZN(new_n1009));
  NOR2_X1   g0809(.A1(new_n1003), .A2(new_n1009), .ZN(new_n1010));
  INV_X1    g0810(.A(new_n744), .ZN(new_n1011));
  AND2_X1   g0811(.A1(new_n1011), .A2(new_n995), .ZN(new_n1012));
  OAI22_X1  g0812(.A1(new_n1008), .A2(new_n1010), .B1(KEYINPUT106), .B2(new_n1012), .ZN(new_n1013));
  NAND2_X1  g0813(.A1(new_n1012), .A2(KEYINPUT106), .ZN(new_n1014));
  NAND2_X1  g0814(.A1(new_n1013), .A2(new_n1014), .ZN(new_n1015));
  OAI211_X1 g0815(.A(KEYINPUT106), .B(new_n1012), .C1(new_n1008), .C2(new_n1010), .ZN(new_n1016));
  XOR2_X1   g0816(.A(new_n750), .B(KEYINPUT41), .Z(new_n1017));
  NAND2_X1  g0817(.A1(new_n995), .A2(new_n748), .ZN(new_n1018));
  XOR2_X1   g0818(.A(new_n1018), .B(KEYINPUT45), .Z(new_n1019));
  NOR2_X1   g0819(.A1(new_n995), .A2(new_n748), .ZN(new_n1020));
  XNOR2_X1  g0820(.A(new_n1020), .B(KEYINPUT44), .ZN(new_n1021));
  NAND2_X1  g0821(.A1(new_n1019), .A2(new_n1021), .ZN(new_n1022));
  NAND2_X1  g0822(.A1(new_n1011), .A2(KEYINPUT107), .ZN(new_n1023));
  XNOR2_X1  g0823(.A(new_n1022), .B(new_n1023), .ZN(new_n1024));
  INV_X1    g0824(.A(new_n746), .ZN(new_n1025));
  OAI21_X1  g0825(.A(new_n1025), .B1(new_n743), .B2(new_n745), .ZN(new_n1026));
  XNOR2_X1  g0826(.A(new_n1026), .B(new_n740), .ZN(new_n1027));
  NAND2_X1  g0827(.A1(new_n786), .A2(new_n1027), .ZN(new_n1028));
  INV_X1    g0828(.A(new_n1028), .ZN(new_n1029));
  NAND2_X1  g0829(.A1(new_n1024), .A2(new_n1029), .ZN(new_n1030));
  AOI21_X1  g0830(.A(new_n1017), .B1(new_n1030), .B2(new_n786), .ZN(new_n1031));
  OAI211_X1 g0831(.A(new_n1015), .B(new_n1016), .C1(new_n790), .C2(new_n1031), .ZN(new_n1032));
  NOR2_X1   g0832(.A1(new_n244), .A2(new_n797), .ZN(new_n1033));
  OAI21_X1  g0833(.A(new_n805), .B1(new_n212), .B2(new_n341), .ZN(new_n1034));
  OAI21_X1  g0834(.A(new_n791), .B1(new_n1033), .B2(new_n1034), .ZN(new_n1035));
  NOR2_X1   g0835(.A1(new_n811), .A2(new_n202), .ZN(new_n1036));
  OAI22_X1  g0836(.A1(new_n819), .A2(new_n843), .B1(new_n839), .B2(new_n881), .ZN(new_n1037));
  AOI211_X1 g0837(.A(new_n1036), .B(new_n1037), .C1(G58), .C2(new_n897), .ZN(new_n1038));
  NAND2_X1  g0838(.A1(new_n834), .A2(G150), .ZN(new_n1039));
  INV_X1    g0839(.A(new_n837), .ZN(new_n1040));
  NAND2_X1  g0840(.A1(new_n1040), .A2(G50), .ZN(new_n1041));
  INV_X1    g0841(.A(G137), .ZN(new_n1042));
  OAI21_X1  g0842(.A(new_n268), .B1(new_n825), .B2(new_n1042), .ZN(new_n1043));
  INV_X1    g0843(.A(new_n829), .ZN(new_n1044));
  AOI21_X1  g0844(.A(new_n1043), .B1(G77), .B2(new_n1044), .ZN(new_n1045));
  NAND4_X1  g0845(.A1(new_n1038), .A2(new_n1039), .A3(new_n1041), .A4(new_n1045), .ZN(new_n1046));
  NAND2_X1  g0846(.A1(new_n897), .A2(G116), .ZN(new_n1047));
  XNOR2_X1  g0847(.A(new_n1047), .B(KEYINPUT46), .ZN(new_n1048));
  OAI221_X1 g0848(.A(new_n1048), .B1(new_n837), .B2(new_n828), .C1(new_n814), .C2(new_n833), .ZN(new_n1049));
  OAI22_X1  g0849(.A1(new_n839), .A2(new_n836), .B1(new_n811), .B2(new_n352), .ZN(new_n1050));
  AOI21_X1  g0850(.A(new_n1050), .B1(G294), .B2(new_n818), .ZN(new_n1051));
  INV_X1    g0851(.A(G317), .ZN(new_n1052));
  OAI221_X1 g0852(.A(new_n282), .B1(new_n825), .B2(new_n1052), .C1(new_n479), .C2(new_n829), .ZN(new_n1053));
  NAND2_X1  g0853(.A1(new_n1053), .A2(KEYINPUT108), .ZN(new_n1054));
  OR2_X1    g0854(.A1(new_n1053), .A2(KEYINPUT108), .ZN(new_n1055));
  NAND3_X1  g0855(.A1(new_n1051), .A2(new_n1054), .A3(new_n1055), .ZN(new_n1056));
  OAI21_X1  g0856(.A(new_n1046), .B1(new_n1049), .B2(new_n1056), .ZN(new_n1057));
  XNOR2_X1  g0857(.A(new_n1057), .B(KEYINPUT47), .ZN(new_n1058));
  AOI21_X1  g0858(.A(new_n1035), .B1(new_n1058), .B2(new_n804), .ZN(new_n1059));
  OAI21_X1  g0859(.A(new_n1059), .B1(new_n852), .B2(new_n1006), .ZN(new_n1060));
  NAND2_X1  g0860(.A1(new_n1032), .A2(new_n1060), .ZN(G387));
  OR2_X1    g0861(.A1(new_n743), .A2(new_n852), .ZN(new_n1062));
  INV_X1    g0862(.A(new_n791), .ZN(new_n1063));
  NOR2_X1   g0863(.A1(new_n240), .A2(new_n431), .ZN(new_n1064));
  INV_X1    g0864(.A(new_n339), .ZN(new_n1065));
  AND3_X1   g0865(.A1(new_n1065), .A2(KEYINPUT50), .A3(new_n220), .ZN(new_n1066));
  AOI21_X1  g0866(.A(KEYINPUT50), .B1(new_n1065), .B2(new_n220), .ZN(new_n1067));
  OR2_X1    g0867(.A1(new_n1066), .A2(new_n1067), .ZN(new_n1068));
  AOI211_X1 g0868(.A(G45), .B(new_n751), .C1(G68), .C2(G77), .ZN(new_n1069));
  AOI211_X1 g0869(.A(new_n797), .B(new_n1064), .C1(new_n1068), .C2(new_n1069), .ZN(new_n1070));
  INV_X1    g0870(.A(KEYINPUT109), .ZN(new_n1071));
  NAND3_X1  g0871(.A1(new_n212), .A2(new_n751), .A3(new_n268), .ZN(new_n1072));
  OAI21_X1  g0872(.A(new_n1072), .B1(G107), .B2(new_n212), .ZN(new_n1073));
  AOI21_X1  g0873(.A(new_n1070), .B1(new_n1071), .B2(new_n1073), .ZN(new_n1074));
  OAI21_X1  g0874(.A(new_n1074), .B1(new_n1071), .B2(new_n1073), .ZN(new_n1075));
  AND2_X1   g0875(.A1(new_n1075), .A2(new_n805), .ZN(new_n1076));
  NOR2_X1   g0876(.A1(new_n811), .A2(new_n341), .ZN(new_n1077));
  OAI22_X1  g0877(.A1(new_n839), .A2(new_n843), .B1(new_n829), .B2(new_n284), .ZN(new_n1078));
  AOI211_X1 g0878(.A(new_n1077), .B(new_n1078), .C1(new_n1065), .C2(new_n818), .ZN(new_n1079));
  NAND2_X1  g0879(.A1(new_n897), .A2(G77), .ZN(new_n1080));
  OAI211_X1 g0880(.A(new_n1080), .B(new_n268), .C1(new_n371), .C2(new_n825), .ZN(new_n1081));
  AOI21_X1  g0881(.A(new_n1081), .B1(new_n1040), .B2(G68), .ZN(new_n1082));
  OAI211_X1 g0882(.A(new_n1079), .B(new_n1082), .C1(new_n220), .C2(new_n833), .ZN(new_n1083));
  XNOR2_X1  g0883(.A(new_n1083), .B(KEYINPUT110), .ZN(new_n1084));
  AOI21_X1  g0884(.A(new_n268), .B1(new_n826), .B2(G326), .ZN(new_n1085));
  OAI22_X1  g0885(.A1(new_n811), .A2(new_n828), .B1(new_n813), .B2(new_n548), .ZN(new_n1086));
  AOI22_X1  g0886(.A1(new_n818), .A2(G311), .B1(new_n822), .B2(G322), .ZN(new_n1087));
  OAI221_X1 g0887(.A(new_n1087), .B1(new_n837), .B2(new_n814), .C1(new_n1052), .C2(new_n833), .ZN(new_n1088));
  INV_X1    g0888(.A(KEYINPUT48), .ZN(new_n1089));
  AOI21_X1  g0889(.A(new_n1086), .B1(new_n1088), .B2(new_n1089), .ZN(new_n1090));
  OAI21_X1  g0890(.A(new_n1090), .B1(new_n1089), .B2(new_n1088), .ZN(new_n1091));
  INV_X1    g0891(.A(KEYINPUT49), .ZN(new_n1092));
  OAI221_X1 g0892(.A(new_n1085), .B1(new_n470), .B2(new_n829), .C1(new_n1091), .C2(new_n1092), .ZN(new_n1093));
  AND2_X1   g0893(.A1(new_n1091), .A2(new_n1092), .ZN(new_n1094));
  OAI21_X1  g0894(.A(new_n1084), .B1(new_n1093), .B2(new_n1094), .ZN(new_n1095));
  AOI211_X1 g0895(.A(new_n1063), .B(new_n1076), .C1(new_n804), .C2(new_n1095), .ZN(new_n1096));
  AOI22_X1  g0896(.A1(new_n1062), .A2(new_n1096), .B1(new_n1027), .B2(new_n790), .ZN(new_n1097));
  NAND2_X1  g0897(.A1(new_n1028), .A2(new_n750), .ZN(new_n1098));
  NOR2_X1   g0898(.A1(new_n786), .A2(new_n1027), .ZN(new_n1099));
  OAI21_X1  g0899(.A(new_n1097), .B1(new_n1098), .B2(new_n1099), .ZN(G393));
  NAND2_X1  g0900(.A1(new_n744), .A2(KEYINPUT111), .ZN(new_n1101));
  NAND2_X1  g0901(.A1(new_n1022), .A2(new_n1101), .ZN(new_n1102));
  NOR2_X1   g0902(.A1(new_n744), .A2(KEYINPUT111), .ZN(new_n1103));
  NAND2_X1  g0903(.A1(new_n1102), .A2(new_n1103), .ZN(new_n1104));
  INV_X1    g0904(.A(new_n1103), .ZN(new_n1105));
  NAND3_X1  g0905(.A1(new_n1022), .A2(new_n1105), .A3(new_n1101), .ZN(new_n1106));
  NAND2_X1  g0906(.A1(new_n1104), .A2(new_n1106), .ZN(new_n1107));
  NAND2_X1  g0907(.A1(new_n1107), .A2(new_n790), .ZN(new_n1108));
  INV_X1    g0908(.A(KEYINPUT115), .ZN(new_n1109));
  OAI22_X1  g0909(.A1(new_n833), .A2(new_n836), .B1(new_n1052), .B2(new_n839), .ZN(new_n1110));
  XOR2_X1   g0910(.A(new_n1110), .B(KEYINPUT113), .Z(new_n1111));
  OR2_X1    g0911(.A1(new_n1111), .A2(KEYINPUT52), .ZN(new_n1112));
  NAND2_X1  g0912(.A1(new_n1111), .A2(KEYINPUT52), .ZN(new_n1113));
  OAI22_X1  g0913(.A1(new_n819), .A2(new_n814), .B1(new_n811), .B2(new_n470), .ZN(new_n1114));
  AOI21_X1  g0914(.A(new_n268), .B1(new_n826), .B2(G322), .ZN(new_n1115));
  OAI221_X1 g0915(.A(new_n1115), .B1(new_n352), .B2(new_n829), .C1(new_n837), .C2(new_n548), .ZN(new_n1116));
  AOI211_X1 g0916(.A(new_n1114), .B(new_n1116), .C1(G283), .C2(new_n897), .ZN(new_n1117));
  NAND3_X1  g0917(.A1(new_n1112), .A2(new_n1113), .A3(new_n1117), .ZN(new_n1118));
  AOI22_X1  g0918(.A1(new_n818), .A2(G50), .B1(new_n810), .B2(G77), .ZN(new_n1119));
  OAI21_X1  g0919(.A(new_n1119), .B1(new_n837), .B2(new_n339), .ZN(new_n1120));
  XOR2_X1   g0920(.A(new_n1120), .B(KEYINPUT112), .Z(new_n1121));
  OAI22_X1  g0921(.A1(new_n833), .A2(new_n843), .B1(new_n371), .B2(new_n839), .ZN(new_n1122));
  XNOR2_X1  g0922(.A(new_n1122), .B(KEYINPUT51), .ZN(new_n1123));
  OAI21_X1  g0923(.A(new_n268), .B1(new_n825), .B2(new_n881), .ZN(new_n1124));
  AOI211_X1 g0924(.A(new_n895), .B(new_n1124), .C1(G68), .C2(new_n897), .ZN(new_n1125));
  NAND3_X1  g0925(.A1(new_n1121), .A2(new_n1123), .A3(new_n1125), .ZN(new_n1126));
  AOI21_X1  g0926(.A(new_n849), .B1(new_n1118), .B2(new_n1126), .ZN(new_n1127));
  NAND2_X1  g0927(.A1(new_n249), .A2(new_n796), .ZN(new_n1128));
  NOR2_X1   g0928(.A1(new_n212), .A2(new_n479), .ZN(new_n1129));
  NOR2_X1   g0929(.A1(new_n1129), .A2(new_n806), .ZN(new_n1130));
  AOI211_X1 g0930(.A(new_n1063), .B(new_n1127), .C1(new_n1128), .C2(new_n1130), .ZN(new_n1131));
  XOR2_X1   g0931(.A(new_n1131), .B(KEYINPUT114), .Z(new_n1132));
  OR2_X1    g0932(.A1(new_n995), .A2(new_n852), .ZN(new_n1133));
  NAND2_X1  g0933(.A1(new_n1132), .A2(new_n1133), .ZN(new_n1134));
  NAND3_X1  g0934(.A1(new_n1108), .A2(new_n1109), .A3(new_n1134), .ZN(new_n1135));
  AOI21_X1  g0935(.A(new_n789), .B1(new_n1104), .B2(new_n1106), .ZN(new_n1136));
  INV_X1    g0936(.A(new_n1134), .ZN(new_n1137));
  OAI21_X1  g0937(.A(KEYINPUT115), .B1(new_n1136), .B2(new_n1137), .ZN(new_n1138));
  NAND2_X1  g0938(.A1(new_n1135), .A2(new_n1138), .ZN(new_n1139));
  OAI211_X1 g0939(.A(new_n1030), .B(new_n750), .C1(new_n1029), .C2(new_n1107), .ZN(new_n1140));
  NAND2_X1  g0940(.A1(new_n1139), .A2(new_n1140), .ZN(G390));
  INV_X1    g0941(.A(new_n875), .ZN(new_n1142));
  OAI21_X1  g0942(.A(new_n1142), .B1(new_n765), .B2(new_n766), .ZN(new_n1143));
  NAND3_X1  g0943(.A1(new_n980), .A2(new_n939), .A3(G330), .ZN(new_n1144));
  NAND3_X1  g0944(.A1(new_n785), .A2(G330), .A3(new_n866), .ZN(new_n1145));
  NAND2_X1  g0945(.A1(new_n1145), .A2(new_n940), .ZN(new_n1146));
  NAND4_X1  g0946(.A1(new_n1143), .A2(new_n957), .A3(new_n1144), .A4(new_n1146), .ZN(new_n1147));
  INV_X1    g0947(.A(new_n1144), .ZN(new_n1148));
  AOI21_X1  g0948(.A(new_n939), .B1(new_n980), .B2(G330), .ZN(new_n1149));
  OAI21_X1  g0949(.A(new_n958), .B1(new_n1148), .B2(new_n1149), .ZN(new_n1150));
  NAND2_X1  g0950(.A1(new_n1147), .A2(new_n1150), .ZN(new_n1151));
  AND3_X1   g0951(.A1(new_n469), .A2(new_n785), .A3(G330), .ZN(new_n1152));
  AOI211_X1 g0952(.A(new_n683), .B(new_n1152), .C1(new_n767), .C2(new_n976), .ZN(new_n1153));
  INV_X1    g0953(.A(KEYINPUT116), .ZN(new_n1154));
  AND3_X1   g0954(.A1(new_n1151), .A2(new_n1153), .A3(new_n1154), .ZN(new_n1155));
  AOI21_X1  g0955(.A(new_n1154), .B1(new_n1151), .B2(new_n1153), .ZN(new_n1156));
  NOR2_X1   g0956(.A1(new_n1155), .A2(new_n1156), .ZN(new_n1157));
  INV_X1    g0957(.A(new_n969), .ZN(new_n1158));
  INV_X1    g0958(.A(new_n970), .ZN(new_n1159));
  NOR2_X1   g0959(.A1(new_n933), .A2(new_n940), .ZN(new_n1160));
  OAI22_X1  g0960(.A1(new_n1158), .A2(new_n1159), .B1(new_n1160), .B2(new_n972), .ZN(new_n1161));
  AOI21_X1  g0961(.A(new_n940), .B1(new_n1143), .B2(new_n957), .ZN(new_n1162));
  OAI22_X1  g0962(.A1(new_n929), .A2(new_n968), .B1(new_n678), .B2(new_n735), .ZN(new_n1163));
  OAI21_X1  g0963(.A(new_n1161), .B1(new_n1162), .B2(new_n1163), .ZN(new_n1164));
  NAND2_X1  g0964(.A1(new_n1164), .A2(new_n1148), .ZN(new_n1165));
  OAI211_X1 g0965(.A(new_n1161), .B(new_n1144), .C1(new_n1162), .C2(new_n1163), .ZN(new_n1166));
  NAND2_X1  g0966(.A1(new_n1165), .A2(new_n1166), .ZN(new_n1167));
  NAND2_X1  g0967(.A1(new_n1157), .A2(new_n1167), .ZN(new_n1168));
  OAI211_X1 g0968(.A(new_n1165), .B(new_n1166), .C1(new_n1155), .C2(new_n1156), .ZN(new_n1169));
  NAND3_X1  g0969(.A1(new_n1168), .A2(new_n750), .A3(new_n1169), .ZN(new_n1170));
  INV_X1    g0970(.A(new_n1167), .ZN(new_n1171));
  OAI21_X1  g0971(.A(new_n801), .B1(new_n1158), .B2(new_n1159), .ZN(new_n1172));
  OAI21_X1  g0972(.A(new_n791), .B1(new_n1065), .B2(new_n877), .ZN(new_n1173));
  XOR2_X1   g0973(.A(KEYINPUT54), .B(G143), .Z(new_n1174));
  NAND2_X1  g0974(.A1(new_n1040), .A2(new_n1174), .ZN(new_n1175));
  NAND2_X1  g0975(.A1(new_n834), .A2(G132), .ZN(new_n1176));
  NAND2_X1  g0976(.A1(new_n1044), .A2(G50), .ZN(new_n1177));
  AOI21_X1  g0977(.A(new_n282), .B1(new_n826), .B2(G125), .ZN(new_n1178));
  NAND4_X1  g0978(.A1(new_n1175), .A2(new_n1176), .A3(new_n1177), .A4(new_n1178), .ZN(new_n1179));
  NOR2_X1   g0979(.A1(new_n813), .A2(new_n371), .ZN(new_n1180));
  XNOR2_X1  g0980(.A(new_n1180), .B(KEYINPUT53), .ZN(new_n1181));
  AOI22_X1  g0981(.A1(new_n822), .A2(G128), .B1(new_n810), .B2(G159), .ZN(new_n1182));
  OAI211_X1 g0982(.A(new_n1181), .B(new_n1182), .C1(new_n1042), .C2(new_n819), .ZN(new_n1183));
  AOI22_X1  g0983(.A1(G68), .A2(new_n1044), .B1(new_n810), .B2(G77), .ZN(new_n1184));
  OAI221_X1 g0984(.A(new_n1184), .B1(new_n839), .B2(new_n828), .C1(new_n352), .C2(new_n819), .ZN(new_n1185));
  OAI21_X1  g0985(.A(new_n282), .B1(new_n825), .B2(new_n548), .ZN(new_n1186));
  AOI21_X1  g0986(.A(new_n1186), .B1(G87), .B2(new_n897), .ZN(new_n1187));
  OAI221_X1 g0987(.A(new_n1187), .B1(new_n837), .B2(new_n479), .C1(new_n470), .C2(new_n833), .ZN(new_n1188));
  OAI22_X1  g0988(.A1(new_n1179), .A2(new_n1183), .B1(new_n1185), .B2(new_n1188), .ZN(new_n1189));
  AOI21_X1  g0989(.A(new_n1173), .B1(new_n1189), .B2(new_n804), .ZN(new_n1190));
  AOI22_X1  g0990(.A1(new_n1171), .A2(new_n790), .B1(new_n1172), .B2(new_n1190), .ZN(new_n1191));
  NAND2_X1  g0991(.A1(new_n1170), .A2(new_n1191), .ZN(G378));
  OAI21_X1  g0992(.A(new_n791), .B1(G50), .B2(new_n877), .ZN(new_n1193));
  OAI21_X1  g0993(.A(new_n377), .B1(new_n389), .B2(new_n384), .ZN(new_n1194));
  NAND2_X1  g0994(.A1(new_n376), .A2(new_n918), .ZN(new_n1195));
  INV_X1    g0995(.A(new_n1195), .ZN(new_n1196));
  AND2_X1   g0996(.A1(new_n1194), .A2(new_n1196), .ZN(new_n1197));
  NOR2_X1   g0997(.A1(new_n1194), .A2(new_n1196), .ZN(new_n1198));
  XNOR2_X1  g0998(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1199));
  INV_X1    g0999(.A(new_n1199), .ZN(new_n1200));
  OR3_X1    g1000(.A1(new_n1197), .A2(new_n1198), .A3(new_n1200), .ZN(new_n1201));
  OAI21_X1  g1001(.A(new_n1200), .B1(new_n1197), .B2(new_n1198), .ZN(new_n1202));
  AND2_X1   g1002(.A1(new_n1201), .A2(new_n1202), .ZN(new_n1203));
  INV_X1    g1003(.A(new_n1203), .ZN(new_n1204));
  NOR2_X1   g1004(.A1(new_n1204), .A2(new_n802), .ZN(new_n1205));
  NOR2_X1   g1005(.A1(new_n268), .A2(G41), .ZN(new_n1206));
  AOI211_X1 g1006(.A(G50), .B(new_n1206), .C1(new_n283), .C2(new_n430), .ZN(new_n1207));
  XNOR2_X1  g1007(.A(new_n1207), .B(KEYINPUT117), .ZN(new_n1208));
  AOI22_X1  g1008(.A1(new_n1040), .A2(new_n621), .B1(new_n834), .B2(G107), .ZN(new_n1209));
  NAND2_X1  g1009(.A1(new_n1044), .A2(G58), .ZN(new_n1210));
  NAND2_X1  g1010(.A1(new_n826), .A2(G283), .ZN(new_n1211));
  NAND4_X1  g1011(.A1(new_n1080), .A2(new_n1210), .A3(new_n1206), .A4(new_n1211), .ZN(new_n1212));
  XOR2_X1   g1012(.A(new_n1212), .B(KEYINPUT118), .Z(new_n1213));
  NAND2_X1  g1013(.A1(new_n818), .A2(G97), .ZN(new_n1214));
  AOI21_X1  g1014(.A(new_n1036), .B1(G116), .B2(new_n822), .ZN(new_n1215));
  NAND4_X1  g1015(.A1(new_n1209), .A2(new_n1213), .A3(new_n1214), .A4(new_n1215), .ZN(new_n1216));
  INV_X1    g1016(.A(KEYINPUT58), .ZN(new_n1217));
  AOI21_X1  g1017(.A(new_n1208), .B1(new_n1216), .B2(new_n1217), .ZN(new_n1218));
  NAND2_X1  g1018(.A1(new_n834), .A2(G128), .ZN(new_n1219));
  NAND2_X1  g1019(.A1(new_n1040), .A2(G137), .ZN(new_n1220));
  AOI22_X1  g1020(.A1(new_n822), .A2(G125), .B1(new_n810), .B2(G150), .ZN(new_n1221));
  AOI22_X1  g1021(.A1(new_n818), .A2(G132), .B1(new_n897), .B2(new_n1174), .ZN(new_n1222));
  NAND4_X1  g1022(.A1(new_n1219), .A2(new_n1220), .A3(new_n1221), .A4(new_n1222), .ZN(new_n1223));
  XOR2_X1   g1023(.A(new_n1223), .B(KEYINPUT119), .Z(new_n1224));
  NAND2_X1  g1024(.A1(new_n1224), .A2(KEYINPUT59), .ZN(new_n1225));
  AOI211_X1 g1025(.A(G33), .B(G41), .C1(new_n826), .C2(G124), .ZN(new_n1226));
  OAI211_X1 g1026(.A(new_n1225), .B(new_n1226), .C1(new_n843), .C2(new_n829), .ZN(new_n1227));
  NOR2_X1   g1027(.A1(new_n1224), .A2(KEYINPUT59), .ZN(new_n1228));
  OAI221_X1 g1028(.A(new_n1218), .B1(new_n1217), .B2(new_n1216), .C1(new_n1227), .C2(new_n1228), .ZN(new_n1229));
  AOI211_X1 g1029(.A(new_n1193), .B(new_n1205), .C1(new_n804), .C2(new_n1229), .ZN(new_n1230));
  INV_X1    g1030(.A(KEYINPUT120), .ZN(new_n1231));
  AOI21_X1  g1031(.A(new_n1204), .B1(new_n985), .B2(G330), .ZN(new_n1232));
  AOI211_X1 g1032(.A(new_n979), .B(new_n1203), .C1(new_n982), .C2(new_n984), .ZN(new_n1233));
  NOR3_X1   g1033(.A1(new_n974), .A2(new_n1232), .A3(new_n1233), .ZN(new_n1234));
  NAND3_X1  g1034(.A1(new_n985), .A2(G330), .A3(new_n1204), .ZN(new_n1235));
  AOI21_X1  g1035(.A(KEYINPUT40), .B1(new_n947), .B2(new_n948), .ZN(new_n1236));
  AND2_X1   g1036(.A1(new_n980), .A2(new_n939), .ZN(new_n1237));
  AOI22_X1  g1037(.A1(KEYINPUT40), .A2(new_n981), .B1(new_n1236), .B2(new_n1237), .ZN(new_n1238));
  OAI21_X1  g1038(.A(new_n1203), .B1(new_n1238), .B2(new_n979), .ZN(new_n1239));
  NAND2_X1  g1039(.A1(new_n959), .A2(new_n942), .ZN(new_n1240));
  AOI22_X1  g1040(.A1(new_n1240), .A2(KEYINPUT103), .B1(new_n971), .B2(new_n972), .ZN(new_n1241));
  AOI22_X1  g1041(.A1(new_n1235), .A2(new_n1239), .B1(new_n1241), .B2(new_n961), .ZN(new_n1242));
  OAI21_X1  g1042(.A(new_n1231), .B1(new_n1234), .B2(new_n1242), .ZN(new_n1243));
  OAI21_X1  g1043(.A(new_n974), .B1(new_n1232), .B2(new_n1233), .ZN(new_n1244));
  NAND4_X1  g1044(.A1(new_n1239), .A2(new_n1241), .A3(new_n1235), .A4(new_n961), .ZN(new_n1245));
  NAND3_X1  g1045(.A1(new_n1244), .A2(new_n1245), .A3(KEYINPUT120), .ZN(new_n1246));
  AND2_X1   g1046(.A1(new_n1243), .A2(new_n1246), .ZN(new_n1247));
  AOI21_X1  g1047(.A(new_n1230), .B1(new_n1247), .B2(new_n790), .ZN(new_n1248));
  OAI21_X1  g1048(.A(new_n1153), .B1(new_n1157), .B2(new_n1167), .ZN(new_n1249));
  AOI21_X1  g1049(.A(KEYINPUT57), .B1(new_n1247), .B2(new_n1249), .ZN(new_n1250));
  NAND2_X1  g1050(.A1(new_n1244), .A2(new_n1245), .ZN(new_n1251));
  NAND3_X1  g1051(.A1(new_n1249), .A2(KEYINPUT57), .A3(new_n1251), .ZN(new_n1252));
  NAND2_X1  g1052(.A1(new_n1252), .A2(new_n750), .ZN(new_n1253));
  OAI21_X1  g1053(.A(new_n1248), .B1(new_n1250), .B2(new_n1253), .ZN(G375));
  NAND2_X1  g1054(.A1(new_n940), .A2(new_n801), .ZN(new_n1255));
  OAI21_X1  g1055(.A(new_n791), .B1(G68), .B2(new_n877), .ZN(new_n1256));
  OAI22_X1  g1056(.A1(new_n819), .A2(new_n470), .B1(new_n839), .B2(new_n548), .ZN(new_n1257));
  AOI211_X1 g1057(.A(new_n1077), .B(new_n1257), .C1(G97), .C2(new_n897), .ZN(new_n1258));
  OAI221_X1 g1058(.A(new_n282), .B1(new_n825), .B2(new_n814), .C1(new_n225), .C2(new_n829), .ZN(new_n1259));
  AOI21_X1  g1059(.A(new_n1259), .B1(new_n1040), .B2(G107), .ZN(new_n1260));
  OAI211_X1 g1060(.A(new_n1258), .B(new_n1260), .C1(new_n828), .C2(new_n833), .ZN(new_n1261));
  NAND2_X1  g1061(.A1(new_n1210), .A2(new_n268), .ZN(new_n1262));
  XNOR2_X1  g1062(.A(new_n1262), .B(KEYINPUT121), .ZN(new_n1263));
  NAND2_X1  g1063(.A1(new_n826), .A2(G128), .ZN(new_n1264));
  OAI21_X1  g1064(.A(new_n1264), .B1(new_n811), .B2(new_n220), .ZN(new_n1265));
  AOI21_X1  g1065(.A(new_n1265), .B1(G159), .B2(new_n897), .ZN(new_n1266));
  OAI211_X1 g1066(.A(new_n1263), .B(new_n1266), .C1(new_n371), .C2(new_n837), .ZN(new_n1267));
  XOR2_X1   g1067(.A(new_n1267), .B(KEYINPUT122), .Z(new_n1268));
  AOI22_X1  g1068(.A1(G132), .A2(new_n822), .B1(new_n818), .B2(new_n1174), .ZN(new_n1269));
  OAI21_X1  g1069(.A(new_n1269), .B1(new_n833), .B2(new_n1042), .ZN(new_n1270));
  OAI21_X1  g1070(.A(new_n1261), .B1(new_n1268), .B2(new_n1270), .ZN(new_n1271));
  AOI21_X1  g1071(.A(new_n1256), .B1(new_n1271), .B2(new_n804), .ZN(new_n1272));
  AOI22_X1  g1072(.A1(new_n1151), .A2(new_n790), .B1(new_n1255), .B2(new_n1272), .ZN(new_n1273));
  OR2_X1    g1073(.A1(new_n1151), .A2(new_n1153), .ZN(new_n1274));
  NAND2_X1  g1074(.A1(new_n1157), .A2(new_n1274), .ZN(new_n1275));
  OAI21_X1  g1075(.A(new_n1273), .B1(new_n1275), .B2(new_n1017), .ZN(G381));
  INV_X1    g1076(.A(G390), .ZN(new_n1277));
  NOR3_X1   g1077(.A1(G393), .A2(G384), .A3(G396), .ZN(new_n1278));
  NAND4_X1  g1078(.A1(new_n1277), .A2(new_n1060), .A3(new_n1032), .A4(new_n1278), .ZN(new_n1279));
  OR4_X1    g1079(.A1(G378), .A2(new_n1279), .A3(G375), .A4(G381), .ZN(G407));
  INV_X1    g1080(.A(G378), .ZN(new_n1281));
  NAND2_X1  g1081(.A1(new_n734), .A2(G213), .ZN(new_n1282));
  INV_X1    g1082(.A(new_n1282), .ZN(new_n1283));
  NAND2_X1  g1083(.A1(new_n1281), .A2(new_n1283), .ZN(new_n1284));
  OAI211_X1 g1084(.A(G407), .B(G213), .C1(G375), .C2(new_n1284), .ZN(G409));
  XOR2_X1   g1085(.A(G393), .B(G396), .Z(new_n1286));
  INV_X1    g1086(.A(new_n1286), .ZN(new_n1287));
  AND3_X1   g1087(.A1(new_n1032), .A2(G390), .A3(new_n1060), .ZN(new_n1288));
  AOI21_X1  g1088(.A(G390), .B1(new_n1032), .B2(new_n1060), .ZN(new_n1289));
  OAI21_X1  g1089(.A(new_n1287), .B1(new_n1288), .B2(new_n1289), .ZN(new_n1290));
  NAND2_X1  g1090(.A1(G387), .A2(new_n1277), .ZN(new_n1291));
  NAND3_X1  g1091(.A1(new_n1032), .A2(G390), .A3(new_n1060), .ZN(new_n1292));
  NAND3_X1  g1092(.A1(new_n1291), .A2(new_n1286), .A3(new_n1292), .ZN(new_n1293));
  NAND2_X1  g1093(.A1(new_n1290), .A2(new_n1293), .ZN(new_n1294));
  INV_X1    g1094(.A(KEYINPUT61), .ZN(new_n1295));
  INV_X1    g1095(.A(new_n1017), .ZN(new_n1296));
  NAND4_X1  g1096(.A1(new_n1249), .A2(new_n1296), .A3(new_n1243), .A4(new_n1246), .ZN(new_n1297));
  NAND2_X1  g1097(.A1(new_n1297), .A2(KEYINPUT123), .ZN(new_n1298));
  AOI21_X1  g1098(.A(new_n1017), .B1(new_n1169), .B2(new_n1153), .ZN(new_n1299));
  INV_X1    g1099(.A(KEYINPUT123), .ZN(new_n1300));
  NAND4_X1  g1100(.A1(new_n1299), .A2(new_n1300), .A3(new_n1246), .A4(new_n1243), .ZN(new_n1301));
  INV_X1    g1101(.A(KEYINPUT124), .ZN(new_n1302));
  AOI21_X1  g1102(.A(new_n789), .B1(new_n1251), .B2(new_n1302), .ZN(new_n1303));
  NAND3_X1  g1103(.A1(new_n1244), .A2(new_n1245), .A3(KEYINPUT124), .ZN(new_n1304));
  AOI21_X1  g1104(.A(new_n1230), .B1(new_n1303), .B2(new_n1304), .ZN(new_n1305));
  NAND3_X1  g1105(.A1(new_n1298), .A2(new_n1301), .A3(new_n1305), .ZN(new_n1306));
  NAND2_X1  g1106(.A1(new_n1306), .A2(new_n1281), .ZN(new_n1307));
  OAI211_X1 g1107(.A(G378), .B(new_n1248), .C1(new_n1250), .C2(new_n1253), .ZN(new_n1308));
  AOI21_X1  g1108(.A(new_n1283), .B1(new_n1307), .B2(new_n1308), .ZN(new_n1309));
  NAND2_X1  g1109(.A1(new_n1283), .A2(G2897), .ZN(new_n1310));
  INV_X1    g1110(.A(new_n1310), .ZN(new_n1311));
  INV_X1    g1111(.A(KEYINPUT60), .ZN(new_n1312));
  NAND2_X1  g1112(.A1(new_n1274), .A2(new_n1312), .ZN(new_n1313));
  NAND2_X1  g1113(.A1(new_n1313), .A2(new_n750), .ZN(new_n1314));
  AOI21_X1  g1114(.A(new_n1314), .B1(new_n1275), .B2(KEYINPUT60), .ZN(new_n1315));
  INV_X1    g1115(.A(new_n1273), .ZN(new_n1316));
  OAI21_X1  g1116(.A(new_n902), .B1(new_n1315), .B2(new_n1316), .ZN(new_n1317));
  INV_X1    g1117(.A(new_n1317), .ZN(new_n1318));
  NOR3_X1   g1118(.A1(new_n1315), .A2(new_n902), .A3(new_n1316), .ZN(new_n1319));
  OAI21_X1  g1119(.A(new_n1311), .B1(new_n1318), .B2(new_n1319), .ZN(new_n1320));
  INV_X1    g1120(.A(new_n1319), .ZN(new_n1321));
  NAND3_X1  g1121(.A1(new_n1321), .A2(new_n1317), .A3(new_n1310), .ZN(new_n1322));
  NAND2_X1  g1122(.A1(new_n1320), .A2(new_n1322), .ZN(new_n1323));
  OAI21_X1  g1123(.A(new_n1295), .B1(new_n1309), .B2(new_n1323), .ZN(new_n1324));
  INV_X1    g1124(.A(KEYINPUT125), .ZN(new_n1325));
  NAND2_X1  g1125(.A1(new_n1324), .A2(new_n1325), .ZN(new_n1326));
  OAI211_X1 g1126(.A(KEYINPUT125), .B(new_n1295), .C1(new_n1309), .C2(new_n1323), .ZN(new_n1327));
  NAND2_X1  g1127(.A1(new_n1326), .A2(new_n1327), .ZN(new_n1328));
  NAND2_X1  g1128(.A1(new_n1307), .A2(new_n1308), .ZN(new_n1329));
  NOR2_X1   g1129(.A1(new_n1318), .A2(new_n1319), .ZN(new_n1330));
  OR2_X1    g1130(.A1(KEYINPUT126), .A2(KEYINPUT62), .ZN(new_n1331));
  NAND4_X1  g1131(.A1(new_n1329), .A2(new_n1282), .A3(new_n1330), .A4(new_n1331), .ZN(new_n1332));
  NAND2_X1  g1132(.A1(KEYINPUT126), .A2(KEYINPUT62), .ZN(new_n1333));
  NAND2_X1  g1133(.A1(new_n1332), .A2(new_n1333), .ZN(new_n1334));
  AOI21_X1  g1134(.A(new_n1331), .B1(new_n1309), .B2(new_n1330), .ZN(new_n1335));
  NOR2_X1   g1135(.A1(new_n1334), .A2(new_n1335), .ZN(new_n1336));
  OAI21_X1  g1136(.A(new_n1294), .B1(new_n1328), .B2(new_n1336), .ZN(new_n1337));
  NAND2_X1  g1137(.A1(new_n1309), .A2(new_n1330), .ZN(new_n1338));
  XNOR2_X1  g1138(.A(new_n1338), .B(KEYINPUT63), .ZN(new_n1339));
  AND2_X1   g1139(.A1(new_n1290), .A2(new_n1293), .ZN(new_n1340));
  INV_X1    g1140(.A(new_n1324), .ZN(new_n1341));
  NAND3_X1  g1141(.A1(new_n1339), .A2(new_n1340), .A3(new_n1341), .ZN(new_n1342));
  NAND2_X1  g1142(.A1(new_n1337), .A2(new_n1342), .ZN(G405));
  XNOR2_X1  g1143(.A(G375), .B(G378), .ZN(new_n1344));
  INV_X1    g1144(.A(new_n1330), .ZN(new_n1345));
  XNOR2_X1  g1145(.A(new_n1344), .B(new_n1345), .ZN(new_n1346));
  XNOR2_X1  g1146(.A(new_n1346), .B(new_n1294), .ZN(G402));
endmodule


