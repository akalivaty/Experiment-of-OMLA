

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
         n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
         n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
         n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
         n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410,
         n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421,
         n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432,
         n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443,
         n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454,
         n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465,
         n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
         n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487,
         n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
         n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
         n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586,
         n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597,
         n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608,
         n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619,
         n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630,
         n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641,
         n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652,
         n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663,
         n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674,
         n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685,
         n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696,
         n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707,
         n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718,
         n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729,
         n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, n740,
         n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, n751,
         n752, n753, n754, n755, n756, n757, n758, n759, n760, n761, n762,
         n763, n764, n765, n766, n767, n768, n769, n770, n771, n772, n773,
         n774, n775, n776, n777, n778, n779, n780, n781, n782, n783, n784,
         n785, n786, n787, n788, n789, n790, n791, n792, n793, n794, n795,
         n796, n797;

  BUF_X1 U379 ( .A(G116), .Z(n356) );
  XOR2_X1 U380 ( .A(n773), .B(n520), .Z(n542) );
  INV_X1 U381 ( .A(G953), .ZN(n783) );
  XNOR2_X1 U382 ( .A(G119), .B(KEYINPUT3), .ZN(n505) );
  XNOR2_X2 U383 ( .A(n517), .B(n516), .ZN(n518) );
  NAND2_X2 U384 ( .A1(n651), .A2(n535), .ZN(n537) );
  AND2_X1 U385 ( .A1(n383), .A2(n616), .ZN(n357) );
  AND2_X2 U386 ( .A1(n456), .A2(n458), .ZN(n455) );
  AND2_X2 U387 ( .A1(n381), .A2(n357), .ZN(n379) );
  XNOR2_X2 U388 ( .A(n545), .B(n544), .ZN(n640) );
  XNOR2_X2 U389 ( .A(n781), .B(n543), .ZN(n756) );
  NOR2_X1 U390 ( .A1(n765), .A2(KEYINPUT2), .ZN(n686) );
  NAND2_X1 U391 ( .A1(n379), .A2(n378), .ZN(n617) );
  INV_X4 U392 ( .A(G116), .ZN(n462) );
  NAND2_X1 U393 ( .A1(n404), .A2(n402), .ZN(n463) );
  NAND2_X1 U394 ( .A1(n403), .A2(n367), .ZN(n402) );
  AND2_X1 U395 ( .A1(n405), .A2(n369), .ZN(n404) );
  NAND2_X1 U396 ( .A1(n470), .A2(n674), .ZN(n469) );
  XNOR2_X1 U397 ( .A(n654), .B(n653), .ZN(n742) );
  XNOR2_X1 U398 ( .A(n408), .B(n407), .ZN(n797) );
  AND2_X1 U399 ( .A1(n485), .A2(n481), .ZN(n480) );
  NAND2_X1 U400 ( .A1(n454), .A2(n457), .ZN(n453) );
  BUF_X1 U401 ( .A(n599), .Z(n706) );
  XNOR2_X1 U402 ( .A(n578), .B(G478), .ZN(n603) );
  XNOR2_X1 U403 ( .A(n563), .B(G472), .ZN(n564) );
  NOR2_X1 U404 ( .A1(n528), .A2(n359), .ZN(n457) );
  XNOR2_X2 U405 ( .A(n462), .B(G113), .ZN(n461) );
  XNOR2_X2 U406 ( .A(n648), .B(KEYINPUT19), .ZN(n651) );
  NAND2_X2 U407 ( .A1(n659), .A2(n694), .ZN(n648) );
  XNOR2_X2 U408 ( .A(n569), .B(n584), .ZN(n538) );
  XNOR2_X2 U409 ( .A(n511), .B(n434), .ZN(n569) );
  XNOR2_X2 U410 ( .A(n425), .B(n460), .ZN(n494) );
  XNOR2_X2 U411 ( .A(n538), .B(n552), .ZN(n781) );
  XNOR2_X2 U412 ( .A(n461), .B(n505), .ZN(n425) );
  XNOR2_X2 U413 ( .A(n432), .B(n605), .ZN(n725) );
  NAND2_X1 U414 ( .A1(n737), .A2(n796), .ZN(n380) );
  XNOR2_X1 U415 ( .A(n414), .B(KEYINPUT67), .ZN(n552) );
  INV_X1 U416 ( .A(G137), .ZN(n414) );
  NAND2_X1 U417 ( .A1(n524), .A2(n523), .ZN(n546) );
  NAND2_X1 U418 ( .A1(n639), .A2(KEYINPUT28), .ZN(n442) );
  AND2_X1 U419 ( .A1(n424), .A2(n446), .ZN(n443) );
  XNOR2_X1 U420 ( .A(KEYINPUT66), .B(G131), .ZN(n584) );
  NOR2_X1 U421 ( .A1(n449), .A2(n504), .ZN(n666) );
  INV_X1 U422 ( .A(KEYINPUT48), .ZN(n474) );
  NAND2_X1 U423 ( .A1(n384), .A2(KEYINPUT84), .ZN(n383) );
  OR2_X2 U424 ( .A1(n793), .A2(n606), .ZN(n607) );
  INV_X1 U425 ( .A(G122), .ZN(n460) );
  INV_X1 U426 ( .A(G134), .ZN(n434) );
  XNOR2_X1 U427 ( .A(n468), .B(KEYINPUT65), .ZN(n520) );
  XNOR2_X1 U428 ( .A(KEYINPUT4), .B(G101), .ZN(n468) );
  NAND2_X1 U429 ( .A1(n604), .A2(n645), .ZN(n432) );
  NOR2_X1 U430 ( .A1(n704), .A2(n703), .ZN(n604) );
  XNOR2_X1 U431 ( .A(n564), .B(n437), .ZN(n636) );
  INV_X1 U432 ( .A(KEYINPUT106), .ZN(n437) );
  XNOR2_X1 U433 ( .A(n564), .B(KEYINPUT6), .ZN(n645) );
  XNOR2_X1 U434 ( .A(n490), .B(n489), .ZN(n599) );
  XNOR2_X1 U435 ( .A(n556), .B(n362), .ZN(n489) );
  OR2_X1 U436 ( .A1(n762), .A2(G902), .ZN(n490) );
  XNOR2_X1 U437 ( .A(n640), .B(KEYINPUT1), .ZN(n704) );
  XNOR2_X1 U438 ( .A(n416), .B(n548), .ZN(n415) );
  XNOR2_X1 U439 ( .A(n547), .B(KEYINPUT23), .ZN(n416) );
  XNOR2_X1 U440 ( .A(n549), .B(n552), .ZN(n413) );
  XNOR2_X1 U441 ( .A(KEYINPUT10), .B(G140), .ZN(n418) );
  XOR2_X1 U442 ( .A(KEYINPUT102), .B(G107), .Z(n574) );
  XNOR2_X1 U443 ( .A(n356), .B(G122), .ZN(n573) );
  NAND2_X1 U444 ( .A1(n676), .A2(n675), .ZN(n397) );
  NOR2_X1 U445 ( .A1(n360), .A2(n469), .ZN(n410) );
  INV_X1 U446 ( .A(n728), .ZN(n430) );
  INV_X1 U447 ( .A(KEYINPUT121), .ZN(n429) );
  XNOR2_X1 U448 ( .A(n635), .B(n634), .ZN(n724) );
  NAND2_X1 U449 ( .A1(n660), .A2(n486), .ZN(n485) );
  NOR2_X1 U450 ( .A1(n482), .A2(n744), .ZN(n481) );
  NAND2_X1 U451 ( .A1(n478), .A2(n483), .ZN(n479) );
  NAND2_X1 U452 ( .A1(n636), .A2(n445), .ZN(n444) );
  NOR2_X1 U453 ( .A1(n643), .A2(KEYINPUT28), .ZN(n445) );
  NAND2_X1 U454 ( .A1(n442), .A2(n652), .ZN(n440) );
  XNOR2_X1 U455 ( .A(KEYINPUT87), .B(KEYINPUT0), .ZN(n536) );
  INV_X1 U456 ( .A(n645), .ZN(n426) );
  BUF_X1 U457 ( .A(n704), .Z(n433) );
  NAND2_X1 U458 ( .A1(n396), .A2(G475), .ZN(n423) );
  AND2_X2 U459 ( .A1(n459), .A2(n397), .ZN(n396) );
  AND2_X1 U460 ( .A1(n691), .A2(n528), .ZN(n459) );
  NAND2_X1 U461 ( .A1(n396), .A2(G210), .ZN(n392) );
  NOR2_X1 U462 ( .A1(n709), .A2(n438), .ZN(n710) );
  NAND2_X1 U463 ( .A1(n528), .A2(n359), .ZN(n458) );
  XNOR2_X1 U464 ( .A(G122), .B(G143), .ZN(n581) );
  XOR2_X1 U465 ( .A(G104), .B(G113), .Z(n582) );
  XNOR2_X1 U466 ( .A(G902), .B(KEYINPUT15), .ZN(n527) );
  XOR2_X1 U467 ( .A(KEYINPUT89), .B(KEYINPUT17), .Z(n515) );
  NAND2_X1 U468 ( .A1(n496), .A2(n495), .ZN(n493) );
  OR2_X1 U469 ( .A1(n666), .A2(n474), .ZN(n470) );
  OR2_X1 U470 ( .A1(n475), .A2(n474), .ZN(n473) );
  NOR2_X1 U471 ( .A1(G237), .A2(G902), .ZN(n529) );
  NOR2_X1 U472 ( .A1(n637), .A2(n627), .ZN(n628) );
  NAND2_X1 U473 ( .A1(G237), .A2(G234), .ZN(n531) );
  XNOR2_X1 U474 ( .A(n406), .B(n509), .ZN(n561) );
  XNOR2_X1 U475 ( .A(n448), .B(n447), .ZN(n406) );
  XNOR2_X1 U476 ( .A(n520), .B(n503), .ZN(n447) );
  NAND2_X1 U477 ( .A1(n361), .A2(n409), .ZN(n436) );
  NOR2_X1 U478 ( .A1(n469), .A2(n411), .ZN(n409) );
  INV_X1 U479 ( .A(n753), .ZN(n411) );
  XNOR2_X1 U480 ( .A(n398), .B(G110), .ZN(n773) );
  XNOR2_X1 U481 ( .A(G107), .B(G104), .ZN(n398) );
  XOR2_X1 U482 ( .A(G146), .B(G140), .Z(n540) );
  NOR2_X1 U483 ( .A1(n680), .A2(n562), .ZN(n477) );
  XNOR2_X1 U484 ( .A(n417), .B(n412), .ZN(n762) );
  XNOR2_X1 U485 ( .A(n553), .B(n779), .ZN(n417) );
  XNOR2_X1 U486 ( .A(n415), .B(n413), .ZN(n412) );
  XNOR2_X1 U487 ( .A(n577), .B(n576), .ZN(n759) );
  XNOR2_X1 U488 ( .A(n575), .B(n502), .ZN(n576) );
  NAND2_X1 U489 ( .A1(n430), .A2(n429), .ZN(n428) );
  INV_X1 U490 ( .A(KEYINPUT42), .ZN(n407) );
  NAND2_X1 U491 ( .A1(n724), .A2(n366), .ZN(n408) );
  XNOR2_X1 U492 ( .A(n488), .B(n487), .ZN(n792) );
  INV_X1 U493 ( .A(KEYINPUT40), .ZN(n487) );
  INV_X1 U494 ( .A(KEYINPUT35), .ZN(n464) );
  AND2_X1 U495 ( .A1(n610), .A2(n426), .ZN(n387) );
  INV_X1 U496 ( .A(KEYINPUT31), .ZN(n376) );
  INV_X1 U497 ( .A(n712), .ZN(n431) );
  INV_X1 U498 ( .A(KEYINPUT75), .ZN(n653) );
  NOR2_X1 U499 ( .A1(n441), .A2(n440), .ZN(n439) );
  AND2_X1 U500 ( .A1(n626), .A2(n564), .ZN(n565) );
  NAND2_X1 U501 ( .A1(n427), .A2(n393), .ZN(n729) );
  AND2_X1 U502 ( .A1(n600), .A2(n426), .ZN(n393) );
  INV_X1 U503 ( .A(KEYINPUT60), .ZN(n419) );
  XNOR2_X1 U504 ( .A(n423), .B(n373), .ZN(n422) );
  AND2_X1 U505 ( .A1(n399), .A2(n421), .ZN(G54) );
  XNOR2_X1 U506 ( .A(n401), .B(n400), .ZN(n399) );
  XNOR2_X1 U507 ( .A(n756), .B(n374), .ZN(n400) );
  INV_X1 U508 ( .A(KEYINPUT56), .ZN(n389) );
  XNOR2_X1 U509 ( .A(n392), .B(n372), .ZN(n391) );
  OR2_X1 U510 ( .A1(n742), .A2(n698), .ZN(n358) );
  AND2_X1 U511 ( .A1(G210), .A2(n530), .ZN(n359) );
  XNOR2_X1 U512 ( .A(KEYINPUT76), .B(n677), .ZN(n360) );
  AND2_X1 U513 ( .A1(n473), .A2(n471), .ZN(n361) );
  XOR2_X1 U514 ( .A(n558), .B(n557), .Z(n362) );
  AND2_X1 U515 ( .A1(n436), .A2(n675), .ZN(n363) );
  AND2_X1 U516 ( .A1(n691), .A2(n429), .ZN(n364) );
  AND2_X1 U517 ( .A1(n443), .A2(n442), .ZN(n365) );
  AND2_X1 U518 ( .A1(n365), .A2(n444), .ZN(n366) );
  AND2_X1 U519 ( .A1(n728), .A2(KEYINPUT121), .ZN(n367) );
  AND2_X1 U520 ( .A1(n485), .A2(n484), .ZN(n368) );
  AND2_X1 U521 ( .A1(n428), .A2(n783), .ZN(n369) );
  XOR2_X1 U522 ( .A(KEYINPUT64), .B(KEYINPUT22), .Z(n370) );
  XOR2_X1 U523 ( .A(KEYINPUT74), .B(KEYINPUT34), .Z(n371) );
  XOR2_X1 U524 ( .A(n754), .B(n755), .Z(n372) );
  XNOR2_X1 U525 ( .A(n757), .B(KEYINPUT59), .ZN(n373) );
  INV_X1 U526 ( .A(KEYINPUT84), .ZN(n614) );
  XNOR2_X1 U527 ( .A(n546), .B(n418), .ZN(n779) );
  XNOR2_X1 U528 ( .A(KEYINPUT57), .B(KEYINPUT58), .ZN(n374) );
  INV_X1 U529 ( .A(G472), .ZN(n562) );
  NOR2_X1 U530 ( .A1(n683), .A2(n764), .ZN(n685) );
  INV_X1 U531 ( .A(n764), .ZN(n421) );
  XNOR2_X2 U532 ( .A(n465), .B(n464), .ZN(n793) );
  XNOR2_X2 U533 ( .A(n375), .B(KEYINPUT96), .ZN(n732) );
  NAND2_X1 U534 ( .A1(n388), .A2(n565), .ZN(n375) );
  XNOR2_X2 U535 ( .A(n377), .B(n376), .ZN(n747) );
  NAND2_X1 U536 ( .A1(n388), .A2(n431), .ZN(n377) );
  NAND2_X1 U537 ( .A1(n422), .A2(n421), .ZN(n420) );
  OR2_X1 U538 ( .A1(n385), .A2(n614), .ZN(n378) );
  XNOR2_X1 U539 ( .A(n609), .B(KEYINPUT85), .ZN(n385) );
  NAND2_X1 U540 ( .A1(n380), .A2(KEYINPUT44), .ZN(n613) );
  NOR2_X1 U541 ( .A1(n380), .A2(KEYINPUT44), .ZN(n615) );
  NAND2_X1 U542 ( .A1(n385), .A2(n382), .ZN(n381) );
  AND2_X1 U543 ( .A1(n613), .A2(n614), .ZN(n382) );
  INV_X1 U544 ( .A(n613), .ZN(n384) );
  XNOR2_X2 U545 ( .A(n386), .B(KEYINPUT32), .ZN(n796) );
  NAND2_X1 U546 ( .A1(n427), .A2(n387), .ZN(n386) );
  NAND2_X1 U547 ( .A1(n388), .A2(n725), .ZN(n467) );
  NAND2_X1 U548 ( .A1(n388), .A2(n597), .ZN(n598) );
  XNOR2_X2 U549 ( .A(n537), .B(n536), .ZN(n388) );
  XNOR2_X1 U550 ( .A(n390), .B(n389), .ZN(G51) );
  NAND2_X1 U551 ( .A1(n391), .A2(n421), .ZN(n390) );
  XNOR2_X2 U552 ( .A(n598), .B(n370), .ZN(n427) );
  NAND2_X1 U553 ( .A1(n394), .A2(n729), .ZN(n601) );
  NAND2_X1 U554 ( .A1(n395), .A2(n658), .ZN(n394) );
  NAND2_X1 U555 ( .A1(n732), .A2(n747), .ZN(n395) );
  NAND2_X1 U556 ( .A1(n396), .A2(G469), .ZN(n401) );
  NAND2_X1 U557 ( .A1(n396), .A2(G217), .ZN(n761) );
  NAND2_X1 U558 ( .A1(n396), .A2(G478), .ZN(n758) );
  NAND2_X1 U559 ( .A1(n476), .A2(n397), .ZN(n681) );
  NAND2_X1 U560 ( .A1(n692), .A2(n691), .ZN(n403) );
  NAND2_X1 U561 ( .A1(n692), .A2(n364), .ZN(n405) );
  XNOR2_X1 U562 ( .A(n467), .B(n371), .ZN(n466) );
  NAND2_X1 U563 ( .A1(n361), .A2(n410), .ZN(n678) );
  XNOR2_X1 U564 ( .A(n420), .B(n419), .ZN(G60) );
  NAND2_X1 U565 ( .A1(n643), .A2(KEYINPUT28), .ZN(n424) );
  NAND2_X1 U566 ( .A1(n638), .A2(n707), .ZN(n643) );
  XNOR2_X1 U567 ( .A(n425), .B(n508), .ZN(n448) );
  NAND2_X1 U568 ( .A1(n427), .A2(n639), .ZN(n611) );
  NAND2_X1 U569 ( .A1(n500), .A2(n499), .ZN(n498) );
  NAND2_X2 U570 ( .A1(n455), .A2(n453), .ZN(n659) );
  NAND2_X1 U571 ( .A1(n765), .A2(n435), .ZN(n676) );
  INV_X1 U572 ( .A(n436), .ZN(n435) );
  XNOR2_X1 U573 ( .A(n436), .B(n785), .ZN(n784) );
  NAND2_X1 U574 ( .A1(n604), .A2(n438), .ZN(n712) );
  INV_X1 U575 ( .A(n564), .ZN(n438) );
  NAND2_X1 U576 ( .A1(n439), .A2(n444), .ZN(n654) );
  INV_X1 U577 ( .A(n443), .ZN(n441) );
  INV_X1 U578 ( .A(n640), .ZN(n446) );
  NAND2_X1 U579 ( .A1(n665), .A2(n450), .ZN(n449) );
  NAND2_X1 U580 ( .A1(n452), .A2(n451), .ZN(n450) );
  INV_X1 U581 ( .A(KEYINPUT47), .ZN(n451) );
  NAND2_X1 U582 ( .A1(n358), .A2(KEYINPUT78), .ZN(n452) );
  INV_X1 U583 ( .A(n754), .ZN(n454) );
  NAND2_X1 U584 ( .A1(n754), .A2(n359), .ZN(n456) );
  NAND2_X1 U585 ( .A1(n679), .A2(n765), .ZN(n691) );
  INV_X1 U586 ( .A(n494), .ZN(n501) );
  XNOR2_X1 U587 ( .A(n463), .B(n491), .ZN(G75) );
  NAND2_X1 U588 ( .A1(n466), .A2(n662), .ZN(n465) );
  NAND2_X1 U589 ( .A1(n472), .A2(n475), .ZN(n471) );
  AND2_X1 U590 ( .A1(n666), .A2(n474), .ZN(n472) );
  XNOR2_X1 U591 ( .A(n642), .B(KEYINPUT46), .ZN(n475) );
  AND2_X1 U592 ( .A1(n691), .A2(n477), .ZN(n476) );
  INV_X1 U593 ( .A(n660), .ZN(n478) );
  NAND2_X1 U594 ( .A1(n368), .A2(n479), .ZN(n641) );
  NAND2_X1 U595 ( .A1(n480), .A2(n479), .ZN(n488) );
  INV_X1 U596 ( .A(n484), .ZN(n482) );
  NOR2_X1 U597 ( .A1(n633), .A2(n486), .ZN(n483) );
  NAND2_X1 U598 ( .A1(n633), .A2(n486), .ZN(n484) );
  INV_X1 U599 ( .A(KEYINPUT39), .ZN(n486) );
  INV_X1 U600 ( .A(KEYINPUT53), .ZN(n491) );
  NAND2_X1 U601 ( .A1(n497), .A2(n492), .ZN(n519) );
  NAND2_X1 U602 ( .A1(n494), .A2(n493), .ZN(n492) );
  NAND2_X1 U603 ( .A1(n511), .A2(n512), .ZN(n495) );
  NAND2_X1 U604 ( .A1(n513), .A2(KEYINPUT16), .ZN(n496) );
  NAND2_X1 U605 ( .A1(n501), .A2(n498), .ZN(n497) );
  NAND2_X1 U606 ( .A1(n511), .A2(KEYINPUT16), .ZN(n499) );
  NAND2_X1 U607 ( .A1(n513), .A2(n512), .ZN(n500) );
  XNOR2_X1 U608 ( .A(n501), .B(KEYINPUT16), .ZN(n772) );
  XNOR2_X1 U609 ( .A(n678), .B(KEYINPUT83), .ZN(n679) );
  XNOR2_X2 U610 ( .A(n526), .B(n525), .ZN(n754) );
  OR2_X1 U611 ( .A1(n748), .A2(n641), .ZN(n753) );
  NOR2_X1 U612 ( .A1(n797), .A2(n792), .ZN(n642) );
  XOR2_X1 U613 ( .A(n574), .B(n573), .Z(n502) );
  AND2_X1 U614 ( .A1(G210), .A2(n586), .ZN(n503) );
  NAND2_X1 U615 ( .A1(n751), .A2(n657), .ZN(n504) );
  INV_X1 U616 ( .A(KEYINPUT16), .ZN(n512) );
  INV_X1 U617 ( .A(KEYINPUT82), .ZN(n687) );
  INV_X1 U618 ( .A(KEYINPUT110), .ZN(n625) );
  INV_X1 U619 ( .A(KEYINPUT94), .ZN(n557) );
  INV_X1 U620 ( .A(n538), .ZN(n509) );
  INV_X1 U621 ( .A(n794), .ZN(n674) );
  XNOR2_X1 U622 ( .A(KEYINPUT100), .B(KEYINPUT7), .ZN(n568) );
  OR2_X1 U623 ( .A1(n603), .A2(n595), .ZN(n748) );
  NOR2_X1 U624 ( .A1(G952), .A2(n783), .ZN(n764) );
  XNOR2_X1 U625 ( .A(KEYINPUT62), .B(KEYINPUT113), .ZN(n510) );
  XOR2_X1 U626 ( .A(KEYINPUT95), .B(KEYINPUT5), .Z(n507) );
  XNOR2_X1 U627 ( .A(G146), .B(G137), .ZN(n506) );
  XNOR2_X1 U628 ( .A(n507), .B(n506), .ZN(n508) );
  NOR2_X1 U629 ( .A1(G953), .A2(G237), .ZN(n586) );
  XOR2_X2 U630 ( .A(G143), .B(G128), .Z(n511) );
  XNOR2_X1 U631 ( .A(n510), .B(n561), .ZN(n682) );
  INV_X1 U632 ( .A(n511), .ZN(n513) );
  NAND2_X1 U633 ( .A1(G224), .A2(n783), .ZN(n514) );
  XOR2_X1 U634 ( .A(n515), .B(n514), .Z(n517) );
  XOR2_X1 U635 ( .A(KEYINPUT73), .B(KEYINPUT18), .Z(n516) );
  XNOR2_X2 U636 ( .A(n519), .B(n518), .ZN(n526) );
  INV_X1 U637 ( .A(G146), .ZN(n521) );
  NAND2_X1 U638 ( .A1(n521), .A2(G125), .ZN(n524) );
  INV_X1 U639 ( .A(G125), .ZN(n522) );
  NAND2_X1 U640 ( .A1(n522), .A2(G146), .ZN(n523) );
  XNOR2_X1 U641 ( .A(n542), .B(n546), .ZN(n525) );
  XNOR2_X1 U642 ( .A(n527), .B(KEYINPUT88), .ZN(n680) );
  INV_X1 U643 ( .A(n680), .ZN(n528) );
  XNOR2_X1 U644 ( .A(n529), .B(KEYINPUT71), .ZN(n530) );
  NAND2_X1 U645 ( .A1(G214), .A2(n530), .ZN(n694) );
  XOR2_X1 U646 ( .A(KEYINPUT14), .B(n531), .Z(n622) );
  NAND2_X1 U647 ( .A1(n783), .A2(G952), .ZN(n621) );
  INV_X1 U648 ( .A(n621), .ZN(n533) );
  NAND2_X1 U649 ( .A1(G953), .A2(G902), .ZN(n618) );
  NOR2_X1 U650 ( .A1(G898), .A2(n618), .ZN(n532) );
  NOR2_X1 U651 ( .A1(n533), .A2(n532), .ZN(n534) );
  NOR2_X1 U652 ( .A1(n622), .A2(n534), .ZN(n535) );
  NAND2_X1 U653 ( .A1(G227), .A2(n783), .ZN(n539) );
  XNOR2_X1 U654 ( .A(n540), .B(n539), .ZN(n541) );
  XNOR2_X1 U655 ( .A(n542), .B(n541), .ZN(n543) );
  NOR2_X1 U656 ( .A1(n756), .A2(G902), .ZN(n545) );
  XNOR2_X1 U657 ( .A(KEYINPUT68), .B(G469), .ZN(n544) );
  XOR2_X1 U658 ( .A(KEYINPUT91), .B(G110), .Z(n548) );
  XNOR2_X1 U659 ( .A(G128), .B(G119), .ZN(n547) );
  XOR2_X1 U660 ( .A(KEYINPUT90), .B(KEYINPUT24), .Z(n549) );
  XOR2_X1 U661 ( .A(KEYINPUT80), .B(KEYINPUT8), .Z(n551) );
  NAND2_X1 U662 ( .A1(G234), .A2(n783), .ZN(n550) );
  XNOR2_X1 U663 ( .A(n551), .B(n550), .ZN(n572) );
  NAND2_X1 U664 ( .A1(G221), .A2(n572), .ZN(n553) );
  NAND2_X1 U665 ( .A1(n680), .A2(G234), .ZN(n555) );
  XNOR2_X1 U666 ( .A(KEYINPUT20), .B(KEYINPUT92), .ZN(n554) );
  XNOR2_X1 U667 ( .A(n555), .B(n554), .ZN(n559) );
  NAND2_X1 U668 ( .A1(G217), .A2(n559), .ZN(n556) );
  XNOR2_X1 U669 ( .A(KEYINPUT93), .B(KEYINPUT25), .ZN(n558) );
  NAND2_X1 U670 ( .A1(G221), .A2(n559), .ZN(n560) );
  XNOR2_X1 U671 ( .A(KEYINPUT21), .B(n560), .ZN(n596) );
  INV_X1 U672 ( .A(n596), .ZN(n707) );
  NAND2_X1 U673 ( .A1(n599), .A2(n707), .ZN(n703) );
  NOR2_X1 U674 ( .A1(n640), .A2(n703), .ZN(n626) );
  NOR2_X1 U675 ( .A1(n561), .A2(G902), .ZN(n563) );
  XOR2_X1 U676 ( .A(KEYINPUT103), .B(KEYINPUT104), .Z(n567) );
  XNOR2_X1 U677 ( .A(KEYINPUT101), .B(KEYINPUT9), .ZN(n566) );
  XNOR2_X1 U678 ( .A(n567), .B(n566), .ZN(n571) );
  XNOR2_X1 U679 ( .A(n569), .B(n568), .ZN(n570) );
  XOR2_X1 U680 ( .A(n571), .B(n570), .Z(n577) );
  NAND2_X1 U681 ( .A1(G217), .A2(n572), .ZN(n575) );
  NOR2_X1 U682 ( .A1(n759), .A2(G902), .ZN(n578) );
  XOR2_X1 U683 ( .A(KEYINPUT13), .B(KEYINPUT99), .Z(n580) );
  XNOR2_X1 U684 ( .A(KEYINPUT98), .B(G475), .ZN(n579) );
  XNOR2_X1 U685 ( .A(n580), .B(n579), .ZN(n594) );
  XNOR2_X1 U686 ( .A(n582), .B(n581), .ZN(n583) );
  XNOR2_X1 U687 ( .A(n779), .B(n583), .ZN(n592) );
  INV_X1 U688 ( .A(n584), .ZN(n585) );
  XNOR2_X1 U689 ( .A(n585), .B(KEYINPUT97), .ZN(n590) );
  XOR2_X1 U690 ( .A(KEYINPUT12), .B(KEYINPUT11), .Z(n588) );
  NAND2_X1 U691 ( .A1(n586), .A2(G214), .ZN(n587) );
  XNOR2_X1 U692 ( .A(n588), .B(n587), .ZN(n589) );
  XNOR2_X1 U693 ( .A(n590), .B(n589), .ZN(n591) );
  XNOR2_X1 U694 ( .A(n592), .B(n591), .ZN(n757) );
  NOR2_X1 U695 ( .A1(G902), .A2(n757), .ZN(n593) );
  XOR2_X1 U696 ( .A(n594), .B(n593), .Z(n602) );
  INV_X1 U697 ( .A(n602), .ZN(n595) );
  NAND2_X1 U698 ( .A1(n603), .A2(n595), .ZN(n744) );
  NAND2_X1 U699 ( .A1(n744), .A2(n748), .ZN(n658) );
  NAND2_X1 U700 ( .A1(n602), .A2(n603), .ZN(n696) );
  NOR2_X1 U701 ( .A1(n596), .A2(n696), .ZN(n597) );
  AND2_X1 U702 ( .A1(n706), .A2(n433), .ZN(n600) );
  XNOR2_X1 U703 ( .A(n601), .B(KEYINPUT105), .ZN(n608) );
  INV_X1 U704 ( .A(KEYINPUT44), .ZN(n606) );
  NOR2_X1 U705 ( .A1(n603), .A2(n602), .ZN(n662) );
  XOR2_X1 U706 ( .A(KEYINPUT33), .B(KEYINPUT69), .Z(n605) );
  NAND2_X1 U707 ( .A1(n607), .A2(n608), .ZN(n609) );
  NOR2_X1 U708 ( .A1(n433), .A2(n706), .ZN(n610) );
  NOR2_X1 U709 ( .A1(n706), .A2(n611), .ZN(n612) );
  NAND2_X1 U710 ( .A1(n612), .A2(n433), .ZN(n737) );
  NAND2_X1 U711 ( .A1(n793), .A2(n615), .ZN(n616) );
  XNOR2_X2 U712 ( .A(n617), .B(KEYINPUT45), .ZN(n765) );
  INV_X1 U713 ( .A(n622), .ZN(n721) );
  NOR2_X1 U714 ( .A1(G900), .A2(n618), .ZN(n619) );
  NAND2_X1 U715 ( .A1(n721), .A2(n619), .ZN(n620) );
  XNOR2_X1 U716 ( .A(n620), .B(KEYINPUT107), .ZN(n624) );
  NOR2_X1 U717 ( .A1(n622), .A2(n621), .ZN(n623) );
  NOR2_X1 U718 ( .A1(n624), .A2(n623), .ZN(n637) );
  XNOR2_X1 U719 ( .A(n626), .B(n625), .ZN(n627) );
  XNOR2_X1 U720 ( .A(n628), .B(KEYINPUT72), .ZN(n631) );
  NAND2_X1 U721 ( .A1(n694), .A2(n636), .ZN(n629) );
  XOR2_X1 U722 ( .A(KEYINPUT30), .B(n629), .Z(n630) );
  NAND2_X1 U723 ( .A1(n631), .A2(n630), .ZN(n660) );
  XOR2_X1 U724 ( .A(KEYINPUT38), .B(KEYINPUT70), .Z(n632) );
  XOR2_X1 U725 ( .A(n659), .B(n632), .Z(n633) );
  INV_X1 U726 ( .A(n633), .ZN(n693) );
  NAND2_X1 U727 ( .A1(n694), .A2(n693), .ZN(n697) );
  NOR2_X1 U728 ( .A1(n696), .A2(n697), .ZN(n635) );
  XNOR2_X1 U729 ( .A(KEYINPUT111), .B(KEYINPUT41), .ZN(n634) );
  INV_X1 U730 ( .A(n636), .ZN(n639) );
  NOR2_X1 U731 ( .A1(n706), .A2(n637), .ZN(n638) );
  NOR2_X1 U732 ( .A1(n744), .A2(n643), .ZN(n644) );
  NAND2_X1 U733 ( .A1(n645), .A2(n644), .ZN(n646) );
  XNOR2_X1 U734 ( .A(KEYINPUT108), .B(n646), .ZN(n667) );
  XNOR2_X1 U735 ( .A(KEYINPUT112), .B(n667), .ZN(n647) );
  NOR2_X1 U736 ( .A1(n648), .A2(n647), .ZN(n649) );
  XNOR2_X1 U737 ( .A(n649), .B(KEYINPUT36), .ZN(n650) );
  INV_X1 U738 ( .A(n433), .ZN(n668) );
  NAND2_X1 U739 ( .A1(n650), .A2(n668), .ZN(n751) );
  BUF_X1 U740 ( .A(n651), .Z(n652) );
  NAND2_X1 U741 ( .A1(n742), .A2(KEYINPUT78), .ZN(n655) );
  NAND2_X1 U742 ( .A1(n655), .A2(n658), .ZN(n656) );
  NAND2_X1 U743 ( .A1(n656), .A2(KEYINPUT47), .ZN(n657) );
  INV_X1 U744 ( .A(n658), .ZN(n698) );
  INV_X1 U745 ( .A(n659), .ZN(n671) );
  NOR2_X1 U746 ( .A1(n671), .A2(n660), .ZN(n661) );
  NAND2_X1 U747 ( .A1(n662), .A2(n661), .ZN(n741) );
  XNOR2_X1 U748 ( .A(n741), .B(KEYINPUT79), .ZN(n664) );
  NOR2_X1 U749 ( .A1(n742), .A2(KEYINPUT78), .ZN(n663) );
  NOR2_X1 U750 ( .A1(n664), .A2(n663), .ZN(n665) );
  NOR2_X1 U751 ( .A1(n668), .A2(n667), .ZN(n669) );
  NAND2_X1 U752 ( .A1(n669), .A2(n694), .ZN(n670) );
  XNOR2_X1 U753 ( .A(n670), .B(KEYINPUT43), .ZN(n672) );
  NAND2_X1 U754 ( .A1(n672), .A2(n671), .ZN(n673) );
  XNOR2_X1 U755 ( .A(KEYINPUT109), .B(n673), .ZN(n794) );
  INV_X1 U756 ( .A(KEYINPUT2), .ZN(n675) );
  NAND2_X1 U757 ( .A1(KEYINPUT2), .A2(n753), .ZN(n677) );
  XOR2_X1 U758 ( .A(n682), .B(n681), .Z(n683) );
  XOR2_X1 U759 ( .A(KEYINPUT86), .B(KEYINPUT63), .Z(n684) );
  XNOR2_X1 U760 ( .A(n685), .B(n684), .ZN(G57) );
  XNOR2_X1 U761 ( .A(n686), .B(KEYINPUT81), .ZN(n689) );
  XNOR2_X1 U762 ( .A(n363), .B(n687), .ZN(n688) );
  NAND2_X1 U763 ( .A1(n689), .A2(n688), .ZN(n690) );
  XNOR2_X1 U764 ( .A(n690), .B(KEYINPUT77), .ZN(n692) );
  INV_X1 U765 ( .A(n725), .ZN(n702) );
  NOR2_X1 U766 ( .A1(n694), .A2(n693), .ZN(n695) );
  NOR2_X1 U767 ( .A1(n696), .A2(n695), .ZN(n700) );
  NOR2_X1 U768 ( .A1(n698), .A2(n697), .ZN(n699) );
  NOR2_X1 U769 ( .A1(n700), .A2(n699), .ZN(n701) );
  NOR2_X1 U770 ( .A1(n702), .A2(n701), .ZN(n719) );
  XNOR2_X1 U771 ( .A(KEYINPUT120), .B(KEYINPUT51), .ZN(n715) );
  NAND2_X1 U772 ( .A1(n433), .A2(n703), .ZN(n705) );
  XNOR2_X1 U773 ( .A(n705), .B(KEYINPUT50), .ZN(n711) );
  NOR2_X1 U774 ( .A1(n707), .A2(n706), .ZN(n708) );
  XOR2_X1 U775 ( .A(KEYINPUT49), .B(n708), .Z(n709) );
  NAND2_X1 U776 ( .A1(n711), .A2(n710), .ZN(n713) );
  NAND2_X1 U777 ( .A1(n713), .A2(n712), .ZN(n714) );
  XNOR2_X1 U778 ( .A(n715), .B(n714), .ZN(n717) );
  INV_X1 U779 ( .A(n724), .ZN(n716) );
  NOR2_X1 U780 ( .A1(n717), .A2(n716), .ZN(n718) );
  NOR2_X1 U781 ( .A1(n719), .A2(n718), .ZN(n720) );
  XNOR2_X1 U782 ( .A(KEYINPUT52), .B(n720), .ZN(n723) );
  NAND2_X1 U783 ( .A1(G952), .A2(n721), .ZN(n722) );
  OR2_X1 U784 ( .A1(n723), .A2(n722), .ZN(n727) );
  NAND2_X1 U785 ( .A1(n725), .A2(n724), .ZN(n726) );
  AND2_X1 U786 ( .A1(n727), .A2(n726), .ZN(n728) );
  XNOR2_X1 U787 ( .A(G101), .B(KEYINPUT114), .ZN(n730) );
  XNOR2_X1 U788 ( .A(n730), .B(n729), .ZN(G3) );
  NOR2_X1 U789 ( .A1(n732), .A2(n744), .ZN(n731) );
  XOR2_X1 U790 ( .A(G104), .B(n731), .Z(G6) );
  NOR2_X1 U791 ( .A1(n732), .A2(n748), .ZN(n734) );
  XNOR2_X1 U792 ( .A(KEYINPUT27), .B(KEYINPUT26), .ZN(n733) );
  XNOR2_X1 U793 ( .A(n734), .B(n733), .ZN(n735) );
  XNOR2_X1 U794 ( .A(G107), .B(n735), .ZN(G9) );
  XOR2_X1 U795 ( .A(G110), .B(KEYINPUT115), .Z(n736) );
  XNOR2_X1 U796 ( .A(n737), .B(n736), .ZN(G12) );
  NOR2_X1 U797 ( .A1(n748), .A2(n742), .ZN(n739) );
  XNOR2_X1 U798 ( .A(KEYINPUT116), .B(KEYINPUT29), .ZN(n738) );
  XNOR2_X1 U799 ( .A(n739), .B(n738), .ZN(n740) );
  XNOR2_X1 U800 ( .A(G128), .B(n740), .ZN(G30) );
  XNOR2_X1 U801 ( .A(G143), .B(n741), .ZN(G45) );
  NOR2_X1 U802 ( .A1(n744), .A2(n742), .ZN(n743) );
  XOR2_X1 U803 ( .A(G146), .B(n743), .Z(G48) );
  NOR2_X1 U804 ( .A1(n744), .A2(n747), .ZN(n746) );
  XNOR2_X1 U805 ( .A(G113), .B(KEYINPUT117), .ZN(n745) );
  XNOR2_X1 U806 ( .A(n746), .B(n745), .ZN(G15) );
  NOR2_X1 U807 ( .A1(n748), .A2(n747), .ZN(n749) );
  XOR2_X1 U808 ( .A(n356), .B(n749), .Z(G18) );
  XOR2_X1 U809 ( .A(KEYINPUT37), .B(KEYINPUT118), .Z(n750) );
  XNOR2_X1 U810 ( .A(n751), .B(n750), .ZN(n752) );
  XNOR2_X1 U811 ( .A(G125), .B(n752), .ZN(G27) );
  XNOR2_X1 U812 ( .A(G134), .B(n753), .ZN(G36) );
  XOR2_X1 U813 ( .A(KEYINPUT54), .B(KEYINPUT55), .Z(n755) );
  XNOR2_X1 U814 ( .A(n759), .B(n758), .ZN(n760) );
  NOR2_X1 U815 ( .A1(n764), .A2(n760), .ZN(G63) );
  XNOR2_X1 U816 ( .A(n762), .B(n761), .ZN(n763) );
  NOR2_X1 U817 ( .A1(n764), .A2(n763), .ZN(G66) );
  NAND2_X1 U818 ( .A1(n765), .A2(n783), .ZN(n771) );
  NAND2_X1 U819 ( .A1(G224), .A2(G953), .ZN(n766) );
  XNOR2_X1 U820 ( .A(n766), .B(KEYINPUT61), .ZN(n767) );
  XNOR2_X1 U821 ( .A(KEYINPUT122), .B(n767), .ZN(n768) );
  NAND2_X1 U822 ( .A1(n768), .A2(G898), .ZN(n769) );
  XOR2_X1 U823 ( .A(KEYINPUT123), .B(n769), .Z(n770) );
  NAND2_X1 U824 ( .A1(n771), .A2(n770), .ZN(n778) );
  XOR2_X1 U825 ( .A(n772), .B(n773), .Z(n774) );
  XNOR2_X1 U826 ( .A(G101), .B(n774), .ZN(n776) );
  NOR2_X1 U827 ( .A1(G898), .A2(n783), .ZN(n775) );
  NOR2_X1 U828 ( .A1(n776), .A2(n775), .ZN(n777) );
  XNOR2_X1 U829 ( .A(n778), .B(n777), .ZN(G69) );
  XOR2_X1 U830 ( .A(KEYINPUT4), .B(KEYINPUT124), .Z(n780) );
  XNOR2_X1 U831 ( .A(n781), .B(n780), .ZN(n782) );
  XOR2_X1 U832 ( .A(n779), .B(n782), .Z(n785) );
  NAND2_X1 U833 ( .A1(n784), .A2(n783), .ZN(n790) );
  XNOR2_X1 U834 ( .A(G227), .B(n785), .ZN(n786) );
  NAND2_X1 U835 ( .A1(n786), .A2(G900), .ZN(n787) );
  XOR2_X1 U836 ( .A(KEYINPUT125), .B(n787), .Z(n788) );
  NAND2_X1 U837 ( .A1(G953), .A2(n788), .ZN(n789) );
  NAND2_X1 U838 ( .A1(n790), .A2(n789), .ZN(G72) );
  XOR2_X1 U839 ( .A(G131), .B(KEYINPUT126), .Z(n791) );
  XNOR2_X1 U840 ( .A(n792), .B(n791), .ZN(G33) );
  XNOR2_X1 U841 ( .A(n793), .B(G122), .ZN(G24) );
  XNOR2_X1 U842 ( .A(G140), .B(n794), .ZN(n795) );
  XNOR2_X1 U843 ( .A(n795), .B(KEYINPUT119), .ZN(G42) );
  XNOR2_X1 U844 ( .A(n796), .B(G119), .ZN(G21) );
  XOR2_X1 U845 ( .A(n797), .B(G137), .Z(G39) );
endmodule

