//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 1 0 1 1 0 0 0 0 0 1 1 0 1 0 0 0 0 0 1 0 1 0 1 1 1 1 0 0 0 1 0 0 0 1 0 1 1 0 1 1 0 0 0 0 1 0 1 1 1 0 1 1 0 0 1 0 0 1 0 0 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:31:39 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n445, new_n447, new_n451, new_n452, new_n453, new_n454, new_n457,
    new_n458, new_n459, new_n460, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n522, new_n523, new_n524, new_n525,
    new_n526, new_n527, new_n528, new_n529, new_n530, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n539, new_n540, new_n541, new_n542,
    new_n543, new_n544, new_n545, new_n546, new_n549, new_n550, new_n551,
    new_n553, new_n554, new_n555, new_n556, new_n557, new_n558, new_n559,
    new_n560, new_n561, new_n562, new_n566, new_n567, new_n568, new_n570,
    new_n571, new_n572, new_n573, new_n574, new_n575, new_n576, new_n577,
    new_n578, new_n579, new_n580, new_n581, new_n583, new_n584, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n600, new_n601, new_n602,
    new_n605, new_n607, new_n608, new_n609, new_n610, new_n612, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1191, new_n1192, new_n1193, new_n1194, new_n1195, new_n1196;
  XNOR2_X1  g000(.A(KEYINPUT64), .B(G452), .ZN(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  XOR2_X1   g007(.A(KEYINPUT65), .B(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  XOR2_X1   g011(.A(KEYINPUT66), .B(G96), .Z(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  XNOR2_X1  g014(.A(KEYINPUT67), .B(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  NAND2_X1  g019(.A1(G94), .A2(G452), .ZN(new_n445));
  XOR2_X1   g020(.A(new_n445), .B(KEYINPUT68), .Z(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g025(.A1(G221), .A2(G220), .A3(G218), .A4(G219), .ZN(new_n451));
  XOR2_X1   g026(.A(new_n451), .B(KEYINPUT2), .Z(new_n452));
  NOR4_X1   g027(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n453));
  INV_X1    g028(.A(new_n453), .ZN(new_n454));
  NOR2_X1   g029(.A1(new_n452), .A2(new_n454), .ZN(G325));
  INV_X1    g030(.A(G325), .ZN(G261));
  NAND2_X1  g031(.A1(new_n452), .A2(G2106), .ZN(new_n457));
  NAND2_X1  g032(.A1(new_n454), .A2(G567), .ZN(new_n458));
  XNOR2_X1  g033(.A(new_n458), .B(KEYINPUT69), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n457), .A2(new_n459), .ZN(new_n460));
  INV_X1    g035(.A(new_n460), .ZN(G319));
  INV_X1    g036(.A(G2105), .ZN(new_n462));
  AND2_X1   g037(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n463));
  NOR2_X1   g038(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n464));
  OAI21_X1  g039(.A(G125), .B1(new_n463), .B2(new_n464), .ZN(new_n465));
  NAND2_X1  g040(.A1(G113), .A2(G2104), .ZN(new_n466));
  AOI21_X1  g041(.A(new_n462), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  OAI211_X1 g042(.A(G137), .B(new_n462), .C1(new_n463), .C2(new_n464), .ZN(new_n468));
  AND2_X1   g043(.A1(new_n462), .A2(G2104), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n469), .A2(G101), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n468), .A2(new_n470), .ZN(new_n471));
  NOR2_X1   g046(.A1(new_n467), .A2(new_n471), .ZN(G160));
  OAI21_X1  g047(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n473));
  INV_X1    g048(.A(G112), .ZN(new_n474));
  AOI21_X1  g049(.A(new_n473), .B1(new_n474), .B2(G2105), .ZN(new_n475));
  OR2_X1    g050(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n476));
  NAND2_X1  g051(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n477));
  AOI21_X1  g052(.A(G2105), .B1(new_n476), .B2(new_n477), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n478), .A2(G136), .ZN(new_n479));
  INV_X1    g054(.A(new_n479), .ZN(new_n480));
  AOI21_X1  g055(.A(new_n462), .B1(new_n476), .B2(new_n477), .ZN(new_n481));
  AOI211_X1 g056(.A(new_n475), .B(new_n480), .C1(G124), .C2(new_n481), .ZN(G162));
  OAI21_X1  g057(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n483));
  INV_X1    g058(.A(new_n483), .ZN(new_n484));
  INV_X1    g059(.A(KEYINPUT70), .ZN(new_n485));
  INV_X1    g060(.A(G114), .ZN(new_n486));
  NAND3_X1  g061(.A1(new_n485), .A2(new_n486), .A3(G2105), .ZN(new_n487));
  OAI21_X1  g062(.A(KEYINPUT70), .B1(new_n462), .B2(G114), .ZN(new_n488));
  NAND3_X1  g063(.A1(new_n484), .A2(new_n487), .A3(new_n488), .ZN(new_n489));
  OAI211_X1 g064(.A(G126), .B(G2105), .C1(new_n463), .C2(new_n464), .ZN(new_n490));
  NAND2_X1  g065(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  INV_X1    g066(.A(G138), .ZN(new_n492));
  NOR2_X1   g067(.A1(new_n492), .A2(G2105), .ZN(new_n493));
  OAI21_X1  g068(.A(new_n493), .B1(new_n463), .B2(new_n464), .ZN(new_n494));
  NAND2_X1  g069(.A1(new_n494), .A2(KEYINPUT4), .ZN(new_n495));
  INV_X1    g070(.A(KEYINPUT4), .ZN(new_n496));
  OAI211_X1 g071(.A(new_n493), .B(new_n496), .C1(new_n464), .C2(new_n463), .ZN(new_n497));
  AOI21_X1  g072(.A(new_n491), .B1(new_n495), .B2(new_n497), .ZN(G164));
  XNOR2_X1  g073(.A(KEYINPUT6), .B(G651), .ZN(new_n499));
  AND2_X1   g074(.A1(new_n499), .A2(G543), .ZN(new_n500));
  NAND2_X1  g075(.A1(new_n500), .A2(G50), .ZN(new_n501));
  INV_X1    g076(.A(KEYINPUT71), .ZN(new_n502));
  INV_X1    g077(.A(KEYINPUT5), .ZN(new_n503));
  OAI21_X1  g078(.A(new_n502), .B1(new_n503), .B2(G543), .ZN(new_n504));
  INV_X1    g079(.A(G543), .ZN(new_n505));
  NAND3_X1  g080(.A1(new_n505), .A2(KEYINPUT71), .A3(KEYINPUT5), .ZN(new_n506));
  NAND2_X1  g081(.A1(new_n504), .A2(new_n506), .ZN(new_n507));
  INV_X1    g082(.A(KEYINPUT72), .ZN(new_n508));
  OAI21_X1  g083(.A(new_n508), .B1(new_n505), .B2(KEYINPUT5), .ZN(new_n509));
  NAND3_X1  g084(.A1(new_n503), .A2(KEYINPUT72), .A3(G543), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  AND3_X1   g086(.A1(new_n507), .A2(new_n511), .A3(new_n499), .ZN(new_n512));
  INV_X1    g087(.A(new_n512), .ZN(new_n513));
  INV_X1    g088(.A(G88), .ZN(new_n514));
  OAI21_X1  g089(.A(new_n501), .B1(new_n513), .B2(new_n514), .ZN(new_n515));
  INV_X1    g090(.A(G651), .ZN(new_n516));
  AND2_X1   g091(.A1(new_n507), .A2(new_n511), .ZN(new_n517));
  NAND2_X1  g092(.A1(new_n517), .A2(G62), .ZN(new_n518));
  NAND2_X1  g093(.A1(G75), .A2(G543), .ZN(new_n519));
  AOI21_X1  g094(.A(new_n516), .B1(new_n518), .B2(new_n519), .ZN(new_n520));
  NOR2_X1   g095(.A1(new_n515), .A2(new_n520), .ZN(G166));
  NAND3_X1  g096(.A1(new_n517), .A2(G63), .A3(G651), .ZN(new_n522));
  XOR2_X1   g097(.A(KEYINPUT73), .B(G51), .Z(new_n523));
  NAND3_X1  g098(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n524));
  NAND2_X1  g099(.A1(new_n524), .A2(KEYINPUT7), .ZN(new_n525));
  OR2_X1    g100(.A1(new_n524), .A2(KEYINPUT7), .ZN(new_n526));
  AOI22_X1  g101(.A1(new_n500), .A2(new_n523), .B1(new_n525), .B2(new_n526), .ZN(new_n527));
  AND2_X1   g102(.A1(new_n522), .A2(new_n527), .ZN(new_n528));
  XOR2_X1   g103(.A(KEYINPUT74), .B(G89), .Z(new_n529));
  NAND2_X1  g104(.A1(new_n512), .A2(new_n529), .ZN(new_n530));
  NAND2_X1  g105(.A1(new_n528), .A2(new_n530), .ZN(G286));
  INV_X1    g106(.A(G286), .ZN(G168));
  AOI22_X1  g107(.A1(new_n517), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n533));
  NOR2_X1   g108(.A1(new_n533), .A2(new_n516), .ZN(new_n534));
  NAND2_X1  g109(.A1(new_n500), .A2(G52), .ZN(new_n535));
  INV_X1    g110(.A(G90), .ZN(new_n536));
  OAI21_X1  g111(.A(new_n535), .B1(new_n513), .B2(new_n536), .ZN(new_n537));
  NOR2_X1   g112(.A1(new_n534), .A2(new_n537), .ZN(G171));
  NAND2_X1  g113(.A1(G68), .A2(G543), .ZN(new_n539));
  NAND2_X1  g114(.A1(new_n507), .A2(new_n511), .ZN(new_n540));
  INV_X1    g115(.A(G56), .ZN(new_n541));
  OAI21_X1  g116(.A(new_n539), .B1(new_n540), .B2(new_n541), .ZN(new_n542));
  NAND2_X1  g117(.A1(new_n542), .A2(G651), .ZN(new_n543));
  AOI22_X1  g118(.A1(new_n512), .A2(G81), .B1(G43), .B2(new_n500), .ZN(new_n544));
  NAND2_X1  g119(.A1(new_n543), .A2(new_n544), .ZN(new_n545));
  INV_X1    g120(.A(new_n545), .ZN(new_n546));
  NAND2_X1  g121(.A1(new_n546), .A2(G860), .ZN(G153));
  NAND4_X1  g122(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g123(.A1(G1), .A2(G3), .ZN(new_n549));
  XNOR2_X1  g124(.A(new_n549), .B(KEYINPUT75), .ZN(new_n550));
  XNOR2_X1  g125(.A(new_n550), .B(KEYINPUT8), .ZN(new_n551));
  NAND4_X1  g126(.A1(G319), .A2(G483), .A3(G661), .A4(new_n551), .ZN(G188));
  NAND3_X1  g127(.A1(new_n499), .A2(G53), .A3(G543), .ZN(new_n553));
  XNOR2_X1  g128(.A(KEYINPUT76), .B(KEYINPUT9), .ZN(new_n554));
  OR3_X1    g129(.A1(new_n553), .A2(KEYINPUT77), .A3(new_n554), .ZN(new_n555));
  OAI21_X1  g130(.A(KEYINPUT77), .B1(new_n553), .B2(new_n554), .ZN(new_n556));
  NAND2_X1  g131(.A1(new_n553), .A2(KEYINPUT9), .ZN(new_n557));
  NAND3_X1  g132(.A1(new_n555), .A2(new_n556), .A3(new_n557), .ZN(new_n558));
  NAND2_X1  g133(.A1(G78), .A2(G543), .ZN(new_n559));
  XOR2_X1   g134(.A(KEYINPUT78), .B(G65), .Z(new_n560));
  OAI21_X1  g135(.A(new_n559), .B1(new_n540), .B2(new_n560), .ZN(new_n561));
  AOI22_X1  g136(.A1(new_n561), .A2(G651), .B1(new_n512), .B2(G91), .ZN(new_n562));
  NAND2_X1  g137(.A1(new_n558), .A2(new_n562), .ZN(G299));
  INV_X1    g138(.A(G171), .ZN(G301));
  INV_X1    g139(.A(G166), .ZN(G303));
  OAI21_X1  g140(.A(G651), .B1(new_n517), .B2(G74), .ZN(new_n566));
  NAND2_X1  g141(.A1(new_n512), .A2(G87), .ZN(new_n567));
  NAND2_X1  g142(.A1(new_n500), .A2(G49), .ZN(new_n568));
  NAND3_X1  g143(.A1(new_n566), .A2(new_n567), .A3(new_n568), .ZN(G288));
  NAND2_X1  g144(.A1(G73), .A2(G543), .ZN(new_n570));
  INV_X1    g145(.A(G61), .ZN(new_n571));
  OAI21_X1  g146(.A(new_n570), .B1(new_n540), .B2(new_n571), .ZN(new_n572));
  INV_X1    g147(.A(KEYINPUT79), .ZN(new_n573));
  AND3_X1   g148(.A1(new_n572), .A2(new_n573), .A3(G651), .ZN(new_n574));
  AOI21_X1  g149(.A(new_n573), .B1(new_n572), .B2(G651), .ZN(new_n575));
  NOR2_X1   g150(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  NAND3_X1  g151(.A1(new_n512), .A2(KEYINPUT80), .A3(G86), .ZN(new_n577));
  NAND4_X1  g152(.A1(new_n507), .A2(new_n511), .A3(G86), .A4(new_n499), .ZN(new_n578));
  INV_X1    g153(.A(KEYINPUT80), .ZN(new_n579));
  NAND2_X1  g154(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  AOI22_X1  g155(.A1(new_n577), .A2(new_n580), .B1(G48), .B2(new_n500), .ZN(new_n581));
  NAND2_X1  g156(.A1(new_n576), .A2(new_n581), .ZN(G305));
  AOI22_X1  g157(.A1(new_n512), .A2(G85), .B1(G47), .B2(new_n500), .ZN(new_n583));
  AOI22_X1  g158(.A1(new_n517), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n584));
  OAI21_X1  g159(.A(new_n583), .B1(new_n584), .B2(new_n516), .ZN(G290));
  NAND2_X1  g160(.A1(G301), .A2(G868), .ZN(new_n586));
  NAND2_X1  g161(.A1(new_n512), .A2(G92), .ZN(new_n587));
  XOR2_X1   g162(.A(new_n587), .B(KEYINPUT81), .Z(new_n588));
  NAND2_X1  g163(.A1(new_n588), .A2(KEYINPUT10), .ZN(new_n589));
  XNOR2_X1  g164(.A(new_n587), .B(KEYINPUT81), .ZN(new_n590));
  INV_X1    g165(.A(KEYINPUT10), .ZN(new_n591));
  NAND2_X1  g166(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  NAND2_X1  g167(.A1(G79), .A2(G543), .ZN(new_n593));
  INV_X1    g168(.A(G66), .ZN(new_n594));
  OAI21_X1  g169(.A(new_n593), .B1(new_n540), .B2(new_n594), .ZN(new_n595));
  AOI22_X1  g170(.A1(new_n595), .A2(G651), .B1(G54), .B2(new_n500), .ZN(new_n596));
  AND3_X1   g171(.A1(new_n589), .A2(new_n592), .A3(new_n596), .ZN(new_n597));
  OAI21_X1  g172(.A(new_n586), .B1(new_n597), .B2(G868), .ZN(G284));
  OAI21_X1  g173(.A(new_n586), .B1(new_n597), .B2(G868), .ZN(G321));
  INV_X1    g174(.A(G868), .ZN(new_n600));
  NAND2_X1  g175(.A1(G299), .A2(new_n600), .ZN(new_n601));
  OAI21_X1  g176(.A(new_n601), .B1(G168), .B2(new_n600), .ZN(new_n602));
  XOR2_X1   g177(.A(new_n602), .B(KEYINPUT82), .Z(G297));
  XOR2_X1   g178(.A(new_n602), .B(KEYINPUT83), .Z(G280));
  INV_X1    g179(.A(G559), .ZN(new_n605));
  OAI21_X1  g180(.A(new_n597), .B1(new_n605), .B2(G860), .ZN(G148));
  NAND3_X1  g181(.A1(new_n589), .A2(new_n592), .A3(new_n596), .ZN(new_n607));
  OR3_X1    g182(.A1(new_n607), .A2(KEYINPUT84), .A3(G559), .ZN(new_n608));
  OAI21_X1  g183(.A(KEYINPUT84), .B1(new_n607), .B2(G559), .ZN(new_n609));
  NAND2_X1  g184(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  MUX2_X1   g185(.A(new_n545), .B(new_n610), .S(G868), .Z(G323));
  XOR2_X1   g186(.A(KEYINPUT85), .B(KEYINPUT11), .Z(new_n612));
  XNOR2_X1  g187(.A(G323), .B(new_n612), .ZN(G282));
  XNOR2_X1  g188(.A(KEYINPUT3), .B(G2104), .ZN(new_n614));
  NAND2_X1  g189(.A1(new_n614), .A2(new_n469), .ZN(new_n615));
  XOR2_X1   g190(.A(new_n615), .B(KEYINPUT12), .Z(new_n616));
  XOR2_X1   g191(.A(new_n616), .B(KEYINPUT13), .Z(new_n617));
  INV_X1    g192(.A(new_n617), .ZN(new_n618));
  OR2_X1    g193(.A1(new_n618), .A2(G2100), .ZN(new_n619));
  NAND2_X1  g194(.A1(new_n478), .A2(G135), .ZN(new_n620));
  XNOR2_X1  g195(.A(new_n620), .B(KEYINPUT86), .ZN(new_n621));
  OAI21_X1  g196(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n622));
  INV_X1    g197(.A(G111), .ZN(new_n623));
  AOI21_X1  g198(.A(new_n622), .B1(new_n623), .B2(G2105), .ZN(new_n624));
  AOI21_X1  g199(.A(new_n624), .B1(new_n481), .B2(G123), .ZN(new_n625));
  AND2_X1   g200(.A1(new_n621), .A2(new_n625), .ZN(new_n626));
  INV_X1    g201(.A(new_n626), .ZN(new_n627));
  OR2_X1    g202(.A1(new_n627), .A2(G2096), .ZN(new_n628));
  NAND2_X1  g203(.A1(new_n618), .A2(G2100), .ZN(new_n629));
  NAND2_X1  g204(.A1(new_n627), .A2(G2096), .ZN(new_n630));
  NAND4_X1  g205(.A1(new_n619), .A2(new_n628), .A3(new_n629), .A4(new_n630), .ZN(G156));
  XNOR2_X1  g206(.A(G2427), .B(G2438), .ZN(new_n632));
  XNOR2_X1  g207(.A(new_n632), .B(G2430), .ZN(new_n633));
  XNOR2_X1  g208(.A(KEYINPUT15), .B(G2435), .ZN(new_n634));
  OR2_X1    g209(.A1(new_n633), .A2(new_n634), .ZN(new_n635));
  NAND2_X1  g210(.A1(new_n633), .A2(new_n634), .ZN(new_n636));
  NAND3_X1  g211(.A1(new_n635), .A2(KEYINPUT14), .A3(new_n636), .ZN(new_n637));
  XNOR2_X1  g212(.A(G2451), .B(G2454), .ZN(new_n638));
  XNOR2_X1  g213(.A(new_n638), .B(KEYINPUT16), .ZN(new_n639));
  XNOR2_X1  g214(.A(new_n637), .B(new_n639), .ZN(new_n640));
  XNOR2_X1  g215(.A(G2443), .B(G2446), .ZN(new_n641));
  XNOR2_X1  g216(.A(new_n640), .B(new_n641), .ZN(new_n642));
  XNOR2_X1  g217(.A(G1341), .B(G1348), .ZN(new_n643));
  NOR2_X1   g218(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  XNOR2_X1  g219(.A(new_n644), .B(KEYINPUT87), .ZN(new_n645));
  INV_X1    g220(.A(G14), .ZN(new_n646));
  AOI21_X1  g221(.A(new_n646), .B1(new_n642), .B2(new_n643), .ZN(new_n647));
  AND2_X1   g222(.A1(new_n645), .A2(new_n647), .ZN(G401));
  XNOR2_X1  g223(.A(G2072), .B(G2078), .ZN(new_n649));
  XNOR2_X1  g224(.A(new_n649), .B(KEYINPUT88), .ZN(new_n650));
  XNOR2_X1  g225(.A(new_n650), .B(KEYINPUT17), .ZN(new_n651));
  XNOR2_X1  g226(.A(G2067), .B(G2678), .ZN(new_n652));
  XNOR2_X1  g227(.A(G2084), .B(G2090), .ZN(new_n653));
  NOR3_X1   g228(.A1(new_n651), .A2(new_n652), .A3(new_n653), .ZN(new_n654));
  OAI21_X1  g229(.A(new_n653), .B1(new_n650), .B2(new_n652), .ZN(new_n655));
  AOI21_X1  g230(.A(new_n655), .B1(new_n651), .B2(new_n652), .ZN(new_n656));
  INV_X1    g231(.A(new_n652), .ZN(new_n657));
  NOR2_X1   g232(.A1(new_n657), .A2(new_n653), .ZN(new_n658));
  NAND2_X1  g233(.A1(new_n650), .A2(new_n658), .ZN(new_n659));
  XNOR2_X1  g234(.A(new_n659), .B(KEYINPUT18), .ZN(new_n660));
  OR3_X1    g235(.A1(new_n654), .A2(new_n656), .A3(new_n660), .ZN(new_n661));
  XNOR2_X1  g236(.A(G2096), .B(G2100), .ZN(new_n662));
  INV_X1    g237(.A(new_n662), .ZN(new_n663));
  OR2_X1    g238(.A1(new_n661), .A2(new_n663), .ZN(new_n664));
  NAND2_X1  g239(.A1(new_n661), .A2(new_n663), .ZN(new_n665));
  NAND2_X1  g240(.A1(new_n664), .A2(new_n665), .ZN(G227));
  XNOR2_X1  g241(.A(G1971), .B(G1976), .ZN(new_n667));
  XNOR2_X1  g242(.A(new_n667), .B(KEYINPUT19), .ZN(new_n668));
  INV_X1    g243(.A(new_n668), .ZN(new_n669));
  XOR2_X1   g244(.A(G1961), .B(G1966), .Z(new_n670));
  XNOR2_X1  g245(.A(new_n670), .B(KEYINPUT89), .ZN(new_n671));
  XNOR2_X1  g246(.A(G1956), .B(G2474), .ZN(new_n672));
  INV_X1    g247(.A(new_n672), .ZN(new_n673));
  NAND3_X1  g248(.A1(new_n669), .A2(new_n671), .A3(new_n673), .ZN(new_n674));
  XNOR2_X1  g249(.A(new_n674), .B(KEYINPUT20), .ZN(new_n675));
  AOI21_X1  g250(.A(new_n669), .B1(new_n671), .B2(new_n673), .ZN(new_n676));
  OR2_X1    g251(.A1(new_n671), .A2(new_n673), .ZN(new_n677));
  NAND2_X1  g252(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  OAI211_X1 g253(.A(new_n675), .B(new_n678), .C1(new_n668), .C2(new_n677), .ZN(new_n679));
  INV_X1    g254(.A(G1981), .ZN(new_n680));
  XNOR2_X1  g255(.A(new_n679), .B(new_n680), .ZN(new_n681));
  OR2_X1    g256(.A1(new_n681), .A2(G1986), .ZN(new_n682));
  XNOR2_X1  g257(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n683));
  XNOR2_X1  g258(.A(new_n683), .B(KEYINPUT90), .ZN(new_n684));
  INV_X1    g259(.A(new_n684), .ZN(new_n685));
  NAND2_X1  g260(.A1(new_n681), .A2(G1986), .ZN(new_n686));
  NAND3_X1  g261(.A1(new_n682), .A2(new_n685), .A3(new_n686), .ZN(new_n687));
  INV_X1    g262(.A(new_n687), .ZN(new_n688));
  XNOR2_X1  g263(.A(G1991), .B(G1996), .ZN(new_n689));
  INV_X1    g264(.A(new_n689), .ZN(new_n690));
  AOI21_X1  g265(.A(new_n685), .B1(new_n682), .B2(new_n686), .ZN(new_n691));
  OR3_X1    g266(.A1(new_n688), .A2(new_n690), .A3(new_n691), .ZN(new_n692));
  OAI21_X1  g267(.A(new_n690), .B1(new_n688), .B2(new_n691), .ZN(new_n693));
  NAND2_X1  g268(.A1(new_n692), .A2(new_n693), .ZN(G229));
  MUX2_X1   g269(.A(G5), .B(G301), .S(G16), .Z(new_n695));
  INV_X1    g270(.A(G1961), .ZN(new_n696));
  XNOR2_X1  g271(.A(new_n695), .B(new_n696), .ZN(new_n697));
  INV_X1    g272(.A(KEYINPUT30), .ZN(new_n698));
  AND2_X1   g273(.A1(new_n698), .A2(G28), .ZN(new_n699));
  INV_X1    g274(.A(G29), .ZN(new_n700));
  OAI21_X1  g275(.A(new_n700), .B1(new_n698), .B2(G28), .ZN(new_n701));
  AND2_X1   g276(.A1(KEYINPUT31), .A2(G11), .ZN(new_n702));
  NOR2_X1   g277(.A1(KEYINPUT31), .A2(G11), .ZN(new_n703));
  OAI22_X1  g278(.A1(new_n699), .A2(new_n701), .B1(new_n702), .B2(new_n703), .ZN(new_n704));
  AOI21_X1  g279(.A(new_n704), .B1(new_n626), .B2(G29), .ZN(new_n705));
  NAND3_X1  g280(.A1(new_n462), .A2(G103), .A3(G2104), .ZN(new_n706));
  XNOR2_X1  g281(.A(new_n706), .B(KEYINPUT25), .ZN(new_n707));
  NAND2_X1  g282(.A1(new_n614), .A2(G127), .ZN(new_n708));
  NAND2_X1  g283(.A1(G115), .A2(G2104), .ZN(new_n709));
  AOI21_X1  g284(.A(new_n462), .B1(new_n708), .B2(new_n709), .ZN(new_n710));
  AOI211_X1 g285(.A(new_n707), .B(new_n710), .C1(G139), .C2(new_n478), .ZN(new_n711));
  NAND2_X1  g286(.A1(new_n711), .A2(G29), .ZN(new_n712));
  NOR2_X1   g287(.A1(G29), .A2(G33), .ZN(new_n713));
  XOR2_X1   g288(.A(new_n713), .B(KEYINPUT101), .Z(new_n714));
  NAND2_X1  g289(.A1(new_n712), .A2(new_n714), .ZN(new_n715));
  INV_X1    g290(.A(G2072), .ZN(new_n716));
  OAI21_X1  g291(.A(new_n705), .B1(new_n715), .B2(new_n716), .ZN(new_n717));
  INV_X1    g292(.A(G1966), .ZN(new_n718));
  INV_X1    g293(.A(G21), .ZN(new_n719));
  NOR2_X1   g294(.A1(new_n719), .A2(G16), .ZN(new_n720));
  AOI21_X1  g295(.A(new_n720), .B1(G286), .B2(G16), .ZN(new_n721));
  AOI21_X1  g296(.A(new_n717), .B1(new_n718), .B2(new_n721), .ZN(new_n722));
  OAI211_X1 g297(.A(new_n697), .B(new_n722), .C1(new_n718), .C2(new_n721), .ZN(new_n723));
  NAND2_X1  g298(.A1(new_n700), .A2(G35), .ZN(new_n724));
  OAI21_X1  g299(.A(new_n724), .B1(G162), .B2(new_n700), .ZN(new_n725));
  XOR2_X1   g300(.A(new_n725), .B(KEYINPUT29), .Z(new_n726));
  INV_X1    g301(.A(new_n726), .ZN(new_n727));
  INV_X1    g302(.A(KEYINPUT103), .ZN(new_n728));
  NAND2_X1  g303(.A1(new_n700), .A2(G27), .ZN(new_n729));
  OAI21_X1  g304(.A(new_n729), .B1(G164), .B2(new_n700), .ZN(new_n730));
  XNOR2_X1  g305(.A(new_n730), .B(G2078), .ZN(new_n731));
  AOI22_X1  g306(.A1(new_n727), .A2(G2090), .B1(new_n728), .B2(new_n731), .ZN(new_n732));
  XOR2_X1   g307(.A(KEYINPUT95), .B(G16), .Z(new_n733));
  NAND2_X1  g308(.A1(new_n733), .A2(G20), .ZN(new_n734));
  XOR2_X1   g309(.A(new_n734), .B(KEYINPUT104), .Z(new_n735));
  XNOR2_X1  g310(.A(new_n735), .B(KEYINPUT23), .ZN(new_n736));
  AOI21_X1  g311(.A(new_n736), .B1(G16), .B2(G299), .ZN(new_n737));
  XNOR2_X1  g312(.A(new_n737), .B(G1956), .ZN(new_n738));
  INV_X1    g313(.A(new_n733), .ZN(new_n739));
  NOR2_X1   g314(.A1(new_n739), .A2(G19), .ZN(new_n740));
  AOI21_X1  g315(.A(new_n740), .B1(new_n546), .B2(new_n739), .ZN(new_n741));
  NAND2_X1  g316(.A1(new_n741), .A2(G1341), .ZN(new_n742));
  NAND3_X1  g317(.A1(new_n732), .A2(new_n738), .A3(new_n742), .ZN(new_n743));
  INV_X1    g318(.A(G34), .ZN(new_n744));
  AND2_X1   g319(.A1(new_n744), .A2(KEYINPUT24), .ZN(new_n745));
  NOR2_X1   g320(.A1(new_n744), .A2(KEYINPUT24), .ZN(new_n746));
  OAI21_X1  g321(.A(new_n700), .B1(new_n745), .B2(new_n746), .ZN(new_n747));
  OAI21_X1  g322(.A(new_n747), .B1(G160), .B2(new_n700), .ZN(new_n748));
  XNOR2_X1  g323(.A(new_n748), .B(G2084), .ZN(new_n749));
  AOI21_X1  g324(.A(new_n749), .B1(new_n715), .B2(new_n716), .ZN(new_n750));
  OAI21_X1  g325(.A(new_n750), .B1(G1341), .B2(new_n741), .ZN(new_n751));
  OAI22_X1  g326(.A1(new_n727), .A2(G2090), .B1(new_n728), .B2(new_n731), .ZN(new_n752));
  NOR4_X1   g327(.A1(new_n723), .A2(new_n743), .A3(new_n751), .A4(new_n752), .ZN(new_n753));
  NAND2_X1  g328(.A1(new_n597), .A2(G16), .ZN(new_n754));
  OAI21_X1  g329(.A(new_n754), .B1(G4), .B2(G16), .ZN(new_n755));
  INV_X1    g330(.A(G1348), .ZN(new_n756));
  OR2_X1    g331(.A1(new_n755), .A2(new_n756), .ZN(new_n757));
  NAND2_X1  g332(.A1(new_n700), .A2(G26), .ZN(new_n758));
  XOR2_X1   g333(.A(new_n758), .B(KEYINPUT28), .Z(new_n759));
  NOR2_X1   g334(.A1(G104), .A2(G2105), .ZN(new_n760));
  XNOR2_X1  g335(.A(new_n760), .B(KEYINPUT97), .ZN(new_n761));
  OAI211_X1 g336(.A(new_n761), .B(G2104), .C1(G116), .C2(new_n462), .ZN(new_n762));
  INV_X1    g337(.A(KEYINPUT98), .ZN(new_n763));
  XNOR2_X1  g338(.A(new_n762), .B(new_n763), .ZN(new_n764));
  AOI22_X1  g339(.A1(G128), .A2(new_n481), .B1(new_n478), .B2(G140), .ZN(new_n765));
  NAND2_X1  g340(.A1(new_n764), .A2(new_n765), .ZN(new_n766));
  OR2_X1    g341(.A1(new_n766), .A2(KEYINPUT99), .ZN(new_n767));
  NAND2_X1  g342(.A1(new_n766), .A2(KEYINPUT99), .ZN(new_n768));
  NAND2_X1  g343(.A1(new_n767), .A2(new_n768), .ZN(new_n769));
  AOI21_X1  g344(.A(new_n759), .B1(new_n769), .B2(G29), .ZN(new_n770));
  XNOR2_X1  g345(.A(KEYINPUT100), .B(G2067), .ZN(new_n771));
  NOR2_X1   g346(.A1(new_n770), .A2(new_n771), .ZN(new_n772));
  NAND2_X1  g347(.A1(new_n770), .A2(new_n771), .ZN(new_n773));
  XOR2_X1   g348(.A(KEYINPUT27), .B(G1996), .Z(new_n774));
  NAND2_X1  g349(.A1(new_n700), .A2(G32), .ZN(new_n775));
  AOI22_X1  g350(.A1(new_n478), .A2(G141), .B1(G105), .B2(new_n469), .ZN(new_n776));
  NAND2_X1  g351(.A1(new_n481), .A2(G129), .ZN(new_n777));
  NAND3_X1  g352(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n778));
  XOR2_X1   g353(.A(new_n778), .B(KEYINPUT26), .Z(new_n779));
  NAND3_X1  g354(.A1(new_n776), .A2(new_n777), .A3(new_n779), .ZN(new_n780));
  INV_X1    g355(.A(new_n780), .ZN(new_n781));
  OAI21_X1  g356(.A(new_n775), .B1(new_n781), .B2(new_n700), .ZN(new_n782));
  INV_X1    g357(.A(KEYINPUT102), .ZN(new_n783));
  AOI21_X1  g358(.A(new_n774), .B1(new_n782), .B2(new_n783), .ZN(new_n784));
  NOR2_X1   g359(.A1(new_n782), .A2(new_n783), .ZN(new_n785));
  XOR2_X1   g360(.A(new_n784), .B(new_n785), .Z(new_n786));
  NAND2_X1  g361(.A1(new_n773), .A2(new_n786), .ZN(new_n787));
  AOI211_X1 g362(.A(new_n772), .B(new_n787), .C1(new_n756), .C2(new_n755), .ZN(new_n788));
  NAND3_X1  g363(.A1(new_n753), .A2(new_n757), .A3(new_n788), .ZN(new_n789));
  NOR2_X1   g364(.A1(new_n739), .A2(G22), .ZN(new_n790));
  AOI21_X1  g365(.A(new_n790), .B1(G166), .B2(new_n739), .ZN(new_n791));
  INV_X1    g366(.A(G1971), .ZN(new_n792));
  XNOR2_X1  g367(.A(new_n791), .B(new_n792), .ZN(new_n793));
  XOR2_X1   g368(.A(KEYINPUT32), .B(G1981), .Z(new_n794));
  INV_X1    g369(.A(G6), .ZN(new_n795));
  NOR2_X1   g370(.A1(new_n795), .A2(G16), .ZN(new_n796));
  AOI21_X1  g371(.A(new_n796), .B1(G305), .B2(G16), .ZN(new_n797));
  AOI22_X1  g372(.A1(new_n793), .A2(KEYINPUT96), .B1(new_n794), .B2(new_n797), .ZN(new_n798));
  OAI21_X1  g373(.A(new_n798), .B1(KEYINPUT96), .B2(new_n793), .ZN(new_n799));
  INV_X1    g374(.A(G23), .ZN(new_n800));
  NOR2_X1   g375(.A1(new_n800), .A2(G16), .ZN(new_n801));
  AOI21_X1  g376(.A(new_n801), .B1(G288), .B2(G16), .ZN(new_n802));
  XOR2_X1   g377(.A(KEYINPUT33), .B(G1976), .Z(new_n803));
  XNOR2_X1  g378(.A(new_n802), .B(new_n803), .ZN(new_n804));
  OAI21_X1  g379(.A(new_n804), .B1(new_n797), .B2(new_n794), .ZN(new_n805));
  OR3_X1    g380(.A1(new_n799), .A2(KEYINPUT34), .A3(new_n805), .ZN(new_n806));
  OAI21_X1  g381(.A(KEYINPUT34), .B1(new_n799), .B2(new_n805), .ZN(new_n807));
  NAND2_X1  g382(.A1(new_n700), .A2(G25), .ZN(new_n808));
  XNOR2_X1  g383(.A(new_n808), .B(KEYINPUT91), .ZN(new_n809));
  NAND2_X1  g384(.A1(new_n478), .A2(G131), .ZN(new_n810));
  INV_X1    g385(.A(KEYINPUT92), .ZN(new_n811));
  XNOR2_X1  g386(.A(new_n810), .B(new_n811), .ZN(new_n812));
  OAI21_X1  g387(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n813));
  INV_X1    g388(.A(G107), .ZN(new_n814));
  AOI21_X1  g389(.A(new_n813), .B1(new_n814), .B2(G2105), .ZN(new_n815));
  AOI21_X1  g390(.A(new_n815), .B1(new_n481), .B2(G119), .ZN(new_n816));
  NAND2_X1  g391(.A1(new_n812), .A2(new_n816), .ZN(new_n817));
  XNOR2_X1  g392(.A(new_n817), .B(KEYINPUT93), .ZN(new_n818));
  OAI21_X1  g393(.A(new_n809), .B1(new_n818), .B2(new_n700), .ZN(new_n819));
  XOR2_X1   g394(.A(KEYINPUT35), .B(G1991), .Z(new_n820));
  XNOR2_X1  g395(.A(new_n820), .B(KEYINPUT94), .ZN(new_n821));
  INV_X1    g396(.A(new_n821), .ZN(new_n822));
  XNOR2_X1  g397(.A(new_n819), .B(new_n822), .ZN(new_n823));
  MUX2_X1   g398(.A(G24), .B(G290), .S(new_n739), .Z(new_n824));
  XOR2_X1   g399(.A(new_n824), .B(G1986), .Z(new_n825));
  NAND4_X1  g400(.A1(new_n806), .A2(new_n807), .A3(new_n823), .A4(new_n825), .ZN(new_n826));
  OR2_X1    g401(.A1(new_n826), .A2(KEYINPUT36), .ZN(new_n827));
  NAND2_X1  g402(.A1(new_n826), .A2(KEYINPUT36), .ZN(new_n828));
  AOI21_X1  g403(.A(new_n789), .B1(new_n827), .B2(new_n828), .ZN(G311));
  INV_X1    g404(.A(G311), .ZN(G150));
  NAND2_X1  g405(.A1(new_n597), .A2(G559), .ZN(new_n831));
  XNOR2_X1  g406(.A(new_n831), .B(KEYINPUT38), .ZN(new_n832));
  NAND2_X1  g407(.A1(new_n500), .A2(G55), .ZN(new_n833));
  INV_X1    g408(.A(G93), .ZN(new_n834));
  OAI21_X1  g409(.A(new_n833), .B1(new_n513), .B2(new_n834), .ZN(new_n835));
  NAND2_X1  g410(.A1(new_n517), .A2(G67), .ZN(new_n836));
  NAND2_X1  g411(.A1(G80), .A2(G543), .ZN(new_n837));
  AOI21_X1  g412(.A(new_n516), .B1(new_n836), .B2(new_n837), .ZN(new_n838));
  NOR2_X1   g413(.A1(new_n835), .A2(new_n838), .ZN(new_n839));
  XNOR2_X1  g414(.A(new_n839), .B(new_n546), .ZN(new_n840));
  XNOR2_X1  g415(.A(new_n832), .B(new_n840), .ZN(new_n841));
  INV_X1    g416(.A(KEYINPUT39), .ZN(new_n842));
  AOI21_X1  g417(.A(G860), .B1(new_n841), .B2(new_n842), .ZN(new_n843));
  OAI21_X1  g418(.A(new_n843), .B1(new_n842), .B2(new_n841), .ZN(new_n844));
  INV_X1    g419(.A(new_n839), .ZN(new_n845));
  NAND2_X1  g420(.A1(new_n845), .A2(G860), .ZN(new_n846));
  XOR2_X1   g421(.A(new_n846), .B(KEYINPUT37), .Z(new_n847));
  NAND2_X1  g422(.A1(new_n844), .A2(new_n847), .ZN(new_n848));
  NAND2_X1  g423(.A1(new_n848), .A2(KEYINPUT105), .ZN(new_n849));
  INV_X1    g424(.A(KEYINPUT105), .ZN(new_n850));
  NAND3_X1  g425(.A1(new_n844), .A2(new_n850), .A3(new_n847), .ZN(new_n851));
  NAND2_X1  g426(.A1(new_n849), .A2(new_n851), .ZN(G145));
  INV_X1    g427(.A(KEYINPUT40), .ZN(new_n853));
  XNOR2_X1  g428(.A(new_n818), .B(KEYINPUT107), .ZN(new_n854));
  NAND2_X1  g429(.A1(new_n854), .A2(new_n616), .ZN(new_n855));
  XNOR2_X1  g430(.A(new_n711), .B(new_n780), .ZN(new_n856));
  INV_X1    g431(.A(new_n856), .ZN(new_n857));
  OR2_X1    g432(.A1(new_n818), .A2(KEYINPUT107), .ZN(new_n858));
  INV_X1    g433(.A(new_n616), .ZN(new_n859));
  NAND2_X1  g434(.A1(new_n818), .A2(KEYINPUT107), .ZN(new_n860));
  NAND3_X1  g435(.A1(new_n858), .A2(new_n859), .A3(new_n860), .ZN(new_n861));
  NAND3_X1  g436(.A1(new_n855), .A2(new_n857), .A3(new_n861), .ZN(new_n862));
  INV_X1    g437(.A(new_n862), .ZN(new_n863));
  AOI21_X1  g438(.A(new_n857), .B1(new_n855), .B2(new_n861), .ZN(new_n864));
  NOR2_X1   g439(.A1(new_n863), .A2(new_n864), .ZN(new_n865));
  INV_X1    g440(.A(new_n769), .ZN(new_n866));
  NAND2_X1  g441(.A1(new_n866), .A2(G164), .ZN(new_n867));
  INV_X1    g442(.A(new_n497), .ZN(new_n868));
  AOI21_X1  g443(.A(new_n496), .B1(new_n614), .B2(new_n493), .ZN(new_n869));
  OAI211_X1 g444(.A(new_n490), .B(new_n489), .C1(new_n868), .C2(new_n869), .ZN(new_n870));
  NAND2_X1  g445(.A1(new_n769), .A2(new_n870), .ZN(new_n871));
  NAND2_X1  g446(.A1(new_n478), .A2(G142), .ZN(new_n872));
  NOR2_X1   g447(.A1(new_n462), .A2(G118), .ZN(new_n873));
  OAI21_X1  g448(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n874));
  AND3_X1   g449(.A1(new_n481), .A2(KEYINPUT106), .A3(G130), .ZN(new_n875));
  AOI21_X1  g450(.A(KEYINPUT106), .B1(new_n481), .B2(G130), .ZN(new_n876));
  OAI221_X1 g451(.A(new_n872), .B1(new_n873), .B2(new_n874), .C1(new_n875), .C2(new_n876), .ZN(new_n877));
  AND3_X1   g452(.A1(new_n867), .A2(new_n871), .A3(new_n877), .ZN(new_n878));
  AOI21_X1  g453(.A(new_n877), .B1(new_n867), .B2(new_n871), .ZN(new_n879));
  NOR2_X1   g454(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  NAND2_X1  g455(.A1(new_n865), .A2(new_n880), .ZN(new_n881));
  XNOR2_X1  g456(.A(G162), .B(G160), .ZN(new_n882));
  XNOR2_X1  g457(.A(new_n882), .B(new_n627), .ZN(new_n883));
  OAI22_X1  g458(.A1(new_n863), .A2(new_n864), .B1(new_n878), .B2(new_n879), .ZN(new_n884));
  NAND3_X1  g459(.A1(new_n881), .A2(new_n883), .A3(new_n884), .ZN(new_n885));
  INV_X1    g460(.A(G37), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n885), .A2(new_n886), .ZN(new_n887));
  AOI21_X1  g462(.A(new_n883), .B1(new_n881), .B2(new_n884), .ZN(new_n888));
  OAI21_X1  g463(.A(new_n853), .B1(new_n887), .B2(new_n888), .ZN(new_n889));
  INV_X1    g464(.A(new_n888), .ZN(new_n890));
  NAND4_X1  g465(.A1(new_n890), .A2(KEYINPUT40), .A3(new_n886), .A4(new_n885), .ZN(new_n891));
  AND2_X1   g466(.A1(new_n889), .A2(new_n891), .ZN(G395));
  XNOR2_X1  g467(.A(new_n607), .B(G299), .ZN(new_n893));
  INV_X1    g468(.A(KEYINPUT41), .ZN(new_n894));
  NAND2_X1  g469(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  OR2_X1    g470(.A1(new_n607), .A2(G299), .ZN(new_n896));
  NAND2_X1  g471(.A1(new_n607), .A2(G299), .ZN(new_n897));
  NAND3_X1  g472(.A1(new_n896), .A2(KEYINPUT41), .A3(new_n897), .ZN(new_n898));
  NAND2_X1  g473(.A1(new_n895), .A2(new_n898), .ZN(new_n899));
  XNOR2_X1  g474(.A(new_n839), .B(new_n545), .ZN(new_n900));
  AOI21_X1  g475(.A(new_n900), .B1(new_n608), .B2(new_n609), .ZN(new_n901));
  INV_X1    g476(.A(new_n901), .ZN(new_n902));
  NAND3_X1  g477(.A1(new_n608), .A2(new_n609), .A3(new_n900), .ZN(new_n903));
  NAND3_X1  g478(.A1(new_n899), .A2(new_n902), .A3(new_n903), .ZN(new_n904));
  INV_X1    g479(.A(new_n903), .ZN(new_n905));
  OAI21_X1  g480(.A(new_n893), .B1(new_n905), .B2(new_n901), .ZN(new_n906));
  NAND2_X1  g481(.A1(new_n904), .A2(new_n906), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n907), .A2(KEYINPUT42), .ZN(new_n908));
  INV_X1    g483(.A(KEYINPUT42), .ZN(new_n909));
  NAND3_X1  g484(.A1(new_n904), .A2(new_n906), .A3(new_n909), .ZN(new_n910));
  XOR2_X1   g485(.A(G305), .B(G290), .Z(new_n911));
  INV_X1    g486(.A(G288), .ZN(new_n912));
  XNOR2_X1  g487(.A(G166), .B(new_n912), .ZN(new_n913));
  XNOR2_X1  g488(.A(new_n911), .B(new_n913), .ZN(new_n914));
  INV_X1    g489(.A(new_n914), .ZN(new_n915));
  NOR2_X1   g490(.A1(new_n915), .A2(KEYINPUT108), .ZN(new_n916));
  AND3_X1   g491(.A1(new_n908), .A2(new_n910), .A3(new_n916), .ZN(new_n917));
  AOI21_X1  g492(.A(new_n916), .B1(new_n908), .B2(new_n910), .ZN(new_n918));
  OAI21_X1  g493(.A(G868), .B1(new_n917), .B2(new_n918), .ZN(new_n919));
  OAI21_X1  g494(.A(new_n919), .B1(G868), .B2(new_n839), .ZN(G295));
  OAI21_X1  g495(.A(new_n919), .B1(G868), .B2(new_n839), .ZN(G331));
  NAND2_X1  g496(.A1(new_n840), .A2(G171), .ZN(new_n922));
  NAND2_X1  g497(.A1(new_n900), .A2(G301), .ZN(new_n923));
  AOI21_X1  g498(.A(G168), .B1(new_n922), .B2(new_n923), .ZN(new_n924));
  INV_X1    g499(.A(new_n924), .ZN(new_n925));
  NAND3_X1  g500(.A1(new_n922), .A2(new_n923), .A3(G168), .ZN(new_n926));
  NAND4_X1  g501(.A1(new_n895), .A2(new_n898), .A3(new_n925), .A4(new_n926), .ZN(new_n927));
  INV_X1    g502(.A(new_n926), .ZN(new_n928));
  OAI211_X1 g503(.A(new_n897), .B(new_n896), .C1(new_n928), .C2(new_n924), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n927), .A2(new_n929), .ZN(new_n930));
  AOI21_X1  g505(.A(G37), .B1(new_n930), .B2(new_n914), .ZN(new_n931));
  NAND3_X1  g506(.A1(new_n927), .A2(new_n915), .A3(new_n929), .ZN(new_n932));
  NAND2_X1  g507(.A1(new_n931), .A2(new_n932), .ZN(new_n933));
  NAND2_X1  g508(.A1(new_n933), .A2(KEYINPUT43), .ZN(new_n934));
  INV_X1    g509(.A(KEYINPUT43), .ZN(new_n935));
  NAND3_X1  g510(.A1(new_n931), .A2(new_n935), .A3(new_n932), .ZN(new_n936));
  NAND2_X1  g511(.A1(new_n934), .A2(new_n936), .ZN(new_n937));
  INV_X1    g512(.A(KEYINPUT44), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n937), .A2(new_n938), .ZN(new_n939));
  NAND3_X1  g514(.A1(new_n934), .A2(KEYINPUT44), .A3(new_n936), .ZN(new_n940));
  NAND2_X1  g515(.A1(new_n939), .A2(new_n940), .ZN(G397));
  INV_X1    g516(.A(KEYINPUT122), .ZN(new_n942));
  INV_X1    g517(.A(KEYINPUT117), .ZN(new_n943));
  INV_X1    g518(.A(G40), .ZN(new_n944));
  NOR3_X1   g519(.A1(new_n467), .A2(new_n471), .A3(new_n944), .ZN(new_n945));
  NOR2_X1   g520(.A1(KEYINPUT50), .A2(G1384), .ZN(new_n946));
  INV_X1    g521(.A(new_n946), .ZN(new_n947));
  OAI21_X1  g522(.A(new_n945), .B1(G164), .B2(new_n947), .ZN(new_n948));
  INV_X1    g523(.A(KEYINPUT50), .ZN(new_n949));
  INV_X1    g524(.A(G1384), .ZN(new_n950));
  AOI21_X1  g525(.A(new_n949), .B1(new_n870), .B2(new_n950), .ZN(new_n951));
  OAI21_X1  g526(.A(new_n943), .B1(new_n948), .B2(new_n951), .ZN(new_n952));
  INV_X1    g527(.A(G125), .ZN(new_n953));
  AOI21_X1  g528(.A(new_n953), .B1(new_n476), .B2(new_n477), .ZN(new_n954));
  INV_X1    g529(.A(new_n466), .ZN(new_n955));
  OAI21_X1  g530(.A(G2105), .B1(new_n954), .B2(new_n955), .ZN(new_n956));
  NAND4_X1  g531(.A1(new_n956), .A2(G40), .A3(new_n470), .A4(new_n468), .ZN(new_n957));
  AOI21_X1  g532(.A(new_n957), .B1(new_n870), .B2(new_n946), .ZN(new_n958));
  OAI21_X1  g533(.A(KEYINPUT50), .B1(G164), .B2(G1384), .ZN(new_n959));
  NAND3_X1  g534(.A1(new_n958), .A2(new_n959), .A3(KEYINPUT117), .ZN(new_n960));
  NAND3_X1  g535(.A1(new_n952), .A2(new_n960), .A3(new_n696), .ZN(new_n961));
  NAND2_X1  g536(.A1(new_n870), .A2(new_n950), .ZN(new_n962));
  INV_X1    g537(.A(KEYINPUT45), .ZN(new_n963));
  AOI21_X1  g538(.A(new_n957), .B1(new_n962), .B2(new_n963), .ZN(new_n964));
  INV_X1    g539(.A(G2078), .ZN(new_n965));
  NAND3_X1  g540(.A1(new_n870), .A2(KEYINPUT45), .A3(new_n950), .ZN(new_n966));
  NAND4_X1  g541(.A1(new_n964), .A2(KEYINPUT53), .A3(new_n965), .A4(new_n966), .ZN(new_n967));
  OAI21_X1  g542(.A(new_n963), .B1(G164), .B2(G1384), .ZN(new_n968));
  NAND4_X1  g543(.A1(new_n968), .A2(new_n965), .A3(new_n945), .A4(new_n966), .ZN(new_n969));
  INV_X1    g544(.A(KEYINPUT53), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n969), .A2(new_n970), .ZN(new_n971));
  NAND3_X1  g546(.A1(new_n961), .A2(new_n967), .A3(new_n971), .ZN(new_n972));
  NAND2_X1  g547(.A1(new_n972), .A2(G171), .ZN(new_n973));
  NAND4_X1  g548(.A1(new_n961), .A2(G301), .A3(new_n971), .A4(new_n967), .ZN(new_n974));
  NAND2_X1  g549(.A1(new_n973), .A2(new_n974), .ZN(new_n975));
  INV_X1    g550(.A(KEYINPUT54), .ZN(new_n976));
  AOI21_X1  g551(.A(new_n976), .B1(new_n974), .B2(KEYINPUT121), .ZN(new_n977));
  NAND2_X1  g552(.A1(new_n975), .A2(new_n977), .ZN(new_n978));
  OAI211_X1 g553(.A(new_n973), .B(new_n974), .C1(KEYINPUT121), .C2(new_n976), .ZN(new_n979));
  NAND2_X1  g554(.A1(new_n978), .A2(new_n979), .ZN(new_n980));
  INV_X1    g555(.A(KEYINPUT49), .ZN(new_n981));
  AOI22_X1  g556(.A1(new_n512), .A2(G86), .B1(G48), .B2(new_n500), .ZN(new_n982));
  AOI21_X1  g557(.A(new_n680), .B1(new_n576), .B2(new_n982), .ZN(new_n983));
  NAND2_X1  g558(.A1(new_n572), .A2(G651), .ZN(new_n984));
  NAND2_X1  g559(.A1(new_n984), .A2(KEYINPUT79), .ZN(new_n985));
  NAND3_X1  g560(.A1(new_n572), .A2(new_n573), .A3(G651), .ZN(new_n986));
  AND4_X1   g561(.A1(new_n680), .A2(new_n581), .A3(new_n985), .A4(new_n986), .ZN(new_n987));
  OAI21_X1  g562(.A(new_n981), .B1(new_n983), .B2(new_n987), .ZN(new_n988));
  NAND3_X1  g563(.A1(new_n576), .A2(new_n680), .A3(new_n581), .ZN(new_n989));
  NAND3_X1  g564(.A1(new_n985), .A2(new_n982), .A3(new_n986), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n990), .A2(G1981), .ZN(new_n991));
  NAND3_X1  g566(.A1(new_n989), .A2(new_n991), .A3(KEYINPUT49), .ZN(new_n992));
  NAND2_X1  g567(.A1(new_n495), .A2(new_n497), .ZN(new_n993));
  AND2_X1   g568(.A1(new_n489), .A2(new_n490), .ZN(new_n994));
  AOI21_X1  g569(.A(G1384), .B1(new_n993), .B2(new_n994), .ZN(new_n995));
  NAND2_X1  g570(.A1(new_n995), .A2(new_n945), .ZN(new_n996));
  NAND2_X1  g571(.A1(new_n996), .A2(G8), .ZN(new_n997));
  INV_X1    g572(.A(new_n997), .ZN(new_n998));
  NAND3_X1  g573(.A1(new_n988), .A2(new_n992), .A3(new_n998), .ZN(new_n999));
  NAND2_X1  g574(.A1(new_n912), .A2(G1976), .ZN(new_n1000));
  NAND3_X1  g575(.A1(new_n998), .A2(KEYINPUT112), .A3(new_n1000), .ZN(new_n1001));
  XNOR2_X1  g576(.A(KEYINPUT111), .B(G1976), .ZN(new_n1002));
  NAND4_X1  g577(.A1(new_n996), .A2(G8), .A3(G288), .A4(new_n1002), .ZN(new_n1003));
  INV_X1    g578(.A(KEYINPUT52), .ZN(new_n1004));
  NAND3_X1  g579(.A1(new_n1001), .A2(new_n1003), .A3(new_n1004), .ZN(new_n1005));
  NAND2_X1  g580(.A1(new_n1003), .A2(new_n1004), .ZN(new_n1006));
  NAND4_X1  g581(.A1(new_n1006), .A2(KEYINPUT112), .A3(new_n998), .A4(new_n1000), .ZN(new_n1007));
  NAND2_X1  g582(.A1(new_n1005), .A2(new_n1007), .ZN(new_n1008));
  AOI21_X1  g583(.A(G1971), .B1(new_n964), .B2(new_n966), .ZN(new_n1009));
  NAND2_X1  g584(.A1(new_n870), .A2(new_n946), .ZN(new_n1010));
  OAI211_X1 g585(.A(new_n1010), .B(new_n945), .C1(new_n995), .C2(new_n949), .ZN(new_n1011));
  NOR2_X1   g586(.A1(new_n1011), .A2(G2090), .ZN(new_n1012));
  OAI21_X1  g587(.A(G8), .B1(new_n1009), .B2(new_n1012), .ZN(new_n1013));
  OAI21_X1  g588(.A(G8), .B1(new_n515), .B2(new_n520), .ZN(new_n1014));
  XNOR2_X1  g589(.A(new_n1014), .B(KEYINPUT55), .ZN(new_n1015));
  NAND2_X1  g590(.A1(new_n1013), .A2(new_n1015), .ZN(new_n1016));
  NAND3_X1  g591(.A1(new_n999), .A2(new_n1008), .A3(new_n1016), .ZN(new_n1017));
  OAI21_X1  g592(.A(new_n945), .B1(new_n995), .B2(KEYINPUT45), .ZN(new_n1018));
  NOR3_X1   g593(.A1(G164), .A2(new_n963), .A3(G1384), .ZN(new_n1019));
  OAI21_X1  g594(.A(new_n792), .B1(new_n1018), .B2(new_n1019), .ZN(new_n1020));
  INV_X1    g595(.A(KEYINPUT110), .ZN(new_n1021));
  INV_X1    g596(.A(G2090), .ZN(new_n1022));
  NOR2_X1   g597(.A1(new_n948), .A2(new_n951), .ZN(new_n1023));
  AOI22_X1  g598(.A1(new_n1020), .A2(new_n1021), .B1(new_n1022), .B2(new_n1023), .ZN(new_n1024));
  NAND2_X1  g599(.A1(new_n1009), .A2(KEYINPUT110), .ZN(new_n1025));
  NAND2_X1  g600(.A1(new_n1024), .A2(new_n1025), .ZN(new_n1026));
  INV_X1    g601(.A(new_n1015), .ZN(new_n1027));
  AND3_X1   g602(.A1(new_n1026), .A2(new_n1027), .A3(G8), .ZN(new_n1028));
  NOR2_X1   g603(.A1(new_n1017), .A2(new_n1028), .ZN(new_n1029));
  INV_X1    g604(.A(G2084), .ZN(new_n1030));
  NAND4_X1  g605(.A1(new_n958), .A2(new_n959), .A3(KEYINPUT113), .A4(new_n1030), .ZN(new_n1031));
  NOR2_X1   g606(.A1(new_n1018), .A2(new_n1019), .ZN(new_n1032));
  OAI21_X1  g607(.A(new_n1031), .B1(new_n1032), .B2(G1966), .ZN(new_n1033));
  AOI21_X1  g608(.A(KEYINPUT113), .B1(new_n1023), .B2(new_n1030), .ZN(new_n1034));
  OAI21_X1  g609(.A(G8), .B1(new_n1033), .B2(new_n1034), .ZN(new_n1035));
  NAND2_X1  g610(.A1(G286), .A2(G8), .ZN(new_n1036));
  INV_X1    g611(.A(KEYINPUT120), .ZN(new_n1037));
  AOI21_X1  g612(.A(KEYINPUT51), .B1(new_n1036), .B2(new_n1037), .ZN(new_n1038));
  INV_X1    g613(.A(new_n1038), .ZN(new_n1039));
  NAND3_X1  g614(.A1(new_n1035), .A2(new_n1036), .A3(new_n1039), .ZN(new_n1040));
  INV_X1    g615(.A(KEYINPUT113), .ZN(new_n1041));
  OAI21_X1  g616(.A(new_n1041), .B1(new_n1011), .B2(G2084), .ZN(new_n1042));
  OAI211_X1 g617(.A(new_n1042), .B(new_n1031), .C1(G1966), .C2(new_n1032), .ZN(new_n1043));
  OAI211_X1 g618(.A(G8), .B(new_n1038), .C1(new_n1043), .C2(G286), .ZN(new_n1044));
  NAND3_X1  g619(.A1(new_n1043), .A2(G8), .A3(G286), .ZN(new_n1045));
  NAND3_X1  g620(.A1(new_n1040), .A2(new_n1044), .A3(new_n1045), .ZN(new_n1046));
  NAND3_X1  g621(.A1(new_n980), .A2(new_n1029), .A3(new_n1046), .ZN(new_n1047));
  XNOR2_X1  g622(.A(KEYINPUT56), .B(G2072), .ZN(new_n1048));
  NAND2_X1  g623(.A1(new_n1032), .A2(new_n1048), .ZN(new_n1049));
  INV_X1    g624(.A(G1956), .ZN(new_n1050));
  OAI211_X1 g625(.A(KEYINPUT115), .B(new_n1050), .C1(new_n948), .C2(new_n951), .ZN(new_n1051));
  INV_X1    g626(.A(new_n1051), .ZN(new_n1052));
  AOI21_X1  g627(.A(KEYINPUT115), .B1(new_n1011), .B2(new_n1050), .ZN(new_n1053));
  OAI21_X1  g628(.A(new_n1049), .B1(new_n1052), .B2(new_n1053), .ZN(new_n1054));
  INV_X1    g629(.A(KEYINPUT57), .ZN(new_n1055));
  AND3_X1   g630(.A1(new_n558), .A2(new_n562), .A3(new_n1055), .ZN(new_n1056));
  AOI21_X1  g631(.A(new_n1055), .B1(new_n558), .B2(new_n562), .ZN(new_n1057));
  NOR2_X1   g632(.A1(new_n1056), .A2(new_n1057), .ZN(new_n1058));
  INV_X1    g633(.A(new_n1058), .ZN(new_n1059));
  NAND2_X1  g634(.A1(new_n1054), .A2(new_n1059), .ZN(new_n1060));
  OAI211_X1 g635(.A(new_n1058), .B(new_n1049), .C1(new_n1052), .C2(new_n1053), .ZN(new_n1061));
  NOR2_X1   g636(.A1(new_n1061), .A2(KEYINPUT116), .ZN(new_n1062));
  INV_X1    g637(.A(KEYINPUT116), .ZN(new_n1063));
  INV_X1    g638(.A(new_n1048), .ZN(new_n1064));
  NOR3_X1   g639(.A1(new_n1018), .A2(new_n1019), .A3(new_n1064), .ZN(new_n1065));
  OAI21_X1  g640(.A(new_n1050), .B1(new_n948), .B2(new_n951), .ZN(new_n1066));
  INV_X1    g641(.A(KEYINPUT115), .ZN(new_n1067));
  NAND2_X1  g642(.A1(new_n1066), .A2(new_n1067), .ZN(new_n1068));
  AOI21_X1  g643(.A(new_n1065), .B1(new_n1068), .B2(new_n1051), .ZN(new_n1069));
  AOI21_X1  g644(.A(new_n1063), .B1(new_n1069), .B2(new_n1058), .ZN(new_n1070));
  OAI21_X1  g645(.A(new_n1060), .B1(new_n1062), .B2(new_n1070), .ZN(new_n1071));
  INV_X1    g646(.A(KEYINPUT61), .ZN(new_n1072));
  NAND2_X1  g647(.A1(new_n1071), .A2(new_n1072), .ZN(new_n1073));
  OAI21_X1  g648(.A(KEYINPUT61), .B1(new_n1069), .B2(new_n1058), .ZN(new_n1074));
  INV_X1    g649(.A(new_n1061), .ZN(new_n1075));
  INV_X1    g650(.A(KEYINPUT59), .ZN(new_n1076));
  INV_X1    g651(.A(G1996), .ZN(new_n1077));
  NAND4_X1  g652(.A1(new_n968), .A2(new_n1077), .A3(new_n945), .A4(new_n966), .ZN(new_n1078));
  XOR2_X1   g653(.A(KEYINPUT58), .B(G1341), .Z(new_n1079));
  NAND2_X1  g654(.A1(new_n996), .A2(new_n1079), .ZN(new_n1080));
  NAND2_X1  g655(.A1(new_n1078), .A2(new_n1080), .ZN(new_n1081));
  AOI211_X1 g656(.A(KEYINPUT118), .B(new_n1076), .C1(new_n1081), .C2(new_n546), .ZN(new_n1082));
  NOR2_X1   g657(.A1(new_n1076), .A2(KEYINPUT118), .ZN(new_n1083));
  AOI211_X1 g658(.A(new_n545), .B(new_n1083), .C1(new_n1078), .C2(new_n1080), .ZN(new_n1084));
  OAI22_X1  g659(.A1(new_n1074), .A2(new_n1075), .B1(new_n1082), .B2(new_n1084), .ZN(new_n1085));
  INV_X1    g660(.A(new_n1085), .ZN(new_n1086));
  NAND3_X1  g661(.A1(new_n952), .A2(new_n960), .A3(new_n756), .ZN(new_n1087));
  INV_X1    g662(.A(G2067), .ZN(new_n1088));
  NAND3_X1  g663(.A1(new_n995), .A2(new_n1088), .A3(new_n945), .ZN(new_n1089));
  NAND2_X1  g664(.A1(new_n1087), .A2(new_n1089), .ZN(new_n1090));
  INV_X1    g665(.A(KEYINPUT60), .ZN(new_n1091));
  NAND2_X1  g666(.A1(new_n1090), .A2(new_n1091), .ZN(new_n1092));
  INV_X1    g667(.A(KEYINPUT119), .ZN(new_n1093));
  NAND3_X1  g668(.A1(new_n1092), .A2(new_n1093), .A3(new_n597), .ZN(new_n1094));
  NOR2_X1   g669(.A1(new_n1090), .A2(new_n1091), .ZN(new_n1095));
  AOI21_X1  g670(.A(KEYINPUT60), .B1(new_n1087), .B2(new_n1089), .ZN(new_n1096));
  OAI21_X1  g671(.A(KEYINPUT119), .B1(new_n1096), .B2(new_n607), .ZN(new_n1097));
  NAND3_X1  g672(.A1(new_n1094), .A2(new_n1095), .A3(new_n1097), .ZN(new_n1098));
  INV_X1    g673(.A(new_n1095), .ZN(new_n1099));
  AOI21_X1  g674(.A(new_n1093), .B1(new_n1092), .B2(new_n597), .ZN(new_n1100));
  NOR3_X1   g675(.A1(new_n1096), .A2(KEYINPUT119), .A3(new_n607), .ZN(new_n1101));
  OAI21_X1  g676(.A(new_n1099), .B1(new_n1100), .B2(new_n1101), .ZN(new_n1102));
  NAND4_X1  g677(.A1(new_n1073), .A2(new_n1086), .A3(new_n1098), .A4(new_n1102), .ZN(new_n1103));
  NOR2_X1   g678(.A1(new_n1062), .A2(new_n1070), .ZN(new_n1104));
  NAND2_X1  g679(.A1(new_n597), .A2(new_n1090), .ZN(new_n1105));
  AOI21_X1  g680(.A(new_n1104), .B1(new_n1105), .B2(new_n1060), .ZN(new_n1106));
  INV_X1    g681(.A(new_n1106), .ZN(new_n1107));
  AOI21_X1  g682(.A(new_n1047), .B1(new_n1103), .B2(new_n1107), .ZN(new_n1108));
  NOR2_X1   g683(.A1(new_n1035), .A2(G286), .ZN(new_n1109));
  AOI21_X1  g684(.A(KEYINPUT63), .B1(new_n1013), .B2(new_n1015), .ZN(new_n1110));
  INV_X1    g685(.A(G8), .ZN(new_n1111));
  AOI21_X1  g686(.A(new_n1111), .B1(new_n1024), .B2(new_n1025), .ZN(new_n1112));
  AOI22_X1  g687(.A1(new_n1109), .A2(new_n1110), .B1(new_n1027), .B2(new_n1112), .ZN(new_n1113));
  NAND2_X1  g688(.A1(new_n989), .A2(new_n991), .ZN(new_n1114));
  AOI21_X1  g689(.A(new_n997), .B1(new_n1114), .B2(new_n981), .ZN(new_n1115));
  AOI22_X1  g690(.A1(new_n1115), .A2(new_n992), .B1(new_n1005), .B2(new_n1007), .ZN(new_n1116));
  INV_X1    g691(.A(new_n1116), .ZN(new_n1117));
  OR2_X1    g692(.A1(new_n1113), .A2(new_n1117), .ZN(new_n1118));
  OR2_X1    g693(.A1(G288), .A2(G1976), .ZN(new_n1119));
  AOI21_X1  g694(.A(new_n1119), .B1(new_n1115), .B2(new_n992), .ZN(new_n1120));
  OAI21_X1  g695(.A(new_n998), .B1(new_n1120), .B2(new_n987), .ZN(new_n1121));
  NAND2_X1  g696(.A1(new_n1116), .A2(new_n1109), .ZN(new_n1122));
  NAND2_X1  g697(.A1(new_n1112), .A2(KEYINPUT114), .ZN(new_n1123));
  NAND2_X1  g698(.A1(new_n1026), .A2(G8), .ZN(new_n1124));
  INV_X1    g699(.A(KEYINPUT114), .ZN(new_n1125));
  AOI21_X1  g700(.A(new_n1027), .B1(new_n1124), .B2(new_n1125), .ZN(new_n1126));
  AOI21_X1  g701(.A(new_n1122), .B1(new_n1123), .B2(new_n1126), .ZN(new_n1127));
  INV_X1    g702(.A(KEYINPUT63), .ZN(new_n1128));
  OAI211_X1 g703(.A(new_n1118), .B(new_n1121), .C1(new_n1127), .C2(new_n1128), .ZN(new_n1129));
  OAI21_X1  g704(.A(new_n942), .B1(new_n1108), .B2(new_n1129), .ZN(new_n1130));
  NAND2_X1  g705(.A1(new_n1126), .A2(new_n1123), .ZN(new_n1131));
  AND3_X1   g706(.A1(new_n1109), .A2(new_n999), .A3(new_n1008), .ZN(new_n1132));
  AOI21_X1  g707(.A(new_n1128), .B1(new_n1131), .B2(new_n1132), .ZN(new_n1133));
  OAI21_X1  g708(.A(new_n1121), .B1(new_n1113), .B2(new_n1117), .ZN(new_n1134));
  NOR2_X1   g709(.A1(new_n1133), .A2(new_n1134), .ZN(new_n1135));
  NOR3_X1   g710(.A1(new_n1100), .A2(new_n1101), .A3(new_n1099), .ZN(new_n1136));
  AOI21_X1  g711(.A(new_n1095), .B1(new_n1094), .B2(new_n1097), .ZN(new_n1137));
  NOR2_X1   g712(.A1(new_n1136), .A2(new_n1137), .ZN(new_n1138));
  AOI21_X1  g713(.A(new_n1085), .B1(new_n1071), .B2(new_n1072), .ZN(new_n1139));
  AOI21_X1  g714(.A(new_n1106), .B1(new_n1138), .B2(new_n1139), .ZN(new_n1140));
  OAI211_X1 g715(.A(new_n1135), .B(KEYINPUT122), .C1(new_n1140), .C2(new_n1047), .ZN(new_n1141));
  INV_X1    g716(.A(KEYINPUT62), .ZN(new_n1142));
  NAND4_X1  g717(.A1(new_n1040), .A2(new_n1044), .A3(new_n1142), .A4(new_n1045), .ZN(new_n1143));
  INV_X1    g718(.A(new_n1143), .ZN(new_n1144));
  NAND2_X1  g719(.A1(new_n1112), .A2(new_n1027), .ZN(new_n1145));
  INV_X1    g720(.A(new_n973), .ZN(new_n1146));
  NAND4_X1  g721(.A1(new_n1116), .A2(new_n1145), .A3(new_n1146), .A4(new_n1016), .ZN(new_n1147));
  OAI21_X1  g722(.A(KEYINPUT123), .B1(new_n1144), .B2(new_n1147), .ZN(new_n1148));
  INV_X1    g723(.A(KEYINPUT123), .ZN(new_n1149));
  NAND4_X1  g724(.A1(new_n1029), .A2(new_n1149), .A3(new_n1143), .A4(new_n1146), .ZN(new_n1150));
  NAND2_X1  g725(.A1(new_n1148), .A2(new_n1150), .ZN(new_n1151));
  AND3_X1   g726(.A1(new_n1046), .A2(KEYINPUT124), .A3(KEYINPUT62), .ZN(new_n1152));
  AOI21_X1  g727(.A(KEYINPUT124), .B1(new_n1046), .B2(KEYINPUT62), .ZN(new_n1153));
  NOR2_X1   g728(.A1(new_n1152), .A2(new_n1153), .ZN(new_n1154));
  OAI21_X1  g729(.A(KEYINPUT125), .B1(new_n1151), .B2(new_n1154), .ZN(new_n1155));
  OR2_X1    g730(.A1(new_n1152), .A2(new_n1153), .ZN(new_n1156));
  INV_X1    g731(.A(KEYINPUT125), .ZN(new_n1157));
  NAND4_X1  g732(.A1(new_n1156), .A2(new_n1157), .A3(new_n1150), .A4(new_n1148), .ZN(new_n1158));
  NAND4_X1  g733(.A1(new_n1130), .A2(new_n1141), .A3(new_n1155), .A4(new_n1158), .ZN(new_n1159));
  NOR2_X1   g734(.A1(new_n968), .A2(new_n957), .ZN(new_n1160));
  NAND2_X1  g735(.A1(new_n1160), .A2(new_n1077), .ZN(new_n1161));
  XOR2_X1   g736(.A(new_n1161), .B(KEYINPUT109), .Z(new_n1162));
  NOR2_X1   g737(.A1(new_n1162), .A2(new_n780), .ZN(new_n1163));
  NAND2_X1  g738(.A1(new_n866), .A2(new_n1088), .ZN(new_n1164));
  NAND2_X1  g739(.A1(new_n769), .A2(G2067), .ZN(new_n1165));
  OAI211_X1 g740(.A(new_n1164), .B(new_n1165), .C1(new_n1077), .C2(new_n781), .ZN(new_n1166));
  AOI21_X1  g741(.A(new_n1163), .B1(new_n1166), .B2(new_n1160), .ZN(new_n1167));
  AND2_X1   g742(.A1(new_n818), .A2(new_n822), .ZN(new_n1168));
  NOR2_X1   g743(.A1(new_n818), .A2(new_n822), .ZN(new_n1169));
  OAI21_X1  g744(.A(new_n1160), .B1(new_n1168), .B2(new_n1169), .ZN(new_n1170));
  NAND2_X1  g745(.A1(new_n1167), .A2(new_n1170), .ZN(new_n1171));
  XNOR2_X1  g746(.A(G290), .B(G1986), .ZN(new_n1172));
  AOI21_X1  g747(.A(new_n1171), .B1(new_n1160), .B2(new_n1172), .ZN(new_n1173));
  NAND2_X1  g748(.A1(new_n1159), .A2(new_n1173), .ZN(new_n1174));
  NAND3_X1  g749(.A1(new_n1164), .A2(new_n781), .A3(new_n1165), .ZN(new_n1175));
  NAND2_X1  g750(.A1(new_n1175), .A2(new_n1160), .ZN(new_n1176));
  AND2_X1   g751(.A1(new_n1162), .A2(KEYINPUT46), .ZN(new_n1177));
  NOR2_X1   g752(.A1(new_n1162), .A2(KEYINPUT46), .ZN(new_n1178));
  OAI21_X1  g753(.A(new_n1176), .B1(new_n1177), .B2(new_n1178), .ZN(new_n1179));
  XNOR2_X1  g754(.A(new_n1179), .B(KEYINPUT47), .ZN(new_n1180));
  NOR2_X1   g755(.A1(G290), .A2(G1986), .ZN(new_n1181));
  NAND2_X1  g756(.A1(new_n1181), .A2(new_n1160), .ZN(new_n1182));
  XNOR2_X1  g757(.A(new_n1182), .B(KEYINPUT126), .ZN(new_n1183));
  XOR2_X1   g758(.A(new_n1183), .B(KEYINPUT48), .Z(new_n1184));
  OAI21_X1  g759(.A(new_n1180), .B1(new_n1171), .B2(new_n1184), .ZN(new_n1185));
  NAND2_X1  g760(.A1(new_n1167), .A2(new_n1168), .ZN(new_n1186));
  NAND2_X1  g761(.A1(new_n1186), .A2(new_n1164), .ZN(new_n1187));
  AOI21_X1  g762(.A(new_n1185), .B1(new_n1160), .B2(new_n1187), .ZN(new_n1188));
  NAND2_X1  g763(.A1(new_n1174), .A2(new_n1188), .ZN(G329));
  assign    G231 = 1'b0;
  NAND3_X1  g764(.A1(new_n664), .A2(G319), .A3(new_n665), .ZN(new_n1191));
  OR2_X1    g765(.A1(new_n1191), .A2(KEYINPUT127), .ZN(new_n1192));
  NAND2_X1  g766(.A1(new_n1191), .A2(KEYINPUT127), .ZN(new_n1193));
  AOI22_X1  g767(.A1(new_n645), .A2(new_n647), .B1(new_n1192), .B2(new_n1193), .ZN(new_n1194));
  AND3_X1   g768(.A1(new_n692), .A2(new_n693), .A3(new_n1194), .ZN(new_n1195));
  NAND3_X1  g769(.A1(new_n890), .A2(new_n886), .A3(new_n885), .ZN(new_n1196));
  NAND3_X1  g770(.A1(new_n937), .A2(new_n1195), .A3(new_n1196), .ZN(G225));
  INV_X1    g771(.A(G225), .ZN(G308));
endmodule


