

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
         n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598,
         n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609,
         n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620,
         n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631,
         n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642,
         n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653,
         n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664,
         n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675,
         n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686,
         n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697,
         n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708,
         n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719,
         n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, n730,
         n731, n732, n733, n734, n735, n736, n737, n738, n739, n740, n741;

  NOR2_X1 U368 ( .A1(n540), .A2(n563), .ZN(n390) );
  XNOR2_X1 U369 ( .A(n397), .B(n410), .ZN(n460) );
  XNOR2_X1 U370 ( .A(n575), .B(n574), .ZN(n738) );
  XNOR2_X2 U371 ( .A(n416), .B(n415), .ZN(n498) );
  NOR2_X2 U372 ( .A1(n347), .A2(n535), .ZN(n639) );
  XNOR2_X2 U373 ( .A(n386), .B(G146), .ZN(n423) );
  XNOR2_X2 U374 ( .A(n507), .B(KEYINPUT22), .ZN(n542) );
  BUF_X1 U375 ( .A(n510), .Z(n346) );
  BUF_X1 U376 ( .A(n510), .Z(n347) );
  XNOR2_X1 U377 ( .A(n464), .B(G472), .ZN(n510) );
  NOR2_X1 U378 ( .A1(G953), .A2(G237), .ZN(n453) );
  OR2_X1 U379 ( .A1(n587), .A2(n648), .ZN(n575) );
  NOR2_X1 U380 ( .A1(n544), .A2(n506), .ZN(n494) );
  INV_X1 U381 ( .A(G125), .ZN(n386) );
  XNOR2_X1 U382 ( .A(G101), .B(KEYINPUT92), .ZN(n398) );
  XNOR2_X1 U383 ( .A(G116), .B(G113), .ZN(n399) );
  OR2_X1 U384 ( .A1(n601), .A2(n589), .ZN(n590) );
  NOR2_X1 U385 ( .A1(n378), .A2(n374), .ZN(n586) );
  XNOR2_X1 U386 ( .A(n375), .B(KEYINPUT46), .ZN(n374) );
  AND2_X1 U387 ( .A1(n367), .A2(n366), .ZN(n364) );
  INV_X1 U388 ( .A(n542), .ZN(n348) );
  XNOR2_X1 U389 ( .A(n411), .B(n460), .ZN(n634) );
  XNOR2_X1 U390 ( .A(n451), .B(n452), .ZN(n469) );
  XNOR2_X1 U391 ( .A(n432), .B(G134), .ZN(n452) );
  XNOR2_X1 U392 ( .A(n400), .B(KEYINPUT4), .ZN(n362) );
  XNOR2_X1 U393 ( .A(n399), .B(n398), .ZN(n397) );
  XNOR2_X1 U394 ( .A(n408), .B(G107), .ZN(n471) );
  XNOR2_X1 U395 ( .A(G104), .B(G110), .ZN(n408) );
  INV_X1 U396 ( .A(KEYINPUT65), .ZN(n400) );
  NAND2_X1 U397 ( .A1(n364), .A2(n363), .ZN(n349) );
  NAND2_X1 U398 ( .A1(n364), .A2(n363), .ZN(n525) );
  XNOR2_X1 U399 ( .A(n368), .B(n395), .ZN(n394) );
  NAND2_X1 U400 ( .A1(n525), .A2(n643), .ZN(n368) );
  XNOR2_X1 U401 ( .A(n686), .B(n539), .ZN(n563) );
  XNOR2_X1 U402 ( .A(n382), .B(n381), .ZN(n686) );
  INV_X1 U403 ( .A(KEYINPUT105), .ZN(n381) );
  NOR2_X1 U404 ( .A1(n651), .A2(n654), .ZN(n382) );
  XOR2_X1 U405 ( .A(G137), .B(G140), .Z(n480) );
  XNOR2_X1 U406 ( .A(n469), .B(n480), .ZN(n727) );
  XNOR2_X1 U407 ( .A(n393), .B(n392), .ZN(n391) );
  INV_X1 U408 ( .A(KEYINPUT44), .ZN(n392) );
  NAND2_X1 U409 ( .A1(n396), .A2(n394), .ZN(n393) );
  NOR2_X1 U410 ( .A1(n584), .A2(n567), .ZN(n380) );
  OR2_X1 U411 ( .A1(n566), .A2(KEYINPUT47), .ZN(n379) );
  NAND2_X1 U412 ( .A1(n377), .A2(n376), .ZN(n375) );
  INV_X1 U413 ( .A(n738), .ZN(n377) );
  XNOR2_X1 U414 ( .A(G101), .B(G146), .ZN(n470) );
  INV_X1 U415 ( .A(KEYINPUT75), .ZN(n472) );
  XNOR2_X1 U416 ( .A(n477), .B(G469), .ZN(n553) );
  XNOR2_X1 U417 ( .A(G119), .B(G110), .ZN(n481) );
  XNOR2_X1 U418 ( .A(n371), .B(n370), .ZN(n369) );
  XNOR2_X1 U419 ( .A(KEYINPUT7), .B(KEYINPUT9), .ZN(n370) );
  XNOR2_X1 U420 ( .A(n372), .B(G107), .ZN(n371) );
  INV_X1 U421 ( .A(KEYINPUT100), .ZN(n372) );
  XNOR2_X1 U422 ( .A(n434), .B(n433), .ZN(n373) );
  XNOR2_X1 U423 ( .A(G116), .B(G122), .ZN(n433) );
  XNOR2_X1 U424 ( .A(KEYINPUT70), .B(KEYINPUT10), .ZN(n422) );
  XNOR2_X1 U425 ( .A(n431), .B(n430), .ZN(n537) );
  XNOR2_X1 U426 ( .A(n429), .B(G475), .ZN(n430) );
  INV_X1 U427 ( .A(KEYINPUT88), .ZN(n395) );
  AND2_X1 U428 ( .A1(n388), .A2(n637), .ZN(n387) );
  XNOR2_X1 U429 ( .A(n390), .B(n389), .ZN(n388) );
  XNOR2_X1 U430 ( .A(G137), .B(G146), .ZN(n457) );
  INV_X1 U431 ( .A(KEYINPUT48), .ZN(n585) );
  AND2_X1 U432 ( .A1(n509), .A2(n361), .ZN(n529) );
  XNOR2_X1 U433 ( .A(G143), .B(G104), .ZN(n418) );
  XNOR2_X1 U434 ( .A(n450), .B(n417), .ZN(n421) );
  XNOR2_X1 U435 ( .A(G113), .B(G122), .ZN(n417) );
  XNOR2_X1 U436 ( .A(n727), .B(n476), .ZN(n709) );
  XNOR2_X1 U437 ( .A(n475), .B(n474), .ZN(n476) );
  NOR2_X1 U438 ( .A1(n517), .A2(n468), .ZN(n569) );
  INV_X1 U439 ( .A(KEYINPUT19), .ZN(n384) );
  XNOR2_X1 U440 ( .A(n487), .B(n486), .ZN(n721) );
  XNOR2_X1 U441 ( .A(n479), .B(n726), .ZN(n487) );
  XNOR2_X1 U442 ( .A(n373), .B(n369), .ZN(n437) );
  AND2_X1 U443 ( .A1(n609), .A2(G953), .ZN(n725) );
  XNOR2_X1 U444 ( .A(n358), .B(n357), .ZN(n396) );
  INV_X1 U445 ( .A(KEYINPUT35), .ZN(n357) );
  XNOR2_X1 U446 ( .A(n527), .B(KEYINPUT34), .ZN(n359) );
  NAND2_X1 U447 ( .A1(n348), .A2(n365), .ZN(n363) );
  NOR2_X1 U448 ( .A1(n514), .A2(n355), .ZN(n365) );
  NAND2_X1 U449 ( .A1(n348), .A2(n352), .ZN(n643) );
  XNOR2_X1 U450 ( .A(n538), .B(n383), .ZN(n654) );
  INV_X1 U451 ( .A(KEYINPUT104), .ZN(n383) );
  XNOR2_X1 U452 ( .A(n360), .B(n356), .ZN(n684) );
  AND2_X1 U453 ( .A1(G217), .A2(n491), .ZN(n350) );
  NAND2_X1 U454 ( .A1(n502), .A2(n501), .ZN(n351) );
  NOR2_X1 U455 ( .A1(n560), .A2(n524), .ZN(n352) );
  AND2_X1 U456 ( .A1(n576), .A2(n674), .ZN(n353) );
  XOR2_X1 U457 ( .A(KEYINPUT68), .B(KEYINPUT0), .Z(n354) );
  XNOR2_X1 U458 ( .A(KEYINPUT66), .B(KEYINPUT32), .ZN(n355) );
  XNOR2_X1 U459 ( .A(KEYINPUT91), .B(n526), .ZN(n356) );
  INV_X1 U460 ( .A(n396), .ZN(n737) );
  NAND2_X1 U461 ( .A1(n359), .A2(n528), .ZN(n358) );
  INV_X1 U462 ( .A(n509), .ZN(n670) );
  NAND2_X1 U463 ( .A1(n529), .A2(n541), .ZN(n360) );
  INV_X1 U464 ( .A(n671), .ZN(n361) );
  XNOR2_X1 U465 ( .A(n362), .B(n423), .ZN(n402) );
  XNOR2_X1 U466 ( .A(n450), .B(n362), .ZN(n451) );
  NAND2_X1 U467 ( .A1(n514), .A2(n355), .ZN(n366) );
  NAND2_X1 U468 ( .A1(n542), .A2(n355), .ZN(n367) );
  INV_X1 U469 ( .A(n533), .ZN(n530) );
  NAND2_X1 U470 ( .A1(n533), .A2(n353), .ZN(n507) );
  XNOR2_X2 U471 ( .A(n504), .B(n354), .ZN(n533) );
  INV_X1 U472 ( .A(n741), .ZN(n376) );
  NAND2_X1 U473 ( .A1(n380), .A2(n379), .ZN(n378) );
  INV_X1 U474 ( .A(n503), .ZN(n555) );
  XNOR2_X1 U475 ( .A(n557), .B(n384), .ZN(n503) );
  XNOR2_X2 U476 ( .A(n385), .B(KEYINPUT89), .ZN(n557) );
  NAND2_X1 U477 ( .A1(n498), .A2(n688), .ZN(n385) );
  NAND2_X1 U478 ( .A1(n391), .A2(n387), .ZN(n549) );
  INV_X1 U479 ( .A(KEYINPUT106), .ZN(n389) );
  BUF_X1 U480 ( .A(n498), .Z(n568) );
  INV_X1 U481 ( .A(KEYINPUT83), .ZN(n539) );
  INV_X1 U482 ( .A(KEYINPUT73), .ZN(n456) );
  XNOR2_X1 U483 ( .A(n457), .B(n456), .ZN(n458) );
  XNOR2_X1 U484 ( .A(n459), .B(n458), .ZN(n461) );
  XNOR2_X1 U485 ( .A(n473), .B(n472), .ZN(n474) );
  BUF_X1 U486 ( .A(n628), .Z(n666) );
  INV_X1 U487 ( .A(KEYINPUT39), .ZN(n572) );
  BUF_X1 U488 ( .A(n715), .Z(n720) );
  XNOR2_X1 U489 ( .A(n573), .B(n572), .ZN(n587) );
  INV_X1 U490 ( .A(KEYINPUT40), .ZN(n574) );
  XNOR2_X2 U491 ( .A(KEYINPUT78), .B(G143), .ZN(n401) );
  XNOR2_X2 U492 ( .A(n401), .B(G128), .ZN(n432) );
  XNOR2_X1 U493 ( .A(n402), .B(n432), .ZN(n407) );
  XOR2_X1 U494 ( .A(KEYINPUT17), .B(KEYINPUT18), .Z(n405) );
  INV_X2 U495 ( .A(G953), .ZN(n730) );
  NAND2_X1 U496 ( .A1(G224), .A2(n730), .ZN(n403) );
  XNOR2_X1 U497 ( .A(n403), .B(KEYINPUT76), .ZN(n404) );
  XNOR2_X1 U498 ( .A(n405), .B(n404), .ZN(n406) );
  XNOR2_X1 U499 ( .A(n407), .B(n406), .ZN(n412) );
  XNOR2_X1 U500 ( .A(KEYINPUT16), .B(G122), .ZN(n409) );
  XNOR2_X1 U501 ( .A(n471), .B(n409), .ZN(n411) );
  XNOR2_X1 U502 ( .A(KEYINPUT3), .B(G119), .ZN(n410) );
  XNOR2_X1 U503 ( .A(n412), .B(n634), .ZN(n604) );
  XNOR2_X1 U504 ( .A(KEYINPUT15), .B(G902), .ZN(n592) );
  INV_X1 U505 ( .A(n592), .ZN(n550) );
  OR2_X2 U506 ( .A1(n604), .A2(n550), .ZN(n416) );
  NOR2_X1 U507 ( .A1(G237), .A2(G902), .ZN(n413) );
  XNOR2_X1 U508 ( .A(n413), .B(KEYINPUT72), .ZN(n466) );
  INV_X1 U509 ( .A(n466), .ZN(n414) );
  AND2_X1 U510 ( .A1(n414), .A2(G210), .ZN(n415) );
  XOR2_X1 U511 ( .A(KEYINPUT71), .B(G131), .Z(n450) );
  XOR2_X1 U512 ( .A(KEYINPUT12), .B(KEYINPUT98), .Z(n419) );
  XNOR2_X1 U513 ( .A(n419), .B(n418), .ZN(n420) );
  XNOR2_X1 U514 ( .A(n421), .B(n420), .ZN(n428) );
  XNOR2_X1 U515 ( .A(n423), .B(n422), .ZN(n726) );
  XOR2_X1 U516 ( .A(G140), .B(KEYINPUT11), .Z(n425) );
  NAND2_X1 U517 ( .A1(G214), .A2(n453), .ZN(n424) );
  XNOR2_X1 U518 ( .A(n425), .B(n424), .ZN(n426) );
  XNOR2_X1 U519 ( .A(n726), .B(n426), .ZN(n427) );
  XNOR2_X1 U520 ( .A(n428), .B(n427), .ZN(n620) );
  NOR2_X1 U521 ( .A1(G902), .A2(n620), .ZN(n431) );
  XNOR2_X1 U522 ( .A(KEYINPUT99), .B(KEYINPUT13), .ZN(n429) );
  INV_X1 U523 ( .A(n537), .ZN(n441) );
  XNOR2_X1 U524 ( .A(KEYINPUT102), .B(KEYINPUT101), .ZN(n434) );
  NAND2_X1 U525 ( .A1(G234), .A2(n730), .ZN(n435) );
  XOR2_X1 U526 ( .A(KEYINPUT8), .B(n435), .Z(n478) );
  NAND2_X1 U527 ( .A1(G217), .A2(n478), .ZN(n436) );
  XNOR2_X1 U528 ( .A(n437), .B(n436), .ZN(n438) );
  XNOR2_X1 U529 ( .A(n452), .B(n438), .ZN(n716) );
  NOR2_X1 U530 ( .A1(G902), .A2(n716), .ZN(n440) );
  XNOR2_X1 U531 ( .A(KEYINPUT103), .B(G478), .ZN(n439) );
  XNOR2_X1 U532 ( .A(n440), .B(n439), .ZN(n536) );
  NAND2_X1 U533 ( .A1(n441), .A2(n536), .ZN(n442) );
  XOR2_X1 U534 ( .A(KEYINPUT108), .B(n442), .Z(n528) );
  NAND2_X1 U535 ( .A1(G234), .A2(G237), .ZN(n443) );
  XNOR2_X1 U536 ( .A(n443), .B(KEYINPUT14), .ZN(n445) );
  NAND2_X1 U537 ( .A1(G952), .A2(n445), .ZN(n444) );
  XNOR2_X1 U538 ( .A(KEYINPUT93), .B(n444), .ZN(n698) );
  NAND2_X1 U539 ( .A1(n698), .A2(n730), .ZN(n502) );
  INV_X1 U540 ( .A(n502), .ZN(n449) );
  NAND2_X1 U541 ( .A1(G902), .A2(n445), .ZN(n499) );
  NOR2_X1 U542 ( .A1(G900), .A2(n499), .ZN(n446) );
  NAND2_X1 U543 ( .A1(G953), .A2(n446), .ZN(n447) );
  XNOR2_X1 U544 ( .A(KEYINPUT109), .B(n447), .ZN(n448) );
  NOR2_X1 U545 ( .A1(n449), .A2(n448), .ZN(n517) );
  XOR2_X1 U546 ( .A(KEYINPUT5), .B(KEYINPUT96), .Z(n455) );
  NAND2_X1 U547 ( .A1(n453), .A2(G210), .ZN(n454) );
  XNOR2_X1 U548 ( .A(n455), .B(n454), .ZN(n459) );
  XNOR2_X1 U549 ( .A(n461), .B(n460), .ZN(n462) );
  XNOR2_X1 U550 ( .A(n469), .B(n462), .ZN(n613) );
  INV_X1 U551 ( .A(G902), .ZN(n463) );
  NAND2_X1 U552 ( .A1(n613), .A2(n463), .ZN(n464) );
  INV_X1 U553 ( .A(G214), .ZN(n465) );
  OR2_X1 U554 ( .A1(n466), .A2(n465), .ZN(n688) );
  NAND2_X1 U555 ( .A1(n346), .A2(n688), .ZN(n467) );
  XNOR2_X1 U556 ( .A(KEYINPUT30), .B(n467), .ZN(n468) );
  XNOR2_X1 U557 ( .A(n471), .B(n470), .ZN(n475) );
  NAND2_X1 U558 ( .A1(G227), .A2(n730), .ZN(n473) );
  NOR2_X1 U559 ( .A1(n709), .A2(G902), .ZN(n477) );
  NAND2_X1 U560 ( .A1(G221), .A2(n478), .ZN(n479) );
  XNOR2_X1 U561 ( .A(n481), .B(n480), .ZN(n485) );
  XOR2_X1 U562 ( .A(KEYINPUT24), .B(KEYINPUT23), .Z(n483) );
  XNOR2_X1 U563 ( .A(G128), .B(KEYINPUT74), .ZN(n482) );
  XNOR2_X1 U564 ( .A(n483), .B(n482), .ZN(n484) );
  XOR2_X1 U565 ( .A(n485), .B(n484), .Z(n486) );
  NOR2_X1 U566 ( .A1(n721), .A2(G902), .ZN(n490) );
  NAND2_X1 U567 ( .A1(G234), .A2(n592), .ZN(n488) );
  XNOR2_X1 U568 ( .A(KEYINPUT20), .B(n488), .ZN(n491) );
  XNOR2_X1 U569 ( .A(KEYINPUT25), .B(n350), .ZN(n489) );
  XNOR2_X2 U570 ( .A(n490), .B(n489), .ZN(n544) );
  AND2_X1 U571 ( .A1(n491), .A2(G221), .ZN(n493) );
  INV_X1 U572 ( .A(KEYINPUT21), .ZN(n492) );
  XNOR2_X1 U573 ( .A(n493), .B(n492), .ZN(n506) );
  XNOR2_X1 U574 ( .A(n494), .B(KEYINPUT69), .ZN(n671) );
  NOR2_X1 U575 ( .A1(n553), .A2(n671), .ZN(n495) );
  XNOR2_X1 U576 ( .A(n495), .B(KEYINPUT94), .ZN(n570) );
  AND2_X1 U577 ( .A1(n569), .A2(n570), .ZN(n496) );
  AND2_X1 U578 ( .A1(n528), .A2(n496), .ZN(n497) );
  NAND2_X1 U579 ( .A1(n568), .A2(n497), .ZN(n580) );
  XNOR2_X1 U580 ( .A(n580), .B(G143), .ZN(G45) );
  INV_X1 U581 ( .A(n499), .ZN(n500) );
  NOR2_X1 U582 ( .A1(G898), .A2(n730), .ZN(n633) );
  NAND2_X1 U583 ( .A1(n500), .A2(n633), .ZN(n501) );
  NAND2_X1 U584 ( .A1(n503), .A2(n351), .ZN(n504) );
  INV_X1 U585 ( .A(n536), .ZN(n505) );
  AND2_X1 U586 ( .A1(n537), .A2(n505), .ZN(n576) );
  INV_X1 U587 ( .A(n506), .ZN(n674) );
  INV_X1 U588 ( .A(KEYINPUT1), .ZN(n508) );
  XNOR2_X1 U589 ( .A(n553), .B(n508), .ZN(n509) );
  INV_X1 U590 ( .A(n670), .ZN(n560) );
  INV_X1 U591 ( .A(KEYINPUT6), .ZN(n511) );
  XNOR2_X1 U592 ( .A(n347), .B(n511), .ZN(n541) );
  XNOR2_X1 U593 ( .A(n541), .B(KEYINPUT77), .ZN(n512) );
  AND2_X1 U594 ( .A1(n512), .A2(n544), .ZN(n513) );
  NAND2_X1 U595 ( .A1(n560), .A2(n513), .ZN(n514) );
  XOR2_X1 U596 ( .A(G119), .B(KEYINPUT127), .Z(n515) );
  XNOR2_X1 U597 ( .A(n349), .B(n515), .ZN(G21) );
  INV_X1 U598 ( .A(n541), .ZN(n519) );
  NAND2_X1 U599 ( .A1(n544), .A2(n674), .ZN(n516) );
  NOR2_X1 U600 ( .A1(n517), .A2(n516), .ZN(n551) );
  OR2_X1 U601 ( .A1(n537), .A2(n536), .ZN(n648) );
  INV_X1 U602 ( .A(n648), .ZN(n651) );
  NAND2_X1 U603 ( .A1(n551), .A2(n651), .ZN(n518) );
  NOR2_X1 U604 ( .A1(n519), .A2(n518), .ZN(n558) );
  NAND2_X1 U605 ( .A1(n558), .A2(n688), .ZN(n520) );
  NOR2_X1 U606 ( .A1(n560), .A2(n520), .ZN(n522) );
  XNOR2_X1 U607 ( .A(KEYINPUT110), .B(KEYINPUT43), .ZN(n521) );
  XNOR2_X1 U608 ( .A(n522), .B(n521), .ZN(n523) );
  OR2_X1 U609 ( .A1(n523), .A2(n568), .ZN(n598) );
  XNOR2_X1 U610 ( .A(n598), .B(G140), .ZN(G42) );
  INV_X1 U611 ( .A(n544), .ZN(n675) );
  OR2_X1 U612 ( .A1(n347), .A2(n675), .ZN(n524) );
  XOR2_X1 U613 ( .A(KEYINPUT107), .B(KEYINPUT33), .Z(n526) );
  NOR2_X1 U614 ( .A1(n684), .A2(n530), .ZN(n527) );
  NAND2_X1 U615 ( .A1(n529), .A2(n347), .ZN(n680) );
  OR2_X1 U616 ( .A1(n680), .A2(n530), .ZN(n532) );
  XOR2_X1 U617 ( .A(KEYINPUT97), .B(KEYINPUT31), .Z(n531) );
  XNOR2_X1 U618 ( .A(n532), .B(n531), .ZN(n653) );
  NAND2_X1 U619 ( .A1(n533), .A2(n570), .ZN(n534) );
  XOR2_X1 U620 ( .A(KEYINPUT95), .B(n534), .Z(n535) );
  NOR2_X1 U621 ( .A1(n653), .A2(n639), .ZN(n540) );
  NAND2_X1 U622 ( .A1(n537), .A2(n536), .ZN(n538) );
  OR2_X1 U623 ( .A1(n542), .A2(n541), .ZN(n543) );
  XNOR2_X1 U624 ( .A(n543), .B(KEYINPUT87), .ZN(n546) );
  NOR2_X1 U625 ( .A1(n560), .A2(n544), .ZN(n545) );
  NAND2_X1 U626 ( .A1(n546), .A2(n545), .ZN(n637) );
  INV_X1 U627 ( .A(KEYINPUT64), .ZN(n547) );
  XNOR2_X1 U628 ( .A(n547), .B(KEYINPUT45), .ZN(n548) );
  XNOR2_X2 U629 ( .A(n549), .B(n548), .ZN(n628) );
  NOR2_X1 U630 ( .A1(n628), .A2(n592), .ZN(n591) );
  AND2_X1 U631 ( .A1(n347), .A2(n551), .ZN(n552) );
  XOR2_X1 U632 ( .A(KEYINPUT28), .B(n552), .Z(n554) );
  OR2_X1 U633 ( .A1(n554), .A2(n553), .ZN(n578) );
  OR2_X1 U634 ( .A1(n578), .A2(n555), .ZN(n649) );
  XNOR2_X1 U635 ( .A(n649), .B(KEYINPUT82), .ZN(n556) );
  NAND2_X1 U636 ( .A1(n556), .A2(KEYINPUT47), .ZN(n562) );
  NAND2_X1 U637 ( .A1(n558), .A2(n557), .ZN(n559) );
  XOR2_X1 U638 ( .A(KEYINPUT36), .B(n559), .Z(n561) );
  NAND2_X1 U639 ( .A1(n561), .A2(n560), .ZN(n656) );
  NAND2_X1 U640 ( .A1(n562), .A2(n656), .ZN(n567) );
  INV_X1 U641 ( .A(KEYINPUT82), .ZN(n565) );
  NOR2_X1 U642 ( .A1(n563), .A2(n649), .ZN(n564) );
  NOR2_X1 U643 ( .A1(n565), .A2(n564), .ZN(n566) );
  XOR2_X1 U644 ( .A(KEYINPUT38), .B(n568), .Z(n689) );
  AND2_X1 U645 ( .A1(n569), .A2(n689), .ZN(n571) );
  NAND2_X1 U646 ( .A1(n571), .A2(n570), .ZN(n573) );
  INV_X1 U647 ( .A(n576), .ZN(n691) );
  NAND2_X1 U648 ( .A1(n689), .A2(n688), .ZN(n685) );
  NOR2_X1 U649 ( .A1(n691), .A2(n685), .ZN(n577) );
  XNOR2_X1 U650 ( .A(n577), .B(KEYINPUT41), .ZN(n703) );
  NOR2_X1 U651 ( .A1(n578), .A2(n703), .ZN(n579) );
  XNOR2_X1 U652 ( .A(n579), .B(KEYINPUT42), .ZN(n741) );
  XNOR2_X1 U653 ( .A(n580), .B(KEYINPUT84), .ZN(n582) );
  NAND2_X1 U654 ( .A1(KEYINPUT47), .A2(n686), .ZN(n581) );
  NAND2_X1 U655 ( .A1(n582), .A2(n581), .ZN(n583) );
  XNOR2_X1 U656 ( .A(KEYINPUT80), .B(n583), .ZN(n584) );
  XNOR2_X1 U657 ( .A(n586), .B(n585), .ZN(n601) );
  INV_X1 U658 ( .A(n654), .ZN(n645) );
  NOR2_X1 U659 ( .A1(n645), .A2(n587), .ZN(n588) );
  XNOR2_X1 U660 ( .A(n588), .B(KEYINPUT111), .ZN(n739) );
  NAND2_X1 U661 ( .A1(n739), .A2(n598), .ZN(n589) );
  INV_X1 U662 ( .A(n590), .ZN(n729) );
  AND2_X1 U663 ( .A1(n591), .A2(n729), .ZN(n596) );
  XOR2_X1 U664 ( .A(KEYINPUT86), .B(n592), .Z(n593) );
  NAND2_X1 U665 ( .A1(n593), .A2(KEYINPUT2), .ZN(n594) );
  XNOR2_X1 U666 ( .A(n594), .B(KEYINPUT67), .ZN(n595) );
  NOR2_X1 U667 ( .A1(n596), .A2(n595), .ZN(n603) );
  NAND2_X1 U668 ( .A1(KEYINPUT2), .A2(n739), .ZN(n597) );
  XNOR2_X1 U669 ( .A(KEYINPUT79), .B(n597), .ZN(n599) );
  NAND2_X1 U670 ( .A1(n599), .A2(n598), .ZN(n600) );
  NOR2_X1 U671 ( .A1(n601), .A2(n600), .ZN(n602) );
  INV_X1 U672 ( .A(n628), .ZN(n660) );
  AND2_X1 U673 ( .A1(n602), .A2(n660), .ZN(n659) );
  NOR2_X4 U674 ( .A1(n603), .A2(n659), .ZN(n715) );
  NAND2_X1 U675 ( .A1(n715), .A2(G210), .ZN(n608) );
  XNOR2_X1 U676 ( .A(KEYINPUT81), .B(KEYINPUT54), .ZN(n605) );
  XNOR2_X1 U677 ( .A(n605), .B(KEYINPUT55), .ZN(n606) );
  XNOR2_X1 U678 ( .A(n604), .B(n606), .ZN(n607) );
  XNOR2_X1 U679 ( .A(n608), .B(n607), .ZN(n610) );
  INV_X1 U680 ( .A(G952), .ZN(n609) );
  NOR2_X1 U681 ( .A1(n610), .A2(n725), .ZN(n612) );
  XOR2_X1 U682 ( .A(KEYINPUT119), .B(KEYINPUT56), .Z(n611) );
  XNOR2_X1 U683 ( .A(n612), .B(n611), .ZN(G51) );
  NAND2_X1 U684 ( .A1(n715), .A2(G472), .ZN(n615) );
  XOR2_X1 U685 ( .A(KEYINPUT62), .B(n613), .Z(n614) );
  XNOR2_X1 U686 ( .A(n615), .B(n614), .ZN(n616) );
  NOR2_X1 U687 ( .A1(n616), .A2(n725), .ZN(n619) );
  XNOR2_X1 U688 ( .A(KEYINPUT112), .B(KEYINPUT63), .ZN(n617) );
  XOR2_X1 U689 ( .A(n617), .B(KEYINPUT90), .Z(n618) );
  XNOR2_X1 U690 ( .A(n619), .B(n618), .ZN(G57) );
  NAND2_X1 U691 ( .A1(n715), .A2(G475), .ZN(n622) );
  XOR2_X1 U692 ( .A(KEYINPUT59), .B(n620), .Z(n621) );
  XNOR2_X1 U693 ( .A(n622), .B(n621), .ZN(n623) );
  NOR2_X1 U694 ( .A1(n623), .A2(n725), .ZN(n624) );
  XNOR2_X1 U695 ( .A(n624), .B(KEYINPUT60), .ZN(G60) );
  NAND2_X1 U696 ( .A1(G953), .A2(G224), .ZN(n625) );
  XNOR2_X1 U697 ( .A(KEYINPUT61), .B(n625), .ZN(n626) );
  NAND2_X1 U698 ( .A1(n626), .A2(G898), .ZN(n627) );
  XNOR2_X1 U699 ( .A(KEYINPUT123), .B(n627), .ZN(n631) );
  NOR2_X1 U700 ( .A1(n666), .A2(G953), .ZN(n629) );
  XNOR2_X1 U701 ( .A(n629), .B(KEYINPUT124), .ZN(n630) );
  NOR2_X1 U702 ( .A1(n631), .A2(n630), .ZN(n632) );
  XOR2_X1 U703 ( .A(KEYINPUT125), .B(n632), .Z(n636) );
  NOR2_X1 U704 ( .A1(n634), .A2(n633), .ZN(n635) );
  XOR2_X1 U705 ( .A(n636), .B(n635), .Z(G69) );
  XNOR2_X1 U706 ( .A(G101), .B(n637), .ZN(G3) );
  NAND2_X1 U707 ( .A1(n639), .A2(n651), .ZN(n638) );
  XNOR2_X1 U708 ( .A(n638), .B(G104), .ZN(G6) );
  XOR2_X1 U709 ( .A(KEYINPUT27), .B(KEYINPUT26), .Z(n641) );
  NAND2_X1 U710 ( .A1(n639), .A2(n654), .ZN(n640) );
  XNOR2_X1 U711 ( .A(n641), .B(n640), .ZN(n642) );
  XNOR2_X1 U712 ( .A(G107), .B(n642), .ZN(G9) );
  INV_X1 U713 ( .A(n643), .ZN(n644) );
  XOR2_X1 U714 ( .A(G110), .B(n644), .Z(G12) );
  NOR2_X1 U715 ( .A1(n649), .A2(n645), .ZN(n647) );
  XNOR2_X1 U716 ( .A(G128), .B(KEYINPUT29), .ZN(n646) );
  XNOR2_X1 U717 ( .A(n647), .B(n646), .ZN(G30) );
  NOR2_X1 U718 ( .A1(n649), .A2(n648), .ZN(n650) );
  XOR2_X1 U719 ( .A(G146), .B(n650), .Z(G48) );
  NAND2_X1 U720 ( .A1(n653), .A2(n651), .ZN(n652) );
  XNOR2_X1 U721 ( .A(n652), .B(G113), .ZN(G15) );
  NAND2_X1 U722 ( .A1(n654), .A2(n653), .ZN(n655) );
  XNOR2_X1 U723 ( .A(n655), .B(G116), .ZN(G18) );
  XNOR2_X1 U724 ( .A(KEYINPUT113), .B(KEYINPUT37), .ZN(n657) );
  XNOR2_X1 U725 ( .A(n657), .B(n656), .ZN(n658) );
  XNOR2_X1 U726 ( .A(G125), .B(n658), .ZN(G27) );
  XOR2_X1 U727 ( .A(KEYINPUT118), .B(KEYINPUT53), .Z(n708) );
  NOR2_X1 U728 ( .A1(n659), .A2(KEYINPUT85), .ZN(n663) );
  NAND2_X1 U729 ( .A1(n660), .A2(n729), .ZN(n661) );
  INV_X1 U730 ( .A(KEYINPUT2), .ZN(n664) );
  NAND2_X1 U731 ( .A1(n661), .A2(n664), .ZN(n662) );
  NAND2_X1 U732 ( .A1(n663), .A2(n662), .ZN(n669) );
  NAND2_X1 U733 ( .A1(KEYINPUT85), .A2(n664), .ZN(n665) );
  NOR2_X1 U734 ( .A1(n590), .A2(n665), .ZN(n667) );
  NAND2_X1 U735 ( .A1(n667), .A2(n666), .ZN(n668) );
  NAND2_X1 U736 ( .A1(n669), .A2(n668), .ZN(n702) );
  NAND2_X1 U737 ( .A1(n671), .A2(n670), .ZN(n672) );
  XOR2_X1 U738 ( .A(KEYINPUT115), .B(n672), .Z(n673) );
  XNOR2_X1 U739 ( .A(n673), .B(KEYINPUT50), .ZN(n679) );
  NOR2_X1 U740 ( .A1(n675), .A2(n674), .ZN(n676) );
  XOR2_X1 U741 ( .A(KEYINPUT49), .B(n676), .Z(n677) );
  NOR2_X1 U742 ( .A1(n347), .A2(n677), .ZN(n678) );
  NAND2_X1 U743 ( .A1(n679), .A2(n678), .ZN(n681) );
  NAND2_X1 U744 ( .A1(n681), .A2(n680), .ZN(n682) );
  XNOR2_X1 U745 ( .A(KEYINPUT51), .B(n682), .ZN(n683) );
  NOR2_X1 U746 ( .A1(n703), .A2(n683), .ZN(n696) );
  NOR2_X1 U747 ( .A1(n686), .A2(n685), .ZN(n687) );
  XNOR2_X1 U748 ( .A(KEYINPUT116), .B(n687), .ZN(n693) );
  NOR2_X1 U749 ( .A1(n689), .A2(n688), .ZN(n690) );
  NOR2_X1 U750 ( .A1(n691), .A2(n690), .ZN(n692) );
  NOR2_X1 U751 ( .A1(n693), .A2(n692), .ZN(n694) );
  NOR2_X1 U752 ( .A1(n684), .A2(n694), .ZN(n695) );
  NOR2_X1 U753 ( .A1(n696), .A2(n695), .ZN(n697) );
  XOR2_X1 U754 ( .A(KEYINPUT52), .B(n697), .Z(n699) );
  NAND2_X1 U755 ( .A1(n699), .A2(n698), .ZN(n700) );
  XNOR2_X1 U756 ( .A(KEYINPUT117), .B(n700), .ZN(n701) );
  NOR2_X1 U757 ( .A1(n702), .A2(n701), .ZN(n706) );
  NOR2_X1 U758 ( .A1(n703), .A2(n684), .ZN(n704) );
  NOR2_X1 U759 ( .A1(G953), .A2(n704), .ZN(n705) );
  NAND2_X1 U760 ( .A1(n706), .A2(n705), .ZN(n707) );
  XNOR2_X1 U761 ( .A(n708), .B(n707), .ZN(G75) );
  XNOR2_X1 U762 ( .A(KEYINPUT58), .B(KEYINPUT120), .ZN(n711) );
  XNOR2_X1 U763 ( .A(n709), .B(KEYINPUT57), .ZN(n710) );
  XNOR2_X1 U764 ( .A(n711), .B(n710), .ZN(n713) );
  NAND2_X1 U765 ( .A1(n715), .A2(G469), .ZN(n712) );
  XOR2_X1 U766 ( .A(n713), .B(n712), .Z(n714) );
  NOR2_X1 U767 ( .A1(n725), .A2(n714), .ZN(G54) );
  NAND2_X1 U768 ( .A1(n720), .A2(G478), .ZN(n718) );
  XOR2_X1 U769 ( .A(n716), .B(KEYINPUT121), .Z(n717) );
  XNOR2_X1 U770 ( .A(n718), .B(n717), .ZN(n719) );
  NOR2_X1 U771 ( .A1(n725), .A2(n719), .ZN(G63) );
  NAND2_X1 U772 ( .A1(n720), .A2(G217), .ZN(n723) );
  XNOR2_X1 U773 ( .A(n721), .B(KEYINPUT122), .ZN(n722) );
  XNOR2_X1 U774 ( .A(n723), .B(n722), .ZN(n724) );
  NOR2_X1 U775 ( .A1(n725), .A2(n724), .ZN(G66) );
  XNOR2_X1 U776 ( .A(n727), .B(n726), .ZN(n728) );
  XOR2_X1 U777 ( .A(n728), .B(KEYINPUT126), .Z(n732) );
  XOR2_X1 U778 ( .A(n732), .B(n729), .Z(n731) );
  NAND2_X1 U779 ( .A1(n731), .A2(n730), .ZN(n736) );
  XNOR2_X1 U780 ( .A(G227), .B(n732), .ZN(n733) );
  NAND2_X1 U781 ( .A1(n733), .A2(G900), .ZN(n734) );
  NAND2_X1 U782 ( .A1(G953), .A2(n734), .ZN(n735) );
  NAND2_X1 U783 ( .A1(n736), .A2(n735), .ZN(G72) );
  XOR2_X1 U784 ( .A(n737), .B(G122), .Z(G24) );
  XOR2_X1 U785 ( .A(G131), .B(n738), .Z(G33) );
  XNOR2_X1 U786 ( .A(G134), .B(KEYINPUT114), .ZN(n740) );
  XNOR2_X1 U787 ( .A(n740), .B(n739), .ZN(G36) );
  XOR2_X1 U788 ( .A(G137), .B(n741), .Z(G39) );
endmodule

