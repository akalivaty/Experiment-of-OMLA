//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 0 0 1 0 0 1 0 0 0 0 1 1 1 1 1 1 0 1 0 0 0 1 0 0 0 0 1 0 1 1 0 0 1 1 1 1 0 1 0 0 0 0 0 1 0 1 0 0 1 1 0 1 0 1 1 0 0 1 0 0 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:34:49 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n442, new_n446, new_n448, new_n452, new_n453, new_n454, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n526,
    new_n527, new_n528, new_n529, new_n530, new_n531, new_n532, new_n533,
    new_n534, new_n535, new_n536, new_n537, new_n538, new_n539, new_n540,
    new_n541, new_n542, new_n543, new_n544, new_n545, new_n546, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n558, new_n559, new_n560, new_n561, new_n562, new_n563,
    new_n564, new_n565, new_n566, new_n567, new_n568, new_n569, new_n570,
    new_n572, new_n574, new_n575, new_n577, new_n578, new_n579, new_n580,
    new_n581, new_n582, new_n583, new_n584, new_n585, new_n586, new_n587,
    new_n588, new_n589, new_n590, new_n591, new_n592, new_n593, new_n594,
    new_n596, new_n597, new_n598, new_n599, new_n600, new_n601, new_n602,
    new_n604, new_n605, new_n606, new_n607, new_n609, new_n610, new_n611,
    new_n612, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n621, new_n622, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n640, new_n641, new_n644, new_n645, new_n647,
    new_n648, new_n649, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n677, new_n678,
    new_n679, new_n680, new_n681, new_n682, new_n683, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n692, new_n693,
    new_n694, new_n695, new_n696, new_n697, new_n698, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n713, new_n714, new_n715,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1200;
  BUF_X1    g000(.A(G452), .Z(G350));
  XNOR2_X1  g001(.A(KEYINPUT64), .B(G452), .ZN(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  XNOR2_X1  g004(.A(KEYINPUT65), .B(G1083), .ZN(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  XNOR2_X1  g014(.A(KEYINPUT66), .B(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  AND2_X1   g016(.A1(G2072), .A2(G2078), .ZN(new_n442));
  NAND3_X1  g017(.A1(new_n442), .A2(G2084), .A3(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  NAND2_X1  g020(.A1(G94), .A2(G452), .ZN(new_n446));
  XNOR2_X1  g021(.A(new_n446), .B(KEYINPUT67), .ZN(G173));
  NAND2_X1  g022(.A1(G7), .A2(G661), .ZN(new_n448));
  XOR2_X1   g023(.A(new_n448), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g024(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g025(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g026(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n452));
  XNOR2_X1  g027(.A(new_n452), .B(KEYINPUT2), .ZN(new_n453));
  NOR4_X1   g028(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n454));
  NAND2_X1  g029(.A1(new_n453), .A2(new_n454), .ZN(G261));
  INV_X1    g030(.A(G261), .ZN(G325));
  INV_X1    g031(.A(new_n453), .ZN(new_n457));
  NAND2_X1  g032(.A1(new_n457), .A2(G2106), .ZN(new_n458));
  INV_X1    g033(.A(G567), .ZN(new_n459));
  OR2_X1    g034(.A1(new_n454), .A2(new_n459), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n458), .A2(new_n460), .ZN(new_n461));
  INV_X1    g036(.A(new_n461), .ZN(G319));
  INV_X1    g037(.A(G2105), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n463), .A2(G2104), .ZN(new_n464));
  XNOR2_X1  g039(.A(new_n464), .B(KEYINPUT69), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n465), .A2(G101), .ZN(new_n466));
  AOI21_X1  g041(.A(KEYINPUT3), .B1(KEYINPUT68), .B2(G2104), .ZN(new_n467));
  INV_X1    g042(.A(new_n467), .ZN(new_n468));
  NAND3_X1  g043(.A1(KEYINPUT68), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n469));
  AOI21_X1  g044(.A(G2105), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n470), .A2(G137), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n466), .A2(new_n471), .ZN(new_n472));
  XNOR2_X1  g047(.A(KEYINPUT3), .B(G2104), .ZN(new_n473));
  AOI22_X1  g048(.A1(new_n473), .A2(G125), .B1(G113), .B2(G2104), .ZN(new_n474));
  NOR2_X1   g049(.A1(new_n474), .A2(new_n463), .ZN(new_n475));
  NOR2_X1   g050(.A1(new_n472), .A2(new_n475), .ZN(G160));
  NAND2_X1  g051(.A1(new_n468), .A2(new_n469), .ZN(new_n477));
  OR2_X1    g052(.A1(new_n477), .A2(KEYINPUT70), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n477), .A2(KEYINPUT70), .ZN(new_n479));
  NAND3_X1  g054(.A1(new_n478), .A2(new_n463), .A3(new_n479), .ZN(new_n480));
  INV_X1    g055(.A(new_n480), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n481), .A2(G136), .ZN(new_n482));
  AND3_X1   g057(.A1(new_n478), .A2(G2105), .A3(new_n479), .ZN(new_n483));
  NAND2_X1  g058(.A1(new_n483), .A2(G124), .ZN(new_n484));
  OR2_X1    g059(.A1(G100), .A2(G2105), .ZN(new_n485));
  OAI211_X1 g060(.A(new_n485), .B(G2104), .C1(G112), .C2(new_n463), .ZN(new_n486));
  NAND3_X1  g061(.A1(new_n482), .A2(new_n484), .A3(new_n486), .ZN(new_n487));
  INV_X1    g062(.A(new_n487), .ZN(G162));
  NAND3_X1  g063(.A1(new_n473), .A2(G138), .A3(new_n463), .ZN(new_n489));
  INV_X1    g064(.A(KEYINPUT4), .ZN(new_n490));
  NAND2_X1  g065(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  AND2_X1   g066(.A1(KEYINPUT4), .A2(G138), .ZN(new_n492));
  NAND2_X1  g067(.A1(new_n470), .A2(new_n492), .ZN(new_n493));
  NAND2_X1  g068(.A1(new_n491), .A2(new_n493), .ZN(new_n494));
  AND2_X1   g069(.A1(G126), .A2(G2105), .ZN(new_n495));
  INV_X1    g070(.A(new_n469), .ZN(new_n496));
  OAI21_X1  g071(.A(new_n495), .B1(new_n496), .B2(new_n467), .ZN(new_n497));
  INV_X1    g072(.A(G114), .ZN(new_n498));
  NAND2_X1  g073(.A1(new_n498), .A2(KEYINPUT71), .ZN(new_n499));
  INV_X1    g074(.A(KEYINPUT71), .ZN(new_n500));
  NAND2_X1  g075(.A1(new_n500), .A2(G114), .ZN(new_n501));
  AOI21_X1  g076(.A(new_n463), .B1(new_n499), .B2(new_n501), .ZN(new_n502));
  OAI21_X1  g077(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n503));
  OAI21_X1  g078(.A(new_n497), .B1(new_n502), .B2(new_n503), .ZN(new_n504));
  NOR2_X1   g079(.A1(new_n494), .A2(new_n504), .ZN(G164));
  INV_X1    g080(.A(G543), .ZN(new_n506));
  NOR2_X1   g081(.A1(new_n506), .A2(KEYINPUT5), .ZN(new_n507));
  INV_X1    g082(.A(KEYINPUT72), .ZN(new_n508));
  INV_X1    g083(.A(KEYINPUT5), .ZN(new_n509));
  OAI21_X1  g084(.A(new_n508), .B1(new_n509), .B2(G543), .ZN(new_n510));
  NAND3_X1  g085(.A1(new_n506), .A2(KEYINPUT72), .A3(KEYINPUT5), .ZN(new_n511));
  AOI21_X1  g086(.A(new_n507), .B1(new_n510), .B2(new_n511), .ZN(new_n512));
  AOI22_X1  g087(.A1(new_n512), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n513));
  INV_X1    g088(.A(G651), .ZN(new_n514));
  NOR2_X1   g089(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  OR2_X1    g090(.A1(KEYINPUT6), .A2(G651), .ZN(new_n516));
  NAND2_X1  g091(.A1(KEYINPUT6), .A2(G651), .ZN(new_n517));
  AOI21_X1  g092(.A(new_n506), .B1(new_n516), .B2(new_n517), .ZN(new_n518));
  NAND2_X1  g093(.A1(new_n518), .A2(G50), .ZN(new_n519));
  XNOR2_X1  g094(.A(KEYINPUT6), .B(G651), .ZN(new_n520));
  NAND2_X1  g095(.A1(new_n512), .A2(new_n520), .ZN(new_n521));
  INV_X1    g096(.A(G88), .ZN(new_n522));
  OAI21_X1  g097(.A(new_n519), .B1(new_n521), .B2(new_n522), .ZN(new_n523));
  OR2_X1    g098(.A1(new_n515), .A2(new_n523), .ZN(G303));
  INV_X1    g099(.A(G303), .ZN(G166));
  NAND2_X1  g100(.A1(new_n509), .A2(G543), .ZN(new_n526));
  AND2_X1   g101(.A1(G63), .A2(G651), .ZN(new_n527));
  AND3_X1   g102(.A1(new_n506), .A2(KEYINPUT72), .A3(KEYINPUT5), .ZN(new_n528));
  AOI21_X1  g103(.A(KEYINPUT72), .B1(new_n506), .B2(KEYINPUT5), .ZN(new_n529));
  OAI211_X1 g104(.A(new_n526), .B(new_n527), .C1(new_n528), .C2(new_n529), .ZN(new_n530));
  NAND3_X1  g105(.A1(new_n520), .A2(G51), .A3(G543), .ZN(new_n531));
  NAND3_X1  g106(.A1(new_n530), .A2(KEYINPUT73), .A3(new_n531), .ZN(new_n532));
  INV_X1    g107(.A(new_n532), .ZN(new_n533));
  AOI21_X1  g108(.A(KEYINPUT73), .B1(new_n530), .B2(new_n531), .ZN(new_n534));
  NAND2_X1  g109(.A1(new_n510), .A2(new_n511), .ZN(new_n535));
  NAND4_X1  g110(.A1(new_n535), .A2(G89), .A3(new_n526), .A4(new_n520), .ZN(new_n536));
  NAND3_X1  g111(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n537));
  INV_X1    g112(.A(new_n537), .ZN(new_n538));
  NAND2_X1  g113(.A1(KEYINPUT74), .A2(KEYINPUT7), .ZN(new_n539));
  INV_X1    g114(.A(new_n539), .ZN(new_n540));
  NOR2_X1   g115(.A1(KEYINPUT74), .A2(KEYINPUT7), .ZN(new_n541));
  OAI21_X1  g116(.A(new_n538), .B1(new_n540), .B2(new_n541), .ZN(new_n542));
  INV_X1    g117(.A(new_n541), .ZN(new_n543));
  NAND3_X1  g118(.A1(new_n543), .A2(new_n537), .A3(new_n539), .ZN(new_n544));
  NAND2_X1  g119(.A1(new_n542), .A2(new_n544), .ZN(new_n545));
  NAND2_X1  g120(.A1(new_n536), .A2(new_n545), .ZN(new_n546));
  NOR3_X1   g121(.A1(new_n533), .A2(new_n534), .A3(new_n546), .ZN(G168));
  NAND3_X1  g122(.A1(new_n535), .A2(G64), .A3(new_n526), .ZN(new_n548));
  NAND2_X1  g123(.A1(G77), .A2(G543), .ZN(new_n549));
  AOI21_X1  g124(.A(new_n514), .B1(new_n548), .B2(new_n549), .ZN(new_n550));
  AND2_X1   g125(.A1(KEYINPUT75), .A2(G90), .ZN(new_n551));
  NOR2_X1   g126(.A1(KEYINPUT75), .A2(G90), .ZN(new_n552));
  NOR2_X1   g127(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  NAND4_X1  g128(.A1(new_n535), .A2(new_n526), .A3(new_n520), .A4(new_n553), .ZN(new_n554));
  NAND2_X1  g129(.A1(new_n518), .A2(G52), .ZN(new_n555));
  NAND2_X1  g130(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  NOR2_X1   g131(.A1(new_n550), .A2(new_n556), .ZN(G171));
  AND2_X1   g132(.A1(new_n512), .A2(new_n520), .ZN(new_n558));
  AOI22_X1  g133(.A1(new_n558), .A2(G81), .B1(G43), .B2(new_n518), .ZN(new_n559));
  NAND2_X1  g134(.A1(G68), .A2(G543), .ZN(new_n560));
  INV_X1    g135(.A(new_n560), .ZN(new_n561));
  AOI21_X1  g136(.A(new_n561), .B1(new_n512), .B2(G56), .ZN(new_n562));
  OAI21_X1  g137(.A(G651), .B1(new_n562), .B2(KEYINPUT76), .ZN(new_n563));
  OAI211_X1 g138(.A(G56), .B(new_n526), .C1(new_n528), .C2(new_n529), .ZN(new_n564));
  NAND2_X1  g139(.A1(new_n564), .A2(new_n560), .ZN(new_n565));
  INV_X1    g140(.A(KEYINPUT76), .ZN(new_n566));
  NOR2_X1   g141(.A1(new_n565), .A2(new_n566), .ZN(new_n567));
  OAI21_X1  g142(.A(new_n559), .B1(new_n563), .B2(new_n567), .ZN(new_n568));
  INV_X1    g143(.A(new_n568), .ZN(new_n569));
  NAND2_X1  g144(.A1(new_n569), .A2(G860), .ZN(new_n570));
  XNOR2_X1  g145(.A(new_n570), .B(KEYINPUT77), .ZN(G153));
  AND3_X1   g146(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n572));
  NAND2_X1  g147(.A1(new_n572), .A2(G36), .ZN(G176));
  NAND2_X1  g148(.A1(G1), .A2(G3), .ZN(new_n574));
  XNOR2_X1  g149(.A(new_n574), .B(KEYINPUT8), .ZN(new_n575));
  NAND2_X1  g150(.A1(new_n572), .A2(new_n575), .ZN(G188));
  INV_X1    g151(.A(new_n517), .ZN(new_n577));
  NOR2_X1   g152(.A1(KEYINPUT6), .A2(G651), .ZN(new_n578));
  OAI211_X1 g153(.A(G53), .B(G543), .C1(new_n577), .C2(new_n578), .ZN(new_n579));
  NAND2_X1  g154(.A1(new_n579), .A2(KEYINPUT9), .ZN(new_n580));
  INV_X1    g155(.A(KEYINPUT9), .ZN(new_n581));
  NAND3_X1  g156(.A1(new_n518), .A2(new_n581), .A3(G53), .ZN(new_n582));
  AOI22_X1  g157(.A1(new_n558), .A2(G91), .B1(new_n580), .B2(new_n582), .ZN(new_n583));
  NAND2_X1  g158(.A1(new_n512), .A2(G65), .ZN(new_n584));
  NAND2_X1  g159(.A1(G78), .A2(G543), .ZN(new_n585));
  NAND2_X1  g160(.A1(new_n584), .A2(new_n585), .ZN(new_n586));
  NAND2_X1  g161(.A1(new_n586), .A2(G651), .ZN(new_n587));
  AOI21_X1  g162(.A(KEYINPUT78), .B1(new_n583), .B2(new_n587), .ZN(new_n588));
  NAND2_X1  g163(.A1(new_n582), .A2(new_n580), .ZN(new_n589));
  NAND3_X1  g164(.A1(new_n512), .A2(G91), .A3(new_n520), .ZN(new_n590));
  NAND2_X1  g165(.A1(new_n589), .A2(new_n590), .ZN(new_n591));
  AOI21_X1  g166(.A(new_n514), .B1(new_n584), .B2(new_n585), .ZN(new_n592));
  INV_X1    g167(.A(KEYINPUT78), .ZN(new_n593));
  NOR3_X1   g168(.A1(new_n591), .A2(new_n592), .A3(new_n593), .ZN(new_n594));
  NOR2_X1   g169(.A1(new_n588), .A2(new_n594), .ZN(G299));
  NAND2_X1  g170(.A1(new_n548), .A2(new_n549), .ZN(new_n596));
  NAND2_X1  g171(.A1(new_n596), .A2(G651), .ZN(new_n597));
  AND2_X1   g172(.A1(new_n554), .A2(new_n555), .ZN(new_n598));
  NAND3_X1  g173(.A1(new_n597), .A2(new_n598), .A3(KEYINPUT79), .ZN(new_n599));
  INV_X1    g174(.A(KEYINPUT79), .ZN(new_n600));
  OAI21_X1  g175(.A(new_n600), .B1(new_n550), .B2(new_n556), .ZN(new_n601));
  NAND2_X1  g176(.A1(new_n599), .A2(new_n601), .ZN(new_n602));
  INV_X1    g177(.A(new_n602), .ZN(G301));
  NAND2_X1  g178(.A1(new_n530), .A2(new_n531), .ZN(new_n604));
  INV_X1    g179(.A(KEYINPUT73), .ZN(new_n605));
  NAND2_X1  g180(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  AND2_X1   g181(.A1(new_n536), .A2(new_n545), .ZN(new_n607));
  NAND3_X1  g182(.A1(new_n606), .A2(new_n607), .A3(new_n532), .ZN(G286));
  NAND2_X1  g183(.A1(new_n518), .A2(G49), .ZN(new_n609));
  XNOR2_X1  g184(.A(new_n609), .B(KEYINPUT80), .ZN(new_n610));
  NAND2_X1  g185(.A1(new_n558), .A2(G87), .ZN(new_n611));
  OAI21_X1  g186(.A(G651), .B1(new_n512), .B2(G74), .ZN(new_n612));
  NAND3_X1  g187(.A1(new_n610), .A2(new_n611), .A3(new_n612), .ZN(G288));
  AOI22_X1  g188(.A1(new_n512), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n614));
  NOR2_X1   g189(.A1(new_n614), .A2(new_n514), .ZN(new_n615));
  NAND2_X1  g190(.A1(new_n518), .A2(G48), .ZN(new_n616));
  INV_X1    g191(.A(G86), .ZN(new_n617));
  OAI21_X1  g192(.A(new_n616), .B1(new_n521), .B2(new_n617), .ZN(new_n618));
  NOR2_X1   g193(.A1(new_n615), .A2(new_n618), .ZN(new_n619));
  INV_X1    g194(.A(new_n619), .ZN(G305));
  AOI22_X1  g195(.A1(new_n558), .A2(G85), .B1(G47), .B2(new_n518), .ZN(new_n621));
  AOI22_X1  g196(.A1(new_n512), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n622));
  OAI21_X1  g197(.A(new_n621), .B1(new_n514), .B2(new_n622), .ZN(G290));
  NAND2_X1  g198(.A1(new_n512), .A2(G66), .ZN(new_n624));
  INV_X1    g199(.A(G79), .ZN(new_n625));
  OAI21_X1  g200(.A(new_n624), .B1(new_n625), .B2(new_n506), .ZN(new_n626));
  INV_X1    g201(.A(new_n518), .ZN(new_n627));
  OR2_X1    g202(.A1(new_n627), .A2(KEYINPUT81), .ZN(new_n628));
  INV_X1    g203(.A(G54), .ZN(new_n629));
  AOI21_X1  g204(.A(new_n629), .B1(new_n627), .B2(KEYINPUT81), .ZN(new_n630));
  AOI22_X1  g205(.A1(new_n626), .A2(G651), .B1(new_n628), .B2(new_n630), .ZN(new_n631));
  NAND3_X1  g206(.A1(new_n558), .A2(KEYINPUT10), .A3(G92), .ZN(new_n632));
  INV_X1    g207(.A(KEYINPUT10), .ZN(new_n633));
  INV_X1    g208(.A(G92), .ZN(new_n634));
  OAI21_X1  g209(.A(new_n633), .B1(new_n521), .B2(new_n634), .ZN(new_n635));
  NAND2_X1  g210(.A1(new_n632), .A2(new_n635), .ZN(new_n636));
  NAND2_X1  g211(.A1(new_n631), .A2(new_n636), .ZN(new_n637));
  MUX2_X1   g212(.A(new_n637), .B(G301), .S(G868), .Z(G284));
  MUX2_X1   g213(.A(new_n637), .B(G301), .S(G868), .Z(G321));
  INV_X1    g214(.A(G868), .ZN(new_n640));
  NAND2_X1  g215(.A1(G299), .A2(new_n640), .ZN(new_n641));
  OAI21_X1  g216(.A(new_n641), .B1(new_n640), .B2(G168), .ZN(G297));
  OAI21_X1  g217(.A(new_n641), .B1(new_n640), .B2(G168), .ZN(G280));
  INV_X1    g218(.A(new_n637), .ZN(new_n644));
  INV_X1    g219(.A(G559), .ZN(new_n645));
  OAI21_X1  g220(.A(new_n644), .B1(new_n645), .B2(G860), .ZN(G148));
  NAND2_X1  g221(.A1(new_n568), .A2(new_n640), .ZN(new_n647));
  NOR2_X1   g222(.A1(new_n637), .A2(G559), .ZN(new_n648));
  OAI21_X1  g223(.A(new_n647), .B1(new_n648), .B2(new_n640), .ZN(new_n649));
  XOR2_X1   g224(.A(new_n649), .B(KEYINPUT82), .Z(G323));
  XNOR2_X1  g225(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g226(.A1(new_n481), .A2(G135), .ZN(new_n652));
  XOR2_X1   g227(.A(new_n652), .B(KEYINPUT84), .Z(new_n653));
  NAND2_X1  g228(.A1(new_n483), .A2(G123), .ZN(new_n654));
  XOR2_X1   g229(.A(new_n654), .B(KEYINPUT85), .Z(new_n655));
  OR2_X1    g230(.A1(G99), .A2(G2105), .ZN(new_n656));
  OAI211_X1 g231(.A(new_n656), .B(G2104), .C1(G111), .C2(new_n463), .ZN(new_n657));
  NAND3_X1  g232(.A1(new_n653), .A2(new_n655), .A3(new_n657), .ZN(new_n658));
  OR2_X1    g233(.A1(new_n658), .A2(G2096), .ZN(new_n659));
  NAND2_X1  g234(.A1(new_n658), .A2(G2096), .ZN(new_n660));
  NAND2_X1  g235(.A1(new_n465), .A2(new_n473), .ZN(new_n661));
  XOR2_X1   g236(.A(new_n661), .B(KEYINPUT12), .Z(new_n662));
  XNOR2_X1  g237(.A(new_n662), .B(KEYINPUT13), .ZN(new_n663));
  OAI21_X1  g238(.A(new_n663), .B1(KEYINPUT83), .B2(G2100), .ZN(new_n664));
  NAND2_X1  g239(.A1(KEYINPUT83), .A2(G2100), .ZN(new_n665));
  NAND2_X1  g240(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  NAND3_X1  g241(.A1(new_n663), .A2(KEYINPUT83), .A3(G2100), .ZN(new_n667));
  NAND4_X1  g242(.A1(new_n659), .A2(new_n660), .A3(new_n666), .A4(new_n667), .ZN(G156));
  XNOR2_X1  g243(.A(G2427), .B(G2438), .ZN(new_n669));
  XNOR2_X1  g244(.A(new_n669), .B(G2430), .ZN(new_n670));
  XNOR2_X1  g245(.A(KEYINPUT15), .B(G2435), .ZN(new_n671));
  OR2_X1    g246(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  NAND2_X1  g247(.A1(new_n670), .A2(new_n671), .ZN(new_n673));
  NAND3_X1  g248(.A1(new_n672), .A2(KEYINPUT14), .A3(new_n673), .ZN(new_n674));
  XNOR2_X1  g249(.A(G2451), .B(G2454), .ZN(new_n675));
  XNOR2_X1  g250(.A(new_n675), .B(KEYINPUT16), .ZN(new_n676));
  XNOR2_X1  g251(.A(new_n674), .B(new_n676), .ZN(new_n677));
  XNOR2_X1  g252(.A(G2443), .B(G2446), .ZN(new_n678));
  XNOR2_X1  g253(.A(new_n677), .B(new_n678), .ZN(new_n679));
  XNOR2_X1  g254(.A(G1341), .B(G1348), .ZN(new_n680));
  NAND2_X1  g255(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  XNOR2_X1  g256(.A(new_n681), .B(KEYINPUT86), .ZN(new_n682));
  OAI21_X1  g257(.A(G14), .B1(new_n679), .B2(new_n680), .ZN(new_n683));
  NOR2_X1   g258(.A1(new_n682), .A2(new_n683), .ZN(G401));
  XNOR2_X1  g259(.A(G2067), .B(G2678), .ZN(new_n685));
  XOR2_X1   g260(.A(new_n685), .B(KEYINPUT87), .Z(new_n686));
  NOR2_X1   g261(.A1(G2072), .A2(G2078), .ZN(new_n687));
  NOR2_X1   g262(.A1(new_n442), .A2(new_n687), .ZN(new_n688));
  NAND2_X1  g263(.A1(new_n686), .A2(new_n688), .ZN(new_n689));
  XOR2_X1   g264(.A(G2084), .B(G2090), .Z(new_n690));
  INV_X1    g265(.A(new_n690), .ZN(new_n691));
  XNOR2_X1  g266(.A(new_n688), .B(KEYINPUT17), .ZN(new_n692));
  OAI211_X1 g267(.A(new_n689), .B(new_n691), .C1(new_n686), .C2(new_n692), .ZN(new_n693));
  OAI211_X1 g268(.A(new_n690), .B(new_n685), .C1(new_n442), .C2(new_n687), .ZN(new_n694));
  XOR2_X1   g269(.A(new_n694), .B(KEYINPUT18), .Z(new_n695));
  NAND3_X1  g270(.A1(new_n686), .A2(new_n692), .A3(new_n690), .ZN(new_n696));
  NAND3_X1  g271(.A1(new_n693), .A2(new_n695), .A3(new_n696), .ZN(new_n697));
  XOR2_X1   g272(.A(G2096), .B(G2100), .Z(new_n698));
  XNOR2_X1  g273(.A(new_n697), .B(new_n698), .ZN(G227));
  XOR2_X1   g274(.A(G1971), .B(G1976), .Z(new_n700));
  XNOR2_X1  g275(.A(new_n700), .B(KEYINPUT19), .ZN(new_n701));
  XOR2_X1   g276(.A(G1956), .B(G2474), .Z(new_n702));
  XOR2_X1   g277(.A(G1961), .B(G1966), .Z(new_n703));
  AND2_X1   g278(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  NAND2_X1  g279(.A1(new_n701), .A2(new_n704), .ZN(new_n705));
  XNOR2_X1  g280(.A(new_n705), .B(KEYINPUT20), .ZN(new_n706));
  NOR2_X1   g281(.A1(new_n702), .A2(new_n703), .ZN(new_n707));
  NOR3_X1   g282(.A1(new_n701), .A2(new_n704), .A3(new_n707), .ZN(new_n708));
  AOI21_X1  g283(.A(new_n708), .B1(new_n701), .B2(new_n707), .ZN(new_n709));
  AND2_X1   g284(.A1(new_n706), .A2(new_n709), .ZN(new_n710));
  XOR2_X1   g285(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n711));
  XNOR2_X1  g286(.A(new_n710), .B(new_n711), .ZN(new_n712));
  XNOR2_X1  g287(.A(G1991), .B(G1996), .ZN(new_n713));
  XNOR2_X1  g288(.A(new_n712), .B(new_n713), .ZN(new_n714));
  XNOR2_X1  g289(.A(G1981), .B(G1986), .ZN(new_n715));
  XNOR2_X1  g290(.A(new_n714), .B(new_n715), .ZN(G229));
  INV_X1    g291(.A(G29), .ZN(new_n717));
  NAND2_X1  g292(.A1(new_n717), .A2(G35), .ZN(new_n718));
  OAI21_X1  g293(.A(new_n718), .B1(G162), .B2(new_n717), .ZN(new_n719));
  XOR2_X1   g294(.A(new_n719), .B(KEYINPUT29), .Z(new_n720));
  INV_X1    g295(.A(G2090), .ZN(new_n721));
  NOR2_X1   g296(.A1(new_n720), .A2(new_n721), .ZN(new_n722));
  XNOR2_X1  g297(.A(new_n722), .B(KEYINPUT99), .ZN(new_n723));
  INV_X1    g298(.A(G27), .ZN(new_n724));
  OR3_X1    g299(.A1(new_n724), .A2(KEYINPUT97), .A3(G29), .ZN(new_n725));
  OAI21_X1  g300(.A(KEYINPUT97), .B1(new_n724), .B2(G29), .ZN(new_n726));
  OAI211_X1 g301(.A(new_n725), .B(new_n726), .C1(G164), .C2(new_n717), .ZN(new_n727));
  XOR2_X1   g302(.A(KEYINPUT98), .B(G2078), .Z(new_n728));
  XNOR2_X1  g303(.A(new_n727), .B(new_n728), .ZN(new_n729));
  INV_X1    g304(.A(G34), .ZN(new_n730));
  AOI21_X1  g305(.A(G29), .B1(new_n730), .B2(KEYINPUT24), .ZN(new_n731));
  NAND2_X1  g306(.A1(new_n731), .A2(KEYINPUT93), .ZN(new_n732));
  OAI21_X1  g307(.A(new_n732), .B1(KEYINPUT24), .B2(new_n730), .ZN(new_n733));
  NOR2_X1   g308(.A1(new_n731), .A2(KEYINPUT93), .ZN(new_n734));
  NOR2_X1   g309(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  AOI21_X1  g310(.A(new_n735), .B1(G160), .B2(G29), .ZN(new_n736));
  NAND2_X1  g311(.A1(new_n736), .A2(G2084), .ZN(new_n737));
  XOR2_X1   g312(.A(KEYINPUT31), .B(G11), .Z(new_n738));
  XOR2_X1   g313(.A(KEYINPUT94), .B(G28), .Z(new_n739));
  AOI21_X1  g314(.A(G29), .B1(new_n739), .B2(KEYINPUT30), .ZN(new_n740));
  INV_X1    g315(.A(KEYINPUT95), .ZN(new_n741));
  OR2_X1    g316(.A1(new_n740), .A2(new_n741), .ZN(new_n742));
  NOR2_X1   g317(.A1(new_n739), .A2(KEYINPUT30), .ZN(new_n743));
  AOI21_X1  g318(.A(new_n743), .B1(new_n740), .B2(new_n741), .ZN(new_n744));
  AOI21_X1  g319(.A(new_n738), .B1(new_n742), .B2(new_n744), .ZN(new_n745));
  NAND3_X1  g320(.A1(new_n729), .A2(new_n737), .A3(new_n745), .ZN(new_n746));
  XOR2_X1   g321(.A(KEYINPUT92), .B(G1348), .Z(new_n747));
  NOR2_X1   g322(.A1(G4), .A2(G16), .ZN(new_n748));
  XNOR2_X1  g323(.A(new_n748), .B(KEYINPUT91), .ZN(new_n749));
  INV_X1    g324(.A(G16), .ZN(new_n750));
  OAI21_X1  g325(.A(new_n749), .B1(new_n637), .B2(new_n750), .ZN(new_n751));
  OAI22_X1  g326(.A1(new_n658), .A2(new_n717), .B1(new_n747), .B2(new_n751), .ZN(new_n752));
  AND2_X1   g327(.A1(new_n717), .A2(G32), .ZN(new_n753));
  NAND2_X1  g328(.A1(new_n481), .A2(G141), .ZN(new_n754));
  NAND2_X1  g329(.A1(new_n483), .A2(G129), .ZN(new_n755));
  NAND3_X1  g330(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n756));
  INV_X1    g331(.A(KEYINPUT26), .ZN(new_n757));
  NAND2_X1  g332(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  OR2_X1    g333(.A1(new_n756), .A2(new_n757), .ZN(new_n759));
  AOI22_X1  g334(.A1(new_n465), .A2(G105), .B1(new_n758), .B2(new_n759), .ZN(new_n760));
  NAND3_X1  g335(.A1(new_n754), .A2(new_n755), .A3(new_n760), .ZN(new_n761));
  AOI21_X1  g336(.A(new_n753), .B1(new_n761), .B2(G29), .ZN(new_n762));
  XNOR2_X1  g337(.A(KEYINPUT27), .B(G1996), .ZN(new_n763));
  AOI211_X1 g338(.A(new_n746), .B(new_n752), .C1(new_n762), .C2(new_n763), .ZN(new_n764));
  NAND2_X1  g339(.A1(new_n750), .A2(G21), .ZN(new_n765));
  OAI21_X1  g340(.A(new_n765), .B1(G168), .B2(new_n750), .ZN(new_n766));
  NOR2_X1   g341(.A1(new_n766), .A2(G1966), .ZN(new_n767));
  AND2_X1   g342(.A1(new_n766), .A2(G1966), .ZN(new_n768));
  AOI211_X1 g343(.A(new_n767), .B(new_n768), .C1(new_n747), .C2(new_n751), .ZN(new_n769));
  XNOR2_X1  g344(.A(KEYINPUT88), .B(G16), .ZN(new_n770));
  INV_X1    g345(.A(new_n770), .ZN(new_n771));
  NOR2_X1   g346(.A1(new_n771), .A2(G19), .ZN(new_n772));
  AOI21_X1  g347(.A(new_n772), .B1(new_n569), .B2(new_n771), .ZN(new_n773));
  XNOR2_X1  g348(.A(new_n773), .B(G1341), .ZN(new_n774));
  AOI21_X1  g349(.A(new_n774), .B1(new_n720), .B2(new_n721), .ZN(new_n775));
  NAND3_X1  g350(.A1(new_n764), .A2(new_n769), .A3(new_n775), .ZN(new_n776));
  NOR2_X1   g351(.A1(G171), .A2(new_n750), .ZN(new_n777));
  AOI21_X1  g352(.A(new_n777), .B1(G5), .B2(new_n750), .ZN(new_n778));
  INV_X1    g353(.A(G1961), .ZN(new_n779));
  NAND2_X1  g354(.A1(new_n778), .A2(new_n779), .ZN(new_n780));
  OAI221_X1 g355(.A(new_n780), .B1(G2084), .B2(new_n736), .C1(new_n762), .C2(new_n763), .ZN(new_n781));
  XNOR2_X1  g356(.A(new_n781), .B(KEYINPUT96), .ZN(new_n782));
  NAND3_X1  g357(.A1(new_n463), .A2(G103), .A3(G2104), .ZN(new_n783));
  XOR2_X1   g358(.A(new_n783), .B(KEYINPUT25), .Z(new_n784));
  AOI22_X1  g359(.A1(new_n473), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n785));
  INV_X1    g360(.A(G139), .ZN(new_n786));
  OAI221_X1 g361(.A(new_n784), .B1(new_n463), .B2(new_n785), .C1(new_n480), .C2(new_n786), .ZN(new_n787));
  MUX2_X1   g362(.A(G33), .B(new_n787), .S(G29), .Z(new_n788));
  NAND2_X1  g363(.A1(new_n788), .A2(G2072), .ZN(new_n789));
  OAI21_X1  g364(.A(new_n789), .B1(new_n779), .B2(new_n778), .ZN(new_n790));
  INV_X1    g365(.A(G1956), .ZN(new_n791));
  NAND2_X1  g366(.A1(G299), .A2(G16), .ZN(new_n792));
  NAND2_X1  g367(.A1(new_n770), .A2(G20), .ZN(new_n793));
  XNOR2_X1  g368(.A(new_n793), .B(KEYINPUT23), .ZN(new_n794));
  AOI21_X1  g369(.A(new_n791), .B1(new_n792), .B2(new_n794), .ZN(new_n795));
  NOR2_X1   g370(.A1(new_n788), .A2(G2072), .ZN(new_n796));
  NOR3_X1   g371(.A1(new_n790), .A2(new_n795), .A3(new_n796), .ZN(new_n797));
  NAND2_X1  g372(.A1(new_n717), .A2(G26), .ZN(new_n798));
  XNOR2_X1  g373(.A(new_n798), .B(KEYINPUT28), .ZN(new_n799));
  NAND2_X1  g374(.A1(new_n481), .A2(G140), .ZN(new_n800));
  NAND2_X1  g375(.A1(new_n483), .A2(G128), .ZN(new_n801));
  OR2_X1    g376(.A1(G104), .A2(G2105), .ZN(new_n802));
  OAI211_X1 g377(.A(new_n802), .B(G2104), .C1(G116), .C2(new_n463), .ZN(new_n803));
  NAND3_X1  g378(.A1(new_n800), .A2(new_n801), .A3(new_n803), .ZN(new_n804));
  INV_X1    g379(.A(new_n804), .ZN(new_n805));
  OAI21_X1  g380(.A(new_n799), .B1(new_n805), .B2(new_n717), .ZN(new_n806));
  INV_X1    g381(.A(G2067), .ZN(new_n807));
  XNOR2_X1  g382(.A(new_n806), .B(new_n807), .ZN(new_n808));
  NAND3_X1  g383(.A1(new_n792), .A2(new_n791), .A3(new_n794), .ZN(new_n809));
  NAND4_X1  g384(.A1(new_n782), .A2(new_n797), .A3(new_n808), .A4(new_n809), .ZN(new_n810));
  NOR3_X1   g385(.A1(new_n723), .A2(new_n776), .A3(new_n810), .ZN(new_n811));
  NAND2_X1  g386(.A1(new_n619), .A2(G16), .ZN(new_n812));
  OAI21_X1  g387(.A(new_n812), .B1(G6), .B2(G16), .ZN(new_n813));
  XOR2_X1   g388(.A(KEYINPUT32), .B(G1981), .Z(new_n814));
  AND2_X1   g389(.A1(new_n750), .A2(G23), .ZN(new_n815));
  AOI21_X1  g390(.A(new_n815), .B1(G288), .B2(G16), .ZN(new_n816));
  XNOR2_X1  g391(.A(KEYINPUT33), .B(G1976), .ZN(new_n817));
  AOI22_X1  g392(.A1(new_n813), .A2(new_n814), .B1(new_n816), .B2(new_n817), .ZN(new_n818));
  OR2_X1    g393(.A1(new_n816), .A2(new_n817), .ZN(new_n819));
  OAI211_X1 g394(.A(new_n818), .B(new_n819), .C1(new_n813), .C2(new_n814), .ZN(new_n820));
  NOR2_X1   g395(.A1(new_n771), .A2(G22), .ZN(new_n821));
  AOI21_X1  g396(.A(new_n821), .B1(G166), .B2(new_n771), .ZN(new_n822));
  XNOR2_X1  g397(.A(new_n822), .B(G1971), .ZN(new_n823));
  NOR2_X1   g398(.A1(new_n820), .A2(new_n823), .ZN(new_n824));
  INV_X1    g399(.A(KEYINPUT34), .ZN(new_n825));
  NOR2_X1   g400(.A1(new_n824), .A2(new_n825), .ZN(new_n826));
  XNOR2_X1  g401(.A(new_n826), .B(KEYINPUT89), .ZN(new_n827));
  AND2_X1   g402(.A1(new_n770), .A2(G24), .ZN(new_n828));
  AOI21_X1  g403(.A(new_n828), .B1(G290), .B2(new_n771), .ZN(new_n829));
  INV_X1    g404(.A(new_n829), .ZN(new_n830));
  AOI21_X1  g405(.A(KEYINPUT90), .B1(new_n830), .B2(G1986), .ZN(new_n831));
  OAI21_X1  g406(.A(new_n831), .B1(G1986), .B2(new_n830), .ZN(new_n832));
  NAND2_X1  g407(.A1(new_n481), .A2(G131), .ZN(new_n833));
  NAND2_X1  g408(.A1(new_n483), .A2(G119), .ZN(new_n834));
  NOR2_X1   g409(.A1(new_n463), .A2(G107), .ZN(new_n835));
  OAI21_X1  g410(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n836));
  OAI211_X1 g411(.A(new_n833), .B(new_n834), .C1(new_n835), .C2(new_n836), .ZN(new_n837));
  MUX2_X1   g412(.A(G25), .B(new_n837), .S(G29), .Z(new_n838));
  XOR2_X1   g413(.A(KEYINPUT35), .B(G1991), .Z(new_n839));
  INV_X1    g414(.A(new_n839), .ZN(new_n840));
  XNOR2_X1  g415(.A(new_n838), .B(new_n840), .ZN(new_n841));
  AOI211_X1 g416(.A(new_n832), .B(new_n841), .C1(new_n824), .C2(new_n825), .ZN(new_n842));
  NAND3_X1  g417(.A1(new_n827), .A2(KEYINPUT36), .A3(new_n842), .ZN(new_n843));
  NAND2_X1  g418(.A1(new_n811), .A2(new_n843), .ZN(new_n844));
  AOI21_X1  g419(.A(KEYINPUT36), .B1(new_n827), .B2(new_n842), .ZN(new_n845));
  NOR2_X1   g420(.A1(new_n844), .A2(new_n845), .ZN(G311));
  INV_X1    g421(.A(G311), .ZN(G150));
  INV_X1    g422(.A(KEYINPUT101), .ZN(new_n848));
  NAND3_X1  g423(.A1(new_n535), .A2(G67), .A3(new_n526), .ZN(new_n849));
  NAND2_X1  g424(.A1(G80), .A2(G543), .ZN(new_n850));
  NAND2_X1  g425(.A1(new_n849), .A2(new_n850), .ZN(new_n851));
  NAND2_X1  g426(.A1(new_n851), .A2(G651), .ZN(new_n852));
  NAND4_X1  g427(.A1(new_n535), .A2(G93), .A3(new_n526), .A4(new_n520), .ZN(new_n853));
  XNOR2_X1  g428(.A(KEYINPUT100), .B(G55), .ZN(new_n854));
  NAND2_X1  g429(.A1(new_n518), .A2(new_n854), .ZN(new_n855));
  NAND2_X1  g430(.A1(new_n853), .A2(new_n855), .ZN(new_n856));
  INV_X1    g431(.A(new_n856), .ZN(new_n857));
  AOI21_X1  g432(.A(new_n848), .B1(new_n852), .B2(new_n857), .ZN(new_n858));
  AOI21_X1  g433(.A(new_n514), .B1(new_n849), .B2(new_n850), .ZN(new_n859));
  NOR3_X1   g434(.A1(new_n859), .A2(new_n856), .A3(KEYINPUT101), .ZN(new_n860));
  OAI21_X1  g435(.A(new_n568), .B1(new_n858), .B2(new_n860), .ZN(new_n861));
  NAND2_X1  g436(.A1(new_n565), .A2(new_n566), .ZN(new_n862));
  NAND2_X1  g437(.A1(new_n562), .A2(KEYINPUT76), .ZN(new_n863));
  NAND3_X1  g438(.A1(new_n862), .A2(new_n863), .A3(G651), .ZN(new_n864));
  NAND4_X1  g439(.A1(new_n864), .A2(new_n559), .A3(new_n852), .A4(new_n857), .ZN(new_n865));
  NAND2_X1  g440(.A1(new_n861), .A2(new_n865), .ZN(new_n866));
  XOR2_X1   g441(.A(new_n866), .B(KEYINPUT38), .Z(new_n867));
  NAND2_X1  g442(.A1(new_n644), .A2(G559), .ZN(new_n868));
  XNOR2_X1  g443(.A(new_n867), .B(new_n868), .ZN(new_n869));
  AND2_X1   g444(.A1(new_n869), .A2(KEYINPUT39), .ZN(new_n870));
  NOR2_X1   g445(.A1(new_n869), .A2(KEYINPUT39), .ZN(new_n871));
  NOR3_X1   g446(.A1(new_n870), .A2(new_n871), .A3(G860), .ZN(new_n872));
  NAND3_X1  g447(.A1(new_n852), .A2(new_n857), .A3(new_n848), .ZN(new_n873));
  OAI21_X1  g448(.A(KEYINPUT101), .B1(new_n859), .B2(new_n856), .ZN(new_n874));
  NAND2_X1  g449(.A1(new_n873), .A2(new_n874), .ZN(new_n875));
  NAND2_X1  g450(.A1(new_n875), .A2(G860), .ZN(new_n876));
  XNOR2_X1  g451(.A(new_n876), .B(KEYINPUT37), .ZN(new_n877));
  OR2_X1    g452(.A1(new_n872), .A2(new_n877), .ZN(G145));
  NAND2_X1  g453(.A1(new_n504), .A2(KEYINPUT102), .ZN(new_n879));
  INV_X1    g454(.A(KEYINPUT102), .ZN(new_n880));
  OAI211_X1 g455(.A(new_n497), .B(new_n880), .C1(new_n502), .C2(new_n503), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n879), .A2(new_n881), .ZN(new_n882));
  AOI22_X1  g457(.A1(new_n490), .A2(new_n489), .B1(new_n470), .B2(new_n492), .ZN(new_n883));
  NAND2_X1  g458(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  INV_X1    g459(.A(KEYINPUT103), .ZN(new_n885));
  NAND2_X1  g460(.A1(new_n884), .A2(new_n885), .ZN(new_n886));
  AOI21_X1  g461(.A(new_n494), .B1(new_n879), .B2(new_n881), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n887), .A2(KEYINPUT103), .ZN(new_n888));
  NAND2_X1  g463(.A1(new_n886), .A2(new_n888), .ZN(new_n889));
  XNOR2_X1  g464(.A(new_n805), .B(new_n889), .ZN(new_n890));
  XNOR2_X1  g465(.A(new_n890), .B(new_n837), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n481), .A2(G142), .ZN(new_n892));
  NAND2_X1  g467(.A1(new_n483), .A2(G130), .ZN(new_n893));
  NOR2_X1   g468(.A1(new_n463), .A2(G118), .ZN(new_n894));
  OAI21_X1  g469(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n895));
  OAI211_X1 g470(.A(new_n892), .B(new_n893), .C1(new_n894), .C2(new_n895), .ZN(new_n896));
  XNOR2_X1  g471(.A(new_n896), .B(new_n662), .ZN(new_n897));
  XNOR2_X1  g472(.A(new_n761), .B(new_n787), .ZN(new_n898));
  XNOR2_X1  g473(.A(new_n897), .B(new_n898), .ZN(new_n899));
  XNOR2_X1  g474(.A(new_n891), .B(new_n899), .ZN(new_n900));
  XNOR2_X1  g475(.A(new_n487), .B(G160), .ZN(new_n901));
  XNOR2_X1  g476(.A(new_n658), .B(new_n901), .ZN(new_n902));
  AOI21_X1  g477(.A(G37), .B1(new_n900), .B2(new_n902), .ZN(new_n903));
  OAI21_X1  g478(.A(new_n903), .B1(new_n902), .B2(new_n900), .ZN(new_n904));
  XOR2_X1   g479(.A(KEYINPUT104), .B(KEYINPUT40), .Z(new_n905));
  XNOR2_X1  g480(.A(new_n904), .B(new_n905), .ZN(G395));
  NAND2_X1  g481(.A1(new_n875), .A2(new_n640), .ZN(new_n907));
  XNOR2_X1  g482(.A(G305), .B(G288), .ZN(new_n908));
  XNOR2_X1  g483(.A(G303), .B(G290), .ZN(new_n909));
  XNOR2_X1  g484(.A(new_n908), .B(new_n909), .ZN(new_n910));
  NOR2_X1   g485(.A1(new_n910), .A2(KEYINPUT42), .ZN(new_n911));
  XOR2_X1   g486(.A(new_n911), .B(KEYINPUT107), .Z(new_n912));
  NAND2_X1  g487(.A1(new_n910), .A2(KEYINPUT42), .ZN(new_n913));
  XNOR2_X1  g488(.A(new_n913), .B(KEYINPUT106), .ZN(new_n914));
  NOR2_X1   g489(.A1(new_n912), .A2(new_n914), .ZN(new_n915));
  XNOR2_X1  g490(.A(new_n866), .B(new_n648), .ZN(new_n916));
  OAI21_X1  g491(.A(new_n593), .B1(new_n591), .B2(new_n592), .ZN(new_n917));
  NAND3_X1  g492(.A1(new_n583), .A2(new_n587), .A3(KEYINPUT78), .ZN(new_n918));
  AND4_X1   g493(.A1(new_n917), .A2(new_n918), .A3(new_n636), .A4(new_n631), .ZN(new_n919));
  AOI22_X1  g494(.A1(new_n917), .A2(new_n918), .B1(new_n631), .B2(new_n636), .ZN(new_n920));
  NOR2_X1   g495(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  NOR2_X1   g496(.A1(new_n916), .A2(new_n921), .ZN(new_n922));
  INV_X1    g497(.A(KEYINPUT41), .ZN(new_n923));
  OAI21_X1  g498(.A(new_n923), .B1(new_n919), .B2(new_n920), .ZN(new_n924));
  OAI21_X1  g499(.A(new_n637), .B1(new_n588), .B2(new_n594), .ZN(new_n925));
  NAND4_X1  g500(.A1(new_n917), .A2(new_n918), .A3(new_n636), .A4(new_n631), .ZN(new_n926));
  XNOR2_X1  g501(.A(KEYINPUT105), .B(KEYINPUT41), .ZN(new_n927));
  INV_X1    g502(.A(new_n927), .ZN(new_n928));
  NAND3_X1  g503(.A1(new_n925), .A2(new_n926), .A3(new_n928), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n924), .A2(new_n929), .ZN(new_n930));
  AOI21_X1  g505(.A(new_n922), .B1(new_n916), .B2(new_n930), .ZN(new_n931));
  XNOR2_X1  g506(.A(new_n915), .B(new_n931), .ZN(new_n932));
  OAI21_X1  g507(.A(new_n907), .B1(new_n932), .B2(new_n640), .ZN(G295));
  OAI21_X1  g508(.A(new_n907), .B1(new_n932), .B2(new_n640), .ZN(G331));
  AOI22_X1  g509(.A1(new_n873), .A2(new_n874), .B1(new_n864), .B2(new_n559), .ZN(new_n935));
  NAND2_X1  g510(.A1(new_n852), .A2(new_n857), .ZN(new_n936));
  NOR2_X1   g511(.A1(new_n568), .A2(new_n936), .ZN(new_n937));
  AOI21_X1  g512(.A(G286), .B1(new_n601), .B2(new_n599), .ZN(new_n938));
  NOR2_X1   g513(.A1(G168), .A2(G171), .ZN(new_n939));
  OAI22_X1  g514(.A1(new_n935), .A2(new_n937), .B1(new_n938), .B2(new_n939), .ZN(new_n940));
  INV_X1    g515(.A(KEYINPUT110), .ZN(new_n941));
  AOI21_X1  g516(.A(KEYINPUT79), .B1(new_n597), .B2(new_n598), .ZN(new_n942));
  NOR3_X1   g517(.A1(new_n550), .A2(new_n556), .A3(new_n600), .ZN(new_n943));
  OAI21_X1  g518(.A(G168), .B1(new_n942), .B2(new_n943), .ZN(new_n944));
  OAI21_X1  g519(.A(G286), .B1(new_n550), .B2(new_n556), .ZN(new_n945));
  NAND4_X1  g520(.A1(new_n861), .A2(new_n944), .A3(new_n865), .A4(new_n945), .ZN(new_n946));
  NAND3_X1  g521(.A1(new_n940), .A2(new_n941), .A3(new_n946), .ZN(new_n947));
  OAI211_X1 g522(.A(new_n866), .B(KEYINPUT110), .C1(new_n938), .C2(new_n939), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n947), .A2(new_n948), .ZN(new_n949));
  INV_X1    g524(.A(new_n921), .ZN(new_n950));
  NAND2_X1  g525(.A1(new_n949), .A2(new_n950), .ZN(new_n951));
  NOR2_X1   g526(.A1(new_n938), .A2(new_n939), .ZN(new_n952));
  INV_X1    g527(.A(KEYINPUT109), .ZN(new_n953));
  NAND4_X1  g528(.A1(new_n952), .A2(new_n953), .A3(new_n861), .A4(new_n865), .ZN(new_n954));
  NAND3_X1  g529(.A1(new_n940), .A2(KEYINPUT109), .A3(new_n946), .ZN(new_n955));
  NAND3_X1  g530(.A1(new_n930), .A2(new_n954), .A3(new_n955), .ZN(new_n956));
  NAND3_X1  g531(.A1(new_n951), .A2(new_n910), .A3(new_n956), .ZN(new_n957));
  INV_X1    g532(.A(G37), .ZN(new_n958));
  NAND2_X1  g533(.A1(new_n957), .A2(new_n958), .ZN(new_n959));
  INV_X1    g534(.A(new_n959), .ZN(new_n960));
  XNOR2_X1  g535(.A(KEYINPUT108), .B(KEYINPUT43), .ZN(new_n961));
  INV_X1    g536(.A(new_n910), .ZN(new_n962));
  NOR3_X1   g537(.A1(new_n919), .A2(new_n920), .A3(KEYINPUT41), .ZN(new_n963));
  AOI21_X1  g538(.A(new_n927), .B1(new_n925), .B2(new_n926), .ZN(new_n964));
  NOR2_X1   g539(.A1(new_n963), .A2(new_n964), .ZN(new_n965));
  AND3_X1   g540(.A1(new_n965), .A2(new_n948), .A3(new_n947), .ZN(new_n966));
  AOI21_X1  g541(.A(new_n921), .B1(new_n955), .B2(new_n954), .ZN(new_n967));
  OAI21_X1  g542(.A(new_n962), .B1(new_n966), .B2(new_n967), .ZN(new_n968));
  NAND3_X1  g543(.A1(new_n960), .A2(new_n961), .A3(new_n968), .ZN(new_n969));
  AND3_X1   g544(.A1(new_n930), .A2(new_n954), .A3(new_n955), .ZN(new_n970));
  AOI21_X1  g545(.A(new_n921), .B1(new_n947), .B2(new_n948), .ZN(new_n971));
  OAI21_X1  g546(.A(new_n962), .B1(new_n970), .B2(new_n971), .ZN(new_n972));
  AND2_X1   g547(.A1(new_n960), .A2(new_n972), .ZN(new_n973));
  OAI21_X1  g548(.A(new_n969), .B1(new_n961), .B2(new_n973), .ZN(new_n974));
  INV_X1    g549(.A(KEYINPUT44), .ZN(new_n975));
  NAND2_X1  g550(.A1(new_n974), .A2(new_n975), .ZN(new_n976));
  INV_X1    g551(.A(new_n967), .ZN(new_n977));
  NAND3_X1  g552(.A1(new_n965), .A2(new_n948), .A3(new_n947), .ZN(new_n978));
  AOI21_X1  g553(.A(new_n910), .B1(new_n977), .B2(new_n978), .ZN(new_n979));
  OAI21_X1  g554(.A(KEYINPUT43), .B1(new_n959), .B2(new_n979), .ZN(new_n980));
  INV_X1    g555(.A(KEYINPUT112), .ZN(new_n981));
  NAND2_X1  g556(.A1(new_n980), .A2(new_n981), .ZN(new_n982));
  OAI211_X1 g557(.A(KEYINPUT112), .B(KEYINPUT43), .C1(new_n959), .C2(new_n979), .ZN(new_n983));
  NAND2_X1  g558(.A1(new_n982), .A2(new_n983), .ZN(new_n984));
  NAND4_X1  g559(.A1(new_n972), .A2(new_n957), .A3(new_n958), .A4(new_n961), .ZN(new_n985));
  XNOR2_X1  g560(.A(new_n985), .B(KEYINPUT111), .ZN(new_n986));
  AND4_X1   g561(.A1(KEYINPUT113), .A2(new_n984), .A3(new_n986), .A4(KEYINPUT44), .ZN(new_n987));
  AOI21_X1  g562(.A(new_n975), .B1(new_n982), .B2(new_n983), .ZN(new_n988));
  AOI21_X1  g563(.A(KEYINPUT113), .B1(new_n988), .B2(new_n986), .ZN(new_n989));
  OAI21_X1  g564(.A(new_n976), .B1(new_n987), .B2(new_n989), .ZN(G397));
  INV_X1    g565(.A(G1384), .ZN(new_n991));
  NAND3_X1  g566(.A1(new_n886), .A2(new_n888), .A3(new_n991), .ZN(new_n992));
  INV_X1    g567(.A(KEYINPUT114), .ZN(new_n993));
  OR2_X1    g568(.A1(new_n992), .A2(new_n993), .ZN(new_n994));
  XOR2_X1   g569(.A(KEYINPUT115), .B(KEYINPUT45), .Z(new_n995));
  INV_X1    g570(.A(new_n995), .ZN(new_n996));
  AOI21_X1  g571(.A(new_n996), .B1(new_n992), .B2(new_n993), .ZN(new_n997));
  AND2_X1   g572(.A1(new_n994), .A2(new_n997), .ZN(new_n998));
  INV_X1    g573(.A(G40), .ZN(new_n999));
  NOR3_X1   g574(.A1(new_n472), .A2(new_n999), .A3(new_n475), .ZN(new_n1000));
  AND2_X1   g575(.A1(new_n998), .A2(new_n1000), .ZN(new_n1001));
  XNOR2_X1  g576(.A(new_n804), .B(new_n807), .ZN(new_n1002));
  INV_X1    g577(.A(G1996), .ZN(new_n1003));
  XNOR2_X1  g578(.A(new_n761), .B(new_n1003), .ZN(new_n1004));
  NAND2_X1  g579(.A1(new_n837), .A2(new_n840), .ZN(new_n1005));
  OR2_X1    g580(.A1(new_n837), .A2(new_n840), .ZN(new_n1006));
  NAND4_X1  g581(.A1(new_n1002), .A2(new_n1004), .A3(new_n1005), .A4(new_n1006), .ZN(new_n1007));
  XNOR2_X1  g582(.A(G290), .B(G1986), .ZN(new_n1008));
  OAI21_X1  g583(.A(new_n1001), .B1(new_n1007), .B2(new_n1008), .ZN(new_n1009));
  NOR2_X1   g584(.A1(new_n591), .A2(new_n592), .ZN(new_n1010));
  XNOR2_X1  g585(.A(new_n1010), .B(KEYINPUT57), .ZN(new_n1011));
  NAND4_X1  g586(.A1(new_n886), .A2(new_n888), .A3(KEYINPUT45), .A4(new_n991), .ZN(new_n1012));
  INV_X1    g587(.A(new_n474), .ZN(new_n1013));
  NAND2_X1  g588(.A1(new_n1013), .A2(G2105), .ZN(new_n1014));
  NAND4_X1  g589(.A1(new_n1014), .A2(G40), .A3(new_n466), .A4(new_n471), .ZN(new_n1015));
  OAI21_X1  g590(.A(new_n991), .B1(new_n494), .B2(new_n504), .ZN(new_n1016));
  AOI21_X1  g591(.A(new_n1015), .B1(new_n1016), .B2(new_n995), .ZN(new_n1017));
  XNOR2_X1  g592(.A(KEYINPUT56), .B(G2072), .ZN(new_n1018));
  NAND3_X1  g593(.A1(new_n1012), .A2(new_n1017), .A3(new_n1018), .ZN(new_n1019));
  INV_X1    g594(.A(new_n504), .ZN(new_n1020));
  AOI21_X1  g595(.A(G1384), .B1(new_n883), .B2(new_n1020), .ZN(new_n1021));
  INV_X1    g596(.A(KEYINPUT50), .ZN(new_n1022));
  AOI21_X1  g597(.A(new_n1015), .B1(new_n1021), .B2(new_n1022), .ZN(new_n1023));
  NOR2_X1   g598(.A1(new_n887), .A2(G1384), .ZN(new_n1024));
  OAI21_X1  g599(.A(new_n1023), .B1(new_n1024), .B2(new_n1022), .ZN(new_n1025));
  NAND2_X1  g600(.A1(new_n1025), .A2(new_n791), .ZN(new_n1026));
  AOI21_X1  g601(.A(new_n1011), .B1(new_n1019), .B2(new_n1026), .ZN(new_n1027));
  NAND3_X1  g602(.A1(new_n1019), .A2(new_n1026), .A3(new_n1011), .ZN(new_n1028));
  AOI21_X1  g603(.A(new_n1015), .B1(KEYINPUT50), .B2(new_n1016), .ZN(new_n1029));
  NAND3_X1  g604(.A1(new_n884), .A2(new_n1022), .A3(new_n991), .ZN(new_n1030));
  AOI21_X1  g605(.A(G1348), .B1(new_n1029), .B2(new_n1030), .ZN(new_n1031));
  NAND3_X1  g606(.A1(new_n884), .A2(new_n1000), .A3(new_n991), .ZN(new_n1032));
  NOR2_X1   g607(.A1(new_n1032), .A2(G2067), .ZN(new_n1033));
  NOR2_X1   g608(.A1(new_n1031), .A2(new_n1033), .ZN(new_n1034));
  NOR2_X1   g609(.A1(new_n1034), .A2(new_n637), .ZN(new_n1035));
  AOI21_X1  g610(.A(new_n1027), .B1(new_n1028), .B2(new_n1035), .ZN(new_n1036));
  INV_X1    g611(.A(KEYINPUT60), .ZN(new_n1037));
  OAI21_X1  g612(.A(new_n1037), .B1(new_n1031), .B2(new_n1033), .ZN(new_n1038));
  INV_X1    g613(.A(KEYINPUT122), .ZN(new_n1039));
  AND3_X1   g614(.A1(new_n1038), .A2(new_n1039), .A3(new_n644), .ZN(new_n1040));
  AOI21_X1  g615(.A(new_n1039), .B1(new_n1038), .B2(new_n644), .ZN(new_n1041));
  NAND2_X1  g616(.A1(new_n1034), .A2(KEYINPUT60), .ZN(new_n1042));
  INV_X1    g617(.A(new_n1042), .ZN(new_n1043));
  NOR3_X1   g618(.A1(new_n1040), .A2(new_n1041), .A3(new_n1043), .ZN(new_n1044));
  NAND2_X1  g619(.A1(new_n1029), .A2(new_n1030), .ZN(new_n1045));
  INV_X1    g620(.A(G1348), .ZN(new_n1046));
  NAND2_X1  g621(.A1(new_n1045), .A2(new_n1046), .ZN(new_n1047));
  INV_X1    g622(.A(new_n1032), .ZN(new_n1048));
  NAND2_X1  g623(.A1(new_n1048), .A2(new_n807), .ZN(new_n1049));
  AOI21_X1  g624(.A(KEYINPUT60), .B1(new_n1047), .B2(new_n1049), .ZN(new_n1050));
  OAI21_X1  g625(.A(KEYINPUT122), .B1(new_n1050), .B2(new_n637), .ZN(new_n1051));
  NAND3_X1  g626(.A1(new_n1038), .A2(new_n1039), .A3(new_n644), .ZN(new_n1052));
  AOI21_X1  g627(.A(new_n1042), .B1(new_n1051), .B2(new_n1052), .ZN(new_n1053));
  NOR2_X1   g628(.A1(new_n1044), .A2(new_n1053), .ZN(new_n1054));
  INV_X1    g629(.A(KEYINPUT121), .ZN(new_n1055));
  INV_X1    g630(.A(KEYINPUT61), .ZN(new_n1056));
  NAND3_X1  g631(.A1(new_n1028), .A2(new_n1055), .A3(new_n1056), .ZN(new_n1057));
  OAI21_X1  g632(.A(new_n1057), .B1(new_n1056), .B2(new_n1028), .ZN(new_n1058));
  NAND3_X1  g633(.A1(new_n1012), .A2(new_n1003), .A3(new_n1017), .ZN(new_n1059));
  XNOR2_X1  g634(.A(KEYINPUT58), .B(G1341), .ZN(new_n1060));
  OAI21_X1  g635(.A(new_n1059), .B1(new_n1048), .B2(new_n1060), .ZN(new_n1061));
  NAND2_X1  g636(.A1(new_n1061), .A2(new_n569), .ZN(new_n1062));
  XNOR2_X1  g637(.A(KEYINPUT120), .B(KEYINPUT59), .ZN(new_n1063));
  INV_X1    g638(.A(new_n1063), .ZN(new_n1064));
  NAND2_X1  g639(.A1(new_n1062), .A2(new_n1064), .ZN(new_n1065));
  NAND3_X1  g640(.A1(new_n1061), .A2(new_n569), .A3(new_n1063), .ZN(new_n1066));
  NAND3_X1  g641(.A1(new_n1058), .A2(new_n1065), .A3(new_n1066), .ZN(new_n1067));
  OAI21_X1  g642(.A(new_n1036), .B1(new_n1054), .B2(new_n1067), .ZN(new_n1068));
  NAND2_X1  g643(.A1(G303), .A2(G8), .ZN(new_n1069));
  XNOR2_X1  g644(.A(new_n1069), .B(KEYINPUT55), .ZN(new_n1070));
  INV_X1    g645(.A(new_n1070), .ZN(new_n1071));
  XOR2_X1   g646(.A(KEYINPUT116), .B(G1971), .Z(new_n1072));
  AOI21_X1  g647(.A(new_n1072), .B1(new_n1012), .B2(new_n1017), .ZN(new_n1073));
  NOR2_X1   g648(.A1(new_n1045), .A2(G2090), .ZN(new_n1074));
  OAI211_X1 g649(.A(new_n1071), .B(G8), .C1(new_n1073), .C2(new_n1074), .ZN(new_n1075));
  OR3_X1    g650(.A1(new_n615), .A2(new_n618), .A3(G1981), .ZN(new_n1076));
  OAI21_X1  g651(.A(G1981), .B1(new_n615), .B2(new_n618), .ZN(new_n1077));
  NAND2_X1  g652(.A1(new_n1076), .A2(new_n1077), .ZN(new_n1078));
  INV_X1    g653(.A(KEYINPUT49), .ZN(new_n1079));
  NAND2_X1  g654(.A1(new_n1078), .A2(new_n1079), .ZN(new_n1080));
  NAND3_X1  g655(.A1(new_n1076), .A2(KEYINPUT49), .A3(new_n1077), .ZN(new_n1081));
  NAND4_X1  g656(.A1(new_n1080), .A2(G8), .A3(new_n1032), .A4(new_n1081), .ZN(new_n1082));
  INV_X1    g657(.A(G288), .ZN(new_n1083));
  NAND2_X1  g658(.A1(new_n1083), .A2(G1976), .ZN(new_n1084));
  NAND3_X1  g659(.A1(new_n1084), .A2(new_n1032), .A3(G8), .ZN(new_n1085));
  NAND2_X1  g660(.A1(new_n1085), .A2(KEYINPUT52), .ZN(new_n1086));
  INV_X1    g661(.A(G1976), .ZN(new_n1087));
  AOI21_X1  g662(.A(KEYINPUT52), .B1(G288), .B2(new_n1087), .ZN(new_n1088));
  NAND4_X1  g663(.A1(new_n1084), .A2(new_n1088), .A3(new_n1032), .A4(G8), .ZN(new_n1089));
  AND3_X1   g664(.A1(new_n1082), .A2(new_n1086), .A3(new_n1089), .ZN(new_n1090));
  NAND2_X1  g665(.A1(new_n1075), .A2(new_n1090), .ZN(new_n1091));
  INV_X1    g666(.A(new_n1073), .ZN(new_n1092));
  NOR2_X1   g667(.A1(new_n1025), .A2(G2090), .ZN(new_n1093));
  INV_X1    g668(.A(new_n1093), .ZN(new_n1094));
  NAND3_X1  g669(.A1(new_n1092), .A2(new_n1094), .A3(KEYINPUT117), .ZN(new_n1095));
  INV_X1    g670(.A(KEYINPUT117), .ZN(new_n1096));
  OAI21_X1  g671(.A(new_n1096), .B1(new_n1073), .B2(new_n1093), .ZN(new_n1097));
  NAND3_X1  g672(.A1(new_n1095), .A2(G8), .A3(new_n1097), .ZN(new_n1098));
  AOI21_X1  g673(.A(new_n1091), .B1(new_n1098), .B2(new_n1070), .ZN(new_n1099));
  INV_X1    g674(.A(G2084), .ZN(new_n1100));
  NAND3_X1  g675(.A1(new_n1029), .A2(new_n1030), .A3(new_n1100), .ZN(new_n1101));
  INV_X1    g676(.A(new_n1101), .ZN(new_n1102));
  AOI21_X1  g677(.A(new_n1015), .B1(new_n1021), .B2(new_n996), .ZN(new_n1103));
  INV_X1    g678(.A(KEYINPUT45), .ZN(new_n1104));
  OAI21_X1  g679(.A(new_n1104), .B1(new_n887), .B2(G1384), .ZN(new_n1105));
  AOI21_X1  g680(.A(G1966), .B1(new_n1103), .B2(new_n1105), .ZN(new_n1106));
  OAI21_X1  g681(.A(G286), .B1(new_n1102), .B2(new_n1106), .ZN(new_n1107));
  INV_X1    g682(.A(G1966), .ZN(new_n1108));
  AOI21_X1  g683(.A(KEYINPUT45), .B1(new_n884), .B2(new_n991), .ZN(new_n1109));
  OAI21_X1  g684(.A(new_n1000), .B1(new_n1016), .B2(new_n995), .ZN(new_n1110));
  OAI21_X1  g685(.A(new_n1108), .B1(new_n1109), .B2(new_n1110), .ZN(new_n1111));
  NAND3_X1  g686(.A1(new_n1111), .A2(G168), .A3(new_n1101), .ZN(new_n1112));
  NAND3_X1  g687(.A1(new_n1107), .A2(new_n1112), .A3(G8), .ZN(new_n1113));
  OAI21_X1  g688(.A(G8), .B1(new_n1102), .B2(new_n1106), .ZN(new_n1114));
  INV_X1    g689(.A(KEYINPUT123), .ZN(new_n1115));
  NAND2_X1  g690(.A1(new_n1114), .A2(new_n1115), .ZN(new_n1116));
  NAND3_X1  g691(.A1(new_n1113), .A2(KEYINPUT51), .A3(new_n1116), .ZN(new_n1117));
  INV_X1    g692(.A(G8), .ZN(new_n1118));
  AOI21_X1  g693(.A(new_n1118), .B1(new_n1111), .B2(new_n1101), .ZN(new_n1119));
  OAI21_X1  g694(.A(KEYINPUT51), .B1(new_n1119), .B2(KEYINPUT123), .ZN(new_n1120));
  NAND3_X1  g695(.A1(new_n1120), .A2(G8), .A3(new_n1112), .ZN(new_n1121));
  INV_X1    g696(.A(KEYINPUT124), .ZN(new_n1122));
  AND3_X1   g697(.A1(new_n1117), .A2(new_n1121), .A3(new_n1122), .ZN(new_n1123));
  AOI21_X1  g698(.A(new_n1122), .B1(new_n1117), .B2(new_n1121), .ZN(new_n1124));
  NOR2_X1   g699(.A1(new_n1123), .A2(new_n1124), .ZN(new_n1125));
  AOI21_X1  g700(.A(G1961), .B1(new_n1029), .B2(new_n1030), .ZN(new_n1126));
  INV_X1    g701(.A(G2078), .ZN(new_n1127));
  NAND3_X1  g702(.A1(new_n1012), .A2(new_n1127), .A3(new_n1017), .ZN(new_n1128));
  INV_X1    g703(.A(KEYINPUT53), .ZN(new_n1129));
  AOI21_X1  g704(.A(new_n1126), .B1(new_n1128), .B2(new_n1129), .ZN(new_n1130));
  NOR2_X1   g705(.A1(new_n1109), .A2(new_n1110), .ZN(new_n1131));
  NOR2_X1   g706(.A1(new_n1129), .A2(G2078), .ZN(new_n1132));
  NAND2_X1  g707(.A1(new_n1131), .A2(new_n1132), .ZN(new_n1133));
  NAND2_X1  g708(.A1(new_n1130), .A2(new_n1133), .ZN(new_n1134));
  NAND2_X1  g709(.A1(new_n1134), .A2(new_n602), .ZN(new_n1135));
  AOI21_X1  g710(.A(new_n463), .B1(new_n1013), .B2(KEYINPUT126), .ZN(new_n1136));
  OAI21_X1  g711(.A(new_n1136), .B1(KEYINPUT126), .B2(new_n1013), .ZN(new_n1137));
  AND3_X1   g712(.A1(new_n1137), .A2(G40), .A3(new_n1132), .ZN(new_n1138));
  XNOR2_X1  g713(.A(new_n472), .B(KEYINPUT125), .ZN(new_n1139));
  NAND3_X1  g714(.A1(new_n1012), .A2(new_n1138), .A3(new_n1139), .ZN(new_n1140));
  OAI21_X1  g715(.A(new_n1130), .B1(new_n998), .B2(new_n1140), .ZN(new_n1141));
  OAI21_X1  g716(.A(new_n1135), .B1(new_n1141), .B2(new_n602), .ZN(new_n1142));
  INV_X1    g717(.A(KEYINPUT54), .ZN(new_n1143));
  AND2_X1   g718(.A1(new_n1130), .A2(new_n1133), .ZN(new_n1144));
  AOI21_X1  g719(.A(new_n1143), .B1(new_n1144), .B2(G301), .ZN(new_n1145));
  NAND2_X1  g720(.A1(new_n1141), .A2(G171), .ZN(new_n1146));
  AOI22_X1  g721(.A1(new_n1142), .A2(new_n1143), .B1(new_n1145), .B2(new_n1146), .ZN(new_n1147));
  NAND4_X1  g722(.A1(new_n1068), .A2(new_n1099), .A3(new_n1125), .A4(new_n1147), .ZN(new_n1148));
  INV_X1    g723(.A(KEYINPUT62), .ZN(new_n1149));
  OAI21_X1  g724(.A(new_n1149), .B1(new_n1123), .B2(new_n1124), .ZN(new_n1150));
  NAND2_X1  g725(.A1(new_n1117), .A2(new_n1121), .ZN(new_n1151));
  NAND2_X1  g726(.A1(new_n1151), .A2(KEYINPUT124), .ZN(new_n1152));
  NAND3_X1  g727(.A1(new_n1117), .A2(new_n1121), .A3(new_n1122), .ZN(new_n1153));
  NAND3_X1  g728(.A1(new_n1152), .A2(KEYINPUT62), .A3(new_n1153), .ZN(new_n1154));
  AOI211_X1 g729(.A(new_n1135), .B(new_n1091), .C1(new_n1070), .C2(new_n1098), .ZN(new_n1155));
  NAND3_X1  g730(.A1(new_n1150), .A2(new_n1154), .A3(new_n1155), .ZN(new_n1156));
  NAND3_X1  g731(.A1(new_n1082), .A2(new_n1087), .A3(new_n1083), .ZN(new_n1157));
  AOI211_X1 g732(.A(new_n1118), .B(new_n1048), .C1(new_n1157), .C2(new_n1076), .ZN(new_n1158));
  INV_X1    g733(.A(new_n1075), .ZN(new_n1159));
  AOI21_X1  g734(.A(new_n1158), .B1(new_n1159), .B2(new_n1090), .ZN(new_n1160));
  NAND3_X1  g735(.A1(new_n1148), .A2(new_n1156), .A3(new_n1160), .ZN(new_n1161));
  NOR2_X1   g736(.A1(new_n1073), .A2(new_n1074), .ZN(new_n1162));
  NOR2_X1   g737(.A1(new_n1162), .A2(new_n1118), .ZN(new_n1163));
  OAI21_X1  g738(.A(new_n1090), .B1(new_n1163), .B2(new_n1071), .ZN(new_n1164));
  NAND2_X1  g739(.A1(new_n1164), .A2(KEYINPUT119), .ZN(new_n1165));
  INV_X1    g740(.A(KEYINPUT119), .ZN(new_n1166));
  OAI211_X1 g741(.A(new_n1166), .B(new_n1090), .C1(new_n1163), .C2(new_n1071), .ZN(new_n1167));
  NOR2_X1   g742(.A1(new_n1114), .A2(G286), .ZN(new_n1168));
  AND3_X1   g743(.A1(new_n1075), .A2(new_n1168), .A3(KEYINPUT63), .ZN(new_n1169));
  NAND3_X1  g744(.A1(new_n1165), .A2(new_n1167), .A3(new_n1169), .ZN(new_n1170));
  AOI21_X1  g745(.A(KEYINPUT63), .B1(new_n1099), .B2(new_n1168), .ZN(new_n1171));
  INV_X1    g746(.A(KEYINPUT118), .ZN(new_n1172));
  OAI21_X1  g747(.A(new_n1170), .B1(new_n1171), .B2(new_n1172), .ZN(new_n1173));
  AOI211_X1 g748(.A(KEYINPUT118), .B(KEYINPUT63), .C1(new_n1099), .C2(new_n1168), .ZN(new_n1174));
  NOR2_X1   g749(.A1(new_n1173), .A2(new_n1174), .ZN(new_n1175));
  OAI21_X1  g750(.A(new_n1009), .B1(new_n1161), .B2(new_n1175), .ZN(new_n1176));
  NAND2_X1  g751(.A1(new_n1002), .A2(new_n1004), .ZN(new_n1177));
  OAI22_X1  g752(.A1(new_n1177), .A2(new_n1006), .B1(G2067), .B2(new_n804), .ZN(new_n1178));
  NAND2_X1  g753(.A1(new_n1001), .A2(new_n1178), .ZN(new_n1179));
  NOR2_X1   g754(.A1(G290), .A2(G1986), .ZN(new_n1180));
  NAND2_X1  g755(.A1(new_n1001), .A2(new_n1180), .ZN(new_n1181));
  XNOR2_X1  g756(.A(KEYINPUT127), .B(KEYINPUT48), .ZN(new_n1182));
  NAND2_X1  g757(.A1(new_n1181), .A2(new_n1182), .ZN(new_n1183));
  NAND2_X1  g758(.A1(new_n1001), .A2(new_n1007), .ZN(new_n1184));
  NAND2_X1  g759(.A1(new_n1183), .A2(new_n1184), .ZN(new_n1185));
  NOR2_X1   g760(.A1(new_n1181), .A2(new_n1182), .ZN(new_n1186));
  OAI21_X1  g761(.A(new_n1179), .B1(new_n1185), .B2(new_n1186), .ZN(new_n1187));
  AND2_X1   g762(.A1(new_n1001), .A2(new_n1003), .ZN(new_n1188));
  OR2_X1    g763(.A1(new_n1188), .A2(KEYINPUT46), .ZN(new_n1189));
  NAND2_X1  g764(.A1(new_n1188), .A2(KEYINPUT46), .ZN(new_n1190));
  INV_X1    g765(.A(new_n1002), .ZN(new_n1191));
  OAI21_X1  g766(.A(new_n1001), .B1(new_n761), .B2(new_n1191), .ZN(new_n1192));
  NAND3_X1  g767(.A1(new_n1189), .A2(new_n1190), .A3(new_n1192), .ZN(new_n1193));
  NAND2_X1  g768(.A1(new_n1193), .A2(KEYINPUT47), .ZN(new_n1194));
  INV_X1    g769(.A(KEYINPUT47), .ZN(new_n1195));
  NAND4_X1  g770(.A1(new_n1189), .A2(new_n1195), .A3(new_n1190), .A4(new_n1192), .ZN(new_n1196));
  AOI21_X1  g771(.A(new_n1187), .B1(new_n1194), .B2(new_n1196), .ZN(new_n1197));
  NAND2_X1  g772(.A1(new_n1176), .A2(new_n1197), .ZN(G329));
  assign    G231 = 1'b0;
  NOR4_X1   g773(.A1(G229), .A2(G401), .A3(new_n461), .A4(G227), .ZN(new_n1200));
  NAND3_X1  g774(.A1(new_n1200), .A2(new_n974), .A3(new_n904), .ZN(G225));
  INV_X1    g775(.A(G225), .ZN(G308));
endmodule


