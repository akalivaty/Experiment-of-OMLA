

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300,
         n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311,
         n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322,
         n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333,
         n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344,
         n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355,
         n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
         n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
         n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
         n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
         n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410,
         n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421,
         n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432,
         n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443,
         n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454,
         n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465,
         n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
         n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487,
         n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
         n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
         n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579;

  NOR2_X2 U322 ( .A1(n514), .A2(n469), .ZN(n470) );
  XNOR2_X1 U323 ( .A(n461), .B(KEYINPUT25), .ZN(n462) );
  XOR2_X2 U324 ( .A(KEYINPUT38), .B(n493), .Z(n499) );
  XOR2_X1 U325 ( .A(n403), .B(n402), .Z(n290) );
  XOR2_X1 U326 ( .A(G71GAT), .B(n438), .Z(n291) );
  XOR2_X1 U327 ( .A(G190GAT), .B(G99GAT), .Z(n292) );
  AND2_X1 U328 ( .A1(n525), .A2(n516), .ZN(n459) );
  XNOR2_X1 U329 ( .A(KEYINPUT45), .B(KEYINPUT64), .ZN(n348) );
  XNOR2_X1 U330 ( .A(n349), .B(n348), .ZN(n367) );
  XNOR2_X1 U331 ( .A(G8GAT), .B(G183GAT), .ZN(n334) );
  XNOR2_X1 U332 ( .A(n334), .B(G211GAT), .ZN(n399) );
  XNOR2_X1 U333 ( .A(n447), .B(n446), .ZN(n448) );
  XNOR2_X1 U334 ( .A(n449), .B(n448), .ZN(n451) );
  XOR2_X1 U335 ( .A(n550), .B(KEYINPUT83), .Z(n534) );
  XNOR2_X1 U336 ( .A(n453), .B(G190GAT), .ZN(n454) );
  XNOR2_X1 U337 ( .A(n455), .B(n454), .ZN(G1351GAT) );
  XNOR2_X1 U338 ( .A(G134GAT), .B(G162GAT), .ZN(n293) );
  XNOR2_X1 U339 ( .A(n293), .B(KEYINPUT82), .ZN(n315) );
  XOR2_X1 U340 ( .A(KEYINPUT9), .B(KEYINPUT10), .Z(n294) );
  XNOR2_X1 U341 ( .A(n315), .B(n294), .ZN(n298) );
  XOR2_X1 U342 ( .A(KEYINPUT81), .B(KEYINPUT11), .Z(n296) );
  NAND2_X1 U343 ( .A1(G232GAT), .A2(G233GAT), .ZN(n295) );
  XNOR2_X1 U344 ( .A(n296), .B(n295), .ZN(n297) );
  XNOR2_X1 U345 ( .A(n298), .B(n297), .ZN(n301) );
  XOR2_X1 U346 ( .A(G92GAT), .B(G218GAT), .Z(n300) );
  XNOR2_X1 U347 ( .A(G36GAT), .B(G190GAT), .ZN(n299) );
  XNOR2_X1 U348 ( .A(n300), .B(n299), .ZN(n402) );
  XOR2_X1 U349 ( .A(n301), .B(n402), .Z(n309) );
  XNOR2_X1 U350 ( .A(G50GAT), .B(KEYINPUT7), .ZN(n302) );
  XNOR2_X1 U351 ( .A(n302), .B(G29GAT), .ZN(n303) );
  XOR2_X1 U352 ( .A(n303), .B(KEYINPUT8), .Z(n305) );
  XNOR2_X1 U353 ( .A(G43GAT), .B(KEYINPUT72), .ZN(n304) );
  XNOR2_X1 U354 ( .A(n305), .B(n304), .ZN(n379) );
  XOR2_X1 U355 ( .A(KEYINPUT78), .B(G85GAT), .Z(n307) );
  XNOR2_X1 U356 ( .A(G99GAT), .B(G106GAT), .ZN(n306) );
  XNOR2_X1 U357 ( .A(n307), .B(n306), .ZN(n362) );
  XNOR2_X1 U358 ( .A(n379), .B(n362), .ZN(n308) );
  XNOR2_X1 U359 ( .A(n309), .B(n308), .ZN(n550) );
  XOR2_X1 U360 ( .A(KEYINPUT0), .B(G127GAT), .Z(n311) );
  XNOR2_X1 U361 ( .A(KEYINPUT88), .B(G120GAT), .ZN(n310) );
  XNOR2_X1 U362 ( .A(n311), .B(n310), .ZN(n312) );
  XNOR2_X1 U363 ( .A(G113GAT), .B(n312), .ZN(n450) );
  INV_X1 U364 ( .A(n450), .ZN(n330) );
  XOR2_X1 U365 ( .A(G148GAT), .B(KEYINPUT3), .Z(n314) );
  XNOR2_X1 U366 ( .A(KEYINPUT96), .B(KEYINPUT2), .ZN(n313) );
  XNOR2_X1 U367 ( .A(n314), .B(n313), .ZN(n423) );
  XNOR2_X1 U368 ( .A(n423), .B(n315), .ZN(n328) );
  XOR2_X1 U369 ( .A(G85GAT), .B(G155GAT), .Z(n317) );
  XNOR2_X1 U370 ( .A(G29GAT), .B(G141GAT), .ZN(n316) );
  XNOR2_X1 U371 ( .A(n317), .B(n316), .ZN(n321) );
  XOR2_X1 U372 ( .A(KEYINPUT4), .B(KEYINPUT6), .Z(n319) );
  XNOR2_X1 U373 ( .A(KEYINPUT1), .B(KEYINPUT5), .ZN(n318) );
  XNOR2_X1 U374 ( .A(n319), .B(n318), .ZN(n320) );
  XOR2_X1 U375 ( .A(n321), .B(n320), .Z(n326) );
  XOR2_X1 U376 ( .A(G57GAT), .B(KEYINPUT99), .Z(n323) );
  NAND2_X1 U377 ( .A1(G225GAT), .A2(G233GAT), .ZN(n322) );
  XNOR2_X1 U378 ( .A(n323), .B(n322), .ZN(n324) );
  XNOR2_X1 U379 ( .A(G1GAT), .B(n324), .ZN(n325) );
  XNOR2_X1 U380 ( .A(n326), .B(n325), .ZN(n327) );
  XNOR2_X1 U381 ( .A(n328), .B(n327), .ZN(n329) );
  XNOR2_X1 U382 ( .A(n330), .B(n329), .ZN(n514) );
  XNOR2_X1 U383 ( .A(G15GAT), .B(G1GAT), .ZN(n331) );
  XNOR2_X1 U384 ( .A(n331), .B(KEYINPUT73), .ZN(n375) );
  XOR2_X1 U385 ( .A(KEYINPUT75), .B(KEYINPUT13), .Z(n333) );
  XNOR2_X1 U386 ( .A(G71GAT), .B(G57GAT), .ZN(n332) );
  XNOR2_X1 U387 ( .A(n333), .B(n332), .ZN(n361) );
  XNOR2_X1 U388 ( .A(n375), .B(n361), .ZN(n347) );
  XOR2_X1 U389 ( .A(G155GAT), .B(G78GAT), .Z(n426) );
  XOR2_X1 U390 ( .A(n399), .B(n426), .Z(n336) );
  XNOR2_X1 U391 ( .A(G22GAT), .B(G127GAT), .ZN(n335) );
  XNOR2_X1 U392 ( .A(n336), .B(n335), .ZN(n340) );
  XOR2_X1 U393 ( .A(KEYINPUT15), .B(KEYINPUT14), .Z(n338) );
  NAND2_X1 U394 ( .A1(G231GAT), .A2(G233GAT), .ZN(n337) );
  XNOR2_X1 U395 ( .A(n338), .B(n337), .ZN(n339) );
  XOR2_X1 U396 ( .A(n340), .B(n339), .Z(n345) );
  XOR2_X1 U397 ( .A(KEYINPUT12), .B(KEYINPUT86), .Z(n342) );
  XNOR2_X1 U398 ( .A(G64GAT), .B(KEYINPUT85), .ZN(n341) );
  XNOR2_X1 U399 ( .A(n342), .B(n341), .ZN(n343) );
  XNOR2_X1 U400 ( .A(n343), .B(KEYINPUT84), .ZN(n344) );
  XNOR2_X1 U401 ( .A(n345), .B(n344), .ZN(n346) );
  XNOR2_X1 U402 ( .A(n347), .B(n346), .ZN(n546) );
  INV_X1 U403 ( .A(n546), .ZN(n574) );
  XNOR2_X1 U404 ( .A(KEYINPUT36), .B(n534), .ZN(n576) );
  NOR2_X1 U405 ( .A1(n574), .A2(n576), .ZN(n349) );
  XOR2_X1 U406 ( .A(G176GAT), .B(G64GAT), .Z(n398) );
  XOR2_X1 U407 ( .A(G92GAT), .B(G78GAT), .Z(n351) );
  XNOR2_X1 U408 ( .A(G120GAT), .B(G148GAT), .ZN(n350) );
  XNOR2_X1 U409 ( .A(n351), .B(n350), .ZN(n352) );
  XOR2_X1 U410 ( .A(n398), .B(n352), .Z(n354) );
  NAND2_X1 U411 ( .A1(G230GAT), .A2(G233GAT), .ZN(n353) );
  XNOR2_X1 U412 ( .A(n354), .B(n353), .ZN(n366) );
  XOR2_X1 U413 ( .A(KEYINPUT80), .B(KEYINPUT32), .Z(n356) );
  XNOR2_X1 U414 ( .A(KEYINPUT31), .B(KEYINPUT79), .ZN(n355) );
  XNOR2_X1 U415 ( .A(n356), .B(n355), .ZN(n360) );
  XOR2_X1 U416 ( .A(KEYINPUT76), .B(KEYINPUT33), .Z(n358) );
  XNOR2_X1 U417 ( .A(G204GAT), .B(KEYINPUT77), .ZN(n357) );
  XNOR2_X1 U418 ( .A(n358), .B(n357), .ZN(n359) );
  XOR2_X1 U419 ( .A(n360), .B(n359), .Z(n364) );
  XNOR2_X1 U420 ( .A(n362), .B(n361), .ZN(n363) );
  XNOR2_X1 U421 ( .A(n364), .B(n363), .ZN(n365) );
  XOR2_X1 U422 ( .A(n366), .B(n365), .Z(n456) );
  INV_X1 U423 ( .A(n456), .ZN(n571) );
  NAND2_X1 U424 ( .A1(n367), .A2(n571), .ZN(n368) );
  XNOR2_X1 U425 ( .A(KEYINPUT117), .B(n368), .ZN(n387) );
  XOR2_X1 U426 ( .A(KEYINPUT71), .B(KEYINPUT67), .Z(n370) );
  XNOR2_X1 U427 ( .A(G169GAT), .B(G197GAT), .ZN(n369) );
  XNOR2_X1 U428 ( .A(n370), .B(n369), .ZN(n374) );
  XOR2_X1 U429 ( .A(KEYINPUT68), .B(KEYINPUT66), .Z(n372) );
  XNOR2_X1 U430 ( .A(KEYINPUT70), .B(KEYINPUT30), .ZN(n371) );
  XNOR2_X1 U431 ( .A(n372), .B(n371), .ZN(n373) );
  XOR2_X1 U432 ( .A(n374), .B(n373), .Z(n381) );
  XOR2_X1 U433 ( .A(G141GAT), .B(G22GAT), .Z(n427) );
  XOR2_X1 U434 ( .A(n375), .B(n427), .Z(n377) );
  XNOR2_X1 U435 ( .A(G36GAT), .B(G113GAT), .ZN(n376) );
  XNOR2_X1 U436 ( .A(n377), .B(n376), .ZN(n378) );
  XNOR2_X1 U437 ( .A(n379), .B(n378), .ZN(n380) );
  XNOR2_X1 U438 ( .A(n381), .B(n380), .ZN(n386) );
  XOR2_X1 U439 ( .A(KEYINPUT29), .B(G8GAT), .Z(n383) );
  NAND2_X1 U440 ( .A1(G229GAT), .A2(G233GAT), .ZN(n382) );
  XNOR2_X1 U441 ( .A(n383), .B(n382), .ZN(n384) );
  XOR2_X1 U442 ( .A(KEYINPUT69), .B(n384), .Z(n385) );
  XNOR2_X1 U443 ( .A(n386), .B(n385), .ZN(n566) );
  XNOR2_X1 U444 ( .A(KEYINPUT74), .B(n566), .ZN(n552) );
  NAND2_X1 U445 ( .A1(n387), .A2(n552), .ZN(n394) );
  XNOR2_X1 U446 ( .A(n456), .B(KEYINPUT41), .ZN(n554) );
  NOR2_X1 U447 ( .A1(n566), .A2(n554), .ZN(n389) );
  XNOR2_X1 U448 ( .A(KEYINPUT116), .B(KEYINPUT46), .ZN(n388) );
  XNOR2_X1 U449 ( .A(n389), .B(n388), .ZN(n391) );
  XNOR2_X1 U450 ( .A(n546), .B(KEYINPUT115), .ZN(n561) );
  NAND2_X1 U451 ( .A1(n550), .A2(n561), .ZN(n390) );
  NOR2_X1 U452 ( .A1(n391), .A2(n390), .ZN(n392) );
  XNOR2_X1 U453 ( .A(KEYINPUT47), .B(n392), .ZN(n393) );
  NAND2_X1 U454 ( .A1(n394), .A2(n393), .ZN(n395) );
  XOR2_X1 U455 ( .A(n395), .B(KEYINPUT48), .Z(n524) );
  INV_X1 U456 ( .A(n524), .ZN(n413) );
  XOR2_X1 U457 ( .A(KEYINPUT103), .B(KEYINPUT101), .Z(n397) );
  XNOR2_X1 U458 ( .A(KEYINPUT100), .B(KEYINPUT102), .ZN(n396) );
  XNOR2_X1 U459 ( .A(n397), .B(n396), .ZN(n411) );
  XOR2_X1 U460 ( .A(n399), .B(n398), .Z(n401) );
  NAND2_X1 U461 ( .A1(G226GAT), .A2(G233GAT), .ZN(n400) );
  XNOR2_X1 U462 ( .A(n401), .B(n400), .ZN(n403) );
  XOR2_X1 U463 ( .A(KEYINPUT17), .B(KEYINPUT19), .Z(n405) );
  XNOR2_X1 U464 ( .A(KEYINPUT18), .B(KEYINPUT92), .ZN(n404) );
  XNOR2_X1 U465 ( .A(n405), .B(n404), .ZN(n406) );
  XOR2_X1 U466 ( .A(G169GAT), .B(n406), .Z(n446) );
  XOR2_X1 U467 ( .A(G204GAT), .B(KEYINPUT95), .Z(n408) );
  XNOR2_X1 U468 ( .A(G197GAT), .B(KEYINPUT21), .ZN(n407) );
  XNOR2_X1 U469 ( .A(n408), .B(n407), .ZN(n422) );
  XNOR2_X1 U470 ( .A(n446), .B(n422), .ZN(n409) );
  XNOR2_X1 U471 ( .A(n290), .B(n409), .ZN(n410) );
  XOR2_X2 U472 ( .A(n411), .B(n410), .Z(n516) );
  XOR2_X1 U473 ( .A(KEYINPUT121), .B(n516), .Z(n412) );
  NAND2_X1 U474 ( .A1(n413), .A2(n412), .ZN(n415) );
  XNOR2_X1 U475 ( .A(KEYINPUT122), .B(KEYINPUT54), .ZN(n414) );
  XNOR2_X1 U476 ( .A(n415), .B(n414), .ZN(n416) );
  NOR2_X1 U477 ( .A1(n514), .A2(n416), .ZN(n564) );
  XOR2_X1 U478 ( .A(KEYINPUT24), .B(G211GAT), .Z(n418) );
  XNOR2_X1 U479 ( .A(KEYINPUT98), .B(KEYINPUT23), .ZN(n417) );
  XNOR2_X1 U480 ( .A(n418), .B(n417), .ZN(n435) );
  XOR2_X1 U481 ( .A(KEYINPUT94), .B(KEYINPUT97), .Z(n420) );
  NAND2_X1 U482 ( .A1(G228GAT), .A2(G233GAT), .ZN(n419) );
  XNOR2_X1 U483 ( .A(n420), .B(n419), .ZN(n421) );
  XOR2_X1 U484 ( .A(n421), .B(KEYINPUT22), .Z(n425) );
  XNOR2_X1 U485 ( .A(n423), .B(n422), .ZN(n424) );
  XNOR2_X1 U486 ( .A(n425), .B(n424), .ZN(n431) );
  XOR2_X1 U487 ( .A(G162GAT), .B(G218GAT), .Z(n429) );
  XNOR2_X1 U488 ( .A(n427), .B(n426), .ZN(n428) );
  XNOR2_X1 U489 ( .A(n429), .B(n428), .ZN(n430) );
  XOR2_X1 U490 ( .A(n431), .B(n430), .Z(n433) );
  XNOR2_X1 U491 ( .A(G50GAT), .B(G106GAT), .ZN(n432) );
  XNOR2_X1 U492 ( .A(n433), .B(n432), .ZN(n434) );
  XNOR2_X1 U493 ( .A(n435), .B(n434), .ZN(n472) );
  NAND2_X1 U494 ( .A1(n564), .A2(n472), .ZN(n436) );
  XNOR2_X1 U495 ( .A(KEYINPUT55), .B(n436), .ZN(n452) );
  XNOR2_X1 U496 ( .A(G43GAT), .B(G134GAT), .ZN(n437) );
  XNOR2_X1 U497 ( .A(n292), .B(n437), .ZN(n438) );
  NAND2_X1 U498 ( .A1(G227GAT), .A2(G233GAT), .ZN(n439) );
  XNOR2_X1 U499 ( .A(n291), .B(n439), .ZN(n449) );
  XOR2_X1 U500 ( .A(KEYINPUT93), .B(G176GAT), .Z(n441) );
  XNOR2_X1 U501 ( .A(KEYINPUT90), .B(KEYINPUT89), .ZN(n440) );
  XNOR2_X1 U502 ( .A(n441), .B(n440), .ZN(n445) );
  XOR2_X1 U503 ( .A(G183GAT), .B(KEYINPUT20), .Z(n443) );
  XNOR2_X1 U504 ( .A(G15GAT), .B(KEYINPUT91), .ZN(n442) );
  XNOR2_X1 U505 ( .A(n443), .B(n442), .ZN(n444) );
  XOR2_X1 U506 ( .A(n445), .B(n444), .Z(n447) );
  XNOR2_X1 U507 ( .A(n451), .B(n450), .ZN(n525) );
  NAND2_X1 U508 ( .A1(n452), .A2(n525), .ZN(n560) );
  NOR2_X1 U509 ( .A1(n534), .A2(n560), .ZN(n455) );
  XNOR2_X1 U510 ( .A(KEYINPUT58), .B(KEYINPUT125), .ZN(n453) );
  NOR2_X1 U511 ( .A1(n552), .A2(n456), .ZN(n492) );
  INV_X1 U512 ( .A(n492), .ZN(n478) );
  NAND2_X1 U513 ( .A1(n546), .A2(n534), .ZN(n457) );
  XNOR2_X1 U514 ( .A(n457), .B(KEYINPUT87), .ZN(n458) );
  XNOR2_X1 U515 ( .A(n458), .B(KEYINPUT16), .ZN(n477) );
  XOR2_X1 U516 ( .A(KEYINPUT106), .B(n459), .Z(n460) );
  NAND2_X1 U517 ( .A1(n472), .A2(n460), .ZN(n461) );
  XNOR2_X1 U518 ( .A(n462), .B(KEYINPUT107), .ZN(n467) );
  NOR2_X1 U519 ( .A1(n525), .A2(n472), .ZN(n464) );
  XNOR2_X1 U520 ( .A(KEYINPUT105), .B(KEYINPUT26), .ZN(n463) );
  XNOR2_X1 U521 ( .A(n464), .B(n463), .ZN(n465) );
  XOR2_X1 U522 ( .A(KEYINPUT104), .B(n465), .Z(n563) );
  XNOR2_X1 U523 ( .A(KEYINPUT27), .B(n516), .ZN(n473) );
  NAND2_X1 U524 ( .A1(n563), .A2(n473), .ZN(n466) );
  NAND2_X1 U525 ( .A1(n467), .A2(n466), .ZN(n468) );
  XOR2_X1 U526 ( .A(KEYINPUT108), .B(n468), .Z(n469) );
  XNOR2_X1 U527 ( .A(KEYINPUT109), .B(n470), .ZN(n476) );
  XOR2_X1 U528 ( .A(KEYINPUT65), .B(KEYINPUT28), .Z(n471) );
  XNOR2_X1 U529 ( .A(n472), .B(n471), .ZN(n527) );
  NAND2_X1 U530 ( .A1(n514), .A2(n473), .ZN(n523) );
  NOR2_X1 U531 ( .A1(n523), .A2(n525), .ZN(n474) );
  NAND2_X1 U532 ( .A1(n527), .A2(n474), .ZN(n475) );
  NAND2_X1 U533 ( .A1(n476), .A2(n475), .ZN(n489) );
  NAND2_X1 U534 ( .A1(n477), .A2(n489), .ZN(n501) );
  NOR2_X1 U535 ( .A1(n478), .A2(n501), .ZN(n486) );
  NAND2_X1 U536 ( .A1(n514), .A2(n486), .ZN(n479) );
  XNOR2_X1 U537 ( .A(n479), .B(KEYINPUT34), .ZN(n480) );
  XNOR2_X1 U538 ( .A(G1GAT), .B(n480), .ZN(G1324GAT) );
  NAND2_X1 U539 ( .A1(n486), .A2(n516), .ZN(n481) );
  XNOR2_X1 U540 ( .A(n481), .B(G8GAT), .ZN(G1325GAT) );
  XOR2_X1 U541 ( .A(KEYINPUT35), .B(KEYINPUT111), .Z(n483) );
  NAND2_X1 U542 ( .A1(n486), .A2(n525), .ZN(n482) );
  XNOR2_X1 U543 ( .A(n483), .B(n482), .ZN(n485) );
  XOR2_X1 U544 ( .A(G15GAT), .B(KEYINPUT110), .Z(n484) );
  XNOR2_X1 U545 ( .A(n485), .B(n484), .ZN(G1326GAT) );
  INV_X1 U546 ( .A(n527), .ZN(n520) );
  NAND2_X1 U547 ( .A1(n520), .A2(n486), .ZN(n487) );
  XNOR2_X1 U548 ( .A(n487), .B(KEYINPUT112), .ZN(n488) );
  XNOR2_X1 U549 ( .A(G22GAT), .B(n488), .ZN(G1327GAT) );
  XOR2_X1 U550 ( .A(G29GAT), .B(KEYINPUT39), .Z(n495) );
  NOR2_X1 U551 ( .A1(n546), .A2(n576), .ZN(n490) );
  NAND2_X1 U552 ( .A1(n490), .A2(n489), .ZN(n491) );
  XNOR2_X1 U553 ( .A(KEYINPUT37), .B(n491), .ZN(n513) );
  NAND2_X1 U554 ( .A1(n513), .A2(n492), .ZN(n493) );
  NAND2_X1 U555 ( .A1(n499), .A2(n514), .ZN(n494) );
  XNOR2_X1 U556 ( .A(n495), .B(n494), .ZN(G1328GAT) );
  NAND2_X1 U557 ( .A1(n499), .A2(n516), .ZN(n496) );
  XNOR2_X1 U558 ( .A(n496), .B(G36GAT), .ZN(G1329GAT) );
  NAND2_X1 U559 ( .A1(n499), .A2(n525), .ZN(n497) );
  XNOR2_X1 U560 ( .A(n497), .B(KEYINPUT40), .ZN(n498) );
  XNOR2_X1 U561 ( .A(n498), .B(G43GAT), .ZN(G1330GAT) );
  NAND2_X1 U562 ( .A1(n520), .A2(n499), .ZN(n500) );
  XNOR2_X1 U563 ( .A(G50GAT), .B(n500), .ZN(G1331GAT) );
  INV_X1 U564 ( .A(n566), .ZN(n541) );
  NOR2_X1 U565 ( .A1(n541), .A2(n554), .ZN(n512) );
  INV_X1 U566 ( .A(n512), .ZN(n502) );
  NOR2_X1 U567 ( .A1(n502), .A2(n501), .ZN(n507) );
  NAND2_X1 U568 ( .A1(n507), .A2(n514), .ZN(n503) );
  XNOR2_X1 U569 ( .A(KEYINPUT42), .B(n503), .ZN(n504) );
  XNOR2_X1 U570 ( .A(G57GAT), .B(n504), .ZN(G1332GAT) );
  NAND2_X1 U571 ( .A1(n507), .A2(n516), .ZN(n505) );
  XNOR2_X1 U572 ( .A(n505), .B(G64GAT), .ZN(G1333GAT) );
  NAND2_X1 U573 ( .A1(n507), .A2(n525), .ZN(n506) );
  XNOR2_X1 U574 ( .A(n506), .B(G71GAT), .ZN(G1334GAT) );
  XOR2_X1 U575 ( .A(KEYINPUT113), .B(KEYINPUT43), .Z(n509) );
  NAND2_X1 U576 ( .A1(n507), .A2(n520), .ZN(n508) );
  XNOR2_X1 U577 ( .A(n509), .B(n508), .ZN(n511) );
  XOR2_X1 U578 ( .A(G78GAT), .B(KEYINPUT114), .Z(n510) );
  XNOR2_X1 U579 ( .A(n511), .B(n510), .ZN(G1335GAT) );
  AND2_X1 U580 ( .A1(n513), .A2(n512), .ZN(n519) );
  NAND2_X1 U581 ( .A1(n519), .A2(n514), .ZN(n515) );
  XNOR2_X1 U582 ( .A(G85GAT), .B(n515), .ZN(G1336GAT) );
  NAND2_X1 U583 ( .A1(n519), .A2(n516), .ZN(n517) );
  XNOR2_X1 U584 ( .A(n517), .B(G92GAT), .ZN(G1337GAT) );
  NAND2_X1 U585 ( .A1(n519), .A2(n525), .ZN(n518) );
  XNOR2_X1 U586 ( .A(n518), .B(G99GAT), .ZN(G1338GAT) );
  NAND2_X1 U587 ( .A1(n520), .A2(n519), .ZN(n521) );
  XNOR2_X1 U588 ( .A(n521), .B(KEYINPUT44), .ZN(n522) );
  XNOR2_X1 U589 ( .A(G106GAT), .B(n522), .ZN(G1339GAT) );
  NOR2_X1 U590 ( .A1(n524), .A2(n523), .ZN(n540) );
  AND2_X1 U591 ( .A1(n525), .A2(n540), .ZN(n526) );
  XNOR2_X1 U592 ( .A(KEYINPUT118), .B(n526), .ZN(n528) );
  NAND2_X1 U593 ( .A1(n528), .A2(n527), .ZN(n535) );
  NOR2_X1 U594 ( .A1(n552), .A2(n535), .ZN(n529) );
  XOR2_X1 U595 ( .A(G113GAT), .B(n529), .Z(G1340GAT) );
  NOR2_X1 U596 ( .A1(n554), .A2(n535), .ZN(n531) );
  XNOR2_X1 U597 ( .A(G120GAT), .B(KEYINPUT49), .ZN(n530) );
  XNOR2_X1 U598 ( .A(n531), .B(n530), .ZN(G1341GAT) );
  NOR2_X1 U599 ( .A1(n561), .A2(n535), .ZN(n532) );
  XOR2_X1 U600 ( .A(KEYINPUT50), .B(n532), .Z(n533) );
  XNOR2_X1 U601 ( .A(G127GAT), .B(n533), .ZN(G1342GAT) );
  NOR2_X1 U602 ( .A1(n535), .A2(n534), .ZN(n539) );
  XOR2_X1 U603 ( .A(KEYINPUT119), .B(KEYINPUT51), .Z(n537) );
  XNOR2_X1 U604 ( .A(G134GAT), .B(KEYINPUT120), .ZN(n536) );
  XNOR2_X1 U605 ( .A(n537), .B(n536), .ZN(n538) );
  XNOR2_X1 U606 ( .A(n539), .B(n538), .ZN(G1343GAT) );
  NAND2_X1 U607 ( .A1(n563), .A2(n540), .ZN(n549) );
  INV_X1 U608 ( .A(n549), .ZN(n547) );
  NAND2_X1 U609 ( .A1(n541), .A2(n547), .ZN(n542) );
  XNOR2_X1 U610 ( .A(G141GAT), .B(n542), .ZN(G1344GAT) );
  XOR2_X1 U611 ( .A(KEYINPUT53), .B(KEYINPUT52), .Z(n544) );
  OR2_X1 U612 ( .A1(n549), .A2(n554), .ZN(n543) );
  XNOR2_X1 U613 ( .A(n544), .B(n543), .ZN(n545) );
  XNOR2_X1 U614 ( .A(G148GAT), .B(n545), .ZN(G1345GAT) );
  NAND2_X1 U615 ( .A1(n547), .A2(n546), .ZN(n548) );
  XNOR2_X1 U616 ( .A(n548), .B(G155GAT), .ZN(G1346GAT) );
  NOR2_X1 U617 ( .A1(n550), .A2(n549), .ZN(n551) );
  XOR2_X1 U618 ( .A(G162GAT), .B(n551), .Z(G1347GAT) );
  NOR2_X1 U619 ( .A1(n552), .A2(n560), .ZN(n553) );
  XOR2_X1 U620 ( .A(G169GAT), .B(n553), .Z(G1348GAT) );
  NOR2_X1 U621 ( .A1(n554), .A2(n560), .ZN(n559) );
  XOR2_X1 U622 ( .A(KEYINPUT57), .B(KEYINPUT124), .Z(n556) );
  XNOR2_X1 U623 ( .A(G176GAT), .B(KEYINPUT56), .ZN(n555) );
  XNOR2_X1 U624 ( .A(n556), .B(n555), .ZN(n557) );
  XNOR2_X1 U625 ( .A(KEYINPUT123), .B(n557), .ZN(n558) );
  XNOR2_X1 U626 ( .A(n559), .B(n558), .ZN(G1349GAT) );
  NOR2_X1 U627 ( .A1(n561), .A2(n560), .ZN(n562) );
  XOR2_X1 U628 ( .A(G183GAT), .B(n562), .Z(G1350GAT) );
  NAND2_X1 U629 ( .A1(n564), .A2(n563), .ZN(n565) );
  XNOR2_X1 U630 ( .A(KEYINPUT126), .B(n565), .ZN(n577) );
  NOR2_X1 U631 ( .A1(n566), .A2(n577), .ZN(n570) );
  XOR2_X1 U632 ( .A(KEYINPUT127), .B(KEYINPUT60), .Z(n568) );
  XNOR2_X1 U633 ( .A(G197GAT), .B(KEYINPUT59), .ZN(n567) );
  XNOR2_X1 U634 ( .A(n568), .B(n567), .ZN(n569) );
  XNOR2_X1 U635 ( .A(n570), .B(n569), .ZN(G1352GAT) );
  NOR2_X1 U636 ( .A1(n577), .A2(n571), .ZN(n573) );
  XNOR2_X1 U637 ( .A(G204GAT), .B(KEYINPUT61), .ZN(n572) );
  XNOR2_X1 U638 ( .A(n573), .B(n572), .ZN(G1353GAT) );
  NOR2_X1 U639 ( .A1(n577), .A2(n574), .ZN(n575) );
  XOR2_X1 U640 ( .A(G211GAT), .B(n575), .Z(G1354GAT) );
  NOR2_X1 U641 ( .A1(n577), .A2(n576), .ZN(n578) );
  XOR2_X1 U642 ( .A(KEYINPUT62), .B(n578), .Z(n579) );
  XNOR2_X1 U643 ( .A(G218GAT), .B(n579), .ZN(G1355GAT) );
endmodule

