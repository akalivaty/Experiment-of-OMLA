

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355,
         n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
         n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
         n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
         n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
         n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410,
         n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421,
         n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432,
         n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443,
         n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454,
         n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465,
         n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
         n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487,
         n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
         n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
         n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586,
         n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597,
         n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608,
         n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619,
         n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630,
         n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641,
         n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652,
         n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663,
         n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674,
         n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685,
         n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696,
         n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707,
         n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718,
         n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729,
         n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, n740,
         n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, n751,
         n752, n753, n754, n755, n756, n757, n758, n759;

  OR2_X1 U367 ( .A1(n637), .A2(n393), .ZN(n649) );
  XNOR2_X1 U368 ( .A(n462), .B(n730), .ZN(n493) );
  XOR2_X1 U369 ( .A(KEYINPUT88), .B(KEYINPUT90), .Z(n345) );
  XOR2_X1 U370 ( .A(n463), .B(n462), .Z(n346) );
  NAND2_X2 U371 ( .A1(n361), .A2(n355), .ZN(n365) );
  NOR2_X2 U372 ( .A1(n571), .A2(n570), .ZN(n572) );
  XNOR2_X2 U373 ( .A(n587), .B(n586), .ZN(n670) );
  XNOR2_X2 U374 ( .A(G101), .B(KEYINPUT66), .ZN(n448) );
  NAND2_X1 U375 ( .A1(n599), .A2(n563), .ZN(n393) );
  NOR2_X1 U376 ( .A1(n750), .A2(n611), .ZN(n616) );
  OR2_X2 U377 ( .A1(n427), .A2(n429), .ZN(n750) );
  NAND2_X1 U378 ( .A1(n405), .A2(n401), .ZN(n562) );
  AND2_X1 U379 ( .A1(n408), .A2(n406), .ZN(n405) );
  NAND2_X1 U380 ( .A1(n373), .A2(n372), .ZN(n703) );
  XNOR2_X1 U381 ( .A(n376), .B(n357), .ZN(n424) );
  NOR2_X1 U382 ( .A1(n542), .A2(n416), .ZN(n415) );
  NOR2_X1 U383 ( .A1(n541), .A2(n546), .ZN(n384) );
  XNOR2_X1 U384 ( .A(n465), .B(n464), .ZN(n552) );
  XNOR2_X1 U385 ( .A(n505), .B(n504), .ZN(n542) );
  XNOR2_X1 U386 ( .A(n444), .B(n442), .ZN(n546) );
  XNOR2_X1 U387 ( .A(n523), .B(n522), .ZN(n541) );
  XNOR2_X1 U388 ( .A(n454), .B(G472), .ZN(n648) );
  XNOR2_X1 U389 ( .A(n366), .B(n346), .ZN(n714) );
  OR2_X1 U390 ( .A1(n718), .A2(G902), .ZN(n444) );
  XNOR2_X1 U391 ( .A(n685), .B(n684), .ZN(n686) );
  XNOR2_X1 U392 ( .A(n411), .B(n524), .ZN(n729) );
  BUF_X1 U393 ( .A(n602), .Z(n347) );
  NAND2_X1 U394 ( .A1(n436), .A2(n380), .ZN(n602) );
  AND2_X2 U395 ( .A1(n417), .A2(n368), .ZN(n721) );
  XNOR2_X2 U396 ( .A(n448), .B(n414), .ZN(n462) );
  XNOR2_X2 U397 ( .A(n744), .B(G146), .ZN(n366) );
  XNOR2_X2 U398 ( .A(n526), .B(n514), .ZN(n744) );
  XNOR2_X2 U399 ( .A(n617), .B(KEYINPUT75), .ZN(n635) );
  XNOR2_X1 U400 ( .A(n384), .B(KEYINPUT102), .ZN(n660) );
  XNOR2_X1 U401 ( .A(n433), .B(G122), .ZN(n524) );
  INV_X1 U402 ( .A(G107), .ZN(n433) );
  INV_X1 U403 ( .A(n491), .ZN(n404) );
  NAND2_X1 U404 ( .A1(n626), .A2(n521), .ZN(n454) );
  OR2_X1 U405 ( .A1(n701), .A2(n369), .ZN(n378) );
  XNOR2_X1 U406 ( .A(n371), .B(n370), .ZN(n369) );
  NOR2_X1 U407 ( .A1(n658), .A2(n703), .ZN(n371) );
  AND2_X1 U408 ( .A1(n581), .A2(n580), .ZN(n582) );
  INV_X1 U409 ( .A(G237), .ZN(n455) );
  XNOR2_X1 U410 ( .A(KEYINPUT68), .B(G131), .ZN(n514) );
  XNOR2_X1 U411 ( .A(G902), .B(KEYINPUT15), .ZN(n613) );
  XNOR2_X1 U412 ( .A(n649), .B(KEYINPUT107), .ZN(n585) );
  AND2_X1 U413 ( .A1(n660), .A2(n657), .ZN(n655) );
  XNOR2_X1 U414 ( .A(n552), .B(KEYINPUT1), .ZN(n637) );
  XNOR2_X1 U415 ( .A(G122), .B(G140), .ZN(n516) );
  XNOR2_X1 U416 ( .A(n508), .B(n507), .ZN(n510) );
  XNOR2_X1 U417 ( .A(G143), .B(KEYINPUT11), .ZN(n507) );
  XOR2_X1 U418 ( .A(KEYINPUT12), .B(KEYINPUT98), .Z(n508) );
  INV_X1 U419 ( .A(KEYINPUT10), .ZN(n474) );
  XNOR2_X1 U420 ( .A(G104), .B(G107), .ZN(n457) );
  XNOR2_X1 U421 ( .A(KEYINPUT17), .B(KEYINPUT18), .ZN(n497) );
  XNOR2_X1 U422 ( .A(G110), .B(KEYINPUT16), .ZN(n412) );
  XNOR2_X1 U423 ( .A(n750), .B(n359), .ZN(n610) );
  INV_X1 U424 ( .A(KEYINPUT74), .ZN(n359) );
  NAND2_X1 U425 ( .A1(n404), .A2(n402), .ZN(n401) );
  XNOR2_X1 U426 ( .A(KEYINPUT71), .B(KEYINPUT34), .ZN(n589) );
  NOR2_X1 U427 ( .A1(n646), .A2(n548), .ZN(n540) );
  XNOR2_X1 U428 ( .A(n443), .B(G478), .ZN(n442) );
  INV_X1 U429 ( .A(KEYINPUT101), .ZN(n443) );
  NOR2_X1 U430 ( .A1(n438), .A2(n437), .ZN(n436) );
  AND2_X1 U431 ( .A1(n588), .A2(n356), .ZN(n435) );
  BUF_X1 U432 ( .A(n637), .Z(n387) );
  INV_X1 U433 ( .A(KEYINPUT79), .ZN(n633) );
  INV_X1 U434 ( .A(n424), .ZN(n423) );
  NOR2_X1 U435 ( .A1(n400), .A2(n399), .ZN(n398) );
  AND2_X1 U436 ( .A1(n759), .A2(KEYINPUT46), .ZN(n400) );
  INV_X1 U437 ( .A(n680), .ZN(n399) );
  INV_X1 U438 ( .A(G902), .ZN(n521) );
  XNOR2_X1 U439 ( .A(G137), .B(G113), .ZN(n449) );
  XOR2_X1 U440 ( .A(KEYINPUT5), .B(KEYINPUT94), .Z(n450) );
  OR2_X1 U441 ( .A1(n603), .A2(n604), .ZN(n374) );
  NOR2_X1 U442 ( .A1(G953), .A2(G237), .ZN(n513) );
  NAND2_X1 U443 ( .A1(G234), .A2(G237), .ZN(n485) );
  NOR2_X1 U444 ( .A1(n492), .A2(n410), .ZN(n409) );
  NOR2_X1 U445 ( .A1(n538), .A2(n599), .ZN(n539) );
  XNOR2_X1 U446 ( .A(n564), .B(KEYINPUT103), .ZN(n573) );
  NOR2_X1 U447 ( .A1(n573), .A2(n356), .ZN(n438) );
  NAND2_X1 U448 ( .A1(n428), .A2(n352), .ZN(n427) );
  XNOR2_X1 U449 ( .A(n512), .B(n475), .ZN(n746) );
  AND2_X1 U450 ( .A1(n615), .A2(n614), .ZN(n417) );
  NAND2_X1 U451 ( .A1(n585), .A2(n584), .ZN(n587) );
  INV_X1 U452 ( .A(n583), .ZN(n584) );
  NOR2_X1 U453 ( .A1(n734), .A2(KEYINPUT2), .ZN(n630) );
  XNOR2_X1 U454 ( .A(n537), .B(n386), .ZN(n672) );
  INV_X1 U455 ( .A(KEYINPUT41), .ZN(n386) );
  BUF_X1 U456 ( .A(n542), .Z(n560) );
  XNOR2_X1 U457 ( .A(n431), .B(KEYINPUT76), .ZN(n491) );
  NAND2_X1 U458 ( .A1(n432), .A2(n490), .ZN(n431) );
  XNOR2_X1 U459 ( .A(n578), .B(KEYINPUT109), .ZN(n432) );
  NAND2_X1 U460 ( .A1(n391), .A2(n392), .ZN(n578) );
  INV_X1 U461 ( .A(n393), .ZN(n391) );
  BUF_X1 U462 ( .A(n648), .Z(n385) );
  INV_X2 U463 ( .A(G953), .ZN(n752) );
  XOR2_X1 U464 ( .A(G116), .B(KEYINPUT9), .Z(n530) );
  XNOR2_X1 U465 ( .A(n520), .B(n519), .ZN(n685) );
  XNOR2_X1 U466 ( .A(n502), .B(n501), .ZN(n620) );
  XNOR2_X1 U467 ( .A(n729), .B(n493), .ZN(n502) );
  AND2_X1 U468 ( .A1(n615), .A2(n367), .ZN(n419) );
  AND2_X1 U469 ( .A1(G210), .A2(n614), .ZN(n367) );
  XNOR2_X1 U470 ( .A(n360), .B(KEYINPUT42), .ZN(n759) );
  NOR2_X1 U471 ( .A1(n672), .A2(n545), .ZN(n360) );
  INV_X1 U472 ( .A(KEYINPUT40), .ZN(n535) );
  INV_X1 U473 ( .A(n545), .ZN(n373) );
  XNOR2_X1 U474 ( .A(n379), .B(KEYINPUT105), .ZN(n683) );
  AND2_X1 U475 ( .A1(n575), .A2(n583), .ZN(n434) );
  AND2_X1 U476 ( .A1(n440), .A2(n439), .ZN(n677) );
  INV_X1 U477 ( .A(G122), .ZN(n681) );
  AND2_X1 U478 ( .A1(G475), .A2(n614), .ZN(n348) );
  INV_X1 U479 ( .A(G146), .ZN(n447) );
  OR2_X1 U480 ( .A1(n491), .A2(n492), .ZN(n349) );
  NAND2_X1 U481 ( .A1(n603), .A2(n604), .ZN(n350) );
  OR2_X1 U482 ( .A1(n678), .A2(KEYINPUT81), .ZN(n351) );
  AND2_X1 U483 ( .A1(n711), .A2(n351), .ZN(n352) );
  AND2_X1 U484 ( .A1(n398), .A2(n394), .ZN(n353) );
  AND2_X1 U485 ( .A1(n678), .A2(KEYINPUT81), .ZN(n354) );
  AND2_X1 U486 ( .A1(n608), .A2(n374), .ZN(n355) );
  XOR2_X1 U487 ( .A(n574), .B(KEYINPUT22), .Z(n356) );
  XOR2_X1 U488 ( .A(n577), .B(KEYINPUT96), .Z(n357) );
  XNOR2_X1 U489 ( .A(n560), .B(KEYINPUT38), .ZN(n657) );
  INV_X1 U490 ( .A(n657), .ZN(n410) );
  XNOR2_X1 U491 ( .A(KEYINPUT62), .B(n626), .ZN(n358) );
  INV_X1 U492 ( .A(n656), .ZN(n416) );
  AND2_X1 U493 ( .A1(n750), .A2(n611), .ZN(n631) );
  NAND2_X1 U494 ( .A1(n363), .A2(n362), .ZN(n361) );
  NAND2_X1 U495 ( .A1(n375), .A2(n350), .ZN(n362) );
  NAND2_X1 U496 ( .A1(n364), .A2(n604), .ZN(n363) );
  INV_X1 U497 ( .A(n375), .ZN(n364) );
  XNOR2_X2 U498 ( .A(n365), .B(n609), .ZN(n734) );
  XNOR2_X1 U499 ( .A(n366), .B(n453), .ZN(n626) );
  AND2_X1 U500 ( .A1(n615), .A2(n348), .ZN(n420) );
  INV_X2 U501 ( .A(n635), .ZN(n368) );
  INV_X1 U502 ( .A(KEYINPUT47), .ZN(n370) );
  INV_X1 U503 ( .A(n571), .ZN(n372) );
  XNOR2_X1 U504 ( .A(n382), .B(KEYINPUT85), .ZN(n375) );
  XNOR2_X1 U505 ( .A(n593), .B(KEYINPUT35), .ZN(n682) );
  XNOR2_X1 U506 ( .A(n383), .B(KEYINPUT106), .ZN(n595) );
  XNOR2_X1 U507 ( .A(n415), .B(KEYINPUT19), .ZN(n571) );
  AND2_X1 U508 ( .A1(n588), .A2(n576), .ZN(n376) );
  XNOR2_X1 U509 ( .A(n511), .B(n512), .ZN(n520) );
  NAND2_X1 U510 ( .A1(n377), .A2(n392), .ZN(n545) );
  XNOR2_X1 U511 ( .A(n540), .B(KEYINPUT28), .ZN(n377) );
  XNOR2_X1 U512 ( .A(n378), .B(KEYINPUT73), .ZN(n397) );
  NAND2_X1 U513 ( .A1(n602), .A2(n434), .ZN(n379) );
  NAND2_X1 U514 ( .A1(n430), .A2(n354), .ZN(n428) );
  NOR2_X1 U515 ( .A1(n723), .A2(G902), .ZN(n480) );
  NAND2_X1 U516 ( .A1(n435), .A2(n573), .ZN(n380) );
  NOR2_X2 U517 ( .A1(n624), .A2(n727), .ZN(n625) );
  NOR2_X2 U518 ( .A1(n688), .A2(n727), .ZN(n689) );
  XNOR2_X2 U519 ( .A(G137), .B(G140), .ZN(n475) );
  BUF_X1 U520 ( .A(n682), .Z(n381) );
  XNOR2_X1 U521 ( .A(n461), .B(n460), .ZN(n463) );
  NAND2_X1 U522 ( .A1(n714), .A2(n521), .ZN(n465) );
  NAND2_X1 U523 ( .A1(n594), .A2(n595), .ZN(n382) );
  NOR2_X2 U524 ( .A1(n683), .A2(n582), .ZN(n383) );
  NOR2_X1 U525 ( .A1(n759), .A2(KEYINPUT46), .ZN(n425) );
  NAND2_X1 U526 ( .A1(n388), .A2(n628), .ZN(n629) );
  XNOR2_X1 U527 ( .A(n627), .B(n358), .ZN(n388) );
  XNOR2_X1 U528 ( .A(n389), .B(n746), .ZN(n723) );
  XNOR2_X1 U529 ( .A(n495), .B(n474), .ZN(n512) );
  XNOR2_X1 U530 ( .A(n390), .B(n473), .ZN(n389) );
  XNOR2_X1 U531 ( .A(n469), .B(n470), .ZN(n390) );
  INV_X1 U532 ( .A(n552), .ZN(n392) );
  NAND2_X1 U533 ( .A1(n387), .A2(n393), .ZN(n639) );
  NAND2_X1 U534 ( .A1(n757), .A2(KEYINPUT46), .ZN(n394) );
  NAND2_X1 U535 ( .A1(n395), .A2(n353), .ZN(n555) );
  AND2_X1 U536 ( .A1(n396), .A2(n397), .ZN(n395) );
  NAND2_X1 U537 ( .A1(n426), .A2(n425), .ZN(n396) );
  AND2_X1 U538 ( .A1(n409), .A2(n403), .ZN(n402) );
  INV_X1 U539 ( .A(n506), .ZN(n403) );
  NAND2_X1 U540 ( .A1(n407), .A2(n506), .ZN(n406) );
  INV_X1 U541 ( .A(n409), .ZN(n407) );
  NAND2_X1 U542 ( .A1(n491), .A2(n506), .ZN(n408) );
  NAND2_X1 U543 ( .A1(n562), .A2(n705), .ZN(n536) );
  XNOR2_X1 U544 ( .A(n509), .B(n412), .ZN(n411) );
  XNOR2_X2 U545 ( .A(n413), .B(G119), .ZN(n730) );
  XNOR2_X2 U546 ( .A(G113), .B(G104), .ZN(n509) );
  XNOR2_X2 U547 ( .A(G116), .B(KEYINPUT3), .ZN(n413) );
  INV_X1 U548 ( .A(KEYINPUT4), .ZN(n414) );
  INV_X1 U549 ( .A(n560), .ZN(n544) );
  NAND2_X1 U550 ( .A1(n418), .A2(n417), .ZN(n627) );
  NOR2_X1 U551 ( .A1(n635), .A2(n421), .ZN(n418) );
  NAND2_X1 U552 ( .A1(n419), .A2(n368), .ZN(n622) );
  NAND2_X1 U553 ( .A1(n420), .A2(n368), .ZN(n687) );
  INV_X1 U554 ( .A(G472), .ZN(n421) );
  NAND2_X1 U555 ( .A1(n423), .A2(n422), .ZN(n581) );
  INV_X1 U556 ( .A(n692), .ZN(n422) );
  NAND2_X1 U557 ( .A1(n424), .A2(n707), .ZN(n708) );
  NAND2_X1 U558 ( .A1(n424), .A2(n705), .ZN(n706) );
  XNOR2_X2 U559 ( .A(n498), .B(G134), .ZN(n526) );
  INV_X1 U560 ( .A(n757), .ZN(n426) );
  XNOR2_X2 U561 ( .A(n536), .B(n535), .ZN(n757) );
  NOR2_X1 U562 ( .A1(n430), .A2(KEYINPUT81), .ZN(n429) );
  XNOR2_X1 U563 ( .A(n555), .B(n554), .ZN(n430) );
  AND2_X1 U564 ( .A1(n347), .A2(n583), .ZN(n597) );
  NOR2_X1 U565 ( .A1(n588), .A2(n356), .ZN(n437) );
  NOR2_X1 U566 ( .A1(n675), .A2(G953), .ZN(n439) );
  NAND2_X1 U567 ( .A1(n441), .A2(n368), .ZN(n440) );
  XNOR2_X1 U568 ( .A(n634), .B(n633), .ZN(n441) );
  XNOR2_X1 U569 ( .A(n723), .B(n722), .ZN(n724) );
  XNOR2_X2 U570 ( .A(n480), .B(n479), .ZN(n599) );
  AND2_X1 U571 ( .A1(n513), .A2(G210), .ZN(n445) );
  XOR2_X1 U572 ( .A(KEYINPUT65), .B(KEYINPUT0), .Z(n446) );
  XNOR2_X1 U573 ( .A(n451), .B(n445), .ZN(n452) );
  XNOR2_X1 U574 ( .A(n493), .B(n452), .ZN(n453) );
  XNOR2_X1 U575 ( .A(n475), .B(n459), .ZN(n460) );
  INV_X1 U576 ( .A(n727), .ZN(n628) );
  XNOR2_X1 U577 ( .A(n725), .B(n724), .ZN(n726) );
  XNOR2_X2 U578 ( .A(G143), .B(G128), .ZN(n498) );
  XNOR2_X1 U579 ( .A(n450), .B(n449), .ZN(n451) );
  NAND2_X1 U580 ( .A1(n521), .A2(n455), .ZN(n503) );
  NAND2_X1 U581 ( .A1(n503), .A2(G214), .ZN(n656) );
  NAND2_X1 U582 ( .A1(n648), .A2(n656), .ZN(n456) );
  XNOR2_X1 U583 ( .A(KEYINPUT30), .B(n456), .ZN(n492) );
  XOR2_X1 U584 ( .A(KEYINPUT77), .B(G110), .Z(n458) );
  XNOR2_X1 U585 ( .A(n458), .B(n457), .ZN(n461) );
  NAND2_X1 U586 ( .A1(G227), .A2(n752), .ZN(n459) );
  XNOR2_X1 U587 ( .A(KEYINPUT69), .B(G469), .ZN(n464) );
  XNOR2_X1 U588 ( .A(KEYINPUT89), .B(G110), .ZN(n467) );
  XNOR2_X1 U589 ( .A(G119), .B(G128), .ZN(n466) );
  XNOR2_X1 U590 ( .A(n467), .B(n466), .ZN(n470) );
  XNOR2_X1 U591 ( .A(KEYINPUT24), .B(KEYINPUT23), .ZN(n468) );
  XNOR2_X1 U592 ( .A(n345), .B(n468), .ZN(n469) );
  NAND2_X1 U593 ( .A1(n752), .A2(G234), .ZN(n472) );
  XNOR2_X1 U594 ( .A(KEYINPUT67), .B(KEYINPUT8), .ZN(n471) );
  XNOR2_X1 U595 ( .A(n472), .B(n471), .ZN(n528) );
  NAND2_X1 U596 ( .A1(G221), .A2(n528), .ZN(n473) );
  XNOR2_X1 U597 ( .A(n447), .B(G125), .ZN(n495) );
  XOR2_X1 U598 ( .A(KEYINPUT25), .B(KEYINPUT91), .Z(n478) );
  NAND2_X1 U599 ( .A1(G234), .A2(n613), .ZN(n476) );
  XNOR2_X1 U600 ( .A(KEYINPUT20), .B(n476), .ZN(n481) );
  NAND2_X1 U601 ( .A1(n481), .A2(G217), .ZN(n477) );
  XNOR2_X1 U602 ( .A(n478), .B(n477), .ZN(n479) );
  XOR2_X1 U603 ( .A(KEYINPUT92), .B(KEYINPUT21), .Z(n483) );
  NAND2_X1 U604 ( .A1(n481), .A2(G221), .ZN(n482) );
  XNOR2_X1 U605 ( .A(n483), .B(n482), .ZN(n641) );
  INV_X1 U606 ( .A(KEYINPUT93), .ZN(n484) );
  XNOR2_X1 U607 ( .A(n641), .B(n484), .ZN(n563) );
  XNOR2_X1 U608 ( .A(n485), .B(KEYINPUT14), .ZN(n486) );
  NAND2_X1 U609 ( .A1(G952), .A2(n486), .ZN(n669) );
  NOR2_X1 U610 ( .A1(n669), .A2(G953), .ZN(n569) );
  NAND2_X1 U611 ( .A1(G902), .A2(n486), .ZN(n565) );
  NOR2_X1 U612 ( .A1(G900), .A2(n565), .ZN(n487) );
  NAND2_X1 U613 ( .A1(G953), .A2(n487), .ZN(n488) );
  XOR2_X1 U614 ( .A(KEYINPUT108), .B(n488), .Z(n489) );
  NOR2_X1 U615 ( .A1(n569), .A2(n489), .ZN(n538) );
  INV_X1 U616 ( .A(n538), .ZN(n490) );
  NAND2_X1 U617 ( .A1(n752), .A2(G224), .ZN(n494) );
  XNOR2_X1 U618 ( .A(n494), .B(KEYINPUT78), .ZN(n496) );
  XNOR2_X1 U619 ( .A(n496), .B(n495), .ZN(n500) );
  XNOR2_X1 U620 ( .A(n498), .B(n497), .ZN(n499) );
  XNOR2_X1 U621 ( .A(n500), .B(n499), .ZN(n501) );
  NAND2_X1 U622 ( .A1(n620), .A2(n613), .ZN(n505) );
  NAND2_X1 U623 ( .A1(n503), .A2(G210), .ZN(n504) );
  XOR2_X1 U624 ( .A(KEYINPUT83), .B(KEYINPUT39), .Z(n506) );
  XNOR2_X1 U625 ( .A(n509), .B(n510), .ZN(n511) );
  NAND2_X1 U626 ( .A1(G214), .A2(n513), .ZN(n515) );
  XNOR2_X1 U627 ( .A(n515), .B(n514), .ZN(n518) );
  XNOR2_X1 U628 ( .A(n516), .B(KEYINPUT97), .ZN(n517) );
  XNOR2_X1 U629 ( .A(n518), .B(n517), .ZN(n519) );
  NAND2_X1 U630 ( .A1(n685), .A2(n521), .ZN(n523) );
  XOR2_X1 U631 ( .A(KEYINPUT13), .B(G475), .Z(n522) );
  XNOR2_X1 U632 ( .A(n541), .B(KEYINPUT99), .ZN(n547) );
  INV_X1 U633 ( .A(n547), .ZN(n534) );
  XOR2_X1 U634 ( .A(KEYINPUT7), .B(KEYINPUT100), .Z(n525) );
  XNOR2_X1 U635 ( .A(n525), .B(n524), .ZN(n527) );
  XOR2_X1 U636 ( .A(n526), .B(n527), .Z(n532) );
  NAND2_X1 U637 ( .A1(G217), .A2(n528), .ZN(n529) );
  XNOR2_X1 U638 ( .A(n530), .B(n529), .ZN(n531) );
  XNOR2_X1 U639 ( .A(n532), .B(n531), .ZN(n718) );
  INV_X1 U640 ( .A(n546), .ZN(n533) );
  NAND2_X1 U641 ( .A1(n534), .A2(n533), .ZN(n702) );
  INV_X1 U642 ( .A(n702), .ZN(n705) );
  NAND2_X1 U643 ( .A1(n655), .A2(n656), .ZN(n537) );
  INV_X1 U644 ( .A(n648), .ZN(n646) );
  NAND2_X1 U645 ( .A1(n641), .A2(n539), .ZN(n548) );
  AND2_X1 U646 ( .A1(n546), .A2(n541), .ZN(n591) );
  NAND2_X1 U647 ( .A1(n591), .A2(n544), .ZN(n543) );
  NOR2_X1 U648 ( .A1(n349), .A2(n543), .ZN(n701) );
  AND2_X1 U649 ( .A1(n547), .A2(n546), .ZN(n707) );
  INV_X1 U650 ( .A(n707), .ZN(n697) );
  NAND2_X1 U651 ( .A1(n702), .A2(n697), .ZN(n580) );
  INV_X1 U652 ( .A(n580), .ZN(n658) );
  NOR2_X1 U653 ( .A1(n702), .A2(n548), .ZN(n549) );
  NAND2_X1 U654 ( .A1(n549), .A2(n656), .ZN(n550) );
  XNOR2_X1 U655 ( .A(n648), .B(KEYINPUT6), .ZN(n583) );
  OR2_X1 U656 ( .A1(n550), .A2(n583), .ZN(n557) );
  NOR2_X1 U657 ( .A1(n557), .A2(n560), .ZN(n551) );
  XNOR2_X1 U658 ( .A(n551), .B(KEYINPUT36), .ZN(n553) );
  INV_X1 U659 ( .A(n387), .ZN(n556) );
  NAND2_X1 U660 ( .A1(n553), .A2(n556), .ZN(n680) );
  XOR2_X1 U661 ( .A(KEYINPUT48), .B(KEYINPUT82), .Z(n554) );
  NOR2_X1 U662 ( .A1(n557), .A2(n556), .ZN(n559) );
  INV_X1 U663 ( .A(KEYINPUT43), .ZN(n558) );
  XNOR2_X1 U664 ( .A(n559), .B(n558), .ZN(n561) );
  NAND2_X1 U665 ( .A1(n561), .A2(n560), .ZN(n678) );
  NAND2_X1 U666 ( .A1(n562), .A2(n707), .ZN(n711) );
  NAND2_X1 U667 ( .A1(n660), .A2(n563), .ZN(n564) );
  NOR2_X1 U668 ( .A1(G898), .A2(n752), .ZN(n733) );
  INV_X1 U669 ( .A(n565), .ZN(n566) );
  NAND2_X1 U670 ( .A1(n733), .A2(n566), .ZN(n567) );
  XNOR2_X1 U671 ( .A(n567), .B(KEYINPUT87), .ZN(n568) );
  NOR2_X1 U672 ( .A1(n569), .A2(n568), .ZN(n570) );
  XNOR2_X2 U673 ( .A(n572), .B(n446), .ZN(n588) );
  INV_X1 U674 ( .A(KEYINPUT72), .ZN(n574) );
  XNOR2_X1 U675 ( .A(n599), .B(KEYINPUT104), .ZN(n640) );
  AND2_X1 U676 ( .A1(n387), .A2(n640), .ZN(n575) );
  NOR2_X1 U677 ( .A1(n649), .A2(n646), .ZN(n576) );
  XOR2_X1 U678 ( .A(KEYINPUT31), .B(KEYINPUT95), .Z(n577) );
  NOR2_X1 U679 ( .A1(n385), .A2(n578), .ZN(n579) );
  AND2_X1 U680 ( .A1(n588), .A2(n579), .ZN(n692) );
  XNOR2_X1 U681 ( .A(KEYINPUT70), .B(KEYINPUT33), .ZN(n586) );
  NAND2_X1 U682 ( .A1(n670), .A2(n588), .ZN(n590) );
  XNOR2_X1 U683 ( .A(n590), .B(n589), .ZN(n592) );
  NAND2_X1 U684 ( .A1(n592), .A2(n591), .ZN(n593) );
  NAND2_X1 U685 ( .A1(n682), .A2(KEYINPUT44), .ZN(n594) );
  NOR2_X1 U686 ( .A1(n387), .A2(n640), .ZN(n596) );
  NAND2_X1 U687 ( .A1(n597), .A2(n596), .ZN(n598) );
  XNOR2_X1 U688 ( .A(n598), .B(KEYINPUT32), .ZN(n756) );
  NOR2_X1 U689 ( .A1(n385), .A2(n599), .ZN(n600) );
  AND2_X1 U690 ( .A1(n600), .A2(n387), .ZN(n601) );
  NAND2_X1 U691 ( .A1(n347), .A2(n601), .ZN(n696) );
  NAND2_X1 U692 ( .A1(n756), .A2(n696), .ZN(n605) );
  NAND2_X1 U693 ( .A1(n605), .A2(KEYINPUT44), .ZN(n603) );
  INV_X1 U694 ( .A(KEYINPUT84), .ZN(n604) );
  NOR2_X1 U695 ( .A1(n605), .A2(KEYINPUT44), .ZN(n607) );
  INV_X1 U696 ( .A(n381), .ZN(n606) );
  NAND2_X1 U697 ( .A1(n607), .A2(n606), .ZN(n608) );
  XNOR2_X1 U698 ( .A(KEYINPUT64), .B(KEYINPUT45), .ZN(n609) );
  NAND2_X1 U699 ( .A1(n610), .A2(n734), .ZN(n612) );
  INV_X1 U700 ( .A(KEYINPUT2), .ZN(n611) );
  NAND2_X1 U701 ( .A1(n612), .A2(n611), .ZN(n615) );
  INV_X1 U702 ( .A(n613), .ZN(n614) );
  NAND2_X1 U703 ( .A1(n616), .A2(n734), .ZN(n617) );
  XOR2_X1 U704 ( .A(KEYINPUT54), .B(KEYINPUT55), .Z(n618) );
  XOR2_X1 U705 ( .A(n618), .B(KEYINPUT86), .Z(n619) );
  XNOR2_X1 U706 ( .A(n620), .B(n619), .ZN(n621) );
  XNOR2_X1 U707 ( .A(n622), .B(n621), .ZN(n624) );
  INV_X1 U708 ( .A(G952), .ZN(n623) );
  AND2_X1 U709 ( .A1(n623), .A2(G953), .ZN(n727) );
  XNOR2_X1 U710 ( .A(n625), .B(KEYINPUT56), .ZN(G51) );
  XNOR2_X1 U711 ( .A(n629), .B(KEYINPUT63), .ZN(G57) );
  XNOR2_X1 U712 ( .A(n630), .B(KEYINPUT80), .ZN(n632) );
  NOR2_X1 U713 ( .A1(n632), .A2(n631), .ZN(n634) );
  XNOR2_X1 U714 ( .A(KEYINPUT51), .B(KEYINPUT117), .ZN(n636) );
  XNOR2_X1 U715 ( .A(n636), .B(KEYINPUT116), .ZN(n653) );
  XOR2_X1 U716 ( .A(KEYINPUT115), .B(KEYINPUT50), .Z(n638) );
  XNOR2_X1 U717 ( .A(n639), .B(n638), .ZN(n645) );
  XNOR2_X1 U718 ( .A(KEYINPUT49), .B(KEYINPUT114), .ZN(n643) );
  NOR2_X1 U719 ( .A1(n641), .A2(n640), .ZN(n642) );
  XNOR2_X1 U720 ( .A(n643), .B(n642), .ZN(n644) );
  NAND2_X1 U721 ( .A1(n645), .A2(n644), .ZN(n647) );
  NAND2_X1 U722 ( .A1(n647), .A2(n646), .ZN(n651) );
  NAND2_X1 U723 ( .A1(n649), .A2(n385), .ZN(n650) );
  NAND2_X1 U724 ( .A1(n651), .A2(n650), .ZN(n652) );
  XNOR2_X1 U725 ( .A(n653), .B(n652), .ZN(n654) );
  NOR2_X1 U726 ( .A1(n672), .A2(n654), .ZN(n666) );
  INV_X1 U727 ( .A(n655), .ZN(n663) );
  NOR2_X1 U728 ( .A1(n658), .A2(n410), .ZN(n659) );
  NOR2_X1 U729 ( .A1(n660), .A2(n659), .ZN(n661) );
  OR2_X1 U730 ( .A1(n416), .A2(n661), .ZN(n662) );
  NAND2_X1 U731 ( .A1(n663), .A2(n662), .ZN(n664) );
  AND2_X1 U732 ( .A1(n670), .A2(n664), .ZN(n665) );
  NOR2_X1 U733 ( .A1(n666), .A2(n665), .ZN(n667) );
  XNOR2_X1 U734 ( .A(n667), .B(KEYINPUT52), .ZN(n668) );
  NOR2_X1 U735 ( .A1(n669), .A2(n668), .ZN(n674) );
  INV_X1 U736 ( .A(n670), .ZN(n671) );
  NOR2_X1 U737 ( .A1(n672), .A2(n671), .ZN(n673) );
  OR2_X1 U738 ( .A1(n674), .A2(n673), .ZN(n675) );
  XNOR2_X1 U739 ( .A(KEYINPUT53), .B(KEYINPUT118), .ZN(n676) );
  XNOR2_X1 U740 ( .A(n677), .B(n676), .ZN(G75) );
  XNOR2_X1 U741 ( .A(n678), .B(G140), .ZN(G42) );
  XOR2_X1 U742 ( .A(G125), .B(KEYINPUT37), .Z(n679) );
  XNOR2_X1 U743 ( .A(n680), .B(n679), .ZN(G27) );
  XNOR2_X1 U744 ( .A(n381), .B(n681), .ZN(G24) );
  XOR2_X1 U745 ( .A(n683), .B(G101), .Z(G3) );
  XNOR2_X1 U746 ( .A(KEYINPUT120), .B(KEYINPUT59), .ZN(n684) );
  XNOR2_X1 U747 ( .A(n687), .B(n686), .ZN(n688) );
  XNOR2_X1 U748 ( .A(n689), .B(KEYINPUT60), .ZN(G60) );
  NAND2_X1 U749 ( .A1(n692), .A2(n705), .ZN(n690) );
  XNOR2_X1 U750 ( .A(n690), .B(KEYINPUT110), .ZN(n691) );
  XNOR2_X1 U751 ( .A(G104), .B(n691), .ZN(G6) );
  XOR2_X1 U752 ( .A(KEYINPUT27), .B(KEYINPUT26), .Z(n694) );
  NAND2_X1 U753 ( .A1(n692), .A2(n707), .ZN(n693) );
  XNOR2_X1 U754 ( .A(n694), .B(n693), .ZN(n695) );
  XNOR2_X1 U755 ( .A(G107), .B(n695), .ZN(G9) );
  XNOR2_X1 U756 ( .A(G110), .B(n696), .ZN(G12) );
  NOR2_X1 U757 ( .A1(n703), .A2(n697), .ZN(n699) );
  XNOR2_X1 U758 ( .A(KEYINPUT29), .B(KEYINPUT111), .ZN(n698) );
  XNOR2_X1 U759 ( .A(n699), .B(n698), .ZN(n700) );
  XOR2_X1 U760 ( .A(G128), .B(n700), .Z(G30) );
  XOR2_X1 U761 ( .A(G143), .B(n701), .Z(G45) );
  NOR2_X1 U762 ( .A1(n703), .A2(n702), .ZN(n704) );
  XOR2_X1 U763 ( .A(G146), .B(n704), .Z(G48) );
  XNOR2_X1 U764 ( .A(n706), .B(G113), .ZN(G15) );
  XOR2_X1 U765 ( .A(KEYINPUT112), .B(KEYINPUT113), .Z(n709) );
  XNOR2_X1 U766 ( .A(n709), .B(n708), .ZN(n710) );
  XNOR2_X1 U767 ( .A(G116), .B(n710), .ZN(G18) );
  XNOR2_X1 U768 ( .A(G134), .B(n711), .ZN(G36) );
  NAND2_X1 U769 ( .A1(n721), .A2(G469), .ZN(n716) );
  XOR2_X1 U770 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n712) );
  XNOR2_X1 U771 ( .A(n712), .B(KEYINPUT119), .ZN(n713) );
  XNOR2_X1 U772 ( .A(n714), .B(n713), .ZN(n715) );
  XNOR2_X1 U773 ( .A(n716), .B(n715), .ZN(n717) );
  NOR2_X1 U774 ( .A1(n727), .A2(n717), .ZN(G54) );
  NAND2_X1 U775 ( .A1(n721), .A2(G478), .ZN(n719) );
  XNOR2_X1 U776 ( .A(n719), .B(n718), .ZN(n720) );
  NOR2_X1 U777 ( .A1(n727), .A2(n720), .ZN(G63) );
  NAND2_X1 U778 ( .A1(n721), .A2(G217), .ZN(n725) );
  INV_X1 U779 ( .A(KEYINPUT121), .ZN(n722) );
  NOR2_X1 U780 ( .A1(n727), .A2(n726), .ZN(G66) );
  XNOR2_X1 U781 ( .A(G101), .B(KEYINPUT125), .ZN(n728) );
  XNOR2_X1 U782 ( .A(n729), .B(n728), .ZN(n731) );
  XNOR2_X1 U783 ( .A(n731), .B(n730), .ZN(n732) );
  NOR2_X1 U784 ( .A1(n733), .A2(n732), .ZN(n743) );
  NAND2_X1 U785 ( .A1(n734), .A2(n752), .ZN(n741) );
  XOR2_X1 U786 ( .A(KEYINPUT123), .B(KEYINPUT61), .Z(n736) );
  NAND2_X1 U787 ( .A1(G224), .A2(G953), .ZN(n735) );
  XNOR2_X1 U788 ( .A(n736), .B(n735), .ZN(n737) );
  XNOR2_X1 U789 ( .A(KEYINPUT122), .B(n737), .ZN(n738) );
  NAND2_X1 U790 ( .A1(n738), .A2(G898), .ZN(n739) );
  XNOR2_X1 U791 ( .A(n739), .B(KEYINPUT124), .ZN(n740) );
  NAND2_X1 U792 ( .A1(n741), .A2(n740), .ZN(n742) );
  XNOR2_X1 U793 ( .A(n743), .B(n742), .ZN(G69) );
  XNOR2_X1 U794 ( .A(n744), .B(KEYINPUT4), .ZN(n745) );
  XNOR2_X1 U795 ( .A(n746), .B(n745), .ZN(n751) );
  XOR2_X1 U796 ( .A(KEYINPUT126), .B(n751), .Z(n747) );
  XNOR2_X1 U797 ( .A(G227), .B(n747), .ZN(n748) );
  NAND2_X1 U798 ( .A1(n748), .A2(G900), .ZN(n749) );
  NAND2_X1 U799 ( .A1(n749), .A2(G953), .ZN(n755) );
  XOR2_X1 U800 ( .A(n751), .B(n750), .Z(n753) );
  NAND2_X1 U801 ( .A1(n753), .A2(n752), .ZN(n754) );
  NAND2_X1 U802 ( .A1(n755), .A2(n754), .ZN(G72) );
  XNOR2_X1 U803 ( .A(G119), .B(n756), .ZN(G21) );
  XNOR2_X1 U804 ( .A(G131), .B(KEYINPUT127), .ZN(n758) );
  XNOR2_X1 U805 ( .A(n758), .B(n757), .ZN(G33) );
  XOR2_X1 U806 ( .A(G137), .B(n759), .Z(G39) );
endmodule

