

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n524, n525, n526, n527,
         n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538,
         n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549,
         n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560,
         n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571,
         n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582,
         n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593,
         n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604,
         n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615,
         n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626,
         n627, n628, n629, n630, n631, n632, n633, n634, n635, n636, n637,
         n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, n648,
         n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659,
         n660, n661, n662, n663, n664, n665, n666, n667, n668, n669, n670,
         n671, n672, n673, n674, n675, n676, n677, n678, n679, n680, n681,
         n682, n683, n684, n685, n686, n687, n688, n689, n690, n691, n692,
         n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, n703,
         n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, n714,
         n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, n725,
         n726, n727, n728, n729, n730, n731, n732, n733, n734, n735, n736,
         n737, n738, n739, n740, n741, n742, n743, n744, n745, n746, n747,
         n748, n749, n750, n751, n752, n753, n754, n755, n756, n757, n758,
         n759, n760, n761, n762, n763, n764, n765, n766, n767, n768, n769,
         n770, n771, n772, n773, n774, n775, n776, n777, n778, n779, n780,
         n781, n782, n783, n784, n785, n786, n787, n788, n789, n790, n791,
         n792, n793, n794, n795, n796, n797, n798, n799, n800, n801, n802,
         n803, n804, n805, n806, n807, n808, n809, n810, n811, n812, n813,
         n814, n815, n816, n817, n818, n819, n820, n821, n822, n823, n824,
         n825, n826, n827, n828, n829, n830, n831, n832, n833, n834, n835,
         n836, n837, n838, n839, n840, n841, n842, n843, n844, n845, n846,
         n847, n848, n849, n850, n851, n852, n853, n854, n855, n856, n857,
         n858, n859, n860, n861, n862, n863, n864, n865, n866, n867, n868,
         n869, n870, n871, n872, n873, n874, n875, n876, n877, n878, n879,
         n880, n881, n882, n883, n884, n885, n886, n887, n888, n889, n890,
         n891, n892, n893, n894, n895, n896, n897, n898, n899, n900, n901,
         n902, n903, n904, n905, n906, n907, n908, n909, n910, n911, n912,
         n913, n914, n915, n916, n917, n918, n919, n920, n921, n922, n923,
         n924, n925, n926, n927, n928, n929, n930, n931, n932, n933, n934,
         n935, n936, n937, n938, n939, n940, n941, n942, n943, n944, n945,
         n946, n947, n948, n949, n950, n951, n952, n953, n954, n955, n956,
         n957, n958, n959, n960, n961, n962, n963, n964, n965, n966, n967,
         n968, n969, n970, n971, n972, n973, n974, n975, n976, n977, n978,
         n979, n980, n981, n982, n983, n984, n985, n986, n987, n988, n989,
         n990, n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000,
         n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010,
         n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020,
         n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030,
         n1031, n1032, n1033, n1034, n1035, n1036;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NOR2_X1 U558 ( .A1(G651), .A2(n588), .ZN(n815) );
  NOR2_X1 U559 ( .A1(n696), .A2(n695), .ZN(n697) );
  NOR2_X2 U560 ( .A1(n731), .A2(n604), .ZN(n655) );
  INV_X1 U561 ( .A(n655), .ZN(n680) );
  AND2_X1 U562 ( .A1(G2105), .A2(G2104), .ZN(n908) );
  XNOR2_X1 U563 ( .A(n528), .B(n527), .ZN(n812) );
  NOR2_X4 U564 ( .A1(G2105), .A2(G2104), .ZN(n544) );
  NOR2_X2 U565 ( .A1(n980), .A2(n642), .ZN(n635) );
  AND2_X1 U566 ( .A1(n655), .A2(G1996), .ZN(n619) );
  XNOR2_X1 U567 ( .A(n680), .B(n606), .ZN(n636) );
  NOR2_X1 U568 ( .A1(G299), .A2(n647), .ZN(n610) );
  NAND2_X1 U569 ( .A1(n671), .A2(n670), .ZN(n678) );
  XNOR2_X1 U570 ( .A(n687), .B(KEYINPUT32), .ZN(n688) );
  NOR2_X2 U571 ( .A1(G2104), .A2(n547), .ZN(n558) );
  AND2_X1 U572 ( .A1(n986), .A2(n768), .ZN(n524) );
  XNOR2_X1 U573 ( .A(n675), .B(n674), .ZN(n676) );
  AND2_X1 U574 ( .A1(n678), .A2(n673), .ZN(n675) );
  NAND2_X2 U575 ( .A1(G160), .A2(G40), .ZN(n731) );
  XOR2_X2 U576 ( .A(KEYINPUT17), .B(n544), .Z(n718) );
  XNOR2_X2 U577 ( .A(n562), .B(n561), .ZN(G160) );
  OR2_X1 U578 ( .A1(n679), .A2(n716), .ZN(n525) );
  XOR2_X1 U579 ( .A(n631), .B(KEYINPUT13), .Z(n526) );
  INV_X1 U580 ( .A(KEYINPUT88), .ZN(n606) );
  INV_X1 U581 ( .A(KEYINPUT96), .ZN(n664) );
  INV_X1 U582 ( .A(KEYINPUT29), .ZN(n652) );
  INV_X1 U583 ( .A(KEYINPUT97), .ZN(n674) );
  INV_X1 U584 ( .A(G2104), .ZN(n542) );
  INV_X1 U585 ( .A(KEYINPUT100), .ZN(n713) );
  NAND2_X1 U586 ( .A1(n812), .A2(G56), .ZN(n623) );
  NOR2_X1 U587 ( .A1(G164), .A2(G1384), .ZN(n733) );
  INV_X1 U588 ( .A(G2105), .ZN(n547) );
  NOR2_X1 U589 ( .A1(n754), .A2(n524), .ZN(n755) );
  NOR2_X2 U590 ( .A1(n588), .A2(n534), .ZN(n816) );
  INV_X1 U591 ( .A(KEYINPUT1), .ZN(n527) );
  INV_X1 U592 ( .A(KEYINPUT66), .ZN(n561) );
  INV_X1 U593 ( .A(G651), .ZN(n534) );
  NOR2_X1 U594 ( .A1(G543), .A2(n534), .ZN(n528) );
  NAND2_X1 U595 ( .A1(G63), .A2(n812), .ZN(n530) );
  XOR2_X1 U596 ( .A(G543), .B(KEYINPUT0), .Z(n588) );
  NAND2_X1 U597 ( .A1(G51), .A2(n815), .ZN(n529) );
  NAND2_X1 U598 ( .A1(n530), .A2(n529), .ZN(n531) );
  XNOR2_X1 U599 ( .A(KEYINPUT6), .B(n531), .ZN(n539) );
  NOR2_X2 U600 ( .A1(G651), .A2(G543), .ZN(n810) );
  NAND2_X1 U601 ( .A1(G89), .A2(n810), .ZN(n532) );
  XOR2_X1 U602 ( .A(KEYINPUT4), .B(n532), .Z(n533) );
  XNOR2_X1 U603 ( .A(n533), .B(KEYINPUT75), .ZN(n536) );
  NAND2_X1 U604 ( .A1(G76), .A2(n816), .ZN(n535) );
  NAND2_X1 U605 ( .A1(n536), .A2(n535), .ZN(n537) );
  XOR2_X1 U606 ( .A(n537), .B(KEYINPUT5), .Z(n538) );
  NOR2_X1 U607 ( .A1(n539), .A2(n538), .ZN(n540) );
  XOR2_X1 U608 ( .A(KEYINPUT76), .B(n540), .Z(n541) );
  XNOR2_X1 U609 ( .A(KEYINPUT7), .B(n541), .ZN(G168) );
  XOR2_X1 U610 ( .A(KEYINPUT8), .B(G168), .Z(G286) );
  NOR2_X1 U611 ( .A1(n542), .A2(G2105), .ZN(n554) );
  BUF_X1 U612 ( .A(n554), .Z(n543) );
  NAND2_X1 U613 ( .A1(G102), .A2(n543), .ZN(n546) );
  NAND2_X1 U614 ( .A1(G138), .A2(n718), .ZN(n545) );
  NAND2_X1 U615 ( .A1(n546), .A2(n545), .ZN(n551) );
  NAND2_X1 U616 ( .A1(G114), .A2(n908), .ZN(n549) );
  NAND2_X1 U617 ( .A1(G126), .A2(n558), .ZN(n548) );
  NAND2_X1 U618 ( .A1(n549), .A2(n548), .ZN(n550) );
  NOR2_X1 U619 ( .A1(n551), .A2(n550), .ZN(G164) );
  NAND2_X1 U620 ( .A1(n718), .A2(G137), .ZN(n553) );
  NAND2_X1 U621 ( .A1(G113), .A2(n908), .ZN(n552) );
  NAND2_X1 U622 ( .A1(n553), .A2(n552), .ZN(n557) );
  AND2_X1 U623 ( .A1(G101), .A2(n554), .ZN(n555) );
  XOR2_X1 U624 ( .A(KEYINPUT23), .B(n555), .Z(n556) );
  NOR2_X1 U625 ( .A1(n557), .A2(n556), .ZN(n560) );
  NAND2_X1 U626 ( .A1(n558), .A2(G125), .ZN(n559) );
  NAND2_X1 U627 ( .A1(n560), .A2(n559), .ZN(n562) );
  NAND2_X1 U628 ( .A1(G65), .A2(n812), .ZN(n564) );
  NAND2_X1 U629 ( .A1(G53), .A2(n815), .ZN(n563) );
  NAND2_X1 U630 ( .A1(n564), .A2(n563), .ZN(n568) );
  NAND2_X1 U631 ( .A1(G91), .A2(n810), .ZN(n566) );
  NAND2_X1 U632 ( .A1(G78), .A2(n816), .ZN(n565) );
  NAND2_X1 U633 ( .A1(n566), .A2(n565), .ZN(n567) );
  NOR2_X1 U634 ( .A1(n568), .A2(n567), .ZN(n569) );
  XOR2_X1 U635 ( .A(KEYINPUT68), .B(n569), .Z(G299) );
  NAND2_X1 U636 ( .A1(G64), .A2(n812), .ZN(n571) );
  NAND2_X1 U637 ( .A1(G52), .A2(n815), .ZN(n570) );
  NAND2_X1 U638 ( .A1(n571), .A2(n570), .ZN(n572) );
  XOR2_X1 U639 ( .A(KEYINPUT67), .B(n572), .Z(n577) );
  NAND2_X1 U640 ( .A1(G90), .A2(n810), .ZN(n574) );
  NAND2_X1 U641 ( .A1(G77), .A2(n816), .ZN(n573) );
  NAND2_X1 U642 ( .A1(n574), .A2(n573), .ZN(n575) );
  XOR2_X1 U643 ( .A(KEYINPUT9), .B(n575), .Z(n576) );
  NOR2_X1 U644 ( .A1(n577), .A2(n576), .ZN(G171) );
  INV_X1 U645 ( .A(G171), .ZN(G301) );
  NAND2_X1 U646 ( .A1(G62), .A2(n812), .ZN(n579) );
  NAND2_X1 U647 ( .A1(G50), .A2(n815), .ZN(n578) );
  NAND2_X1 U648 ( .A1(n579), .A2(n578), .ZN(n583) );
  NAND2_X1 U649 ( .A1(G88), .A2(n810), .ZN(n581) );
  NAND2_X1 U650 ( .A1(G75), .A2(n816), .ZN(n580) );
  NAND2_X1 U651 ( .A1(n581), .A2(n580), .ZN(n582) );
  NOR2_X1 U652 ( .A1(n583), .A2(n582), .ZN(n584) );
  XOR2_X1 U653 ( .A(KEYINPUT79), .B(n584), .Z(G166) );
  INV_X1 U654 ( .A(G166), .ZN(G303) );
  NAND2_X1 U655 ( .A1(G49), .A2(n815), .ZN(n586) );
  NAND2_X1 U656 ( .A1(G74), .A2(G651), .ZN(n585) );
  NAND2_X1 U657 ( .A1(n586), .A2(n585), .ZN(n587) );
  NOR2_X1 U658 ( .A1(n812), .A2(n587), .ZN(n590) );
  NAND2_X1 U659 ( .A1(n588), .A2(G87), .ZN(n589) );
  NAND2_X1 U660 ( .A1(n590), .A2(n589), .ZN(G288) );
  NAND2_X1 U661 ( .A1(G61), .A2(n812), .ZN(n592) );
  NAND2_X1 U662 ( .A1(G48), .A2(n815), .ZN(n591) );
  NAND2_X1 U663 ( .A1(n592), .A2(n591), .ZN(n595) );
  NAND2_X1 U664 ( .A1(n816), .A2(G73), .ZN(n593) );
  XOR2_X1 U665 ( .A(KEYINPUT2), .B(n593), .Z(n594) );
  NOR2_X1 U666 ( .A1(n595), .A2(n594), .ZN(n597) );
  NAND2_X1 U667 ( .A1(n810), .A2(G86), .ZN(n596) );
  NAND2_X1 U668 ( .A1(n597), .A2(n596), .ZN(G305) );
  NAND2_X1 U669 ( .A1(G60), .A2(n812), .ZN(n599) );
  NAND2_X1 U670 ( .A1(G47), .A2(n815), .ZN(n598) );
  NAND2_X1 U671 ( .A1(n599), .A2(n598), .ZN(n603) );
  NAND2_X1 U672 ( .A1(G85), .A2(n810), .ZN(n601) );
  NAND2_X1 U673 ( .A1(G72), .A2(n816), .ZN(n600) );
  NAND2_X1 U674 ( .A1(n601), .A2(n600), .ZN(n602) );
  OR2_X1 U675 ( .A1(n603), .A2(n602), .ZN(G290) );
  INV_X1 U676 ( .A(n733), .ZN(n604) );
  NOR2_X1 U677 ( .A1(G2084), .A2(n680), .ZN(n660) );
  NAND2_X1 U678 ( .A1(G8), .A2(n660), .ZN(n677) );
  XNOR2_X1 U679 ( .A(KEYINPUT88), .B(n680), .ZN(n654) );
  XOR2_X1 U680 ( .A(G1956), .B(KEYINPUT89), .Z(n1015) );
  NAND2_X1 U681 ( .A1(n654), .A2(n1015), .ZN(n605) );
  XNOR2_X1 U682 ( .A(KEYINPUT90), .B(n605), .ZN(n609) );
  AND2_X1 U683 ( .A1(G2072), .A2(n636), .ZN(n607) );
  XNOR2_X1 U684 ( .A(n607), .B(KEYINPUT27), .ZN(n608) );
  NAND2_X1 U685 ( .A1(n609), .A2(n608), .ZN(n647) );
  XNOR2_X1 U686 ( .A(n610), .B(KEYINPUT95), .ZN(n646) );
  NAND2_X1 U687 ( .A1(G92), .A2(n810), .ZN(n612) );
  NAND2_X1 U688 ( .A1(G79), .A2(n816), .ZN(n611) );
  NAND2_X1 U689 ( .A1(n612), .A2(n611), .ZN(n616) );
  NAND2_X1 U690 ( .A1(G66), .A2(n812), .ZN(n614) );
  NAND2_X1 U691 ( .A1(G54), .A2(n815), .ZN(n613) );
  NAND2_X1 U692 ( .A1(n614), .A2(n613), .ZN(n615) );
  NOR2_X1 U693 ( .A1(n616), .A2(n615), .ZN(n617) );
  XNOR2_X1 U694 ( .A(n617), .B(KEYINPUT15), .ZN(n980) );
  XNOR2_X1 U695 ( .A(KEYINPUT65), .B(KEYINPUT26), .ZN(n618) );
  XNOR2_X1 U696 ( .A(n619), .B(n618), .ZN(n621) );
  NAND2_X1 U697 ( .A1(n680), .A2(G1341), .ZN(n620) );
  NAND2_X1 U698 ( .A1(n621), .A2(n620), .ZN(n622) );
  XOR2_X1 U699 ( .A(n622), .B(KEYINPUT92), .Z(n634) );
  XNOR2_X1 U700 ( .A(n623), .B(KEYINPUT14), .ZN(n625) );
  NAND2_X1 U701 ( .A1(G43), .A2(n815), .ZN(n624) );
  NAND2_X1 U702 ( .A1(n625), .A2(n624), .ZN(n632) );
  XOR2_X1 U703 ( .A(KEYINPUT12), .B(KEYINPUT71), .Z(n627) );
  NAND2_X1 U704 ( .A1(G81), .A2(n810), .ZN(n626) );
  XNOR2_X1 U705 ( .A(n627), .B(n626), .ZN(n628) );
  XNOR2_X1 U706 ( .A(KEYINPUT70), .B(n628), .ZN(n630) );
  NAND2_X1 U707 ( .A1(n816), .A2(G68), .ZN(n629) );
  NAND2_X1 U708 ( .A1(n630), .A2(n629), .ZN(n631) );
  NOR2_X1 U709 ( .A1(n632), .A2(n526), .ZN(n633) );
  XNOR2_X1 U710 ( .A(KEYINPUT72), .B(n633), .ZN(n978) );
  NAND2_X1 U711 ( .A1(n634), .A2(n978), .ZN(n642) );
  XNOR2_X1 U712 ( .A(n635), .B(KEYINPUT93), .ZN(n641) );
  NAND2_X1 U713 ( .A1(G2067), .A2(n636), .ZN(n638) );
  NAND2_X1 U714 ( .A1(G1348), .A2(n680), .ZN(n637) );
  NAND2_X1 U715 ( .A1(n638), .A2(n637), .ZN(n639) );
  XNOR2_X1 U716 ( .A(KEYINPUT94), .B(n639), .ZN(n640) );
  NAND2_X1 U717 ( .A1(n641), .A2(n640), .ZN(n644) );
  NAND2_X1 U718 ( .A1(n980), .A2(n642), .ZN(n643) );
  NAND2_X1 U719 ( .A1(n644), .A2(n643), .ZN(n645) );
  NAND2_X1 U720 ( .A1(n646), .A2(n645), .ZN(n651) );
  XOR2_X1 U721 ( .A(KEYINPUT91), .B(KEYINPUT28), .Z(n649) );
  NAND2_X1 U722 ( .A1(G299), .A2(n647), .ZN(n648) );
  XNOR2_X1 U723 ( .A(n649), .B(n648), .ZN(n650) );
  NAND2_X1 U724 ( .A1(n651), .A2(n650), .ZN(n653) );
  XNOR2_X1 U725 ( .A(n653), .B(n652), .ZN(n659) );
  XOR2_X1 U726 ( .A(G2078), .B(KEYINPUT25), .Z(n961) );
  NOR2_X1 U727 ( .A1(n961), .A2(n654), .ZN(n657) );
  NOR2_X1 U728 ( .A1(n655), .A2(G1961), .ZN(n656) );
  NOR2_X1 U729 ( .A1(n657), .A2(n656), .ZN(n666) );
  OR2_X1 U730 ( .A1(n666), .A2(G301), .ZN(n658) );
  NAND2_X1 U731 ( .A1(n659), .A2(n658), .ZN(n671) );
  NAND2_X1 U732 ( .A1(G8), .A2(n680), .ZN(n679) );
  NOR2_X1 U733 ( .A1(G1966), .A2(n679), .ZN(n672) );
  NOR2_X1 U734 ( .A1(n660), .A2(n672), .ZN(n661) );
  NAND2_X1 U735 ( .A1(G8), .A2(n661), .ZN(n662) );
  XNOR2_X1 U736 ( .A(KEYINPUT30), .B(n662), .ZN(n663) );
  NOR2_X1 U737 ( .A1(G168), .A2(n663), .ZN(n665) );
  XNOR2_X1 U738 ( .A(n665), .B(n664), .ZN(n668) );
  NAND2_X1 U739 ( .A1(n666), .A2(G301), .ZN(n667) );
  NAND2_X1 U740 ( .A1(n668), .A2(n667), .ZN(n669) );
  XNOR2_X1 U741 ( .A(KEYINPUT31), .B(n669), .ZN(n670) );
  INV_X1 U742 ( .A(n672), .ZN(n673) );
  NAND2_X1 U743 ( .A1(n677), .A2(n676), .ZN(n689) );
  NAND2_X1 U744 ( .A1(n678), .A2(G286), .ZN(n685) );
  NOR2_X1 U745 ( .A1(G1971), .A2(n679), .ZN(n682) );
  NOR2_X1 U746 ( .A1(G2090), .A2(n680), .ZN(n681) );
  NOR2_X1 U747 ( .A1(n682), .A2(n681), .ZN(n683) );
  NAND2_X1 U748 ( .A1(n683), .A2(G303), .ZN(n684) );
  NAND2_X1 U749 ( .A1(n685), .A2(n684), .ZN(n686) );
  NAND2_X1 U750 ( .A1(n686), .A2(G8), .ZN(n687) );
  NAND2_X1 U751 ( .A1(n689), .A2(n688), .ZN(n708) );
  NOR2_X1 U752 ( .A1(G1976), .A2(G288), .ZN(n700) );
  NOR2_X1 U753 ( .A1(G1971), .A2(G303), .ZN(n690) );
  NOR2_X1 U754 ( .A1(n700), .A2(n690), .ZN(n991) );
  NAND2_X1 U755 ( .A1(n708), .A2(n991), .ZN(n693) );
  NAND2_X1 U756 ( .A1(G288), .A2(G1976), .ZN(n691) );
  XOR2_X1 U757 ( .A(KEYINPUT98), .B(n691), .Z(n990) );
  NOR2_X1 U758 ( .A1(n679), .A2(n990), .ZN(n692) );
  NAND2_X1 U759 ( .A1(n693), .A2(n692), .ZN(n694) );
  XNOR2_X1 U760 ( .A(n694), .B(KEYINPUT64), .ZN(n696) );
  INV_X1 U761 ( .A(KEYINPUT99), .ZN(n699) );
  NOR2_X1 U762 ( .A1(n679), .A2(n699), .ZN(n695) );
  NOR2_X1 U763 ( .A1(n697), .A2(KEYINPUT33), .ZN(n705) );
  NAND2_X1 U764 ( .A1(n700), .A2(KEYINPUT33), .ZN(n698) );
  NAND2_X1 U765 ( .A1(n699), .A2(n698), .ZN(n702) );
  NAND2_X1 U766 ( .A1(n700), .A2(KEYINPUT99), .ZN(n701) );
  NAND2_X1 U767 ( .A1(n702), .A2(n701), .ZN(n703) );
  NOR2_X1 U768 ( .A1(n679), .A2(n703), .ZN(n704) );
  NOR2_X1 U769 ( .A1(n705), .A2(n704), .ZN(n706) );
  XOR2_X1 U770 ( .A(G1981), .B(G305), .Z(n996) );
  NAND2_X1 U771 ( .A1(n706), .A2(n996), .ZN(n712) );
  NOR2_X1 U772 ( .A1(G2090), .A2(G303), .ZN(n707) );
  NAND2_X1 U773 ( .A1(G8), .A2(n707), .ZN(n709) );
  NAND2_X1 U774 ( .A1(n709), .A2(n708), .ZN(n710) );
  NAND2_X1 U775 ( .A1(n710), .A2(n679), .ZN(n711) );
  NAND2_X1 U776 ( .A1(n712), .A2(n711), .ZN(n714) );
  XNOR2_X1 U777 ( .A(n714), .B(n713), .ZN(n717) );
  NOR2_X1 U778 ( .A1(G1981), .A2(G305), .ZN(n715) );
  XOR2_X1 U779 ( .A(n715), .B(KEYINPUT24), .Z(n716) );
  NAND2_X1 U780 ( .A1(n717), .A2(n525), .ZN(n756) );
  NAND2_X1 U781 ( .A1(G104), .A2(n543), .ZN(n720) );
  BUF_X1 U782 ( .A(n718), .Z(n905) );
  NAND2_X1 U783 ( .A1(G140), .A2(n905), .ZN(n719) );
  NAND2_X1 U784 ( .A1(n720), .A2(n719), .ZN(n721) );
  XNOR2_X1 U785 ( .A(KEYINPUT34), .B(n721), .ZN(n727) );
  NAND2_X1 U786 ( .A1(n908), .A2(G116), .ZN(n722) );
  XOR2_X1 U787 ( .A(KEYINPUT81), .B(n722), .Z(n724) );
  NAND2_X1 U788 ( .A1(n558), .A2(G128), .ZN(n723) );
  NAND2_X1 U789 ( .A1(n724), .A2(n723), .ZN(n725) );
  XOR2_X1 U790 ( .A(n725), .B(KEYINPUT35), .Z(n726) );
  NOR2_X1 U791 ( .A1(n727), .A2(n726), .ZN(n728) );
  XOR2_X1 U792 ( .A(KEYINPUT36), .B(n728), .Z(n729) );
  XOR2_X1 U793 ( .A(KEYINPUT82), .B(n729), .Z(n918) );
  XNOR2_X1 U794 ( .A(G2067), .B(KEYINPUT37), .ZN(n766) );
  OR2_X1 U795 ( .A1(n918), .A2(n766), .ZN(n730) );
  XNOR2_X1 U796 ( .A(n730), .B(KEYINPUT83), .ZN(n951) );
  BUF_X1 U797 ( .A(n731), .Z(n732) );
  NOR2_X1 U798 ( .A1(n733), .A2(n732), .ZN(n768) );
  NAND2_X1 U799 ( .A1(n951), .A2(n768), .ZN(n734) );
  XNOR2_X1 U800 ( .A(n734), .B(KEYINPUT84), .ZN(n764) );
  XOR2_X1 U801 ( .A(KEYINPUT38), .B(KEYINPUT86), .Z(n736) );
  NAND2_X1 U802 ( .A1(G105), .A2(n543), .ZN(n735) );
  XNOR2_X1 U803 ( .A(n736), .B(n735), .ZN(n740) );
  NAND2_X1 U804 ( .A1(G141), .A2(n905), .ZN(n738) );
  NAND2_X1 U805 ( .A1(G117), .A2(n908), .ZN(n737) );
  NAND2_X1 U806 ( .A1(n738), .A2(n737), .ZN(n739) );
  NOR2_X1 U807 ( .A1(n740), .A2(n739), .ZN(n742) );
  NAND2_X1 U808 ( .A1(n558), .A2(G129), .ZN(n741) );
  NAND2_X1 U809 ( .A1(n742), .A2(n741), .ZN(n898) );
  NAND2_X1 U810 ( .A1(G1996), .A2(n898), .ZN(n751) );
  NAND2_X1 U811 ( .A1(G95), .A2(n543), .ZN(n744) );
  NAND2_X1 U812 ( .A1(G131), .A2(n905), .ZN(n743) );
  NAND2_X1 U813 ( .A1(n744), .A2(n743), .ZN(n747) );
  NAND2_X1 U814 ( .A1(G107), .A2(n908), .ZN(n745) );
  XNOR2_X1 U815 ( .A(KEYINPUT85), .B(n745), .ZN(n746) );
  NOR2_X1 U816 ( .A1(n747), .A2(n746), .ZN(n749) );
  NAND2_X1 U817 ( .A1(n558), .A2(G119), .ZN(n748) );
  NAND2_X1 U818 ( .A1(n749), .A2(n748), .ZN(n915) );
  NAND2_X1 U819 ( .A1(G1991), .A2(n915), .ZN(n750) );
  NAND2_X1 U820 ( .A1(n751), .A2(n750), .ZN(n752) );
  XNOR2_X1 U821 ( .A(KEYINPUT87), .B(n752), .ZN(n934) );
  INV_X1 U822 ( .A(n934), .ZN(n753) );
  NAND2_X1 U823 ( .A1(n753), .A2(n768), .ZN(n757) );
  NAND2_X1 U824 ( .A1(n764), .A2(n757), .ZN(n754) );
  XNOR2_X1 U825 ( .A(G1986), .B(G290), .ZN(n986) );
  NAND2_X1 U826 ( .A1(n756), .A2(n755), .ZN(n771) );
  NOR2_X1 U827 ( .A1(G1996), .A2(n898), .ZN(n944) );
  INV_X1 U828 ( .A(n757), .ZN(n760) );
  NOR2_X1 U829 ( .A1(G1991), .A2(n915), .ZN(n936) );
  NOR2_X1 U830 ( .A1(G1986), .A2(G290), .ZN(n758) );
  NOR2_X1 U831 ( .A1(n936), .A2(n758), .ZN(n759) );
  NOR2_X1 U832 ( .A1(n760), .A2(n759), .ZN(n761) );
  XOR2_X1 U833 ( .A(KEYINPUT101), .B(n761), .Z(n762) );
  NOR2_X1 U834 ( .A1(n944), .A2(n762), .ZN(n763) );
  XNOR2_X1 U835 ( .A(n763), .B(KEYINPUT39), .ZN(n765) );
  NAND2_X1 U836 ( .A1(n765), .A2(n764), .ZN(n767) );
  NAND2_X1 U837 ( .A1(n918), .A2(n766), .ZN(n941) );
  NAND2_X1 U838 ( .A1(n767), .A2(n941), .ZN(n769) );
  NAND2_X1 U839 ( .A1(n769), .A2(n768), .ZN(n770) );
  NAND2_X1 U840 ( .A1(n771), .A2(n770), .ZN(n772) );
  XNOR2_X1 U841 ( .A(n772), .B(KEYINPUT40), .ZN(G329) );
  XOR2_X1 U842 ( .A(G2451), .B(G2454), .Z(n774) );
  XNOR2_X1 U843 ( .A(G2430), .B(KEYINPUT102), .ZN(n773) );
  XNOR2_X1 U844 ( .A(n774), .B(n773), .ZN(n775) );
  XOR2_X1 U845 ( .A(n775), .B(G2446), .Z(n777) );
  XNOR2_X1 U846 ( .A(G1341), .B(G1348), .ZN(n776) );
  XNOR2_X1 U847 ( .A(n777), .B(n776), .ZN(n781) );
  XOR2_X1 U848 ( .A(G2438), .B(G2427), .Z(n779) );
  XNOR2_X1 U849 ( .A(G2443), .B(G2435), .ZN(n778) );
  XNOR2_X1 U850 ( .A(n779), .B(n778), .ZN(n780) );
  XOR2_X1 U851 ( .A(n781), .B(n780), .Z(n782) );
  AND2_X1 U852 ( .A1(G14), .A2(n782), .ZN(G401) );
  AND2_X1 U853 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U854 ( .A(G132), .ZN(G219) );
  INV_X1 U855 ( .A(G82), .ZN(G220) );
  INV_X1 U856 ( .A(G57), .ZN(G237) );
  XOR2_X1 U857 ( .A(KEYINPUT69), .B(KEYINPUT10), .Z(n784) );
  NAND2_X1 U858 ( .A1(G7), .A2(G661), .ZN(n783) );
  XNOR2_X1 U859 ( .A(n784), .B(n783), .ZN(G223) );
  INV_X1 U860 ( .A(G223), .ZN(n846) );
  NAND2_X1 U861 ( .A1(n846), .A2(G567), .ZN(n785) );
  XOR2_X1 U862 ( .A(KEYINPUT11), .B(n785), .Z(G234) );
  XOR2_X1 U863 ( .A(G860), .B(KEYINPUT73), .Z(n792) );
  NAND2_X1 U864 ( .A1(n792), .A2(n978), .ZN(G153) );
  INV_X1 U865 ( .A(G868), .ZN(n830) );
  NAND2_X1 U866 ( .A1(n980), .A2(n830), .ZN(n786) );
  XNOR2_X1 U867 ( .A(n786), .B(KEYINPUT74), .ZN(n788) );
  NAND2_X1 U868 ( .A1(G868), .A2(G301), .ZN(n787) );
  NAND2_X1 U869 ( .A1(n788), .A2(n787), .ZN(G284) );
  NAND2_X1 U870 ( .A1(G868), .A2(G286), .ZN(n790) );
  NAND2_X1 U871 ( .A1(G299), .A2(n830), .ZN(n789) );
  NAND2_X1 U872 ( .A1(n790), .A2(n789), .ZN(G297) );
  INV_X1 U873 ( .A(G559), .ZN(n791) );
  NOR2_X1 U874 ( .A1(n792), .A2(n791), .ZN(n793) );
  NOR2_X1 U875 ( .A1(n980), .A2(n793), .ZN(n794) );
  XOR2_X1 U876 ( .A(KEYINPUT16), .B(n794), .Z(G148) );
  INV_X1 U877 ( .A(n980), .ZN(n808) );
  NAND2_X1 U878 ( .A1(n808), .A2(G868), .ZN(n795) );
  NOR2_X1 U879 ( .A1(G559), .A2(n795), .ZN(n797) );
  AND2_X1 U880 ( .A1(n978), .A2(n830), .ZN(n796) );
  NOR2_X1 U881 ( .A1(n797), .A2(n796), .ZN(G282) );
  NAND2_X1 U882 ( .A1(G99), .A2(n543), .ZN(n799) );
  NAND2_X1 U883 ( .A1(G111), .A2(n908), .ZN(n798) );
  NAND2_X1 U884 ( .A1(n799), .A2(n798), .ZN(n800) );
  XNOR2_X1 U885 ( .A(n800), .B(KEYINPUT77), .ZN(n802) );
  NAND2_X1 U886 ( .A1(G135), .A2(n905), .ZN(n801) );
  NAND2_X1 U887 ( .A1(n802), .A2(n801), .ZN(n805) );
  NAND2_X1 U888 ( .A1(n558), .A2(G123), .ZN(n803) );
  XOR2_X1 U889 ( .A(KEYINPUT18), .B(n803), .Z(n804) );
  NOR2_X1 U890 ( .A1(n805), .A2(n804), .ZN(n932) );
  XNOR2_X1 U891 ( .A(n932), .B(G2096), .ZN(n807) );
  INV_X1 U892 ( .A(G2100), .ZN(n806) );
  NAND2_X1 U893 ( .A1(n807), .A2(n806), .ZN(G156) );
  NAND2_X1 U894 ( .A1(G559), .A2(n808), .ZN(n809) );
  XOR2_X1 U895 ( .A(n978), .B(n809), .Z(n827) );
  NOR2_X1 U896 ( .A1(G860), .A2(n827), .ZN(n821) );
  NAND2_X1 U897 ( .A1(G93), .A2(n810), .ZN(n811) );
  XNOR2_X1 U898 ( .A(n811), .B(KEYINPUT78), .ZN(n814) );
  NAND2_X1 U899 ( .A1(n812), .A2(G67), .ZN(n813) );
  NAND2_X1 U900 ( .A1(n814), .A2(n813), .ZN(n820) );
  NAND2_X1 U901 ( .A1(G55), .A2(n815), .ZN(n818) );
  NAND2_X1 U902 ( .A1(G80), .A2(n816), .ZN(n817) );
  NAND2_X1 U903 ( .A1(n818), .A2(n817), .ZN(n819) );
  OR2_X1 U904 ( .A1(n820), .A2(n819), .ZN(n829) );
  XOR2_X1 U905 ( .A(n821), .B(n829), .Z(G145) );
  XNOR2_X1 U906 ( .A(KEYINPUT19), .B(G288), .ZN(n826) );
  XNOR2_X1 U907 ( .A(G299), .B(G305), .ZN(n822) );
  XNOR2_X1 U908 ( .A(n822), .B(G303), .ZN(n823) );
  XOR2_X1 U909 ( .A(n829), .B(n823), .Z(n824) );
  XNOR2_X1 U910 ( .A(n824), .B(G290), .ZN(n825) );
  XNOR2_X1 U911 ( .A(n826), .B(n825), .ZN(n855) );
  XNOR2_X1 U912 ( .A(n827), .B(n855), .ZN(n828) );
  NAND2_X1 U913 ( .A1(n828), .A2(G868), .ZN(n832) );
  NAND2_X1 U914 ( .A1(n830), .A2(n829), .ZN(n831) );
  NAND2_X1 U915 ( .A1(n832), .A2(n831), .ZN(G295) );
  NAND2_X1 U916 ( .A1(G2084), .A2(G2078), .ZN(n833) );
  XOR2_X1 U917 ( .A(KEYINPUT20), .B(n833), .Z(n834) );
  NAND2_X1 U918 ( .A1(G2090), .A2(n834), .ZN(n835) );
  XNOR2_X1 U919 ( .A(KEYINPUT21), .B(n835), .ZN(n836) );
  NAND2_X1 U920 ( .A1(n836), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U921 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NAND2_X1 U922 ( .A1(G120), .A2(G69), .ZN(n837) );
  XNOR2_X1 U923 ( .A(KEYINPUT80), .B(n837), .ZN(n838) );
  NOR2_X1 U924 ( .A1(G237), .A2(n838), .ZN(n839) );
  NAND2_X1 U925 ( .A1(G108), .A2(n839), .ZN(n852) );
  NAND2_X1 U926 ( .A1(n852), .A2(G567), .ZN(n844) );
  NOR2_X1 U927 ( .A1(G220), .A2(G219), .ZN(n840) );
  XOR2_X1 U928 ( .A(KEYINPUT22), .B(n840), .Z(n841) );
  NOR2_X1 U929 ( .A1(G218), .A2(n841), .ZN(n842) );
  NAND2_X1 U930 ( .A1(G96), .A2(n842), .ZN(n853) );
  NAND2_X1 U931 ( .A1(n853), .A2(G2106), .ZN(n843) );
  NAND2_X1 U932 ( .A1(n844), .A2(n843), .ZN(n930) );
  NAND2_X1 U933 ( .A1(G483), .A2(G661), .ZN(n845) );
  NOR2_X1 U934 ( .A1(n930), .A2(n845), .ZN(n851) );
  NAND2_X1 U935 ( .A1(n851), .A2(G36), .ZN(G176) );
  NAND2_X1 U936 ( .A1(G2106), .A2(n846), .ZN(G217) );
  NAND2_X1 U937 ( .A1(G15), .A2(G2), .ZN(n848) );
  INV_X1 U938 ( .A(G661), .ZN(n847) );
  NOR2_X1 U939 ( .A1(n848), .A2(n847), .ZN(n849) );
  XNOR2_X1 U940 ( .A(n849), .B(KEYINPUT103), .ZN(G259) );
  NAND2_X1 U941 ( .A1(G3), .A2(G1), .ZN(n850) );
  NAND2_X1 U942 ( .A1(n851), .A2(n850), .ZN(G188) );
  XOR2_X1 U943 ( .A(G120), .B(KEYINPUT104), .Z(G236) );
  XNOR2_X1 U944 ( .A(G69), .B(KEYINPUT105), .ZN(G235) );
  XNOR2_X1 U945 ( .A(G108), .B(KEYINPUT119), .ZN(G238) );
  INV_X1 U947 ( .A(G96), .ZN(G221) );
  NOR2_X1 U948 ( .A1(n853), .A2(n852), .ZN(G325) );
  INV_X1 U949 ( .A(G325), .ZN(G261) );
  XNOR2_X1 U950 ( .A(G171), .B(n980), .ZN(n854) );
  XNOR2_X1 U951 ( .A(n854), .B(G286), .ZN(n857) );
  XOR2_X1 U952 ( .A(n978), .B(n855), .Z(n856) );
  XNOR2_X1 U953 ( .A(n857), .B(n856), .ZN(n858) );
  NOR2_X1 U954 ( .A1(G37), .A2(n858), .ZN(G397) );
  XNOR2_X1 U955 ( .A(G1956), .B(KEYINPUT41), .ZN(n868) );
  XOR2_X1 U956 ( .A(G1976), .B(G1971), .Z(n860) );
  XNOR2_X1 U957 ( .A(G1986), .B(G1961), .ZN(n859) );
  XNOR2_X1 U958 ( .A(n860), .B(n859), .ZN(n864) );
  XOR2_X1 U959 ( .A(G1966), .B(G1981), .Z(n862) );
  XNOR2_X1 U960 ( .A(G1996), .B(G1991), .ZN(n861) );
  XNOR2_X1 U961 ( .A(n862), .B(n861), .ZN(n863) );
  XOR2_X1 U962 ( .A(n864), .B(n863), .Z(n866) );
  XNOR2_X1 U963 ( .A(KEYINPUT108), .B(G2474), .ZN(n865) );
  XNOR2_X1 U964 ( .A(n866), .B(n865), .ZN(n867) );
  XNOR2_X1 U965 ( .A(n868), .B(n867), .ZN(G229) );
  XOR2_X1 U966 ( .A(KEYINPUT43), .B(G2678), .Z(n870) );
  XNOR2_X1 U967 ( .A(KEYINPUT107), .B(KEYINPUT106), .ZN(n869) );
  XNOR2_X1 U968 ( .A(n870), .B(n869), .ZN(n874) );
  XOR2_X1 U969 ( .A(KEYINPUT42), .B(G2072), .Z(n872) );
  XNOR2_X1 U970 ( .A(G2067), .B(G2090), .ZN(n871) );
  XNOR2_X1 U971 ( .A(n872), .B(n871), .ZN(n873) );
  XOR2_X1 U972 ( .A(n874), .B(n873), .Z(n876) );
  XNOR2_X1 U973 ( .A(G2096), .B(G2100), .ZN(n875) );
  XNOR2_X1 U974 ( .A(n876), .B(n875), .ZN(n878) );
  XOR2_X1 U975 ( .A(G2084), .B(G2078), .Z(n877) );
  XNOR2_X1 U976 ( .A(n878), .B(n877), .ZN(G227) );
  NAND2_X1 U977 ( .A1(G100), .A2(n543), .ZN(n880) );
  NAND2_X1 U978 ( .A1(G112), .A2(n908), .ZN(n879) );
  NAND2_X1 U979 ( .A1(n880), .A2(n879), .ZN(n881) );
  XNOR2_X1 U980 ( .A(KEYINPUT110), .B(n881), .ZN(n887) );
  NAND2_X1 U981 ( .A1(G124), .A2(n558), .ZN(n882) );
  XOR2_X1 U982 ( .A(KEYINPUT44), .B(n882), .Z(n883) );
  XNOR2_X1 U983 ( .A(n883), .B(KEYINPUT109), .ZN(n885) );
  NAND2_X1 U984 ( .A1(G136), .A2(n905), .ZN(n884) );
  NAND2_X1 U985 ( .A1(n885), .A2(n884), .ZN(n886) );
  NOR2_X1 U986 ( .A1(n887), .A2(n886), .ZN(G162) );
  NAND2_X1 U987 ( .A1(G106), .A2(n543), .ZN(n889) );
  NAND2_X1 U988 ( .A1(G142), .A2(n905), .ZN(n888) );
  NAND2_X1 U989 ( .A1(n889), .A2(n888), .ZN(n890) );
  XNOR2_X1 U990 ( .A(n890), .B(KEYINPUT45), .ZN(n892) );
  NAND2_X1 U991 ( .A1(G130), .A2(n558), .ZN(n891) );
  NAND2_X1 U992 ( .A1(n892), .A2(n891), .ZN(n895) );
  NAND2_X1 U993 ( .A1(G118), .A2(n908), .ZN(n893) );
  XNOR2_X1 U994 ( .A(KEYINPUT111), .B(n893), .ZN(n894) );
  NOR2_X1 U995 ( .A1(n895), .A2(n894), .ZN(n896) );
  XOR2_X1 U996 ( .A(n932), .B(n896), .Z(n897) );
  XNOR2_X1 U997 ( .A(n898), .B(n897), .ZN(n902) );
  XOR2_X1 U998 ( .A(KEYINPUT46), .B(KEYINPUT112), .Z(n900) );
  XNOR2_X1 U999 ( .A(KEYINPUT114), .B(KEYINPUT48), .ZN(n899) );
  XNOR2_X1 U1000 ( .A(n900), .B(n899), .ZN(n901) );
  XOR2_X1 U1001 ( .A(n902), .B(n901), .Z(n904) );
  XNOR2_X1 U1002 ( .A(G164), .B(G162), .ZN(n903) );
  XNOR2_X1 U1003 ( .A(n904), .B(n903), .ZN(n920) );
  NAND2_X1 U1004 ( .A1(G103), .A2(n543), .ZN(n907) );
  NAND2_X1 U1005 ( .A1(G139), .A2(n905), .ZN(n906) );
  NAND2_X1 U1006 ( .A1(n907), .A2(n906), .ZN(n914) );
  NAND2_X1 U1007 ( .A1(G115), .A2(n908), .ZN(n910) );
  NAND2_X1 U1008 ( .A1(G127), .A2(n558), .ZN(n909) );
  NAND2_X1 U1009 ( .A1(n910), .A2(n909), .ZN(n911) );
  XNOR2_X1 U1010 ( .A(KEYINPUT47), .B(n911), .ZN(n912) );
  XNOR2_X1 U1011 ( .A(KEYINPUT113), .B(n912), .ZN(n913) );
  NOR2_X1 U1012 ( .A1(n914), .A2(n913), .ZN(n937) );
  XNOR2_X1 U1013 ( .A(n937), .B(G160), .ZN(n916) );
  XNOR2_X1 U1014 ( .A(n916), .B(n915), .ZN(n917) );
  XOR2_X1 U1015 ( .A(n918), .B(n917), .Z(n919) );
  XNOR2_X1 U1016 ( .A(n920), .B(n919), .ZN(n921) );
  NOR2_X1 U1017 ( .A1(G37), .A2(n921), .ZN(n922) );
  XOR2_X1 U1018 ( .A(KEYINPUT115), .B(n922), .Z(G395) );
  NOR2_X1 U1019 ( .A1(G401), .A2(n930), .ZN(n927) );
  NOR2_X1 U1020 ( .A1(G229), .A2(G227), .ZN(n924) );
  XNOR2_X1 U1021 ( .A(KEYINPUT116), .B(KEYINPUT49), .ZN(n923) );
  XNOR2_X1 U1022 ( .A(n924), .B(n923), .ZN(n925) );
  NOR2_X1 U1023 ( .A1(G397), .A2(n925), .ZN(n926) );
  NAND2_X1 U1024 ( .A1(n927), .A2(n926), .ZN(n928) );
  NOR2_X1 U1025 ( .A1(n928), .A2(G395), .ZN(n929) );
  XNOR2_X1 U1026 ( .A(n929), .B(KEYINPUT117), .ZN(G225) );
  XOR2_X1 U1027 ( .A(KEYINPUT118), .B(G225), .Z(G308) );
  INV_X1 U1028 ( .A(n930), .ZN(G319) );
  XOR2_X1 U1029 ( .A(G2084), .B(G160), .Z(n931) );
  NOR2_X1 U1030 ( .A1(n932), .A2(n931), .ZN(n933) );
  NAND2_X1 U1031 ( .A1(n934), .A2(n933), .ZN(n935) );
  NOR2_X1 U1032 ( .A1(n936), .A2(n935), .ZN(n949) );
  XOR2_X1 U1033 ( .A(G2072), .B(n937), .Z(n939) );
  XOR2_X1 U1034 ( .A(G164), .B(G2078), .Z(n938) );
  NOR2_X1 U1035 ( .A1(n939), .A2(n938), .ZN(n940) );
  XNOR2_X1 U1036 ( .A(n940), .B(KEYINPUT50), .ZN(n942) );
  NAND2_X1 U1037 ( .A1(n942), .A2(n941), .ZN(n947) );
  XOR2_X1 U1038 ( .A(G2090), .B(G162), .Z(n943) );
  NOR2_X1 U1039 ( .A1(n944), .A2(n943), .ZN(n945) );
  XNOR2_X1 U1040 ( .A(n945), .B(KEYINPUT51), .ZN(n946) );
  NOR2_X1 U1041 ( .A1(n947), .A2(n946), .ZN(n948) );
  NAND2_X1 U1042 ( .A1(n949), .A2(n948), .ZN(n950) );
  NOR2_X1 U1043 ( .A1(n951), .A2(n950), .ZN(n952) );
  XNOR2_X1 U1044 ( .A(KEYINPUT52), .B(n952), .ZN(n953) );
  INV_X1 U1045 ( .A(KEYINPUT55), .ZN(n974) );
  NAND2_X1 U1046 ( .A1(n953), .A2(n974), .ZN(n954) );
  NAND2_X1 U1047 ( .A1(n954), .A2(G29), .ZN(n1035) );
  XNOR2_X1 U1048 ( .A(G2090), .B(G35), .ZN(n969) );
  XNOR2_X1 U1049 ( .A(G2067), .B(G26), .ZN(n956) );
  XNOR2_X1 U1050 ( .A(G33), .B(G2072), .ZN(n955) );
  NOR2_X1 U1051 ( .A1(n956), .A2(n955), .ZN(n960) );
  XOR2_X1 U1052 ( .A(G1991), .B(G25), .Z(n957) );
  NAND2_X1 U1053 ( .A1(n957), .A2(G28), .ZN(n958) );
  XOR2_X1 U1054 ( .A(KEYINPUT120), .B(n958), .Z(n959) );
  NAND2_X1 U1055 ( .A1(n960), .A2(n959), .ZN(n966) );
  XNOR2_X1 U1056 ( .A(G1996), .B(G32), .ZN(n963) );
  XNOR2_X1 U1057 ( .A(n961), .B(G27), .ZN(n962) );
  NOR2_X1 U1058 ( .A1(n963), .A2(n962), .ZN(n964) );
  XNOR2_X1 U1059 ( .A(n964), .B(KEYINPUT121), .ZN(n965) );
  NOR2_X1 U1060 ( .A1(n966), .A2(n965), .ZN(n967) );
  XNOR2_X1 U1061 ( .A(KEYINPUT53), .B(n967), .ZN(n968) );
  NOR2_X1 U1062 ( .A1(n969), .A2(n968), .ZN(n972) );
  XOR2_X1 U1063 ( .A(G2084), .B(KEYINPUT54), .Z(n970) );
  XNOR2_X1 U1064 ( .A(G34), .B(n970), .ZN(n971) );
  NAND2_X1 U1065 ( .A1(n972), .A2(n971), .ZN(n973) );
  XNOR2_X1 U1066 ( .A(n974), .B(n973), .ZN(n976) );
  INV_X1 U1067 ( .A(G29), .ZN(n975) );
  NAND2_X1 U1068 ( .A1(n976), .A2(n975), .ZN(n977) );
  NAND2_X1 U1069 ( .A1(G11), .A2(n977), .ZN(n1033) );
  XNOR2_X1 U1070 ( .A(G16), .B(KEYINPUT56), .ZN(n1003) );
  XNOR2_X1 U1071 ( .A(G1341), .B(n978), .ZN(n984) );
  XOR2_X1 U1072 ( .A(G1348), .B(KEYINPUT123), .Z(n979) );
  XNOR2_X1 U1073 ( .A(n980), .B(n979), .ZN(n982) );
  XOR2_X1 U1074 ( .A(G1961), .B(G171), .Z(n981) );
  NOR2_X1 U1075 ( .A1(n982), .A2(n981), .ZN(n983) );
  NAND2_X1 U1076 ( .A1(n984), .A2(n983), .ZN(n995) );
  XOR2_X1 U1077 ( .A(G299), .B(G1956), .Z(n988) );
  AND2_X1 U1078 ( .A1(G303), .A2(G1971), .ZN(n985) );
  NOR2_X1 U1079 ( .A1(n986), .A2(n985), .ZN(n987) );
  NAND2_X1 U1080 ( .A1(n988), .A2(n987), .ZN(n989) );
  NOR2_X1 U1081 ( .A1(n990), .A2(n989), .ZN(n992) );
  NAND2_X1 U1082 ( .A1(n992), .A2(n991), .ZN(n993) );
  XNOR2_X1 U1083 ( .A(KEYINPUT124), .B(n993), .ZN(n994) );
  NOR2_X1 U1084 ( .A1(n995), .A2(n994), .ZN(n1001) );
  XNOR2_X1 U1085 ( .A(KEYINPUT122), .B(KEYINPUT57), .ZN(n999) );
  XNOR2_X1 U1086 ( .A(G1966), .B(G168), .ZN(n997) );
  NAND2_X1 U1087 ( .A1(n997), .A2(n996), .ZN(n998) );
  XNOR2_X1 U1088 ( .A(n999), .B(n998), .ZN(n1000) );
  NAND2_X1 U1089 ( .A1(n1001), .A2(n1000), .ZN(n1002) );
  NAND2_X1 U1090 ( .A1(n1003), .A2(n1002), .ZN(n1031) );
  INV_X1 U1091 ( .A(G16), .ZN(n1029) );
  XOR2_X1 U1092 ( .A(G1986), .B(G24), .Z(n1005) );
  XOR2_X1 U1093 ( .A(G1971), .B(G22), .Z(n1004) );
  NAND2_X1 U1094 ( .A1(n1005), .A2(n1004), .ZN(n1007) );
  XNOR2_X1 U1095 ( .A(G23), .B(G1976), .ZN(n1006) );
  NOR2_X1 U1096 ( .A1(n1007), .A2(n1006), .ZN(n1008) );
  XOR2_X1 U1097 ( .A(KEYINPUT58), .B(n1008), .Z(n1026) );
  XOR2_X1 U1098 ( .A(G1961), .B(KEYINPUT125), .Z(n1009) );
  XNOR2_X1 U1099 ( .A(G5), .B(n1009), .ZN(n1023) );
  XNOR2_X1 U1100 ( .A(G1348), .B(KEYINPUT59), .ZN(n1010) );
  XNOR2_X1 U1101 ( .A(n1010), .B(G4), .ZN(n1014) );
  XNOR2_X1 U1102 ( .A(G1981), .B(G6), .ZN(n1012) );
  XNOR2_X1 U1103 ( .A(G19), .B(G1341), .ZN(n1011) );
  NOR2_X1 U1104 ( .A1(n1012), .A2(n1011), .ZN(n1013) );
  NAND2_X1 U1105 ( .A1(n1014), .A2(n1013), .ZN(n1017) );
  XNOR2_X1 U1106 ( .A(G20), .B(n1015), .ZN(n1016) );
  NOR2_X1 U1107 ( .A1(n1017), .A2(n1016), .ZN(n1018) );
  XOR2_X1 U1108 ( .A(KEYINPUT60), .B(n1018), .Z(n1020) );
  XNOR2_X1 U1109 ( .A(G1966), .B(G21), .ZN(n1019) );
  NOR2_X1 U1110 ( .A1(n1020), .A2(n1019), .ZN(n1021) );
  XOR2_X1 U1111 ( .A(KEYINPUT126), .B(n1021), .Z(n1022) );
  NOR2_X1 U1112 ( .A1(n1023), .A2(n1022), .ZN(n1024) );
  XNOR2_X1 U1113 ( .A(KEYINPUT127), .B(n1024), .ZN(n1025) );
  NOR2_X1 U1114 ( .A1(n1026), .A2(n1025), .ZN(n1027) );
  XNOR2_X1 U1115 ( .A(KEYINPUT61), .B(n1027), .ZN(n1028) );
  NAND2_X1 U1116 ( .A1(n1029), .A2(n1028), .ZN(n1030) );
  NAND2_X1 U1117 ( .A1(n1031), .A2(n1030), .ZN(n1032) );
  NOR2_X1 U1118 ( .A1(n1033), .A2(n1032), .ZN(n1034) );
  NAND2_X1 U1119 ( .A1(n1035), .A2(n1034), .ZN(n1036) );
  XOR2_X1 U1120 ( .A(KEYINPUT62), .B(n1036), .Z(G311) );
  INV_X1 U1121 ( .A(G311), .ZN(G150) );
endmodule

