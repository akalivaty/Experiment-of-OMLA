//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 0 0 1 0 0 1 0 1 0 1 1 0 1 0 1 0 1 1 0 0 0 1 1 1 1 0 0 1 1 1 0 1 0 1 1 0 0 0 1 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 0 0 1 0 1 1 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:24:58 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n624, new_n625, new_n626, new_n628, new_n629, new_n630,
    new_n631, new_n632, new_n633, new_n634, new_n635, new_n636, new_n637,
    new_n638, new_n639, new_n640, new_n641, new_n643, new_n644, new_n645,
    new_n646, new_n647, new_n648, new_n649, new_n650, new_n651, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n674, new_n675,
    new_n676, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n685, new_n687, new_n688, new_n689, new_n690, new_n691, new_n692,
    new_n693, new_n694, new_n695, new_n696, new_n698, new_n699, new_n700,
    new_n701, new_n702, new_n703, new_n704, new_n706, new_n707, new_n708,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n720, new_n721, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n879, new_n880, new_n881, new_n882, new_n883, new_n884,
    new_n885, new_n886, new_n887, new_n888, new_n889, new_n890, new_n891,
    new_n893, new_n894, new_n895, new_n896, new_n897, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n909, new_n910, new_n911, new_n912, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n935, new_n936, new_n937, new_n938,
    new_n939, new_n940, new_n941, new_n942, new_n943, new_n944;
  INV_X1    g000(.A(G478), .ZN(new_n187));
  NOR2_X1   g001(.A1(new_n187), .A2(KEYINPUT15), .ZN(new_n188));
  INV_X1    g002(.A(G107), .ZN(new_n189));
  INV_X1    g003(.A(G122), .ZN(new_n190));
  NAND2_X1  g004(.A1(new_n190), .A2(G116), .ZN(new_n191));
  AOI21_X1  g005(.A(new_n189), .B1(new_n191), .B2(KEYINPUT14), .ZN(new_n192));
  XNOR2_X1  g006(.A(G116), .B(G122), .ZN(new_n193));
  XNOR2_X1  g007(.A(new_n192), .B(new_n193), .ZN(new_n194));
  INV_X1    g008(.A(KEYINPUT71), .ZN(new_n195));
  INV_X1    g009(.A(G128), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n195), .A2(new_n196), .ZN(new_n197));
  NAND2_X1  g011(.A1(KEYINPUT71), .A2(G128), .ZN(new_n198));
  NAND3_X1  g012(.A1(new_n197), .A2(G143), .A3(new_n198), .ZN(new_n199));
  INV_X1    g013(.A(KEYINPUT95), .ZN(new_n200));
  INV_X1    g014(.A(G143), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n201), .A2(G128), .ZN(new_n202));
  NAND3_X1  g016(.A1(new_n199), .A2(new_n200), .A3(new_n202), .ZN(new_n203));
  INV_X1    g017(.A(new_n203), .ZN(new_n204));
  AOI21_X1  g018(.A(new_n200), .B1(new_n199), .B2(new_n202), .ZN(new_n205));
  NOR3_X1   g019(.A1(new_n204), .A2(new_n205), .A3(G134), .ZN(new_n206));
  INV_X1    g020(.A(G134), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n199), .A2(new_n202), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n208), .A2(KEYINPUT95), .ZN(new_n209));
  AOI21_X1  g023(.A(new_n207), .B1(new_n209), .B2(new_n203), .ZN(new_n210));
  OAI21_X1  g024(.A(new_n194), .B1(new_n206), .B2(new_n210), .ZN(new_n211));
  NAND3_X1  g025(.A1(new_n209), .A2(new_n207), .A3(new_n203), .ZN(new_n212));
  XNOR2_X1  g026(.A(new_n193), .B(new_n189), .ZN(new_n213));
  OR2_X1    g027(.A1(KEYINPUT94), .A2(KEYINPUT13), .ZN(new_n214));
  NAND2_X1  g028(.A1(KEYINPUT94), .A2(KEYINPUT13), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n214), .A2(new_n215), .ZN(new_n216));
  NAND3_X1  g030(.A1(new_n216), .A2(G128), .A3(new_n201), .ZN(new_n217));
  NAND3_X1  g031(.A1(new_n214), .A2(new_n202), .A3(new_n215), .ZN(new_n218));
  AND3_X1   g032(.A1(new_n217), .A2(new_n199), .A3(new_n218), .ZN(new_n219));
  OAI211_X1 g033(.A(new_n212), .B(new_n213), .C1(new_n207), .C2(new_n219), .ZN(new_n220));
  XNOR2_X1  g034(.A(KEYINPUT9), .B(G234), .ZN(new_n221));
  INV_X1    g035(.A(G217), .ZN(new_n222));
  NOR3_X1   g036(.A1(new_n221), .A2(new_n222), .A3(G953), .ZN(new_n223));
  NAND3_X1  g037(.A1(new_n211), .A2(new_n220), .A3(new_n223), .ZN(new_n224));
  NAND2_X1  g038(.A1(new_n224), .A2(KEYINPUT96), .ZN(new_n225));
  INV_X1    g039(.A(KEYINPUT96), .ZN(new_n226));
  NAND4_X1  g040(.A1(new_n211), .A2(new_n220), .A3(new_n226), .A4(new_n223), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n211), .A2(new_n220), .ZN(new_n228));
  INV_X1    g042(.A(new_n223), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n228), .A2(new_n229), .ZN(new_n230));
  NAND3_X1  g044(.A1(new_n225), .A2(new_n227), .A3(new_n230), .ZN(new_n231));
  INV_X1    g045(.A(G902), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n231), .A2(new_n232), .ZN(new_n233));
  INV_X1    g047(.A(KEYINPUT97), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n233), .A2(new_n234), .ZN(new_n235));
  NAND3_X1  g049(.A1(new_n231), .A2(KEYINPUT97), .A3(new_n232), .ZN(new_n236));
  AOI21_X1  g050(.A(new_n188), .B1(new_n235), .B2(new_n236), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n236), .A2(new_n188), .ZN(new_n238));
  INV_X1    g052(.A(new_n238), .ZN(new_n239));
  OAI21_X1  g053(.A(KEYINPUT98), .B1(new_n237), .B2(new_n239), .ZN(new_n240));
  INV_X1    g054(.A(new_n188), .ZN(new_n241));
  AND3_X1   g055(.A1(new_n231), .A2(KEYINPUT97), .A3(new_n232), .ZN(new_n242));
  AOI21_X1  g056(.A(KEYINPUT97), .B1(new_n231), .B2(new_n232), .ZN(new_n243));
  OAI21_X1  g057(.A(new_n241), .B1(new_n242), .B2(new_n243), .ZN(new_n244));
  INV_X1    g058(.A(KEYINPUT98), .ZN(new_n245));
  NAND3_X1  g059(.A1(new_n244), .A2(new_n245), .A3(new_n238), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n240), .A2(new_n246), .ZN(new_n247));
  INV_X1    g061(.A(new_n247), .ZN(new_n248));
  INV_X1    g062(.A(G104), .ZN(new_n249));
  OAI21_X1  g063(.A(KEYINPUT3), .B1(new_n249), .B2(G107), .ZN(new_n250));
  INV_X1    g064(.A(KEYINPUT3), .ZN(new_n251));
  NAND3_X1  g065(.A1(new_n251), .A2(new_n189), .A3(G104), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n249), .A2(G107), .ZN(new_n253));
  NAND3_X1  g067(.A1(new_n250), .A2(new_n252), .A3(new_n253), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n254), .A2(G101), .ZN(new_n255));
  INV_X1    g069(.A(G101), .ZN(new_n256));
  NAND4_X1  g070(.A1(new_n250), .A2(new_n252), .A3(new_n256), .A4(new_n253), .ZN(new_n257));
  NAND3_X1  g071(.A1(new_n255), .A2(KEYINPUT4), .A3(new_n257), .ZN(new_n258));
  INV_X1    g072(.A(new_n258), .ZN(new_n259));
  INV_X1    g073(.A(KEYINPUT4), .ZN(new_n260));
  NAND3_X1  g074(.A1(new_n254), .A2(new_n260), .A3(G101), .ZN(new_n261));
  INV_X1    g075(.A(G146), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n262), .A2(G143), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n201), .A2(G146), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n263), .A2(new_n264), .ZN(new_n265));
  INV_X1    g079(.A(KEYINPUT64), .ZN(new_n266));
  NAND2_X1  g080(.A1(KEYINPUT0), .A2(G128), .ZN(new_n267));
  OR2_X1    g081(.A1(KEYINPUT0), .A2(G128), .ZN(new_n268));
  NAND4_X1  g082(.A1(new_n265), .A2(new_n266), .A3(new_n267), .A4(new_n268), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n268), .A2(new_n267), .ZN(new_n270));
  XNOR2_X1  g084(.A(G143), .B(G146), .ZN(new_n271));
  OAI21_X1  g085(.A(KEYINPUT64), .B1(new_n270), .B2(new_n271), .ZN(new_n272));
  NAND3_X1  g086(.A1(new_n271), .A2(KEYINPUT0), .A3(G128), .ZN(new_n273));
  NAND4_X1  g087(.A1(new_n261), .A2(new_n269), .A3(new_n272), .A4(new_n273), .ZN(new_n274));
  OAI21_X1  g088(.A(KEYINPUT82), .B1(new_n259), .B2(new_n274), .ZN(new_n275));
  NAND3_X1  g089(.A1(new_n272), .A2(new_n269), .A3(new_n273), .ZN(new_n276));
  INV_X1    g090(.A(new_n276), .ZN(new_n277));
  INV_X1    g091(.A(KEYINPUT82), .ZN(new_n278));
  NAND4_X1  g092(.A1(new_n277), .A2(new_n278), .A3(new_n258), .A4(new_n261), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n275), .A2(new_n279), .ZN(new_n280));
  NOR3_X1   g094(.A1(new_n265), .A2(KEYINPUT1), .A3(new_n196), .ZN(new_n281));
  INV_X1    g095(.A(KEYINPUT1), .ZN(new_n282));
  AOI21_X1  g096(.A(new_n282), .B1(G143), .B2(new_n262), .ZN(new_n283));
  INV_X1    g097(.A(KEYINPUT70), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n283), .A2(new_n284), .ZN(new_n285));
  OAI21_X1  g099(.A(KEYINPUT1), .B1(new_n201), .B2(G146), .ZN(new_n286));
  NAND2_X1  g100(.A1(new_n286), .A2(KEYINPUT70), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n197), .A2(new_n198), .ZN(new_n288));
  NAND3_X1  g102(.A1(new_n285), .A2(new_n287), .A3(new_n288), .ZN(new_n289));
  AOI21_X1  g103(.A(new_n281), .B1(new_n289), .B2(new_n265), .ZN(new_n290));
  INV_X1    g104(.A(KEYINPUT10), .ZN(new_n291));
  NOR2_X1   g105(.A1(new_n290), .A2(new_n291), .ZN(new_n292));
  NOR2_X1   g106(.A1(new_n249), .A2(G107), .ZN(new_n293));
  NOR2_X1   g107(.A1(new_n189), .A2(G104), .ZN(new_n294));
  OAI21_X1  g108(.A(G101), .B1(new_n293), .B2(new_n294), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n257), .A2(new_n295), .ZN(new_n296));
  XNOR2_X1  g110(.A(new_n296), .B(KEYINPUT85), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n292), .A2(new_n297), .ZN(new_n298));
  INV_X1    g112(.A(KEYINPUT83), .ZN(new_n299));
  OAI21_X1  g113(.A(G128), .B1(new_n286), .B2(new_n299), .ZN(new_n300));
  NOR2_X1   g114(.A1(new_n283), .A2(KEYINPUT83), .ZN(new_n301));
  OAI21_X1  g115(.A(new_n265), .B1(new_n300), .B2(new_n301), .ZN(new_n302));
  INV_X1    g116(.A(new_n281), .ZN(new_n303));
  AOI21_X1  g117(.A(new_n296), .B1(new_n302), .B2(new_n303), .ZN(new_n304));
  OAI21_X1  g118(.A(KEYINPUT84), .B1(new_n304), .B2(KEYINPUT10), .ZN(new_n305));
  INV_X1    g119(.A(KEYINPUT84), .ZN(new_n306));
  AOI21_X1  g120(.A(new_n196), .B1(new_n283), .B2(KEYINPUT83), .ZN(new_n307));
  OAI21_X1  g121(.A(new_n307), .B1(KEYINPUT83), .B2(new_n283), .ZN(new_n308));
  AOI21_X1  g122(.A(new_n281), .B1(new_n308), .B2(new_n265), .ZN(new_n309));
  OAI211_X1 g123(.A(new_n306), .B(new_n291), .C1(new_n309), .C2(new_n296), .ZN(new_n310));
  NAND4_X1  g124(.A1(new_n280), .A2(new_n298), .A3(new_n305), .A4(new_n310), .ZN(new_n311));
  XNOR2_X1  g125(.A(KEYINPUT67), .B(G131), .ZN(new_n312));
  AND2_X1   g126(.A1(KEYINPUT11), .A2(G134), .ZN(new_n313));
  INV_X1    g127(.A(KEYINPUT11), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n314), .A2(new_n207), .ZN(new_n315));
  INV_X1    g129(.A(G137), .ZN(new_n316));
  AOI21_X1  g130(.A(new_n313), .B1(new_n315), .B2(new_n316), .ZN(new_n317));
  INV_X1    g131(.A(new_n317), .ZN(new_n318));
  XNOR2_X1  g132(.A(KEYINPUT65), .B(G137), .ZN(new_n319));
  AOI21_X1  g133(.A(KEYINPUT66), .B1(new_n319), .B2(new_n313), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n316), .A2(KEYINPUT65), .ZN(new_n321));
  INV_X1    g135(.A(KEYINPUT65), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n322), .A2(G137), .ZN(new_n323));
  AND4_X1   g137(.A1(KEYINPUT66), .A2(new_n321), .A3(new_n323), .A4(new_n313), .ZN(new_n324));
  OAI211_X1 g138(.A(new_n312), .B(new_n318), .C1(new_n320), .C2(new_n324), .ZN(new_n325));
  INV_X1    g139(.A(G131), .ZN(new_n326));
  NAND3_X1  g140(.A1(new_n321), .A2(new_n323), .A3(new_n313), .ZN(new_n327));
  INV_X1    g141(.A(KEYINPUT66), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n327), .A2(new_n328), .ZN(new_n329));
  NAND4_X1  g143(.A1(new_n321), .A2(new_n323), .A3(new_n313), .A4(KEYINPUT66), .ZN(new_n330));
  AOI21_X1  g144(.A(new_n317), .B1(new_n329), .B2(new_n330), .ZN(new_n331));
  OAI21_X1  g145(.A(new_n325), .B1(new_n326), .B2(new_n331), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n311), .A2(new_n332), .ZN(new_n333));
  AOI22_X1  g147(.A1(new_n275), .A2(new_n279), .B1(new_n292), .B2(new_n297), .ZN(new_n334));
  INV_X1    g148(.A(new_n332), .ZN(new_n335));
  NAND4_X1  g149(.A1(new_n334), .A2(new_n335), .A3(new_n305), .A4(new_n310), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n333), .A2(new_n336), .ZN(new_n337));
  XNOR2_X1  g151(.A(G110), .B(G140), .ZN(new_n338));
  INV_X1    g152(.A(G953), .ZN(new_n339));
  AND2_X1   g153(.A1(new_n339), .A2(G227), .ZN(new_n340));
  XNOR2_X1  g154(.A(new_n338), .B(new_n340), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n337), .A2(new_n341), .ZN(new_n342));
  INV_X1    g156(.A(new_n341), .ZN(new_n343));
  NAND3_X1  g157(.A1(new_n336), .A2(KEYINPUT86), .A3(new_n343), .ZN(new_n344));
  AND2_X1   g158(.A1(new_n290), .A2(new_n296), .ZN(new_n345));
  OAI21_X1  g159(.A(new_n332), .B1(new_n345), .B2(new_n304), .ZN(new_n346));
  INV_X1    g160(.A(KEYINPUT12), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n346), .A2(new_n347), .ZN(new_n348));
  OAI211_X1 g162(.A(KEYINPUT12), .B(new_n332), .C1(new_n345), .C2(new_n304), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n348), .A2(new_n349), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n344), .A2(new_n350), .ZN(new_n351));
  AOI21_X1  g165(.A(KEYINPUT86), .B1(new_n336), .B2(new_n343), .ZN(new_n352));
  OAI21_X1  g166(.A(new_n342), .B1(new_n351), .B2(new_n352), .ZN(new_n353));
  INV_X1    g167(.A(G469), .ZN(new_n354));
  NAND3_X1  g168(.A1(new_n353), .A2(new_n354), .A3(new_n232), .ZN(new_n355));
  AOI21_X1  g169(.A(new_n343), .B1(new_n350), .B2(new_n336), .ZN(new_n356));
  AND2_X1   g170(.A1(new_n336), .A2(new_n343), .ZN(new_n357));
  AOI21_X1  g171(.A(new_n356), .B1(new_n333), .B2(new_n357), .ZN(new_n358));
  OAI21_X1  g172(.A(G469), .B1(new_n358), .B2(G902), .ZN(new_n359));
  NAND2_X1  g173(.A1(new_n355), .A2(new_n359), .ZN(new_n360));
  OAI21_X1  g174(.A(G221), .B1(new_n221), .B2(G902), .ZN(new_n361));
  OAI21_X1  g175(.A(G214), .B1(G237), .B2(G902), .ZN(new_n362));
  INV_X1    g176(.A(new_n362), .ZN(new_n363));
  OAI21_X1  g177(.A(G210), .B1(G237), .B2(G902), .ZN(new_n364));
  INV_X1    g178(.A(new_n364), .ZN(new_n365));
  INV_X1    g179(.A(KEYINPUT5), .ZN(new_n366));
  INV_X1    g180(.A(G119), .ZN(new_n367));
  NAND3_X1  g181(.A1(new_n366), .A2(new_n367), .A3(G116), .ZN(new_n368));
  XNOR2_X1  g182(.A(G116), .B(G119), .ZN(new_n369));
  INV_X1    g183(.A(new_n369), .ZN(new_n370));
  OAI211_X1 g184(.A(G113), .B(new_n368), .C1(new_n370), .C2(new_n366), .ZN(new_n371));
  XNOR2_X1  g185(.A(KEYINPUT2), .B(G113), .ZN(new_n372));
  INV_X1    g186(.A(new_n372), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n373), .A2(new_n369), .ZN(new_n374));
  AND2_X1   g188(.A1(new_n371), .A2(new_n374), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n297), .A2(new_n375), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n370), .A2(new_n372), .ZN(new_n377));
  NAND3_X1  g191(.A1(new_n377), .A2(new_n374), .A3(KEYINPUT73), .ZN(new_n378));
  OR3_X1    g192(.A1(new_n373), .A2(KEYINPUT73), .A3(new_n369), .ZN(new_n379));
  NAND4_X1  g193(.A1(new_n378), .A2(new_n258), .A3(new_n379), .A4(new_n261), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n376), .A2(new_n380), .ZN(new_n381));
  XNOR2_X1  g195(.A(G110), .B(G122), .ZN(new_n382));
  INV_X1    g196(.A(new_n382), .ZN(new_n383));
  NAND2_X1  g197(.A1(new_n381), .A2(new_n383), .ZN(new_n384));
  NAND3_X1  g198(.A1(new_n376), .A2(new_n382), .A3(new_n380), .ZN(new_n385));
  NAND3_X1  g199(.A1(new_n384), .A2(KEYINPUT6), .A3(new_n385), .ZN(new_n386));
  INV_X1    g200(.A(G125), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n290), .A2(new_n387), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n276), .A2(G125), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n388), .A2(new_n389), .ZN(new_n390));
  XOR2_X1   g204(.A(KEYINPUT87), .B(G224), .Z(new_n391));
  NOR2_X1   g205(.A1(new_n391), .A2(G953), .ZN(new_n392));
  XNOR2_X1  g206(.A(new_n390), .B(new_n392), .ZN(new_n393));
  INV_X1    g207(.A(KEYINPUT6), .ZN(new_n394));
  NAND3_X1  g208(.A1(new_n381), .A2(new_n394), .A3(new_n383), .ZN(new_n395));
  NAND3_X1  g209(.A1(new_n386), .A2(new_n393), .A3(new_n395), .ZN(new_n396));
  INV_X1    g210(.A(new_n396), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n390), .A2(new_n392), .ZN(new_n398));
  AND2_X1   g212(.A1(new_n375), .A2(new_n296), .ZN(new_n399));
  XNOR2_X1  g213(.A(new_n382), .B(KEYINPUT8), .ZN(new_n400));
  OAI21_X1  g214(.A(new_n400), .B1(new_n375), .B2(new_n296), .ZN(new_n401));
  INV_X1    g215(.A(new_n390), .ZN(new_n402));
  OAI221_X1 g216(.A(new_n398), .B1(new_n399), .B2(new_n401), .C1(new_n402), .C2(KEYINPUT7), .ZN(new_n403));
  INV_X1    g217(.A(new_n392), .ZN(new_n404));
  NAND3_X1  g218(.A1(new_n402), .A2(KEYINPUT7), .A3(new_n404), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n405), .A2(new_n385), .ZN(new_n406));
  OAI21_X1  g220(.A(new_n232), .B1(new_n403), .B2(new_n406), .ZN(new_n407));
  OAI21_X1  g221(.A(new_n365), .B1(new_n397), .B2(new_n407), .ZN(new_n408));
  INV_X1    g222(.A(new_n407), .ZN(new_n409));
  NAND3_X1  g223(.A1(new_n409), .A2(new_n364), .A3(new_n396), .ZN(new_n410));
  AOI21_X1  g224(.A(new_n363), .B1(new_n408), .B2(new_n410), .ZN(new_n411));
  NAND3_X1  g225(.A1(new_n360), .A2(new_n361), .A3(new_n411), .ZN(new_n412));
  XNOR2_X1  g226(.A(G125), .B(G140), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n413), .A2(new_n262), .ZN(new_n414));
  XNOR2_X1  g228(.A(new_n414), .B(KEYINPUT78), .ZN(new_n415));
  OAI21_X1  g229(.A(new_n415), .B1(new_n262), .B2(new_n413), .ZN(new_n416));
  INV_X1    g230(.A(G214), .ZN(new_n417));
  NOR3_X1   g231(.A1(new_n417), .A2(G237), .A3(G953), .ZN(new_n418));
  INV_X1    g232(.A(KEYINPUT88), .ZN(new_n419));
  OAI21_X1  g233(.A(new_n418), .B1(new_n419), .B2(G143), .ZN(new_n420));
  XNOR2_X1  g234(.A(KEYINPUT88), .B(G143), .ZN(new_n421));
  OAI21_X1  g235(.A(new_n420), .B1(new_n418), .B2(new_n421), .ZN(new_n422));
  NAND2_X1  g236(.A1(KEYINPUT18), .A2(G131), .ZN(new_n423));
  XNOR2_X1  g237(.A(new_n422), .B(new_n423), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n416), .A2(new_n424), .ZN(new_n425));
  INV_X1    g239(.A(KEYINPUT91), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n413), .A2(KEYINPUT16), .ZN(new_n427));
  OR3_X1    g241(.A1(new_n387), .A2(KEYINPUT16), .A3(G140), .ZN(new_n428));
  NAND3_X1  g242(.A1(new_n427), .A2(G146), .A3(new_n428), .ZN(new_n429));
  INV_X1    g243(.A(new_n429), .ZN(new_n430));
  AOI21_X1  g244(.A(G146), .B1(new_n427), .B2(new_n428), .ZN(new_n431));
  OAI21_X1  g245(.A(new_n426), .B1(new_n430), .B2(new_n431), .ZN(new_n432));
  INV_X1    g246(.A(new_n431), .ZN(new_n433));
  NAND3_X1  g247(.A1(new_n433), .A2(KEYINPUT91), .A3(new_n429), .ZN(new_n434));
  INV_X1    g248(.A(KEYINPUT17), .ZN(new_n435));
  XOR2_X1   g249(.A(KEYINPUT67), .B(G131), .Z(new_n436));
  NOR2_X1   g250(.A1(new_n421), .A2(new_n418), .ZN(new_n437));
  NAND2_X1  g251(.A1(new_n201), .A2(KEYINPUT88), .ZN(new_n438));
  AND2_X1   g252(.A1(new_n418), .A2(new_n438), .ZN(new_n439));
  OAI21_X1  g253(.A(new_n436), .B1(new_n437), .B2(new_n439), .ZN(new_n440));
  OAI211_X1 g254(.A(new_n432), .B(new_n434), .C1(new_n435), .C2(new_n440), .ZN(new_n441));
  OAI211_X1 g255(.A(new_n420), .B(new_n312), .C1(new_n418), .C2(new_n421), .ZN(new_n442));
  NAND3_X1  g256(.A1(new_n440), .A2(new_n435), .A3(new_n442), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n443), .A2(KEYINPUT92), .ZN(new_n444));
  INV_X1    g258(.A(KEYINPUT92), .ZN(new_n445));
  NAND4_X1  g259(.A1(new_n440), .A2(new_n442), .A3(new_n445), .A4(new_n435), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n444), .A2(new_n446), .ZN(new_n447));
  OAI21_X1  g261(.A(new_n425), .B1(new_n441), .B2(new_n447), .ZN(new_n448));
  XOR2_X1   g262(.A(G113), .B(G122), .Z(new_n449));
  XOR2_X1   g263(.A(KEYINPUT90), .B(G104), .Z(new_n450));
  XOR2_X1   g264(.A(new_n449), .B(new_n450), .Z(new_n451));
  NAND2_X1  g265(.A1(new_n448), .A2(new_n451), .ZN(new_n452));
  XOR2_X1   g266(.A(new_n413), .B(KEYINPUT19), .Z(new_n453));
  OAI21_X1  g267(.A(new_n429), .B1(new_n453), .B2(G146), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n454), .A2(KEYINPUT89), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n440), .A2(new_n442), .ZN(new_n456));
  INV_X1    g270(.A(KEYINPUT89), .ZN(new_n457));
  OAI211_X1 g271(.A(new_n429), .B(new_n457), .C1(new_n453), .C2(G146), .ZN(new_n458));
  NAND3_X1  g272(.A1(new_n455), .A2(new_n456), .A3(new_n458), .ZN(new_n459));
  AOI21_X1  g273(.A(new_n451), .B1(new_n416), .B2(new_n424), .ZN(new_n460));
  NAND2_X1  g274(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  NOR2_X1   g275(.A1(G475), .A2(G902), .ZN(new_n462));
  NAND3_X1  g276(.A1(new_n452), .A2(new_n461), .A3(new_n462), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n463), .A2(KEYINPUT20), .ZN(new_n464));
  AOI22_X1  g278(.A1(new_n448), .A2(new_n451), .B1(new_n459), .B2(new_n460), .ZN(new_n465));
  INV_X1    g279(.A(KEYINPUT20), .ZN(new_n466));
  NAND3_X1  g280(.A1(new_n465), .A2(new_n466), .A3(new_n462), .ZN(new_n467));
  NAND2_X1  g281(.A1(new_n464), .A2(new_n467), .ZN(new_n468));
  INV_X1    g282(.A(new_n451), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n469), .A2(KEYINPUT93), .ZN(new_n470));
  AND2_X1   g284(.A1(new_n448), .A2(new_n470), .ZN(new_n471));
  OAI21_X1  g285(.A(new_n232), .B1(new_n448), .B2(new_n470), .ZN(new_n472));
  OAI21_X1  g286(.A(G475), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n468), .A2(new_n473), .ZN(new_n474));
  INV_X1    g288(.A(new_n474), .ZN(new_n475));
  NAND2_X1  g289(.A1(G234), .A2(G237), .ZN(new_n476));
  AND3_X1   g290(.A1(new_n476), .A2(G952), .A3(new_n339), .ZN(new_n477));
  AND3_X1   g291(.A1(new_n476), .A2(G902), .A3(G953), .ZN(new_n478));
  XNOR2_X1  g292(.A(KEYINPUT21), .B(G898), .ZN(new_n479));
  AOI21_X1  g293(.A(new_n477), .B1(new_n478), .B2(new_n479), .ZN(new_n480));
  INV_X1    g294(.A(new_n480), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n475), .A2(new_n481), .ZN(new_n482));
  NOR3_X1   g296(.A1(new_n248), .A2(new_n412), .A3(new_n482), .ZN(new_n483));
  AOI211_X1 g297(.A(new_n436), .B(new_n317), .C1(new_n329), .C2(new_n330), .ZN(new_n484));
  NOR2_X1   g298(.A1(new_n207), .A2(G137), .ZN(new_n485));
  XNOR2_X1  g299(.A(new_n485), .B(KEYINPUT69), .ZN(new_n486));
  OR2_X1    g300(.A1(new_n319), .A2(G134), .ZN(new_n487));
  AOI21_X1  g301(.A(new_n326), .B1(new_n486), .B2(new_n487), .ZN(new_n488));
  OR3_X1    g302(.A1(new_n484), .A2(new_n290), .A3(new_n488), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n329), .A2(new_n330), .ZN(new_n490));
  AOI21_X1  g304(.A(new_n326), .B1(new_n490), .B2(new_n318), .ZN(new_n491));
  OAI21_X1  g305(.A(new_n277), .B1(new_n491), .B2(new_n484), .ZN(new_n492));
  NAND3_X1  g306(.A1(new_n489), .A2(KEYINPUT30), .A3(new_n492), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n378), .A2(new_n379), .ZN(new_n494));
  INV_X1    g308(.A(new_n494), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n493), .A2(new_n495), .ZN(new_n496));
  INV_X1    g310(.A(KEYINPUT72), .ZN(new_n497));
  NOR3_X1   g311(.A1(new_n484), .A2(new_n290), .A3(new_n488), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n492), .A2(KEYINPUT68), .ZN(new_n499));
  INV_X1    g313(.A(KEYINPUT68), .ZN(new_n500));
  NAND3_X1  g314(.A1(new_n332), .A2(new_n500), .A3(new_n277), .ZN(new_n501));
  AOI21_X1  g315(.A(new_n498), .B1(new_n499), .B2(new_n501), .ZN(new_n502));
  OAI21_X1  g316(.A(new_n497), .B1(new_n502), .B2(KEYINPUT30), .ZN(new_n503));
  OAI21_X1  g317(.A(new_n318), .B1(new_n320), .B2(new_n324), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n504), .A2(G131), .ZN(new_n505));
  AOI211_X1 g319(.A(KEYINPUT68), .B(new_n276), .C1(new_n505), .C2(new_n325), .ZN(new_n506));
  AOI21_X1  g320(.A(new_n500), .B1(new_n332), .B2(new_n277), .ZN(new_n507));
  OAI21_X1  g321(.A(new_n489), .B1(new_n506), .B2(new_n507), .ZN(new_n508));
  INV_X1    g322(.A(KEYINPUT30), .ZN(new_n509));
  NAND3_X1  g323(.A1(new_n508), .A2(KEYINPUT72), .A3(new_n509), .ZN(new_n510));
  AOI21_X1  g324(.A(new_n496), .B1(new_n503), .B2(new_n510), .ZN(new_n511));
  NAND3_X1  g325(.A1(new_n489), .A2(new_n492), .A3(new_n494), .ZN(new_n512));
  INV_X1    g326(.A(new_n512), .ZN(new_n513));
  INV_X1    g327(.A(G237), .ZN(new_n514));
  NAND3_X1  g328(.A1(new_n514), .A2(new_n339), .A3(G210), .ZN(new_n515));
  XNOR2_X1  g329(.A(new_n515), .B(KEYINPUT27), .ZN(new_n516));
  XNOR2_X1  g330(.A(KEYINPUT26), .B(G101), .ZN(new_n517));
  XNOR2_X1  g331(.A(new_n516), .B(new_n517), .ZN(new_n518));
  INV_X1    g332(.A(new_n518), .ZN(new_n519));
  NOR2_X1   g333(.A1(new_n513), .A2(new_n519), .ZN(new_n520));
  INV_X1    g334(.A(new_n520), .ZN(new_n521));
  OAI21_X1  g335(.A(KEYINPUT31), .B1(new_n511), .B2(new_n521), .ZN(new_n522));
  INV_X1    g336(.A(new_n496), .ZN(new_n523));
  NOR3_X1   g337(.A1(new_n502), .A2(new_n497), .A3(KEYINPUT30), .ZN(new_n524));
  AOI21_X1  g338(.A(KEYINPUT72), .B1(new_n508), .B2(new_n509), .ZN(new_n525));
  OAI21_X1  g339(.A(new_n523), .B1(new_n524), .B2(new_n525), .ZN(new_n526));
  INV_X1    g340(.A(KEYINPUT31), .ZN(new_n527));
  NAND3_X1  g341(.A1(new_n526), .A2(new_n527), .A3(new_n520), .ZN(new_n528));
  NOR2_X1   g342(.A1(new_n513), .A2(KEYINPUT28), .ZN(new_n529));
  OAI21_X1  g343(.A(KEYINPUT74), .B1(new_n502), .B2(new_n494), .ZN(new_n530));
  INV_X1    g344(.A(KEYINPUT74), .ZN(new_n531));
  NAND3_X1  g345(.A1(new_n508), .A2(new_n531), .A3(new_n495), .ZN(new_n532));
  NAND3_X1  g346(.A1(new_n530), .A2(new_n512), .A3(new_n532), .ZN(new_n533));
  AOI21_X1  g347(.A(new_n529), .B1(new_n533), .B2(KEYINPUT28), .ZN(new_n534));
  OAI211_X1 g348(.A(new_n522), .B(new_n528), .C1(new_n534), .C2(new_n518), .ZN(new_n535));
  INV_X1    g349(.A(KEYINPUT32), .ZN(new_n536));
  NOR2_X1   g350(.A1(G472), .A2(G902), .ZN(new_n537));
  AND3_X1   g351(.A1(new_n535), .A2(new_n536), .A3(new_n537), .ZN(new_n538));
  AOI21_X1  g352(.A(new_n536), .B1(new_n535), .B2(new_n537), .ZN(new_n539));
  INV_X1    g353(.A(KEYINPUT75), .ZN(new_n540));
  INV_X1    g354(.A(KEYINPUT28), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n489), .A2(new_n492), .ZN(new_n542));
  NAND2_X1  g356(.A1(new_n542), .A2(new_n495), .ZN(new_n543));
  AOI21_X1  g357(.A(new_n541), .B1(new_n543), .B2(new_n512), .ZN(new_n544));
  NOR2_X1   g358(.A1(new_n544), .A2(new_n529), .ZN(new_n545));
  NAND2_X1  g359(.A1(new_n518), .A2(KEYINPUT29), .ZN(new_n546));
  INV_X1    g360(.A(new_n546), .ZN(new_n547));
  AOI21_X1  g361(.A(new_n540), .B1(new_n545), .B2(new_n547), .ZN(new_n548));
  NOR4_X1   g362(.A1(new_n544), .A2(new_n529), .A3(KEYINPUT75), .A4(new_n546), .ZN(new_n549));
  OAI21_X1  g363(.A(new_n232), .B1(new_n548), .B2(new_n549), .ZN(new_n550));
  INV_X1    g364(.A(KEYINPUT29), .ZN(new_n551));
  NAND3_X1  g365(.A1(new_n526), .A2(new_n512), .A3(new_n519), .ZN(new_n552));
  OAI21_X1  g366(.A(new_n552), .B1(new_n534), .B2(new_n519), .ZN(new_n553));
  AOI21_X1  g367(.A(new_n550), .B1(new_n551), .B2(new_n553), .ZN(new_n554));
  INV_X1    g368(.A(G472), .ZN(new_n555));
  OAI22_X1  g369(.A1(new_n538), .A2(new_n539), .B1(new_n554), .B2(new_n555), .ZN(new_n556));
  XNOR2_X1  g370(.A(KEYINPUT24), .B(G110), .ZN(new_n557));
  XNOR2_X1  g371(.A(new_n557), .B(KEYINPUT76), .ZN(new_n558));
  NAND3_X1  g372(.A1(new_n197), .A2(G119), .A3(new_n198), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n367), .A2(G128), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n559), .A2(new_n560), .ZN(new_n561));
  INV_X1    g375(.A(KEYINPUT77), .ZN(new_n562));
  NAND3_X1  g376(.A1(new_n558), .A2(new_n561), .A3(new_n562), .ZN(new_n563));
  INV_X1    g377(.A(KEYINPUT23), .ZN(new_n564));
  OAI21_X1  g378(.A(new_n564), .B1(new_n367), .B2(G128), .ZN(new_n565));
  OAI211_X1 g379(.A(new_n565), .B(new_n560), .C1(new_n559), .C2(new_n564), .ZN(new_n566));
  OAI21_X1  g380(.A(new_n563), .B1(G110), .B2(new_n566), .ZN(new_n567));
  AOI21_X1  g381(.A(new_n562), .B1(new_n558), .B2(new_n561), .ZN(new_n568));
  OAI211_X1 g382(.A(new_n429), .B(new_n415), .C1(new_n567), .C2(new_n568), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n566), .A2(G110), .ZN(new_n570));
  OAI221_X1 g384(.A(new_n570), .B1(new_n558), .B2(new_n561), .C1(new_n430), .C2(new_n431), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n569), .A2(new_n571), .ZN(new_n572));
  XNOR2_X1  g386(.A(KEYINPUT22), .B(G137), .ZN(new_n573));
  NAND3_X1  g387(.A1(new_n339), .A2(G221), .A3(G234), .ZN(new_n574));
  XNOR2_X1  g388(.A(new_n573), .B(new_n574), .ZN(new_n575));
  XOR2_X1   g389(.A(new_n575), .B(KEYINPUT79), .Z(new_n576));
  INV_X1    g390(.A(new_n576), .ZN(new_n577));
  NAND2_X1  g391(.A1(new_n572), .A2(new_n577), .ZN(new_n578));
  NAND3_X1  g392(.A1(new_n569), .A2(new_n571), .A3(new_n575), .ZN(new_n579));
  INV_X1    g393(.A(KEYINPUT80), .ZN(new_n580));
  INV_X1    g394(.A(KEYINPUT25), .ZN(new_n581));
  AOI21_X1  g395(.A(G902), .B1(new_n580), .B2(new_n581), .ZN(new_n582));
  NAND3_X1  g396(.A1(new_n578), .A2(new_n579), .A3(new_n582), .ZN(new_n583));
  NOR2_X1   g397(.A1(new_n580), .A2(new_n581), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  INV_X1    g399(.A(new_n584), .ZN(new_n586));
  NAND4_X1  g400(.A1(new_n578), .A2(new_n586), .A3(new_n579), .A4(new_n582), .ZN(new_n587));
  AOI21_X1  g401(.A(new_n222), .B1(G234), .B2(new_n232), .ZN(new_n588));
  NAND3_X1  g402(.A1(new_n585), .A2(new_n587), .A3(new_n588), .ZN(new_n589));
  NAND2_X1  g403(.A1(new_n589), .A2(KEYINPUT81), .ZN(new_n590));
  INV_X1    g404(.A(KEYINPUT81), .ZN(new_n591));
  NAND4_X1  g405(.A1(new_n585), .A2(new_n591), .A3(new_n587), .A4(new_n588), .ZN(new_n592));
  AND2_X1   g406(.A1(new_n578), .A2(new_n579), .ZN(new_n593));
  NOR2_X1   g407(.A1(new_n588), .A2(G902), .ZN(new_n594));
  NAND2_X1  g408(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  AND3_X1   g409(.A1(new_n590), .A2(new_n592), .A3(new_n595), .ZN(new_n596));
  NAND3_X1  g410(.A1(new_n483), .A2(new_n556), .A3(new_n596), .ZN(new_n597));
  XNOR2_X1  g411(.A(KEYINPUT99), .B(G101), .ZN(new_n598));
  XNOR2_X1  g412(.A(new_n597), .B(new_n598), .ZN(G3));
  NAND2_X1  g413(.A1(new_n411), .A2(new_n481), .ZN(new_n600));
  INV_X1    g414(.A(new_n600), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n233), .A2(new_n187), .ZN(new_n602));
  INV_X1    g416(.A(KEYINPUT33), .ZN(new_n603));
  NAND2_X1  g417(.A1(new_n231), .A2(new_n603), .ZN(new_n604));
  NAND3_X1  g418(.A1(new_n230), .A2(KEYINPUT33), .A3(new_n224), .ZN(new_n605));
  NAND2_X1  g419(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  NOR2_X1   g420(.A1(new_n187), .A2(G902), .ZN(new_n607));
  INV_X1    g421(.A(new_n607), .ZN(new_n608));
  OAI21_X1  g422(.A(new_n602), .B1(new_n606), .B2(new_n608), .ZN(new_n609));
  AND2_X1   g423(.A1(new_n474), .A2(new_n609), .ZN(new_n610));
  NAND3_X1  g424(.A1(new_n601), .A2(KEYINPUT100), .A3(new_n610), .ZN(new_n611));
  INV_X1    g425(.A(KEYINPUT100), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n474), .A2(new_n609), .ZN(new_n613));
  OAI21_X1  g427(.A(new_n612), .B1(new_n600), .B2(new_n613), .ZN(new_n614));
  NAND2_X1  g428(.A1(new_n611), .A2(new_n614), .ZN(new_n615));
  AOI21_X1  g429(.A(new_n555), .B1(new_n535), .B2(new_n232), .ZN(new_n616));
  AOI21_X1  g430(.A(new_n616), .B1(new_n537), .B2(new_n535), .ZN(new_n617));
  INV_X1    g431(.A(new_n596), .ZN(new_n618));
  NAND2_X1  g432(.A1(new_n360), .A2(new_n361), .ZN(new_n619));
  NOR2_X1   g433(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  NAND3_X1  g434(.A1(new_n615), .A2(new_n617), .A3(new_n620), .ZN(new_n621));
  XOR2_X1   g435(.A(KEYINPUT34), .B(G104), .Z(new_n622));
  XNOR2_X1  g436(.A(new_n621), .B(new_n622), .ZN(G6));
  NOR3_X1   g437(.A1(new_n247), .A2(new_n600), .A3(new_n474), .ZN(new_n624));
  NAND3_X1  g438(.A1(new_n617), .A2(new_n620), .A3(new_n624), .ZN(new_n625));
  XOR2_X1   g439(.A(KEYINPUT35), .B(G107), .Z(new_n626));
  XNOR2_X1  g440(.A(new_n625), .B(new_n626), .ZN(G9));
  NAND2_X1  g441(.A1(new_n535), .A2(new_n232), .ZN(new_n628));
  NAND2_X1  g442(.A1(new_n628), .A2(G472), .ZN(new_n629));
  NAND2_X1  g443(.A1(new_n535), .A2(new_n537), .ZN(new_n630));
  NOR2_X1   g444(.A1(new_n577), .A2(KEYINPUT36), .ZN(new_n631));
  XNOR2_X1  g445(.A(new_n572), .B(new_n631), .ZN(new_n632));
  NAND2_X1  g446(.A1(new_n632), .A2(new_n594), .ZN(new_n633));
  NAND3_X1  g447(.A1(new_n590), .A2(new_n592), .A3(new_n633), .ZN(new_n634));
  NAND3_X1  g448(.A1(new_n629), .A2(new_n630), .A3(new_n634), .ZN(new_n635));
  INV_X1    g449(.A(KEYINPUT101), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n635), .A2(new_n636), .ZN(new_n637));
  NAND4_X1  g451(.A1(new_n629), .A2(KEYINPUT101), .A3(new_n630), .A4(new_n634), .ZN(new_n638));
  NAND3_X1  g452(.A1(new_n637), .A2(new_n483), .A3(new_n638), .ZN(new_n639));
  XNOR2_X1  g453(.A(new_n639), .B(KEYINPUT102), .ZN(new_n640));
  XNOR2_X1  g454(.A(KEYINPUT37), .B(G110), .ZN(new_n641));
  XNOR2_X1  g455(.A(new_n640), .B(new_n641), .ZN(G12));
  NAND2_X1  g456(.A1(new_n556), .A2(new_n634), .ZN(new_n643));
  INV_X1    g457(.A(new_n643), .ZN(new_n644));
  INV_X1    g458(.A(G900), .ZN(new_n645));
  AOI21_X1  g459(.A(new_n477), .B1(new_n478), .B2(new_n645), .ZN(new_n646));
  INV_X1    g460(.A(new_n646), .ZN(new_n647));
  NAND4_X1  g461(.A1(new_n240), .A2(new_n475), .A3(new_n246), .A4(new_n647), .ZN(new_n648));
  NOR2_X1   g462(.A1(new_n412), .A2(new_n648), .ZN(new_n649));
  NAND2_X1  g463(.A1(new_n644), .A2(new_n649), .ZN(new_n650));
  XOR2_X1   g464(.A(KEYINPUT103), .B(G128), .Z(new_n651));
  XNOR2_X1  g465(.A(new_n650), .B(new_n651), .ZN(G30));
  AOI21_X1  g466(.A(new_n519), .B1(new_n526), .B2(new_n512), .ZN(new_n653));
  NAND3_X1  g467(.A1(new_n543), .A2(new_n512), .A3(new_n519), .ZN(new_n654));
  NAND2_X1  g468(.A1(new_n654), .A2(new_n232), .ZN(new_n655));
  OAI21_X1  g469(.A(G472), .B1(new_n653), .B2(new_n655), .ZN(new_n656));
  OAI21_X1  g470(.A(new_n656), .B1(new_n538), .B2(new_n539), .ZN(new_n657));
  INV_X1    g471(.A(new_n657), .ZN(new_n658));
  INV_X1    g472(.A(new_n634), .ZN(new_n659));
  AOI21_X1  g473(.A(new_n363), .B1(new_n468), .B2(new_n473), .ZN(new_n660));
  NAND3_X1  g474(.A1(new_n248), .A2(new_n659), .A3(new_n660), .ZN(new_n661));
  AOI21_X1  g475(.A(new_n658), .B1(new_n661), .B2(KEYINPUT104), .ZN(new_n662));
  INV_X1    g476(.A(new_n361), .ZN(new_n663));
  AOI21_X1  g477(.A(new_n663), .B1(new_n355), .B2(new_n359), .ZN(new_n664));
  XOR2_X1   g478(.A(new_n646), .B(KEYINPUT39), .Z(new_n665));
  NAND2_X1  g479(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  XOR2_X1   g480(.A(new_n666), .B(KEYINPUT40), .Z(new_n667));
  NOR2_X1   g481(.A1(new_n661), .A2(KEYINPUT104), .ZN(new_n668));
  NAND2_X1  g482(.A1(new_n408), .A2(new_n410), .ZN(new_n669));
  XOR2_X1   g483(.A(new_n669), .B(KEYINPUT38), .Z(new_n670));
  NOR2_X1   g484(.A1(new_n668), .A2(new_n670), .ZN(new_n671));
  NAND3_X1  g485(.A1(new_n662), .A2(new_n667), .A3(new_n671), .ZN(new_n672));
  XNOR2_X1  g486(.A(new_n672), .B(G143), .ZN(G45));
  NAND2_X1  g487(.A1(new_n610), .A2(new_n647), .ZN(new_n674));
  NOR2_X1   g488(.A1(new_n412), .A2(new_n674), .ZN(new_n675));
  NAND2_X1  g489(.A1(new_n644), .A2(new_n675), .ZN(new_n676));
  XNOR2_X1  g490(.A(new_n676), .B(G146), .ZN(G48));
  NAND2_X1  g491(.A1(new_n353), .A2(new_n232), .ZN(new_n678));
  NAND2_X1  g492(.A1(new_n678), .A2(G469), .ZN(new_n679));
  NAND2_X1  g493(.A1(new_n679), .A2(new_n355), .ZN(new_n680));
  NOR2_X1   g494(.A1(new_n680), .A2(new_n663), .ZN(new_n681));
  NAND4_X1  g495(.A1(new_n615), .A2(new_n556), .A3(new_n596), .A4(new_n681), .ZN(new_n682));
  XNOR2_X1  g496(.A(KEYINPUT41), .B(G113), .ZN(new_n683));
  XNOR2_X1  g497(.A(new_n682), .B(new_n683), .ZN(G15));
  NAND4_X1  g498(.A1(new_n556), .A2(new_n624), .A3(new_n596), .A4(new_n681), .ZN(new_n685));
  XNOR2_X1  g499(.A(new_n685), .B(G116), .ZN(G18));
  AND3_X1   g500(.A1(new_n353), .A2(new_n354), .A3(new_n232), .ZN(new_n687));
  AOI21_X1  g501(.A(new_n354), .B1(new_n353), .B2(new_n232), .ZN(new_n688));
  NOR2_X1   g502(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  INV_X1    g503(.A(KEYINPUT105), .ZN(new_n690));
  NAND4_X1  g504(.A1(new_n689), .A2(new_n690), .A3(new_n361), .A4(new_n411), .ZN(new_n691));
  NAND4_X1  g505(.A1(new_n679), .A2(new_n411), .A3(new_n361), .A4(new_n355), .ZN(new_n692));
  NAND2_X1  g506(.A1(new_n692), .A2(KEYINPUT105), .ZN(new_n693));
  NAND2_X1  g507(.A1(new_n691), .A2(new_n693), .ZN(new_n694));
  NOR2_X1   g508(.A1(new_n248), .A2(new_n482), .ZN(new_n695));
  NAND4_X1  g509(.A1(new_n694), .A2(new_n556), .A3(new_n695), .A4(new_n634), .ZN(new_n696));
  XNOR2_X1  g510(.A(new_n696), .B(G119), .ZN(G21));
  NAND4_X1  g511(.A1(new_n240), .A2(new_n669), .A3(new_n246), .A4(new_n660), .ZN(new_n698));
  INV_X1    g512(.A(KEYINPUT106), .ZN(new_n699));
  XNOR2_X1  g513(.A(new_n698), .B(new_n699), .ZN(new_n700));
  OAI211_X1 g514(.A(new_n522), .B(new_n528), .C1(new_n518), .C2(new_n545), .ZN(new_n701));
  AND2_X1   g515(.A1(new_n701), .A2(new_n537), .ZN(new_n702));
  NOR3_X1   g516(.A1(new_n618), .A2(new_n702), .A3(new_n616), .ZN(new_n703));
  NAND4_X1  g517(.A1(new_n700), .A2(new_n481), .A3(new_n681), .A4(new_n703), .ZN(new_n704));
  XNOR2_X1  g518(.A(new_n704), .B(G122), .ZN(G24));
  NOR3_X1   g519(.A1(new_n702), .A2(new_n616), .A3(new_n659), .ZN(new_n706));
  INV_X1    g520(.A(new_n674), .ZN(new_n707));
  NAND3_X1  g521(.A1(new_n694), .A2(new_n706), .A3(new_n707), .ZN(new_n708));
  XNOR2_X1  g522(.A(new_n708), .B(G125), .ZN(G27));
  NOR2_X1   g523(.A1(new_n669), .A2(new_n363), .ZN(new_n710));
  AND2_X1   g524(.A1(new_n664), .A2(new_n710), .ZN(new_n711));
  NAND4_X1  g525(.A1(new_n556), .A2(new_n596), .A3(new_n707), .A4(new_n711), .ZN(new_n712));
  XNOR2_X1  g526(.A(KEYINPUT107), .B(KEYINPUT42), .ZN(new_n713));
  INV_X1    g527(.A(new_n713), .ZN(new_n714));
  NAND2_X1  g528(.A1(new_n712), .A2(new_n714), .ZN(new_n715));
  INV_X1    g529(.A(KEYINPUT107), .ZN(new_n716));
  NOR2_X1   g530(.A1(new_n716), .A2(KEYINPUT42), .ZN(new_n717));
  OAI21_X1  g531(.A(new_n715), .B1(new_n712), .B2(new_n717), .ZN(new_n718));
  XNOR2_X1  g532(.A(new_n718), .B(G131), .ZN(G33));
  INV_X1    g533(.A(new_n648), .ZN(new_n720));
  AND4_X1   g534(.A1(new_n556), .A2(new_n720), .A3(new_n596), .A4(new_n711), .ZN(new_n721));
  XNOR2_X1  g535(.A(new_n721), .B(new_n207), .ZN(G36));
  AND3_X1   g536(.A1(new_n609), .A2(new_n473), .A3(new_n468), .ZN(new_n723));
  OAI21_X1  g537(.A(new_n723), .B1(KEYINPUT108), .B2(KEYINPUT43), .ZN(new_n724));
  XOR2_X1   g538(.A(KEYINPUT108), .B(KEYINPUT43), .Z(new_n725));
  OAI21_X1  g539(.A(new_n724), .B1(new_n723), .B2(new_n725), .ZN(new_n726));
  NOR2_X1   g540(.A1(new_n617), .A2(new_n659), .ZN(new_n727));
  NAND2_X1  g541(.A1(new_n727), .A2(KEYINPUT109), .ZN(new_n728));
  INV_X1    g542(.A(new_n728), .ZN(new_n729));
  NOR2_X1   g543(.A1(new_n727), .A2(KEYINPUT109), .ZN(new_n730));
  OAI21_X1  g544(.A(new_n726), .B1(new_n729), .B2(new_n730), .ZN(new_n731));
  INV_X1    g545(.A(KEYINPUT44), .ZN(new_n732));
  NAND2_X1  g546(.A1(new_n731), .A2(new_n732), .ZN(new_n733));
  OR2_X1    g547(.A1(new_n358), .A2(KEYINPUT45), .ZN(new_n734));
  NAND2_X1  g548(.A1(new_n358), .A2(KEYINPUT45), .ZN(new_n735));
  NAND3_X1  g549(.A1(new_n734), .A2(G469), .A3(new_n735), .ZN(new_n736));
  NAND2_X1  g550(.A1(G469), .A2(G902), .ZN(new_n737));
  AOI21_X1  g551(.A(KEYINPUT46), .B1(new_n736), .B2(new_n737), .ZN(new_n738));
  NOR2_X1   g552(.A1(new_n738), .A2(new_n687), .ZN(new_n739));
  NAND3_X1  g553(.A1(new_n736), .A2(KEYINPUT46), .A3(new_n737), .ZN(new_n740));
  AOI21_X1  g554(.A(new_n663), .B1(new_n739), .B2(new_n740), .ZN(new_n741));
  NAND4_X1  g555(.A1(new_n733), .A2(new_n665), .A3(new_n710), .A4(new_n741), .ZN(new_n742));
  NOR2_X1   g556(.A1(new_n731), .A2(new_n732), .ZN(new_n743));
  NOR2_X1   g557(.A1(new_n742), .A2(new_n743), .ZN(new_n744));
  XNOR2_X1  g558(.A(new_n744), .B(new_n316), .ZN(G39));
  AND2_X1   g559(.A1(KEYINPUT110), .A2(KEYINPUT47), .ZN(new_n746));
  NOR2_X1   g560(.A1(KEYINPUT110), .A2(KEYINPUT47), .ZN(new_n747));
  NOR2_X1   g561(.A1(new_n746), .A2(new_n747), .ZN(new_n748));
  MUX2_X1   g562(.A(new_n748), .B(new_n746), .S(new_n741), .Z(new_n749));
  NAND3_X1  g563(.A1(new_n707), .A2(new_n618), .A3(new_n710), .ZN(new_n750));
  NOR2_X1   g564(.A1(new_n556), .A2(new_n750), .ZN(new_n751));
  NAND2_X1  g565(.A1(new_n749), .A2(new_n751), .ZN(new_n752));
  XNOR2_X1  g566(.A(new_n752), .B(G140), .ZN(G42));
  NOR2_X1   g567(.A1(new_n663), .A2(new_n363), .ZN(new_n754));
  NAND4_X1  g568(.A1(new_n670), .A2(new_n596), .A3(new_n723), .A4(new_n754), .ZN(new_n755));
  AOI21_X1  g569(.A(new_n755), .B1(KEYINPUT49), .B2(new_n680), .ZN(new_n756));
  NOR2_X1   g570(.A1(new_n680), .A2(KEYINPUT49), .ZN(new_n757));
  XNOR2_X1  g571(.A(new_n757), .B(KEYINPUT111), .ZN(new_n758));
  NAND3_X1  g572(.A1(new_n756), .A2(new_n658), .A3(new_n758), .ZN(new_n759));
  INV_X1    g573(.A(KEYINPUT113), .ZN(new_n760));
  NOR3_X1   g574(.A1(new_n619), .A2(new_n634), .A3(new_n646), .ZN(new_n761));
  NAND2_X1  g575(.A1(new_n657), .A2(new_n761), .ZN(new_n762));
  XNOR2_X1  g576(.A(new_n698), .B(KEYINPUT106), .ZN(new_n763));
  OAI21_X1  g577(.A(new_n760), .B1(new_n762), .B2(new_n763), .ZN(new_n764));
  NAND4_X1  g578(.A1(new_n700), .A2(KEYINPUT113), .A3(new_n657), .A4(new_n761), .ZN(new_n765));
  NAND2_X1  g579(.A1(new_n764), .A2(new_n765), .ZN(new_n766));
  OAI211_X1 g580(.A(new_n556), .B(new_n634), .C1(new_n675), .C2(new_n649), .ZN(new_n767));
  AND2_X1   g581(.A1(new_n767), .A2(new_n708), .ZN(new_n768));
  NAND2_X1  g582(.A1(new_n766), .A2(new_n768), .ZN(new_n769));
  INV_X1    g583(.A(KEYINPUT52), .ZN(new_n770));
  NAND2_X1  g584(.A1(new_n769), .A2(new_n770), .ZN(new_n771));
  INV_X1    g585(.A(KEYINPUT114), .ZN(new_n772));
  NAND3_X1  g586(.A1(new_n766), .A2(new_n768), .A3(KEYINPUT52), .ZN(new_n773));
  NAND3_X1  g587(.A1(new_n771), .A2(new_n772), .A3(new_n773), .ZN(new_n774));
  NAND4_X1  g588(.A1(new_n639), .A2(new_n682), .A3(new_n696), .A4(new_n685), .ZN(new_n775));
  INV_X1    g589(.A(new_n775), .ZN(new_n776));
  NOR2_X1   g590(.A1(new_n237), .A2(new_n239), .ZN(new_n777));
  OAI21_X1  g591(.A(new_n613), .B1(new_n777), .B2(new_n474), .ZN(new_n778));
  NAND4_X1  g592(.A1(new_n617), .A2(new_n620), .A3(new_n601), .A4(new_n778), .ZN(new_n779));
  NAND3_X1  g593(.A1(new_n704), .A2(new_n779), .A3(new_n597), .ZN(new_n780));
  INV_X1    g594(.A(new_n780), .ZN(new_n781));
  NAND2_X1  g595(.A1(new_n706), .A2(new_n707), .ZN(new_n782));
  NAND3_X1  g596(.A1(new_n475), .A2(new_n777), .A3(new_n647), .ZN(new_n783));
  XNOR2_X1  g597(.A(new_n783), .B(KEYINPUT112), .ZN(new_n784));
  OAI21_X1  g598(.A(new_n782), .B1(new_n643), .B2(new_n784), .ZN(new_n785));
  AOI21_X1  g599(.A(new_n721), .B1(new_n785), .B2(new_n711), .ZN(new_n786));
  AND4_X1   g600(.A1(new_n718), .A2(new_n776), .A3(new_n781), .A4(new_n786), .ZN(new_n787));
  AOI21_X1  g601(.A(KEYINPUT52), .B1(new_n766), .B2(new_n768), .ZN(new_n788));
  NAND2_X1  g602(.A1(new_n788), .A2(KEYINPUT114), .ZN(new_n789));
  NAND4_X1  g603(.A1(new_n774), .A2(new_n787), .A3(KEYINPUT53), .A4(new_n789), .ZN(new_n790));
  INV_X1    g604(.A(KEYINPUT53), .ZN(new_n791));
  AND3_X1   g605(.A1(new_n766), .A2(new_n768), .A3(KEYINPUT52), .ZN(new_n792));
  NOR2_X1   g606(.A1(new_n792), .A2(new_n788), .ZN(new_n793));
  NOR2_X1   g607(.A1(new_n775), .A2(new_n780), .ZN(new_n794));
  NAND3_X1  g608(.A1(new_n794), .A2(new_n718), .A3(new_n786), .ZN(new_n795));
  OAI21_X1  g609(.A(new_n791), .B1(new_n793), .B2(new_n795), .ZN(new_n796));
  NAND2_X1  g610(.A1(new_n790), .A2(new_n796), .ZN(new_n797));
  NOR2_X1   g611(.A1(new_n797), .A2(KEYINPUT54), .ZN(new_n798));
  AOI211_X1 g612(.A(new_n772), .B(KEYINPUT52), .C1(new_n766), .C2(new_n768), .ZN(new_n799));
  AOI21_X1  g613(.A(new_n799), .B1(new_n793), .B2(new_n772), .ZN(new_n800));
  AOI21_X1  g614(.A(KEYINPUT53), .B1(new_n800), .B2(new_n787), .ZN(new_n801));
  AND2_X1   g615(.A1(new_n786), .A2(new_n718), .ZN(new_n802));
  OAI211_X1 g616(.A(new_n802), .B(new_n794), .C1(new_n788), .C2(new_n792), .ZN(new_n803));
  NOR2_X1   g617(.A1(new_n803), .A2(new_n791), .ZN(new_n804));
  OR2_X1    g618(.A1(new_n801), .A2(new_n804), .ZN(new_n805));
  AOI21_X1  g619(.A(new_n798), .B1(new_n805), .B2(KEYINPUT54), .ZN(new_n806));
  INV_X1    g620(.A(KEYINPUT51), .ZN(new_n807));
  NAND3_X1  g621(.A1(new_n703), .A2(new_n477), .A3(new_n726), .ZN(new_n808));
  NAND3_X1  g622(.A1(new_n670), .A2(new_n681), .A3(new_n363), .ZN(new_n809));
  NOR2_X1   g623(.A1(new_n808), .A2(new_n809), .ZN(new_n810));
  XNOR2_X1  g624(.A(new_n810), .B(KEYINPUT50), .ZN(new_n811));
  NAND2_X1  g625(.A1(new_n681), .A2(new_n710), .ZN(new_n812));
  NAND2_X1  g626(.A1(new_n596), .A2(new_n477), .ZN(new_n813));
  NOR3_X1   g627(.A1(new_n812), .A2(new_n657), .A3(new_n813), .ZN(new_n814));
  NOR2_X1   g628(.A1(new_n474), .A2(new_n609), .ZN(new_n815));
  NAND2_X1  g629(.A1(new_n814), .A2(new_n815), .ZN(new_n816));
  AND2_X1   g630(.A1(new_n811), .A2(new_n816), .ZN(new_n817));
  INV_X1    g631(.A(new_n808), .ZN(new_n818));
  NOR2_X1   g632(.A1(new_n680), .A2(new_n361), .ZN(new_n819));
  OAI211_X1 g633(.A(new_n710), .B(new_n818), .C1(new_n749), .C2(new_n819), .ZN(new_n820));
  NAND2_X1  g634(.A1(new_n817), .A2(new_n820), .ZN(new_n821));
  NAND2_X1  g635(.A1(new_n726), .A2(new_n477), .ZN(new_n822));
  OR3_X1    g636(.A1(new_n822), .A2(new_n812), .A3(KEYINPUT115), .ZN(new_n823));
  OAI21_X1  g637(.A(KEYINPUT115), .B1(new_n822), .B2(new_n812), .ZN(new_n824));
  NAND2_X1  g638(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  NAND2_X1  g639(.A1(new_n825), .A2(new_n706), .ZN(new_n826));
  XNOR2_X1  g640(.A(new_n826), .B(KEYINPUT116), .ZN(new_n827));
  OAI21_X1  g641(.A(new_n807), .B1(new_n821), .B2(new_n827), .ZN(new_n828));
  INV_X1    g642(.A(KEYINPUT116), .ZN(new_n829));
  XNOR2_X1  g643(.A(new_n826), .B(new_n829), .ZN(new_n830));
  NAND4_X1  g644(.A1(new_n830), .A2(new_n817), .A3(KEYINPUT51), .A4(new_n820), .ZN(new_n831));
  NAND2_X1  g645(.A1(new_n556), .A2(new_n596), .ZN(new_n832));
  INV_X1    g646(.A(new_n832), .ZN(new_n833));
  INV_X1    g647(.A(KEYINPUT48), .ZN(new_n834));
  AOI22_X1  g648(.A1(new_n825), .A2(new_n833), .B1(KEYINPUT117), .B2(new_n834), .ZN(new_n835));
  OAI21_X1  g649(.A(new_n835), .B1(KEYINPUT117), .B2(new_n834), .ZN(new_n836));
  INV_X1    g650(.A(KEYINPUT117), .ZN(new_n837));
  NAND4_X1  g651(.A1(new_n825), .A2(new_n837), .A3(KEYINPUT48), .A4(new_n833), .ZN(new_n838));
  NAND2_X1  g652(.A1(new_n818), .A2(new_n694), .ZN(new_n839));
  NAND2_X1  g653(.A1(new_n339), .A2(G952), .ZN(new_n840));
  AOI21_X1  g654(.A(new_n840), .B1(new_n814), .B2(new_n610), .ZN(new_n841));
  AND4_X1   g655(.A1(new_n836), .A2(new_n838), .A3(new_n839), .A4(new_n841), .ZN(new_n842));
  NAND3_X1  g656(.A1(new_n828), .A2(new_n831), .A3(new_n842), .ZN(new_n843));
  NAND2_X1  g657(.A1(new_n843), .A2(KEYINPUT118), .ZN(new_n844));
  OR2_X1    g658(.A1(new_n843), .A2(KEYINPUT118), .ZN(new_n845));
  AND3_X1   g659(.A1(new_n806), .A2(new_n844), .A3(new_n845), .ZN(new_n846));
  NOR2_X1   g660(.A1(G952), .A2(G953), .ZN(new_n847));
  OAI21_X1  g661(.A(new_n759), .B1(new_n846), .B2(new_n847), .ZN(G75));
  NOR2_X1   g662(.A1(new_n339), .A2(G952), .ZN(new_n849));
  INV_X1    g663(.A(new_n849), .ZN(new_n850));
  NOR2_X1   g664(.A1(new_n795), .A2(new_n791), .ZN(new_n851));
  AOI22_X1  g665(.A1(new_n800), .A2(new_n851), .B1(new_n791), .B2(new_n803), .ZN(new_n852));
  NOR2_X1   g666(.A1(new_n852), .A2(new_n232), .ZN(new_n853));
  AOI21_X1  g667(.A(KEYINPUT56), .B1(new_n853), .B2(G210), .ZN(new_n854));
  NAND2_X1  g668(.A1(new_n386), .A2(new_n395), .ZN(new_n855));
  XNOR2_X1  g669(.A(new_n855), .B(new_n393), .ZN(new_n856));
  XNOR2_X1  g670(.A(new_n856), .B(KEYINPUT55), .ZN(new_n857));
  OAI21_X1  g671(.A(new_n850), .B1(new_n854), .B2(new_n857), .ZN(new_n858));
  INV_X1    g672(.A(KEYINPUT119), .ZN(new_n859));
  AOI21_X1  g673(.A(new_n859), .B1(new_n797), .B2(G902), .ZN(new_n860));
  AOI211_X1 g674(.A(KEYINPUT119), .B(new_n232), .C1(new_n790), .C2(new_n796), .ZN(new_n861));
  NOR2_X1   g675(.A1(new_n860), .A2(new_n861), .ZN(new_n862));
  NAND2_X1  g676(.A1(new_n862), .A2(new_n365), .ZN(new_n863));
  INV_X1    g677(.A(KEYINPUT56), .ZN(new_n864));
  AND2_X1   g678(.A1(new_n857), .A2(new_n864), .ZN(new_n865));
  AOI21_X1  g679(.A(new_n858), .B1(new_n863), .B2(new_n865), .ZN(G51));
  INV_X1    g680(.A(KEYINPUT120), .ZN(new_n867));
  INV_X1    g681(.A(KEYINPUT54), .ZN(new_n868));
  NAND3_X1  g682(.A1(new_n852), .A2(new_n867), .A3(new_n868), .ZN(new_n869));
  OAI21_X1  g683(.A(KEYINPUT120), .B1(new_n797), .B2(KEYINPUT54), .ZN(new_n870));
  OAI211_X1 g684(.A(new_n869), .B(new_n870), .C1(new_n868), .C2(new_n852), .ZN(new_n871));
  XOR2_X1   g685(.A(new_n737), .B(KEYINPUT57), .Z(new_n872));
  NAND2_X1  g686(.A1(new_n871), .A2(new_n872), .ZN(new_n873));
  XOR2_X1   g687(.A(new_n353), .B(KEYINPUT121), .Z(new_n874));
  NAND2_X1  g688(.A1(new_n873), .A2(new_n874), .ZN(new_n875));
  INV_X1    g689(.A(new_n736), .ZN(new_n876));
  NAND2_X1  g690(.A1(new_n862), .A2(new_n876), .ZN(new_n877));
  AOI21_X1  g691(.A(new_n849), .B1(new_n875), .B2(new_n877), .ZN(G54));
  INV_X1    g692(.A(KEYINPUT122), .ZN(new_n879));
  AND2_X1   g693(.A1(KEYINPUT58), .A2(G475), .ZN(new_n880));
  AOI21_X1  g694(.A(new_n465), .B1(new_n862), .B2(new_n880), .ZN(new_n881));
  OAI21_X1  g695(.A(KEYINPUT119), .B1(new_n852), .B2(new_n232), .ZN(new_n882));
  NAND3_X1  g696(.A1(new_n797), .A2(new_n859), .A3(G902), .ZN(new_n883));
  AND2_X1   g697(.A1(new_n465), .A2(new_n880), .ZN(new_n884));
  NAND3_X1  g698(.A1(new_n882), .A2(new_n883), .A3(new_n884), .ZN(new_n885));
  NAND2_X1  g699(.A1(new_n885), .A2(new_n850), .ZN(new_n886));
  OAI21_X1  g700(.A(new_n879), .B1(new_n881), .B2(new_n886), .ZN(new_n887));
  NAND3_X1  g701(.A1(new_n882), .A2(new_n883), .A3(new_n880), .ZN(new_n888));
  INV_X1    g702(.A(new_n465), .ZN(new_n889));
  NAND2_X1  g703(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  NAND4_X1  g704(.A1(new_n890), .A2(KEYINPUT122), .A3(new_n850), .A4(new_n885), .ZN(new_n891));
  NAND2_X1  g705(.A1(new_n887), .A2(new_n891), .ZN(G60));
  NAND2_X1  g706(.A1(G478), .A2(G902), .ZN(new_n893));
  XOR2_X1   g707(.A(new_n893), .B(KEYINPUT59), .Z(new_n894));
  OAI21_X1  g708(.A(new_n606), .B1(new_n806), .B2(new_n894), .ZN(new_n895));
  NOR2_X1   g709(.A1(new_n606), .A2(new_n894), .ZN(new_n896));
  NAND2_X1  g710(.A1(new_n871), .A2(new_n896), .ZN(new_n897));
  AND3_X1   g711(.A1(new_n895), .A2(new_n850), .A3(new_n897), .ZN(G63));
  NAND2_X1  g712(.A1(G217), .A2(G902), .ZN(new_n899));
  XNOR2_X1  g713(.A(new_n899), .B(KEYINPUT124), .ZN(new_n900));
  XOR2_X1   g714(.A(KEYINPUT123), .B(KEYINPUT60), .Z(new_n901));
  XNOR2_X1  g715(.A(new_n900), .B(new_n901), .ZN(new_n902));
  NOR2_X1   g716(.A1(new_n852), .A2(new_n902), .ZN(new_n903));
  XNOR2_X1  g717(.A(new_n632), .B(KEYINPUT125), .ZN(new_n904));
  NAND2_X1  g718(.A1(new_n903), .A2(new_n904), .ZN(new_n905));
  OAI211_X1 g719(.A(new_n905), .B(new_n850), .C1(new_n593), .C2(new_n903), .ZN(new_n906));
  INV_X1    g720(.A(KEYINPUT61), .ZN(new_n907));
  XNOR2_X1  g721(.A(new_n906), .B(new_n907), .ZN(G66));
  OAI21_X1  g722(.A(G953), .B1(new_n391), .B2(new_n479), .ZN(new_n909));
  OAI21_X1  g723(.A(new_n909), .B1(new_n794), .B2(G953), .ZN(new_n910));
  OAI21_X1  g724(.A(new_n855), .B1(G898), .B2(new_n339), .ZN(new_n911));
  XOR2_X1   g725(.A(new_n911), .B(KEYINPUT126), .Z(new_n912));
  XNOR2_X1  g726(.A(new_n910), .B(new_n912), .ZN(G69));
  OAI21_X1  g727(.A(new_n493), .B1(new_n524), .B2(new_n525), .ZN(new_n914));
  XOR2_X1   g728(.A(new_n914), .B(KEYINPUT127), .Z(new_n915));
  XNOR2_X1  g729(.A(new_n915), .B(new_n453), .ZN(new_n916));
  INV_X1    g730(.A(new_n916), .ZN(new_n917));
  NAND2_X1  g731(.A1(new_n778), .A2(new_n710), .ZN(new_n918));
  OR3_X1    g732(.A1(new_n832), .A2(new_n666), .A3(new_n918), .ZN(new_n919));
  OAI211_X1 g733(.A(new_n752), .B(new_n919), .C1(new_n742), .C2(new_n743), .ZN(new_n920));
  NAND2_X1  g734(.A1(new_n672), .A2(new_n768), .ZN(new_n921));
  XNOR2_X1  g735(.A(new_n921), .B(KEYINPUT62), .ZN(new_n922));
  OAI211_X1 g736(.A(new_n339), .B(new_n917), .C1(new_n920), .C2(new_n922), .ZN(new_n923));
  NOR2_X1   g737(.A1(new_n645), .A2(new_n339), .ZN(new_n924));
  OAI21_X1  g738(.A(new_n752), .B1(new_n742), .B2(new_n743), .ZN(new_n925));
  INV_X1    g739(.A(new_n721), .ZN(new_n926));
  NAND4_X1  g740(.A1(new_n833), .A2(new_n741), .A3(new_n665), .A4(new_n700), .ZN(new_n927));
  AND4_X1   g741(.A1(new_n718), .A2(new_n926), .A3(new_n768), .A4(new_n927), .ZN(new_n928));
  INV_X1    g742(.A(new_n928), .ZN(new_n929));
  NOR2_X1   g743(.A1(new_n925), .A2(new_n929), .ZN(new_n930));
  AOI21_X1  g744(.A(new_n924), .B1(new_n930), .B2(new_n339), .ZN(new_n931));
  OAI21_X1  g745(.A(new_n923), .B1(new_n931), .B2(new_n917), .ZN(new_n932));
  AOI21_X1  g746(.A(new_n339), .B1(G227), .B2(G900), .ZN(new_n933));
  XOR2_X1   g747(.A(new_n932), .B(new_n933), .Z(G72));
  INV_X1    g748(.A(new_n794), .ZN(new_n935));
  NOR3_X1   g749(.A1(new_n920), .A2(new_n922), .A3(new_n935), .ZN(new_n936));
  NAND2_X1  g750(.A1(G472), .A2(G902), .ZN(new_n937));
  XNOR2_X1  g751(.A(new_n937), .B(KEYINPUT63), .ZN(new_n938));
  OAI21_X1  g752(.A(new_n653), .B1(new_n936), .B2(new_n938), .ZN(new_n939));
  INV_X1    g753(.A(new_n552), .ZN(new_n940));
  NOR3_X1   g754(.A1(new_n925), .A2(new_n935), .A3(new_n929), .ZN(new_n941));
  OAI21_X1  g755(.A(new_n940), .B1(new_n941), .B2(new_n938), .ZN(new_n942));
  NAND3_X1  g756(.A1(new_n939), .A2(new_n942), .A3(new_n850), .ZN(new_n943));
  NOR3_X1   g757(.A1(new_n940), .A2(new_n653), .A3(new_n938), .ZN(new_n944));
  AOI21_X1  g758(.A(new_n943), .B1(new_n805), .B2(new_n944), .ZN(G57));
endmodule


