//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 0 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 0 0 0 0 0 1 1 1 1 0 1 1 1 0 0 0 0 0 0 1 0 0 1 0 0 1 1 0 1 0 1 0 1 1 1 0 0 1 0 1 1 0 0 1 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:42:07 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n202, new_n203, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1032, new_n1033, new_n1034,
    new_n1035, new_n1036, new_n1037, new_n1038, new_n1039, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1055, new_n1056, new_n1057, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1107, new_n1108,
    new_n1109, new_n1110, new_n1111, new_n1112, new_n1113, new_n1114,
    new_n1115, new_n1116, new_n1117, new_n1118, new_n1119, new_n1120,
    new_n1121, new_n1122, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1173, new_n1174, new_n1175,
    new_n1176, new_n1177, new_n1178, new_n1179, new_n1180, new_n1181,
    new_n1182, new_n1183, new_n1184, new_n1185, new_n1186, new_n1187,
    new_n1188, new_n1189, new_n1190, new_n1191, new_n1192, new_n1193,
    new_n1194, new_n1195, new_n1196, new_n1197, new_n1198, new_n1199,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1214, new_n1215, new_n1216, new_n1217, new_n1218, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1279, new_n1280;
  NOR4_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .A4(G77), .ZN(G353));
  NOR2_X1   g0001(.A1(G97), .A2(G107), .ZN(new_n202));
  INV_X1    g0002(.A(new_n202), .ZN(new_n203));
  NAND2_X1  g0003(.A1(new_n203), .A2(G87), .ZN(G355));
  NAND2_X1  g0004(.A1(G1), .A2(G20), .ZN(new_n205));
  AOI22_X1  g0005(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n206));
  INV_X1    g0006(.A(G68), .ZN(new_n207));
  INV_X1    g0007(.A(G238), .ZN(new_n208));
  INV_X1    g0008(.A(G107), .ZN(new_n209));
  INV_X1    g0009(.A(G264), .ZN(new_n210));
  OAI221_X1 g0010(.A(new_n206), .B1(new_n207), .B2(new_n208), .C1(new_n209), .C2(new_n210), .ZN(new_n211));
  AOI21_X1  g0011(.A(new_n211), .B1(G116), .B2(G270), .ZN(new_n212));
  INV_X1    g0012(.A(G50), .ZN(new_n213));
  INV_X1    g0013(.A(G226), .ZN(new_n214));
  INV_X1    g0014(.A(G77), .ZN(new_n215));
  INV_X1    g0015(.A(G244), .ZN(new_n216));
  OAI221_X1 g0016(.A(new_n212), .B1(new_n213), .B2(new_n214), .C1(new_n215), .C2(new_n216), .ZN(new_n217));
  INV_X1    g0017(.A(G58), .ZN(new_n218));
  INV_X1    g0018(.A(G232), .ZN(new_n219));
  NOR2_X1   g0019(.A1(new_n218), .A2(new_n219), .ZN(new_n220));
  OAI21_X1  g0020(.A(new_n205), .B1(new_n217), .B2(new_n220), .ZN(new_n221));
  NAND2_X1  g0021(.A1(new_n221), .A2(KEYINPUT1), .ZN(new_n222));
  XNOR2_X1  g0022(.A(new_n222), .B(KEYINPUT65), .ZN(new_n223));
  NOR2_X1   g0023(.A1(new_n205), .A2(G13), .ZN(new_n224));
  OAI211_X1 g0024(.A(new_n224), .B(G250), .C1(G257), .C2(G264), .ZN(new_n225));
  XNOR2_X1  g0025(.A(new_n225), .B(KEYINPUT0), .ZN(new_n226));
  OAI211_X1 g0026(.A(new_n223), .B(new_n226), .C1(KEYINPUT1), .C2(new_n221), .ZN(new_n227));
  NAND2_X1  g0027(.A1(G1), .A2(G13), .ZN(new_n228));
  INV_X1    g0028(.A(G20), .ZN(new_n229));
  NOR2_X1   g0029(.A1(new_n228), .A2(new_n229), .ZN(new_n230));
  OAI21_X1  g0030(.A(G50), .B1(G58), .B2(G68), .ZN(new_n231));
  XOR2_X1   g0031(.A(new_n231), .B(KEYINPUT64), .Z(new_n232));
  AOI21_X1  g0032(.A(new_n227), .B1(new_n230), .B2(new_n232), .ZN(G361));
  XNOR2_X1  g0033(.A(KEYINPUT2), .B(G226), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n234), .B(new_n219), .ZN(new_n235));
  XNOR2_X1  g0035(.A(G238), .B(G244), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XNOR2_X1  g0037(.A(G250), .B(G257), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n238), .B(new_n210), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n239), .B(G270), .ZN(new_n240));
  XOR2_X1   g0040(.A(new_n237), .B(new_n240), .Z(G358));
  XOR2_X1   g0041(.A(G68), .B(G77), .Z(new_n242));
  XNOR2_X1  g0042(.A(G50), .B(G58), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XOR2_X1   g0044(.A(G107), .B(G116), .Z(new_n245));
  XNOR2_X1  g0045(.A(G87), .B(G97), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n245), .B(new_n246), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n244), .B(new_n247), .ZN(G351));
  NAND3_X1  g0048(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n249));
  NAND2_X1  g0049(.A1(new_n249), .A2(new_n228), .ZN(new_n250));
  XNOR2_X1  g0050(.A(KEYINPUT8), .B(G58), .ZN(new_n251));
  NAND2_X1  g0051(.A1(new_n229), .A2(G33), .ZN(new_n252));
  NOR2_X1   g0052(.A1(new_n251), .A2(new_n252), .ZN(new_n253));
  NOR3_X1   g0053(.A1(G50), .A2(G58), .A3(G68), .ZN(new_n254));
  INV_X1    g0054(.A(G33), .ZN(new_n255));
  NAND2_X1  g0055(.A1(new_n229), .A2(new_n255), .ZN(new_n256));
  INV_X1    g0056(.A(G150), .ZN(new_n257));
  OAI22_X1  g0057(.A1(new_n254), .A2(new_n229), .B1(new_n256), .B2(new_n257), .ZN(new_n258));
  OAI21_X1  g0058(.A(new_n250), .B1(new_n253), .B2(new_n258), .ZN(new_n259));
  XOR2_X1   g0059(.A(new_n259), .B(KEYINPUT66), .Z(new_n260));
  INV_X1    g0060(.A(G1), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n261), .A2(G20), .ZN(new_n262));
  NAND2_X1  g0062(.A1(new_n262), .A2(G50), .ZN(new_n263));
  XOR2_X1   g0063(.A(new_n263), .B(KEYINPUT67), .Z(new_n264));
  INV_X1    g0064(.A(G13), .ZN(new_n265));
  NOR3_X1   g0065(.A1(new_n265), .A2(new_n229), .A3(G1), .ZN(new_n266));
  NOR2_X1   g0066(.A1(new_n266), .A2(new_n250), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n264), .A2(new_n267), .ZN(new_n268));
  INV_X1    g0068(.A(new_n266), .ZN(new_n269));
  OAI211_X1 g0069(.A(new_n260), .B(new_n268), .C1(G50), .C2(new_n269), .ZN(new_n270));
  INV_X1    g0070(.A(KEYINPUT9), .ZN(new_n271));
  NOR2_X1   g0071(.A1(new_n270), .A2(new_n271), .ZN(new_n272));
  INV_X1    g0072(.A(KEYINPUT68), .ZN(new_n273));
  XNOR2_X1  g0073(.A(new_n272), .B(new_n273), .ZN(new_n274));
  INV_X1    g0074(.A(KEYINPUT3), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n275), .A2(new_n255), .ZN(new_n276));
  NAND2_X1  g0076(.A1(KEYINPUT3), .A2(G33), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n276), .A2(new_n277), .ZN(new_n278));
  INV_X1    g0078(.A(G1698), .ZN(new_n279));
  NAND2_X1  g0079(.A1(new_n279), .A2(G222), .ZN(new_n280));
  NAND2_X1  g0080(.A1(G223), .A2(G1698), .ZN(new_n281));
  NAND3_X1  g0081(.A1(new_n278), .A2(new_n280), .A3(new_n281), .ZN(new_n282));
  INV_X1    g0082(.A(G41), .ZN(new_n283));
  OAI211_X1 g0083(.A(G1), .B(G13), .C1(new_n255), .C2(new_n283), .ZN(new_n284));
  INV_X1    g0084(.A(new_n284), .ZN(new_n285));
  OAI211_X1 g0085(.A(new_n282), .B(new_n285), .C1(G77), .C2(new_n278), .ZN(new_n286));
  OAI21_X1  g0086(.A(new_n261), .B1(G41), .B2(G45), .ZN(new_n287));
  INV_X1    g0087(.A(G274), .ZN(new_n288));
  NOR2_X1   g0088(.A1(new_n287), .A2(new_n288), .ZN(new_n289));
  INV_X1    g0089(.A(new_n289), .ZN(new_n290));
  NAND2_X1  g0090(.A1(new_n284), .A2(new_n287), .ZN(new_n291));
  OAI211_X1 g0091(.A(new_n286), .B(new_n290), .C1(new_n214), .C2(new_n291), .ZN(new_n292));
  INV_X1    g0092(.A(G190), .ZN(new_n293));
  NOR2_X1   g0093(.A1(new_n292), .A2(new_n293), .ZN(new_n294));
  AOI21_X1  g0094(.A(new_n294), .B1(new_n270), .B2(new_n271), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n292), .A2(G200), .ZN(new_n296));
  OR2_X1    g0096(.A1(new_n296), .A2(KEYINPUT69), .ZN(new_n297));
  AND2_X1   g0097(.A1(new_n295), .A2(new_n297), .ZN(new_n298));
  INV_X1    g0098(.A(KEYINPUT10), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n296), .A2(KEYINPUT69), .ZN(new_n300));
  NAND4_X1  g0100(.A1(new_n274), .A2(new_n298), .A3(new_n299), .A4(new_n300), .ZN(new_n301));
  AND2_X1   g0101(.A1(new_n295), .A2(new_n296), .ZN(new_n302));
  AND2_X1   g0102(.A1(new_n274), .A2(new_n302), .ZN(new_n303));
  OAI21_X1  g0103(.A(new_n301), .B1(new_n303), .B2(new_n299), .ZN(new_n304));
  INV_X1    g0104(.A(G169), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n292), .A2(new_n305), .ZN(new_n306));
  OR2_X1    g0106(.A1(new_n292), .A2(G179), .ZN(new_n307));
  NAND3_X1  g0107(.A1(new_n270), .A2(new_n306), .A3(new_n307), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n304), .A2(new_n308), .ZN(new_n309));
  INV_X1    g0109(.A(new_n309), .ZN(new_n310));
  INV_X1    g0110(.A(new_n250), .ZN(new_n311));
  INV_X1    g0111(.A(KEYINPUT75), .ZN(new_n312));
  INV_X1    g0112(.A(G159), .ZN(new_n313));
  OAI21_X1  g0113(.A(new_n312), .B1(new_n256), .B2(new_n313), .ZN(new_n314));
  NOR2_X1   g0114(.A1(G20), .A2(G33), .ZN(new_n315));
  NAND3_X1  g0115(.A1(new_n315), .A2(KEYINPUT75), .A3(G159), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n314), .A2(new_n316), .ZN(new_n317));
  XNOR2_X1  g0117(.A(G58), .B(G68), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n318), .A2(G20), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n317), .A2(new_n319), .ZN(new_n320));
  NAND2_X1  g0120(.A1(new_n275), .A2(KEYINPUT74), .ZN(new_n321));
  INV_X1    g0121(.A(KEYINPUT74), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n322), .A2(KEYINPUT3), .ZN(new_n323));
  NAND3_X1  g0123(.A1(new_n321), .A2(new_n323), .A3(G33), .ZN(new_n324));
  INV_X1    g0124(.A(KEYINPUT7), .ZN(new_n325));
  NAND4_X1  g0125(.A1(new_n324), .A2(new_n325), .A3(new_n229), .A4(new_n276), .ZN(new_n326));
  AND2_X1   g0126(.A1(new_n326), .A2(G68), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n324), .A2(new_n276), .ZN(new_n328));
  OAI21_X1  g0128(.A(KEYINPUT7), .B1(new_n328), .B2(G20), .ZN(new_n329));
  AOI21_X1  g0129(.A(new_n320), .B1(new_n327), .B2(new_n329), .ZN(new_n330));
  AOI21_X1  g0130(.A(new_n311), .B1(new_n330), .B2(KEYINPUT16), .ZN(new_n331));
  AOI21_X1  g0131(.A(G20), .B1(KEYINPUT3), .B2(G33), .ZN(new_n332));
  XNOR2_X1  g0132(.A(KEYINPUT74), .B(KEYINPUT3), .ZN(new_n333));
  OAI211_X1 g0133(.A(KEYINPUT7), .B(new_n332), .C1(new_n333), .C2(G33), .ZN(new_n334));
  NAND3_X1  g0134(.A1(new_n276), .A2(new_n229), .A3(new_n277), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n335), .A2(new_n325), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n334), .A2(new_n336), .ZN(new_n337));
  AOI21_X1  g0137(.A(KEYINPUT76), .B1(new_n337), .B2(G68), .ZN(new_n338));
  INV_X1    g0138(.A(KEYINPUT76), .ZN(new_n339));
  AOI211_X1 g0139(.A(new_n339), .B(new_n207), .C1(new_n334), .C2(new_n336), .ZN(new_n340));
  NOR3_X1   g0140(.A1(new_n338), .A2(new_n340), .A3(new_n320), .ZN(new_n341));
  OAI21_X1  g0141(.A(new_n331), .B1(new_n341), .B2(KEYINPUT16), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n251), .A2(new_n266), .ZN(new_n343));
  NAND2_X1  g0143(.A1(new_n311), .A2(new_n262), .ZN(new_n344));
  OAI21_X1  g0144(.A(new_n343), .B1(new_n344), .B2(new_n251), .ZN(new_n345));
  XNOR2_X1  g0145(.A(new_n345), .B(KEYINPUT77), .ZN(new_n346));
  INV_X1    g0146(.A(new_n346), .ZN(new_n347));
  OAI21_X1  g0147(.A(new_n290), .B1(new_n291), .B2(new_n219), .ZN(new_n348));
  INV_X1    g0148(.A(new_n348), .ZN(new_n349));
  AOI22_X1  g0149(.A1(new_n324), .A2(new_n276), .B1(new_n214), .B2(G1698), .ZN(new_n350));
  OR2_X1    g0150(.A1(G223), .A2(G1698), .ZN(new_n351));
  AOI22_X1  g0151(.A1(new_n350), .A2(new_n351), .B1(G33), .B2(G87), .ZN(new_n352));
  OAI21_X1  g0152(.A(new_n349), .B1(new_n352), .B2(new_n284), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n353), .A2(G200), .ZN(new_n354));
  OR2_X1    g0154(.A1(new_n353), .A2(new_n293), .ZN(new_n355));
  NAND4_X1  g0155(.A1(new_n342), .A2(new_n347), .A3(new_n354), .A4(new_n355), .ZN(new_n356));
  INV_X1    g0156(.A(KEYINPUT17), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n356), .A2(new_n357), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n321), .A2(new_n323), .ZN(new_n359));
  AOI21_X1  g0159(.A(new_n325), .B1(new_n359), .B2(new_n255), .ZN(new_n360));
  AOI22_X1  g0160(.A1(new_n360), .A2(new_n332), .B1(new_n325), .B2(new_n335), .ZN(new_n361));
  OAI21_X1  g0161(.A(new_n339), .B1(new_n361), .B2(new_n207), .ZN(new_n362));
  AND2_X1   g0162(.A1(new_n317), .A2(new_n319), .ZN(new_n363));
  NAND3_X1  g0163(.A1(new_n337), .A2(KEYINPUT76), .A3(G68), .ZN(new_n364));
  NAND3_X1  g0164(.A1(new_n362), .A2(new_n363), .A3(new_n364), .ZN(new_n365));
  INV_X1    g0165(.A(KEYINPUT16), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n365), .A2(new_n366), .ZN(new_n367));
  AOI21_X1  g0167(.A(new_n346), .B1(new_n367), .B2(new_n331), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n353), .A2(G169), .ZN(new_n369));
  OAI211_X1 g0169(.A(G179), .B(new_n349), .C1(new_n352), .C2(new_n284), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n369), .A2(new_n370), .ZN(new_n371));
  INV_X1    g0171(.A(new_n371), .ZN(new_n372));
  OAI21_X1  g0172(.A(KEYINPUT18), .B1(new_n368), .B2(new_n372), .ZN(new_n373));
  NAND4_X1  g0173(.A1(new_n368), .A2(KEYINPUT17), .A3(new_n354), .A4(new_n355), .ZN(new_n374));
  INV_X1    g0174(.A(KEYINPUT18), .ZN(new_n375));
  INV_X1    g0175(.A(new_n276), .ZN(new_n376));
  AOI21_X1  g0176(.A(new_n376), .B1(new_n333), .B2(G33), .ZN(new_n377));
  AOI21_X1  g0177(.A(new_n325), .B1(new_n377), .B2(new_n229), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n326), .A2(G68), .ZN(new_n379));
  OAI211_X1 g0179(.A(KEYINPUT16), .B(new_n363), .C1(new_n378), .C2(new_n379), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n380), .A2(new_n250), .ZN(new_n381));
  AOI21_X1  g0181(.A(new_n381), .B1(new_n366), .B2(new_n365), .ZN(new_n382));
  OAI211_X1 g0182(.A(new_n375), .B(new_n371), .C1(new_n382), .C2(new_n346), .ZN(new_n383));
  NAND4_X1  g0183(.A1(new_n358), .A2(new_n373), .A3(new_n374), .A4(new_n383), .ZN(new_n384));
  NOR2_X1   g0184(.A1(new_n265), .A2(G1), .ZN(new_n385));
  NAND3_X1  g0185(.A1(new_n385), .A2(G20), .A3(new_n207), .ZN(new_n386));
  INV_X1    g0186(.A(KEYINPUT12), .ZN(new_n387));
  NOR2_X1   g0187(.A1(new_n386), .A2(new_n387), .ZN(new_n388));
  INV_X1    g0188(.A(new_n388), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n386), .A2(new_n387), .ZN(new_n390));
  INV_X1    g0190(.A(KEYINPUT72), .ZN(new_n391));
  INV_X1    g0191(.A(new_n344), .ZN(new_n392));
  AOI21_X1  g0192(.A(new_n391), .B1(new_n392), .B2(G68), .ZN(new_n393));
  NOR3_X1   g0193(.A1(new_n344), .A2(KEYINPUT72), .A3(new_n207), .ZN(new_n394));
  OAI211_X1 g0194(.A(new_n389), .B(new_n390), .C1(new_n393), .C2(new_n394), .ZN(new_n395));
  NOR2_X1   g0195(.A1(new_n255), .A2(G20), .ZN(new_n396));
  AOI22_X1  g0196(.A1(new_n396), .A2(G77), .B1(G20), .B2(new_n207), .ZN(new_n397));
  XNOR2_X1  g0197(.A(new_n397), .B(KEYINPUT71), .ZN(new_n398));
  OAI21_X1  g0198(.A(new_n398), .B1(new_n213), .B2(new_n256), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n399), .A2(new_n250), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n400), .A2(KEYINPUT11), .ZN(new_n401));
  INV_X1    g0201(.A(KEYINPUT11), .ZN(new_n402));
  NAND3_X1  g0202(.A1(new_n399), .A2(new_n402), .A3(new_n250), .ZN(new_n403));
  AOI21_X1  g0203(.A(new_n395), .B1(new_n401), .B2(new_n403), .ZN(new_n404));
  NAND2_X1  g0204(.A1(G33), .A2(G97), .ZN(new_n405));
  OAI21_X1  g0205(.A(new_n278), .B1(G232), .B2(new_n279), .ZN(new_n406));
  NOR2_X1   g0206(.A1(G226), .A2(G1698), .ZN(new_n407));
  OAI21_X1  g0207(.A(new_n405), .B1(new_n406), .B2(new_n407), .ZN(new_n408));
  AOI21_X1  g0208(.A(new_n289), .B1(new_n408), .B2(new_n285), .ZN(new_n409));
  INV_X1    g0209(.A(KEYINPUT13), .ZN(new_n410));
  INV_X1    g0210(.A(KEYINPUT70), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n291), .A2(new_n411), .ZN(new_n412));
  NAND3_X1  g0212(.A1(new_n284), .A2(KEYINPUT70), .A3(new_n287), .ZN(new_n413));
  NAND3_X1  g0213(.A1(new_n412), .A2(G238), .A3(new_n413), .ZN(new_n414));
  NAND3_X1  g0214(.A1(new_n409), .A2(new_n410), .A3(new_n414), .ZN(new_n415));
  INV_X1    g0215(.A(new_n415), .ZN(new_n416));
  AOI21_X1  g0216(.A(new_n410), .B1(new_n409), .B2(new_n414), .ZN(new_n417));
  OAI21_X1  g0217(.A(G200), .B1(new_n416), .B2(new_n417), .ZN(new_n418));
  INV_X1    g0218(.A(new_n417), .ZN(new_n419));
  NAND3_X1  g0219(.A1(new_n419), .A2(G190), .A3(new_n415), .ZN(new_n420));
  AND3_X1   g0220(.A1(new_n404), .A2(new_n418), .A3(new_n420), .ZN(new_n421));
  NOR2_X1   g0221(.A1(new_n416), .A2(new_n417), .ZN(new_n422));
  OAI21_X1  g0222(.A(KEYINPUT14), .B1(new_n422), .B2(new_n305), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n422), .A2(G179), .ZN(new_n424));
  INV_X1    g0224(.A(KEYINPUT14), .ZN(new_n425));
  OAI211_X1 g0225(.A(new_n425), .B(G169), .C1(new_n416), .C2(new_n417), .ZN(new_n426));
  NAND3_X1  g0226(.A1(new_n423), .A2(new_n424), .A3(new_n426), .ZN(new_n427));
  INV_X1    g0227(.A(new_n404), .ZN(new_n428));
  AOI21_X1  g0228(.A(new_n421), .B1(new_n427), .B2(new_n428), .ZN(new_n429));
  AOI21_X1  g0229(.A(new_n384), .B1(new_n429), .B2(KEYINPUT73), .ZN(new_n430));
  INV_X1    g0230(.A(new_n251), .ZN(new_n431));
  AOI22_X1  g0231(.A1(new_n431), .A2(new_n315), .B1(G20), .B2(G77), .ZN(new_n432));
  XOR2_X1   g0232(.A(KEYINPUT15), .B(G87), .Z(new_n433));
  INV_X1    g0233(.A(new_n433), .ZN(new_n434));
  OAI21_X1  g0234(.A(new_n432), .B1(new_n252), .B2(new_n434), .ZN(new_n435));
  AOI22_X1  g0235(.A1(new_n435), .A2(new_n250), .B1(G77), .B2(new_n392), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n266), .A2(new_n215), .ZN(new_n437));
  NAND2_X1  g0237(.A1(new_n436), .A2(new_n437), .ZN(new_n438));
  NAND2_X1  g0238(.A1(G238), .A2(G1698), .ZN(new_n439));
  OAI211_X1 g0239(.A(new_n278), .B(new_n439), .C1(new_n219), .C2(G1698), .ZN(new_n440));
  OAI211_X1 g0240(.A(new_n440), .B(new_n285), .C1(G107), .C2(new_n278), .ZN(new_n441));
  OAI211_X1 g0241(.A(new_n441), .B(new_n290), .C1(new_n216), .C2(new_n291), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n442), .A2(new_n305), .ZN(new_n443));
  OAI211_X1 g0243(.A(new_n438), .B(new_n443), .C1(G179), .C2(new_n442), .ZN(new_n444));
  OR2_X1    g0244(.A1(new_n442), .A2(new_n293), .ZN(new_n445));
  NAND2_X1  g0245(.A1(new_n442), .A2(G200), .ZN(new_n446));
  NAND4_X1  g0246(.A1(new_n445), .A2(new_n437), .A3(new_n436), .A4(new_n446), .ZN(new_n447));
  OAI211_X1 g0247(.A(new_n444), .B(new_n447), .C1(new_n429), .C2(KEYINPUT73), .ZN(new_n448));
  INV_X1    g0248(.A(new_n448), .ZN(new_n449));
  AND3_X1   g0249(.A1(new_n310), .A2(new_n430), .A3(new_n449), .ZN(new_n450));
  INV_X1    g0250(.A(new_n450), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n261), .A2(G33), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n267), .A2(new_n452), .ZN(new_n453));
  INV_X1    g0253(.A(new_n453), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n454), .A2(G116), .ZN(new_n455));
  NOR2_X1   g0255(.A1(new_n269), .A2(G116), .ZN(new_n456));
  INV_X1    g0256(.A(new_n456), .ZN(new_n457));
  NAND2_X1  g0257(.A1(G33), .A2(G283), .ZN(new_n458));
  INV_X1    g0258(.A(KEYINPUT78), .ZN(new_n459));
  XNOR2_X1  g0259(.A(new_n458), .B(new_n459), .ZN(new_n460));
  AOI21_X1  g0260(.A(G20), .B1(new_n255), .B2(G97), .ZN(new_n461));
  NAND2_X1  g0261(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  INV_X1    g0262(.A(G116), .ZN(new_n463));
  AOI22_X1  g0263(.A1(new_n249), .A2(new_n228), .B1(G20), .B2(new_n463), .ZN(new_n464));
  NAND3_X1  g0264(.A1(new_n462), .A2(KEYINPUT20), .A3(new_n464), .ZN(new_n465));
  INV_X1    g0265(.A(new_n465), .ZN(new_n466));
  AOI21_X1  g0266(.A(KEYINPUT20), .B1(new_n462), .B2(new_n464), .ZN(new_n467));
  OAI211_X1 g0267(.A(new_n455), .B(new_n457), .C1(new_n466), .C2(new_n467), .ZN(new_n468));
  INV_X1    g0268(.A(G45), .ZN(new_n469));
  NOR2_X1   g0269(.A1(new_n469), .A2(G1), .ZN(new_n470));
  AND2_X1   g0270(.A1(KEYINPUT5), .A2(G41), .ZN(new_n471));
  NOR2_X1   g0271(.A1(KEYINPUT5), .A2(G41), .ZN(new_n472));
  OAI21_X1  g0272(.A(new_n470), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n473), .A2(new_n284), .ZN(new_n474));
  INV_X1    g0274(.A(new_n474), .ZN(new_n475));
  INV_X1    g0275(.A(new_n473), .ZN(new_n476));
  AOI22_X1  g0276(.A1(new_n475), .A2(G270), .B1(G274), .B2(new_n476), .ZN(new_n477));
  INV_X1    g0277(.A(G303), .ZN(new_n478));
  NOR2_X1   g0278(.A1(new_n278), .A2(new_n478), .ZN(new_n479));
  AOI22_X1  g0279(.A1(new_n324), .A2(new_n276), .B1(new_n210), .B2(G1698), .ZN(new_n480));
  OR2_X1    g0280(.A1(G257), .A2(G1698), .ZN(new_n481));
  AOI21_X1  g0281(.A(new_n479), .B1(new_n480), .B2(new_n481), .ZN(new_n482));
  OAI21_X1  g0282(.A(new_n477), .B1(new_n284), .B2(new_n482), .ZN(new_n483));
  NAND3_X1  g0283(.A1(new_n468), .A2(new_n483), .A3(G169), .ZN(new_n484));
  INV_X1    g0284(.A(KEYINPUT21), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n484), .A2(new_n485), .ZN(new_n486));
  AND2_X1   g0286(.A1(new_n480), .A2(new_n481), .ZN(new_n487));
  OAI21_X1  g0287(.A(new_n285), .B1(new_n487), .B2(new_n479), .ZN(new_n488));
  AOI21_X1  g0288(.A(new_n305), .B1(new_n488), .B2(new_n477), .ZN(new_n489));
  NAND3_X1  g0289(.A1(new_n489), .A2(KEYINPUT21), .A3(new_n468), .ZN(new_n490));
  INV_X1    g0290(.A(G179), .ZN(new_n491));
  NOR2_X1   g0291(.A1(new_n483), .A2(new_n491), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n492), .A2(new_n468), .ZN(new_n493));
  AND3_X1   g0293(.A1(new_n486), .A2(new_n490), .A3(new_n493), .ZN(new_n494));
  INV_X1    g0294(.A(KEYINPUT84), .ZN(new_n495));
  INV_X1    g0295(.A(new_n468), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n483), .A2(G200), .ZN(new_n497));
  OAI211_X1 g0297(.A(new_n496), .B(new_n497), .C1(new_n293), .C2(new_n483), .ZN(new_n498));
  NAND3_X1  g0298(.A1(new_n494), .A2(new_n495), .A3(new_n498), .ZN(new_n499));
  NAND4_X1  g0299(.A1(new_n498), .A2(new_n486), .A3(new_n490), .A4(new_n493), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n500), .A2(KEYINPUT84), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n499), .A2(new_n501), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n454), .A2(new_n433), .ZN(new_n503));
  NAND3_X1  g0303(.A1(new_n328), .A2(new_n229), .A3(G68), .ZN(new_n504));
  INV_X1    g0304(.A(KEYINPUT19), .ZN(new_n505));
  NAND3_X1  g0305(.A1(new_n396), .A2(new_n505), .A3(G97), .ZN(new_n506));
  AOI21_X1  g0306(.A(G20), .B1(G33), .B2(G97), .ZN(new_n507));
  INV_X1    g0307(.A(G87), .ZN(new_n508));
  AOI21_X1  g0308(.A(new_n507), .B1(new_n508), .B2(new_n202), .ZN(new_n509));
  OAI21_X1  g0309(.A(new_n506), .B1(new_n509), .B2(new_n505), .ZN(new_n510));
  AOI21_X1  g0310(.A(new_n311), .B1(new_n504), .B2(new_n510), .ZN(new_n511));
  NOR2_X1   g0311(.A1(new_n269), .A2(new_n433), .ZN(new_n512));
  NOR3_X1   g0312(.A1(new_n511), .A2(KEYINPUT81), .A3(new_n512), .ZN(new_n513));
  INV_X1    g0313(.A(KEYINPUT81), .ZN(new_n514));
  AOI211_X1 g0314(.A(G20), .B(new_n207), .C1(new_n324), .C2(new_n276), .ZN(new_n515));
  INV_X1    g0315(.A(G97), .ZN(new_n516));
  NOR3_X1   g0316(.A1(new_n252), .A2(KEYINPUT19), .A3(new_n516), .ZN(new_n517));
  INV_X1    g0317(.A(new_n507), .ZN(new_n518));
  OAI21_X1  g0318(.A(new_n518), .B1(new_n203), .B2(G87), .ZN(new_n519));
  AOI21_X1  g0319(.A(new_n517), .B1(new_n519), .B2(KEYINPUT19), .ZN(new_n520));
  OAI21_X1  g0320(.A(new_n250), .B1(new_n515), .B2(new_n520), .ZN(new_n521));
  INV_X1    g0321(.A(new_n512), .ZN(new_n522));
  AOI21_X1  g0322(.A(new_n514), .B1(new_n521), .B2(new_n522), .ZN(new_n523));
  OAI21_X1  g0323(.A(new_n503), .B1(new_n513), .B2(new_n523), .ZN(new_n524));
  INV_X1    g0324(.A(new_n470), .ZN(new_n525));
  OAI21_X1  g0325(.A(new_n284), .B1(new_n525), .B2(G274), .ZN(new_n526));
  INV_X1    g0326(.A(G250), .ZN(new_n527));
  AOI21_X1  g0327(.A(new_n526), .B1(new_n527), .B2(new_n525), .ZN(new_n528));
  AOI21_X1  g0328(.A(new_n216), .B1(new_n324), .B2(new_n276), .ZN(new_n529));
  AOI22_X1  g0329(.A1(new_n529), .A2(G1698), .B1(G33), .B2(G116), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n279), .A2(G238), .ZN(new_n531));
  OAI21_X1  g0331(.A(KEYINPUT80), .B1(new_n377), .B2(new_n531), .ZN(new_n532));
  INV_X1    g0332(.A(KEYINPUT80), .ZN(new_n533));
  INV_X1    g0333(.A(new_n531), .ZN(new_n534));
  NAND3_X1  g0334(.A1(new_n328), .A2(new_n533), .A3(new_n534), .ZN(new_n535));
  NAND3_X1  g0335(.A1(new_n530), .A2(new_n532), .A3(new_n535), .ZN(new_n536));
  AOI21_X1  g0336(.A(new_n528), .B1(new_n536), .B2(new_n285), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n537), .A2(new_n491), .ZN(new_n538));
  AOI21_X1  g0338(.A(new_n533), .B1(new_n328), .B2(new_n534), .ZN(new_n539));
  AOI211_X1 g0339(.A(KEYINPUT80), .B(new_n531), .C1(new_n324), .C2(new_n276), .ZN(new_n540));
  NOR2_X1   g0340(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  AOI21_X1  g0341(.A(new_n284), .B1(new_n541), .B2(new_n530), .ZN(new_n542));
  OAI21_X1  g0342(.A(new_n305), .B1(new_n542), .B2(new_n528), .ZN(new_n543));
  NAND3_X1  g0343(.A1(new_n524), .A2(new_n538), .A3(new_n543), .ZN(new_n544));
  OAI21_X1  g0344(.A(KEYINPUT81), .B1(new_n511), .B2(new_n512), .ZN(new_n545));
  NAND3_X1  g0345(.A1(new_n521), .A2(new_n514), .A3(new_n522), .ZN(new_n546));
  NOR2_X1   g0346(.A1(new_n453), .A2(new_n508), .ZN(new_n547));
  OR2_X1    g0347(.A1(new_n547), .A2(KEYINPUT82), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n547), .A2(KEYINPUT82), .ZN(new_n549));
  AOI22_X1  g0349(.A1(new_n545), .A2(new_n546), .B1(new_n548), .B2(new_n549), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n537), .A2(G190), .ZN(new_n551));
  OAI21_X1  g0351(.A(G200), .B1(new_n542), .B2(new_n528), .ZN(new_n552));
  NAND3_X1  g0352(.A1(new_n550), .A2(new_n551), .A3(new_n552), .ZN(new_n553));
  AND3_X1   g0353(.A1(new_n544), .A2(new_n553), .A3(KEYINPUT83), .ZN(new_n554));
  AOI21_X1  g0354(.A(KEYINPUT83), .B1(new_n544), .B2(new_n553), .ZN(new_n555));
  NOR2_X1   g0355(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n502), .A2(new_n556), .ZN(new_n557));
  NOR2_X1   g0357(.A1(new_n453), .A2(new_n516), .ZN(new_n558));
  NOR2_X1   g0358(.A1(new_n256), .A2(new_n215), .ZN(new_n559));
  INV_X1    g0359(.A(new_n559), .ZN(new_n560));
  INV_X1    g0360(.A(KEYINPUT6), .ZN(new_n561));
  NOR2_X1   g0361(.A1(new_n516), .A2(new_n209), .ZN(new_n562));
  OAI21_X1  g0362(.A(new_n561), .B1(new_n562), .B2(new_n202), .ZN(new_n563));
  NAND3_X1  g0363(.A1(new_n209), .A2(KEYINPUT6), .A3(G97), .ZN(new_n564));
  AND2_X1   g0364(.A1(new_n563), .A2(new_n564), .ZN(new_n565));
  OAI221_X1 g0365(.A(new_n560), .B1(new_n565), .B2(new_n229), .C1(new_n361), .C2(new_n209), .ZN(new_n566));
  AOI21_X1  g0366(.A(new_n558), .B1(new_n566), .B2(new_n250), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n266), .A2(new_n516), .ZN(new_n568));
  NAND3_X1  g0368(.A1(new_n567), .A2(KEYINPUT79), .A3(new_n568), .ZN(new_n569));
  NOR2_X1   g0369(.A1(KEYINPUT4), .A2(G1698), .ZN(new_n570));
  NAND3_X1  g0370(.A1(new_n278), .A2(G244), .A3(new_n279), .ZN(new_n571));
  AOI22_X1  g0371(.A1(new_n529), .A2(new_n570), .B1(new_n571), .B2(KEYINPUT4), .ZN(new_n572));
  NAND3_X1  g0372(.A1(new_n278), .A2(G250), .A3(G1698), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n573), .A2(new_n460), .ZN(new_n574));
  OAI21_X1  g0374(.A(new_n285), .B1(new_n572), .B2(new_n574), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n476), .A2(G274), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n475), .A2(G257), .ZN(new_n577));
  NAND3_X1  g0377(.A1(new_n575), .A2(new_n576), .A3(new_n577), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n578), .A2(G169), .ZN(new_n579));
  NAND4_X1  g0379(.A1(new_n575), .A2(G179), .A3(new_n576), .A4(new_n577), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  INV_X1    g0381(.A(new_n558), .ZN(new_n582));
  AOI21_X1  g0382(.A(new_n229), .B1(new_n563), .B2(new_n564), .ZN(new_n583));
  AOI211_X1 g0383(.A(new_n559), .B(new_n583), .C1(G107), .C2(new_n337), .ZN(new_n584));
  OAI211_X1 g0384(.A(new_n568), .B(new_n582), .C1(new_n584), .C2(new_n311), .ZN(new_n585));
  INV_X1    g0385(.A(KEYINPUT79), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  NAND3_X1  g0387(.A1(new_n569), .A2(new_n581), .A3(new_n587), .ZN(new_n588));
  INV_X1    g0388(.A(new_n585), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n578), .A2(G200), .ZN(new_n590));
  OAI211_X1 g0390(.A(new_n589), .B(new_n590), .C1(new_n293), .C2(new_n578), .ZN(new_n591));
  AND2_X1   g0391(.A1(new_n588), .A2(new_n591), .ZN(new_n592));
  NAND3_X1  g0392(.A1(new_n229), .A2(G33), .A3(G116), .ZN(new_n593));
  NOR2_X1   g0393(.A1(new_n229), .A2(G107), .ZN(new_n594));
  OR2_X1    g0394(.A1(KEYINPUT86), .A2(KEYINPUT23), .ZN(new_n595));
  NAND2_X1  g0395(.A1(KEYINPUT86), .A2(KEYINPUT23), .ZN(new_n596));
  NAND3_X1  g0396(.A1(new_n594), .A2(new_n595), .A3(new_n596), .ZN(new_n597));
  OAI21_X1  g0397(.A(new_n597), .B1(new_n594), .B2(new_n595), .ZN(new_n598));
  NAND2_X1  g0398(.A1(KEYINPUT22), .A2(G87), .ZN(new_n599));
  AOI211_X1 g0399(.A(G20), .B(new_n599), .C1(new_n324), .C2(new_n276), .ZN(new_n600));
  AOI21_X1  g0400(.A(G20), .B1(new_n276), .B2(new_n277), .ZN(new_n601));
  AOI21_X1  g0401(.A(KEYINPUT22), .B1(new_n601), .B2(G87), .ZN(new_n602));
  NOR3_X1   g0402(.A1(new_n600), .A2(KEYINPUT85), .A3(new_n602), .ZN(new_n603));
  INV_X1    g0403(.A(KEYINPUT85), .ZN(new_n604));
  NAND4_X1  g0404(.A1(new_n328), .A2(KEYINPUT22), .A3(new_n229), .A4(G87), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n601), .A2(G87), .ZN(new_n606));
  INV_X1    g0406(.A(KEYINPUT22), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  AOI21_X1  g0408(.A(new_n604), .B1(new_n605), .B2(new_n608), .ZN(new_n609));
  OAI211_X1 g0409(.A(new_n593), .B(new_n598), .C1(new_n603), .C2(new_n609), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n610), .A2(KEYINPUT24), .ZN(new_n611));
  OAI21_X1  g0411(.A(KEYINPUT85), .B1(new_n600), .B2(new_n602), .ZN(new_n612));
  NAND3_X1  g0412(.A1(new_n605), .A2(new_n604), .A3(new_n608), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n612), .A2(new_n613), .ZN(new_n614));
  INV_X1    g0414(.A(KEYINPUT24), .ZN(new_n615));
  NAND4_X1  g0415(.A1(new_n614), .A2(new_n615), .A3(new_n593), .A4(new_n598), .ZN(new_n616));
  AOI21_X1  g0416(.A(new_n311), .B1(new_n611), .B2(new_n616), .ZN(new_n617));
  INV_X1    g0417(.A(new_n617), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n266), .A2(new_n209), .ZN(new_n619));
  XOR2_X1   g0419(.A(KEYINPUT87), .B(KEYINPUT25), .Z(new_n620));
  XNOR2_X1  g0420(.A(new_n619), .B(new_n620), .ZN(new_n621));
  OAI21_X1  g0421(.A(new_n621), .B1(new_n209), .B2(new_n453), .ZN(new_n622));
  INV_X1    g0422(.A(new_n622), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n527), .A2(new_n279), .ZN(new_n624));
  OAI211_X1 g0424(.A(new_n328), .B(new_n624), .C1(G257), .C2(new_n279), .ZN(new_n625));
  NAND2_X1  g0425(.A1(G33), .A2(G294), .ZN(new_n626));
  AOI21_X1  g0426(.A(new_n284), .B1(new_n625), .B2(new_n626), .ZN(new_n627));
  OAI21_X1  g0427(.A(new_n576), .B1(new_n210), .B2(new_n474), .ZN(new_n628));
  NOR2_X1   g0428(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n629), .A2(new_n293), .ZN(new_n630));
  OAI21_X1  g0430(.A(new_n630), .B1(G200), .B2(new_n629), .ZN(new_n631));
  NAND3_X1  g0431(.A1(new_n618), .A2(new_n623), .A3(new_n631), .ZN(new_n632));
  NOR2_X1   g0432(.A1(new_n629), .A2(G169), .ZN(new_n633));
  AOI21_X1  g0433(.A(new_n633), .B1(new_n491), .B2(new_n629), .ZN(new_n634));
  OAI21_X1  g0434(.A(new_n634), .B1(new_n617), .B2(new_n622), .ZN(new_n635));
  NAND3_X1  g0435(.A1(new_n592), .A2(new_n632), .A3(new_n635), .ZN(new_n636));
  NOR3_X1   g0436(.A1(new_n451), .A2(new_n557), .A3(new_n636), .ZN(G372));
  INV_X1    g0437(.A(new_n308), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n427), .A2(new_n428), .ZN(new_n639));
  OAI21_X1  g0439(.A(new_n639), .B1(new_n421), .B2(new_n444), .ZN(new_n640));
  XNOR2_X1  g0440(.A(new_n640), .B(KEYINPUT90), .ZN(new_n641));
  AND2_X1   g0441(.A1(new_n358), .A2(new_n374), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  AND3_X1   g0443(.A1(new_n373), .A2(KEYINPUT89), .A3(new_n383), .ZN(new_n644));
  AOI21_X1  g0444(.A(KEYINPUT89), .B1(new_n373), .B2(new_n383), .ZN(new_n645));
  NOR2_X1   g0445(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  INV_X1    g0446(.A(new_n646), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n643), .A2(new_n647), .ZN(new_n648));
  AOI21_X1  g0448(.A(new_n638), .B1(new_n648), .B2(new_n304), .ZN(new_n649));
  INV_X1    g0449(.A(KEYINPUT88), .ZN(new_n650));
  INV_X1    g0450(.A(G200), .ZN(new_n651));
  OAI21_X1  g0451(.A(new_n650), .B1(new_n537), .B2(new_n651), .ZN(new_n652));
  OAI211_X1 g0452(.A(KEYINPUT88), .B(G200), .C1(new_n542), .C2(new_n528), .ZN(new_n653));
  NAND4_X1  g0453(.A1(new_n652), .A2(new_n653), .A3(new_n550), .A4(new_n551), .ZN(new_n654));
  AOI22_X1  g0454(.A1(new_n579), .A2(new_n580), .B1(new_n567), .B2(new_n568), .ZN(new_n655));
  INV_X1    g0455(.A(KEYINPUT26), .ZN(new_n656));
  NAND4_X1  g0456(.A1(new_n654), .A2(new_n655), .A3(new_n544), .A4(new_n656), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n657), .A2(new_n544), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n544), .A2(new_n553), .ZN(new_n659));
  INV_X1    g0459(.A(KEYINPUT83), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  NAND3_X1  g0461(.A1(new_n544), .A2(new_n553), .A3(KEYINPUT83), .ZN(new_n662));
  INV_X1    g0462(.A(new_n588), .ZN(new_n663));
  NAND3_X1  g0463(.A1(new_n661), .A2(new_n662), .A3(new_n663), .ZN(new_n664));
  AOI21_X1  g0464(.A(new_n658), .B1(new_n664), .B2(KEYINPUT26), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n635), .A2(new_n494), .ZN(new_n666));
  AND2_X1   g0466(.A1(new_n654), .A2(new_n544), .ZN(new_n667));
  NAND4_X1  g0467(.A1(new_n666), .A2(new_n592), .A3(new_n632), .A4(new_n667), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n665), .A2(new_n668), .ZN(new_n669));
  INV_X1    g0469(.A(new_n669), .ZN(new_n670));
  OAI21_X1  g0470(.A(new_n649), .B1(new_n451), .B2(new_n670), .ZN(G369));
  NAND2_X1  g0471(.A1(new_n618), .A2(new_n623), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n385), .A2(new_n229), .ZN(new_n673));
  OR2_X1    g0473(.A1(new_n673), .A2(KEYINPUT27), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n673), .A2(KEYINPUT27), .ZN(new_n675));
  NAND3_X1  g0475(.A1(new_n674), .A2(G213), .A3(new_n675), .ZN(new_n676));
  INV_X1    g0476(.A(G343), .ZN(new_n677));
  NOR2_X1   g0477(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  INV_X1    g0478(.A(new_n678), .ZN(new_n679));
  NAND3_X1  g0479(.A1(new_n672), .A2(new_n634), .A3(new_n679), .ZN(new_n680));
  INV_X1    g0480(.A(new_n680), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n672), .A2(new_n678), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n682), .A2(new_n632), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n683), .A2(new_n635), .ZN(new_n684));
  NOR2_X1   g0484(.A1(new_n494), .A2(new_n678), .ZN(new_n685));
  AOI21_X1  g0485(.A(new_n681), .B1(new_n684), .B2(new_n685), .ZN(new_n686));
  XNOR2_X1  g0486(.A(new_n502), .B(KEYINPUT91), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n468), .A2(new_n678), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  NAND3_X1  g0489(.A1(new_n494), .A2(new_n468), .A3(new_n678), .ZN(new_n690));
  NAND3_X1  g0490(.A1(new_n689), .A2(G330), .A3(new_n690), .ZN(new_n691));
  AOI21_X1  g0491(.A(new_n681), .B1(new_n635), .B2(new_n683), .ZN(new_n692));
  INV_X1    g0492(.A(new_n692), .ZN(new_n693));
  OAI21_X1  g0493(.A(new_n686), .B1(new_n691), .B2(new_n693), .ZN(G399));
  INV_X1    g0494(.A(new_n224), .ZN(new_n695));
  NOR2_X1   g0495(.A1(new_n695), .A2(G41), .ZN(new_n696));
  INV_X1    g0496(.A(new_n696), .ZN(new_n697));
  NOR3_X1   g0497(.A1(new_n203), .A2(G87), .A3(G116), .ZN(new_n698));
  NAND3_X1  g0498(.A1(new_n697), .A2(G1), .A3(new_n698), .ZN(new_n699));
  OAI21_X1  g0499(.A(new_n699), .B1(new_n231), .B2(new_n697), .ZN(new_n700));
  XNOR2_X1  g0500(.A(new_n700), .B(KEYINPUT28), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n669), .A2(new_n679), .ZN(new_n702));
  NOR2_X1   g0502(.A1(new_n702), .A2(KEYINPUT29), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n667), .A2(new_n655), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n704), .A2(KEYINPUT26), .ZN(new_n705));
  XNOR2_X1  g0505(.A(new_n544), .B(KEYINPUT93), .ZN(new_n706));
  NAND3_X1  g0506(.A1(new_n668), .A2(new_n705), .A3(new_n706), .ZN(new_n707));
  NOR2_X1   g0507(.A1(new_n664), .A2(KEYINPUT26), .ZN(new_n708));
  OAI21_X1  g0508(.A(new_n679), .B1(new_n707), .B2(new_n708), .ZN(new_n709));
  AND2_X1   g0509(.A1(new_n709), .A2(KEYINPUT29), .ZN(new_n710));
  NOR3_X1   g0510(.A1(new_n557), .A2(new_n636), .A3(new_n678), .ZN(new_n711));
  NAND2_X1  g0511(.A1(new_n492), .A2(new_n537), .ZN(new_n712));
  NAND3_X1  g0512(.A1(new_n629), .A2(new_n577), .A3(new_n575), .ZN(new_n713));
  INV_X1    g0513(.A(KEYINPUT30), .ZN(new_n714));
  OR3_X1    g0514(.A1(new_n712), .A2(new_n713), .A3(new_n714), .ZN(new_n715));
  OAI21_X1  g0515(.A(new_n714), .B1(new_n712), .B2(new_n713), .ZN(new_n716));
  INV_X1    g0516(.A(new_n629), .ZN(new_n717));
  NAND4_X1  g0517(.A1(new_n717), .A2(new_n578), .A3(new_n491), .A4(new_n483), .ZN(new_n718));
  OAI211_X1 g0518(.A(new_n715), .B(new_n716), .C1(new_n537), .C2(new_n718), .ZN(new_n719));
  NAND2_X1  g0519(.A1(new_n719), .A2(new_n678), .ZN(new_n720));
  INV_X1    g0520(.A(KEYINPUT31), .ZN(new_n721));
  NAND2_X1  g0521(.A1(new_n720), .A2(new_n721), .ZN(new_n722));
  NAND3_X1  g0522(.A1(new_n719), .A2(KEYINPUT31), .A3(new_n678), .ZN(new_n723));
  NAND2_X1  g0523(.A1(new_n722), .A2(new_n723), .ZN(new_n724));
  OAI21_X1  g0524(.A(G330), .B1(new_n711), .B2(new_n724), .ZN(new_n725));
  NAND2_X1  g0525(.A1(new_n725), .A2(KEYINPUT92), .ZN(new_n726));
  INV_X1    g0526(.A(KEYINPUT92), .ZN(new_n727));
  OAI211_X1 g0527(.A(new_n727), .B(G330), .C1(new_n711), .C2(new_n724), .ZN(new_n728));
  AOI211_X1 g0528(.A(new_n703), .B(new_n710), .C1(new_n726), .C2(new_n728), .ZN(new_n729));
  OAI21_X1  g0529(.A(new_n701), .B1(new_n729), .B2(G1), .ZN(G364));
  NAND2_X1  g0530(.A1(new_n689), .A2(new_n690), .ZN(new_n731));
  XNOR2_X1  g0531(.A(new_n731), .B(G330), .ZN(new_n732));
  NOR2_X1   g0532(.A1(new_n265), .A2(G20), .ZN(new_n733));
  NAND2_X1  g0533(.A1(new_n733), .A2(G45), .ZN(new_n734));
  NAND3_X1  g0534(.A1(new_n697), .A2(G1), .A3(new_n734), .ZN(new_n735));
  NAND2_X1  g0535(.A1(new_n232), .A2(new_n469), .ZN(new_n736));
  NOR2_X1   g0536(.A1(new_n328), .A2(new_n695), .ZN(new_n737));
  OAI211_X1 g0537(.A(new_n736), .B(new_n737), .C1(new_n244), .C2(new_n469), .ZN(new_n738));
  INV_X1    g0538(.A(G355), .ZN(new_n739));
  NAND2_X1  g0539(.A1(new_n278), .A2(new_n224), .ZN(new_n740));
  OAI221_X1 g0540(.A(new_n738), .B1(G116), .B2(new_n224), .C1(new_n739), .C2(new_n740), .ZN(new_n741));
  NOR2_X1   g0541(.A1(G13), .A2(G33), .ZN(new_n742));
  INV_X1    g0542(.A(new_n742), .ZN(new_n743));
  NOR2_X1   g0543(.A1(new_n743), .A2(G20), .ZN(new_n744));
  AOI21_X1  g0544(.A(new_n228), .B1(G20), .B2(new_n305), .ZN(new_n745));
  NOR2_X1   g0545(.A1(new_n744), .A2(new_n745), .ZN(new_n746));
  AOI21_X1  g0546(.A(new_n735), .B1(new_n741), .B2(new_n746), .ZN(new_n747));
  XNOR2_X1  g0547(.A(new_n747), .B(KEYINPUT94), .ZN(new_n748));
  NOR2_X1   g0548(.A1(new_n229), .A2(G179), .ZN(new_n749));
  NOR2_X1   g0549(.A1(G190), .A2(G200), .ZN(new_n750));
  AND2_X1   g0550(.A1(new_n749), .A2(new_n750), .ZN(new_n751));
  OR2_X1    g0551(.A1(new_n751), .A2(KEYINPUT96), .ZN(new_n752));
  NAND2_X1  g0552(.A1(new_n751), .A2(KEYINPUT96), .ZN(new_n753));
  NAND2_X1  g0553(.A1(new_n752), .A2(new_n753), .ZN(new_n754));
  NOR2_X1   g0554(.A1(new_n754), .A2(new_n313), .ZN(new_n755));
  XNOR2_X1  g0555(.A(new_n755), .B(KEYINPUT32), .ZN(new_n756));
  INV_X1    g0556(.A(new_n278), .ZN(new_n757));
  NOR2_X1   g0557(.A1(new_n229), .A2(new_n491), .ZN(new_n758));
  INV_X1    g0558(.A(new_n758), .ZN(new_n759));
  NOR3_X1   g0559(.A1(new_n759), .A2(new_n293), .A3(G200), .ZN(new_n760));
  INV_X1    g0560(.A(new_n760), .ZN(new_n761));
  NAND3_X1  g0561(.A1(new_n749), .A2(new_n293), .A3(G200), .ZN(new_n762));
  OAI22_X1  g0562(.A1(new_n761), .A2(new_n218), .B1(new_n209), .B2(new_n762), .ZN(new_n763));
  NAND2_X1  g0563(.A1(new_n758), .A2(G200), .ZN(new_n764));
  NOR2_X1   g0564(.A1(new_n764), .A2(G190), .ZN(new_n765));
  AOI211_X1 g0565(.A(new_n757), .B(new_n763), .C1(G68), .C2(new_n765), .ZN(new_n766));
  NOR3_X1   g0566(.A1(new_n293), .A2(G179), .A3(G200), .ZN(new_n767));
  NOR2_X1   g0567(.A1(new_n767), .A2(new_n229), .ZN(new_n768));
  NOR2_X1   g0568(.A1(new_n768), .A2(new_n516), .ZN(new_n769));
  INV_X1    g0569(.A(new_n769), .ZN(new_n770));
  NAND2_X1  g0570(.A1(new_n758), .A2(new_n750), .ZN(new_n771));
  XNOR2_X1  g0571(.A(new_n771), .B(KEYINPUT95), .ZN(new_n772));
  INV_X1    g0572(.A(new_n772), .ZN(new_n773));
  OAI21_X1  g0573(.A(new_n770), .B1(new_n773), .B2(new_n215), .ZN(new_n774));
  NOR2_X1   g0574(.A1(new_n764), .A2(new_n293), .ZN(new_n775));
  AOI21_X1  g0575(.A(new_n774), .B1(G50), .B2(new_n775), .ZN(new_n776));
  NAND3_X1  g0576(.A1(new_n749), .A2(G190), .A3(G200), .ZN(new_n777));
  INV_X1    g0577(.A(new_n777), .ZN(new_n778));
  NAND2_X1  g0578(.A1(new_n778), .A2(G87), .ZN(new_n779));
  NAND4_X1  g0579(.A1(new_n756), .A2(new_n766), .A3(new_n776), .A4(new_n779), .ZN(new_n780));
  OAI21_X1  g0580(.A(new_n757), .B1(new_n777), .B2(new_n478), .ZN(new_n781));
  INV_X1    g0581(.A(new_n771), .ZN(new_n782));
  NAND2_X1  g0582(.A1(new_n782), .A2(G311), .ZN(new_n783));
  INV_X1    g0583(.A(G294), .ZN(new_n784));
  INV_X1    g0584(.A(new_n775), .ZN(new_n785));
  INV_X1    g0585(.A(G326), .ZN(new_n786));
  OAI221_X1 g0586(.A(new_n783), .B1(new_n784), .B2(new_n768), .C1(new_n785), .C2(new_n786), .ZN(new_n787));
  XOR2_X1   g0587(.A(new_n787), .B(KEYINPUT97), .Z(new_n788));
  INV_X1    g0588(.A(new_n754), .ZN(new_n789));
  AOI211_X1 g0589(.A(new_n781), .B(new_n788), .C1(G329), .C2(new_n789), .ZN(new_n790));
  INV_X1    g0590(.A(G283), .ZN(new_n791));
  INV_X1    g0591(.A(G322), .ZN(new_n792));
  OAI221_X1 g0592(.A(new_n790), .B1(new_n791), .B2(new_n762), .C1(new_n792), .C2(new_n761), .ZN(new_n793));
  INV_X1    g0593(.A(new_n765), .ZN(new_n794));
  XOR2_X1   g0594(.A(KEYINPUT33), .B(G317), .Z(new_n795));
  NOR2_X1   g0595(.A1(new_n794), .A2(new_n795), .ZN(new_n796));
  OAI21_X1  g0596(.A(new_n780), .B1(new_n793), .B2(new_n796), .ZN(new_n797));
  AOI22_X1  g0597(.A1(new_n731), .A2(new_n744), .B1(new_n745), .B2(new_n797), .ZN(new_n798));
  AOI22_X1  g0598(.A1(new_n732), .A2(new_n735), .B1(new_n748), .B2(new_n798), .ZN(new_n799));
  INV_X1    g0599(.A(new_n799), .ZN(G396));
  NAND2_X1  g0600(.A1(new_n726), .A2(new_n728), .ZN(new_n801));
  NAND2_X1  g0601(.A1(new_n438), .A2(new_n678), .ZN(new_n802));
  NAND2_X1  g0602(.A1(new_n447), .A2(new_n802), .ZN(new_n803));
  NAND2_X1  g0603(.A1(new_n803), .A2(new_n444), .ZN(new_n804));
  NOR2_X1   g0604(.A1(new_n444), .A2(new_n678), .ZN(new_n805));
  INV_X1    g0605(.A(new_n805), .ZN(new_n806));
  NAND2_X1  g0606(.A1(new_n804), .A2(new_n806), .ZN(new_n807));
  INV_X1    g0607(.A(new_n807), .ZN(new_n808));
  XNOR2_X1  g0608(.A(new_n702), .B(new_n808), .ZN(new_n809));
  XNOR2_X1  g0609(.A(new_n801), .B(new_n809), .ZN(new_n810));
  NAND2_X1  g0610(.A1(new_n810), .A2(new_n735), .ZN(new_n811));
  AOI22_X1  g0611(.A1(new_n775), .A2(G303), .B1(new_n778), .B2(G107), .ZN(new_n812));
  OAI221_X1 g0612(.A(new_n812), .B1(new_n791), .B2(new_n794), .C1(new_n773), .C2(new_n463), .ZN(new_n813));
  INV_X1    g0613(.A(new_n762), .ZN(new_n814));
  AOI21_X1  g0614(.A(new_n813), .B1(G87), .B2(new_n814), .ZN(new_n815));
  NAND2_X1  g0615(.A1(new_n789), .A2(G311), .ZN(new_n816));
  NAND3_X1  g0616(.A1(new_n815), .A2(new_n770), .A3(new_n816), .ZN(new_n817));
  AOI211_X1 g0617(.A(new_n278), .B(new_n817), .C1(G294), .C2(new_n760), .ZN(new_n818));
  AOI22_X1  g0618(.A1(new_n772), .A2(G159), .B1(G150), .B2(new_n765), .ZN(new_n819));
  NAND2_X1  g0619(.A1(new_n775), .A2(G137), .ZN(new_n820));
  INV_X1    g0620(.A(G143), .ZN(new_n821));
  OAI211_X1 g0621(.A(new_n819), .B(new_n820), .C1(new_n821), .C2(new_n761), .ZN(new_n822));
  XOR2_X1   g0622(.A(new_n822), .B(KEYINPUT34), .Z(new_n823));
  OAI22_X1  g0623(.A1(new_n762), .A2(new_n207), .B1(new_n777), .B2(new_n213), .ZN(new_n824));
  XOR2_X1   g0624(.A(new_n824), .B(KEYINPUT98), .Z(new_n825));
  INV_X1    g0625(.A(G132), .ZN(new_n826));
  OAI221_X1 g0626(.A(new_n328), .B1(new_n218), .B2(new_n768), .C1(new_n754), .C2(new_n826), .ZN(new_n827));
  NOR3_X1   g0627(.A1(new_n823), .A2(new_n825), .A3(new_n827), .ZN(new_n828));
  OAI21_X1  g0628(.A(new_n745), .B1(new_n818), .B2(new_n828), .ZN(new_n829));
  INV_X1    g0629(.A(new_n735), .ZN(new_n830));
  NAND2_X1  g0630(.A1(new_n807), .A2(new_n742), .ZN(new_n831));
  NOR2_X1   g0631(.A1(new_n745), .A2(new_n742), .ZN(new_n832));
  NAND2_X1  g0632(.A1(new_n832), .A2(new_n215), .ZN(new_n833));
  NAND4_X1  g0633(.A1(new_n829), .A2(new_n830), .A3(new_n831), .A4(new_n833), .ZN(new_n834));
  NAND2_X1  g0634(.A1(new_n811), .A2(new_n834), .ZN(G384));
  INV_X1    g0635(.A(new_n724), .ZN(new_n836));
  INV_X1    g0636(.A(new_n636), .ZN(new_n837));
  NAND4_X1  g0637(.A1(new_n837), .A2(new_n556), .A3(new_n502), .A4(new_n679), .ZN(new_n838));
  NAND2_X1  g0638(.A1(new_n836), .A2(new_n838), .ZN(new_n839));
  NAND2_X1  g0639(.A1(new_n450), .A2(new_n839), .ZN(new_n840));
  XNOR2_X1  g0640(.A(new_n840), .B(KEYINPUT103), .ZN(new_n841));
  OAI21_X1  g0641(.A(new_n642), .B1(new_n644), .B2(new_n645), .ZN(new_n842));
  NOR2_X1   g0642(.A1(new_n368), .A2(new_n676), .ZN(new_n843));
  NAND3_X1  g0643(.A1(new_n369), .A2(new_n370), .A3(new_n676), .ZN(new_n844));
  OAI21_X1  g0644(.A(new_n844), .B1(new_n382), .B2(new_n346), .ZN(new_n845));
  INV_X1    g0645(.A(KEYINPUT37), .ZN(new_n846));
  NAND3_X1  g0646(.A1(new_n356), .A2(new_n845), .A3(new_n846), .ZN(new_n847));
  INV_X1    g0647(.A(KEYINPUT99), .ZN(new_n848));
  NAND2_X1  g0648(.A1(new_n847), .A2(new_n848), .ZN(new_n849));
  NAND4_X1  g0649(.A1(new_n356), .A2(new_n845), .A3(KEYINPUT99), .A4(new_n846), .ZN(new_n850));
  NAND2_X1  g0650(.A1(new_n849), .A2(new_n850), .ZN(new_n851));
  NAND2_X1  g0651(.A1(new_n356), .A2(new_n845), .ZN(new_n852));
  NAND2_X1  g0652(.A1(new_n852), .A2(KEYINPUT37), .ZN(new_n853));
  AOI22_X1  g0653(.A1(new_n842), .A2(new_n843), .B1(new_n851), .B2(new_n853), .ZN(new_n854));
  OR2_X1    g0654(.A1(new_n854), .A2(KEYINPUT38), .ZN(new_n855));
  NOR2_X1   g0655(.A1(new_n330), .A2(KEYINPUT16), .ZN(new_n856));
  OAI221_X1 g0656(.A(new_n343), .B1(new_n251), .B2(new_n344), .C1(new_n856), .C2(new_n381), .ZN(new_n857));
  NAND2_X1  g0657(.A1(new_n857), .A2(new_n844), .ZN(new_n858));
  AOI21_X1  g0658(.A(new_n846), .B1(new_n858), .B2(new_n356), .ZN(new_n859));
  INV_X1    g0659(.A(new_n859), .ZN(new_n860));
  NAND2_X1  g0660(.A1(new_n851), .A2(new_n860), .ZN(new_n861));
  INV_X1    g0661(.A(new_n676), .ZN(new_n862));
  NAND3_X1  g0662(.A1(new_n384), .A2(new_n862), .A3(new_n857), .ZN(new_n863));
  NAND3_X1  g0663(.A1(new_n861), .A2(KEYINPUT38), .A3(new_n863), .ZN(new_n864));
  NAND2_X1  g0664(.A1(new_n855), .A2(new_n864), .ZN(new_n865));
  NOR2_X1   g0665(.A1(new_n404), .A2(new_n679), .ZN(new_n866));
  INV_X1    g0666(.A(new_n866), .ZN(new_n867));
  NOR2_X1   g0667(.A1(new_n429), .A2(new_n867), .ZN(new_n868));
  AOI211_X1 g0668(.A(new_n866), .B(new_n421), .C1(new_n427), .C2(new_n428), .ZN(new_n869));
  OAI21_X1  g0669(.A(new_n808), .B1(new_n868), .B2(new_n869), .ZN(new_n870));
  AOI21_X1  g0670(.A(new_n870), .B1(new_n836), .B2(new_n838), .ZN(new_n871));
  NAND3_X1  g0671(.A1(new_n865), .A2(KEYINPUT40), .A3(new_n871), .ZN(new_n872));
  INV_X1    g0672(.A(KEYINPUT38), .ZN(new_n873));
  AND3_X1   g0673(.A1(new_n384), .A2(new_n862), .A3(new_n857), .ZN(new_n874));
  AOI21_X1  g0674(.A(new_n859), .B1(new_n849), .B2(new_n850), .ZN(new_n875));
  OAI21_X1  g0675(.A(new_n873), .B1(new_n874), .B2(new_n875), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n876), .A2(new_n864), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n871), .A2(new_n877), .ZN(new_n878));
  INV_X1    g0678(.A(KEYINPUT40), .ZN(new_n879));
  AOI21_X1  g0679(.A(KEYINPUT102), .B1(new_n878), .B2(new_n879), .ZN(new_n880));
  INV_X1    g0680(.A(KEYINPUT102), .ZN(new_n881));
  AOI211_X1 g0681(.A(new_n881), .B(KEYINPUT40), .C1(new_n871), .C2(new_n877), .ZN(new_n882));
  OAI21_X1  g0682(.A(new_n872), .B1(new_n880), .B2(new_n882), .ZN(new_n883));
  XNOR2_X1  g0683(.A(new_n841), .B(new_n883), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n884), .A2(G330), .ZN(new_n885));
  NOR2_X1   g0685(.A1(new_n868), .A2(new_n869), .ZN(new_n886));
  INV_X1    g0686(.A(new_n886), .ZN(new_n887));
  AOI211_X1 g0687(.A(new_n678), .B(new_n807), .C1(new_n665), .C2(new_n668), .ZN(new_n888));
  OAI211_X1 g0688(.A(new_n877), .B(new_n887), .C1(new_n888), .C2(new_n805), .ZN(new_n889));
  NOR2_X1   g0689(.A1(new_n647), .A2(new_n862), .ZN(new_n890));
  INV_X1    g0690(.A(new_n890), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n889), .A2(new_n891), .ZN(new_n892));
  NOR2_X1   g0692(.A1(new_n639), .A2(new_n678), .ZN(new_n893));
  INV_X1    g0693(.A(new_n893), .ZN(new_n894));
  NOR3_X1   g0694(.A1(new_n874), .A2(new_n875), .A3(new_n873), .ZN(new_n895));
  AOI21_X1  g0695(.A(KEYINPUT38), .B1(new_n861), .B2(new_n863), .ZN(new_n896));
  OAI21_X1  g0696(.A(KEYINPUT39), .B1(new_n895), .B2(new_n896), .ZN(new_n897));
  XNOR2_X1  g0697(.A(KEYINPUT100), .B(KEYINPUT39), .ZN(new_n898));
  OAI211_X1 g0698(.A(new_n864), .B(new_n898), .C1(new_n854), .C2(KEYINPUT38), .ZN(new_n899));
  AOI21_X1  g0699(.A(new_n894), .B1(new_n897), .B2(new_n899), .ZN(new_n900));
  INV_X1    g0700(.A(KEYINPUT101), .ZN(new_n901));
  NOR3_X1   g0701(.A1(new_n892), .A2(new_n900), .A3(new_n901), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n897), .A2(new_n899), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n903), .A2(new_n893), .ZN(new_n904));
  INV_X1    g0704(.A(new_n658), .ZN(new_n905));
  NOR3_X1   g0705(.A1(new_n554), .A2(new_n555), .A3(new_n588), .ZN(new_n906));
  OAI21_X1  g0706(.A(new_n905), .B1(new_n906), .B2(new_n656), .ZN(new_n907));
  AND4_X1   g0707(.A1(new_n592), .A2(new_n666), .A3(new_n632), .A4(new_n667), .ZN(new_n908));
  OAI211_X1 g0708(.A(new_n679), .B(new_n808), .C1(new_n907), .C2(new_n908), .ZN(new_n909));
  AOI21_X1  g0709(.A(new_n886), .B1(new_n909), .B2(new_n806), .ZN(new_n910));
  AOI21_X1  g0710(.A(new_n890), .B1(new_n910), .B2(new_n877), .ZN(new_n911));
  AOI21_X1  g0711(.A(KEYINPUT101), .B1(new_n904), .B2(new_n911), .ZN(new_n912));
  NOR2_X1   g0712(.A1(new_n902), .A2(new_n912), .ZN(new_n913));
  XNOR2_X1  g0713(.A(new_n885), .B(new_n913), .ZN(new_n914));
  OAI21_X1  g0714(.A(new_n450), .B1(new_n710), .B2(new_n703), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n915), .A2(new_n649), .ZN(new_n916));
  XOR2_X1   g0716(.A(new_n914), .B(new_n916), .Z(new_n917));
  OAI21_X1  g0717(.A(new_n917), .B1(new_n261), .B2(new_n733), .ZN(new_n918));
  INV_X1    g0718(.A(KEYINPUT35), .ZN(new_n919));
  AOI211_X1 g0719(.A(new_n229), .B(new_n228), .C1(new_n565), .C2(new_n919), .ZN(new_n920));
  OAI211_X1 g0720(.A(new_n920), .B(G116), .C1(new_n919), .C2(new_n565), .ZN(new_n921));
  XNOR2_X1  g0721(.A(new_n921), .B(KEYINPUT36), .ZN(new_n922));
  OAI21_X1  g0722(.A(G77), .B1(new_n218), .B2(new_n207), .ZN(new_n923));
  OAI22_X1  g0723(.A1(new_n923), .A2(new_n231), .B1(G50), .B2(new_n207), .ZN(new_n924));
  NAND3_X1  g0724(.A1(new_n924), .A2(G1), .A3(new_n265), .ZN(new_n925));
  NAND3_X1  g0725(.A1(new_n918), .A2(new_n922), .A3(new_n925), .ZN(G367));
  NAND2_X1  g0726(.A1(new_n734), .A2(G1), .ZN(new_n927));
  OR2_X1    g0727(.A1(new_n691), .A2(KEYINPUT106), .ZN(new_n928));
  XOR2_X1   g0728(.A(new_n692), .B(new_n685), .Z(new_n929));
  NAND2_X1  g0729(.A1(new_n691), .A2(KEYINPUT106), .ZN(new_n930));
  NAND3_X1  g0730(.A1(new_n928), .A2(new_n929), .A3(new_n930), .ZN(new_n931));
  OAI21_X1  g0731(.A(new_n931), .B1(new_n929), .B2(new_n928), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n932), .A2(new_n729), .ZN(new_n933));
  OAI21_X1  g0733(.A(new_n592), .B1(new_n589), .B2(new_n679), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n655), .A2(new_n678), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n934), .A2(new_n935), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n686), .A2(new_n936), .ZN(new_n937));
  XNOR2_X1  g0737(.A(new_n937), .B(KEYINPUT45), .ZN(new_n938));
  OR3_X1    g0738(.A1(new_n686), .A2(KEYINPUT44), .A3(new_n936), .ZN(new_n939));
  OAI21_X1  g0739(.A(KEYINPUT44), .B1(new_n686), .B2(new_n936), .ZN(new_n940));
  NAND2_X1  g0740(.A1(new_n939), .A2(new_n940), .ZN(new_n941));
  NOR2_X1   g0741(.A1(new_n691), .A2(new_n693), .ZN(new_n942));
  OR3_X1    g0742(.A1(new_n938), .A2(new_n941), .A3(new_n942), .ZN(new_n943));
  OAI21_X1  g0743(.A(new_n942), .B1(new_n938), .B2(new_n941), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n943), .A2(new_n944), .ZN(new_n945));
  OAI21_X1  g0745(.A(new_n729), .B1(new_n933), .B2(new_n945), .ZN(new_n946));
  XNOR2_X1  g0746(.A(new_n696), .B(KEYINPUT41), .ZN(new_n947));
  AOI21_X1  g0747(.A(new_n927), .B1(new_n946), .B2(new_n947), .ZN(new_n948));
  NAND3_X1  g0748(.A1(new_n692), .A2(new_n685), .A3(new_n936), .ZN(new_n949));
  OR2_X1    g0749(.A1(new_n949), .A2(KEYINPUT42), .ZN(new_n950));
  NAND2_X1  g0750(.A1(new_n936), .A2(new_n681), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n663), .A2(new_n679), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n949), .A2(KEYINPUT42), .ZN(new_n953));
  NAND4_X1  g0753(.A1(new_n950), .A2(new_n951), .A3(new_n952), .A4(new_n953), .ZN(new_n954));
  OAI21_X1  g0754(.A(new_n667), .B1(new_n550), .B2(new_n679), .ZN(new_n955));
  OR3_X1    g0755(.A1(new_n544), .A2(new_n550), .A3(new_n679), .ZN(new_n956));
  NAND2_X1  g0756(.A1(new_n955), .A2(new_n956), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n957), .A2(KEYINPUT43), .ZN(new_n958));
  NAND2_X1  g0758(.A1(new_n954), .A2(new_n958), .ZN(new_n959));
  NAND2_X1  g0759(.A1(new_n959), .A2(KEYINPUT104), .ZN(new_n960));
  INV_X1    g0760(.A(KEYINPUT104), .ZN(new_n961));
  NAND3_X1  g0761(.A1(new_n954), .A2(new_n961), .A3(new_n958), .ZN(new_n962));
  NAND2_X1  g0762(.A1(new_n960), .A2(new_n962), .ZN(new_n963));
  OAI21_X1  g0763(.A(new_n963), .B1(KEYINPUT43), .B2(new_n957), .ZN(new_n964));
  NAND2_X1  g0764(.A1(new_n942), .A2(new_n936), .ZN(new_n965));
  OR2_X1    g0765(.A1(new_n965), .A2(KEYINPUT105), .ZN(new_n966));
  NOR2_X1   g0766(.A1(new_n957), .A2(KEYINPUT43), .ZN(new_n967));
  NAND3_X1  g0767(.A1(new_n960), .A2(new_n967), .A3(new_n962), .ZN(new_n968));
  AND3_X1   g0768(.A1(new_n964), .A2(new_n966), .A3(new_n968), .ZN(new_n969));
  NAND2_X1  g0769(.A1(new_n965), .A2(KEYINPUT105), .ZN(new_n970));
  AOI22_X1  g0770(.A1(new_n964), .A2(new_n968), .B1(new_n966), .B2(new_n970), .ZN(new_n971));
  NOR3_X1   g0771(.A1(new_n948), .A2(new_n969), .A3(new_n971), .ZN(new_n972));
  NAND3_X1  g0772(.A1(new_n955), .A2(new_n744), .A3(new_n956), .ZN(new_n973));
  OAI221_X1 g0773(.A(new_n278), .B1(new_n218), .B2(new_n777), .C1(new_n785), .C2(new_n821), .ZN(new_n974));
  AOI21_X1  g0774(.A(new_n974), .B1(G137), .B2(new_n789), .ZN(new_n975));
  INV_X1    g0775(.A(new_n768), .ZN(new_n976));
  AOI22_X1  g0776(.A1(G150), .A2(new_n760), .B1(new_n976), .B2(G68), .ZN(new_n977));
  XNOR2_X1  g0777(.A(new_n977), .B(KEYINPUT108), .ZN(new_n978));
  NAND2_X1  g0778(.A1(new_n772), .A2(G50), .ZN(new_n979));
  AOI22_X1  g0779(.A1(new_n765), .A2(G159), .B1(new_n814), .B2(G77), .ZN(new_n980));
  NAND4_X1  g0780(.A1(new_n975), .A2(new_n978), .A3(new_n979), .A4(new_n980), .ZN(new_n981));
  AOI22_X1  g0781(.A1(new_n760), .A2(G303), .B1(new_n775), .B2(G311), .ZN(new_n982));
  XNOR2_X1  g0782(.A(new_n982), .B(KEYINPUT107), .ZN(new_n983));
  NAND2_X1  g0783(.A1(new_n976), .A2(G107), .ZN(new_n984));
  AOI21_X1  g0784(.A(KEYINPUT46), .B1(new_n778), .B2(G116), .ZN(new_n985));
  AOI211_X1 g0785(.A(new_n328), .B(new_n985), .C1(new_n772), .C2(G283), .ZN(new_n986));
  NAND2_X1  g0786(.A1(new_n814), .A2(G97), .ZN(new_n987));
  OAI21_X1  g0787(.A(new_n987), .B1(new_n794), .B2(new_n784), .ZN(new_n988));
  AOI21_X1  g0788(.A(new_n988), .B1(new_n789), .B2(G317), .ZN(new_n989));
  NAND4_X1  g0789(.A1(new_n983), .A2(new_n984), .A3(new_n986), .A4(new_n989), .ZN(new_n990));
  AND3_X1   g0790(.A1(new_n778), .A2(KEYINPUT46), .A3(G116), .ZN(new_n991));
  OAI21_X1  g0791(.A(new_n981), .B1(new_n990), .B2(new_n991), .ZN(new_n992));
  XNOR2_X1  g0792(.A(new_n992), .B(KEYINPUT47), .ZN(new_n993));
  NAND2_X1  g0793(.A1(new_n993), .A2(new_n745), .ZN(new_n994));
  INV_X1    g0794(.A(new_n737), .ZN(new_n995));
  OAI221_X1 g0795(.A(new_n746), .B1(new_n224), .B2(new_n434), .C1(new_n240), .C2(new_n995), .ZN(new_n996));
  NAND4_X1  g0796(.A1(new_n973), .A2(new_n830), .A3(new_n994), .A4(new_n996), .ZN(new_n997));
  XNOR2_X1  g0797(.A(new_n997), .B(KEYINPUT109), .ZN(new_n998));
  OR2_X1    g0798(.A1(new_n972), .A2(new_n998), .ZN(G387));
  OR2_X1    g0799(.A1(new_n932), .A2(new_n729), .ZN(new_n1000));
  NAND3_X1  g0800(.A1(new_n1000), .A2(new_n696), .A3(new_n933), .ZN(new_n1001));
  INV_X1    g0801(.A(new_n744), .ZN(new_n1002));
  OAI21_X1  g0802(.A(new_n830), .B1(new_n692), .B2(new_n1002), .ZN(new_n1003));
  INV_X1    g0803(.A(new_n745), .ZN(new_n1004));
  AOI22_X1  g0804(.A1(new_n772), .A2(G303), .B1(G311), .B2(new_n765), .ZN(new_n1005));
  OAI21_X1  g0805(.A(new_n1005), .B1(new_n792), .B2(new_n785), .ZN(new_n1006));
  AOI21_X1  g0806(.A(new_n1006), .B1(G317), .B2(new_n760), .ZN(new_n1007));
  XOR2_X1   g0807(.A(new_n1007), .B(KEYINPUT48), .Z(new_n1008));
  OAI221_X1 g0808(.A(new_n1008), .B1(new_n791), .B2(new_n768), .C1(new_n784), .C2(new_n777), .ZN(new_n1009));
  XNOR2_X1  g0809(.A(new_n1009), .B(KEYINPUT49), .ZN(new_n1010));
  AOI21_X1  g0810(.A(new_n328), .B1(G116), .B2(new_n814), .ZN(new_n1011));
  OAI211_X1 g0811(.A(new_n1010), .B(new_n1011), .C1(new_n786), .C2(new_n754), .ZN(new_n1012));
  NOR2_X1   g0812(.A1(new_n434), .A2(new_n768), .ZN(new_n1013));
  AOI22_X1  g0813(.A1(G159), .A2(new_n775), .B1(new_n765), .B2(new_n431), .ZN(new_n1014));
  OAI221_X1 g0814(.A(new_n1014), .B1(new_n215), .B2(new_n777), .C1(new_n754), .C2(new_n257), .ZN(new_n1015));
  AOI211_X1 g0815(.A(new_n1013), .B(new_n1015), .C1(G68), .C2(new_n782), .ZN(new_n1016));
  NAND2_X1  g0816(.A1(new_n760), .A2(G50), .ZN(new_n1017));
  NAND4_X1  g0817(.A1(new_n1016), .A2(new_n328), .A3(new_n987), .A4(new_n1017), .ZN(new_n1018));
  AOI21_X1  g0818(.A(new_n1004), .B1(new_n1012), .B2(new_n1018), .ZN(new_n1019));
  NAND2_X1  g0819(.A1(new_n237), .A2(G45), .ZN(new_n1020));
  XNOR2_X1  g0820(.A(new_n1020), .B(KEYINPUT110), .ZN(new_n1021));
  NAND2_X1  g0821(.A1(new_n431), .A2(new_n213), .ZN(new_n1022));
  XNOR2_X1  g0822(.A(new_n1022), .B(KEYINPUT111), .ZN(new_n1023));
  XNOR2_X1  g0823(.A(new_n1023), .B(KEYINPUT50), .ZN(new_n1024));
  AOI21_X1  g0824(.A(G45), .B1(G68), .B2(G77), .ZN(new_n1025));
  NAND3_X1  g0825(.A1(new_n1024), .A2(new_n698), .A3(new_n1025), .ZN(new_n1026));
  NAND3_X1  g0826(.A1(new_n1021), .A2(new_n737), .A3(new_n1026), .ZN(new_n1027));
  OAI221_X1 g0827(.A(new_n1027), .B1(G107), .B2(new_n224), .C1(new_n698), .C2(new_n740), .ZN(new_n1028));
  AOI211_X1 g0828(.A(new_n1003), .B(new_n1019), .C1(new_n746), .C2(new_n1028), .ZN(new_n1029));
  AOI21_X1  g0829(.A(new_n1029), .B1(new_n932), .B2(new_n927), .ZN(new_n1030));
  NAND2_X1  g0830(.A1(new_n1001), .A2(new_n1030), .ZN(G393));
  AOI21_X1  g0831(.A(new_n697), .B1(new_n933), .B2(new_n945), .ZN(new_n1032));
  OAI21_X1  g0832(.A(new_n1032), .B1(new_n945), .B2(new_n933), .ZN(new_n1033));
  NAND3_X1  g0833(.A1(new_n934), .A2(new_n744), .A3(new_n935), .ZN(new_n1034));
  AOI22_X1  g0834(.A1(G116), .A2(new_n976), .B1(new_n765), .B2(G303), .ZN(new_n1035));
  OAI221_X1 g0835(.A(new_n1035), .B1(new_n209), .B2(new_n762), .C1(new_n784), .C2(new_n771), .ZN(new_n1036));
  AOI22_X1  g0836(.A1(new_n760), .A2(G311), .B1(new_n775), .B2(G317), .ZN(new_n1037));
  XOR2_X1   g0837(.A(new_n1037), .B(KEYINPUT52), .Z(new_n1038));
  OAI211_X1 g0838(.A(new_n1038), .B(new_n757), .C1(new_n792), .C2(new_n754), .ZN(new_n1039));
  AOI211_X1 g0839(.A(new_n1036), .B(new_n1039), .C1(G283), .C2(new_n778), .ZN(new_n1040));
  OAI22_X1  g0840(.A1(new_n761), .A2(new_n313), .B1(new_n785), .B2(new_n257), .ZN(new_n1041));
  INV_X1    g0841(.A(KEYINPUT51), .ZN(new_n1042));
  AOI22_X1  g0842(.A1(new_n1041), .A2(new_n1042), .B1(G87), .B2(new_n814), .ZN(new_n1043));
  OAI21_X1  g0843(.A(new_n1043), .B1(new_n1042), .B2(new_n1041), .ZN(new_n1044));
  AOI21_X1  g0844(.A(new_n377), .B1(new_n772), .B2(new_n431), .ZN(new_n1045));
  OAI221_X1 g0845(.A(new_n1045), .B1(new_n213), .B2(new_n794), .C1(new_n821), .C2(new_n754), .ZN(new_n1046));
  NOR2_X1   g0846(.A1(new_n768), .A2(new_n215), .ZN(new_n1047));
  NOR2_X1   g0847(.A1(new_n777), .A2(new_n207), .ZN(new_n1048));
  NOR4_X1   g0848(.A1(new_n1044), .A2(new_n1046), .A3(new_n1047), .A4(new_n1048), .ZN(new_n1049));
  OAI21_X1  g0849(.A(new_n745), .B1(new_n1040), .B2(new_n1049), .ZN(new_n1050));
  OAI221_X1 g0850(.A(new_n746), .B1(new_n516), .B2(new_n224), .C1(new_n995), .C2(new_n247), .ZN(new_n1051));
  NAND4_X1  g0851(.A1(new_n1034), .A2(new_n830), .A3(new_n1050), .A4(new_n1051), .ZN(new_n1052));
  INV_X1    g0852(.A(new_n927), .ZN(new_n1053));
  OAI211_X1 g0853(.A(new_n1033), .B(new_n1052), .C1(new_n1053), .C2(new_n945), .ZN(G390));
  NOR2_X1   g0854(.A1(new_n725), .A2(new_n870), .ZN(new_n1055));
  INV_X1    g0855(.A(new_n804), .ZN(new_n1056));
  NOR2_X1   g0856(.A1(new_n709), .A2(new_n1056), .ZN(new_n1057));
  NOR2_X1   g0857(.A1(new_n1057), .A2(new_n805), .ZN(new_n1058));
  OAI211_X1 g0858(.A(new_n894), .B(new_n865), .C1(new_n1058), .C2(new_n886), .ZN(new_n1059));
  OAI211_X1 g0859(.A(new_n897), .B(new_n899), .C1(new_n910), .C2(new_n893), .ZN(new_n1060));
  AOI21_X1  g0860(.A(new_n1055), .B1(new_n1059), .B2(new_n1060), .ZN(new_n1061));
  AND2_X1   g0861(.A1(new_n1059), .A2(new_n1060), .ZN(new_n1062));
  NAND3_X1  g0862(.A1(new_n726), .A2(new_n728), .A3(new_n808), .ZN(new_n1063));
  NOR2_X1   g0863(.A1(new_n1063), .A2(new_n886), .ZN(new_n1064));
  AOI21_X1  g0864(.A(new_n1061), .B1(new_n1062), .B2(new_n1064), .ZN(new_n1065));
  OAI21_X1  g0865(.A(new_n886), .B1(new_n725), .B2(new_n807), .ZN(new_n1066));
  OAI211_X1 g0866(.A(new_n1058), .B(new_n1066), .C1(new_n1063), .C2(new_n886), .ZN(new_n1067));
  AOI21_X1  g0867(.A(new_n1055), .B1(new_n1063), .B2(new_n886), .ZN(new_n1068));
  NOR2_X1   g0868(.A1(new_n888), .A2(new_n805), .ZN(new_n1069));
  OAI21_X1  g0869(.A(new_n1067), .B1(new_n1068), .B2(new_n1069), .ZN(new_n1070));
  INV_X1    g0870(.A(KEYINPUT112), .ZN(new_n1071));
  NAND3_X1  g0871(.A1(new_n450), .A2(G330), .A3(new_n839), .ZN(new_n1072));
  AND3_X1   g0872(.A1(new_n915), .A2(new_n1072), .A3(new_n649), .ZN(new_n1073));
  AND3_X1   g0873(.A1(new_n1070), .A2(new_n1071), .A3(new_n1073), .ZN(new_n1074));
  AOI21_X1  g0874(.A(new_n1071), .B1(new_n1070), .B2(new_n1073), .ZN(new_n1075));
  OAI21_X1  g0875(.A(new_n1065), .B1(new_n1074), .B2(new_n1075), .ZN(new_n1076));
  NAND2_X1  g0876(.A1(new_n1062), .A2(new_n1064), .ZN(new_n1077));
  OAI21_X1  g0877(.A(new_n1077), .B1(new_n1062), .B2(new_n1055), .ZN(new_n1078));
  NAND2_X1  g0878(.A1(new_n1070), .A2(new_n1073), .ZN(new_n1079));
  INV_X1    g0879(.A(new_n1079), .ZN(new_n1080));
  NAND2_X1  g0880(.A1(new_n1078), .A2(new_n1080), .ZN(new_n1081));
  NAND3_X1  g0881(.A1(new_n1076), .A2(new_n1081), .A3(new_n696), .ZN(new_n1082));
  NAND2_X1  g0882(.A1(new_n1078), .A2(new_n927), .ZN(new_n1083));
  INV_X1    g0883(.A(new_n903), .ZN(new_n1084));
  NAND2_X1  g0884(.A1(new_n832), .A2(new_n251), .ZN(new_n1085));
  AOI21_X1  g0885(.A(new_n278), .B1(new_n765), .B2(G107), .ZN(new_n1086));
  OAI211_X1 g0886(.A(new_n1086), .B(new_n779), .C1(new_n463), .C2(new_n761), .ZN(new_n1087));
  AOI21_X1  g0887(.A(new_n1047), .B1(G283), .B2(new_n775), .ZN(new_n1088));
  OAI221_X1 g0888(.A(new_n1088), .B1(new_n207), .B2(new_n762), .C1(new_n754), .C2(new_n784), .ZN(new_n1089));
  AOI211_X1 g0889(.A(new_n1087), .B(new_n1089), .C1(G97), .C2(new_n772), .ZN(new_n1090));
  XOR2_X1   g0890(.A(KEYINPUT54), .B(G143), .Z(new_n1091));
  AOI21_X1  g0891(.A(new_n757), .B1(new_n772), .B2(new_n1091), .ZN(new_n1092));
  OAI21_X1  g0892(.A(new_n1092), .B1(new_n313), .B2(new_n768), .ZN(new_n1093));
  AOI22_X1  g0893(.A1(new_n760), .A2(G132), .B1(new_n775), .B2(G128), .ZN(new_n1094));
  XOR2_X1   g0894(.A(new_n1094), .B(KEYINPUT113), .Z(new_n1095));
  NAND2_X1  g0895(.A1(new_n789), .A2(G125), .ZN(new_n1096));
  NOR2_X1   g0896(.A1(new_n777), .A2(new_n257), .ZN(new_n1097));
  XNOR2_X1  g0897(.A(new_n1097), .B(KEYINPUT53), .ZN(new_n1098));
  NAND3_X1  g0898(.A1(new_n1095), .A2(new_n1096), .A3(new_n1098), .ZN(new_n1099));
  AOI211_X1 g0899(.A(new_n1093), .B(new_n1099), .C1(G50), .C2(new_n814), .ZN(new_n1100));
  NAND2_X1  g0900(.A1(new_n765), .A2(G137), .ZN(new_n1101));
  AOI21_X1  g0901(.A(new_n1090), .B1(new_n1100), .B2(new_n1101), .ZN(new_n1102));
  OAI211_X1 g0902(.A(new_n830), .B(new_n1085), .C1(new_n1102), .C2(new_n1004), .ZN(new_n1103));
  AOI22_X1  g0903(.A1(new_n1084), .A2(new_n742), .B1(KEYINPUT114), .B2(new_n1103), .ZN(new_n1104));
  OAI21_X1  g0904(.A(new_n1104), .B1(KEYINPUT114), .B2(new_n1103), .ZN(new_n1105));
  NAND3_X1  g0905(.A1(new_n1082), .A2(new_n1083), .A3(new_n1105), .ZN(G378));
  OAI21_X1  g0906(.A(new_n1073), .B1(new_n1065), .B2(new_n1079), .ZN(new_n1107));
  OAI21_X1  g0907(.A(new_n901), .B1(new_n892), .B2(new_n900), .ZN(new_n1108));
  NAND3_X1  g0908(.A1(new_n904), .A2(new_n911), .A3(KEYINPUT101), .ZN(new_n1109));
  NAND2_X1  g0909(.A1(new_n270), .A2(new_n862), .ZN(new_n1110));
  XOR2_X1   g0910(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1111));
  NAND2_X1  g0911(.A1(new_n309), .A2(new_n1111), .ZN(new_n1112));
  INV_X1    g0912(.A(new_n1112), .ZN(new_n1113));
  NOR2_X1   g0913(.A1(new_n309), .A2(new_n1111), .ZN(new_n1114));
  OAI21_X1  g0914(.A(new_n1110), .B1(new_n1113), .B2(new_n1114), .ZN(new_n1115));
  INV_X1    g0915(.A(new_n1114), .ZN(new_n1116));
  INV_X1    g0916(.A(new_n1110), .ZN(new_n1117));
  NAND3_X1  g0917(.A1(new_n1116), .A2(new_n1117), .A3(new_n1112), .ZN(new_n1118));
  NAND2_X1  g0918(.A1(new_n1115), .A2(new_n1118), .ZN(new_n1119));
  AND3_X1   g0919(.A1(new_n1108), .A2(new_n1109), .A3(new_n1119), .ZN(new_n1120));
  AOI21_X1  g0920(.A(new_n1119), .B1(new_n1108), .B2(new_n1109), .ZN(new_n1121));
  OAI211_X1 g0921(.A(G330), .B(new_n872), .C1(new_n880), .C2(new_n882), .ZN(new_n1122));
  NOR3_X1   g0922(.A1(new_n1120), .A2(new_n1121), .A3(new_n1122), .ZN(new_n1123));
  INV_X1    g0923(.A(new_n1122), .ZN(new_n1124));
  INV_X1    g0924(.A(new_n1119), .ZN(new_n1125));
  OAI21_X1  g0925(.A(new_n1125), .B1(new_n902), .B2(new_n912), .ZN(new_n1126));
  NAND3_X1  g0926(.A1(new_n1108), .A2(new_n1109), .A3(new_n1119), .ZN(new_n1127));
  AOI21_X1  g0927(.A(new_n1124), .B1(new_n1126), .B2(new_n1127), .ZN(new_n1128));
  OAI211_X1 g0928(.A(new_n1107), .B(KEYINPUT57), .C1(new_n1123), .C2(new_n1128), .ZN(new_n1129));
  INV_X1    g0929(.A(KEYINPUT118), .ZN(new_n1130));
  OAI21_X1  g0930(.A(new_n1130), .B1(new_n1123), .B2(new_n1128), .ZN(new_n1131));
  OAI21_X1  g0931(.A(new_n1122), .B1(new_n1120), .B2(new_n1121), .ZN(new_n1132));
  NAND3_X1  g0932(.A1(new_n1126), .A2(new_n1124), .A3(new_n1127), .ZN(new_n1133));
  NAND3_X1  g0933(.A1(new_n1132), .A2(KEYINPUT118), .A3(new_n1133), .ZN(new_n1134));
  AOI22_X1  g0934(.A1(new_n1131), .A2(new_n1134), .B1(new_n1081), .B2(new_n1073), .ZN(new_n1135));
  OAI211_X1 g0935(.A(new_n696), .B(new_n1129), .C1(new_n1135), .C2(KEYINPUT57), .ZN(new_n1136));
  AOI21_X1  g0936(.A(new_n1053), .B1(new_n1131), .B2(new_n1134), .ZN(new_n1137));
  INV_X1    g0937(.A(KEYINPUT119), .ZN(new_n1138));
  NOR2_X1   g0938(.A1(new_n1125), .A2(new_n743), .ZN(new_n1139));
  AOI22_X1  g0939(.A1(new_n765), .A2(G97), .B1(new_n782), .B2(new_n433), .ZN(new_n1140));
  XNOR2_X1  g0940(.A(new_n1140), .B(KEYINPUT116), .ZN(new_n1141));
  AOI22_X1  g0941(.A1(new_n760), .A2(G107), .B1(G58), .B2(new_n814), .ZN(new_n1142));
  OAI211_X1 g0942(.A(new_n1141), .B(new_n1142), .C1(new_n207), .C2(new_n768), .ZN(new_n1143));
  AOI21_X1  g0943(.A(new_n1143), .B1(G116), .B2(new_n775), .ZN(new_n1144));
  AOI211_X1 g0944(.A(G41), .B(new_n328), .C1(G77), .C2(new_n778), .ZN(new_n1145));
  OAI211_X1 g0945(.A(new_n1144), .B(new_n1145), .C1(new_n791), .C2(new_n754), .ZN(new_n1146));
  XNOR2_X1  g0946(.A(new_n1146), .B(KEYINPUT58), .ZN(new_n1147));
  AOI22_X1  g0947(.A1(G150), .A2(new_n976), .B1(new_n775), .B2(G125), .ZN(new_n1148));
  NAND2_X1  g0948(.A1(new_n760), .A2(G128), .ZN(new_n1149));
  NAND2_X1  g0949(.A1(new_n782), .A2(G137), .ZN(new_n1150));
  AOI22_X1  g0950(.A1(new_n765), .A2(G132), .B1(new_n778), .B2(new_n1091), .ZN(new_n1151));
  NAND4_X1  g0951(.A1(new_n1148), .A2(new_n1149), .A3(new_n1150), .A4(new_n1151), .ZN(new_n1152));
  NOR2_X1   g0952(.A1(new_n1152), .A2(KEYINPUT59), .ZN(new_n1153));
  NOR2_X1   g0953(.A1(new_n1153), .A2(G33), .ZN(new_n1154));
  NAND2_X1  g0954(.A1(new_n1152), .A2(KEYINPUT59), .ZN(new_n1155));
  NAND2_X1  g0955(.A1(new_n814), .A2(G159), .ZN(new_n1156));
  AOI21_X1  g0956(.A(G41), .B1(new_n789), .B2(G124), .ZN(new_n1157));
  NAND4_X1  g0957(.A1(new_n1154), .A2(new_n1155), .A3(new_n1156), .A4(new_n1157), .ZN(new_n1158));
  AOI21_X1  g0958(.A(G50), .B1(new_n324), .B2(new_n283), .ZN(new_n1159));
  XOR2_X1   g0959(.A(new_n1159), .B(KEYINPUT115), .Z(new_n1160));
  NAND3_X1  g0960(.A1(new_n1147), .A2(new_n1158), .A3(new_n1160), .ZN(new_n1161));
  AND2_X1   g0961(.A1(new_n1161), .A2(new_n745), .ZN(new_n1162));
  AOI21_X1  g0962(.A(new_n735), .B1(new_n213), .B2(new_n832), .ZN(new_n1163));
  XNOR2_X1  g0963(.A(new_n1163), .B(KEYINPUT117), .ZN(new_n1164));
  NOR3_X1   g0964(.A1(new_n1139), .A2(new_n1162), .A3(new_n1164), .ZN(new_n1165));
  NOR3_X1   g0965(.A1(new_n1137), .A2(new_n1138), .A3(new_n1165), .ZN(new_n1166));
  AND3_X1   g0966(.A1(new_n1132), .A2(KEYINPUT118), .A3(new_n1133), .ZN(new_n1167));
  AOI21_X1  g0967(.A(KEYINPUT118), .B1(new_n1132), .B2(new_n1133), .ZN(new_n1168));
  OAI21_X1  g0968(.A(new_n927), .B1(new_n1167), .B2(new_n1168), .ZN(new_n1169));
  INV_X1    g0969(.A(new_n1165), .ZN(new_n1170));
  AOI21_X1  g0970(.A(KEYINPUT119), .B1(new_n1169), .B2(new_n1170), .ZN(new_n1171));
  OAI21_X1  g0971(.A(new_n1136), .B1(new_n1166), .B2(new_n1171), .ZN(G375));
  XOR2_X1   g0972(.A(new_n927), .B(KEYINPUT120), .Z(new_n1173));
  NAND2_X1  g0973(.A1(new_n1070), .A2(new_n1173), .ZN(new_n1174));
  XNOR2_X1  g0974(.A(new_n1174), .B(KEYINPUT121), .ZN(new_n1175));
  OAI21_X1  g0975(.A(new_n757), .B1(new_n794), .B2(new_n463), .ZN(new_n1176));
  AOI21_X1  g0976(.A(new_n1013), .B1(G283), .B2(new_n760), .ZN(new_n1177));
  XNOR2_X1  g0977(.A(new_n1177), .B(KEYINPUT122), .ZN(new_n1178));
  OAI221_X1 g0978(.A(new_n1178), .B1(new_n215), .B2(new_n762), .C1(new_n209), .C2(new_n773), .ZN(new_n1179));
  AOI211_X1 g0979(.A(new_n1176), .B(new_n1179), .C1(G303), .C2(new_n789), .ZN(new_n1180));
  OAI221_X1 g0980(.A(new_n1180), .B1(new_n516), .B2(new_n777), .C1(new_n784), .C2(new_n785), .ZN(new_n1181));
  AOI22_X1  g0981(.A1(new_n789), .A2(G128), .B1(G159), .B2(new_n778), .ZN(new_n1182));
  XNOR2_X1  g0982(.A(new_n1182), .B(KEYINPUT123), .ZN(new_n1183));
  AOI21_X1  g0983(.A(new_n1183), .B1(G58), .B2(new_n814), .ZN(new_n1184));
  AOI21_X1  g0984(.A(new_n377), .B1(new_n976), .B2(G50), .ZN(new_n1185));
  OAI211_X1 g0985(.A(new_n1184), .B(new_n1185), .C1(new_n257), .C2(new_n771), .ZN(new_n1186));
  XNOR2_X1  g0986(.A(new_n1186), .B(KEYINPUT124), .ZN(new_n1187));
  NAND2_X1  g0987(.A1(new_n765), .A2(new_n1091), .ZN(new_n1188));
  NAND2_X1  g0988(.A1(new_n760), .A2(G137), .ZN(new_n1189));
  NAND3_X1  g0989(.A1(new_n1187), .A2(new_n1188), .A3(new_n1189), .ZN(new_n1190));
  NOR2_X1   g0990(.A1(new_n785), .A2(new_n826), .ZN(new_n1191));
  OAI21_X1  g0991(.A(new_n1181), .B1(new_n1190), .B2(new_n1191), .ZN(new_n1192));
  AOI22_X1  g0992(.A1(new_n1192), .A2(new_n745), .B1(new_n207), .B2(new_n832), .ZN(new_n1193));
  OAI211_X1 g0993(.A(new_n1193), .B(new_n830), .C1(new_n743), .C2(new_n887), .ZN(new_n1194));
  NAND2_X1  g0994(.A1(new_n1175), .A2(new_n1194), .ZN(new_n1195));
  OR2_X1    g0995(.A1(new_n1074), .A2(new_n1075), .ZN(new_n1196));
  OR2_X1    g0996(.A1(new_n1070), .A2(new_n1073), .ZN(new_n1197));
  AND2_X1   g0997(.A1(new_n1196), .A2(new_n1197), .ZN(new_n1198));
  AOI21_X1  g0998(.A(new_n1195), .B1(new_n1198), .B2(new_n947), .ZN(new_n1199));
  INV_X1    g0999(.A(new_n1199), .ZN(G381));
  OAI21_X1  g1000(.A(new_n1107), .B1(new_n1167), .B2(new_n1168), .ZN(new_n1201));
  INV_X1    g1001(.A(KEYINPUT57), .ZN(new_n1202));
  AOI21_X1  g1002(.A(new_n697), .B1(new_n1201), .B2(new_n1202), .ZN(new_n1203));
  OAI21_X1  g1003(.A(new_n1138), .B1(new_n1137), .B2(new_n1165), .ZN(new_n1204));
  NAND3_X1  g1004(.A1(new_n1169), .A2(KEYINPUT119), .A3(new_n1170), .ZN(new_n1205));
  AOI22_X1  g1005(.A1(new_n1129), .A2(new_n1203), .B1(new_n1204), .B2(new_n1205), .ZN(new_n1206));
  INV_X1    g1006(.A(G378), .ZN(new_n1207));
  NAND2_X1  g1007(.A1(new_n1206), .A2(new_n1207), .ZN(new_n1208));
  INV_X1    g1008(.A(new_n1208), .ZN(new_n1209));
  INV_X1    g1009(.A(G384), .ZN(new_n1210));
  OR3_X1    g1010(.A1(new_n972), .A2(G390), .A3(new_n998), .ZN(new_n1211));
  NOR3_X1   g1011(.A1(new_n1211), .A2(G396), .A3(G393), .ZN(new_n1212));
  NAND4_X1  g1012(.A1(new_n1209), .A2(new_n1210), .A3(new_n1199), .A4(new_n1212), .ZN(G407));
  NAND2_X1  g1013(.A1(new_n677), .A2(G213), .ZN(new_n1214));
  INV_X1    g1014(.A(new_n1214), .ZN(new_n1215));
  NAND3_X1  g1015(.A1(new_n1209), .A2(KEYINPUT125), .A3(new_n1215), .ZN(new_n1216));
  INV_X1    g1016(.A(KEYINPUT125), .ZN(new_n1217));
  OAI21_X1  g1017(.A(new_n1217), .B1(new_n1208), .B2(new_n1214), .ZN(new_n1218));
  NAND4_X1  g1018(.A1(G407), .A2(new_n1216), .A3(G213), .A4(new_n1218), .ZN(G409));
  INV_X1    g1019(.A(KEYINPUT127), .ZN(new_n1220));
  NAND2_X1  g1020(.A1(G387), .A2(G390), .ZN(new_n1221));
  XNOR2_X1  g1021(.A(G393), .B(G396), .ZN(new_n1222));
  AND3_X1   g1022(.A1(new_n1221), .A2(new_n1211), .A3(new_n1222), .ZN(new_n1223));
  AOI21_X1  g1023(.A(new_n1222), .B1(new_n1221), .B2(new_n1211), .ZN(new_n1224));
  NOR2_X1   g1024(.A1(new_n1223), .A2(new_n1224), .ZN(new_n1225));
  AND2_X1   g1025(.A1(new_n1175), .A2(new_n1194), .ZN(new_n1226));
  INV_X1    g1026(.A(KEYINPUT60), .ZN(new_n1227));
  NAND2_X1  g1027(.A1(new_n1197), .A2(new_n1227), .ZN(new_n1228));
  OR3_X1    g1028(.A1(new_n1070), .A2(new_n1073), .A3(new_n1227), .ZN(new_n1229));
  NAND4_X1  g1029(.A1(new_n1228), .A2(new_n696), .A3(new_n1079), .A4(new_n1229), .ZN(new_n1230));
  AOI21_X1  g1030(.A(G384), .B1(new_n1226), .B2(new_n1230), .ZN(new_n1231));
  AND4_X1   g1031(.A1(G384), .A2(new_n1230), .A3(new_n1194), .A4(new_n1175), .ZN(new_n1232));
  OAI21_X1  g1032(.A(KEYINPUT126), .B1(new_n1231), .B2(new_n1232), .ZN(new_n1233));
  INV_X1    g1033(.A(new_n1230), .ZN(new_n1234));
  OAI21_X1  g1034(.A(new_n1210), .B1(new_n1234), .B2(new_n1195), .ZN(new_n1235));
  NAND3_X1  g1035(.A1(new_n1226), .A2(G384), .A3(new_n1230), .ZN(new_n1236));
  INV_X1    g1036(.A(KEYINPUT126), .ZN(new_n1237));
  NAND3_X1  g1037(.A1(new_n1235), .A2(new_n1236), .A3(new_n1237), .ZN(new_n1238));
  AOI22_X1  g1038(.A1(new_n1233), .A2(new_n1238), .B1(G2897), .B2(new_n1215), .ZN(new_n1239));
  AOI21_X1  g1039(.A(new_n1215), .B1(G375), .B2(G378), .ZN(new_n1240));
  NAND2_X1  g1040(.A1(new_n1135), .A2(new_n947), .ZN(new_n1241));
  OAI21_X1  g1041(.A(new_n1173), .B1(new_n1123), .B2(new_n1128), .ZN(new_n1242));
  NAND4_X1  g1042(.A1(new_n1207), .A2(new_n1241), .A3(new_n1170), .A4(new_n1242), .ZN(new_n1243));
  AOI21_X1  g1043(.A(new_n1239), .B1(new_n1240), .B2(new_n1243), .ZN(new_n1244));
  NAND3_X1  g1044(.A1(new_n1238), .A2(G2897), .A3(new_n1215), .ZN(new_n1245));
  NAND2_X1  g1045(.A1(G375), .A2(G378), .ZN(new_n1246));
  NAND2_X1  g1046(.A1(new_n1235), .A2(new_n1236), .ZN(new_n1247));
  INV_X1    g1047(.A(new_n1247), .ZN(new_n1248));
  NAND4_X1  g1048(.A1(new_n1246), .A2(new_n1214), .A3(new_n1248), .A4(new_n1243), .ZN(new_n1249));
  AOI22_X1  g1049(.A1(new_n1244), .A2(new_n1245), .B1(new_n1249), .B2(KEYINPUT62), .ZN(new_n1250));
  NAND2_X1  g1050(.A1(new_n1204), .A2(new_n1205), .ZN(new_n1251));
  AOI21_X1  g1051(.A(new_n1207), .B1(new_n1251), .B2(new_n1136), .ZN(new_n1252));
  AND4_X1   g1052(.A1(new_n1207), .A2(new_n1241), .A3(new_n1170), .A4(new_n1242), .ZN(new_n1253));
  NOR4_X1   g1053(.A1(new_n1252), .A2(new_n1253), .A3(new_n1215), .A4(new_n1247), .ZN(new_n1254));
  INV_X1    g1054(.A(KEYINPUT62), .ZN(new_n1255));
  AOI21_X1  g1055(.A(KEYINPUT61), .B1(new_n1254), .B2(new_n1255), .ZN(new_n1256));
  AOI21_X1  g1056(.A(new_n1225), .B1(new_n1250), .B2(new_n1256), .ZN(new_n1257));
  OAI211_X1 g1057(.A(new_n1214), .B(new_n1243), .C1(new_n1206), .C2(new_n1207), .ZN(new_n1258));
  NAND2_X1  g1058(.A1(new_n1233), .A2(new_n1238), .ZN(new_n1259));
  NAND2_X1  g1059(.A1(new_n1215), .A2(G2897), .ZN(new_n1260));
  NAND2_X1  g1060(.A1(new_n1259), .A2(new_n1260), .ZN(new_n1261));
  NAND3_X1  g1061(.A1(new_n1258), .A2(new_n1245), .A3(new_n1261), .ZN(new_n1262));
  AOI21_X1  g1062(.A(new_n1254), .B1(new_n1262), .B2(KEYINPUT63), .ZN(new_n1263));
  NAND4_X1  g1063(.A1(new_n1240), .A2(KEYINPUT63), .A3(new_n1248), .A4(new_n1243), .ZN(new_n1264));
  INV_X1    g1064(.A(KEYINPUT61), .ZN(new_n1265));
  NAND3_X1  g1065(.A1(new_n1264), .A2(new_n1225), .A3(new_n1265), .ZN(new_n1266));
  NOR2_X1   g1066(.A1(new_n1263), .A2(new_n1266), .ZN(new_n1267));
  OAI21_X1  g1067(.A(new_n1220), .B1(new_n1257), .B2(new_n1267), .ZN(new_n1268));
  AND3_X1   g1068(.A1(new_n1264), .A2(new_n1265), .A3(new_n1225), .ZN(new_n1269));
  AND2_X1   g1069(.A1(new_n1262), .A2(KEYINPUT63), .ZN(new_n1270));
  OAI21_X1  g1070(.A(new_n1269), .B1(new_n1270), .B2(new_n1254), .ZN(new_n1271));
  NAND2_X1  g1071(.A1(new_n1249), .A2(KEYINPUT62), .ZN(new_n1272));
  NAND4_X1  g1072(.A1(new_n1240), .A2(new_n1255), .A3(new_n1248), .A4(new_n1243), .ZN(new_n1273));
  NAND4_X1  g1073(.A1(new_n1272), .A2(new_n1262), .A3(new_n1265), .A4(new_n1273), .ZN(new_n1274));
  INV_X1    g1074(.A(new_n1225), .ZN(new_n1275));
  NAND2_X1  g1075(.A1(new_n1274), .A2(new_n1275), .ZN(new_n1276));
  NAND3_X1  g1076(.A1(new_n1271), .A2(new_n1276), .A3(KEYINPUT127), .ZN(new_n1277));
  NAND2_X1  g1077(.A1(new_n1268), .A2(new_n1277), .ZN(G405));
  NAND2_X1  g1078(.A1(new_n1208), .A2(new_n1246), .ZN(new_n1279));
  XNOR2_X1  g1079(.A(new_n1225), .B(new_n1279), .ZN(new_n1280));
  XNOR2_X1  g1080(.A(new_n1280), .B(new_n1248), .ZN(G402));
endmodule


