//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 0 0 0 1 1 0 0 1 0 0 1 0 1 0 0 1 1 0 1 0 1 1 0 0 0 1 1 1 1 0 1 1 0 0 1 1 1 0 1 1 0 0 1 0 1 1 1 1 1 0 1 1 1 0 0 1 1 1 0 0 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:26:11 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n691, new_n692,
    new_n693, new_n694, new_n695, new_n696, new_n697, new_n699, new_n700,
    new_n701, new_n702, new_n703, new_n704, new_n705, new_n706, new_n707,
    new_n708, new_n709, new_n710, new_n711, new_n712, new_n713, new_n714,
    new_n716, new_n717, new_n718, new_n719, new_n720, new_n721, new_n722,
    new_n723, new_n724, new_n725, new_n726, new_n727, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n746, new_n747, new_n748, new_n749, new_n750, new_n751, new_n752,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n760, new_n762,
    new_n763, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n793, new_n794, new_n795, new_n796, new_n797, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n819, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n966,
    new_n967, new_n968, new_n969, new_n970, new_n971, new_n972, new_n973,
    new_n974, new_n975, new_n976, new_n977, new_n978, new_n979, new_n980,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1014, new_n1015, new_n1016,
    new_n1017, new_n1018, new_n1019, new_n1020, new_n1021, new_n1022,
    new_n1023, new_n1024, new_n1025, new_n1027, new_n1028, new_n1029,
    new_n1030, new_n1031, new_n1033, new_n1034, new_n1035, new_n1036,
    new_n1037, new_n1038, new_n1039, new_n1040, new_n1041, new_n1042,
    new_n1043, new_n1044, new_n1045, new_n1046, new_n1047, new_n1048,
    new_n1049, new_n1050, new_n1051, new_n1053, new_n1054, new_n1055,
    new_n1056, new_n1057, new_n1058, new_n1059, new_n1060, new_n1061,
    new_n1062, new_n1063, new_n1064, new_n1065, new_n1066;
  NOR2_X1   g000(.A1(G472), .A2(G902), .ZN(new_n187));
  XNOR2_X1  g001(.A(KEYINPUT2), .B(G113), .ZN(new_n188));
  INV_X1    g002(.A(KEYINPUT64), .ZN(new_n189));
  INV_X1    g003(.A(G116), .ZN(new_n190));
  NOR2_X1   g004(.A1(new_n190), .A2(G119), .ZN(new_n191));
  INV_X1    g005(.A(G119), .ZN(new_n192));
  NOR2_X1   g006(.A1(new_n192), .A2(G116), .ZN(new_n193));
  OAI211_X1 g007(.A(new_n188), .B(new_n189), .C1(new_n191), .C2(new_n193), .ZN(new_n194));
  INV_X1    g008(.A(G113), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n195), .A2(KEYINPUT2), .ZN(new_n196));
  INV_X1    g010(.A(KEYINPUT2), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n197), .A2(G113), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n196), .A2(new_n198), .ZN(new_n199));
  XNOR2_X1  g013(.A(G116), .B(G119), .ZN(new_n200));
  OAI21_X1  g014(.A(new_n199), .B1(new_n200), .B2(KEYINPUT64), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n194), .A2(new_n201), .ZN(new_n202));
  INV_X1    g016(.A(G146), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n203), .A2(G143), .ZN(new_n204));
  INV_X1    g018(.A(G143), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n205), .A2(G146), .ZN(new_n206));
  AND2_X1   g020(.A1(KEYINPUT0), .A2(G128), .ZN(new_n207));
  NAND3_X1  g021(.A1(new_n204), .A2(new_n206), .A3(new_n207), .ZN(new_n208));
  XNOR2_X1  g022(.A(G143), .B(G146), .ZN(new_n209));
  XNOR2_X1  g023(.A(KEYINPUT0), .B(G128), .ZN(new_n210));
  OAI21_X1  g024(.A(new_n208), .B1(new_n209), .B2(new_n210), .ZN(new_n211));
  INV_X1    g025(.A(KEYINPUT11), .ZN(new_n212));
  INV_X1    g026(.A(G134), .ZN(new_n213));
  OAI21_X1  g027(.A(new_n212), .B1(new_n213), .B2(G137), .ZN(new_n214));
  INV_X1    g028(.A(G137), .ZN(new_n215));
  NAND3_X1  g029(.A1(new_n215), .A2(KEYINPUT11), .A3(G134), .ZN(new_n216));
  INV_X1    g030(.A(G131), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n213), .A2(G137), .ZN(new_n218));
  NAND4_X1  g032(.A1(new_n214), .A2(new_n216), .A3(new_n217), .A4(new_n218), .ZN(new_n219));
  NAND3_X1  g033(.A1(new_n214), .A2(new_n216), .A3(new_n218), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n220), .A2(G131), .ZN(new_n221));
  AOI21_X1  g035(.A(new_n211), .B1(new_n219), .B2(new_n221), .ZN(new_n222));
  OAI21_X1  g036(.A(KEYINPUT1), .B1(new_n205), .B2(G146), .ZN(new_n223));
  NOR2_X1   g037(.A1(new_n205), .A2(G146), .ZN(new_n224));
  NOR2_X1   g038(.A1(new_n203), .A2(G143), .ZN(new_n225));
  OAI211_X1 g039(.A(G128), .B(new_n223), .C1(new_n224), .C2(new_n225), .ZN(new_n226));
  INV_X1    g040(.A(G128), .ZN(new_n227));
  OAI211_X1 g041(.A(new_n204), .B(new_n206), .C1(KEYINPUT1), .C2(new_n227), .ZN(new_n228));
  NOR2_X1   g042(.A1(new_n213), .A2(G137), .ZN(new_n229));
  NOR2_X1   g043(.A1(new_n215), .A2(G134), .ZN(new_n230));
  OAI21_X1  g044(.A(G131), .B1(new_n229), .B2(new_n230), .ZN(new_n231));
  AND4_X1   g045(.A1(new_n219), .A2(new_n226), .A3(new_n228), .A4(new_n231), .ZN(new_n232));
  NOR3_X1   g046(.A1(new_n222), .A2(new_n232), .A3(KEYINPUT30), .ZN(new_n233));
  INV_X1    g047(.A(KEYINPUT30), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n221), .A2(new_n219), .ZN(new_n235));
  INV_X1    g049(.A(new_n211), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n235), .A2(new_n236), .ZN(new_n237));
  NAND4_X1  g051(.A1(new_n226), .A2(new_n219), .A3(new_n231), .A4(new_n228), .ZN(new_n238));
  AOI21_X1  g052(.A(new_n234), .B1(new_n237), .B2(new_n238), .ZN(new_n239));
  OAI21_X1  g053(.A(new_n202), .B1(new_n233), .B2(new_n239), .ZN(new_n240));
  INV_X1    g054(.A(G237), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n241), .A2(KEYINPUT65), .ZN(new_n242));
  INV_X1    g056(.A(KEYINPUT65), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n243), .A2(G237), .ZN(new_n244));
  AOI21_X1  g058(.A(G953), .B1(new_n242), .B2(new_n244), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n245), .A2(G210), .ZN(new_n246));
  XNOR2_X1  g060(.A(new_n246), .B(KEYINPUT27), .ZN(new_n247));
  XNOR2_X1  g061(.A(KEYINPUT26), .B(G101), .ZN(new_n248));
  INV_X1    g062(.A(new_n248), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n247), .A2(new_n249), .ZN(new_n250));
  OR2_X1    g064(.A1(new_n246), .A2(KEYINPUT27), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n246), .A2(KEYINPUT27), .ZN(new_n252));
  NAND3_X1  g066(.A1(new_n251), .A2(new_n252), .A3(new_n248), .ZN(new_n253));
  AND2_X1   g067(.A1(new_n250), .A2(new_n253), .ZN(new_n254));
  INV_X1    g068(.A(new_n202), .ZN(new_n255));
  NAND3_X1  g069(.A1(new_n237), .A2(new_n238), .A3(new_n255), .ZN(new_n256));
  NAND3_X1  g070(.A1(new_n240), .A2(new_n254), .A3(new_n256), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n257), .A2(KEYINPUT31), .ZN(new_n258));
  NOR3_X1   g072(.A1(new_n222), .A2(new_n232), .A3(new_n202), .ZN(new_n259));
  OAI21_X1  g073(.A(KEYINPUT30), .B1(new_n222), .B2(new_n232), .ZN(new_n260));
  NAND3_X1  g074(.A1(new_n237), .A2(new_n234), .A3(new_n238), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n260), .A2(new_n261), .ZN(new_n262));
  AOI21_X1  g076(.A(new_n259), .B1(new_n262), .B2(new_n202), .ZN(new_n263));
  INV_X1    g077(.A(KEYINPUT31), .ZN(new_n264));
  NAND3_X1  g078(.A1(new_n263), .A2(new_n264), .A3(new_n254), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n258), .A2(new_n265), .ZN(new_n266));
  NOR2_X1   g080(.A1(new_n259), .A2(KEYINPUT28), .ZN(new_n267));
  INV_X1    g081(.A(KEYINPUT66), .ZN(new_n268));
  INV_X1    g082(.A(KEYINPUT28), .ZN(new_n269));
  OAI21_X1  g083(.A(new_n202), .B1(new_n222), .B2(new_n232), .ZN(new_n270));
  AOI21_X1  g084(.A(new_n269), .B1(new_n270), .B2(new_n256), .ZN(new_n271));
  AOI21_X1  g085(.A(new_n267), .B1(new_n268), .B2(new_n271), .ZN(new_n272));
  NAND2_X1  g086(.A1(new_n270), .A2(new_n256), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n273), .A2(KEYINPUT28), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n274), .A2(KEYINPUT66), .ZN(new_n275));
  AOI21_X1  g089(.A(new_n254), .B1(new_n272), .B2(new_n275), .ZN(new_n276));
  OAI21_X1  g090(.A(new_n187), .B1(new_n266), .B2(new_n276), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n277), .A2(KEYINPUT67), .ZN(new_n278));
  INV_X1    g092(.A(KEYINPUT32), .ZN(new_n279));
  INV_X1    g093(.A(new_n254), .ZN(new_n280));
  NAND3_X1  g094(.A1(new_n273), .A2(new_n268), .A3(KEYINPUT28), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n256), .A2(new_n269), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n281), .A2(new_n282), .ZN(new_n283));
  NOR2_X1   g097(.A1(new_n271), .A2(new_n268), .ZN(new_n284));
  OAI21_X1  g098(.A(new_n280), .B1(new_n283), .B2(new_n284), .ZN(new_n285));
  NAND3_X1  g099(.A1(new_n285), .A2(new_n258), .A3(new_n265), .ZN(new_n286));
  INV_X1    g100(.A(KEYINPUT67), .ZN(new_n287));
  NAND3_X1  g101(.A1(new_n286), .A2(new_n287), .A3(new_n187), .ZN(new_n288));
  NAND3_X1  g102(.A1(new_n278), .A2(new_n279), .A3(new_n288), .ZN(new_n289));
  INV_X1    g103(.A(KEYINPUT68), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n289), .A2(new_n290), .ZN(new_n291));
  NAND4_X1  g105(.A1(new_n278), .A2(new_n288), .A3(KEYINPUT68), .A4(new_n279), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n291), .A2(new_n292), .ZN(new_n293));
  NAND3_X1  g107(.A1(new_n286), .A2(KEYINPUT32), .A3(new_n187), .ZN(new_n294));
  INV_X1    g108(.A(KEYINPUT70), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n294), .A2(new_n295), .ZN(new_n296));
  NAND3_X1  g110(.A1(new_n250), .A2(new_n253), .A3(KEYINPUT29), .ZN(new_n297));
  NOR3_X1   g111(.A1(new_n267), .A2(new_n271), .A3(new_n297), .ZN(new_n298));
  OAI21_X1  g112(.A(KEYINPUT69), .B1(new_n298), .B2(G902), .ZN(new_n299));
  INV_X1    g113(.A(KEYINPUT69), .ZN(new_n300));
  INV_X1    g114(.A(G902), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n274), .A2(new_n282), .ZN(new_n302));
  OAI211_X1 g116(.A(new_n300), .B(new_n301), .C1(new_n302), .C2(new_n297), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n299), .A2(new_n303), .ZN(new_n304));
  INV_X1    g118(.A(KEYINPUT29), .ZN(new_n305));
  OAI21_X1  g119(.A(new_n305), .B1(new_n263), .B2(new_n254), .ZN(new_n306));
  NOR2_X1   g120(.A1(new_n283), .A2(new_n284), .ZN(new_n307));
  AOI21_X1  g121(.A(new_n306), .B1(new_n307), .B2(new_n254), .ZN(new_n308));
  OAI21_X1  g122(.A(G472), .B1(new_n304), .B2(new_n308), .ZN(new_n309));
  NAND4_X1  g123(.A1(new_n286), .A2(KEYINPUT70), .A3(KEYINPUT32), .A4(new_n187), .ZN(new_n310));
  NAND3_X1  g124(.A1(new_n296), .A2(new_n309), .A3(new_n310), .ZN(new_n311));
  INV_X1    g125(.A(new_n311), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n293), .A2(new_n312), .ZN(new_n313));
  INV_X1    g127(.A(KEYINPUT78), .ZN(new_n314));
  XNOR2_X1  g128(.A(G110), .B(G140), .ZN(new_n315));
  INV_X1    g129(.A(G227), .ZN(new_n316));
  NOR2_X1   g130(.A1(new_n316), .A2(G953), .ZN(new_n317));
  XNOR2_X1  g131(.A(new_n315), .B(new_n317), .ZN(new_n318));
  INV_X1    g132(.A(new_n235), .ZN(new_n319));
  INV_X1    g133(.A(G104), .ZN(new_n320));
  NOR3_X1   g134(.A1(new_n320), .A2(KEYINPUT3), .A3(G107), .ZN(new_n321));
  INV_X1    g135(.A(G107), .ZN(new_n322));
  NOR2_X1   g136(.A1(new_n322), .A2(G104), .ZN(new_n323));
  NOR2_X1   g137(.A1(new_n321), .A2(new_n323), .ZN(new_n324));
  INV_X1    g138(.A(G101), .ZN(new_n325));
  OAI21_X1  g139(.A(KEYINPUT3), .B1(new_n320), .B2(G107), .ZN(new_n326));
  NAND4_X1  g140(.A1(new_n324), .A2(KEYINPUT75), .A3(new_n325), .A4(new_n326), .ZN(new_n327));
  INV_X1    g141(.A(KEYINPUT3), .ZN(new_n328));
  NAND3_X1  g142(.A1(new_n328), .A2(new_n322), .A3(G104), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n320), .A2(G107), .ZN(new_n330));
  NAND4_X1  g144(.A1(new_n326), .A2(new_n329), .A3(new_n325), .A4(new_n330), .ZN(new_n331));
  INV_X1    g145(.A(KEYINPUT75), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n331), .A2(new_n332), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n327), .A2(new_n333), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n322), .A2(G104), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n335), .A2(new_n330), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n336), .A2(G101), .ZN(new_n337));
  NAND3_X1  g151(.A1(new_n226), .A2(new_n337), .A3(new_n228), .ZN(new_n338));
  INV_X1    g152(.A(new_n338), .ZN(new_n339));
  AND3_X1   g153(.A1(new_n334), .A2(new_n339), .A3(KEYINPUT10), .ZN(new_n340));
  AOI21_X1  g154(.A(KEYINPUT10), .B1(new_n334), .B2(new_n339), .ZN(new_n341));
  NOR2_X1   g155(.A1(new_n340), .A2(new_n341), .ZN(new_n342));
  INV_X1    g156(.A(KEYINPUT4), .ZN(new_n343));
  NAND3_X1  g157(.A1(new_n326), .A2(new_n329), .A3(new_n330), .ZN(new_n344));
  AOI21_X1  g158(.A(new_n343), .B1(new_n344), .B2(G101), .ZN(new_n345));
  AND2_X1   g159(.A1(new_n331), .A2(new_n332), .ZN(new_n346));
  NOR2_X1   g160(.A1(new_n331), .A2(new_n332), .ZN(new_n347));
  OAI21_X1  g161(.A(new_n345), .B1(new_n346), .B2(new_n347), .ZN(new_n348));
  NAND3_X1  g162(.A1(new_n344), .A2(new_n343), .A3(G101), .ZN(new_n349));
  NAND3_X1  g163(.A1(new_n348), .A2(new_n236), .A3(new_n349), .ZN(new_n350));
  AOI21_X1  g164(.A(new_n319), .B1(new_n342), .B2(new_n350), .ZN(new_n351));
  INV_X1    g165(.A(KEYINPUT10), .ZN(new_n352));
  NOR2_X1   g166(.A1(new_n346), .A2(new_n347), .ZN(new_n353));
  OAI21_X1  g167(.A(new_n352), .B1(new_n353), .B2(new_n338), .ZN(new_n354));
  NAND3_X1  g168(.A1(new_n334), .A2(new_n339), .A3(KEYINPUT10), .ZN(new_n355));
  AND4_X1   g169(.A1(new_n319), .A2(new_n350), .A3(new_n354), .A4(new_n355), .ZN(new_n356));
  OAI21_X1  g170(.A(new_n318), .B1(new_n351), .B2(new_n356), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n357), .A2(KEYINPUT77), .ZN(new_n358));
  NAND4_X1  g172(.A1(new_n350), .A2(new_n354), .A3(new_n319), .A4(new_n355), .ZN(new_n359));
  INV_X1    g173(.A(new_n318), .ZN(new_n360));
  NAND2_X1  g174(.A1(new_n359), .A2(new_n360), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n361), .A2(KEYINPUT76), .ZN(new_n362));
  INV_X1    g176(.A(new_n337), .ZN(new_n363));
  AOI21_X1  g177(.A(new_n363), .B1(new_n327), .B2(new_n333), .ZN(new_n364));
  AND2_X1   g178(.A1(new_n226), .A2(new_n228), .ZN(new_n365));
  OAI22_X1  g179(.A1(new_n353), .A2(new_n338), .B1(new_n364), .B2(new_n365), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n366), .A2(new_n235), .ZN(new_n367));
  INV_X1    g181(.A(KEYINPUT12), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n367), .A2(new_n368), .ZN(new_n369));
  NAND3_X1  g183(.A1(new_n366), .A2(KEYINPUT12), .A3(new_n235), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n369), .A2(new_n370), .ZN(new_n371));
  INV_X1    g185(.A(KEYINPUT76), .ZN(new_n372));
  NAND3_X1  g186(.A1(new_n359), .A2(new_n372), .A3(new_n360), .ZN(new_n373));
  NAND3_X1  g187(.A1(new_n362), .A2(new_n371), .A3(new_n373), .ZN(new_n374));
  INV_X1    g188(.A(KEYINPUT77), .ZN(new_n375));
  OAI211_X1 g189(.A(new_n375), .B(new_n318), .C1(new_n351), .C2(new_n356), .ZN(new_n376));
  NAND3_X1  g190(.A1(new_n358), .A2(new_n374), .A3(new_n376), .ZN(new_n377));
  INV_X1    g191(.A(G469), .ZN(new_n378));
  NAND3_X1  g192(.A1(new_n377), .A2(new_n378), .A3(new_n301), .ZN(new_n379));
  NOR2_X1   g193(.A1(new_n361), .A2(new_n351), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n371), .A2(new_n359), .ZN(new_n381));
  XOR2_X1   g195(.A(new_n318), .B(KEYINPUT74), .Z(new_n382));
  AOI21_X1  g196(.A(new_n380), .B1(new_n381), .B2(new_n382), .ZN(new_n383));
  OAI21_X1  g197(.A(G469), .B1(new_n383), .B2(G902), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n379), .A2(new_n384), .ZN(new_n385));
  INV_X1    g199(.A(G221), .ZN(new_n386));
  XNOR2_X1  g200(.A(KEYINPUT9), .B(G234), .ZN(new_n387));
  INV_X1    g201(.A(new_n387), .ZN(new_n388));
  AOI21_X1  g202(.A(new_n386), .B1(new_n388), .B2(new_n301), .ZN(new_n389));
  INV_X1    g203(.A(new_n389), .ZN(new_n390));
  AOI21_X1  g204(.A(new_n314), .B1(new_n385), .B2(new_n390), .ZN(new_n391));
  AOI211_X1 g205(.A(KEYINPUT78), .B(new_n389), .C1(new_n379), .C2(new_n384), .ZN(new_n392));
  NOR2_X1   g206(.A1(new_n391), .A2(new_n392), .ZN(new_n393));
  INV_X1    g207(.A(G234), .ZN(new_n394));
  OAI21_X1  g208(.A(G217), .B1(new_n394), .B2(G902), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n395), .A2(new_n301), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n192), .A2(G128), .ZN(new_n397));
  NAND3_X1  g211(.A1(new_n227), .A2(KEYINPUT23), .A3(G119), .ZN(new_n398));
  NOR2_X1   g212(.A1(new_n192), .A2(G128), .ZN(new_n399));
  OAI211_X1 g213(.A(new_n397), .B(new_n398), .C1(new_n399), .C2(KEYINPUT23), .ZN(new_n400));
  XOR2_X1   g214(.A(KEYINPUT24), .B(G110), .Z(new_n401));
  XNOR2_X1  g215(.A(G119), .B(G128), .ZN(new_n402));
  AOI22_X1  g216(.A1(new_n400), .A2(G110), .B1(new_n401), .B2(new_n402), .ZN(new_n403));
  INV_X1    g217(.A(G140), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n404), .A2(G125), .ZN(new_n405));
  INV_X1    g219(.A(G125), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n406), .A2(G140), .ZN(new_n407));
  NAND3_X1  g221(.A1(new_n405), .A2(new_n407), .A3(KEYINPUT16), .ZN(new_n408));
  OR3_X1    g222(.A1(new_n406), .A2(KEYINPUT16), .A3(G140), .ZN(new_n409));
  NAND2_X1  g223(.A1(new_n408), .A2(new_n409), .ZN(new_n410));
  NOR2_X1   g224(.A1(new_n410), .A2(new_n203), .ZN(new_n411));
  AOI21_X1  g225(.A(G146), .B1(new_n408), .B2(new_n409), .ZN(new_n412));
  OAI21_X1  g226(.A(new_n403), .B1(new_n411), .B2(new_n412), .ZN(new_n413));
  AND3_X1   g227(.A1(new_n405), .A2(new_n407), .A3(new_n203), .ZN(new_n414));
  NOR3_X1   g228(.A1(new_n406), .A2(KEYINPUT16), .A3(G140), .ZN(new_n415));
  XNOR2_X1  g229(.A(G125), .B(G140), .ZN(new_n416));
  AOI21_X1  g230(.A(new_n415), .B1(new_n416), .B2(KEYINPUT16), .ZN(new_n417));
  AOI21_X1  g231(.A(new_n414), .B1(new_n417), .B2(G146), .ZN(new_n418));
  OAI22_X1  g232(.A1(new_n400), .A2(G110), .B1(new_n401), .B2(new_n402), .ZN(new_n419));
  NAND2_X1  g233(.A1(new_n418), .A2(new_n419), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n413), .A2(new_n420), .ZN(new_n421));
  XNOR2_X1  g235(.A(KEYINPUT22), .B(G137), .ZN(new_n422));
  INV_X1    g236(.A(G953), .ZN(new_n423));
  NAND3_X1  g237(.A1(new_n423), .A2(G221), .A3(G234), .ZN(new_n424));
  INV_X1    g238(.A(new_n424), .ZN(new_n425));
  OR2_X1    g239(.A1(new_n422), .A2(new_n425), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n422), .A2(new_n425), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n426), .A2(new_n427), .ZN(new_n428));
  INV_X1    g242(.A(KEYINPUT71), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n428), .A2(new_n429), .ZN(new_n430));
  XNOR2_X1  g244(.A(new_n422), .B(new_n424), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n431), .A2(KEYINPUT71), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n430), .A2(new_n432), .ZN(new_n433));
  INV_X1    g247(.A(KEYINPUT72), .ZN(new_n434));
  NAND3_X1  g248(.A1(new_n421), .A2(new_n433), .A3(new_n434), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n417), .A2(G146), .ZN(new_n436));
  NAND2_X1  g250(.A1(new_n410), .A2(new_n203), .ZN(new_n437));
  NAND2_X1  g251(.A1(new_n436), .A2(new_n437), .ZN(new_n438));
  AOI22_X1  g252(.A1(new_n438), .A2(new_n403), .B1(new_n418), .B2(new_n419), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n439), .A2(new_n431), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n435), .A2(new_n440), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n421), .A2(new_n433), .ZN(new_n442));
  AOI211_X1 g256(.A(new_n396), .B(new_n441), .C1(KEYINPUT72), .C2(new_n442), .ZN(new_n443));
  AND3_X1   g257(.A1(new_n426), .A2(new_n427), .A3(KEYINPUT71), .ZN(new_n444));
  AOI21_X1  g258(.A(KEYINPUT71), .B1(new_n426), .B2(new_n427), .ZN(new_n445));
  NOR2_X1   g259(.A1(new_n444), .A2(new_n445), .ZN(new_n446));
  OAI21_X1  g260(.A(KEYINPUT72), .B1(new_n439), .B2(new_n446), .ZN(new_n447));
  NAND4_X1  g261(.A1(new_n447), .A2(new_n301), .A3(new_n435), .A4(new_n440), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n448), .A2(KEYINPUT73), .ZN(new_n449));
  INV_X1    g263(.A(KEYINPUT25), .ZN(new_n450));
  AOI21_X1  g264(.A(new_n395), .B1(new_n449), .B2(new_n450), .ZN(new_n451));
  NAND3_X1  g265(.A1(new_n448), .A2(KEYINPUT73), .A3(KEYINPUT25), .ZN(new_n452));
  AOI21_X1  g266(.A(new_n443), .B1(new_n451), .B2(new_n452), .ZN(new_n453));
  OAI21_X1  g267(.A(G214), .B1(G237), .B2(G902), .ZN(new_n454));
  XNOR2_X1  g268(.A(G110), .B(G122), .ZN(new_n455));
  INV_X1    g269(.A(new_n455), .ZN(new_n456));
  AND2_X1   g270(.A1(new_n344), .A2(G101), .ZN(new_n457));
  AOI22_X1  g271(.A1(new_n457), .A2(new_n343), .B1(new_n194), .B2(new_n201), .ZN(new_n458));
  AND3_X1   g272(.A1(new_n348), .A2(new_n458), .A3(KEYINPUT79), .ZN(new_n459));
  AOI21_X1  g273(.A(KEYINPUT79), .B1(new_n348), .B2(new_n458), .ZN(new_n460));
  NOR2_X1   g274(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n200), .A2(KEYINPUT5), .ZN(new_n462));
  INV_X1    g276(.A(KEYINPUT5), .ZN(new_n463));
  AOI21_X1  g277(.A(new_n195), .B1(new_n191), .B2(new_n463), .ZN(new_n464));
  AOI22_X1  g278(.A1(new_n462), .A2(new_n464), .B1(new_n199), .B2(new_n200), .ZN(new_n465));
  NAND2_X1  g279(.A1(new_n364), .A2(new_n465), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n466), .A2(KEYINPUT80), .ZN(new_n467));
  INV_X1    g281(.A(KEYINPUT80), .ZN(new_n468));
  NAND3_X1  g282(.A1(new_n364), .A2(new_n468), .A3(new_n465), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n467), .A2(new_n469), .ZN(new_n470));
  OAI21_X1  g284(.A(new_n456), .B1(new_n461), .B2(new_n470), .ZN(new_n471));
  INV_X1    g285(.A(KEYINPUT79), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n344), .A2(G101), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n473), .A2(KEYINPUT4), .ZN(new_n474));
  AOI21_X1  g288(.A(new_n474), .B1(new_n333), .B2(new_n327), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n202), .A2(new_n349), .ZN(new_n476));
  OAI21_X1  g290(.A(new_n472), .B1(new_n475), .B2(new_n476), .ZN(new_n477));
  NAND3_X1  g291(.A1(new_n348), .A2(new_n458), .A3(KEYINPUT79), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  AND3_X1   g293(.A1(new_n364), .A2(new_n468), .A3(new_n465), .ZN(new_n480));
  AOI21_X1  g294(.A(new_n468), .B1(new_n364), .B2(new_n465), .ZN(new_n481));
  NOR2_X1   g295(.A1(new_n480), .A2(new_n481), .ZN(new_n482));
  NAND3_X1  g296(.A1(new_n479), .A2(new_n482), .A3(new_n455), .ZN(new_n483));
  NAND3_X1  g297(.A1(new_n471), .A2(KEYINPUT6), .A3(new_n483), .ZN(new_n484));
  OR3_X1    g298(.A1(new_n236), .A2(KEYINPUT83), .A3(new_n406), .ZN(new_n485));
  OAI21_X1  g299(.A(KEYINPUT83), .B1(new_n236), .B2(new_n406), .ZN(new_n486));
  OAI211_X1 g300(.A(new_n485), .B(new_n486), .C1(G125), .C2(new_n365), .ZN(new_n487));
  INV_X1    g301(.A(G224), .ZN(new_n488));
  NOR2_X1   g302(.A1(new_n488), .A2(G953), .ZN(new_n489));
  XNOR2_X1  g303(.A(new_n489), .B(KEYINPUT84), .ZN(new_n490));
  XNOR2_X1  g304(.A(new_n487), .B(new_n490), .ZN(new_n491));
  INV_X1    g305(.A(KEYINPUT6), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n492), .A2(KEYINPUT81), .ZN(new_n493));
  OR2_X1    g307(.A1(new_n492), .A2(KEYINPUT81), .ZN(new_n494));
  AOI21_X1  g308(.A(new_n455), .B1(new_n493), .B2(new_n494), .ZN(new_n495));
  INV_X1    g309(.A(new_n495), .ZN(new_n496));
  AOI211_X1 g310(.A(KEYINPUT82), .B(new_n496), .C1(new_n479), .C2(new_n482), .ZN(new_n497));
  INV_X1    g311(.A(KEYINPUT82), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n479), .A2(new_n482), .ZN(new_n499));
  AOI21_X1  g313(.A(new_n498), .B1(new_n499), .B2(new_n495), .ZN(new_n500));
  OAI211_X1 g314(.A(new_n484), .B(new_n491), .C1(new_n497), .C2(new_n500), .ZN(new_n501));
  OAI21_X1  g315(.A(KEYINPUT7), .B1(new_n488), .B2(G953), .ZN(new_n502));
  NOR2_X1   g316(.A1(new_n365), .A2(G125), .ZN(new_n503));
  NOR2_X1   g317(.A1(new_n236), .A2(new_n406), .ZN(new_n504));
  OAI21_X1  g318(.A(new_n502), .B1(new_n503), .B2(new_n504), .ZN(new_n505));
  OAI21_X1  g319(.A(new_n505), .B1(new_n487), .B2(new_n502), .ZN(new_n506));
  NOR2_X1   g320(.A1(new_n461), .A2(new_n470), .ZN(new_n507));
  AOI21_X1  g321(.A(new_n506), .B1(new_n507), .B2(new_n455), .ZN(new_n508));
  XNOR2_X1  g322(.A(new_n455), .B(KEYINPUT8), .ZN(new_n509));
  NOR2_X1   g323(.A1(new_n364), .A2(new_n465), .ZN(new_n510));
  INV_X1    g324(.A(KEYINPUT85), .ZN(new_n511));
  AOI21_X1  g325(.A(new_n510), .B1(new_n511), .B2(new_n466), .ZN(new_n512));
  NOR3_X1   g326(.A1(new_n364), .A2(KEYINPUT85), .A3(new_n465), .ZN(new_n513));
  OAI21_X1  g327(.A(new_n509), .B1(new_n512), .B2(new_n513), .ZN(new_n514));
  AOI21_X1  g328(.A(G902), .B1(new_n508), .B2(new_n514), .ZN(new_n515));
  OAI21_X1  g329(.A(G210), .B1(G237), .B2(G902), .ZN(new_n516));
  AND3_X1   g330(.A1(new_n501), .A2(new_n515), .A3(new_n516), .ZN(new_n517));
  AOI21_X1  g331(.A(new_n516), .B1(new_n501), .B2(new_n515), .ZN(new_n518));
  OAI21_X1  g332(.A(new_n454), .B1(new_n517), .B2(new_n518), .ZN(new_n519));
  NAND3_X1  g333(.A1(new_n388), .A2(G217), .A3(new_n423), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n190), .A2(G122), .ZN(new_n521));
  NOR2_X1   g335(.A1(new_n521), .A2(KEYINPUT14), .ZN(new_n522));
  INV_X1    g336(.A(KEYINPUT14), .ZN(new_n523));
  OAI21_X1  g337(.A(new_n523), .B1(new_n190), .B2(G122), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n524), .A2(new_n521), .ZN(new_n525));
  AOI21_X1  g339(.A(new_n522), .B1(new_n525), .B2(KEYINPUT95), .ZN(new_n526));
  INV_X1    g340(.A(KEYINPUT95), .ZN(new_n527));
  NAND3_X1  g341(.A1(new_n524), .A2(new_n527), .A3(new_n521), .ZN(new_n528));
  AOI21_X1  g342(.A(new_n322), .B1(new_n526), .B2(new_n528), .ZN(new_n529));
  INV_X1    g343(.A(G122), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n530), .A2(G116), .ZN(new_n531));
  NAND3_X1  g345(.A1(new_n531), .A2(new_n521), .A3(new_n322), .ZN(new_n532));
  INV_X1    g346(.A(KEYINPUT94), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  NAND4_X1  g348(.A1(new_n531), .A2(new_n521), .A3(KEYINPUT94), .A4(new_n322), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n205), .A2(G128), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n227), .A2(G143), .ZN(new_n537));
  NAND3_X1  g351(.A1(new_n536), .A2(new_n537), .A3(new_n213), .ZN(new_n538));
  INV_X1    g352(.A(new_n538), .ZN(new_n539));
  AOI21_X1  g353(.A(new_n213), .B1(new_n536), .B2(new_n537), .ZN(new_n540));
  OAI211_X1 g354(.A(new_n534), .B(new_n535), .C1(new_n539), .C2(new_n540), .ZN(new_n541));
  NOR2_X1   g355(.A1(new_n529), .A2(new_n541), .ZN(new_n542));
  INV_X1    g356(.A(new_n532), .ZN(new_n543));
  AOI21_X1  g357(.A(new_n322), .B1(new_n531), .B2(new_n521), .ZN(new_n544));
  OAI21_X1  g358(.A(new_n538), .B1(new_n543), .B2(new_n544), .ZN(new_n545));
  INV_X1    g359(.A(new_n537), .ZN(new_n546));
  AND2_X1   g360(.A1(KEYINPUT92), .A2(KEYINPUT13), .ZN(new_n547));
  NOR2_X1   g361(.A1(KEYINPUT92), .A2(KEYINPUT13), .ZN(new_n548));
  NOR2_X1   g362(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  AOI21_X1  g363(.A(new_n546), .B1(new_n549), .B2(new_n536), .ZN(new_n550));
  NOR2_X1   g364(.A1(new_n227), .A2(G143), .ZN(new_n551));
  OAI21_X1  g365(.A(new_n551), .B1(new_n547), .B2(new_n548), .ZN(new_n552));
  INV_X1    g366(.A(KEYINPUT93), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n552), .A2(new_n553), .ZN(new_n554));
  OAI211_X1 g368(.A(new_n551), .B(KEYINPUT93), .C1(new_n548), .C2(new_n547), .ZN(new_n555));
  NAND3_X1  g369(.A1(new_n550), .A2(new_n554), .A3(new_n555), .ZN(new_n556));
  AOI21_X1  g370(.A(new_n545), .B1(new_n556), .B2(G134), .ZN(new_n557));
  OAI21_X1  g371(.A(new_n520), .B1(new_n542), .B2(new_n557), .ZN(new_n558));
  INV_X1    g372(.A(new_n548), .ZN(new_n559));
  NAND2_X1  g373(.A1(KEYINPUT92), .A2(KEYINPUT13), .ZN(new_n560));
  NAND3_X1  g374(.A1(new_n559), .A2(new_n536), .A3(new_n560), .ZN(new_n561));
  NAND3_X1  g375(.A1(new_n555), .A2(new_n561), .A3(new_n537), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n559), .A2(new_n560), .ZN(new_n563));
  AOI21_X1  g377(.A(KEYINPUT93), .B1(new_n563), .B2(new_n551), .ZN(new_n564));
  OAI21_X1  g378(.A(G134), .B1(new_n562), .B2(new_n564), .ZN(new_n565));
  INV_X1    g379(.A(new_n545), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n565), .A2(new_n566), .ZN(new_n567));
  AOI21_X1  g381(.A(KEYINPUT14), .B1(new_n530), .B2(G116), .ZN(new_n568));
  NOR2_X1   g382(.A1(new_n530), .A2(G116), .ZN(new_n569));
  OAI21_X1  g383(.A(KEYINPUT95), .B1(new_n568), .B2(new_n569), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n569), .A2(new_n523), .ZN(new_n571));
  NAND3_X1  g385(.A1(new_n570), .A2(new_n528), .A3(new_n571), .ZN(new_n572));
  NAND2_X1  g386(.A1(new_n572), .A2(G107), .ZN(new_n573));
  INV_X1    g387(.A(new_n540), .ZN(new_n574));
  AOI22_X1  g388(.A1(new_n574), .A2(new_n538), .B1(new_n533), .B2(new_n532), .ZN(new_n575));
  NAND3_X1  g389(.A1(new_n573), .A2(new_n575), .A3(new_n535), .ZN(new_n576));
  INV_X1    g390(.A(new_n520), .ZN(new_n577));
  NAND3_X1  g391(.A1(new_n567), .A2(new_n576), .A3(new_n577), .ZN(new_n578));
  NAND3_X1  g392(.A1(new_n558), .A2(KEYINPUT96), .A3(new_n578), .ZN(new_n579));
  INV_X1    g393(.A(KEYINPUT96), .ZN(new_n580));
  NAND4_X1  g394(.A1(new_n567), .A2(new_n576), .A3(new_n580), .A4(new_n577), .ZN(new_n581));
  NAND3_X1  g395(.A1(new_n579), .A2(new_n301), .A3(new_n581), .ZN(new_n582));
  NAND2_X1  g396(.A1(new_n582), .A2(KEYINPUT97), .ZN(new_n583));
  INV_X1    g397(.A(KEYINPUT97), .ZN(new_n584));
  NAND4_X1  g398(.A1(new_n579), .A2(new_n584), .A3(new_n301), .A4(new_n581), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n583), .A2(new_n585), .ZN(new_n586));
  INV_X1    g400(.A(G478), .ZN(new_n587));
  NOR2_X1   g401(.A1(new_n587), .A2(KEYINPUT15), .ZN(new_n588));
  NAND2_X1  g402(.A1(new_n586), .A2(new_n588), .ZN(new_n589));
  AOI21_X1  g403(.A(new_n588), .B1(new_n582), .B2(KEYINPUT97), .ZN(new_n590));
  INV_X1    g404(.A(new_n590), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n589), .A2(new_n591), .ZN(new_n592));
  AND2_X1   g406(.A1(new_n423), .A2(G952), .ZN(new_n593));
  NAND2_X1  g407(.A1(G234), .A2(G237), .ZN(new_n594));
  NAND2_X1  g408(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  INV_X1    g409(.A(new_n595), .ZN(new_n596));
  NAND3_X1  g410(.A1(new_n594), .A2(G902), .A3(G953), .ZN(new_n597));
  INV_X1    g411(.A(new_n597), .ZN(new_n598));
  XNOR2_X1  g412(.A(KEYINPUT21), .B(G898), .ZN(new_n599));
  AOI21_X1  g413(.A(new_n596), .B1(new_n598), .B2(new_n599), .ZN(new_n600));
  OR2_X1    g414(.A1(new_n592), .A2(new_n600), .ZN(new_n601));
  INV_X1    g415(.A(KEYINPUT20), .ZN(new_n602));
  NOR2_X1   g416(.A1(G475), .A2(G902), .ZN(new_n603));
  XOR2_X1   g417(.A(G113), .B(G122), .Z(new_n604));
  XOR2_X1   g418(.A(KEYINPUT88), .B(G104), .Z(new_n605));
  XOR2_X1   g419(.A(new_n604), .B(new_n605), .Z(new_n606));
  NOR2_X1   g420(.A1(new_n243), .A2(G237), .ZN(new_n607));
  NOR2_X1   g421(.A1(new_n241), .A2(KEYINPUT65), .ZN(new_n608));
  OAI211_X1 g422(.A(G214), .B(new_n423), .C1(new_n607), .C2(new_n608), .ZN(new_n609));
  NOR2_X1   g423(.A1(new_n609), .A2(new_n205), .ZN(new_n610));
  AOI21_X1  g424(.A(G143), .B1(new_n245), .B2(G214), .ZN(new_n611));
  OAI211_X1 g425(.A(KEYINPUT18), .B(G131), .C1(new_n610), .C2(new_n611), .ZN(new_n612));
  INV_X1    g426(.A(KEYINPUT86), .ZN(new_n613));
  AOI21_X1  g427(.A(new_n613), .B1(new_n416), .B2(new_n203), .ZN(new_n614));
  NOR2_X1   g428(.A1(new_n416), .A2(new_n203), .ZN(new_n615));
  XNOR2_X1  g429(.A(new_n614), .B(new_n615), .ZN(new_n616));
  NAND2_X1  g430(.A1(new_n609), .A2(new_n205), .ZN(new_n617));
  NAND3_X1  g431(.A1(new_n245), .A2(G143), .A3(G214), .ZN(new_n618));
  NAND2_X1  g432(.A1(KEYINPUT18), .A2(G131), .ZN(new_n619));
  NAND3_X1  g433(.A1(new_n617), .A2(new_n618), .A3(new_n619), .ZN(new_n620));
  AND3_X1   g434(.A1(new_n612), .A2(new_n616), .A3(new_n620), .ZN(new_n621));
  OAI211_X1 g435(.A(KEYINPUT17), .B(G131), .C1(new_n610), .C2(new_n611), .ZN(new_n622));
  INV_X1    g436(.A(KEYINPUT89), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  NAND2_X1  g438(.A1(new_n617), .A2(new_n618), .ZN(new_n625));
  NAND4_X1  g439(.A1(new_n625), .A2(KEYINPUT89), .A3(KEYINPUT17), .A4(G131), .ZN(new_n626));
  AOI21_X1  g440(.A(new_n438), .B1(new_n624), .B2(new_n626), .ZN(new_n627));
  INV_X1    g441(.A(KEYINPUT87), .ZN(new_n628));
  OAI21_X1  g442(.A(new_n628), .B1(new_n625), .B2(G131), .ZN(new_n629));
  INV_X1    g443(.A(KEYINPUT17), .ZN(new_n630));
  NAND4_X1  g444(.A1(new_n617), .A2(KEYINPUT87), .A3(new_n618), .A4(new_n217), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n625), .A2(G131), .ZN(new_n632));
  NAND4_X1  g446(.A1(new_n629), .A2(new_n630), .A3(new_n631), .A4(new_n632), .ZN(new_n633));
  AOI211_X1 g447(.A(new_n606), .B(new_n621), .C1(new_n627), .C2(new_n633), .ZN(new_n634));
  INV_X1    g448(.A(new_n606), .ZN(new_n635));
  NAND3_X1  g449(.A1(new_n629), .A2(new_n631), .A3(new_n632), .ZN(new_n636));
  XNOR2_X1  g450(.A(new_n416), .B(KEYINPUT19), .ZN(new_n637));
  AOI21_X1  g451(.A(new_n411), .B1(new_n637), .B2(new_n203), .ZN(new_n638));
  NAND2_X1  g452(.A1(new_n636), .A2(new_n638), .ZN(new_n639));
  INV_X1    g453(.A(new_n621), .ZN(new_n640));
  AOI21_X1  g454(.A(new_n635), .B1(new_n639), .B2(new_n640), .ZN(new_n641));
  OAI211_X1 g455(.A(new_n602), .B(new_n603), .C1(new_n634), .C2(new_n641), .ZN(new_n642));
  NAND2_X1  g456(.A1(new_n642), .A2(KEYINPUT90), .ZN(new_n643));
  NAND2_X1  g457(.A1(new_n639), .A2(new_n640), .ZN(new_n644));
  NAND2_X1  g458(.A1(new_n644), .A2(new_n606), .ZN(new_n645));
  NAND2_X1  g459(.A1(new_n627), .A2(new_n633), .ZN(new_n646));
  NAND3_X1  g460(.A1(new_n646), .A2(new_n640), .A3(new_n635), .ZN(new_n647));
  NAND2_X1  g461(.A1(new_n645), .A2(new_n647), .ZN(new_n648));
  INV_X1    g462(.A(KEYINPUT90), .ZN(new_n649));
  NAND4_X1  g463(.A1(new_n648), .A2(new_n649), .A3(new_n602), .A4(new_n603), .ZN(new_n650));
  OAI21_X1  g464(.A(new_n603), .B1(new_n634), .B2(new_n641), .ZN(new_n651));
  NAND2_X1  g465(.A1(new_n651), .A2(KEYINPUT20), .ZN(new_n652));
  NAND3_X1  g466(.A1(new_n643), .A2(new_n650), .A3(new_n652), .ZN(new_n653));
  AOI21_X1  g467(.A(new_n635), .B1(new_n646), .B2(new_n640), .ZN(new_n654));
  INV_X1    g468(.A(KEYINPUT91), .ZN(new_n655));
  NOR3_X1   g469(.A1(new_n654), .A2(new_n634), .A3(new_n655), .ZN(new_n656));
  NAND2_X1  g470(.A1(new_n646), .A2(new_n640), .ZN(new_n657));
  NAND3_X1  g471(.A1(new_n657), .A2(new_n655), .A3(new_n606), .ZN(new_n658));
  NAND2_X1  g472(.A1(new_n658), .A2(new_n301), .ZN(new_n659));
  OAI21_X1  g473(.A(G475), .B1(new_n656), .B2(new_n659), .ZN(new_n660));
  NAND2_X1  g474(.A1(new_n653), .A2(new_n660), .ZN(new_n661));
  NOR3_X1   g475(.A1(new_n519), .A2(new_n601), .A3(new_n661), .ZN(new_n662));
  NAND4_X1  g476(.A1(new_n313), .A2(new_n393), .A3(new_n453), .A4(new_n662), .ZN(new_n663));
  XNOR2_X1  g477(.A(new_n663), .B(G101), .ZN(G3));
  INV_X1    g478(.A(new_n582), .ZN(new_n665));
  XNOR2_X1  g479(.A(KEYINPUT100), .B(G478), .ZN(new_n666));
  NOR2_X1   g480(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  NAND2_X1  g481(.A1(new_n579), .A2(new_n581), .ZN(new_n668));
  INV_X1    g482(.A(KEYINPUT33), .ZN(new_n669));
  NAND2_X1  g483(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  INV_X1    g484(.A(new_n558), .ZN(new_n671));
  INV_X1    g485(.A(KEYINPUT99), .ZN(new_n672));
  NAND2_X1  g486(.A1(new_n578), .A2(new_n672), .ZN(new_n673));
  XNOR2_X1  g487(.A(new_n671), .B(new_n673), .ZN(new_n674));
  OAI21_X1  g488(.A(new_n670), .B1(new_n674), .B2(new_n669), .ZN(new_n675));
  NOR2_X1   g489(.A1(new_n587), .A2(G902), .ZN(new_n676));
  AOI21_X1  g490(.A(new_n667), .B1(new_n675), .B2(new_n676), .ZN(new_n677));
  AOI21_X1  g491(.A(new_n677), .B1(new_n653), .B2(new_n660), .ZN(new_n678));
  INV_X1    g492(.A(new_n678), .ZN(new_n679));
  NOR3_X1   g493(.A1(new_n679), .A2(new_n519), .A3(new_n600), .ZN(new_n680));
  NAND2_X1  g494(.A1(new_n286), .A2(new_n301), .ZN(new_n681));
  AND2_X1   g495(.A1(new_n681), .A2(KEYINPUT98), .ZN(new_n682));
  OAI21_X1  g496(.A(G472), .B1(new_n681), .B2(KEYINPUT98), .ZN(new_n683));
  NOR2_X1   g497(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  NAND2_X1  g498(.A1(new_n278), .A2(new_n288), .ZN(new_n685));
  INV_X1    g499(.A(new_n453), .ZN(new_n686));
  NOR3_X1   g500(.A1(new_n684), .A2(new_n685), .A3(new_n686), .ZN(new_n687));
  NAND3_X1  g501(.A1(new_n680), .A2(new_n687), .A3(new_n393), .ZN(new_n688));
  XOR2_X1   g502(.A(KEYINPUT34), .B(G104), .Z(new_n689));
  XNOR2_X1  g503(.A(new_n688), .B(new_n689), .ZN(G6));
  XOR2_X1   g504(.A(new_n600), .B(KEYINPUT101), .Z(new_n691));
  OAI211_X1 g505(.A(new_n454), .B(new_n691), .C1(new_n517), .C2(new_n518), .ZN(new_n692));
  NAND2_X1  g506(.A1(new_n652), .A2(new_n642), .ZN(new_n693));
  NAND3_X1  g507(.A1(new_n592), .A2(new_n660), .A3(new_n693), .ZN(new_n694));
  NOR2_X1   g508(.A1(new_n692), .A2(new_n694), .ZN(new_n695));
  NAND3_X1  g509(.A1(new_n687), .A2(new_n393), .A3(new_n695), .ZN(new_n696));
  XOR2_X1   g510(.A(KEYINPUT35), .B(G107), .Z(new_n697));
  XNOR2_X1  g511(.A(new_n696), .B(new_n697), .ZN(G9));
  INV_X1    g512(.A(new_n452), .ZN(new_n699));
  AOI21_X1  g513(.A(KEYINPUT25), .B1(new_n448), .B2(KEYINPUT73), .ZN(new_n700));
  NOR3_X1   g514(.A1(new_n699), .A2(new_n700), .A3(new_n395), .ZN(new_n701));
  NOR2_X1   g515(.A1(new_n433), .A2(KEYINPUT36), .ZN(new_n702));
  XNOR2_X1  g516(.A(new_n702), .B(new_n421), .ZN(new_n703));
  NAND3_X1  g517(.A1(new_n703), .A2(new_n301), .A3(new_n395), .ZN(new_n704));
  INV_X1    g518(.A(new_n704), .ZN(new_n705));
  OAI21_X1  g519(.A(KEYINPUT102), .B1(new_n701), .B2(new_n705), .ZN(new_n706));
  NAND2_X1  g520(.A1(new_n451), .A2(new_n452), .ZN(new_n707));
  INV_X1    g521(.A(KEYINPUT102), .ZN(new_n708));
  NAND3_X1  g522(.A1(new_n707), .A2(new_n708), .A3(new_n704), .ZN(new_n709));
  NAND2_X1  g523(.A1(new_n706), .A2(new_n709), .ZN(new_n710));
  INV_X1    g524(.A(new_n710), .ZN(new_n711));
  NOR3_X1   g525(.A1(new_n711), .A2(new_n684), .A3(new_n685), .ZN(new_n712));
  NAND3_X1  g526(.A1(new_n712), .A2(new_n393), .A3(new_n662), .ZN(new_n713));
  XOR2_X1   g527(.A(KEYINPUT37), .B(G110), .Z(new_n714));
  XNOR2_X1  g528(.A(new_n713), .B(new_n714), .ZN(G12));
  INV_X1    g529(.A(new_n454), .ZN(new_n716));
  NAND2_X1  g530(.A1(new_n501), .A2(new_n515), .ZN(new_n717));
  INV_X1    g531(.A(new_n516), .ZN(new_n718));
  NAND2_X1  g532(.A1(new_n717), .A2(new_n718), .ZN(new_n719));
  NAND3_X1  g533(.A1(new_n501), .A2(new_n515), .A3(new_n516), .ZN(new_n720));
  AOI21_X1  g534(.A(new_n716), .B1(new_n719), .B2(new_n720), .ZN(new_n721));
  INV_X1    g535(.A(G900), .ZN(new_n722));
  NAND2_X1  g536(.A1(new_n598), .A2(new_n722), .ZN(new_n723));
  NAND2_X1  g537(.A1(new_n723), .A2(new_n595), .ZN(new_n724));
  AND4_X1   g538(.A1(new_n660), .A2(new_n592), .A3(new_n693), .A4(new_n724), .ZN(new_n725));
  AND3_X1   g539(.A1(new_n721), .A2(new_n710), .A3(new_n725), .ZN(new_n726));
  NAND3_X1  g540(.A1(new_n313), .A2(new_n726), .A3(new_n393), .ZN(new_n727));
  XNOR2_X1  g541(.A(new_n727), .B(G128), .ZN(G30));
  XNOR2_X1  g542(.A(new_n724), .B(KEYINPUT39), .ZN(new_n729));
  NAND2_X1  g543(.A1(new_n393), .A2(new_n729), .ZN(new_n730));
  OR2_X1    g544(.A1(new_n730), .A2(KEYINPUT40), .ZN(new_n731));
  NAND2_X1  g545(.A1(new_n730), .A2(KEYINPUT40), .ZN(new_n732));
  NOR2_X1   g546(.A1(new_n517), .A2(new_n518), .ZN(new_n733));
  XNOR2_X1  g547(.A(KEYINPUT103), .B(KEYINPUT38), .ZN(new_n734));
  XNOR2_X1  g548(.A(new_n733), .B(new_n734), .ZN(new_n735));
  NOR2_X1   g549(.A1(new_n263), .A2(new_n280), .ZN(new_n736));
  OAI21_X1  g550(.A(new_n301), .B1(new_n254), .B2(new_n273), .ZN(new_n737));
  OAI21_X1  g551(.A(G472), .B1(new_n736), .B2(new_n737), .ZN(new_n738));
  AND3_X1   g552(.A1(new_n296), .A2(new_n310), .A3(new_n738), .ZN(new_n739));
  NAND2_X1  g553(.A1(new_n293), .A2(new_n739), .ZN(new_n740));
  NAND2_X1  g554(.A1(new_n661), .A2(new_n592), .ZN(new_n741));
  NOR3_X1   g555(.A1(new_n741), .A2(new_n716), .A3(new_n710), .ZN(new_n742));
  AND3_X1   g556(.A1(new_n735), .A2(new_n740), .A3(new_n742), .ZN(new_n743));
  NAND3_X1  g557(.A1(new_n731), .A2(new_n732), .A3(new_n743), .ZN(new_n744));
  XNOR2_X1  g558(.A(new_n744), .B(G143), .ZN(G45));
  AOI21_X1  g559(.A(new_n311), .B1(new_n291), .B2(new_n292), .ZN(new_n746));
  NOR2_X1   g560(.A1(new_n746), .A2(new_n711), .ZN(new_n747));
  NAND2_X1  g561(.A1(new_n678), .A2(new_n724), .ZN(new_n748));
  OAI21_X1  g562(.A(KEYINPUT104), .B1(new_n748), .B2(new_n519), .ZN(new_n749));
  INV_X1    g563(.A(KEYINPUT104), .ZN(new_n750));
  NAND4_X1  g564(.A1(new_n721), .A2(new_n750), .A3(new_n678), .A4(new_n724), .ZN(new_n751));
  NAND4_X1  g565(.A1(new_n747), .A2(new_n393), .A3(new_n749), .A4(new_n751), .ZN(new_n752));
  XNOR2_X1  g566(.A(new_n752), .B(G146), .ZN(G48));
  AND3_X1   g567(.A1(new_n377), .A2(new_n378), .A3(new_n301), .ZN(new_n754));
  AOI21_X1  g568(.A(new_n378), .B1(new_n377), .B2(new_n301), .ZN(new_n755));
  NOR3_X1   g569(.A1(new_n754), .A2(new_n755), .A3(new_n389), .ZN(new_n756));
  NAND4_X1  g570(.A1(new_n313), .A2(new_n680), .A3(new_n453), .A4(new_n756), .ZN(new_n757));
  XNOR2_X1  g571(.A(KEYINPUT41), .B(G113), .ZN(new_n758));
  XNOR2_X1  g572(.A(new_n757), .B(new_n758), .ZN(G15));
  NAND4_X1  g573(.A1(new_n313), .A2(new_n453), .A3(new_n695), .A4(new_n756), .ZN(new_n760));
  XNOR2_X1  g574(.A(new_n760), .B(G116), .ZN(G18));
  NAND4_X1  g575(.A1(new_n313), .A2(new_n662), .A3(new_n710), .A4(new_n756), .ZN(new_n762));
  XNOR2_X1  g576(.A(KEYINPUT105), .B(G119), .ZN(new_n763));
  XNOR2_X1  g577(.A(new_n762), .B(new_n763), .ZN(G21));
  INV_X1    g578(.A(KEYINPUT106), .ZN(new_n765));
  AOI21_X1  g579(.A(new_n254), .B1(new_n274), .B2(new_n282), .ZN(new_n766));
  OAI21_X1  g580(.A(new_n187), .B1(new_n266), .B2(new_n766), .ZN(new_n767));
  AND4_X1   g581(.A1(new_n264), .A2(new_n240), .A3(new_n254), .A4(new_n256), .ZN(new_n768));
  AOI21_X1  g582(.A(new_n264), .B1(new_n263), .B2(new_n254), .ZN(new_n769));
  NOR2_X1   g583(.A1(new_n768), .A2(new_n769), .ZN(new_n770));
  AOI21_X1  g584(.A(G902), .B1(new_n770), .B2(new_n285), .ZN(new_n771));
  INV_X1    g585(.A(G472), .ZN(new_n772));
  OAI211_X1 g586(.A(new_n453), .B(new_n767), .C1(new_n771), .C2(new_n772), .ZN(new_n773));
  INV_X1    g587(.A(new_n691), .ZN(new_n774));
  NOR2_X1   g588(.A1(new_n773), .A2(new_n774), .ZN(new_n775));
  NAND2_X1  g589(.A1(new_n756), .A2(new_n775), .ZN(new_n776));
  NAND2_X1  g590(.A1(new_n719), .A2(new_n720), .ZN(new_n777));
  AOI21_X1  g591(.A(new_n590), .B1(new_n586), .B2(new_n588), .ZN(new_n778));
  AOI21_X1  g592(.A(new_n778), .B1(new_n653), .B2(new_n660), .ZN(new_n779));
  NAND3_X1  g593(.A1(new_n777), .A2(new_n779), .A3(new_n454), .ZN(new_n780));
  OAI21_X1  g594(.A(new_n765), .B1(new_n776), .B2(new_n780), .ZN(new_n781));
  NOR2_X1   g595(.A1(new_n741), .A2(new_n519), .ZN(new_n782));
  NAND2_X1  g596(.A1(new_n377), .A2(new_n301), .ZN(new_n783));
  NAND2_X1  g597(.A1(new_n783), .A2(G469), .ZN(new_n784));
  NAND3_X1  g598(.A1(new_n784), .A2(new_n390), .A3(new_n379), .ZN(new_n785));
  NAND2_X1  g599(.A1(new_n681), .A2(G472), .ZN(new_n786));
  NAND4_X1  g600(.A1(new_n786), .A2(new_n453), .A3(new_n691), .A4(new_n767), .ZN(new_n787));
  NOR2_X1   g601(.A1(new_n785), .A2(new_n787), .ZN(new_n788));
  NAND3_X1  g602(.A1(new_n782), .A2(new_n788), .A3(KEYINPUT106), .ZN(new_n789));
  NAND2_X1  g603(.A1(new_n781), .A2(new_n789), .ZN(new_n790));
  XOR2_X1   g604(.A(KEYINPUT107), .B(G122), .Z(new_n791));
  XNOR2_X1  g605(.A(new_n790), .B(new_n791), .ZN(G24));
  NAND2_X1  g606(.A1(new_n756), .A2(new_n721), .ZN(new_n793));
  OR2_X1    g607(.A1(new_n266), .A2(new_n766), .ZN(new_n794));
  AOI22_X1  g608(.A1(G472), .A2(new_n681), .B1(new_n794), .B2(new_n187), .ZN(new_n795));
  NAND4_X1  g609(.A1(new_n678), .A2(new_n710), .A3(new_n724), .A4(new_n795), .ZN(new_n796));
  NOR2_X1   g610(.A1(new_n793), .A2(new_n796), .ZN(new_n797));
  XNOR2_X1  g611(.A(new_n797), .B(new_n406), .ZN(G27));
  AOI21_X1  g612(.A(new_n389), .B1(new_n379), .B2(new_n384), .ZN(new_n799));
  NAND4_X1  g613(.A1(new_n733), .A2(new_n799), .A3(new_n453), .A4(new_n454), .ZN(new_n800));
  NAND2_X1  g614(.A1(new_n277), .A2(new_n279), .ZN(new_n801));
  NAND3_X1  g615(.A1(new_n309), .A2(new_n801), .A3(new_n294), .ZN(new_n802));
  NAND4_X1  g616(.A1(new_n678), .A2(KEYINPUT42), .A3(new_n724), .A4(new_n802), .ZN(new_n803));
  NOR2_X1   g617(.A1(new_n800), .A2(new_n803), .ZN(new_n804));
  INV_X1    g618(.A(new_n804), .ZN(new_n805));
  NOR3_X1   g619(.A1(new_n746), .A2(new_n800), .A3(new_n748), .ZN(new_n806));
  XNOR2_X1  g620(.A(KEYINPUT108), .B(KEYINPUT42), .ZN(new_n807));
  OAI21_X1  g621(.A(new_n805), .B1(new_n806), .B2(new_n807), .ZN(new_n808));
  NAND2_X1  g622(.A1(new_n808), .A2(KEYINPUT109), .ZN(new_n809));
  AND4_X1   g623(.A1(new_n453), .A2(new_n733), .A3(new_n799), .A4(new_n454), .ZN(new_n810));
  INV_X1    g624(.A(new_n748), .ZN(new_n811));
  NAND3_X1  g625(.A1(new_n313), .A2(new_n810), .A3(new_n811), .ZN(new_n812));
  INV_X1    g626(.A(new_n807), .ZN(new_n813));
  NAND2_X1  g627(.A1(new_n812), .A2(new_n813), .ZN(new_n814));
  INV_X1    g628(.A(KEYINPUT109), .ZN(new_n815));
  NAND3_X1  g629(.A1(new_n814), .A2(new_n815), .A3(new_n805), .ZN(new_n816));
  NAND2_X1  g630(.A1(new_n809), .A2(new_n816), .ZN(new_n817));
  XNOR2_X1  g631(.A(new_n817), .B(new_n217), .ZN(G33));
  NAND3_X1  g632(.A1(new_n313), .A2(new_n810), .A3(new_n725), .ZN(new_n819));
  XNOR2_X1  g633(.A(new_n819), .B(G134), .ZN(G36));
  NAND3_X1  g634(.A1(new_n719), .A2(new_n454), .A3(new_n720), .ZN(new_n821));
  OR2_X1    g635(.A1(new_n383), .A2(KEYINPUT45), .ZN(new_n822));
  NAND2_X1  g636(.A1(new_n383), .A2(KEYINPUT45), .ZN(new_n823));
  NAND3_X1  g637(.A1(new_n822), .A2(G469), .A3(new_n823), .ZN(new_n824));
  NAND2_X1  g638(.A1(G469), .A2(G902), .ZN(new_n825));
  AOI21_X1  g639(.A(KEYINPUT46), .B1(new_n824), .B2(new_n825), .ZN(new_n826));
  NOR2_X1   g640(.A1(new_n826), .A2(new_n754), .ZN(new_n827));
  NAND3_X1  g641(.A1(new_n824), .A2(KEYINPUT46), .A3(new_n825), .ZN(new_n828));
  NAND2_X1  g642(.A1(new_n827), .A2(new_n828), .ZN(new_n829));
  NAND3_X1  g643(.A1(new_n829), .A2(new_n390), .A3(new_n729), .ZN(new_n830));
  INV_X1    g644(.A(new_n661), .ZN(new_n831));
  INV_X1    g645(.A(KEYINPUT110), .ZN(new_n832));
  AOI21_X1  g646(.A(KEYINPUT43), .B1(new_n831), .B2(new_n832), .ZN(new_n833));
  INV_X1    g647(.A(new_n677), .ZN(new_n834));
  NAND2_X1  g648(.A1(new_n831), .A2(new_n834), .ZN(new_n835));
  NAND2_X1  g649(.A1(new_n833), .A2(new_n835), .ZN(new_n836));
  OAI211_X1 g650(.A(new_n831), .B(new_n834), .C1(new_n832), .C2(KEYINPUT43), .ZN(new_n837));
  NAND2_X1  g651(.A1(new_n836), .A2(new_n837), .ZN(new_n838));
  OAI211_X1 g652(.A(new_n838), .B(new_n710), .C1(new_n685), .C2(new_n684), .ZN(new_n839));
  INV_X1    g653(.A(KEYINPUT44), .ZN(new_n840));
  AOI211_X1 g654(.A(new_n821), .B(new_n830), .C1(new_n839), .C2(new_n840), .ZN(new_n841));
  OAI21_X1  g655(.A(new_n841), .B1(new_n840), .B2(new_n839), .ZN(new_n842));
  XNOR2_X1  g656(.A(new_n842), .B(G137), .ZN(G39));
  INV_X1    g657(.A(new_n821), .ZN(new_n844));
  NAND4_X1  g658(.A1(new_n746), .A2(new_n811), .A3(new_n686), .A4(new_n844), .ZN(new_n845));
  NOR2_X1   g659(.A1(new_n845), .A2(KEYINPUT112), .ZN(new_n846));
  AOI21_X1  g660(.A(new_n389), .B1(new_n827), .B2(new_n828), .ZN(new_n847));
  XNOR2_X1  g661(.A(KEYINPUT111), .B(KEYINPUT47), .ZN(new_n848));
  NOR2_X1   g662(.A1(new_n847), .A2(new_n848), .ZN(new_n849));
  INV_X1    g663(.A(new_n849), .ZN(new_n850));
  NAND3_X1  g664(.A1(new_n829), .A2(new_n390), .A3(new_n848), .ZN(new_n851));
  AOI21_X1  g665(.A(new_n846), .B1(new_n850), .B2(new_n851), .ZN(new_n852));
  NAND2_X1  g666(.A1(new_n845), .A2(KEYINPUT112), .ZN(new_n853));
  NAND2_X1  g667(.A1(new_n852), .A2(new_n853), .ZN(new_n854));
  XNOR2_X1  g668(.A(new_n854), .B(G140), .ZN(G42));
  AND2_X1   g669(.A1(new_n710), .A2(new_n795), .ZN(new_n856));
  NOR2_X1   g670(.A1(new_n785), .A2(new_n821), .ZN(new_n857));
  AOI21_X1  g671(.A(KEYINPUT117), .B1(new_n838), .B2(new_n596), .ZN(new_n858));
  INV_X1    g672(.A(KEYINPUT117), .ZN(new_n859));
  AOI211_X1 g673(.A(new_n859), .B(new_n595), .C1(new_n836), .C2(new_n837), .ZN(new_n860));
  OAI211_X1 g674(.A(new_n856), .B(new_n857), .C1(new_n858), .C2(new_n860), .ZN(new_n861));
  INV_X1    g675(.A(new_n740), .ZN(new_n862));
  NAND4_X1  g676(.A1(new_n862), .A2(new_n453), .A3(new_n596), .A4(new_n857), .ZN(new_n863));
  INV_X1    g677(.A(KEYINPUT120), .ZN(new_n864));
  XNOR2_X1  g678(.A(new_n863), .B(new_n864), .ZN(new_n865));
  NOR2_X1   g679(.A1(new_n661), .A2(new_n834), .ZN(new_n866));
  INV_X1    g680(.A(new_n866), .ZN(new_n867));
  OAI21_X1  g681(.A(new_n861), .B1(new_n865), .B2(new_n867), .ZN(new_n868));
  INV_X1    g682(.A(new_n773), .ZN(new_n869));
  NOR3_X1   g683(.A1(new_n735), .A2(new_n454), .A3(new_n785), .ZN(new_n870));
  OAI211_X1 g684(.A(new_n869), .B(new_n870), .C1(new_n858), .C2(new_n860), .ZN(new_n871));
  INV_X1    g685(.A(KEYINPUT50), .ZN(new_n872));
  OR2_X1    g686(.A1(new_n871), .A2(new_n872), .ZN(new_n873));
  NAND2_X1  g687(.A1(new_n871), .A2(new_n872), .ZN(new_n874));
  AOI21_X1  g688(.A(new_n868), .B1(new_n873), .B2(new_n874), .ZN(new_n875));
  INV_X1    g689(.A(KEYINPUT51), .ZN(new_n876));
  INV_X1    g690(.A(new_n858), .ZN(new_n877));
  INV_X1    g691(.A(new_n860), .ZN(new_n878));
  AOI211_X1 g692(.A(new_n773), .B(new_n821), .C1(new_n877), .C2(new_n878), .ZN(new_n879));
  NOR2_X1   g693(.A1(new_n754), .A2(new_n755), .ZN(new_n880));
  XNOR2_X1  g694(.A(new_n880), .B(KEYINPUT114), .ZN(new_n881));
  NAND2_X1  g695(.A1(new_n881), .A2(new_n389), .ZN(new_n882));
  NAND3_X1  g696(.A1(new_n850), .A2(new_n851), .A3(new_n882), .ZN(new_n883));
  AOI21_X1  g697(.A(new_n876), .B1(new_n879), .B2(new_n883), .ZN(new_n884));
  NAND2_X1  g698(.A1(new_n875), .A2(new_n884), .ZN(new_n885));
  INV_X1    g699(.A(new_n793), .ZN(new_n886));
  OAI211_X1 g700(.A(new_n869), .B(new_n886), .C1(new_n858), .C2(new_n860), .ZN(new_n887));
  OAI211_X1 g701(.A(new_n887), .B(new_n593), .C1(new_n865), .C2(new_n679), .ZN(new_n888));
  NAND2_X1  g702(.A1(new_n877), .A2(new_n878), .ZN(new_n889));
  AND2_X1   g703(.A1(new_n802), .A2(new_n453), .ZN(new_n890));
  NAND3_X1  g704(.A1(new_n889), .A2(new_n857), .A3(new_n890), .ZN(new_n891));
  NAND2_X1  g705(.A1(new_n891), .A2(KEYINPUT48), .ZN(new_n892));
  INV_X1    g706(.A(KEYINPUT48), .ZN(new_n893));
  NAND4_X1  g707(.A1(new_n889), .A2(new_n893), .A3(new_n857), .A4(new_n890), .ZN(new_n894));
  AOI21_X1  g708(.A(new_n888), .B1(new_n892), .B2(new_n894), .ZN(new_n895));
  XOR2_X1   g709(.A(new_n882), .B(KEYINPUT119), .Z(new_n896));
  AND3_X1   g710(.A1(new_n850), .A2(KEYINPUT118), .A3(new_n851), .ZN(new_n897));
  AOI21_X1  g711(.A(KEYINPUT118), .B1(new_n850), .B2(new_n851), .ZN(new_n898));
  OAI21_X1  g712(.A(new_n896), .B1(new_n897), .B2(new_n898), .ZN(new_n899));
  NAND2_X1  g713(.A1(new_n899), .A2(new_n879), .ZN(new_n900));
  AND2_X1   g714(.A1(new_n875), .A2(new_n900), .ZN(new_n901));
  OAI211_X1 g715(.A(new_n885), .B(new_n895), .C1(new_n901), .C2(KEYINPUT51), .ZN(new_n902));
  AND3_X1   g716(.A1(new_n790), .A2(new_n757), .A3(new_n760), .ZN(new_n903));
  NAND3_X1  g717(.A1(new_n653), .A2(new_n660), .A3(new_n592), .ZN(new_n904));
  NOR2_X1   g718(.A1(new_n692), .A2(new_n904), .ZN(new_n905));
  NAND3_X1  g719(.A1(new_n687), .A2(new_n393), .A3(new_n905), .ZN(new_n906));
  AND3_X1   g720(.A1(new_n762), .A2(new_n713), .A3(new_n906), .ZN(new_n907));
  NOR3_X1   g721(.A1(new_n679), .A2(new_n519), .A3(new_n774), .ZN(new_n908));
  NAND3_X1  g722(.A1(new_n908), .A2(new_n687), .A3(new_n393), .ZN(new_n909));
  INV_X1    g723(.A(KEYINPUT115), .ZN(new_n910));
  NAND3_X1  g724(.A1(new_n663), .A2(new_n909), .A3(new_n910), .ZN(new_n911));
  INV_X1    g725(.A(new_n911), .ZN(new_n912));
  AOI21_X1  g726(.A(new_n910), .B1(new_n663), .B2(new_n909), .ZN(new_n913));
  OAI211_X1 g727(.A(new_n903), .B(new_n907), .C1(new_n912), .C2(new_n913), .ZN(new_n914));
  NAND4_X1  g728(.A1(new_n660), .A2(new_n693), .A3(new_n778), .A4(new_n724), .ZN(new_n915));
  NOR2_X1   g729(.A1(new_n821), .A2(new_n915), .ZN(new_n916));
  NAND4_X1  g730(.A1(new_n313), .A2(new_n393), .A3(new_n710), .A4(new_n916), .ZN(new_n917));
  NAND4_X1  g731(.A1(new_n811), .A2(new_n799), .A3(new_n856), .A4(new_n844), .ZN(new_n918));
  AND3_X1   g732(.A1(new_n917), .A2(new_n819), .A3(new_n918), .ZN(new_n919));
  NAND3_X1  g733(.A1(new_n809), .A2(new_n816), .A3(new_n919), .ZN(new_n920));
  NOR2_X1   g734(.A1(new_n914), .A2(new_n920), .ZN(new_n921));
  INV_X1    g735(.A(KEYINPUT53), .ZN(new_n922));
  INV_X1    g736(.A(new_n752), .ZN(new_n923));
  INV_X1    g737(.A(new_n797), .ZN(new_n924));
  AND4_X1   g738(.A1(new_n707), .A2(new_n799), .A3(new_n704), .A4(new_n724), .ZN(new_n925));
  NAND3_X1  g739(.A1(new_n740), .A2(new_n782), .A3(new_n925), .ZN(new_n926));
  NAND3_X1  g740(.A1(new_n727), .A2(new_n924), .A3(new_n926), .ZN(new_n927));
  OAI21_X1  g741(.A(KEYINPUT52), .B1(new_n923), .B2(new_n927), .ZN(new_n928));
  NAND3_X1  g742(.A1(new_n721), .A2(new_n725), .A3(new_n710), .ZN(new_n929));
  NOR2_X1   g743(.A1(new_n746), .A2(new_n929), .ZN(new_n930));
  AOI21_X1  g744(.A(new_n797), .B1(new_n930), .B2(new_n393), .ZN(new_n931));
  INV_X1    g745(.A(KEYINPUT52), .ZN(new_n932));
  NAND4_X1  g746(.A1(new_n931), .A2(new_n752), .A3(new_n932), .A4(new_n926), .ZN(new_n933));
  AND3_X1   g747(.A1(new_n928), .A2(KEYINPUT116), .A3(new_n933), .ZN(new_n934));
  AOI21_X1  g748(.A(KEYINPUT116), .B1(new_n928), .B2(new_n933), .ZN(new_n935));
  OAI211_X1 g749(.A(new_n921), .B(new_n922), .C1(new_n934), .C2(new_n935), .ZN(new_n936));
  AOI21_X1  g750(.A(new_n815), .B1(new_n814), .B2(new_n805), .ZN(new_n937));
  AOI211_X1 g751(.A(KEYINPUT109), .B(new_n804), .C1(new_n812), .C2(new_n813), .ZN(new_n938));
  NOR2_X1   g752(.A1(new_n937), .A2(new_n938), .ZN(new_n939));
  NAND2_X1  g753(.A1(new_n663), .A2(new_n909), .ZN(new_n940));
  NAND2_X1  g754(.A1(new_n940), .A2(KEYINPUT115), .ZN(new_n941));
  NAND2_X1  g755(.A1(new_n941), .A2(new_n911), .ZN(new_n942));
  NAND3_X1  g756(.A1(new_n790), .A2(new_n757), .A3(new_n760), .ZN(new_n943));
  NAND3_X1  g757(.A1(new_n762), .A2(new_n713), .A3(new_n906), .ZN(new_n944));
  NOR2_X1   g758(.A1(new_n943), .A2(new_n944), .ZN(new_n945));
  NAND4_X1  g759(.A1(new_n939), .A2(new_n942), .A3(new_n945), .A4(new_n919), .ZN(new_n946));
  NAND2_X1  g760(.A1(new_n928), .A2(new_n933), .ZN(new_n947));
  OAI21_X1  g761(.A(KEYINPUT53), .B1(new_n946), .B2(new_n947), .ZN(new_n948));
  NAND3_X1  g762(.A1(new_n936), .A2(new_n948), .A3(KEYINPUT54), .ZN(new_n949));
  OAI21_X1  g763(.A(new_n922), .B1(new_n946), .B2(new_n947), .ZN(new_n950));
  INV_X1    g764(.A(KEYINPUT54), .ZN(new_n951));
  AOI21_X1  g765(.A(new_n922), .B1(new_n814), .B2(new_n805), .ZN(new_n952));
  NAND2_X1  g766(.A1(new_n952), .A2(new_n919), .ZN(new_n953));
  NOR2_X1   g767(.A1(new_n914), .A2(new_n953), .ZN(new_n954));
  OAI21_X1  g768(.A(new_n954), .B1(new_n934), .B2(new_n935), .ZN(new_n955));
  NAND3_X1  g769(.A1(new_n950), .A2(new_n951), .A3(new_n955), .ZN(new_n956));
  NAND2_X1  g770(.A1(new_n949), .A2(new_n956), .ZN(new_n957));
  OAI22_X1  g771(.A1(new_n902), .A2(new_n957), .B1(G952), .B2(G953), .ZN(new_n958));
  NAND3_X1  g772(.A1(new_n453), .A2(new_n390), .A3(new_n454), .ZN(new_n959));
  XNOR2_X1  g773(.A(new_n959), .B(KEYINPUT113), .ZN(new_n960));
  NOR3_X1   g774(.A1(new_n735), .A2(new_n835), .A3(new_n960), .ZN(new_n961));
  INV_X1    g775(.A(KEYINPUT49), .ZN(new_n962));
  AOI21_X1  g776(.A(new_n740), .B1(new_n881), .B2(new_n962), .ZN(new_n963));
  OAI211_X1 g777(.A(new_n961), .B(new_n963), .C1(new_n962), .C2(new_n881), .ZN(new_n964));
  NAND2_X1  g778(.A1(new_n958), .A2(new_n964), .ZN(G75));
  NOR2_X1   g779(.A1(new_n423), .A2(G952), .ZN(new_n966));
  XOR2_X1   g780(.A(new_n966), .B(KEYINPUT122), .Z(new_n967));
  INV_X1    g781(.A(new_n967), .ZN(new_n968));
  INV_X1    g782(.A(KEYINPUT121), .ZN(new_n969));
  NOR2_X1   g783(.A1(new_n969), .A2(KEYINPUT56), .ZN(new_n970));
  NAND2_X1  g784(.A1(new_n950), .A2(new_n955), .ZN(new_n971));
  NAND2_X1  g785(.A1(new_n971), .A2(G902), .ZN(new_n972));
  INV_X1    g786(.A(G210), .ZN(new_n973));
  OAI21_X1  g787(.A(new_n970), .B1(new_n972), .B2(new_n973), .ZN(new_n974));
  OAI21_X1  g788(.A(new_n484), .B1(new_n500), .B2(new_n497), .ZN(new_n975));
  XNOR2_X1  g789(.A(new_n975), .B(new_n491), .ZN(new_n976));
  XNOR2_X1  g790(.A(new_n976), .B(KEYINPUT55), .ZN(new_n977));
  NAND2_X1  g791(.A1(new_n974), .A2(new_n977), .ZN(new_n978));
  INV_X1    g792(.A(new_n977), .ZN(new_n979));
  OAI211_X1 g793(.A(new_n979), .B(new_n970), .C1(new_n972), .C2(new_n973), .ZN(new_n980));
  AOI21_X1  g794(.A(new_n968), .B1(new_n978), .B2(new_n980), .ZN(G51));
  INV_X1    g795(.A(new_n947), .ZN(new_n982));
  AOI21_X1  g796(.A(KEYINPUT53), .B1(new_n921), .B2(new_n982), .ZN(new_n983));
  NAND4_X1  g797(.A1(new_n942), .A2(new_n945), .A3(new_n919), .A4(new_n952), .ZN(new_n984));
  INV_X1    g798(.A(KEYINPUT116), .ZN(new_n985));
  AND3_X1   g799(.A1(new_n727), .A2(new_n924), .A3(new_n926), .ZN(new_n986));
  AOI21_X1  g800(.A(new_n932), .B1(new_n986), .B2(new_n752), .ZN(new_n987));
  AND4_X1   g801(.A1(new_n932), .A2(new_n931), .A3(new_n752), .A4(new_n926), .ZN(new_n988));
  OAI21_X1  g802(.A(new_n985), .B1(new_n987), .B2(new_n988), .ZN(new_n989));
  NAND3_X1  g803(.A1(new_n928), .A2(KEYINPUT116), .A3(new_n933), .ZN(new_n990));
  AOI21_X1  g804(.A(new_n984), .B1(new_n989), .B2(new_n990), .ZN(new_n991));
  OAI21_X1  g805(.A(KEYINPUT54), .B1(new_n983), .B2(new_n991), .ZN(new_n992));
  NAND3_X1  g806(.A1(new_n992), .A2(new_n956), .A3(KEYINPUT123), .ZN(new_n993));
  INV_X1    g807(.A(KEYINPUT123), .ZN(new_n994));
  NAND3_X1  g808(.A1(new_n971), .A2(new_n994), .A3(KEYINPUT54), .ZN(new_n995));
  XOR2_X1   g809(.A(new_n825), .B(KEYINPUT57), .Z(new_n996));
  NAND3_X1  g810(.A1(new_n993), .A2(new_n995), .A3(new_n996), .ZN(new_n997));
  NAND2_X1  g811(.A1(new_n997), .A2(new_n377), .ZN(new_n998));
  OR2_X1    g812(.A1(new_n972), .A2(new_n824), .ZN(new_n999));
  AOI21_X1  g813(.A(new_n966), .B1(new_n998), .B2(new_n999), .ZN(G54));
  NAND2_X1  g814(.A1(KEYINPUT58), .A2(G475), .ZN(new_n1001));
  NOR2_X1   g815(.A1(new_n972), .A2(new_n1001), .ZN(new_n1002));
  NOR2_X1   g816(.A1(new_n1002), .A2(new_n648), .ZN(new_n1003));
  INV_X1    g817(.A(new_n648), .ZN(new_n1004));
  NOR3_X1   g818(.A1(new_n972), .A2(new_n1004), .A3(new_n1001), .ZN(new_n1005));
  NOR3_X1   g819(.A1(new_n1003), .A2(new_n966), .A3(new_n1005), .ZN(G60));
  NAND2_X1  g820(.A1(G478), .A2(G902), .ZN(new_n1007));
  XOR2_X1   g821(.A(new_n1007), .B(KEYINPUT59), .Z(new_n1008));
  INV_X1    g822(.A(new_n1008), .ZN(new_n1009));
  AND4_X1   g823(.A1(new_n675), .A2(new_n993), .A3(new_n995), .A4(new_n1009), .ZN(new_n1010));
  AOI21_X1  g824(.A(new_n1008), .B1(new_n949), .B2(new_n956), .ZN(new_n1011));
  OAI21_X1  g825(.A(new_n967), .B1(new_n1011), .B2(new_n675), .ZN(new_n1012));
  NOR2_X1   g826(.A1(new_n1010), .A2(new_n1012), .ZN(G63));
  NAND2_X1  g827(.A1(G217), .A2(G902), .ZN(new_n1014));
  XNOR2_X1  g828(.A(new_n1014), .B(KEYINPUT124), .ZN(new_n1015));
  XNOR2_X1  g829(.A(new_n1015), .B(KEYINPUT60), .ZN(new_n1016));
  INV_X1    g830(.A(new_n1016), .ZN(new_n1017));
  AOI21_X1  g831(.A(new_n1017), .B1(new_n950), .B2(new_n955), .ZN(new_n1018));
  NAND2_X1  g832(.A1(new_n1018), .A2(new_n703), .ZN(new_n1019));
  AOI21_X1  g833(.A(new_n441), .B1(KEYINPUT72), .B2(new_n442), .ZN(new_n1020));
  OAI211_X1 g834(.A(new_n1019), .B(new_n967), .C1(new_n1020), .C2(new_n1018), .ZN(new_n1021));
  INV_X1    g835(.A(KEYINPUT61), .ZN(new_n1022));
  NAND2_X1  g836(.A1(new_n1021), .A2(new_n1022), .ZN(new_n1023));
  OR2_X1    g837(.A1(new_n1018), .A2(new_n1020), .ZN(new_n1024));
  NAND4_X1  g838(.A1(new_n1024), .A2(KEYINPUT61), .A3(new_n967), .A4(new_n1019), .ZN(new_n1025));
  NAND2_X1  g839(.A1(new_n1023), .A2(new_n1025), .ZN(G66));
  INV_X1    g840(.A(new_n599), .ZN(new_n1027));
  AOI21_X1  g841(.A(new_n423), .B1(new_n1027), .B2(G224), .ZN(new_n1028));
  AOI21_X1  g842(.A(new_n1028), .B1(new_n914), .B2(new_n423), .ZN(new_n1029));
  OAI21_X1  g843(.A(new_n975), .B1(G898), .B2(new_n423), .ZN(new_n1030));
  XNOR2_X1  g844(.A(new_n1030), .B(KEYINPUT125), .ZN(new_n1031));
  XNOR2_X1  g845(.A(new_n1029), .B(new_n1031), .ZN(G69));
  AND2_X1   g846(.A1(new_n931), .A2(new_n752), .ZN(new_n1033));
  NAND2_X1  g847(.A1(new_n1033), .A2(new_n744), .ZN(new_n1034));
  INV_X1    g848(.A(KEYINPUT62), .ZN(new_n1035));
  XNOR2_X1  g849(.A(new_n1034), .B(new_n1035), .ZN(new_n1036));
  NAND2_X1  g850(.A1(new_n679), .A2(new_n904), .ZN(new_n1037));
  AOI21_X1  g851(.A(new_n730), .B1(KEYINPUT126), .B2(new_n1037), .ZN(new_n1038));
  NOR3_X1   g852(.A1(new_n746), .A2(new_n686), .A3(new_n821), .ZN(new_n1039));
  OAI211_X1 g853(.A(new_n1038), .B(new_n1039), .C1(KEYINPUT126), .C2(new_n1037), .ZN(new_n1040));
  NAND4_X1  g854(.A1(new_n1036), .A2(new_n842), .A3(new_n854), .A4(new_n1040), .ZN(new_n1041));
  NAND2_X1  g855(.A1(new_n1041), .A2(new_n423), .ZN(new_n1042));
  XOR2_X1   g856(.A(new_n262), .B(new_n637), .Z(new_n1043));
  NAND2_X1  g857(.A1(new_n782), .A2(new_n890), .ZN(new_n1044));
  OAI211_X1 g858(.A(new_n1033), .B(new_n819), .C1(new_n830), .C2(new_n1044), .ZN(new_n1045));
  NOR2_X1   g859(.A1(new_n1045), .A2(new_n817), .ZN(new_n1046));
  NAND3_X1  g860(.A1(new_n1046), .A2(new_n842), .A3(new_n854), .ZN(new_n1047));
  OR2_X1    g861(.A1(new_n1047), .A2(G953), .ZN(new_n1048));
  AOI21_X1  g862(.A(new_n1043), .B1(G900), .B2(G953), .ZN(new_n1049));
  AOI22_X1  g863(.A1(new_n1042), .A2(new_n1043), .B1(new_n1048), .B2(new_n1049), .ZN(new_n1050));
  OAI21_X1  g864(.A(G953), .B1(new_n316), .B2(new_n722), .ZN(new_n1051));
  XNOR2_X1  g865(.A(new_n1050), .B(new_n1051), .ZN(G72));
  NAND2_X1  g866(.A1(G472), .A2(G902), .ZN(new_n1053));
  XOR2_X1   g867(.A(new_n1053), .B(KEYINPUT63), .Z(new_n1054));
  OAI21_X1  g868(.A(new_n1054), .B1(new_n1041), .B2(new_n914), .ZN(new_n1055));
  NAND2_X1  g869(.A1(new_n1055), .A2(new_n736), .ZN(new_n1056));
  OAI21_X1  g870(.A(new_n1054), .B1(new_n1047), .B2(new_n914), .ZN(new_n1057));
  NAND2_X1  g871(.A1(new_n263), .A2(new_n280), .ZN(new_n1058));
  INV_X1    g872(.A(new_n1058), .ZN(new_n1059));
  AOI21_X1  g873(.A(new_n966), .B1(new_n1057), .B2(new_n1059), .ZN(new_n1060));
  NAND2_X1  g874(.A1(new_n1056), .A2(new_n1060), .ZN(new_n1061));
  INV_X1    g875(.A(new_n1054), .ZN(new_n1062));
  NOR3_X1   g876(.A1(new_n1059), .A2(new_n736), .A3(new_n1062), .ZN(new_n1063));
  NAND3_X1  g877(.A1(new_n936), .A2(new_n948), .A3(new_n1063), .ZN(new_n1064));
  OR2_X1    g878(.A1(new_n1064), .A2(KEYINPUT127), .ZN(new_n1065));
  NAND2_X1  g879(.A1(new_n1064), .A2(KEYINPUT127), .ZN(new_n1066));
  AOI21_X1  g880(.A(new_n1061), .B1(new_n1065), .B2(new_n1066), .ZN(G57));
endmodule


