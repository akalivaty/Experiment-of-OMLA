//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 0 0 0 1 1 1 1 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 0 0 0 1 1 0 1 1 0 0 0 0 0 0 1 1 0 1 1 1 0 1 0 1 0 0 1 0 0 0 1 1 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:26:59 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n584, new_n585, new_n586, new_n587,
    new_n589, new_n590, new_n591, new_n592, new_n593, new_n594, new_n595,
    new_n597, new_n598, new_n599, new_n600, new_n601, new_n602, new_n603,
    new_n604, new_n605, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n622, new_n623, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n643, new_n645, new_n646, new_n647, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n656, new_n657, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n684, new_n685, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n865, new_n866, new_n868, new_n869, new_n870, new_n871,
    new_n872, new_n873, new_n874, new_n875, new_n876, new_n877, new_n878,
    new_n879, new_n880, new_n881, new_n882, new_n883, new_n884, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n903, new_n904, new_n905, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n929, new_n930, new_n931,
    new_n932, new_n933, new_n934, new_n935, new_n936, new_n937, new_n938,
    new_n939, new_n940;
  INV_X1    g000(.A(G475), .ZN(new_n187));
  INV_X1    g001(.A(G902), .ZN(new_n188));
  INV_X1    g002(.A(G125), .ZN(new_n189));
  NOR3_X1   g003(.A1(new_n189), .A2(KEYINPUT16), .A3(G140), .ZN(new_n190));
  XNOR2_X1  g004(.A(G125), .B(G140), .ZN(new_n191));
  AOI21_X1  g005(.A(new_n190), .B1(new_n191), .B2(KEYINPUT16), .ZN(new_n192));
  OAI21_X1  g006(.A(KEYINPUT71), .B1(new_n192), .B2(G146), .ZN(new_n193));
  INV_X1    g007(.A(new_n190), .ZN(new_n194));
  INV_X1    g008(.A(G140), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n195), .A2(G125), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n189), .A2(G140), .ZN(new_n197));
  NAND3_X1  g011(.A1(new_n196), .A2(new_n197), .A3(KEYINPUT16), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n194), .A2(new_n198), .ZN(new_n199));
  INV_X1    g013(.A(KEYINPUT71), .ZN(new_n200));
  INV_X1    g014(.A(G146), .ZN(new_n201));
  NAND3_X1  g015(.A1(new_n199), .A2(new_n200), .A3(new_n201), .ZN(new_n202));
  AND2_X1   g016(.A1(new_n193), .A2(new_n202), .ZN(new_n203));
  INV_X1    g017(.A(G237), .ZN(new_n204));
  INV_X1    g018(.A(G953), .ZN(new_n205));
  NAND3_X1  g019(.A1(new_n204), .A2(new_n205), .A3(G214), .ZN(new_n206));
  INV_X1    g020(.A(KEYINPUT86), .ZN(new_n207));
  INV_X1    g021(.A(G143), .ZN(new_n208));
  NAND3_X1  g022(.A1(new_n206), .A2(new_n207), .A3(new_n208), .ZN(new_n209));
  INV_X1    g023(.A(G131), .ZN(new_n210));
  NOR2_X1   g024(.A1(G237), .A2(G953), .ZN(new_n211));
  OAI211_X1 g025(.A(new_n211), .B(G214), .C1(KEYINPUT86), .C2(G143), .ZN(new_n212));
  NAND3_X1  g026(.A1(new_n209), .A2(new_n210), .A3(new_n212), .ZN(new_n213));
  INV_X1    g027(.A(KEYINPUT88), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n213), .A2(new_n214), .ZN(new_n215));
  AOI21_X1  g029(.A(new_n210), .B1(new_n209), .B2(new_n212), .ZN(new_n216));
  INV_X1    g030(.A(new_n216), .ZN(new_n217));
  INV_X1    g031(.A(KEYINPUT17), .ZN(new_n218));
  NAND4_X1  g032(.A1(new_n209), .A2(KEYINPUT88), .A3(new_n212), .A4(new_n210), .ZN(new_n219));
  NAND4_X1  g033(.A1(new_n215), .A2(new_n217), .A3(new_n218), .A4(new_n219), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n192), .A2(G146), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n216), .A2(KEYINPUT17), .ZN(new_n222));
  NAND4_X1  g036(.A1(new_n203), .A2(new_n220), .A3(new_n221), .A4(new_n222), .ZN(new_n223));
  XNOR2_X1  g037(.A(new_n191), .B(new_n201), .ZN(new_n224));
  NAND2_X1  g038(.A1(KEYINPUT18), .A2(G131), .ZN(new_n225));
  NAND3_X1  g039(.A1(new_n209), .A2(new_n212), .A3(new_n225), .ZN(new_n226));
  AND3_X1   g040(.A1(new_n216), .A2(KEYINPUT87), .A3(KEYINPUT18), .ZN(new_n227));
  AOI21_X1  g041(.A(KEYINPUT87), .B1(new_n216), .B2(KEYINPUT18), .ZN(new_n228));
  OAI211_X1 g042(.A(new_n224), .B(new_n226), .C1(new_n227), .C2(new_n228), .ZN(new_n229));
  XNOR2_X1  g043(.A(G113), .B(G122), .ZN(new_n230));
  INV_X1    g044(.A(G104), .ZN(new_n231));
  XNOR2_X1  g045(.A(new_n230), .B(new_n231), .ZN(new_n232));
  AND3_X1   g046(.A1(new_n223), .A2(new_n229), .A3(new_n232), .ZN(new_n233));
  NAND3_X1  g047(.A1(new_n215), .A2(new_n217), .A3(new_n219), .ZN(new_n234));
  INV_X1    g048(.A(KEYINPUT89), .ZN(new_n235));
  INV_X1    g049(.A(new_n191), .ZN(new_n236));
  OAI21_X1  g050(.A(new_n235), .B1(new_n236), .B2(KEYINPUT19), .ZN(new_n237));
  INV_X1    g051(.A(KEYINPUT19), .ZN(new_n238));
  NAND3_X1  g052(.A1(new_n191), .A2(KEYINPUT89), .A3(new_n238), .ZN(new_n239));
  OAI211_X1 g053(.A(new_n237), .B(new_n239), .C1(new_n238), .C2(new_n191), .ZN(new_n240));
  OAI211_X1 g054(.A(new_n234), .B(new_n221), .C1(G146), .C2(new_n240), .ZN(new_n241));
  AOI21_X1  g055(.A(new_n232), .B1(new_n241), .B2(new_n229), .ZN(new_n242));
  OAI211_X1 g056(.A(new_n187), .B(new_n188), .C1(new_n233), .C2(new_n242), .ZN(new_n243));
  INV_X1    g057(.A(KEYINPUT20), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n243), .A2(new_n244), .ZN(new_n245));
  NAND3_X1  g059(.A1(new_n223), .A2(new_n229), .A3(new_n232), .ZN(new_n246));
  AND2_X1   g060(.A1(new_n241), .A2(new_n229), .ZN(new_n247));
  OAI21_X1  g061(.A(new_n246), .B1(new_n247), .B2(new_n232), .ZN(new_n248));
  NAND4_X1  g062(.A1(new_n248), .A2(KEYINPUT20), .A3(new_n187), .A4(new_n188), .ZN(new_n249));
  AOI21_X1  g063(.A(new_n232), .B1(new_n223), .B2(new_n229), .ZN(new_n250));
  OAI21_X1  g064(.A(new_n188), .B1(new_n233), .B2(new_n250), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n251), .A2(G475), .ZN(new_n252));
  NAND3_X1  g066(.A1(new_n245), .A2(new_n249), .A3(new_n252), .ZN(new_n253));
  INV_X1    g067(.A(KEYINPUT90), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n253), .A2(new_n254), .ZN(new_n255));
  NAND4_X1  g069(.A1(new_n245), .A2(new_n252), .A3(new_n249), .A4(KEYINPUT90), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n255), .A2(new_n256), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n208), .A2(G128), .ZN(new_n258));
  XNOR2_X1  g072(.A(new_n258), .B(KEYINPUT91), .ZN(new_n259));
  OAI21_X1  g073(.A(new_n259), .B1(G128), .B2(new_n208), .ZN(new_n260));
  XNOR2_X1  g074(.A(new_n260), .B(G134), .ZN(new_n261));
  INV_X1    g075(.A(G116), .ZN(new_n262));
  NOR2_X1   g076(.A1(new_n262), .A2(G122), .ZN(new_n263));
  INV_X1    g077(.A(G122), .ZN(new_n264));
  NOR2_X1   g078(.A1(new_n264), .A2(G116), .ZN(new_n265));
  NOR2_X1   g079(.A1(new_n263), .A2(new_n265), .ZN(new_n266));
  INV_X1    g080(.A(G107), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n266), .A2(new_n267), .ZN(new_n268));
  INV_X1    g082(.A(KEYINPUT14), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n265), .A2(new_n269), .ZN(new_n270));
  AOI21_X1  g084(.A(new_n263), .B1(new_n270), .B2(KEYINPUT92), .ZN(new_n271));
  OAI21_X1  g085(.A(new_n271), .B1(KEYINPUT92), .B2(new_n270), .ZN(new_n272));
  NOR2_X1   g086(.A1(new_n265), .A2(new_n269), .ZN(new_n273));
  OAI21_X1  g087(.A(G107), .B1(new_n272), .B2(new_n273), .ZN(new_n274));
  NAND3_X1  g088(.A1(new_n261), .A2(new_n268), .A3(new_n274), .ZN(new_n275));
  INV_X1    g089(.A(KEYINPUT13), .ZN(new_n276));
  OAI22_X1  g090(.A1(new_n259), .A2(new_n276), .B1(G128), .B2(new_n208), .ZN(new_n277));
  AND2_X1   g091(.A1(new_n259), .A2(new_n276), .ZN(new_n278));
  OAI21_X1  g092(.A(G134), .B1(new_n277), .B2(new_n278), .ZN(new_n279));
  XNOR2_X1  g093(.A(new_n266), .B(new_n267), .ZN(new_n280));
  OAI211_X1 g094(.A(new_n279), .B(new_n280), .C1(G134), .C2(new_n260), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n275), .A2(new_n281), .ZN(new_n282));
  XOR2_X1   g096(.A(KEYINPUT9), .B(G234), .Z(new_n283));
  INV_X1    g097(.A(new_n283), .ZN(new_n284));
  INV_X1    g098(.A(G217), .ZN(new_n285));
  NOR3_X1   g099(.A1(new_n284), .A2(new_n285), .A3(G953), .ZN(new_n286));
  INV_X1    g100(.A(new_n286), .ZN(new_n287));
  NOR2_X1   g101(.A1(new_n282), .A2(new_n287), .ZN(new_n288));
  AOI21_X1  g102(.A(new_n286), .B1(new_n275), .B2(new_n281), .ZN(new_n289));
  OAI211_X1 g103(.A(KEYINPUT93), .B(new_n188), .C1(new_n288), .C2(new_n289), .ZN(new_n290));
  INV_X1    g104(.A(KEYINPUT15), .ZN(new_n291));
  NAND3_X1  g105(.A1(new_n290), .A2(new_n291), .A3(G478), .ZN(new_n292));
  XNOR2_X1  g106(.A(new_n282), .B(new_n287), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n291), .A2(G478), .ZN(new_n294));
  NAND4_X1  g108(.A1(new_n293), .A2(KEYINPUT93), .A3(new_n188), .A4(new_n294), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n292), .A2(new_n295), .ZN(new_n296));
  INV_X1    g110(.A(G952), .ZN(new_n297));
  NOR2_X1   g111(.A1(new_n297), .A2(G953), .ZN(new_n298));
  NAND2_X1  g112(.A1(G234), .A2(G237), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n298), .A2(new_n299), .ZN(new_n300));
  XOR2_X1   g114(.A(KEYINPUT21), .B(G898), .Z(new_n301));
  NAND3_X1  g115(.A1(new_n299), .A2(G902), .A3(G953), .ZN(new_n302));
  OAI21_X1  g116(.A(new_n300), .B1(new_n301), .B2(new_n302), .ZN(new_n303));
  INV_X1    g117(.A(new_n303), .ZN(new_n304));
  NOR3_X1   g118(.A1(new_n257), .A2(new_n296), .A3(new_n304), .ZN(new_n305));
  XNOR2_X1  g119(.A(G143), .B(G146), .ZN(new_n306));
  NAND3_X1  g120(.A1(new_n306), .A2(KEYINPUT0), .A3(G128), .ZN(new_n307));
  XNOR2_X1  g121(.A(KEYINPUT0), .B(G128), .ZN(new_n308));
  OAI21_X1  g122(.A(new_n307), .B1(new_n306), .B2(new_n308), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n309), .A2(G125), .ZN(new_n310));
  INV_X1    g124(.A(G128), .ZN(new_n311));
  NOR2_X1   g125(.A1(new_n311), .A2(KEYINPUT1), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n201), .A2(G143), .ZN(new_n313));
  NAND2_X1  g127(.A1(new_n208), .A2(G146), .ZN(new_n314));
  NAND3_X1  g128(.A1(new_n312), .A2(new_n313), .A3(new_n314), .ZN(new_n315));
  NAND3_X1  g129(.A1(new_n208), .A2(KEYINPUT1), .A3(G146), .ZN(new_n316));
  OAI211_X1 g130(.A(new_n315), .B(new_n316), .C1(G128), .C2(new_n306), .ZN(new_n317));
  OAI21_X1  g131(.A(new_n310), .B1(G125), .B2(new_n317), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n205), .A2(G224), .ZN(new_n319));
  XOR2_X1   g133(.A(new_n318), .B(new_n319), .Z(new_n320));
  INV_X1    g134(.A(KEYINPUT76), .ZN(new_n321));
  OAI21_X1  g135(.A(new_n321), .B1(new_n267), .B2(G104), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n267), .A2(G104), .ZN(new_n323));
  NAND3_X1  g137(.A1(new_n231), .A2(KEYINPUT76), .A3(G107), .ZN(new_n324));
  NAND3_X1  g138(.A1(new_n322), .A2(new_n323), .A3(new_n324), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n325), .A2(G101), .ZN(new_n326));
  INV_X1    g140(.A(G101), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n231), .A2(G107), .ZN(new_n328));
  AND3_X1   g142(.A1(new_n267), .A2(KEYINPUT3), .A3(G104), .ZN(new_n329));
  AOI21_X1  g143(.A(KEYINPUT3), .B1(new_n267), .B2(G104), .ZN(new_n330));
  OAI211_X1 g144(.A(new_n327), .B(new_n328), .C1(new_n329), .C2(new_n330), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n326), .A2(new_n331), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n332), .A2(KEYINPUT77), .ZN(new_n333));
  XOR2_X1   g147(.A(G116), .B(G119), .Z(new_n334));
  XNOR2_X1  g148(.A(KEYINPUT2), .B(G113), .ZN(new_n335));
  NOR2_X1   g149(.A1(new_n334), .A2(new_n335), .ZN(new_n336));
  NOR3_X1   g150(.A1(new_n262), .A2(KEYINPUT5), .A3(G119), .ZN(new_n337));
  XNOR2_X1  g151(.A(G116), .B(G119), .ZN(new_n338));
  AOI21_X1  g152(.A(new_n337), .B1(new_n338), .B2(KEYINPUT5), .ZN(new_n339));
  AOI21_X1  g153(.A(new_n336), .B1(G113), .B2(new_n339), .ZN(new_n340));
  AOI21_X1  g154(.A(KEYINPUT77), .B1(new_n325), .B2(G101), .ZN(new_n341));
  INV_X1    g155(.A(new_n341), .ZN(new_n342));
  NAND3_X1  g156(.A1(new_n333), .A2(new_n340), .A3(new_n342), .ZN(new_n343));
  OAI21_X1  g157(.A(new_n328), .B1(new_n329), .B2(new_n330), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n344), .A2(G101), .ZN(new_n345));
  NAND3_X1  g159(.A1(new_n345), .A2(KEYINPUT4), .A3(new_n331), .ZN(new_n346));
  XNOR2_X1  g160(.A(new_n334), .B(new_n335), .ZN(new_n347));
  INV_X1    g161(.A(KEYINPUT4), .ZN(new_n348));
  NAND3_X1  g162(.A1(new_n344), .A2(new_n348), .A3(G101), .ZN(new_n349));
  NAND3_X1  g163(.A1(new_n346), .A2(new_n347), .A3(new_n349), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n343), .A2(new_n350), .ZN(new_n351));
  XNOR2_X1  g165(.A(G110), .B(G122), .ZN(new_n352));
  XNOR2_X1  g166(.A(new_n352), .B(KEYINPUT83), .ZN(new_n353));
  NAND2_X1  g167(.A1(new_n351), .A2(new_n353), .ZN(new_n354));
  NAND3_X1  g168(.A1(new_n343), .A2(new_n350), .A3(new_n352), .ZN(new_n355));
  NAND3_X1  g169(.A1(new_n354), .A2(KEYINPUT6), .A3(new_n355), .ZN(new_n356));
  INV_X1    g170(.A(KEYINPUT84), .ZN(new_n357));
  INV_X1    g171(.A(KEYINPUT6), .ZN(new_n358));
  AND4_X1   g172(.A1(new_n357), .A2(new_n351), .A3(new_n358), .A4(new_n353), .ZN(new_n359));
  INV_X1    g173(.A(new_n353), .ZN(new_n360));
  AOI21_X1  g174(.A(new_n360), .B1(new_n343), .B2(new_n350), .ZN(new_n361));
  AOI21_X1  g175(.A(new_n357), .B1(new_n361), .B2(new_n358), .ZN(new_n362));
  OAI211_X1 g176(.A(new_n320), .B(new_n356), .C1(new_n359), .C2(new_n362), .ZN(new_n363));
  AND2_X1   g177(.A1(new_n319), .A2(KEYINPUT7), .ZN(new_n364));
  XNOR2_X1  g178(.A(new_n318), .B(new_n364), .ZN(new_n365));
  AOI21_X1  g179(.A(new_n341), .B1(new_n332), .B2(KEYINPUT77), .ZN(new_n366));
  XOR2_X1   g180(.A(new_n366), .B(new_n340), .Z(new_n367));
  XOR2_X1   g181(.A(new_n352), .B(KEYINPUT8), .Z(new_n368));
  OAI211_X1 g182(.A(new_n365), .B(new_n355), .C1(new_n367), .C2(new_n368), .ZN(new_n369));
  NAND3_X1  g183(.A1(new_n363), .A2(new_n188), .A3(new_n369), .ZN(new_n370));
  OAI21_X1  g184(.A(G210), .B1(G237), .B2(G902), .ZN(new_n371));
  INV_X1    g185(.A(new_n371), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n370), .A2(new_n372), .ZN(new_n373));
  NAND4_X1  g187(.A1(new_n363), .A2(new_n188), .A3(new_n371), .A4(new_n369), .ZN(new_n374));
  NAND3_X1  g188(.A1(new_n373), .A2(KEYINPUT85), .A3(new_n374), .ZN(new_n375));
  OR2_X1    g189(.A1(new_n374), .A2(KEYINPUT85), .ZN(new_n376));
  OAI21_X1  g190(.A(G214), .B1(G237), .B2(G902), .ZN(new_n377));
  AND3_X1   g191(.A1(new_n375), .A2(new_n376), .A3(new_n377), .ZN(new_n378));
  AND2_X1   g192(.A1(new_n305), .A2(new_n378), .ZN(new_n379));
  AOI21_X1  g193(.A(new_n285), .B1(G234), .B2(new_n188), .ZN(new_n380));
  NOR2_X1   g194(.A1(KEYINPUT74), .A2(KEYINPUT25), .ZN(new_n381));
  INV_X1    g195(.A(new_n381), .ZN(new_n382));
  NAND3_X1  g196(.A1(new_n193), .A2(new_n221), .A3(new_n202), .ZN(new_n383));
  INV_X1    g197(.A(KEYINPUT23), .ZN(new_n384));
  INV_X1    g198(.A(G119), .ZN(new_n385));
  OAI21_X1  g199(.A(new_n384), .B1(new_n385), .B2(G128), .ZN(new_n386));
  NAND2_X1  g200(.A1(new_n385), .A2(G128), .ZN(new_n387));
  NAND3_X1  g201(.A1(new_n311), .A2(KEYINPUT23), .A3(G119), .ZN(new_n388));
  NAND3_X1  g202(.A1(new_n386), .A2(new_n387), .A3(new_n388), .ZN(new_n389));
  INV_X1    g203(.A(KEYINPUT70), .ZN(new_n390));
  OR2_X1    g204(.A1(new_n389), .A2(new_n390), .ZN(new_n391));
  NAND2_X1  g205(.A1(new_n389), .A2(new_n390), .ZN(new_n392));
  NAND3_X1  g206(.A1(new_n391), .A2(new_n392), .A3(G110), .ZN(new_n393));
  XOR2_X1   g207(.A(KEYINPUT24), .B(G110), .Z(new_n394));
  XNOR2_X1  g208(.A(G119), .B(G128), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n394), .A2(new_n395), .ZN(new_n396));
  NAND3_X1  g210(.A1(new_n383), .A2(new_n393), .A3(new_n396), .ZN(new_n397));
  INV_X1    g211(.A(KEYINPUT72), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n397), .A2(new_n398), .ZN(new_n399));
  NAND4_X1  g213(.A1(new_n383), .A2(KEYINPUT72), .A3(new_n393), .A4(new_n396), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n399), .A2(new_n400), .ZN(new_n401));
  OAI22_X1  g215(.A1(new_n389), .A2(G110), .B1(new_n394), .B2(new_n395), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n191), .A2(new_n201), .ZN(new_n403));
  NAND3_X1  g217(.A1(new_n221), .A2(new_n402), .A3(new_n403), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n401), .A2(new_n404), .ZN(new_n405));
  INV_X1    g219(.A(KEYINPUT73), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n405), .A2(new_n406), .ZN(new_n407));
  NAND3_X1  g221(.A1(new_n205), .A2(G221), .A3(G234), .ZN(new_n408));
  XNOR2_X1  g222(.A(new_n408), .B(KEYINPUT22), .ZN(new_n409));
  XNOR2_X1  g223(.A(new_n409), .B(G137), .ZN(new_n410));
  INV_X1    g224(.A(new_n404), .ZN(new_n411));
  AOI21_X1  g225(.A(new_n411), .B1(new_n399), .B2(new_n400), .ZN(new_n412));
  AOI21_X1  g226(.A(new_n410), .B1(new_n412), .B2(KEYINPUT73), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n407), .A2(new_n413), .ZN(new_n414));
  NAND3_X1  g228(.A1(new_n405), .A2(new_n406), .A3(new_n410), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n414), .A2(new_n415), .ZN(new_n416));
  AOI21_X1  g230(.A(new_n382), .B1(new_n416), .B2(new_n188), .ZN(new_n417));
  AOI211_X1 g231(.A(G902), .B(new_n381), .C1(new_n414), .C2(new_n415), .ZN(new_n418));
  OAI21_X1  g232(.A(new_n380), .B1(new_n417), .B2(new_n418), .ZN(new_n419));
  INV_X1    g233(.A(KEYINPUT75), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n419), .A2(new_n420), .ZN(new_n421));
  OAI211_X1 g235(.A(KEYINPUT75), .B(new_n380), .C1(new_n417), .C2(new_n418), .ZN(new_n422));
  NOR2_X1   g236(.A1(new_n380), .A2(G902), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n416), .A2(new_n423), .ZN(new_n424));
  AND3_X1   g238(.A1(new_n421), .A2(new_n422), .A3(new_n424), .ZN(new_n425));
  OAI21_X1  g239(.A(G221), .B1(new_n284), .B2(G902), .ZN(new_n426));
  INV_X1    g240(.A(new_n426), .ZN(new_n427));
  INV_X1    g241(.A(G469), .ZN(new_n428));
  NOR2_X1   g242(.A1(new_n428), .A2(new_n188), .ZN(new_n429));
  NOR2_X1   g243(.A1(new_n366), .A2(new_n317), .ZN(new_n430));
  NAND3_X1  g244(.A1(new_n333), .A2(new_n342), .A3(new_n317), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n431), .A2(KEYINPUT78), .ZN(new_n432));
  INV_X1    g246(.A(KEYINPUT78), .ZN(new_n433));
  NAND3_X1  g247(.A1(new_n366), .A2(new_n433), .A3(new_n317), .ZN(new_n434));
  AOI21_X1  g248(.A(new_n430), .B1(new_n432), .B2(new_n434), .ZN(new_n435));
  INV_X1    g249(.A(KEYINPUT64), .ZN(new_n436));
  INV_X1    g250(.A(G134), .ZN(new_n437));
  OAI21_X1  g251(.A(new_n436), .B1(new_n437), .B2(G137), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n438), .A2(KEYINPUT11), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n437), .A2(G137), .ZN(new_n440));
  INV_X1    g254(.A(KEYINPUT11), .ZN(new_n441));
  OAI211_X1 g255(.A(new_n436), .B(new_n441), .C1(new_n437), .C2(G137), .ZN(new_n442));
  NAND3_X1  g256(.A1(new_n439), .A2(new_n440), .A3(new_n442), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n443), .A2(G131), .ZN(new_n444));
  NAND4_X1  g258(.A1(new_n439), .A2(new_n210), .A3(new_n440), .A4(new_n442), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n444), .A2(new_n445), .ZN(new_n446));
  INV_X1    g260(.A(new_n446), .ZN(new_n447));
  OAI21_X1  g261(.A(KEYINPUT12), .B1(new_n435), .B2(new_n447), .ZN(new_n448));
  INV_X1    g262(.A(KEYINPUT10), .ZN(new_n449));
  AOI21_X1  g263(.A(new_n433), .B1(new_n366), .B2(new_n317), .ZN(new_n450));
  INV_X1    g264(.A(KEYINPUT77), .ZN(new_n451));
  AOI21_X1  g265(.A(new_n451), .B1(new_n326), .B2(new_n331), .ZN(new_n452));
  AND3_X1   g266(.A1(new_n312), .A2(new_n313), .A3(new_n314), .ZN(new_n453));
  AOI21_X1  g267(.A(G128), .B1(new_n313), .B2(new_n314), .ZN(new_n454));
  INV_X1    g268(.A(new_n316), .ZN(new_n455));
  NOR3_X1   g269(.A1(new_n453), .A2(new_n454), .A3(new_n455), .ZN(new_n456));
  NOR4_X1   g270(.A1(new_n452), .A2(new_n456), .A3(KEYINPUT78), .A4(new_n341), .ZN(new_n457));
  OAI21_X1  g271(.A(new_n449), .B1(new_n450), .B2(new_n457), .ZN(new_n458));
  AND2_X1   g272(.A1(new_n346), .A2(new_n349), .ZN(new_n459));
  INV_X1    g273(.A(new_n309), .ZN(new_n460));
  NOR3_X1   g274(.A1(new_n452), .A2(new_n341), .A3(new_n456), .ZN(new_n461));
  AOI22_X1  g275(.A1(new_n459), .A2(new_n460), .B1(new_n461), .B2(KEYINPUT10), .ZN(new_n462));
  NAND3_X1  g276(.A1(new_n458), .A2(new_n447), .A3(new_n462), .ZN(new_n463));
  XNOR2_X1  g277(.A(G110), .B(G140), .ZN(new_n464));
  INV_X1    g278(.A(G227), .ZN(new_n465));
  NOR2_X1   g279(.A1(new_n465), .A2(G953), .ZN(new_n466));
  XOR2_X1   g280(.A(new_n464), .B(new_n466), .Z(new_n467));
  OAI22_X1  g281(.A1(new_n450), .A2(new_n457), .B1(new_n366), .B2(new_n317), .ZN(new_n468));
  INV_X1    g282(.A(KEYINPUT12), .ZN(new_n469));
  NAND3_X1  g283(.A1(new_n468), .A2(new_n469), .A3(new_n446), .ZN(new_n470));
  NAND4_X1  g284(.A1(new_n448), .A2(new_n463), .A3(new_n467), .A4(new_n470), .ZN(new_n471));
  INV_X1    g285(.A(KEYINPUT82), .ZN(new_n472));
  XNOR2_X1  g286(.A(new_n471), .B(new_n472), .ZN(new_n473));
  INV_X1    g287(.A(new_n467), .ZN(new_n474));
  INV_X1    g288(.A(KEYINPUT80), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n458), .A2(new_n462), .ZN(new_n476));
  AOI21_X1  g290(.A(new_n475), .B1(new_n476), .B2(new_n446), .ZN(new_n477));
  AOI211_X1 g291(.A(KEYINPUT80), .B(new_n447), .C1(new_n458), .C2(new_n462), .ZN(new_n478));
  NOR2_X1   g292(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  INV_X1    g293(.A(new_n463), .ZN(new_n480));
  OAI21_X1  g294(.A(new_n474), .B1(new_n479), .B2(new_n480), .ZN(new_n481));
  AOI21_X1  g295(.A(G902), .B1(new_n473), .B2(new_n481), .ZN(new_n482));
  AOI21_X1  g296(.A(new_n429), .B1(new_n482), .B2(new_n428), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n463), .A2(new_n467), .ZN(new_n484));
  NAND2_X1  g298(.A1(new_n484), .A2(KEYINPUT79), .ZN(new_n485));
  INV_X1    g299(.A(KEYINPUT79), .ZN(new_n486));
  NAND3_X1  g300(.A1(new_n463), .A2(new_n486), .A3(new_n467), .ZN(new_n487));
  OAI211_X1 g301(.A(new_n485), .B(new_n487), .C1(new_n478), .C2(new_n477), .ZN(new_n488));
  NAND3_X1  g302(.A1(new_n448), .A2(new_n463), .A3(new_n470), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n489), .A2(new_n474), .ZN(new_n490));
  NAND3_X1  g304(.A1(new_n488), .A2(KEYINPUT81), .A3(new_n490), .ZN(new_n491));
  INV_X1    g305(.A(new_n491), .ZN(new_n492));
  AOI21_X1  g306(.A(KEYINPUT81), .B1(new_n488), .B2(new_n490), .ZN(new_n493));
  OAI21_X1  g307(.A(G469), .B1(new_n492), .B2(new_n493), .ZN(new_n494));
  AOI21_X1  g308(.A(new_n427), .B1(new_n483), .B2(new_n494), .ZN(new_n495));
  INV_X1    g309(.A(KEYINPUT66), .ZN(new_n496));
  INV_X1    g310(.A(new_n347), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n446), .A2(new_n460), .ZN(new_n498));
  INV_X1    g312(.A(new_n440), .ZN(new_n499));
  NOR2_X1   g313(.A1(new_n437), .A2(G137), .ZN(new_n500));
  OAI21_X1  g314(.A(G131), .B1(new_n499), .B2(new_n500), .ZN(new_n501));
  AND3_X1   g315(.A1(new_n317), .A2(new_n445), .A3(new_n501), .ZN(new_n502));
  INV_X1    g316(.A(new_n502), .ZN(new_n503));
  AOI21_X1  g317(.A(new_n497), .B1(new_n498), .B2(new_n503), .ZN(new_n504));
  AOI21_X1  g318(.A(new_n309), .B1(new_n444), .B2(new_n445), .ZN(new_n505));
  NOR3_X1   g319(.A1(new_n505), .A2(new_n502), .A3(new_n347), .ZN(new_n506));
  OAI211_X1 g320(.A(new_n496), .B(KEYINPUT28), .C1(new_n504), .C2(new_n506), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n211), .A2(G210), .ZN(new_n508));
  XNOR2_X1  g322(.A(new_n508), .B(KEYINPUT27), .ZN(new_n509));
  NAND2_X1  g323(.A1(new_n509), .A2(KEYINPUT26), .ZN(new_n510));
  INV_X1    g324(.A(KEYINPUT27), .ZN(new_n511));
  XNOR2_X1  g325(.A(new_n508), .B(new_n511), .ZN(new_n512));
  INV_X1    g326(.A(KEYINPUT26), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  AOI21_X1  g328(.A(G101), .B1(new_n510), .B2(new_n514), .ZN(new_n515));
  INV_X1    g329(.A(new_n515), .ZN(new_n516));
  NAND3_X1  g330(.A1(new_n510), .A2(new_n514), .A3(G101), .ZN(new_n517));
  NAND3_X1  g331(.A1(new_n516), .A2(KEYINPUT65), .A3(new_n517), .ZN(new_n518));
  INV_X1    g332(.A(KEYINPUT65), .ZN(new_n519));
  INV_X1    g333(.A(new_n517), .ZN(new_n520));
  OAI21_X1  g334(.A(new_n519), .B1(new_n520), .B2(new_n515), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n518), .A2(new_n521), .ZN(new_n522));
  INV_X1    g336(.A(KEYINPUT28), .ZN(new_n523));
  NAND3_X1  g337(.A1(new_n498), .A2(new_n503), .A3(new_n497), .ZN(new_n524));
  OAI21_X1  g338(.A(new_n347), .B1(new_n505), .B2(new_n502), .ZN(new_n525));
  AOI21_X1  g339(.A(new_n523), .B1(new_n524), .B2(new_n525), .ZN(new_n526));
  OAI21_X1  g340(.A(KEYINPUT66), .B1(new_n506), .B2(KEYINPUT28), .ZN(new_n527));
  OAI211_X1 g341(.A(new_n507), .B(new_n522), .C1(new_n526), .C2(new_n527), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n528), .A2(KEYINPUT67), .ZN(new_n529));
  NAND3_X1  g343(.A1(new_n498), .A2(new_n503), .A3(KEYINPUT30), .ZN(new_n530));
  INV_X1    g344(.A(KEYINPUT30), .ZN(new_n531));
  OAI21_X1  g345(.A(new_n531), .B1(new_n505), .B2(new_n502), .ZN(new_n532));
  NAND3_X1  g346(.A1(new_n530), .A2(new_n347), .A3(new_n532), .ZN(new_n533));
  NOR2_X1   g347(.A1(new_n520), .A2(new_n515), .ZN(new_n534));
  NAND3_X1  g348(.A1(new_n533), .A2(new_n524), .A3(new_n534), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n535), .A2(KEYINPUT31), .ZN(new_n536));
  OR2_X1    g350(.A1(new_n535), .A2(KEYINPUT31), .ZN(new_n537));
  OAI21_X1  g351(.A(KEYINPUT28), .B1(new_n504), .B2(new_n506), .ZN(new_n538));
  AOI21_X1  g352(.A(new_n496), .B1(new_n524), .B2(new_n523), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n538), .A2(new_n539), .ZN(new_n540));
  INV_X1    g354(.A(KEYINPUT67), .ZN(new_n541));
  NAND4_X1  g355(.A1(new_n540), .A2(new_n541), .A3(new_n522), .A4(new_n507), .ZN(new_n542));
  NAND4_X1  g356(.A1(new_n529), .A2(new_n536), .A3(new_n537), .A4(new_n542), .ZN(new_n543));
  NOR2_X1   g357(.A1(G472), .A2(G902), .ZN(new_n544));
  NAND2_X1  g358(.A1(new_n543), .A2(new_n544), .ZN(new_n545));
  INV_X1    g359(.A(KEYINPUT68), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n545), .A2(new_n546), .ZN(new_n547));
  AND3_X1   g361(.A1(new_n543), .A2(KEYINPUT32), .A3(new_n544), .ZN(new_n548));
  AOI21_X1  g362(.A(KEYINPUT32), .B1(new_n543), .B2(new_n544), .ZN(new_n549));
  OAI21_X1  g363(.A(new_n547), .B1(new_n548), .B2(new_n549), .ZN(new_n550));
  AOI21_X1  g364(.A(new_n522), .B1(new_n540), .B2(new_n507), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n533), .A2(new_n524), .ZN(new_n552));
  INV_X1    g366(.A(new_n534), .ZN(new_n553));
  AOI211_X1 g367(.A(KEYINPUT29), .B(new_n551), .C1(new_n552), .C2(new_n553), .ZN(new_n554));
  OAI21_X1  g368(.A(KEYINPUT69), .B1(new_n506), .B2(KEYINPUT28), .ZN(new_n555));
  OR2_X1    g369(.A1(new_n526), .A2(new_n555), .ZN(new_n556));
  OAI21_X1  g370(.A(new_n556), .B1(KEYINPUT69), .B2(new_n538), .ZN(new_n557));
  NAND3_X1  g371(.A1(new_n557), .A2(KEYINPUT29), .A3(new_n534), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n558), .A2(new_n188), .ZN(new_n559));
  OAI21_X1  g373(.A(G472), .B1(new_n554), .B2(new_n559), .ZN(new_n560));
  NAND3_X1  g374(.A1(new_n545), .A2(new_n546), .A3(KEYINPUT32), .ZN(new_n561));
  NAND3_X1  g375(.A1(new_n550), .A2(new_n560), .A3(new_n561), .ZN(new_n562));
  AND4_X1   g376(.A1(new_n379), .A2(new_n425), .A3(new_n495), .A4(new_n562), .ZN(new_n563));
  XNOR2_X1  g377(.A(new_n563), .B(new_n327), .ZN(G3));
  NAND2_X1  g378(.A1(new_n543), .A2(new_n188), .ZN(new_n565));
  AOI22_X1  g379(.A1(new_n565), .A2(G472), .B1(new_n544), .B2(new_n543), .ZN(new_n566));
  NAND3_X1  g380(.A1(new_n425), .A2(new_n495), .A3(new_n566), .ZN(new_n567));
  INV_X1    g381(.A(new_n567), .ZN(new_n568));
  INV_X1    g382(.A(KEYINPUT33), .ZN(new_n569));
  XNOR2_X1  g383(.A(new_n293), .B(new_n569), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n188), .A2(G478), .ZN(new_n571));
  AND2_X1   g385(.A1(new_n293), .A2(new_n188), .ZN(new_n572));
  OAI22_X1  g386(.A1(new_n570), .A2(new_n571), .B1(G478), .B2(new_n572), .ZN(new_n573));
  NAND2_X1  g387(.A1(new_n573), .A2(new_n257), .ZN(new_n574));
  INV_X1    g388(.A(new_n377), .ZN(new_n575));
  AOI21_X1  g389(.A(new_n575), .B1(new_n373), .B2(new_n374), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n576), .A2(new_n303), .ZN(new_n577));
  NOR2_X1   g391(.A1(new_n574), .A2(new_n577), .ZN(new_n578));
  NAND2_X1  g392(.A1(new_n568), .A2(new_n578), .ZN(new_n579));
  XOR2_X1   g393(.A(KEYINPUT34), .B(G104), .Z(new_n580));
  XNOR2_X1  g394(.A(new_n579), .B(new_n580), .ZN(new_n581));
  XNOR2_X1  g395(.A(KEYINPUT94), .B(KEYINPUT95), .ZN(new_n582));
  XNOR2_X1  g396(.A(new_n581), .B(new_n582), .ZN(G6));
  XNOR2_X1  g397(.A(new_n290), .B(new_n294), .ZN(new_n584));
  NOR3_X1   g398(.A1(new_n577), .A2(new_n253), .A3(new_n584), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n568), .A2(new_n585), .ZN(new_n586));
  XOR2_X1   g400(.A(KEYINPUT35), .B(G107), .Z(new_n587));
  XNOR2_X1  g401(.A(new_n586), .B(new_n587), .ZN(G9));
  INV_X1    g402(.A(KEYINPUT36), .ZN(new_n589));
  NAND2_X1  g403(.A1(new_n410), .A2(new_n589), .ZN(new_n590));
  XNOR2_X1  g404(.A(new_n412), .B(new_n590), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n591), .A2(new_n423), .ZN(new_n592));
  NAND3_X1  g406(.A1(new_n421), .A2(new_n422), .A3(new_n592), .ZN(new_n593));
  NAND4_X1  g407(.A1(new_n495), .A2(new_n379), .A3(new_n566), .A4(new_n593), .ZN(new_n594));
  XOR2_X1   g408(.A(new_n594), .B(KEYINPUT37), .Z(new_n595));
  XNOR2_X1  g409(.A(new_n595), .B(G110), .ZN(G12));
  AND2_X1   g410(.A1(new_n593), .A2(new_n562), .ZN(new_n597));
  XNOR2_X1  g411(.A(new_n300), .B(KEYINPUT96), .ZN(new_n598));
  INV_X1    g412(.A(new_n598), .ZN(new_n599));
  OAI21_X1  g413(.A(new_n599), .B1(G900), .B2(new_n302), .ZN(new_n600));
  INV_X1    g414(.A(new_n600), .ZN(new_n601));
  NOR2_X1   g415(.A1(new_n253), .A2(new_n601), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n602), .A2(new_n296), .ZN(new_n603));
  INV_X1    g417(.A(new_n603), .ZN(new_n604));
  NAND4_X1  g418(.A1(new_n597), .A2(new_n495), .A3(new_n576), .A4(new_n604), .ZN(new_n605));
  XNOR2_X1  g419(.A(new_n605), .B(G128), .ZN(G30));
  NAND2_X1  g420(.A1(new_n375), .A2(new_n376), .ZN(new_n607));
  XNOR2_X1  g421(.A(new_n607), .B(KEYINPUT38), .ZN(new_n608));
  XOR2_X1   g422(.A(new_n600), .B(KEYINPUT39), .Z(new_n609));
  INV_X1    g423(.A(new_n609), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n495), .A2(new_n610), .ZN(new_n611));
  AOI211_X1 g425(.A(new_n593), .B(new_n608), .C1(new_n611), .C2(KEYINPUT40), .ZN(new_n612));
  OAI21_X1  g426(.A(new_n522), .B1(new_n506), .B2(new_n504), .ZN(new_n613));
  AND2_X1   g427(.A1(new_n613), .A2(new_n535), .ZN(new_n614));
  OAI21_X1  g428(.A(G472), .B1(new_n614), .B2(G902), .ZN(new_n615));
  NAND3_X1  g429(.A1(new_n550), .A2(new_n561), .A3(new_n615), .ZN(new_n616));
  INV_X1    g430(.A(new_n616), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n257), .A2(new_n296), .ZN(new_n618));
  NOR3_X1   g432(.A1(new_n617), .A2(new_n575), .A3(new_n618), .ZN(new_n619));
  OAI211_X1 g433(.A(new_n612), .B(new_n619), .C1(KEYINPUT40), .C2(new_n611), .ZN(new_n620));
  XNOR2_X1  g434(.A(new_n620), .B(G143), .ZN(G45));
  NOR2_X1   g435(.A1(new_n574), .A2(new_n601), .ZN(new_n622));
  NAND4_X1  g436(.A1(new_n597), .A2(new_n495), .A3(new_n576), .A4(new_n622), .ZN(new_n623));
  XNOR2_X1  g437(.A(new_n623), .B(G146), .ZN(G48));
  NAND3_X1  g438(.A1(new_n346), .A2(new_n460), .A3(new_n349), .ZN(new_n625));
  OAI21_X1  g439(.A(new_n625), .B1(new_n431), .B2(new_n449), .ZN(new_n626));
  NAND2_X1  g440(.A1(new_n432), .A2(new_n434), .ZN(new_n627));
  AOI21_X1  g441(.A(new_n626), .B1(new_n627), .B2(new_n449), .ZN(new_n628));
  AOI21_X1  g442(.A(new_n474), .B1(new_n628), .B2(new_n447), .ZN(new_n629));
  NAND4_X1  g443(.A1(new_n629), .A2(new_n472), .A3(new_n448), .A4(new_n470), .ZN(new_n630));
  NAND2_X1  g444(.A1(new_n471), .A2(KEYINPUT82), .ZN(new_n631));
  OAI21_X1  g445(.A(KEYINPUT80), .B1(new_n628), .B2(new_n447), .ZN(new_n632));
  NAND3_X1  g446(.A1(new_n476), .A2(new_n475), .A3(new_n446), .ZN(new_n633));
  AOI21_X1  g447(.A(new_n480), .B1(new_n632), .B2(new_n633), .ZN(new_n634));
  OAI211_X1 g448(.A(new_n630), .B(new_n631), .C1(new_n634), .C2(new_n467), .ZN(new_n635));
  NAND3_X1  g449(.A1(new_n635), .A2(new_n428), .A3(new_n188), .ZN(new_n636));
  INV_X1    g450(.A(new_n636), .ZN(new_n637));
  AOI21_X1  g451(.A(new_n428), .B1(new_n635), .B2(new_n188), .ZN(new_n638));
  NOR3_X1   g452(.A1(new_n637), .A2(new_n638), .A3(new_n427), .ZN(new_n639));
  NAND4_X1  g453(.A1(new_n425), .A2(new_n562), .A3(new_n578), .A4(new_n639), .ZN(new_n640));
  XNOR2_X1  g454(.A(KEYINPUT41), .B(G113), .ZN(new_n641));
  XNOR2_X1  g455(.A(new_n640), .B(new_n641), .ZN(G15));
  NAND4_X1  g456(.A1(new_n425), .A2(new_n585), .A3(new_n562), .A4(new_n639), .ZN(new_n643));
  XNOR2_X1  g457(.A(new_n643), .B(G116), .ZN(G18));
  INV_X1    g458(.A(new_n576), .ZN(new_n645));
  NOR4_X1   g459(.A1(new_n637), .A2(new_n638), .A3(new_n645), .A4(new_n427), .ZN(new_n646));
  NAND4_X1  g460(.A1(new_n646), .A2(new_n305), .A3(new_n562), .A4(new_n593), .ZN(new_n647));
  XNOR2_X1  g461(.A(new_n647), .B(G119), .ZN(G21));
  INV_X1    g462(.A(new_n522), .ZN(new_n649));
  OAI211_X1 g463(.A(new_n536), .B(new_n537), .C1(new_n557), .C2(new_n649), .ZN(new_n650));
  AOI22_X1  g464(.A1(new_n565), .A2(G472), .B1(new_n544), .B2(new_n650), .ZN(new_n651));
  AND4_X1   g465(.A1(new_n421), .A2(new_n422), .A3(new_n424), .A4(new_n651), .ZN(new_n652));
  NOR2_X1   g466(.A1(new_n577), .A2(new_n584), .ZN(new_n653));
  NAND4_X1  g467(.A1(new_n652), .A2(new_n257), .A3(new_n653), .A4(new_n639), .ZN(new_n654));
  XNOR2_X1  g468(.A(new_n654), .B(G122), .ZN(G24));
  AND3_X1   g469(.A1(new_n593), .A2(new_n622), .A3(new_n651), .ZN(new_n656));
  NAND2_X1  g470(.A1(new_n656), .A2(new_n646), .ZN(new_n657));
  XNOR2_X1  g471(.A(new_n657), .B(G125), .ZN(G27));
  INV_X1    g472(.A(KEYINPUT98), .ZN(new_n659));
  INV_X1    g473(.A(new_n429), .ZN(new_n660));
  NAND3_X1  g474(.A1(new_n488), .A2(G469), .A3(new_n490), .ZN(new_n661));
  NAND3_X1  g475(.A1(new_n636), .A2(new_n660), .A3(new_n661), .ZN(new_n662));
  AND2_X1   g476(.A1(new_n662), .A2(new_n426), .ZN(new_n663));
  INV_X1    g477(.A(KEYINPUT97), .ZN(new_n664));
  AOI21_X1  g478(.A(new_n664), .B1(new_n607), .B2(new_n377), .ZN(new_n665));
  AOI211_X1 g479(.A(KEYINPUT97), .B(new_n575), .C1(new_n375), .C2(new_n376), .ZN(new_n666));
  NOR2_X1   g480(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  NAND4_X1  g481(.A1(new_n425), .A2(new_n663), .A3(new_n667), .A4(new_n562), .ZN(new_n668));
  INV_X1    g482(.A(new_n622), .ZN(new_n669));
  OAI21_X1  g483(.A(new_n659), .B1(new_n668), .B2(new_n669), .ZN(new_n670));
  XNOR2_X1  g484(.A(KEYINPUT99), .B(KEYINPUT42), .ZN(new_n671));
  INV_X1    g485(.A(new_n562), .ZN(new_n672));
  NAND3_X1  g486(.A1(new_n421), .A2(new_n422), .A3(new_n424), .ZN(new_n673));
  NOR2_X1   g487(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  NAND2_X1  g488(.A1(new_n662), .A2(new_n426), .ZN(new_n675));
  NOR3_X1   g489(.A1(new_n675), .A2(new_n666), .A3(new_n665), .ZN(new_n676));
  NAND4_X1  g490(.A1(new_n674), .A2(new_n676), .A3(KEYINPUT98), .A4(new_n622), .ZN(new_n677));
  NAND3_X1  g491(.A1(new_n670), .A2(new_n671), .A3(new_n677), .ZN(new_n678));
  NOR2_X1   g492(.A1(new_n548), .A2(new_n549), .ZN(new_n679));
  AOI21_X1  g493(.A(new_n673), .B1(new_n679), .B2(new_n560), .ZN(new_n680));
  NAND4_X1  g494(.A1(new_n680), .A2(KEYINPUT42), .A3(new_n676), .A4(new_n622), .ZN(new_n681));
  NAND2_X1  g495(.A1(new_n678), .A2(new_n681), .ZN(new_n682));
  XNOR2_X1  g496(.A(new_n682), .B(G131), .ZN(G33));
  NOR2_X1   g497(.A1(new_n668), .A2(new_n603), .ZN(new_n684));
  XOR2_X1   g498(.A(KEYINPUT100), .B(G134), .Z(new_n685));
  XNOR2_X1  g499(.A(new_n684), .B(new_n685), .ZN(G36));
  NAND3_X1  g500(.A1(new_n488), .A2(KEYINPUT45), .A3(new_n490), .ZN(new_n687));
  NAND2_X1  g501(.A1(new_n485), .A2(new_n487), .ZN(new_n688));
  OAI21_X1  g502(.A(new_n490), .B1(new_n688), .B2(new_n479), .ZN(new_n689));
  INV_X1    g503(.A(KEYINPUT81), .ZN(new_n690));
  NAND2_X1  g504(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  NAND2_X1  g505(.A1(new_n691), .A2(new_n491), .ZN(new_n692));
  OAI211_X1 g506(.A(G469), .B(new_n687), .C1(new_n692), .C2(KEYINPUT45), .ZN(new_n693));
  XNOR2_X1  g507(.A(new_n693), .B(KEYINPUT101), .ZN(new_n694));
  NAND2_X1  g508(.A1(new_n694), .A2(new_n660), .ZN(new_n695));
  INV_X1    g509(.A(KEYINPUT46), .ZN(new_n696));
  OAI21_X1  g510(.A(new_n636), .B1(new_n695), .B2(new_n696), .ZN(new_n697));
  INV_X1    g511(.A(KEYINPUT102), .ZN(new_n698));
  NAND2_X1  g512(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  NAND2_X1  g513(.A1(new_n695), .A2(new_n696), .ZN(new_n700));
  OAI211_X1 g514(.A(KEYINPUT102), .B(new_n636), .C1(new_n695), .C2(new_n696), .ZN(new_n701));
  NAND3_X1  g515(.A1(new_n699), .A2(new_n700), .A3(new_n701), .ZN(new_n702));
  NAND2_X1  g516(.A1(new_n702), .A2(new_n426), .ZN(new_n703));
  NOR2_X1   g517(.A1(new_n703), .A2(new_n609), .ZN(new_n704));
  NAND3_X1  g518(.A1(new_n573), .A2(new_n255), .A3(new_n256), .ZN(new_n705));
  XOR2_X1   g519(.A(new_n705), .B(KEYINPUT43), .Z(new_n706));
  INV_X1    g520(.A(new_n706), .ZN(new_n707));
  INV_X1    g521(.A(new_n593), .ZN(new_n708));
  NOR3_X1   g522(.A1(new_n707), .A2(new_n566), .A3(new_n708), .ZN(new_n709));
  XOR2_X1   g523(.A(new_n709), .B(KEYINPUT44), .Z(new_n710));
  NAND3_X1  g524(.A1(new_n704), .A2(new_n667), .A3(new_n710), .ZN(new_n711));
  XNOR2_X1  g525(.A(new_n711), .B(G137), .ZN(G39));
  OR2_X1    g526(.A1(new_n703), .A2(KEYINPUT47), .ZN(new_n713));
  NAND2_X1  g527(.A1(new_n703), .A2(KEYINPUT47), .ZN(new_n714));
  NAND2_X1  g528(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  INV_X1    g529(.A(new_n667), .ZN(new_n716));
  NOR3_X1   g530(.A1(new_n715), .A2(new_n669), .A3(new_n716), .ZN(new_n717));
  NOR2_X1   g531(.A1(new_n425), .A2(new_n562), .ZN(new_n718));
  NAND2_X1  g532(.A1(new_n717), .A2(new_n718), .ZN(new_n719));
  XNOR2_X1  g533(.A(new_n719), .B(G140), .ZN(G42));
  NAND2_X1  g534(.A1(new_n297), .A2(new_n205), .ZN(new_n721));
  XNOR2_X1  g535(.A(new_n721), .B(KEYINPUT112), .ZN(new_n722));
  NAND2_X1  g536(.A1(new_n706), .A2(new_n598), .ZN(new_n723));
  INV_X1    g537(.A(new_n723), .ZN(new_n724));
  NAND2_X1  g538(.A1(new_n724), .A2(new_n652), .ZN(new_n725));
  INV_X1    g539(.A(new_n639), .ZN(new_n726));
  NOR2_X1   g540(.A1(new_n725), .A2(new_n726), .ZN(new_n727));
  NAND3_X1  g541(.A1(new_n727), .A2(new_n575), .A3(new_n608), .ZN(new_n728));
  INV_X1    g542(.A(KEYINPUT50), .ZN(new_n729));
  XNOR2_X1  g543(.A(new_n728), .B(new_n729), .ZN(new_n730));
  NOR2_X1   g544(.A1(new_n716), .A2(new_n726), .ZN(new_n731));
  NAND4_X1  g545(.A1(new_n724), .A2(new_n593), .A3(new_n651), .A4(new_n731), .ZN(new_n732));
  NOR2_X1   g546(.A1(new_n673), .A2(new_n300), .ZN(new_n733));
  NAND3_X1  g547(.A1(new_n731), .A2(new_n617), .A3(new_n733), .ZN(new_n734));
  OR3_X1    g548(.A1(new_n734), .A2(new_n257), .A3(new_n573), .ZN(new_n735));
  AND3_X1   g549(.A1(new_n730), .A2(new_n732), .A3(new_n735), .ZN(new_n736));
  NAND2_X1  g550(.A1(new_n736), .A2(KEYINPUT110), .ZN(new_n737));
  NAND4_X1  g551(.A1(new_n730), .A2(KEYINPUT51), .A3(new_n732), .A4(new_n735), .ZN(new_n738));
  INV_X1    g552(.A(KEYINPUT110), .ZN(new_n739));
  NAND2_X1  g553(.A1(new_n738), .A2(new_n739), .ZN(new_n740));
  NOR3_X1   g554(.A1(new_n637), .A2(new_n638), .A3(new_n426), .ZN(new_n741));
  AOI21_X1  g555(.A(new_n741), .B1(new_n713), .B2(new_n714), .ZN(new_n742));
  NOR2_X1   g556(.A1(new_n725), .A2(new_n716), .ZN(new_n743));
  INV_X1    g557(.A(new_n743), .ZN(new_n744));
  OAI211_X1 g558(.A(new_n737), .B(new_n740), .C1(new_n742), .C2(new_n744), .ZN(new_n745));
  NAND3_X1  g559(.A1(new_n724), .A2(new_n680), .A3(new_n731), .ZN(new_n746));
  OR2_X1    g560(.A1(KEYINPUT111), .A2(KEYINPUT48), .ZN(new_n747));
  NAND2_X1  g561(.A1(KEYINPUT111), .A2(KEYINPUT48), .ZN(new_n748));
  NAND3_X1  g562(.A1(new_n746), .A2(new_n747), .A3(new_n748), .ZN(new_n749));
  OR2_X1    g563(.A1(new_n746), .A2(new_n748), .ZN(new_n750));
  OR2_X1    g564(.A1(new_n734), .A2(new_n574), .ZN(new_n751));
  AND3_X1   g565(.A1(new_n750), .A2(new_n298), .A3(new_n751), .ZN(new_n752));
  NAND3_X1  g566(.A1(new_n745), .A2(new_n749), .A3(new_n752), .ZN(new_n753));
  NAND3_X1  g567(.A1(new_n257), .A2(new_n296), .A3(new_n576), .ZN(new_n754));
  NOR2_X1   g568(.A1(new_n675), .A2(new_n754), .ZN(new_n755));
  NAND4_X1  g569(.A1(new_n755), .A2(new_n708), .A3(new_n600), .A4(new_n616), .ZN(new_n756));
  NAND4_X1  g570(.A1(new_n605), .A2(new_n623), .A3(new_n657), .A4(new_n756), .ZN(new_n757));
  INV_X1    g571(.A(KEYINPUT52), .ZN(new_n758));
  NAND2_X1  g572(.A1(new_n757), .A2(new_n758), .ZN(new_n759));
  NAND3_X1  g573(.A1(new_n593), .A2(new_n562), .A3(new_n576), .ZN(new_n760));
  NAND2_X1  g574(.A1(new_n636), .A2(new_n660), .ZN(new_n761));
  AOI21_X1  g575(.A(new_n428), .B1(new_n691), .B2(new_n491), .ZN(new_n762));
  OAI21_X1  g576(.A(new_n426), .B1(new_n761), .B2(new_n762), .ZN(new_n763));
  NOR2_X1   g577(.A1(new_n760), .A2(new_n763), .ZN(new_n764));
  AOI22_X1  g578(.A1(new_n764), .A2(new_n622), .B1(new_n646), .B2(new_n656), .ZN(new_n765));
  NAND4_X1  g579(.A1(new_n765), .A2(KEYINPUT52), .A3(new_n605), .A4(new_n756), .ZN(new_n766));
  NAND2_X1  g580(.A1(new_n759), .A2(new_n766), .ZN(new_n767));
  AOI21_X1  g581(.A(new_n684), .B1(new_n678), .B2(new_n681), .ZN(new_n768));
  NAND3_X1  g582(.A1(new_n667), .A2(new_n562), .A3(new_n602), .ZN(new_n769));
  NOR4_X1   g583(.A1(new_n769), .A2(new_n708), .A3(new_n296), .A4(new_n763), .ZN(new_n770));
  INV_X1    g584(.A(new_n770), .ZN(new_n771));
  AND3_X1   g585(.A1(new_n767), .A2(new_n768), .A3(new_n771), .ZN(new_n772));
  OAI211_X1 g586(.A(new_n566), .B(new_n426), .C1(new_n761), .C2(new_n762), .ZN(new_n773));
  NAND4_X1  g587(.A1(new_n375), .A2(new_n376), .A3(new_n377), .A4(new_n303), .ZN(new_n774));
  NOR4_X1   g588(.A1(new_n773), .A2(new_n673), .A3(new_n574), .A4(new_n774), .ZN(new_n775));
  NOR2_X1   g589(.A1(new_n563), .A2(new_n775), .ZN(new_n776));
  AND4_X1   g590(.A1(new_n640), .A2(new_n654), .A3(new_n643), .A4(new_n647), .ZN(new_n777));
  INV_X1    g591(.A(KEYINPUT104), .ZN(new_n778));
  AND3_X1   g592(.A1(new_n255), .A2(new_n296), .A3(new_n256), .ZN(new_n779));
  NAND4_X1  g593(.A1(new_n378), .A2(KEYINPUT103), .A3(new_n303), .A4(new_n779), .ZN(new_n780));
  INV_X1    g594(.A(KEYINPUT103), .ZN(new_n781));
  NAND3_X1  g595(.A1(new_n255), .A2(new_n296), .A3(new_n256), .ZN(new_n782));
  OAI21_X1  g596(.A(new_n781), .B1(new_n774), .B2(new_n782), .ZN(new_n783));
  NAND2_X1  g597(.A1(new_n780), .A2(new_n783), .ZN(new_n784));
  OAI211_X1 g598(.A(new_n594), .B(new_n778), .C1(new_n567), .C2(new_n784), .ZN(new_n785));
  INV_X1    g599(.A(new_n785), .ZN(new_n786));
  AND2_X1   g600(.A1(new_n780), .A2(new_n783), .ZN(new_n787));
  INV_X1    g601(.A(new_n773), .ZN(new_n788));
  NAND3_X1  g602(.A1(new_n787), .A2(new_n788), .A3(new_n425), .ZN(new_n789));
  AOI21_X1  g603(.A(new_n778), .B1(new_n789), .B2(new_n594), .ZN(new_n790));
  OAI211_X1 g604(.A(new_n776), .B(new_n777), .C1(new_n786), .C2(new_n790), .ZN(new_n791));
  NAND2_X1  g605(.A1(new_n656), .A2(new_n676), .ZN(new_n792));
  INV_X1    g606(.A(new_n792), .ZN(new_n793));
  NOR2_X1   g607(.A1(new_n791), .A2(new_n793), .ZN(new_n794));
  NAND4_X1  g608(.A1(new_n772), .A2(KEYINPUT107), .A3(KEYINPUT53), .A4(new_n794), .ZN(new_n795));
  AOI211_X1 g609(.A(new_n684), .B(new_n770), .C1(new_n678), .C2(new_n681), .ZN(new_n796));
  NAND4_X1  g610(.A1(new_n794), .A2(new_n796), .A3(KEYINPUT53), .A4(new_n767), .ZN(new_n797));
  INV_X1    g611(.A(KEYINPUT107), .ZN(new_n798));
  NAND2_X1  g612(.A1(new_n797), .A2(new_n798), .ZN(new_n799));
  NAND2_X1  g613(.A1(new_n795), .A2(new_n799), .ZN(new_n800));
  INV_X1    g614(.A(KEYINPUT54), .ZN(new_n801));
  NAND3_X1  g615(.A1(new_n794), .A2(new_n767), .A3(new_n796), .ZN(new_n802));
  INV_X1    g616(.A(KEYINPUT53), .ZN(new_n803));
  AOI21_X1  g617(.A(KEYINPUT106), .B1(new_n802), .B2(new_n803), .ZN(new_n804));
  AND3_X1   g618(.A1(new_n802), .A2(KEYINPUT106), .A3(new_n803), .ZN(new_n805));
  OAI211_X1 g619(.A(new_n800), .B(new_n801), .C1(new_n804), .C2(new_n805), .ZN(new_n806));
  INV_X1    g620(.A(KEYINPUT108), .ZN(new_n807));
  NAND2_X1  g621(.A1(new_n806), .A2(new_n807), .ZN(new_n808));
  NAND3_X1  g622(.A1(new_n767), .A2(new_n768), .A3(new_n771), .ZN(new_n809));
  OR2_X1    g623(.A1(new_n786), .A2(new_n790), .ZN(new_n810));
  NAND4_X1  g624(.A1(new_n810), .A2(new_n792), .A3(new_n776), .A4(new_n777), .ZN(new_n811));
  OAI21_X1  g625(.A(new_n803), .B1(new_n809), .B2(new_n811), .ZN(new_n812));
  AOI21_X1  g626(.A(new_n801), .B1(new_n812), .B2(new_n797), .ZN(new_n813));
  XNOR2_X1  g627(.A(new_n813), .B(KEYINPUT105), .ZN(new_n814));
  INV_X1    g628(.A(KEYINPUT106), .ZN(new_n815));
  NAND2_X1  g629(.A1(new_n812), .A2(new_n815), .ZN(new_n816));
  NAND3_X1  g630(.A1(new_n802), .A2(KEYINPUT106), .A3(new_n803), .ZN(new_n817));
  AOI22_X1  g631(.A1(new_n816), .A2(new_n817), .B1(new_n795), .B2(new_n799), .ZN(new_n818));
  NAND3_X1  g632(.A1(new_n818), .A2(KEYINPUT108), .A3(new_n801), .ZN(new_n819));
  NAND3_X1  g633(.A1(new_n808), .A2(new_n814), .A3(new_n819), .ZN(new_n820));
  XOR2_X1   g634(.A(new_n741), .B(KEYINPUT109), .Z(new_n821));
  NAND2_X1  g635(.A1(new_n715), .A2(new_n821), .ZN(new_n822));
  NAND2_X1  g636(.A1(new_n822), .A2(new_n743), .ZN(new_n823));
  AOI21_X1  g637(.A(KEYINPUT51), .B1(new_n823), .B2(new_n736), .ZN(new_n824));
  OR3_X1    g638(.A1(new_n753), .A2(new_n820), .A3(new_n824), .ZN(new_n825));
  NOR3_X1   g639(.A1(new_n725), .A2(new_n645), .A3(new_n726), .ZN(new_n826));
  OAI21_X1  g640(.A(new_n722), .B1(new_n825), .B2(new_n826), .ZN(new_n827));
  NOR3_X1   g641(.A1(new_n705), .A2(new_n575), .A3(new_n427), .ZN(new_n828));
  NAND4_X1  g642(.A1(new_n425), .A2(new_n617), .A3(new_n828), .A4(new_n608), .ZN(new_n829));
  NOR2_X1   g643(.A1(new_n637), .A2(new_n638), .ZN(new_n830));
  XOR2_X1   g644(.A(new_n830), .B(KEYINPUT49), .Z(new_n831));
  OAI21_X1  g645(.A(new_n827), .B1(new_n829), .B2(new_n831), .ZN(G75));
  OAI21_X1  g646(.A(new_n356), .B1(new_n359), .B2(new_n362), .ZN(new_n833));
  XNOR2_X1  g647(.A(new_n833), .B(new_n320), .ZN(new_n834));
  XOR2_X1   g648(.A(new_n834), .B(KEYINPUT55), .Z(new_n835));
  OAI21_X1  g649(.A(new_n800), .B1(new_n804), .B2(new_n805), .ZN(new_n836));
  NAND3_X1  g650(.A1(new_n836), .A2(G210), .A3(G902), .ZN(new_n837));
  INV_X1    g651(.A(KEYINPUT113), .ZN(new_n838));
  NAND2_X1  g652(.A1(new_n837), .A2(new_n838), .ZN(new_n839));
  INV_X1    g653(.A(KEYINPUT56), .ZN(new_n840));
  NAND2_X1  g654(.A1(new_n839), .A2(new_n840), .ZN(new_n841));
  NOR2_X1   g655(.A1(new_n837), .A2(new_n838), .ZN(new_n842));
  OAI21_X1  g656(.A(new_n835), .B1(new_n841), .B2(new_n842), .ZN(new_n843));
  NOR2_X1   g657(.A1(new_n205), .A2(G952), .ZN(new_n844));
  INV_X1    g658(.A(new_n844), .ZN(new_n845));
  AOI21_X1  g659(.A(KEYINPUT56), .B1(new_n837), .B2(KEYINPUT114), .ZN(new_n846));
  INV_X1    g660(.A(new_n835), .ZN(new_n847));
  OAI211_X1 g661(.A(new_n846), .B(new_n847), .C1(KEYINPUT114), .C2(new_n837), .ZN(new_n848));
  NAND3_X1  g662(.A1(new_n843), .A2(new_n845), .A3(new_n848), .ZN(new_n849));
  INV_X1    g663(.A(KEYINPUT115), .ZN(new_n850));
  NAND2_X1  g664(.A1(new_n849), .A2(new_n850), .ZN(new_n851));
  NAND4_X1  g665(.A1(new_n843), .A2(KEYINPUT115), .A3(new_n848), .A4(new_n845), .ZN(new_n852));
  NAND2_X1  g666(.A1(new_n851), .A2(new_n852), .ZN(G51));
  OAI21_X1  g667(.A(KEYINPUT116), .B1(new_n818), .B2(new_n801), .ZN(new_n854));
  INV_X1    g668(.A(KEYINPUT116), .ZN(new_n855));
  NOR2_X1   g669(.A1(new_n805), .A2(new_n804), .ZN(new_n856));
  XNOR2_X1  g670(.A(new_n797), .B(KEYINPUT107), .ZN(new_n857));
  OAI211_X1 g671(.A(new_n855), .B(KEYINPUT54), .C1(new_n856), .C2(new_n857), .ZN(new_n858));
  NAND3_X1  g672(.A1(new_n854), .A2(new_n858), .A3(new_n806), .ZN(new_n859));
  XNOR2_X1  g673(.A(new_n429), .B(KEYINPUT57), .ZN(new_n860));
  NAND2_X1  g674(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  NAND2_X1  g675(.A1(new_n861), .A2(new_n635), .ZN(new_n862));
  OR3_X1    g676(.A1(new_n818), .A2(new_n188), .A3(new_n694), .ZN(new_n863));
  AOI21_X1  g677(.A(new_n844), .B1(new_n862), .B2(new_n863), .ZN(G54));
  NAND4_X1  g678(.A1(new_n836), .A2(KEYINPUT58), .A3(G475), .A4(G902), .ZN(new_n865));
  XOR2_X1   g679(.A(new_n865), .B(new_n248), .Z(new_n866));
  NOR2_X1   g680(.A1(new_n866), .A2(new_n844), .ZN(G60));
  XNOR2_X1  g681(.A(KEYINPUT118), .B(KEYINPUT59), .ZN(new_n868));
  NAND2_X1  g682(.A1(G478), .A2(G902), .ZN(new_n869));
  XOR2_X1   g683(.A(new_n868), .B(new_n869), .Z(new_n870));
  NAND2_X1  g684(.A1(new_n820), .A2(new_n870), .ZN(new_n871));
  XNOR2_X1  g685(.A(new_n570), .B(KEYINPUT117), .ZN(new_n872));
  NAND2_X1  g686(.A1(new_n871), .A2(new_n872), .ZN(new_n873));
  INV_X1    g687(.A(new_n870), .ZN(new_n874));
  NOR2_X1   g688(.A1(new_n872), .A2(new_n874), .ZN(new_n875));
  NAND2_X1  g689(.A1(new_n859), .A2(new_n875), .ZN(new_n876));
  NAND2_X1  g690(.A1(new_n876), .A2(KEYINPUT119), .ZN(new_n877));
  INV_X1    g691(.A(KEYINPUT119), .ZN(new_n878));
  NAND3_X1  g692(.A1(new_n859), .A2(new_n878), .A3(new_n875), .ZN(new_n879));
  NAND4_X1  g693(.A1(new_n873), .A2(new_n877), .A3(new_n845), .A4(new_n879), .ZN(new_n880));
  INV_X1    g694(.A(KEYINPUT120), .ZN(new_n881));
  NAND2_X1  g695(.A1(new_n880), .A2(new_n881), .ZN(new_n882));
  AOI21_X1  g696(.A(new_n844), .B1(new_n871), .B2(new_n872), .ZN(new_n883));
  NAND4_X1  g697(.A1(new_n883), .A2(KEYINPUT120), .A3(new_n877), .A4(new_n879), .ZN(new_n884));
  NAND2_X1  g698(.A1(new_n882), .A2(new_n884), .ZN(G63));
  INV_X1    g699(.A(KEYINPUT61), .ZN(new_n886));
  NAND2_X1  g700(.A1(G217), .A2(G902), .ZN(new_n887));
  XNOR2_X1  g701(.A(new_n887), .B(KEYINPUT122), .ZN(new_n888));
  XOR2_X1   g702(.A(KEYINPUT121), .B(KEYINPUT60), .Z(new_n889));
  XNOR2_X1  g703(.A(new_n888), .B(new_n889), .ZN(new_n890));
  NAND2_X1  g704(.A1(new_n836), .A2(new_n890), .ZN(new_n891));
  NAND3_X1  g705(.A1(new_n891), .A2(new_n415), .A3(new_n414), .ZN(new_n892));
  NAND3_X1  g706(.A1(new_n892), .A2(KEYINPUT123), .A3(new_n845), .ZN(new_n893));
  NAND3_X1  g707(.A1(new_n836), .A2(new_n591), .A3(new_n890), .ZN(new_n894));
  NAND2_X1  g708(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  AOI21_X1  g709(.A(KEYINPUT123), .B1(new_n892), .B2(new_n845), .ZN(new_n896));
  OAI21_X1  g710(.A(new_n886), .B1(new_n895), .B2(new_n896), .ZN(new_n897));
  INV_X1    g711(.A(KEYINPUT124), .ZN(new_n898));
  OR2_X1    g712(.A1(new_n892), .A2(new_n898), .ZN(new_n899));
  AOI21_X1  g713(.A(new_n886), .B1(new_n892), .B2(new_n898), .ZN(new_n900));
  NAND4_X1  g714(.A1(new_n899), .A2(new_n900), .A3(new_n845), .A4(new_n894), .ZN(new_n901));
  NAND2_X1  g715(.A1(new_n897), .A2(new_n901), .ZN(G66));
  AOI21_X1  g716(.A(new_n205), .B1(new_n301), .B2(G224), .ZN(new_n903));
  AOI21_X1  g717(.A(new_n903), .B1(new_n791), .B2(new_n205), .ZN(new_n904));
  OAI21_X1  g718(.A(new_n833), .B1(G898), .B2(new_n205), .ZN(new_n905));
  XOR2_X1   g719(.A(new_n904), .B(new_n905), .Z(G69));
  INV_X1    g720(.A(new_n754), .ZN(new_n907));
  NAND3_X1  g721(.A1(new_n704), .A2(new_n680), .A3(new_n907), .ZN(new_n908));
  NAND2_X1  g722(.A1(new_n765), .A2(new_n605), .ZN(new_n909));
  INV_X1    g723(.A(new_n909), .ZN(new_n910));
  AND2_X1   g724(.A1(new_n768), .A2(new_n910), .ZN(new_n911));
  NAND4_X1  g725(.A1(new_n719), .A2(new_n711), .A3(new_n908), .A4(new_n911), .ZN(new_n912));
  NAND2_X1  g726(.A1(new_n912), .A2(new_n205), .ZN(new_n913));
  NAND3_X1  g727(.A1(new_n465), .A2(G900), .A3(G953), .ZN(new_n914));
  NAND2_X1  g728(.A1(new_n913), .A2(new_n914), .ZN(new_n915));
  NAND2_X1  g729(.A1(new_n530), .A2(new_n532), .ZN(new_n916));
  XNOR2_X1  g730(.A(new_n240), .B(KEYINPUT125), .ZN(new_n917));
  XNOR2_X1  g731(.A(new_n916), .B(new_n917), .ZN(new_n918));
  INV_X1    g732(.A(new_n611), .ZN(new_n919));
  NAND2_X1  g733(.A1(new_n574), .A2(new_n782), .ZN(new_n920));
  NAND4_X1  g734(.A1(new_n919), .A2(new_n674), .A3(new_n667), .A4(new_n920), .ZN(new_n921));
  NAND2_X1  g735(.A1(new_n910), .A2(new_n620), .ZN(new_n922));
  XOR2_X1   g736(.A(new_n922), .B(KEYINPUT62), .Z(new_n923));
  NAND4_X1  g737(.A1(new_n719), .A2(new_n711), .A3(new_n921), .A4(new_n923), .ZN(new_n924));
  AOI21_X1  g738(.A(new_n918), .B1(new_n924), .B2(new_n205), .ZN(new_n925));
  INV_X1    g739(.A(G900), .ZN(new_n926));
  OAI21_X1  g740(.A(G953), .B1(new_n465), .B2(new_n926), .ZN(new_n927));
  AOI22_X1  g741(.A1(new_n915), .A2(new_n918), .B1(new_n925), .B2(new_n927), .ZN(G72));
  NAND2_X1  g742(.A1(G472), .A2(G902), .ZN(new_n929));
  XOR2_X1   g743(.A(new_n929), .B(KEYINPUT127), .Z(new_n930));
  XNOR2_X1  g744(.A(new_n930), .B(KEYINPUT126), .ZN(new_n931));
  XNOR2_X1  g745(.A(new_n931), .B(KEYINPUT63), .ZN(new_n932));
  OAI21_X1  g746(.A(new_n932), .B1(new_n912), .B2(new_n791), .ZN(new_n933));
  NAND4_X1  g747(.A1(new_n933), .A2(new_n524), .A3(new_n533), .A4(new_n553), .ZN(new_n934));
  OAI21_X1  g748(.A(new_n932), .B1(new_n924), .B2(new_n791), .ZN(new_n935));
  NAND3_X1  g749(.A1(new_n935), .A2(new_n552), .A3(new_n534), .ZN(new_n936));
  NAND2_X1  g750(.A1(new_n812), .A2(new_n797), .ZN(new_n937));
  NAND2_X1  g751(.A1(new_n552), .A2(new_n553), .ZN(new_n938));
  NAND2_X1  g752(.A1(new_n938), .A2(new_n535), .ZN(new_n939));
  NAND3_X1  g753(.A1(new_n937), .A2(new_n932), .A3(new_n939), .ZN(new_n940));
  AND4_X1   g754(.A1(new_n845), .A2(new_n934), .A3(new_n936), .A4(new_n940), .ZN(G57));
endmodule


