

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300,
         n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311,
         n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322,
         n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333,
         n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344,
         n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355,
         n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
         n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
         n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
         n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
         n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410,
         n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421,
         n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432,
         n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443,
         n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454,
         n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465,
         n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
         n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487,
         n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
         n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
         n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583, n584, n585;

  XOR2_X1 U322 ( .A(KEYINPUT91), .B(n331), .Z(n290) );
  XOR2_X1 U323 ( .A(n338), .B(n429), .Z(n291) );
  XOR2_X1 U324 ( .A(n333), .B(KEYINPUT22), .Z(n292) );
  XNOR2_X1 U325 ( .A(KEYINPUT87), .B(KEYINPUT24), .ZN(n328) );
  XNOR2_X1 U326 ( .A(n463), .B(n462), .ZN(n464) );
  INV_X1 U327 ( .A(KEYINPUT9), .ZN(n403) );
  NOR2_X1 U328 ( .A1(n527), .A2(n384), .ZN(n385) );
  XNOR2_X1 U329 ( .A(n404), .B(n403), .ZN(n405) );
  XNOR2_X1 U330 ( .A(n345), .B(n372), .ZN(n472) );
  XNOR2_X1 U331 ( .A(n406), .B(n405), .ZN(n415) );
  XOR2_X1 U332 ( .A(KEYINPUT78), .B(n555), .Z(n562) );
  NOR2_X1 U333 ( .A1(n475), .A2(n517), .ZN(n563) );
  XOR2_X1 U334 ( .A(KEYINPUT38), .B(n454), .Z(n496) );
  XNOR2_X1 U335 ( .A(n477), .B(n476), .ZN(n478) );
  XNOR2_X1 U336 ( .A(G43GAT), .B(KEYINPUT40), .ZN(n455) );
  XNOR2_X1 U337 ( .A(n479), .B(n478), .ZN(G1349GAT) );
  XNOR2_X1 U338 ( .A(n456), .B(n455), .ZN(G1330GAT) );
  XOR2_X1 U339 ( .A(G78GAT), .B(G64GAT), .Z(n294) );
  XNOR2_X1 U340 ( .A(G22GAT), .B(G71GAT), .ZN(n293) );
  XNOR2_X1 U341 ( .A(n294), .B(n293), .ZN(n307) );
  XOR2_X1 U342 ( .A(KEYINPUT13), .B(G57GAT), .Z(n430) );
  XOR2_X1 U343 ( .A(G155GAT), .B(n430), .Z(n296) );
  NAND2_X1 U344 ( .A1(G231GAT), .A2(G233GAT), .ZN(n295) );
  XNOR2_X1 U345 ( .A(n296), .B(n295), .ZN(n300) );
  XOR2_X1 U346 ( .A(KEYINPUT14), .B(G211GAT), .Z(n298) );
  XNOR2_X1 U347 ( .A(G183GAT), .B(KEYINPUT15), .ZN(n297) );
  XNOR2_X1 U348 ( .A(n298), .B(n297), .ZN(n299) );
  XOR2_X1 U349 ( .A(n300), .B(n299), .Z(n305) );
  XOR2_X1 U350 ( .A(G15GAT), .B(G127GAT), .Z(n324) );
  XOR2_X1 U351 ( .A(KEYINPUT79), .B(KEYINPUT12), .Z(n302) );
  XNOR2_X1 U352 ( .A(G8GAT), .B(G1GAT), .ZN(n301) );
  XNOR2_X1 U353 ( .A(n302), .B(n301), .ZN(n303) );
  XNOR2_X1 U354 ( .A(n324), .B(n303), .ZN(n304) );
  XNOR2_X1 U355 ( .A(n305), .B(n304), .ZN(n306) );
  XOR2_X1 U356 ( .A(n307), .B(n306), .Z(n577) );
  XOR2_X1 U357 ( .A(KEYINPUT17), .B(G183GAT), .Z(n309) );
  XNOR2_X1 U358 ( .A(KEYINPUT19), .B(KEYINPUT18), .ZN(n308) );
  XNOR2_X1 U359 ( .A(n309), .B(n308), .ZN(n310) );
  XOR2_X1 U360 ( .A(KEYINPUT85), .B(n310), .Z(n380) );
  XOR2_X1 U361 ( .A(G99GAT), .B(G190GAT), .Z(n312) );
  XNOR2_X1 U362 ( .A(G43GAT), .B(G134GAT), .ZN(n311) );
  XNOR2_X1 U363 ( .A(n312), .B(n311), .ZN(n316) );
  XOR2_X1 U364 ( .A(KEYINPUT86), .B(KEYINPUT83), .Z(n314) );
  XNOR2_X1 U365 ( .A(G169GAT), .B(G176GAT), .ZN(n313) );
  XNOR2_X1 U366 ( .A(n314), .B(n313), .ZN(n315) );
  XOR2_X1 U367 ( .A(n316), .B(n315), .Z(n321) );
  XOR2_X1 U368 ( .A(KEYINPUT82), .B(KEYINPUT20), .Z(n318) );
  NAND2_X1 U369 ( .A1(G227GAT), .A2(G233GAT), .ZN(n317) );
  XNOR2_X1 U370 ( .A(n318), .B(n317), .ZN(n319) );
  XNOR2_X1 U371 ( .A(KEYINPUT84), .B(n319), .ZN(n320) );
  XNOR2_X1 U372 ( .A(n321), .B(n320), .ZN(n323) );
  XNOR2_X1 U373 ( .A(G113GAT), .B(KEYINPUT0), .ZN(n322) );
  XNOR2_X1 U374 ( .A(n322), .B(KEYINPUT81), .ZN(n363) );
  XOR2_X1 U375 ( .A(n323), .B(n363), .Z(n326) );
  XOR2_X1 U376 ( .A(G120GAT), .B(G71GAT), .Z(n423) );
  XNOR2_X1 U377 ( .A(n423), .B(n324), .ZN(n325) );
  XNOR2_X1 U378 ( .A(n326), .B(n325), .ZN(n327) );
  XNOR2_X1 U379 ( .A(n380), .B(n327), .ZN(n517) );
  INV_X1 U380 ( .A(n517), .ZN(n527) );
  INV_X1 U381 ( .A(n328), .ZN(n330) );
  XNOR2_X1 U382 ( .A(KEYINPUT23), .B(KEYINPUT92), .ZN(n329) );
  XNOR2_X1 U383 ( .A(n330), .B(n329), .ZN(n331) );
  NAND2_X1 U384 ( .A1(G228GAT), .A2(G233GAT), .ZN(n332) );
  XNOR2_X1 U385 ( .A(n290), .B(n332), .ZN(n333) );
  XOR2_X1 U386 ( .A(KEYINPUT90), .B(KEYINPUT89), .Z(n335) );
  XNOR2_X1 U387 ( .A(G155GAT), .B(KEYINPUT2), .ZN(n334) );
  XNOR2_X1 U388 ( .A(n335), .B(n334), .ZN(n336) );
  XOR2_X1 U389 ( .A(KEYINPUT3), .B(n336), .Z(n349) );
  XNOR2_X1 U390 ( .A(G106GAT), .B(n349), .ZN(n337) );
  XNOR2_X1 U391 ( .A(n292), .B(n337), .ZN(n338) );
  XOR2_X1 U392 ( .A(G78GAT), .B(G148GAT), .Z(n429) );
  XOR2_X1 U393 ( .A(G141GAT), .B(G22GAT), .Z(n447) );
  XOR2_X1 U394 ( .A(G162GAT), .B(KEYINPUT76), .Z(n340) );
  XNOR2_X1 U395 ( .A(G50GAT), .B(G218GAT), .ZN(n339) );
  XNOR2_X1 U396 ( .A(n340), .B(n339), .ZN(n402) );
  XNOR2_X1 U397 ( .A(n447), .B(n402), .ZN(n341) );
  XNOR2_X1 U398 ( .A(n291), .B(n341), .ZN(n345) );
  XOR2_X1 U399 ( .A(KEYINPUT88), .B(KEYINPUT21), .Z(n343) );
  XNOR2_X1 U400 ( .A(G197GAT), .B(G204GAT), .ZN(n342) );
  XNOR2_X1 U401 ( .A(n343), .B(n342), .ZN(n344) );
  XNOR2_X1 U402 ( .A(G211GAT), .B(n344), .ZN(n372) );
  XNOR2_X1 U403 ( .A(n472), .B(KEYINPUT65), .ZN(n346) );
  XNOR2_X1 U404 ( .A(n346), .B(KEYINPUT28), .ZN(n530) );
  XOR2_X1 U405 ( .A(KEYINPUT4), .B(KEYINPUT95), .Z(n348) );
  XNOR2_X1 U406 ( .A(KEYINPUT93), .B(KEYINPUT5), .ZN(n347) );
  XNOR2_X1 U407 ( .A(n348), .B(n347), .ZN(n350) );
  XOR2_X1 U408 ( .A(n350), .B(n349), .Z(n358) );
  XOR2_X1 U409 ( .A(KEYINPUT94), .B(KEYINPUT96), .Z(n352) );
  XNOR2_X1 U410 ( .A(KEYINPUT97), .B(KEYINPUT6), .ZN(n351) );
  XNOR2_X1 U411 ( .A(n352), .B(n351), .ZN(n356) );
  XOR2_X1 U412 ( .A(KEYINPUT1), .B(KEYINPUT98), .Z(n354) );
  XNOR2_X1 U413 ( .A(G127GAT), .B(KEYINPUT99), .ZN(n353) );
  XNOR2_X1 U414 ( .A(n354), .B(n353), .ZN(n355) );
  XNOR2_X1 U415 ( .A(n356), .B(n355), .ZN(n357) );
  XNOR2_X1 U416 ( .A(n358), .B(n357), .ZN(n362) );
  XOR2_X1 U417 ( .A(G85GAT), .B(G162GAT), .Z(n360) );
  XNOR2_X1 U418 ( .A(G29GAT), .B(G120GAT), .ZN(n359) );
  XNOR2_X1 U419 ( .A(n360), .B(n359), .ZN(n361) );
  XOR2_X1 U420 ( .A(n362), .B(n361), .Z(n371) );
  XOR2_X1 U421 ( .A(G134GAT), .B(KEYINPUT77), .Z(n399) );
  XOR2_X1 U422 ( .A(n399), .B(n363), .Z(n365) );
  NAND2_X1 U423 ( .A1(G225GAT), .A2(G233GAT), .ZN(n364) );
  XNOR2_X1 U424 ( .A(n365), .B(n364), .ZN(n369) );
  XOR2_X1 U425 ( .A(G148GAT), .B(G57GAT), .Z(n367) );
  XNOR2_X1 U426 ( .A(G141GAT), .B(G1GAT), .ZN(n366) );
  XNOR2_X1 U427 ( .A(n367), .B(n366), .ZN(n368) );
  XNOR2_X1 U428 ( .A(n369), .B(n368), .ZN(n370) );
  XNOR2_X1 U429 ( .A(n371), .B(n370), .ZN(n501) );
  INV_X1 U430 ( .A(n372), .ZN(n373) );
  XOR2_X1 U431 ( .A(n373), .B(G92GAT), .Z(n375) );
  XOR2_X1 U432 ( .A(G169GAT), .B(G8GAT), .Z(n443) );
  XNOR2_X1 U433 ( .A(n443), .B(G218GAT), .ZN(n374) );
  XNOR2_X1 U434 ( .A(n375), .B(n374), .ZN(n379) );
  XOR2_X1 U435 ( .A(G176GAT), .B(G64GAT), .Z(n421) );
  XOR2_X1 U436 ( .A(n421), .B(KEYINPUT100), .Z(n377) );
  NAND2_X1 U437 ( .A1(G226GAT), .A2(G233GAT), .ZN(n376) );
  XNOR2_X1 U438 ( .A(n377), .B(n376), .ZN(n378) );
  XOR2_X1 U439 ( .A(n379), .B(n378), .Z(n382) );
  XOR2_X1 U440 ( .A(G36GAT), .B(G190GAT), .Z(n411) );
  XNOR2_X1 U441 ( .A(n380), .B(n411), .ZN(n381) );
  XNOR2_X1 U442 ( .A(n382), .B(n381), .ZN(n515) );
  XOR2_X1 U443 ( .A(n515), .B(KEYINPUT27), .Z(n387) );
  NAND2_X1 U444 ( .A1(n501), .A2(n387), .ZN(n525) );
  NOR2_X1 U445 ( .A1(n530), .A2(n525), .ZN(n383) );
  XNOR2_X1 U446 ( .A(n383), .B(KEYINPUT101), .ZN(n384) );
  XNOR2_X1 U447 ( .A(n385), .B(KEYINPUT102), .ZN(n396) );
  NOR2_X1 U448 ( .A1(n472), .A2(n527), .ZN(n386) );
  XNOR2_X1 U449 ( .A(n386), .B(KEYINPUT26), .ZN(n568) );
  NAND2_X1 U450 ( .A1(n387), .A2(n568), .ZN(n388) );
  XNOR2_X1 U451 ( .A(KEYINPUT103), .B(n388), .ZN(n393) );
  INV_X1 U452 ( .A(n515), .ZN(n504) );
  NAND2_X1 U453 ( .A1(n504), .A2(n527), .ZN(n389) );
  NAND2_X1 U454 ( .A1(n389), .A2(n472), .ZN(n390) );
  XNOR2_X1 U455 ( .A(n390), .B(KEYINPUT25), .ZN(n391) );
  XNOR2_X1 U456 ( .A(n391), .B(KEYINPUT104), .ZN(n392) );
  NOR2_X1 U457 ( .A1(n393), .A2(n392), .ZN(n394) );
  NOR2_X1 U458 ( .A1(n501), .A2(n394), .ZN(n395) );
  NOR2_X1 U459 ( .A1(n396), .A2(n395), .ZN(n483) );
  NOR2_X1 U460 ( .A1(n577), .A2(n483), .ZN(n416) );
  XOR2_X1 U461 ( .A(G85GAT), .B(G92GAT), .Z(n398) );
  XNOR2_X1 U462 ( .A(G99GAT), .B(G106GAT), .ZN(n397) );
  XNOR2_X1 U463 ( .A(n398), .B(n397), .ZN(n422) );
  XOR2_X1 U464 ( .A(n422), .B(n399), .Z(n401) );
  NAND2_X1 U465 ( .A1(G232GAT), .A2(G233GAT), .ZN(n400) );
  XNOR2_X1 U466 ( .A(n401), .B(n400), .ZN(n406) );
  XNOR2_X1 U467 ( .A(n402), .B(KEYINPUT64), .ZN(n404) );
  XOR2_X1 U468 ( .A(KEYINPUT11), .B(KEYINPUT10), .Z(n413) );
  XOR2_X1 U469 ( .A(G29GAT), .B(KEYINPUT70), .Z(n408) );
  XNOR2_X1 U470 ( .A(KEYINPUT8), .B(G43GAT), .ZN(n407) );
  XNOR2_X1 U471 ( .A(n408), .B(n407), .ZN(n410) );
  XOR2_X1 U472 ( .A(KEYINPUT7), .B(KEYINPUT71), .Z(n409) );
  XOR2_X1 U473 ( .A(n410), .B(n409), .Z(n453) );
  XNOR2_X1 U474 ( .A(n453), .B(n411), .ZN(n412) );
  XNOR2_X1 U475 ( .A(n413), .B(n412), .ZN(n414) );
  XOR2_X1 U476 ( .A(n415), .B(n414), .Z(n555) );
  XNOR2_X1 U477 ( .A(KEYINPUT36), .B(n562), .ZN(n580) );
  NAND2_X1 U478 ( .A1(n416), .A2(n580), .ZN(n417) );
  XNOR2_X1 U479 ( .A(KEYINPUT37), .B(n417), .ZN(n512) );
  XOR2_X1 U480 ( .A(G204GAT), .B(KEYINPUT75), .Z(n419) );
  XNOR2_X1 U481 ( .A(KEYINPUT74), .B(KEYINPUT73), .ZN(n418) );
  XNOR2_X1 U482 ( .A(n419), .B(n418), .ZN(n420) );
  XOR2_X1 U483 ( .A(n421), .B(n420), .Z(n425) );
  XNOR2_X1 U484 ( .A(n423), .B(n422), .ZN(n424) );
  XNOR2_X1 U485 ( .A(n425), .B(n424), .ZN(n434) );
  XOR2_X1 U486 ( .A(KEYINPUT33), .B(KEYINPUT32), .Z(n427) );
  NAND2_X1 U487 ( .A1(G230GAT), .A2(G233GAT), .ZN(n426) );
  XNOR2_X1 U488 ( .A(n427), .B(n426), .ZN(n428) );
  XOR2_X1 U489 ( .A(n428), .B(KEYINPUT31), .Z(n432) );
  XNOR2_X1 U490 ( .A(n430), .B(n429), .ZN(n431) );
  XNOR2_X1 U491 ( .A(n432), .B(n431), .ZN(n433) );
  XOR2_X1 U492 ( .A(n434), .B(n433), .Z(n574) );
  XOR2_X1 U493 ( .A(KEYINPUT66), .B(KEYINPUT67), .Z(n436) );
  XNOR2_X1 U494 ( .A(G197GAT), .B(G113GAT), .ZN(n435) );
  XNOR2_X1 U495 ( .A(n436), .B(n435), .ZN(n451) );
  XOR2_X1 U496 ( .A(KEYINPUT30), .B(G15GAT), .Z(n438) );
  XNOR2_X1 U497 ( .A(G50GAT), .B(G36GAT), .ZN(n437) );
  XNOR2_X1 U498 ( .A(n438), .B(n437), .ZN(n442) );
  XOR2_X1 U499 ( .A(KEYINPUT29), .B(G1GAT), .Z(n440) );
  XNOR2_X1 U500 ( .A(KEYINPUT72), .B(KEYINPUT69), .ZN(n439) );
  XNOR2_X1 U501 ( .A(n440), .B(n439), .ZN(n441) );
  XOR2_X1 U502 ( .A(n442), .B(n441), .Z(n449) );
  XOR2_X1 U503 ( .A(n443), .B(KEYINPUT68), .Z(n445) );
  NAND2_X1 U504 ( .A1(G229GAT), .A2(G233GAT), .ZN(n444) );
  XNOR2_X1 U505 ( .A(n445), .B(n444), .ZN(n446) );
  XNOR2_X1 U506 ( .A(n447), .B(n446), .ZN(n448) );
  XNOR2_X1 U507 ( .A(n449), .B(n448), .ZN(n450) );
  XOR2_X1 U508 ( .A(n451), .B(n450), .Z(n452) );
  XNOR2_X1 U509 ( .A(n453), .B(n452), .ZN(n570) );
  NOR2_X1 U510 ( .A1(n574), .A2(n570), .ZN(n484) );
  NAND2_X1 U511 ( .A1(n512), .A2(n484), .ZN(n454) );
  NAND2_X1 U512 ( .A1(n496), .A2(n527), .ZN(n456) );
  XNOR2_X1 U513 ( .A(KEYINPUT122), .B(KEYINPUT55), .ZN(n474) );
  INV_X1 U514 ( .A(KEYINPUT54), .ZN(n470) );
  XOR2_X1 U515 ( .A(KEYINPUT47), .B(KEYINPUT111), .Z(n461) );
  XNOR2_X1 U516 ( .A(KEYINPUT41), .B(n574), .ZN(n548) );
  NOR2_X1 U517 ( .A1(n570), .A2(n548), .ZN(n457) );
  XNOR2_X1 U518 ( .A(n457), .B(KEYINPUT46), .ZN(n458) );
  NOR2_X1 U519 ( .A1(n577), .A2(n458), .ZN(n459) );
  NAND2_X1 U520 ( .A1(n459), .A2(n555), .ZN(n460) );
  XNOR2_X1 U521 ( .A(n461), .B(n460), .ZN(n467) );
  NAND2_X1 U522 ( .A1(n577), .A2(n580), .ZN(n463) );
  XOR2_X1 U523 ( .A(KEYINPUT45), .B(KEYINPUT112), .Z(n462) );
  NAND2_X1 U524 ( .A1(n464), .A2(n570), .ZN(n465) );
  NOR2_X1 U525 ( .A1(n574), .A2(n465), .ZN(n466) );
  NOR2_X1 U526 ( .A1(n467), .A2(n466), .ZN(n468) );
  XNOR2_X1 U527 ( .A(n468), .B(KEYINPUT48), .ZN(n526) );
  NOR2_X1 U528 ( .A1(n515), .A2(n526), .ZN(n469) );
  XNOR2_X1 U529 ( .A(n470), .B(n469), .ZN(n471) );
  NOR2_X1 U530 ( .A1(n471), .A2(n501), .ZN(n569) );
  AND2_X1 U531 ( .A1(n569), .A2(n472), .ZN(n473) );
  XNOR2_X1 U532 ( .A(n474), .B(n473), .ZN(n475) );
  INV_X1 U533 ( .A(n548), .ZN(n533) );
  NAND2_X1 U534 ( .A1(n563), .A2(n533), .ZN(n479) );
  XOR2_X1 U535 ( .A(G176GAT), .B(KEYINPUT57), .Z(n477) );
  XOR2_X1 U536 ( .A(KEYINPUT123), .B(KEYINPUT56), .Z(n476) );
  INV_X1 U537 ( .A(n501), .ZN(n513) );
  INV_X1 U538 ( .A(n577), .ZN(n551) );
  NOR2_X1 U539 ( .A1(n562), .A2(n551), .ZN(n480) );
  XOR2_X1 U540 ( .A(KEYINPUT80), .B(n480), .Z(n481) );
  XNOR2_X1 U541 ( .A(KEYINPUT16), .B(n481), .ZN(n482) );
  NOR2_X1 U542 ( .A1(n483), .A2(n482), .ZN(n499) );
  NAND2_X1 U543 ( .A1(n484), .A2(n499), .ZN(n490) );
  NOR2_X1 U544 ( .A1(n513), .A2(n490), .ZN(n485) );
  XOR2_X1 U545 ( .A(G1GAT), .B(n485), .Z(n486) );
  XNOR2_X1 U546 ( .A(KEYINPUT34), .B(n486), .ZN(G1324GAT) );
  NOR2_X1 U547 ( .A1(n515), .A2(n490), .ZN(n487) );
  XOR2_X1 U548 ( .A(G8GAT), .B(n487), .Z(G1325GAT) );
  NOR2_X1 U549 ( .A1(n517), .A2(n490), .ZN(n489) );
  XNOR2_X1 U550 ( .A(G15GAT), .B(KEYINPUT35), .ZN(n488) );
  XNOR2_X1 U551 ( .A(n489), .B(n488), .ZN(G1326GAT) );
  INV_X1 U552 ( .A(n530), .ZN(n521) );
  NOR2_X1 U553 ( .A1(n521), .A2(n490), .ZN(n491) );
  XOR2_X1 U554 ( .A(G22GAT), .B(n491), .Z(G1327GAT) );
  NAND2_X1 U555 ( .A1(n501), .A2(n496), .ZN(n493) );
  XOR2_X1 U556 ( .A(G29GAT), .B(KEYINPUT39), .Z(n492) );
  XNOR2_X1 U557 ( .A(n493), .B(n492), .ZN(G1328GAT) );
  XOR2_X1 U558 ( .A(G36GAT), .B(KEYINPUT105), .Z(n495) );
  NAND2_X1 U559 ( .A1(n496), .A2(n504), .ZN(n494) );
  XNOR2_X1 U560 ( .A(n495), .B(n494), .ZN(G1329GAT) );
  NAND2_X1 U561 ( .A1(n496), .A2(n530), .ZN(n497) );
  XNOR2_X1 U562 ( .A(n497), .B(KEYINPUT106), .ZN(n498) );
  XNOR2_X1 U563 ( .A(G50GAT), .B(n498), .ZN(G1331GAT) );
  XNOR2_X1 U564 ( .A(G57GAT), .B(KEYINPUT42), .ZN(n503) );
  INV_X1 U565 ( .A(n570), .ZN(n559) );
  NOR2_X1 U566 ( .A1(n559), .A2(n548), .ZN(n511) );
  NAND2_X1 U567 ( .A1(n511), .A2(n499), .ZN(n500) );
  XNOR2_X1 U568 ( .A(KEYINPUT107), .B(n500), .ZN(n507) );
  NAND2_X1 U569 ( .A1(n501), .A2(n507), .ZN(n502) );
  XNOR2_X1 U570 ( .A(n503), .B(n502), .ZN(G1332GAT) );
  NAND2_X1 U571 ( .A1(n504), .A2(n507), .ZN(n505) );
  XNOR2_X1 U572 ( .A(n505), .B(G64GAT), .ZN(G1333GAT) );
  NAND2_X1 U573 ( .A1(n507), .A2(n527), .ZN(n506) );
  XNOR2_X1 U574 ( .A(n506), .B(G71GAT), .ZN(G1334GAT) );
  XOR2_X1 U575 ( .A(KEYINPUT108), .B(KEYINPUT43), .Z(n509) );
  NAND2_X1 U576 ( .A1(n507), .A2(n530), .ZN(n508) );
  XNOR2_X1 U577 ( .A(n509), .B(n508), .ZN(n510) );
  XNOR2_X1 U578 ( .A(G78GAT), .B(n510), .ZN(G1335GAT) );
  NAND2_X1 U579 ( .A1(n512), .A2(n511), .ZN(n520) );
  NOR2_X1 U580 ( .A1(n513), .A2(n520), .ZN(n514) );
  XOR2_X1 U581 ( .A(G85GAT), .B(n514), .Z(G1336GAT) );
  NOR2_X1 U582 ( .A1(n515), .A2(n520), .ZN(n516) );
  XOR2_X1 U583 ( .A(G92GAT), .B(n516), .Z(G1337GAT) );
  NOR2_X1 U584 ( .A1(n517), .A2(n520), .ZN(n519) );
  XNOR2_X1 U585 ( .A(G99GAT), .B(KEYINPUT109), .ZN(n518) );
  XNOR2_X1 U586 ( .A(n519), .B(n518), .ZN(G1338GAT) );
  NOR2_X1 U587 ( .A1(n521), .A2(n520), .ZN(n523) );
  XNOR2_X1 U588 ( .A(KEYINPUT44), .B(KEYINPUT110), .ZN(n522) );
  XNOR2_X1 U589 ( .A(n523), .B(n522), .ZN(n524) );
  XOR2_X1 U590 ( .A(G106GAT), .B(n524), .Z(G1339GAT) );
  NOR2_X1 U591 ( .A1(n526), .A2(n525), .ZN(n543) );
  NAND2_X1 U592 ( .A1(n527), .A2(n543), .ZN(n528) );
  XOR2_X1 U593 ( .A(KEYINPUT113), .B(n528), .Z(n529) );
  NOR2_X1 U594 ( .A1(n530), .A2(n529), .ZN(n539) );
  NAND2_X1 U595 ( .A1(n539), .A2(n559), .ZN(n531) );
  XNOR2_X1 U596 ( .A(n531), .B(KEYINPUT114), .ZN(n532) );
  XNOR2_X1 U597 ( .A(G113GAT), .B(n532), .ZN(G1340GAT) );
  XOR2_X1 U598 ( .A(G120GAT), .B(KEYINPUT49), .Z(n535) );
  NAND2_X1 U599 ( .A1(n539), .A2(n533), .ZN(n534) );
  XNOR2_X1 U600 ( .A(n535), .B(n534), .ZN(G1341GAT) );
  XOR2_X1 U601 ( .A(KEYINPUT115), .B(KEYINPUT50), .Z(n537) );
  NAND2_X1 U602 ( .A1(n539), .A2(n577), .ZN(n536) );
  XNOR2_X1 U603 ( .A(n537), .B(n536), .ZN(n538) );
  XNOR2_X1 U604 ( .A(G127GAT), .B(n538), .ZN(G1342GAT) );
  XOR2_X1 U605 ( .A(KEYINPUT116), .B(KEYINPUT51), .Z(n541) );
  NAND2_X1 U606 ( .A1(n539), .A2(n562), .ZN(n540) );
  XNOR2_X1 U607 ( .A(n541), .B(n540), .ZN(n542) );
  XNOR2_X1 U608 ( .A(G134GAT), .B(n542), .ZN(G1343GAT) );
  NAND2_X1 U609 ( .A1(n543), .A2(n568), .ZN(n554) );
  NOR2_X1 U610 ( .A1(n570), .A2(n554), .ZN(n545) );
  XNOR2_X1 U611 ( .A(G141GAT), .B(KEYINPUT117), .ZN(n544) );
  XNOR2_X1 U612 ( .A(n545), .B(n544), .ZN(G1344GAT) );
  XOR2_X1 U613 ( .A(KEYINPUT52), .B(KEYINPUT118), .Z(n547) );
  XNOR2_X1 U614 ( .A(G148GAT), .B(KEYINPUT53), .ZN(n546) );
  XNOR2_X1 U615 ( .A(n547), .B(n546), .ZN(n550) );
  NOR2_X1 U616 ( .A1(n548), .A2(n554), .ZN(n549) );
  XOR2_X1 U617 ( .A(n550), .B(n549), .Z(G1345GAT) );
  NOR2_X1 U618 ( .A1(n551), .A2(n554), .ZN(n553) );
  XNOR2_X1 U619 ( .A(G155GAT), .B(KEYINPUT119), .ZN(n552) );
  XNOR2_X1 U620 ( .A(n553), .B(n552), .ZN(G1346GAT) );
  NOR2_X1 U621 ( .A1(n555), .A2(n554), .ZN(n557) );
  XNOR2_X1 U622 ( .A(KEYINPUT120), .B(KEYINPUT121), .ZN(n556) );
  XNOR2_X1 U623 ( .A(n557), .B(n556), .ZN(n558) );
  XNOR2_X1 U624 ( .A(G162GAT), .B(n558), .ZN(G1347GAT) );
  NAND2_X1 U625 ( .A1(n563), .A2(n559), .ZN(n560) );
  XNOR2_X1 U626 ( .A(n560), .B(G169GAT), .ZN(G1348GAT) );
  NAND2_X1 U627 ( .A1(n563), .A2(n577), .ZN(n561) );
  XNOR2_X1 U628 ( .A(n561), .B(G183GAT), .ZN(G1350GAT) );
  NAND2_X1 U629 ( .A1(n563), .A2(n562), .ZN(n564) );
  XNOR2_X1 U630 ( .A(n564), .B(KEYINPUT58), .ZN(n565) );
  XNOR2_X1 U631 ( .A(G190GAT), .B(n565), .ZN(G1351GAT) );
  XOR2_X1 U632 ( .A(KEYINPUT124), .B(KEYINPUT59), .Z(n567) );
  XNOR2_X1 U633 ( .A(G197GAT), .B(KEYINPUT60), .ZN(n566) );
  XNOR2_X1 U634 ( .A(n567), .B(n566), .ZN(n572) );
  NAND2_X1 U635 ( .A1(n569), .A2(n568), .ZN(n573) );
  NOR2_X1 U636 ( .A1(n570), .A2(n573), .ZN(n571) );
  XOR2_X1 U637 ( .A(n572), .B(n571), .Z(G1352GAT) );
  XOR2_X1 U638 ( .A(G204GAT), .B(KEYINPUT61), .Z(n576) );
  INV_X1 U639 ( .A(n573), .ZN(n581) );
  NAND2_X1 U640 ( .A1(n581), .A2(n574), .ZN(n575) );
  XNOR2_X1 U641 ( .A(n576), .B(n575), .ZN(G1353GAT) );
  XOR2_X1 U642 ( .A(G211GAT), .B(KEYINPUT125), .Z(n579) );
  NAND2_X1 U643 ( .A1(n581), .A2(n577), .ZN(n578) );
  XNOR2_X1 U644 ( .A(n579), .B(n578), .ZN(G1354GAT) );
  XNOR2_X1 U645 ( .A(G218GAT), .B(KEYINPUT126), .ZN(n585) );
  XOR2_X1 U646 ( .A(KEYINPUT127), .B(KEYINPUT62), .Z(n583) );
  NAND2_X1 U647 ( .A1(n581), .A2(n580), .ZN(n582) );
  XNOR2_X1 U648 ( .A(n583), .B(n582), .ZN(n584) );
  XNOR2_X1 U649 ( .A(n585), .B(n584), .ZN(G1355GAT) );
endmodule

