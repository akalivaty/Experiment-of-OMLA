//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 1 0 1 0 1 1 1 1 1 0 0 0 1 0 1 0 0 1 1 0 0 1 1 1 1 0 0 0 1 1 0 0 0 1 1 1 1 1 1 1 1 1 1 0 0 1 1 1 1 0 0 0 1 0 1 1 0 1 0 0 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:33:04 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n455, new_n456, new_n457,
    new_n458, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n488, new_n489,
    new_n490, new_n491, new_n492, new_n493, new_n494, new_n495, new_n496,
    new_n497, new_n498, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n508, new_n509, new_n510, new_n511, new_n512,
    new_n513, new_n514, new_n515, new_n516, new_n517, new_n520, new_n521,
    new_n522, new_n523, new_n524, new_n525, new_n526, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n540, new_n541, new_n542, new_n544, new_n545, new_n546, new_n547,
    new_n548, new_n549, new_n550, new_n551, new_n552, new_n553, new_n554,
    new_n555, new_n556, new_n557, new_n558, new_n559, new_n560, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n570,
    new_n571, new_n572, new_n573, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n596, new_n597, new_n600, new_n602, new_n603, new_n605, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n653, new_n654, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n823, new_n824,
    new_n825, new_n826, new_n827, new_n828, new_n829, new_n830, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1090, new_n1091;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  XNOR2_X1  g009(.A(KEYINPUT64), .B(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G219), .A2(G220), .A3(G218), .A4(G221), .ZN(new_n450));
  XOR2_X1   g025(.A(new_n450), .B(KEYINPUT2), .Z(new_n451));
  NAND4_X1  g026(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n452));
  NOR2_X1   g027(.A1(new_n451), .A2(new_n452), .ZN(G325));
  INV_X1    g028(.A(G325), .ZN(G261));
  NAND2_X1  g029(.A1(new_n451), .A2(G2106), .ZN(new_n455));
  NAND2_X1  g030(.A1(new_n452), .A2(G567), .ZN(new_n456));
  XOR2_X1   g031(.A(new_n456), .B(KEYINPUT65), .Z(new_n457));
  NAND2_X1  g032(.A1(new_n455), .A2(new_n457), .ZN(new_n458));
  INV_X1    g033(.A(new_n458), .ZN(G319));
  AND2_X1   g034(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n460));
  NOR2_X1   g035(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n461));
  NOR2_X1   g036(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  INV_X1    g037(.A(new_n462), .ZN(new_n463));
  AND2_X1   g038(.A1(new_n463), .A2(G125), .ZN(new_n464));
  AND2_X1   g039(.A1(G113), .A2(G2104), .ZN(new_n465));
  OAI21_X1  g040(.A(G2105), .B1(new_n464), .B2(new_n465), .ZN(new_n466));
  NOR2_X1   g041(.A1(new_n462), .A2(G2105), .ZN(new_n467));
  INV_X1    g042(.A(G2104), .ZN(new_n468));
  NOR2_X1   g043(.A1(new_n468), .A2(G2105), .ZN(new_n469));
  AOI22_X1  g044(.A1(new_n467), .A2(G137), .B1(G101), .B2(new_n469), .ZN(new_n470));
  AND2_X1   g045(.A1(new_n466), .A2(new_n470), .ZN(G160));
  OAI21_X1  g046(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n472));
  INV_X1    g047(.A(G112), .ZN(new_n473));
  AOI21_X1  g048(.A(new_n472), .B1(new_n473), .B2(G2105), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n467), .A2(G136), .ZN(new_n475));
  XOR2_X1   g050(.A(new_n475), .B(KEYINPUT66), .Z(new_n476));
  INV_X1    g051(.A(G2105), .ZN(new_n477));
  NOR2_X1   g052(.A1(new_n462), .A2(new_n477), .ZN(new_n478));
  AOI211_X1 g053(.A(new_n474), .B(new_n476), .C1(G124), .C2(new_n478), .ZN(G162));
  NAND2_X1  g054(.A1(new_n467), .A2(G138), .ZN(new_n480));
  XNOR2_X1  g055(.A(new_n480), .B(KEYINPUT4), .ZN(new_n481));
  OAI21_X1  g056(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n482));
  INV_X1    g057(.A(G114), .ZN(new_n483));
  AOI21_X1  g058(.A(new_n482), .B1(new_n483), .B2(G2105), .ZN(new_n484));
  AOI21_X1  g059(.A(new_n484), .B1(new_n478), .B2(G126), .ZN(new_n485));
  NAND2_X1  g060(.A1(new_n481), .A2(new_n485), .ZN(new_n486));
  INV_X1    g061(.A(new_n486), .ZN(G164));
  XNOR2_X1  g062(.A(KEYINPUT5), .B(G543), .ZN(new_n488));
  AOI22_X1  g063(.A1(new_n488), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n489));
  INV_X1    g064(.A(new_n489), .ZN(new_n490));
  AND2_X1   g065(.A1(KEYINPUT6), .A2(G651), .ZN(new_n491));
  NOR2_X1   g066(.A1(KEYINPUT6), .A2(G651), .ZN(new_n492));
  NOR2_X1   g067(.A1(new_n491), .A2(new_n492), .ZN(new_n493));
  INV_X1    g068(.A(G543), .ZN(new_n494));
  NOR2_X1   g069(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  AOI22_X1  g070(.A1(new_n490), .A2(G651), .B1(G50), .B2(new_n495), .ZN(new_n496));
  INV_X1    g071(.A(G88), .ZN(new_n497));
  INV_X1    g072(.A(KEYINPUT67), .ZN(new_n498));
  AND2_X1   g073(.A1(KEYINPUT5), .A2(G543), .ZN(new_n499));
  NOR2_X1   g074(.A1(KEYINPUT5), .A2(G543), .ZN(new_n500));
  NOR2_X1   g075(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  OAI21_X1  g076(.A(new_n498), .B1(new_n501), .B2(new_n493), .ZN(new_n502));
  XNOR2_X1  g077(.A(KEYINPUT6), .B(G651), .ZN(new_n503));
  NAND3_X1  g078(.A1(new_n488), .A2(new_n503), .A3(KEYINPUT67), .ZN(new_n504));
  NAND2_X1  g079(.A1(new_n502), .A2(new_n504), .ZN(new_n505));
  OAI21_X1  g080(.A(new_n496), .B1(new_n497), .B2(new_n505), .ZN(G303));
  INV_X1    g081(.A(G303), .ZN(G166));
  AND2_X1   g082(.A1(G76), .A2(G543), .ZN(new_n508));
  AOI21_X1  g083(.A(KEYINPUT7), .B1(new_n508), .B2(G651), .ZN(new_n509));
  INV_X1    g084(.A(G651), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n488), .A2(G63), .ZN(new_n511));
  NAND2_X1  g086(.A1(new_n508), .A2(KEYINPUT7), .ZN(new_n512));
  AOI21_X1  g087(.A(new_n510), .B1(new_n511), .B2(new_n512), .ZN(new_n513));
  XNOR2_X1  g088(.A(KEYINPUT68), .B(G51), .ZN(new_n514));
  AOI211_X1 g089(.A(new_n509), .B(new_n513), .C1(new_n495), .C2(new_n514), .ZN(new_n515));
  INV_X1    g090(.A(new_n505), .ZN(new_n516));
  NAND2_X1  g091(.A1(new_n516), .A2(G89), .ZN(new_n517));
  NAND2_X1  g092(.A1(new_n515), .A2(new_n517), .ZN(G286));
  INV_X1    g093(.A(G286), .ZN(G168));
  NAND2_X1  g094(.A1(new_n516), .A2(G90), .ZN(new_n520));
  NAND2_X1  g095(.A1(G77), .A2(G543), .ZN(new_n521));
  INV_X1    g096(.A(G64), .ZN(new_n522));
  OAI21_X1  g097(.A(new_n521), .B1(new_n501), .B2(new_n522), .ZN(new_n523));
  AOI21_X1  g098(.A(new_n510), .B1(new_n523), .B2(KEYINPUT69), .ZN(new_n524));
  OAI21_X1  g099(.A(new_n524), .B1(KEYINPUT69), .B2(new_n523), .ZN(new_n525));
  NAND2_X1  g100(.A1(new_n495), .A2(G52), .ZN(new_n526));
  NAND3_X1  g101(.A1(new_n520), .A2(new_n525), .A3(new_n526), .ZN(G301));
  INV_X1    g102(.A(G301), .ZN(G171));
  NAND2_X1  g103(.A1(new_n495), .A2(G43), .ZN(new_n529));
  INV_X1    g104(.A(G81), .ZN(new_n530));
  OAI21_X1  g105(.A(new_n529), .B1(new_n505), .B2(new_n530), .ZN(new_n531));
  INV_X1    g106(.A(KEYINPUT70), .ZN(new_n532));
  XNOR2_X1  g107(.A(new_n531), .B(new_n532), .ZN(new_n533));
  AOI22_X1  g108(.A1(new_n488), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n534));
  OR2_X1    g109(.A1(new_n534), .A2(new_n510), .ZN(new_n535));
  NAND2_X1  g110(.A1(new_n533), .A2(new_n535), .ZN(new_n536));
  INV_X1    g111(.A(new_n536), .ZN(new_n537));
  NAND2_X1  g112(.A1(new_n537), .A2(G860), .ZN(G153));
  NAND4_X1  g113(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g114(.A1(G1), .A2(G3), .ZN(new_n540));
  XNOR2_X1  g115(.A(new_n540), .B(KEYINPUT8), .ZN(new_n541));
  NAND4_X1  g116(.A1(G319), .A2(G483), .A3(G661), .A4(new_n541), .ZN(new_n542));
  XNOR2_X1  g117(.A(new_n542), .B(KEYINPUT71), .ZN(G188));
  AND3_X1   g118(.A1(new_n488), .A2(new_n503), .A3(KEYINPUT67), .ZN(new_n544));
  AOI21_X1  g119(.A(KEYINPUT67), .B1(new_n488), .B2(new_n503), .ZN(new_n545));
  OAI21_X1  g120(.A(KEYINPUT73), .B1(new_n544), .B2(new_n545), .ZN(new_n546));
  INV_X1    g121(.A(KEYINPUT73), .ZN(new_n547));
  NAND3_X1  g122(.A1(new_n502), .A2(new_n547), .A3(new_n504), .ZN(new_n548));
  NAND3_X1  g123(.A1(new_n546), .A2(G91), .A3(new_n548), .ZN(new_n549));
  INV_X1    g124(.A(KEYINPUT9), .ZN(new_n550));
  NAND2_X1  g125(.A1(new_n503), .A2(G543), .ZN(new_n551));
  INV_X1    g126(.A(G53), .ZN(new_n552));
  OAI211_X1 g127(.A(KEYINPUT72), .B(new_n550), .C1(new_n551), .C2(new_n552), .ZN(new_n553));
  XNOR2_X1  g128(.A(KEYINPUT72), .B(KEYINPUT9), .ZN(new_n554));
  NAND3_X1  g129(.A1(new_n495), .A2(G53), .A3(new_n554), .ZN(new_n555));
  NAND2_X1  g130(.A1(G78), .A2(G543), .ZN(new_n556));
  INV_X1    g131(.A(G65), .ZN(new_n557));
  OAI21_X1  g132(.A(new_n556), .B1(new_n501), .B2(new_n557), .ZN(new_n558));
  NAND2_X1  g133(.A1(new_n558), .A2(G651), .ZN(new_n559));
  AND3_X1   g134(.A1(new_n553), .A2(new_n555), .A3(new_n559), .ZN(new_n560));
  NAND2_X1  g135(.A1(new_n549), .A2(new_n560), .ZN(G299));
  AND2_X1   g136(.A1(new_n546), .A2(new_n548), .ZN(new_n562));
  NAND2_X1  g137(.A1(new_n562), .A2(G87), .ZN(new_n563));
  INV_X1    g138(.A(G49), .ZN(new_n564));
  OR3_X1    g139(.A1(new_n551), .A2(KEYINPUT74), .A3(new_n564), .ZN(new_n565));
  OAI21_X1  g140(.A(KEYINPUT74), .B1(new_n551), .B2(new_n564), .ZN(new_n566));
  OR2_X1    g141(.A1(new_n488), .A2(G74), .ZN(new_n567));
  AOI22_X1  g142(.A1(new_n565), .A2(new_n566), .B1(G651), .B2(new_n567), .ZN(new_n568));
  NAND2_X1  g143(.A1(new_n563), .A2(new_n568), .ZN(G288));
  NAND2_X1  g144(.A1(new_n562), .A2(G86), .ZN(new_n570));
  AOI22_X1  g145(.A1(new_n488), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n571));
  INV_X1    g146(.A(new_n571), .ZN(new_n572));
  AOI22_X1  g147(.A1(new_n572), .A2(G651), .B1(G48), .B2(new_n495), .ZN(new_n573));
  NAND2_X1  g148(.A1(new_n570), .A2(new_n573), .ZN(G305));
  NAND2_X1  g149(.A1(new_n495), .A2(G47), .ZN(new_n575));
  AOI22_X1  g150(.A1(new_n488), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n576));
  INV_X1    g151(.A(G85), .ZN(new_n577));
  OAI221_X1 g152(.A(new_n575), .B1(new_n510), .B2(new_n576), .C1(new_n505), .C2(new_n577), .ZN(new_n578));
  XNOR2_X1  g153(.A(new_n578), .B(KEYINPUT75), .ZN(new_n579));
  INV_X1    g154(.A(new_n579), .ZN(G290));
  INV_X1    g155(.A(G868), .ZN(new_n581));
  NOR2_X1   g156(.A1(G301), .A2(new_n581), .ZN(new_n582));
  NAND3_X1  g157(.A1(new_n546), .A2(G92), .A3(new_n548), .ZN(new_n583));
  INV_X1    g158(.A(KEYINPUT10), .ZN(new_n584));
  NAND2_X1  g159(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  NAND4_X1  g160(.A1(new_n546), .A2(KEYINPUT10), .A3(G92), .A4(new_n548), .ZN(new_n586));
  NAND2_X1  g161(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  AOI22_X1  g162(.A1(new_n488), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n588));
  INV_X1    g163(.A(G54), .ZN(new_n589));
  OAI22_X1  g164(.A1(new_n588), .A2(new_n510), .B1(new_n589), .B2(new_n551), .ZN(new_n590));
  INV_X1    g165(.A(new_n590), .ZN(new_n591));
  NAND2_X1  g166(.A1(new_n587), .A2(new_n591), .ZN(new_n592));
  XNOR2_X1  g167(.A(new_n592), .B(KEYINPUT76), .ZN(new_n593));
  AOI21_X1  g168(.A(new_n582), .B1(new_n593), .B2(new_n581), .ZN(G284));
  XOR2_X1   g169(.A(G284), .B(KEYINPUT77), .Z(G321));
  NOR2_X1   g170(.A1(G286), .A2(new_n581), .ZN(new_n596));
  XOR2_X1   g171(.A(G299), .B(KEYINPUT78), .Z(new_n597));
  AOI21_X1  g172(.A(new_n596), .B1(new_n597), .B2(new_n581), .ZN(G297));
  AOI21_X1  g173(.A(new_n596), .B1(new_n597), .B2(new_n581), .ZN(G280));
  INV_X1    g174(.A(G559), .ZN(new_n600));
  OAI21_X1  g175(.A(new_n593), .B1(new_n600), .B2(G860), .ZN(G148));
  NAND2_X1  g176(.A1(new_n536), .A2(new_n581), .ZN(new_n602));
  AND2_X1   g177(.A1(new_n593), .A2(new_n600), .ZN(new_n603));
  OAI21_X1  g178(.A(new_n602), .B1(new_n603), .B2(new_n581), .ZN(G323));
  XOR2_X1   g179(.A(KEYINPUT79), .B(KEYINPUT11), .Z(new_n605));
  XNOR2_X1  g180(.A(G323), .B(new_n605), .ZN(G282));
  NAND2_X1  g181(.A1(new_n463), .A2(new_n469), .ZN(new_n607));
  XOR2_X1   g182(.A(KEYINPUT80), .B(KEYINPUT12), .Z(new_n608));
  XNOR2_X1  g183(.A(new_n607), .B(new_n608), .ZN(new_n609));
  XOR2_X1   g184(.A(KEYINPUT81), .B(KEYINPUT13), .Z(new_n610));
  XNOR2_X1  g185(.A(new_n609), .B(new_n610), .ZN(new_n611));
  INV_X1    g186(.A(new_n611), .ZN(new_n612));
  XNOR2_X1  g187(.A(KEYINPUT82), .B(G2100), .ZN(new_n613));
  OR2_X1    g188(.A1(new_n612), .A2(new_n613), .ZN(new_n614));
  NAND2_X1  g189(.A1(new_n612), .A2(new_n613), .ZN(new_n615));
  NAND2_X1  g190(.A1(new_n467), .A2(G135), .ZN(new_n616));
  NAND2_X1  g191(.A1(new_n478), .A2(G123), .ZN(new_n617));
  OR2_X1    g192(.A1(G99), .A2(G2105), .ZN(new_n618));
  OAI211_X1 g193(.A(new_n618), .B(G2104), .C1(G111), .C2(new_n477), .ZN(new_n619));
  NAND3_X1  g194(.A1(new_n616), .A2(new_n617), .A3(new_n619), .ZN(new_n620));
  XOR2_X1   g195(.A(new_n620), .B(G2096), .Z(new_n621));
  NAND3_X1  g196(.A1(new_n614), .A2(new_n615), .A3(new_n621), .ZN(G156));
  XOR2_X1   g197(.A(G2451), .B(G2454), .Z(new_n623));
  XNOR2_X1  g198(.A(new_n623), .B(KEYINPUT16), .ZN(new_n624));
  XNOR2_X1  g199(.A(G1341), .B(G1348), .ZN(new_n625));
  XNOR2_X1  g200(.A(new_n625), .B(KEYINPUT83), .ZN(new_n626));
  XNOR2_X1  g201(.A(new_n624), .B(new_n626), .ZN(new_n627));
  INV_X1    g202(.A(KEYINPUT14), .ZN(new_n628));
  XNOR2_X1  g203(.A(G2427), .B(G2438), .ZN(new_n629));
  XNOR2_X1  g204(.A(new_n629), .B(G2430), .ZN(new_n630));
  XNOR2_X1  g205(.A(KEYINPUT15), .B(G2435), .ZN(new_n631));
  AOI21_X1  g206(.A(new_n628), .B1(new_n630), .B2(new_n631), .ZN(new_n632));
  OAI21_X1  g207(.A(new_n632), .B1(new_n631), .B2(new_n630), .ZN(new_n633));
  XOR2_X1   g208(.A(new_n627), .B(new_n633), .Z(new_n634));
  INV_X1    g209(.A(new_n634), .ZN(new_n635));
  XNOR2_X1  g210(.A(G2443), .B(G2446), .ZN(new_n636));
  INV_X1    g211(.A(new_n636), .ZN(new_n637));
  OAI21_X1  g212(.A(G14), .B1(new_n635), .B2(new_n637), .ZN(new_n638));
  AOI21_X1  g213(.A(new_n638), .B1(new_n637), .B2(new_n635), .ZN(G401));
  XOR2_X1   g214(.A(G2072), .B(G2078), .Z(new_n640));
  XOR2_X1   g215(.A(G2084), .B(G2090), .Z(new_n641));
  XNOR2_X1  g216(.A(G2067), .B(G2678), .ZN(new_n642));
  NAND2_X1  g217(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  AOI21_X1  g218(.A(new_n640), .B1(new_n643), .B2(KEYINPUT18), .ZN(new_n644));
  XNOR2_X1  g219(.A(new_n644), .B(KEYINPUT84), .ZN(new_n645));
  XNOR2_X1  g220(.A(new_n645), .B(G2100), .ZN(new_n646));
  INV_X1    g221(.A(KEYINPUT18), .ZN(new_n647));
  NAND2_X1  g222(.A1(new_n643), .A2(KEYINPUT17), .ZN(new_n648));
  NOR2_X1   g223(.A1(new_n641), .A2(new_n642), .ZN(new_n649));
  OAI21_X1  g224(.A(new_n647), .B1(new_n648), .B2(new_n649), .ZN(new_n650));
  XNOR2_X1  g225(.A(new_n650), .B(G2096), .ZN(new_n651));
  XNOR2_X1  g226(.A(new_n646), .B(new_n651), .ZN(G227));
  XOR2_X1   g227(.A(G1971), .B(G1976), .Z(new_n653));
  XNOR2_X1  g228(.A(new_n653), .B(KEYINPUT19), .ZN(new_n654));
  XNOR2_X1  g229(.A(G1956), .B(G2474), .ZN(new_n655));
  XNOR2_X1  g230(.A(G1961), .B(G1966), .ZN(new_n656));
  NOR2_X1   g231(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  NAND2_X1  g232(.A1(new_n654), .A2(new_n657), .ZN(new_n658));
  XOR2_X1   g233(.A(new_n658), .B(KEYINPUT20), .Z(new_n659));
  AND2_X1   g234(.A1(new_n655), .A2(new_n656), .ZN(new_n660));
  NAND2_X1  g235(.A1(new_n654), .A2(new_n660), .ZN(new_n661));
  XNOR2_X1  g236(.A(new_n661), .B(KEYINPUT85), .ZN(new_n662));
  NOR3_X1   g237(.A1(new_n654), .A2(new_n657), .A3(new_n660), .ZN(new_n663));
  NOR3_X1   g238(.A1(new_n659), .A2(new_n662), .A3(new_n663), .ZN(new_n664));
  XNOR2_X1  g239(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n665));
  XOR2_X1   g240(.A(new_n664), .B(new_n665), .Z(new_n666));
  XNOR2_X1  g241(.A(G1991), .B(G1996), .ZN(new_n667));
  XNOR2_X1  g242(.A(new_n667), .B(KEYINPUT86), .ZN(new_n668));
  XNOR2_X1  g243(.A(new_n666), .B(new_n668), .ZN(new_n669));
  INV_X1    g244(.A(new_n669), .ZN(new_n670));
  XNOR2_X1  g245(.A(G1981), .B(G1986), .ZN(new_n671));
  OR2_X1    g246(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  NAND2_X1  g247(.A1(new_n670), .A2(new_n671), .ZN(new_n673));
  NAND2_X1  g248(.A1(new_n672), .A2(new_n673), .ZN(G229));
  INV_X1    g249(.A(G16), .ZN(new_n675));
  NAND2_X1  g250(.A1(new_n675), .A2(G21), .ZN(new_n676));
  OAI21_X1  g251(.A(new_n676), .B1(G168), .B2(new_n675), .ZN(new_n677));
  XNOR2_X1  g252(.A(new_n677), .B(KEYINPUT94), .ZN(new_n678));
  NAND2_X1  g253(.A1(new_n678), .A2(G1966), .ZN(new_n679));
  XOR2_X1   g254(.A(new_n679), .B(KEYINPUT95), .Z(new_n680));
  AOI22_X1  g255(.A1(new_n467), .A2(G141), .B1(G105), .B2(new_n469), .ZN(new_n681));
  NAND2_X1  g256(.A1(new_n478), .A2(G129), .ZN(new_n682));
  NAND3_X1  g257(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n683));
  XOR2_X1   g258(.A(new_n683), .B(KEYINPUT26), .Z(new_n684));
  NAND3_X1  g259(.A1(new_n681), .A2(new_n682), .A3(new_n684), .ZN(new_n685));
  INV_X1    g260(.A(new_n685), .ZN(new_n686));
  INV_X1    g261(.A(G29), .ZN(new_n687));
  NOR2_X1   g262(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  AOI21_X1  g263(.A(new_n688), .B1(new_n687), .B2(G32), .ZN(new_n689));
  XOR2_X1   g264(.A(KEYINPUT27), .B(G1996), .Z(new_n690));
  XNOR2_X1  g265(.A(new_n690), .B(KEYINPUT93), .ZN(new_n691));
  NOR2_X1   g266(.A1(new_n689), .A2(new_n691), .ZN(new_n692));
  NOR2_X1   g267(.A1(G29), .A2(G33), .ZN(new_n693));
  XOR2_X1   g268(.A(new_n693), .B(KEYINPUT92), .Z(new_n694));
  AND2_X1   g269(.A1(new_n463), .A2(G127), .ZN(new_n695));
  AND2_X1   g270(.A1(G115), .A2(G2104), .ZN(new_n696));
  OAI21_X1  g271(.A(G2105), .B1(new_n695), .B2(new_n696), .ZN(new_n697));
  INV_X1    g272(.A(KEYINPUT25), .ZN(new_n698));
  NAND2_X1  g273(.A1(G103), .A2(G2104), .ZN(new_n699));
  OAI21_X1  g274(.A(new_n698), .B1(new_n699), .B2(G2105), .ZN(new_n700));
  NAND4_X1  g275(.A1(new_n477), .A2(KEYINPUT25), .A3(G103), .A4(G2104), .ZN(new_n701));
  AOI22_X1  g276(.A1(new_n467), .A2(G139), .B1(new_n700), .B2(new_n701), .ZN(new_n702));
  AND2_X1   g277(.A1(new_n697), .A2(new_n702), .ZN(new_n703));
  AOI21_X1  g278(.A(new_n694), .B1(new_n703), .B2(G29), .ZN(new_n704));
  AOI21_X1  g279(.A(new_n692), .B1(G2072), .B2(new_n704), .ZN(new_n705));
  OAI21_X1  g280(.A(new_n705), .B1(G2072), .B2(new_n704), .ZN(new_n706));
  INV_X1    g281(.A(KEYINPUT24), .ZN(new_n707));
  OAI21_X1  g282(.A(new_n687), .B1(new_n707), .B2(G34), .ZN(new_n708));
  AOI21_X1  g283(.A(new_n708), .B1(new_n707), .B2(G34), .ZN(new_n709));
  AOI21_X1  g284(.A(new_n709), .B1(G160), .B2(G29), .ZN(new_n710));
  NAND2_X1  g285(.A1(new_n710), .A2(G2084), .ZN(new_n711));
  OR2_X1    g286(.A1(KEYINPUT30), .A2(G28), .ZN(new_n712));
  NAND2_X1  g287(.A1(KEYINPUT30), .A2(G28), .ZN(new_n713));
  AOI21_X1  g288(.A(G29), .B1(new_n712), .B2(new_n713), .ZN(new_n714));
  XOR2_X1   g289(.A(KEYINPUT31), .B(G11), .Z(new_n715));
  NOR2_X1   g290(.A1(new_n714), .A2(new_n715), .ZN(new_n716));
  OAI211_X1 g291(.A(new_n711), .B(new_n716), .C1(new_n687), .C2(new_n620), .ZN(new_n717));
  NAND2_X1  g292(.A1(new_n689), .A2(new_n691), .ZN(new_n718));
  OAI21_X1  g293(.A(new_n718), .B1(G2084), .B2(new_n710), .ZN(new_n719));
  NOR3_X1   g294(.A1(new_n706), .A2(new_n717), .A3(new_n719), .ZN(new_n720));
  NOR2_X1   g295(.A1(G171), .A2(new_n675), .ZN(new_n721));
  AOI21_X1  g296(.A(new_n721), .B1(G5), .B2(new_n675), .ZN(new_n722));
  XNOR2_X1  g297(.A(KEYINPUT96), .B(G1961), .ZN(new_n723));
  OR2_X1    g298(.A1(new_n722), .A2(new_n723), .ZN(new_n724));
  NAND2_X1  g299(.A1(new_n687), .A2(G27), .ZN(new_n725));
  OAI21_X1  g300(.A(new_n725), .B1(G164), .B2(new_n687), .ZN(new_n726));
  XNOR2_X1  g301(.A(new_n726), .B(G2078), .ZN(new_n727));
  AOI21_X1  g302(.A(new_n727), .B1(new_n722), .B2(new_n723), .ZN(new_n728));
  OR2_X1    g303(.A1(new_n678), .A2(G1966), .ZN(new_n729));
  NAND4_X1  g304(.A1(new_n720), .A2(new_n724), .A3(new_n728), .A4(new_n729), .ZN(new_n730));
  NOR2_X1   g305(.A1(new_n680), .A2(new_n730), .ZN(new_n731));
  XOR2_X1   g306(.A(new_n731), .B(KEYINPUT97), .Z(new_n732));
  NAND2_X1  g307(.A1(new_n675), .A2(G19), .ZN(new_n733));
  XNOR2_X1  g308(.A(new_n733), .B(KEYINPUT90), .ZN(new_n734));
  OAI21_X1  g309(.A(new_n734), .B1(new_n537), .B2(new_n675), .ZN(new_n735));
  XOR2_X1   g310(.A(new_n735), .B(G1341), .Z(new_n736));
  NAND2_X1  g311(.A1(new_n687), .A2(G35), .ZN(new_n737));
  OAI21_X1  g312(.A(new_n737), .B1(G162), .B2(new_n687), .ZN(new_n738));
  XOR2_X1   g313(.A(KEYINPUT29), .B(G2090), .Z(new_n739));
  XNOR2_X1  g314(.A(new_n738), .B(new_n739), .ZN(new_n740));
  NAND2_X1  g315(.A1(new_n675), .A2(G20), .ZN(new_n741));
  XOR2_X1   g316(.A(new_n741), .B(KEYINPUT23), .Z(new_n742));
  AOI21_X1  g317(.A(new_n742), .B1(G299), .B2(G16), .ZN(new_n743));
  XNOR2_X1  g318(.A(new_n743), .B(G1956), .ZN(new_n744));
  NAND2_X1  g319(.A1(new_n687), .A2(G26), .ZN(new_n745));
  XOR2_X1   g320(.A(new_n745), .B(KEYINPUT28), .Z(new_n746));
  NAND2_X1  g321(.A1(new_n478), .A2(G128), .ZN(new_n747));
  XOR2_X1   g322(.A(new_n747), .B(KEYINPUT91), .Z(new_n748));
  NAND2_X1  g323(.A1(new_n467), .A2(G140), .ZN(new_n749));
  NOR2_X1   g324(.A1(new_n477), .A2(G116), .ZN(new_n750));
  OAI21_X1  g325(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n751));
  OAI211_X1 g326(.A(new_n748), .B(new_n749), .C1(new_n750), .C2(new_n751), .ZN(new_n752));
  AOI21_X1  g327(.A(new_n746), .B1(new_n752), .B2(G29), .ZN(new_n753));
  XNOR2_X1  g328(.A(new_n753), .B(G2067), .ZN(new_n754));
  NAND4_X1  g329(.A1(new_n736), .A2(new_n740), .A3(new_n744), .A4(new_n754), .ZN(new_n755));
  INV_X1    g330(.A(G1348), .ZN(new_n756));
  NOR2_X1   g331(.A1(new_n593), .A2(new_n675), .ZN(new_n757));
  AOI21_X1  g332(.A(new_n757), .B1(G4), .B2(new_n675), .ZN(new_n758));
  AOI21_X1  g333(.A(new_n755), .B1(new_n756), .B2(new_n758), .ZN(new_n759));
  OAI211_X1 g334(.A(new_n732), .B(new_n759), .C1(new_n756), .C2(new_n758), .ZN(new_n760));
  INV_X1    g335(.A(G288), .ZN(new_n761));
  NOR2_X1   g336(.A1(new_n761), .A2(new_n675), .ZN(new_n762));
  AOI21_X1  g337(.A(new_n762), .B1(new_n675), .B2(G23), .ZN(new_n763));
  XNOR2_X1  g338(.A(KEYINPUT33), .B(G1976), .ZN(new_n764));
  XOR2_X1   g339(.A(KEYINPUT32), .B(G1981), .Z(new_n765));
  AND2_X1   g340(.A1(new_n675), .A2(G6), .ZN(new_n766));
  AOI21_X1  g341(.A(new_n766), .B1(G305), .B2(G16), .ZN(new_n767));
  AOI22_X1  g342(.A1(new_n763), .A2(new_n764), .B1(new_n765), .B2(new_n767), .ZN(new_n768));
  OAI21_X1  g343(.A(new_n768), .B1(new_n763), .B2(new_n764), .ZN(new_n769));
  NAND2_X1  g344(.A1(new_n675), .A2(G22), .ZN(new_n770));
  OAI21_X1  g345(.A(new_n770), .B1(G166), .B2(new_n675), .ZN(new_n771));
  INV_X1    g346(.A(G1971), .ZN(new_n772));
  XNOR2_X1  g347(.A(new_n771), .B(new_n772), .ZN(new_n773));
  OAI21_X1  g348(.A(new_n773), .B1(new_n765), .B2(new_n767), .ZN(new_n774));
  NOR2_X1   g349(.A1(new_n769), .A2(new_n774), .ZN(new_n775));
  INV_X1    g350(.A(KEYINPUT34), .ZN(new_n776));
  NOR2_X1   g351(.A1(new_n775), .A2(new_n776), .ZN(new_n777));
  XOR2_X1   g352(.A(new_n777), .B(KEYINPUT88), .Z(new_n778));
  NAND2_X1  g353(.A1(new_n675), .A2(G24), .ZN(new_n779));
  OAI21_X1  g354(.A(new_n779), .B1(new_n579), .B2(new_n675), .ZN(new_n780));
  INV_X1    g355(.A(G1986), .ZN(new_n781));
  XNOR2_X1  g356(.A(new_n780), .B(new_n781), .ZN(new_n782));
  NAND2_X1  g357(.A1(new_n467), .A2(G131), .ZN(new_n783));
  NAND2_X1  g358(.A1(new_n478), .A2(G119), .ZN(new_n784));
  NOR2_X1   g359(.A1(new_n477), .A2(G107), .ZN(new_n785));
  OAI21_X1  g360(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n786));
  OAI211_X1 g361(.A(new_n783), .B(new_n784), .C1(new_n785), .C2(new_n786), .ZN(new_n787));
  XNOR2_X1  g362(.A(new_n787), .B(KEYINPUT87), .ZN(new_n788));
  MUX2_X1   g363(.A(G25), .B(new_n788), .S(G29), .Z(new_n789));
  XOR2_X1   g364(.A(KEYINPUT35), .B(G1991), .Z(new_n790));
  XNOR2_X1  g365(.A(new_n789), .B(new_n790), .ZN(new_n791));
  NAND3_X1  g366(.A1(new_n782), .A2(KEYINPUT89), .A3(new_n791), .ZN(new_n792));
  AOI21_X1  g367(.A(new_n792), .B1(new_n775), .B2(new_n776), .ZN(new_n793));
  NAND3_X1  g368(.A1(new_n778), .A2(KEYINPUT36), .A3(new_n793), .ZN(new_n794));
  INV_X1    g369(.A(new_n794), .ZN(new_n795));
  AOI21_X1  g370(.A(KEYINPUT36), .B1(new_n778), .B2(new_n793), .ZN(new_n796));
  NOR3_X1   g371(.A1(new_n760), .A2(new_n795), .A3(new_n796), .ZN(G311));
  INV_X1    g372(.A(G311), .ZN(G150));
  AOI22_X1  g373(.A1(new_n488), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n799));
  NOR2_X1   g374(.A1(new_n799), .A2(new_n510), .ZN(new_n800));
  OR2_X1    g375(.A1(new_n800), .A2(KEYINPUT99), .ZN(new_n801));
  NAND2_X1  g376(.A1(new_n516), .A2(G93), .ZN(new_n802));
  AOI22_X1  g377(.A1(new_n800), .A2(KEYINPUT99), .B1(G55), .B2(new_n495), .ZN(new_n803));
  NAND3_X1  g378(.A1(new_n801), .A2(new_n802), .A3(new_n803), .ZN(new_n804));
  NAND2_X1  g379(.A1(new_n804), .A2(G860), .ZN(new_n805));
  XOR2_X1   g380(.A(new_n805), .B(KEYINPUT37), .Z(new_n806));
  NAND2_X1  g381(.A1(new_n593), .A2(G559), .ZN(new_n807));
  XOR2_X1   g382(.A(KEYINPUT98), .B(KEYINPUT38), .Z(new_n808));
  XNOR2_X1  g383(.A(new_n807), .B(new_n808), .ZN(new_n809));
  NOR2_X1   g384(.A1(new_n536), .A2(new_n804), .ZN(new_n810));
  INV_X1    g385(.A(new_n810), .ZN(new_n811));
  INV_X1    g386(.A(new_n804), .ZN(new_n812));
  AOI21_X1  g387(.A(new_n812), .B1(new_n533), .B2(new_n535), .ZN(new_n813));
  INV_X1    g388(.A(new_n813), .ZN(new_n814));
  NAND2_X1  g389(.A1(new_n811), .A2(new_n814), .ZN(new_n815));
  XNOR2_X1  g390(.A(new_n809), .B(new_n815), .ZN(new_n816));
  INV_X1    g391(.A(KEYINPUT39), .ZN(new_n817));
  NAND2_X1  g392(.A1(new_n816), .A2(new_n817), .ZN(new_n818));
  XOR2_X1   g393(.A(new_n818), .B(KEYINPUT100), .Z(new_n819));
  INV_X1    g394(.A(G860), .ZN(new_n820));
  OAI21_X1  g395(.A(new_n820), .B1(new_n816), .B2(new_n817), .ZN(new_n821));
  OAI21_X1  g396(.A(new_n806), .B1(new_n819), .B2(new_n821), .ZN(G145));
  XNOR2_X1  g397(.A(new_n752), .B(new_n486), .ZN(new_n823));
  XNOR2_X1  g398(.A(new_n823), .B(new_n609), .ZN(new_n824));
  NAND2_X1  g399(.A1(new_n703), .A2(KEYINPUT101), .ZN(new_n825));
  XNOR2_X1  g400(.A(new_n825), .B(new_n685), .ZN(new_n826));
  NAND2_X1  g401(.A1(new_n478), .A2(G130), .ZN(new_n827));
  NOR2_X1   g402(.A1(new_n477), .A2(G118), .ZN(new_n828));
  OAI21_X1  g403(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n829));
  OAI21_X1  g404(.A(new_n827), .B1(new_n828), .B2(new_n829), .ZN(new_n830));
  AOI21_X1  g405(.A(new_n830), .B1(G142), .B2(new_n467), .ZN(new_n831));
  XNOR2_X1  g406(.A(new_n831), .B(new_n787), .ZN(new_n832));
  XNOR2_X1  g407(.A(new_n826), .B(new_n832), .ZN(new_n833));
  XNOR2_X1  g408(.A(new_n824), .B(new_n833), .ZN(new_n834));
  XNOR2_X1  g409(.A(G160), .B(new_n620), .ZN(new_n835));
  XNOR2_X1  g410(.A(G162), .B(new_n835), .ZN(new_n836));
  AOI21_X1  g411(.A(G37), .B1(new_n834), .B2(new_n836), .ZN(new_n837));
  OAI21_X1  g412(.A(new_n837), .B1(new_n836), .B2(new_n834), .ZN(new_n838));
  XNOR2_X1  g413(.A(new_n838), .B(KEYINPUT40), .ZN(G395));
  NAND2_X1  g414(.A1(new_n804), .A2(new_n581), .ZN(new_n840));
  INV_X1    g415(.A(G299), .ZN(new_n841));
  NAND2_X1  g416(.A1(new_n592), .A2(new_n841), .ZN(new_n842));
  INV_X1    g417(.A(KEYINPUT103), .ZN(new_n843));
  AOI21_X1  g418(.A(new_n590), .B1(new_n549), .B2(new_n560), .ZN(new_n844));
  AND3_X1   g419(.A1(new_n587), .A2(new_n843), .A3(new_n844), .ZN(new_n845));
  AOI21_X1  g420(.A(new_n843), .B1(new_n587), .B2(new_n844), .ZN(new_n846));
  OAI21_X1  g421(.A(new_n842), .B1(new_n845), .B2(new_n846), .ZN(new_n847));
  INV_X1    g422(.A(KEYINPUT104), .ZN(new_n848));
  NOR2_X1   g423(.A1(new_n845), .A2(new_n846), .ZN(new_n849));
  AOI21_X1  g424(.A(new_n590), .B1(new_n585), .B2(new_n586), .ZN(new_n850));
  OAI21_X1  g425(.A(KEYINPUT41), .B1(new_n850), .B2(G299), .ZN(new_n851));
  OAI21_X1  g426(.A(new_n848), .B1(new_n849), .B2(new_n851), .ZN(new_n852));
  INV_X1    g427(.A(KEYINPUT41), .ZN(new_n853));
  NAND2_X1  g428(.A1(new_n847), .A2(new_n853), .ZN(new_n854));
  AOI21_X1  g429(.A(new_n853), .B1(new_n592), .B2(new_n841), .ZN(new_n855));
  OAI211_X1 g430(.A(new_n855), .B(KEYINPUT104), .C1(new_n846), .C2(new_n845), .ZN(new_n856));
  NAND3_X1  g431(.A1(new_n852), .A2(new_n854), .A3(new_n856), .ZN(new_n857));
  XNOR2_X1  g432(.A(new_n815), .B(KEYINPUT102), .ZN(new_n858));
  XNOR2_X1  g433(.A(new_n858), .B(new_n603), .ZN(new_n859));
  MUX2_X1   g434(.A(new_n847), .B(new_n857), .S(new_n859), .Z(new_n860));
  XNOR2_X1  g435(.A(new_n579), .B(G166), .ZN(new_n861));
  XNOR2_X1  g436(.A(G288), .B(G305), .ZN(new_n862));
  XNOR2_X1  g437(.A(new_n861), .B(new_n862), .ZN(new_n863));
  XNOR2_X1  g438(.A(new_n863), .B(KEYINPUT42), .ZN(new_n864));
  XNOR2_X1  g439(.A(new_n860), .B(new_n864), .ZN(new_n865));
  OAI21_X1  g440(.A(new_n840), .B1(new_n865), .B2(new_n581), .ZN(G295));
  OAI21_X1  g441(.A(new_n840), .B1(new_n865), .B2(new_n581), .ZN(G331));
  INV_X1    g442(.A(KEYINPUT44), .ZN(new_n868));
  XOR2_X1   g443(.A(new_n863), .B(KEYINPUT108), .Z(new_n869));
  XNOR2_X1  g444(.A(G286), .B(G301), .ZN(new_n870));
  INV_X1    g445(.A(new_n870), .ZN(new_n871));
  NAND3_X1  g446(.A1(new_n811), .A2(new_n871), .A3(new_n814), .ZN(new_n872));
  OAI21_X1  g447(.A(new_n870), .B1(new_n810), .B2(new_n813), .ZN(new_n873));
  NAND3_X1  g448(.A1(new_n872), .A2(new_n847), .A3(new_n873), .ZN(new_n874));
  INV_X1    g449(.A(KEYINPUT106), .ZN(new_n875));
  NAND2_X1  g450(.A1(new_n873), .A2(new_n875), .ZN(new_n876));
  OAI211_X1 g451(.A(new_n870), .B(KEYINPUT106), .C1(new_n810), .C2(new_n813), .ZN(new_n877));
  AND3_X1   g452(.A1(new_n876), .A2(new_n872), .A3(new_n877), .ZN(new_n878));
  NOR2_X1   g453(.A1(new_n849), .A2(new_n851), .ZN(new_n879));
  AOI21_X1  g454(.A(new_n879), .B1(new_n853), .B2(new_n847), .ZN(new_n880));
  OAI21_X1  g455(.A(new_n874), .B1(new_n878), .B2(new_n880), .ZN(new_n881));
  AOI21_X1  g456(.A(G37), .B1(new_n869), .B2(new_n881), .ZN(new_n882));
  NAND2_X1  g457(.A1(new_n876), .A2(new_n877), .ZN(new_n883));
  NAND2_X1  g458(.A1(new_n872), .A2(new_n847), .ZN(new_n884));
  NOR2_X1   g459(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  NAND2_X1  g460(.A1(new_n872), .A2(new_n873), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n857), .A2(new_n886), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n887), .A2(KEYINPUT105), .ZN(new_n888));
  INV_X1    g463(.A(KEYINPUT105), .ZN(new_n889));
  NAND3_X1  g464(.A1(new_n857), .A2(new_n889), .A3(new_n886), .ZN(new_n890));
  AOI21_X1  g465(.A(new_n885), .B1(new_n888), .B2(new_n890), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n891), .A2(new_n863), .ZN(new_n892));
  NAND2_X1  g467(.A1(new_n882), .A2(new_n892), .ZN(new_n893));
  NAND2_X1  g468(.A1(new_n893), .A2(KEYINPUT43), .ZN(new_n894));
  INV_X1    g469(.A(G37), .ZN(new_n895));
  AOI21_X1  g470(.A(KEYINPUT43), .B1(new_n891), .B2(new_n863), .ZN(new_n896));
  OAI21_X1  g471(.A(new_n869), .B1(new_n891), .B2(KEYINPUT107), .ZN(new_n897));
  INV_X1    g472(.A(new_n885), .ZN(new_n898));
  INV_X1    g473(.A(new_n890), .ZN(new_n899));
  AOI21_X1  g474(.A(new_n889), .B1(new_n857), .B2(new_n886), .ZN(new_n900));
  OAI211_X1 g475(.A(new_n898), .B(KEYINPUT107), .C1(new_n899), .C2(new_n900), .ZN(new_n901));
  INV_X1    g476(.A(new_n901), .ZN(new_n902));
  OAI211_X1 g477(.A(new_n895), .B(new_n896), .C1(new_n897), .C2(new_n902), .ZN(new_n903));
  AOI21_X1  g478(.A(new_n868), .B1(new_n894), .B2(new_n903), .ZN(new_n904));
  OAI211_X1 g479(.A(new_n895), .B(new_n892), .C1(new_n897), .C2(new_n902), .ZN(new_n905));
  INV_X1    g480(.A(KEYINPUT109), .ZN(new_n906));
  AND3_X1   g481(.A1(new_n905), .A2(new_n906), .A3(KEYINPUT43), .ZN(new_n907));
  AOI21_X1  g482(.A(new_n906), .B1(new_n905), .B2(KEYINPUT43), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n882), .A2(new_n896), .ZN(new_n909));
  INV_X1    g484(.A(new_n909), .ZN(new_n910));
  NOR3_X1   g485(.A1(new_n907), .A2(new_n908), .A3(new_n910), .ZN(new_n911));
  AOI21_X1  g486(.A(new_n904), .B1(new_n911), .B2(new_n868), .ZN(G397));
  INV_X1    g487(.A(G2067), .ZN(new_n913));
  XNOR2_X1  g488(.A(new_n752), .B(new_n913), .ZN(new_n914));
  INV_X1    g489(.A(G1996), .ZN(new_n915));
  XNOR2_X1  g490(.A(new_n685), .B(new_n915), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n914), .A2(new_n916), .ZN(new_n917));
  INV_X1    g492(.A(new_n790), .ZN(new_n918));
  XNOR2_X1  g493(.A(new_n787), .B(new_n918), .ZN(new_n919));
  NOR2_X1   g494(.A1(new_n917), .A2(new_n919), .ZN(new_n920));
  INV_X1    g495(.A(G1384), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n486), .A2(new_n921), .ZN(new_n922));
  INV_X1    g497(.A(KEYINPUT45), .ZN(new_n923));
  NAND2_X1  g498(.A1(new_n922), .A2(new_n923), .ZN(new_n924));
  NAND2_X1  g499(.A1(G160), .A2(G40), .ZN(new_n925));
  NOR2_X1   g500(.A1(new_n924), .A2(new_n925), .ZN(new_n926));
  INV_X1    g501(.A(new_n926), .ZN(new_n927));
  NOR2_X1   g502(.A1(new_n920), .A2(new_n927), .ZN(new_n928));
  NOR3_X1   g503(.A1(new_n927), .A2(G1986), .A3(G290), .ZN(new_n929));
  AOI21_X1  g504(.A(new_n928), .B1(KEYINPUT48), .B2(new_n929), .ZN(new_n930));
  OAI21_X1  g505(.A(new_n930), .B1(KEYINPUT48), .B2(new_n929), .ZN(new_n931));
  NOR3_X1   g506(.A1(new_n917), .A2(new_n788), .A3(new_n918), .ZN(new_n932));
  NOR2_X1   g507(.A1(new_n752), .A2(G2067), .ZN(new_n933));
  OAI21_X1  g508(.A(new_n926), .B1(new_n932), .B2(new_n933), .ZN(new_n934));
  NOR2_X1   g509(.A1(new_n927), .A2(G1996), .ZN(new_n935));
  NAND2_X1  g510(.A1(new_n935), .A2(KEYINPUT46), .ZN(new_n936));
  XOR2_X1   g511(.A(new_n936), .B(KEYINPUT125), .Z(new_n937));
  AOI21_X1  g512(.A(new_n927), .B1(new_n686), .B2(new_n914), .ZN(new_n938));
  XOR2_X1   g513(.A(new_n938), .B(KEYINPUT126), .Z(new_n939));
  OAI211_X1 g514(.A(new_n937), .B(new_n939), .C1(KEYINPUT46), .C2(new_n935), .ZN(new_n940));
  INV_X1    g515(.A(KEYINPUT47), .ZN(new_n941));
  OAI211_X1 g516(.A(new_n931), .B(new_n934), .C1(new_n940), .C2(new_n941), .ZN(new_n942));
  AOI21_X1  g517(.A(new_n942), .B1(new_n941), .B2(new_n940), .ZN(new_n943));
  INV_X1    g518(.A(KEYINPUT52), .ZN(new_n944));
  INV_X1    g519(.A(new_n922), .ZN(new_n945));
  INV_X1    g520(.A(new_n925), .ZN(new_n946));
  NAND2_X1  g521(.A1(new_n945), .A2(new_n946), .ZN(new_n947));
  NAND2_X1  g522(.A1(new_n947), .A2(G8), .ZN(new_n948));
  AOI21_X1  g523(.A(new_n948), .B1(G1976), .B2(new_n761), .ZN(new_n949));
  AOI21_X1  g524(.A(new_n944), .B1(new_n949), .B2(KEYINPUT112), .ZN(new_n950));
  OAI21_X1  g525(.A(new_n950), .B1(KEYINPUT112), .B2(new_n949), .ZN(new_n951));
  INV_X1    g526(.A(KEYINPUT49), .ZN(new_n952));
  AND2_X1   g527(.A1(new_n516), .A2(G86), .ZN(new_n953));
  INV_X1    g528(.A(new_n573), .ZN(new_n954));
  OAI21_X1  g529(.A(G1981), .B1(new_n953), .B2(new_n954), .ZN(new_n955));
  OAI21_X1  g530(.A(new_n955), .B1(G305), .B2(G1981), .ZN(new_n956));
  AOI21_X1  g531(.A(new_n948), .B1(new_n952), .B2(new_n956), .ZN(new_n957));
  OAI21_X1  g532(.A(new_n957), .B1(new_n952), .B2(new_n956), .ZN(new_n958));
  XOR2_X1   g533(.A(KEYINPUT113), .B(G1976), .Z(new_n959));
  AOI21_X1  g534(.A(KEYINPUT52), .B1(G288), .B2(new_n959), .ZN(new_n960));
  NAND2_X1  g535(.A1(new_n949), .A2(new_n960), .ZN(new_n961));
  AND2_X1   g536(.A1(new_n961), .A2(KEYINPUT114), .ZN(new_n962));
  NOR2_X1   g537(.A1(new_n961), .A2(KEYINPUT114), .ZN(new_n963));
  OAI211_X1 g538(.A(new_n951), .B(new_n958), .C1(new_n962), .C2(new_n963), .ZN(new_n964));
  INV_X1    g539(.A(G8), .ZN(new_n965));
  NAND2_X1  g540(.A1(new_n922), .A2(KEYINPUT50), .ZN(new_n966));
  XOR2_X1   g541(.A(new_n966), .B(KEYINPUT110), .Z(new_n967));
  INV_X1    g542(.A(G2090), .ZN(new_n968));
  INV_X1    g543(.A(KEYINPUT50), .ZN(new_n969));
  AOI21_X1  g544(.A(new_n925), .B1(new_n945), .B2(new_n969), .ZN(new_n970));
  NAND3_X1  g545(.A1(new_n967), .A2(new_n968), .A3(new_n970), .ZN(new_n971));
  NAND2_X1  g546(.A1(new_n945), .A2(KEYINPUT45), .ZN(new_n972));
  NAND3_X1  g547(.A1(new_n972), .A2(new_n924), .A3(new_n946), .ZN(new_n973));
  NAND2_X1  g548(.A1(new_n973), .A2(new_n772), .ZN(new_n974));
  AOI21_X1  g549(.A(new_n965), .B1(new_n971), .B2(new_n974), .ZN(new_n975));
  NAND2_X1  g550(.A1(G303), .A2(G8), .ZN(new_n976));
  XOR2_X1   g551(.A(new_n976), .B(KEYINPUT55), .Z(new_n977));
  XNOR2_X1  g552(.A(new_n977), .B(KEYINPUT111), .ZN(new_n978));
  NAND2_X1  g553(.A1(new_n975), .A2(new_n978), .ZN(new_n979));
  NOR2_X1   g554(.A1(G305), .A2(G1981), .ZN(new_n980));
  NOR2_X1   g555(.A1(G288), .A2(G1976), .ZN(new_n981));
  AOI21_X1  g556(.A(new_n980), .B1(new_n958), .B2(new_n981), .ZN(new_n982));
  OAI22_X1  g557(.A1(new_n964), .A2(new_n979), .B1(new_n948), .B2(new_n982), .ZN(new_n983));
  INV_X1    g558(.A(new_n983), .ZN(new_n984));
  NAND2_X1  g559(.A1(new_n970), .A2(new_n966), .ZN(new_n985));
  OAI21_X1  g560(.A(new_n974), .B1(G2090), .B2(new_n985), .ZN(new_n986));
  OR2_X1    g561(.A1(new_n986), .A2(KEYINPUT115), .ZN(new_n987));
  AOI21_X1  g562(.A(new_n965), .B1(new_n986), .B2(KEYINPUT115), .ZN(new_n988));
  AOI21_X1  g563(.A(new_n977), .B1(new_n987), .B2(new_n988), .ZN(new_n989));
  AOI211_X1 g564(.A(new_n989), .B(new_n964), .C1(new_n975), .C2(new_n978), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n967), .A2(new_n970), .ZN(new_n991));
  INV_X1    g566(.A(new_n991), .ZN(new_n992));
  INV_X1    g567(.A(G2084), .ZN(new_n993));
  INV_X1    g568(.A(G1966), .ZN(new_n994));
  AOI22_X1  g569(.A1(new_n992), .A2(new_n993), .B1(new_n994), .B2(new_n973), .ZN(new_n995));
  NOR3_X1   g570(.A1(new_n995), .A2(new_n965), .A3(G286), .ZN(new_n996));
  AOI21_X1  g571(.A(KEYINPUT63), .B1(new_n990), .B2(new_n996), .ZN(new_n997));
  NAND3_X1  g572(.A1(new_n996), .A2(KEYINPUT63), .A3(new_n979), .ZN(new_n998));
  INV_X1    g573(.A(KEYINPUT116), .ZN(new_n999));
  OR2_X1    g574(.A1(new_n975), .A2(new_n999), .ZN(new_n1000));
  AOI21_X1  g575(.A(new_n977), .B1(new_n975), .B2(new_n999), .ZN(new_n1001));
  NAND2_X1  g576(.A1(new_n1000), .A2(new_n1001), .ZN(new_n1002));
  INV_X1    g577(.A(new_n1002), .ZN(new_n1003));
  OAI21_X1  g578(.A(KEYINPUT117), .B1(new_n1003), .B2(new_n964), .ZN(new_n1004));
  INV_X1    g579(.A(new_n964), .ZN(new_n1005));
  INV_X1    g580(.A(KEYINPUT117), .ZN(new_n1006));
  NAND3_X1  g581(.A1(new_n1005), .A2(new_n1002), .A3(new_n1006), .ZN(new_n1007));
  AOI21_X1  g582(.A(new_n998), .B1(new_n1004), .B2(new_n1007), .ZN(new_n1008));
  OAI21_X1  g583(.A(new_n984), .B1(new_n997), .B2(new_n1008), .ZN(new_n1009));
  INV_X1    g584(.A(new_n973), .ZN(new_n1010));
  XNOR2_X1  g585(.A(KEYINPUT56), .B(G2072), .ZN(new_n1011));
  XOR2_X1   g586(.A(KEYINPUT118), .B(G1956), .Z(new_n1012));
  AOI22_X1  g587(.A1(new_n1010), .A2(new_n1011), .B1(new_n985), .B2(new_n1012), .ZN(new_n1013));
  XOR2_X1   g588(.A(G299), .B(KEYINPUT57), .Z(new_n1014));
  AND2_X1   g589(.A1(new_n1013), .A2(new_n1014), .ZN(new_n1015));
  XNOR2_X1  g590(.A(new_n947), .B(KEYINPUT119), .ZN(new_n1016));
  AOI22_X1  g591(.A1(new_n991), .A2(new_n756), .B1(new_n1016), .B2(new_n913), .ZN(new_n1017));
  NOR3_X1   g592(.A1(new_n1015), .A2(new_n1017), .A3(new_n592), .ZN(new_n1018));
  NOR2_X1   g593(.A1(new_n1013), .A2(new_n1014), .ZN(new_n1019));
  NOR2_X1   g594(.A1(new_n1018), .A2(new_n1019), .ZN(new_n1020));
  XNOR2_X1  g595(.A(KEYINPUT58), .B(G1341), .ZN(new_n1021));
  OR2_X1    g596(.A1(new_n1016), .A2(new_n1021), .ZN(new_n1022));
  NAND2_X1  g597(.A1(new_n1010), .A2(new_n915), .ZN(new_n1023));
  AOI21_X1  g598(.A(new_n536), .B1(new_n1022), .B2(new_n1023), .ZN(new_n1024));
  OR2_X1    g599(.A1(new_n1024), .A2(KEYINPUT59), .ZN(new_n1025));
  INV_X1    g600(.A(KEYINPUT61), .ZN(new_n1026));
  OR3_X1    g601(.A1(new_n1015), .A2(new_n1019), .A3(new_n1026), .ZN(new_n1027));
  OAI21_X1  g602(.A(new_n1026), .B1(new_n1015), .B2(new_n1019), .ZN(new_n1028));
  NAND2_X1  g603(.A1(new_n1024), .A2(KEYINPUT59), .ZN(new_n1029));
  NAND4_X1  g604(.A1(new_n1025), .A2(new_n1027), .A3(new_n1028), .A4(new_n1029), .ZN(new_n1030));
  AND3_X1   g605(.A1(new_n1017), .A2(KEYINPUT60), .A3(new_n850), .ZN(new_n1031));
  AOI21_X1  g606(.A(new_n850), .B1(new_n1017), .B2(KEYINPUT60), .ZN(new_n1032));
  NOR2_X1   g607(.A1(new_n1017), .A2(KEYINPUT60), .ZN(new_n1033));
  NOR3_X1   g608(.A1(new_n1031), .A2(new_n1032), .A3(new_n1033), .ZN(new_n1034));
  OAI21_X1  g609(.A(new_n1020), .B1(new_n1030), .B2(new_n1034), .ZN(new_n1035));
  XNOR2_X1  g610(.A(KEYINPUT121), .B(KEYINPUT54), .ZN(new_n1036));
  INV_X1    g611(.A(G1961), .ZN(new_n1037));
  NAND2_X1  g612(.A1(new_n991), .A2(new_n1037), .ZN(new_n1038));
  INV_X1    g613(.A(G2078), .ZN(new_n1039));
  NAND3_X1  g614(.A1(new_n1010), .A2(KEYINPUT53), .A3(new_n1039), .ZN(new_n1040));
  INV_X1    g615(.A(KEYINPUT53), .ZN(new_n1041));
  OAI21_X1  g616(.A(new_n1041), .B1(new_n973), .B2(G2078), .ZN(new_n1042));
  NAND3_X1  g617(.A1(new_n1038), .A2(new_n1040), .A3(new_n1042), .ZN(new_n1043));
  NAND2_X1  g618(.A1(new_n1043), .A2(G171), .ZN(new_n1044));
  NAND4_X1  g619(.A1(new_n1038), .A2(G301), .A3(new_n1040), .A4(new_n1042), .ZN(new_n1045));
  AOI21_X1  g620(.A(new_n1036), .B1(new_n1044), .B2(new_n1045), .ZN(new_n1046));
  NAND2_X1  g621(.A1(new_n973), .A2(new_n994), .ZN(new_n1047));
  OAI211_X1 g622(.A(G168), .B(new_n1047), .C1(new_n991), .C2(G2084), .ZN(new_n1048));
  AOI21_X1  g623(.A(KEYINPUT51), .B1(new_n1048), .B2(G8), .ZN(new_n1049));
  INV_X1    g624(.A(KEYINPUT120), .ZN(new_n1050));
  NOR2_X1   g625(.A1(new_n1049), .A2(new_n1050), .ZN(new_n1051));
  NAND3_X1  g626(.A1(new_n1048), .A2(KEYINPUT51), .A3(G8), .ZN(new_n1052));
  NAND2_X1  g627(.A1(new_n1051), .A2(new_n1052), .ZN(new_n1053));
  NOR2_X1   g628(.A1(new_n995), .A2(new_n965), .ZN(new_n1054));
  AOI22_X1  g629(.A1(new_n1054), .A2(G286), .B1(new_n1049), .B2(new_n1050), .ZN(new_n1055));
  AOI21_X1  g630(.A(new_n1046), .B1(new_n1053), .B2(new_n1055), .ZN(new_n1056));
  NAND2_X1  g631(.A1(new_n1044), .A2(KEYINPUT122), .ZN(new_n1057));
  AND2_X1   g632(.A1(new_n1045), .A2(KEYINPUT54), .ZN(new_n1058));
  INV_X1    g633(.A(KEYINPUT122), .ZN(new_n1059));
  NAND3_X1  g634(.A1(new_n1043), .A2(new_n1059), .A3(G171), .ZN(new_n1060));
  NAND3_X1  g635(.A1(new_n1057), .A2(new_n1058), .A3(new_n1060), .ZN(new_n1061));
  AND2_X1   g636(.A1(new_n1061), .A2(KEYINPUT123), .ZN(new_n1062));
  NOR2_X1   g637(.A1(new_n1061), .A2(KEYINPUT123), .ZN(new_n1063));
  OAI211_X1 g638(.A(new_n1035), .B(new_n1056), .C1(new_n1062), .C2(new_n1063), .ZN(new_n1064));
  INV_X1    g639(.A(new_n1044), .ZN(new_n1065));
  INV_X1    g640(.A(KEYINPUT62), .ZN(new_n1066));
  NAND3_X1  g641(.A1(new_n1053), .A2(new_n1055), .A3(new_n1066), .ZN(new_n1067));
  AOI21_X1  g642(.A(new_n1066), .B1(new_n1053), .B2(new_n1055), .ZN(new_n1068));
  INV_X1    g643(.A(KEYINPUT124), .ZN(new_n1069));
  OAI211_X1 g644(.A(new_n1065), .B(new_n1067), .C1(new_n1068), .C2(new_n1069), .ZN(new_n1070));
  AND2_X1   g645(.A1(new_n1068), .A2(new_n1069), .ZN(new_n1071));
  OAI21_X1  g646(.A(new_n1064), .B1(new_n1070), .B2(new_n1071), .ZN(new_n1072));
  AOI21_X1  g647(.A(new_n1009), .B1(new_n1072), .B2(new_n990), .ZN(new_n1073));
  XNOR2_X1  g648(.A(new_n579), .B(G1986), .ZN(new_n1074));
  AOI21_X1  g649(.A(new_n927), .B1(new_n920), .B2(new_n1074), .ZN(new_n1075));
  OAI21_X1  g650(.A(new_n943), .B1(new_n1073), .B2(new_n1075), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g651(.A(KEYINPUT127), .ZN(new_n1078));
  NOR3_X1   g652(.A1(G401), .A2(new_n458), .A3(G227), .ZN(new_n1079));
  NAND4_X1  g653(.A1(new_n838), .A2(new_n673), .A3(new_n672), .A4(new_n1079), .ZN(new_n1080));
  NAND2_X1  g654(.A1(new_n905), .A2(KEYINPUT43), .ZN(new_n1081));
  AOI21_X1  g655(.A(new_n910), .B1(new_n1081), .B2(KEYINPUT109), .ZN(new_n1082));
  NAND3_X1  g656(.A1(new_n905), .A2(new_n906), .A3(KEYINPUT43), .ZN(new_n1083));
  AOI211_X1 g657(.A(new_n1078), .B(new_n1080), .C1(new_n1082), .C2(new_n1083), .ZN(new_n1084));
  NAND2_X1  g658(.A1(new_n1081), .A2(KEYINPUT109), .ZN(new_n1085));
  NAND3_X1  g659(.A1(new_n1085), .A2(new_n1083), .A3(new_n909), .ZN(new_n1086));
  INV_X1    g660(.A(new_n1080), .ZN(new_n1087));
  AOI21_X1  g661(.A(KEYINPUT127), .B1(new_n1086), .B2(new_n1087), .ZN(new_n1088));
  NOR2_X1   g662(.A1(new_n1084), .A2(new_n1088), .ZN(G308));
  OAI21_X1  g663(.A(new_n1078), .B1(new_n911), .B2(new_n1080), .ZN(new_n1090));
  NAND3_X1  g664(.A1(new_n1086), .A2(KEYINPUT127), .A3(new_n1087), .ZN(new_n1091));
  NAND2_X1  g665(.A1(new_n1090), .A2(new_n1091), .ZN(G225));
endmodule


