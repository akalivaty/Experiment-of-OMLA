//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 0 1 1 0 1 1 0 0 0 1 0 0 0 1 1 1 0 0 1 0 1 1 0 1 1 1 1 1 0 1 0 0 1 1 1 0 0 1 0 0 1 1 0 0 0 0 1 1 1 1 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:19:37 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n701, new_n702, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n709, new_n710, new_n711, new_n713, new_n714, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n764, new_n765, new_n766,
    new_n767, new_n768, new_n769, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n783, new_n784, new_n785, new_n786, new_n787, new_n788, new_n790,
    new_n791, new_n792, new_n793, new_n795, new_n796, new_n797, new_n799,
    new_n800, new_n801, new_n802, new_n803, new_n804, new_n805, new_n807,
    new_n809, new_n810, new_n811, new_n812, new_n813, new_n814, new_n815,
    new_n816, new_n817, new_n818, new_n819, new_n820, new_n821, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n832, new_n833, new_n834, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n894, new_n895, new_n897, new_n898,
    new_n899, new_n901, new_n902, new_n903, new_n904, new_n905, new_n906,
    new_n907, new_n908, new_n909, new_n910, new_n911, new_n912, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n939, new_n940, new_n941, new_n942,
    new_n943, new_n944, new_n945, new_n946, new_n947, new_n948, new_n949,
    new_n950, new_n951, new_n952, new_n953, new_n954, new_n955, new_n956,
    new_n957, new_n958, new_n959, new_n960, new_n961, new_n962, new_n963,
    new_n964, new_n965, new_n966, new_n968, new_n969, new_n970, new_n971,
    new_n972, new_n973, new_n974, new_n975, new_n976, new_n977, new_n978,
    new_n979, new_n980, new_n981, new_n982, new_n983, new_n984, new_n985,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n993, new_n994,
    new_n995, new_n996, new_n997, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1021,
    new_n1022, new_n1023, new_n1025, new_n1026, new_n1027, new_n1029,
    new_n1030, new_n1031, new_n1032, new_n1033, new_n1034, new_n1035,
    new_n1037, new_n1038, new_n1039, new_n1040, new_n1041, new_n1042,
    new_n1043, new_n1045, new_n1046, new_n1047, new_n1048, new_n1050,
    new_n1051;
  NAND2_X1  g000(.A1(G229gat), .A2(G233gat), .ZN(new_n202));
  XNOR2_X1  g001(.A(new_n202), .B(KEYINPUT92), .ZN(new_n203));
  XNOR2_X1  g002(.A(new_n203), .B(KEYINPUT13), .ZN(new_n204));
  INV_X1    g003(.A(new_n204), .ZN(new_n205));
  INV_X1    g004(.A(KEYINPUT89), .ZN(new_n206));
  OR2_X1    g005(.A1(KEYINPUT14), .A2(G29gat), .ZN(new_n207));
  NAND2_X1  g006(.A1(KEYINPUT14), .A2(G29gat), .ZN(new_n208));
  AOI21_X1  g007(.A(G36gat), .B1(new_n207), .B2(new_n208), .ZN(new_n209));
  INV_X1    g008(.A(G29gat), .ZN(new_n210));
  AND3_X1   g009(.A1(new_n210), .A2(KEYINPUT14), .A3(G36gat), .ZN(new_n211));
  OAI21_X1  g010(.A(new_n206), .B1(new_n209), .B2(new_n211), .ZN(new_n212));
  INV_X1    g011(.A(G43gat), .ZN(new_n213));
  INV_X1    g012(.A(G50gat), .ZN(new_n214));
  NAND2_X1  g013(.A1(new_n213), .A2(new_n214), .ZN(new_n215));
  INV_X1    g014(.A(KEYINPUT15), .ZN(new_n216));
  NAND2_X1  g015(.A1(G43gat), .A2(G50gat), .ZN(new_n217));
  NAND3_X1  g016(.A1(new_n215), .A2(new_n216), .A3(new_n217), .ZN(new_n218));
  OAI21_X1  g017(.A(new_n218), .B1(new_n209), .B2(new_n211), .ZN(new_n219));
  AOI21_X1  g018(.A(new_n216), .B1(new_n215), .B2(new_n217), .ZN(new_n220));
  INV_X1    g019(.A(new_n220), .ZN(new_n221));
  NAND3_X1  g020(.A1(new_n212), .A2(new_n219), .A3(new_n221), .ZN(new_n222));
  OAI221_X1 g021(.A(new_n218), .B1(new_n220), .B2(new_n206), .C1(new_n209), .C2(new_n211), .ZN(new_n223));
  AOI21_X1  g022(.A(KEYINPUT90), .B1(new_n222), .B2(new_n223), .ZN(new_n224));
  INV_X1    g023(.A(new_n224), .ZN(new_n225));
  NAND3_X1  g024(.A1(new_n222), .A2(new_n223), .A3(KEYINPUT90), .ZN(new_n226));
  XNOR2_X1  g025(.A(G15gat), .B(G22gat), .ZN(new_n227));
  INV_X1    g026(.A(G1gat), .ZN(new_n228));
  NAND2_X1  g027(.A1(new_n228), .A2(KEYINPUT16), .ZN(new_n229));
  AND2_X1   g028(.A1(new_n227), .A2(new_n229), .ZN(new_n230));
  NOR2_X1   g029(.A1(new_n227), .A2(G1gat), .ZN(new_n231));
  OAI21_X1  g030(.A(G8gat), .B1(new_n230), .B2(new_n231), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n227), .A2(new_n229), .ZN(new_n233));
  INV_X1    g032(.A(G8gat), .ZN(new_n234));
  OAI211_X1 g033(.A(new_n233), .B(new_n234), .C1(G1gat), .C2(new_n227), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n232), .A2(new_n235), .ZN(new_n236));
  INV_X1    g035(.A(new_n236), .ZN(new_n237));
  NAND3_X1  g036(.A1(new_n225), .A2(new_n226), .A3(new_n237), .ZN(new_n238));
  INV_X1    g037(.A(new_n226), .ZN(new_n239));
  OAI21_X1  g038(.A(new_n236), .B1(new_n239), .B2(new_n224), .ZN(new_n240));
  AOI21_X1  g039(.A(new_n205), .B1(new_n238), .B2(new_n240), .ZN(new_n241));
  INV_X1    g040(.A(new_n203), .ZN(new_n242));
  AOI21_X1  g041(.A(KEYINPUT17), .B1(new_n225), .B2(new_n226), .ZN(new_n243));
  AND3_X1   g042(.A1(new_n232), .A2(KEYINPUT91), .A3(new_n235), .ZN(new_n244));
  AOI21_X1  g043(.A(KEYINPUT91), .B1(new_n232), .B2(new_n235), .ZN(new_n245));
  NOR2_X1   g044(.A1(new_n244), .A2(new_n245), .ZN(new_n246));
  NAND2_X1  g045(.A1(new_n222), .A2(new_n223), .ZN(new_n247));
  NAND2_X1  g046(.A1(new_n247), .A2(KEYINPUT17), .ZN(new_n248));
  NAND2_X1  g047(.A1(new_n246), .A2(new_n248), .ZN(new_n249));
  OAI211_X1 g048(.A(new_n242), .B(new_n240), .C1(new_n243), .C2(new_n249), .ZN(new_n250));
  INV_X1    g049(.A(KEYINPUT18), .ZN(new_n251));
  AOI21_X1  g050(.A(new_n241), .B1(new_n250), .B2(new_n251), .ZN(new_n252));
  INV_X1    g051(.A(KEYINPUT17), .ZN(new_n253));
  OAI21_X1  g052(.A(new_n253), .B1(new_n239), .B2(new_n224), .ZN(new_n254));
  NAND3_X1  g053(.A1(new_n254), .A2(new_n248), .A3(new_n246), .ZN(new_n255));
  NAND4_X1  g054(.A1(new_n255), .A2(KEYINPUT18), .A3(new_n242), .A4(new_n240), .ZN(new_n256));
  NAND2_X1  g055(.A1(new_n252), .A2(new_n256), .ZN(new_n257));
  XNOR2_X1  g056(.A(G113gat), .B(G141gat), .ZN(new_n258));
  XNOR2_X1  g057(.A(new_n258), .B(G197gat), .ZN(new_n259));
  XOR2_X1   g058(.A(KEYINPUT11), .B(G169gat), .Z(new_n260));
  XNOR2_X1  g059(.A(new_n259), .B(new_n260), .ZN(new_n261));
  XNOR2_X1  g060(.A(new_n261), .B(KEYINPUT12), .ZN(new_n262));
  INV_X1    g061(.A(new_n262), .ZN(new_n263));
  NAND2_X1  g062(.A1(new_n257), .A2(new_n263), .ZN(new_n264));
  NAND3_X1  g063(.A1(new_n252), .A2(new_n262), .A3(new_n256), .ZN(new_n265));
  NAND2_X1  g064(.A1(new_n264), .A2(new_n265), .ZN(new_n266));
  INV_X1    g065(.A(new_n266), .ZN(new_n267));
  XNOR2_X1  g066(.A(G15gat), .B(G43gat), .ZN(new_n268));
  XNOR2_X1  g067(.A(G71gat), .B(G99gat), .ZN(new_n269));
  XNOR2_X1  g068(.A(new_n268), .B(new_n269), .ZN(new_n270));
  XNOR2_X1  g069(.A(KEYINPUT27), .B(G183gat), .ZN(new_n271));
  INV_X1    g070(.A(G190gat), .ZN(new_n272));
  NAND3_X1  g071(.A1(new_n271), .A2(KEYINPUT28), .A3(new_n272), .ZN(new_n273));
  INV_X1    g072(.A(G183gat), .ZN(new_n274));
  NOR2_X1   g073(.A1(new_n274), .A2(KEYINPUT27), .ZN(new_n275));
  AOI21_X1  g074(.A(G190gat), .B1(new_n275), .B2(KEYINPUT69), .ZN(new_n276));
  INV_X1    g075(.A(KEYINPUT68), .ZN(new_n277));
  NAND3_X1  g076(.A1(new_n277), .A2(KEYINPUT69), .A3(G183gat), .ZN(new_n278));
  NAND2_X1  g077(.A1(new_n274), .A2(KEYINPUT68), .ZN(new_n279));
  NAND3_X1  g078(.A1(new_n278), .A2(KEYINPUT27), .A3(new_n279), .ZN(new_n280));
  NAND3_X1  g079(.A1(new_n276), .A2(new_n280), .A3(KEYINPUT70), .ZN(new_n281));
  INV_X1    g080(.A(KEYINPUT28), .ZN(new_n282));
  NAND2_X1  g081(.A1(new_n281), .A2(new_n282), .ZN(new_n283));
  AOI21_X1  g082(.A(KEYINPUT70), .B1(new_n276), .B2(new_n280), .ZN(new_n284));
  OAI21_X1  g083(.A(new_n273), .B1(new_n283), .B2(new_n284), .ZN(new_n285));
  NOR2_X1   g084(.A1(G169gat), .A2(G176gat), .ZN(new_n286));
  NAND2_X1  g085(.A1(new_n286), .A2(KEYINPUT26), .ZN(new_n287));
  OAI21_X1  g086(.A(new_n287), .B1(new_n274), .B2(new_n272), .ZN(new_n288));
  NAND2_X1  g087(.A1(G169gat), .A2(G176gat), .ZN(new_n289));
  NOR2_X1   g088(.A1(new_n286), .A2(KEYINPUT26), .ZN(new_n290));
  AOI21_X1  g089(.A(new_n288), .B1(new_n289), .B2(new_n290), .ZN(new_n291));
  NAND2_X1  g090(.A1(new_n285), .A2(new_n291), .ZN(new_n292));
  NAND2_X1  g091(.A1(new_n286), .A2(KEYINPUT23), .ZN(new_n293));
  INV_X1    g092(.A(KEYINPUT23), .ZN(new_n294));
  OAI21_X1  g093(.A(new_n294), .B1(G169gat), .B2(G176gat), .ZN(new_n295));
  NAND3_X1  g094(.A1(new_n293), .A2(new_n289), .A3(new_n295), .ZN(new_n296));
  INV_X1    g095(.A(new_n296), .ZN(new_n297));
  AOI21_X1  g096(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n298));
  XOR2_X1   g097(.A(new_n298), .B(KEYINPUT67), .Z(new_n299));
  AND2_X1   g098(.A1(KEYINPUT24), .A2(G183gat), .ZN(new_n300));
  NAND2_X1  g099(.A1(new_n300), .A2(G190gat), .ZN(new_n301));
  NAND2_X1  g100(.A1(new_n277), .A2(G183gat), .ZN(new_n302));
  NAND2_X1  g101(.A1(new_n279), .A2(new_n302), .ZN(new_n303));
  OAI21_X1  g102(.A(new_n301), .B1(new_n303), .B2(G190gat), .ZN(new_n304));
  OAI211_X1 g103(.A(KEYINPUT25), .B(new_n297), .C1(new_n299), .C2(new_n304), .ZN(new_n305));
  XOR2_X1   g104(.A(KEYINPUT64), .B(KEYINPUT25), .Z(new_n306));
  INV_X1    g105(.A(new_n306), .ZN(new_n307));
  INV_X1    g106(.A(KEYINPUT65), .ZN(new_n308));
  NOR2_X1   g107(.A1(G183gat), .A2(G190gat), .ZN(new_n309));
  AOI21_X1  g108(.A(new_n309), .B1(new_n300), .B2(G190gat), .ZN(new_n310));
  INV_X1    g109(.A(new_n298), .ZN(new_n311));
  AOI22_X1  g110(.A1(new_n296), .A2(new_n308), .B1(new_n310), .B2(new_n311), .ZN(new_n312));
  NAND4_X1  g111(.A1(new_n293), .A2(KEYINPUT65), .A3(new_n295), .A4(new_n289), .ZN(new_n313));
  AOI21_X1  g112(.A(new_n307), .B1(new_n312), .B2(new_n313), .ZN(new_n314));
  OAI21_X1  g113(.A(new_n305), .B1(new_n314), .B2(KEYINPUT66), .ZN(new_n315));
  NAND2_X1  g114(.A1(new_n295), .A2(new_n289), .ZN(new_n316));
  NOR3_X1   g115(.A1(new_n294), .A2(G169gat), .A3(G176gat), .ZN(new_n317));
  OAI21_X1  g116(.A(new_n308), .B1(new_n316), .B2(new_n317), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n310), .A2(new_n311), .ZN(new_n319));
  NAND3_X1  g118(.A1(new_n318), .A2(new_n313), .A3(new_n319), .ZN(new_n320));
  NAND3_X1  g119(.A1(new_n320), .A2(KEYINPUT66), .A3(new_n306), .ZN(new_n321));
  INV_X1    g120(.A(new_n321), .ZN(new_n322));
  OAI21_X1  g121(.A(new_n292), .B1(new_n315), .B2(new_n322), .ZN(new_n323));
  XNOR2_X1  g122(.A(KEYINPUT71), .B(G134gat), .ZN(new_n324));
  NAND2_X1  g123(.A1(new_n324), .A2(G127gat), .ZN(new_n325));
  OR2_X1    g124(.A1(KEYINPUT72), .A2(G127gat), .ZN(new_n326));
  NAND2_X1  g125(.A1(KEYINPUT72), .A2(G127gat), .ZN(new_n327));
  NAND3_X1  g126(.A1(new_n326), .A2(G134gat), .A3(new_n327), .ZN(new_n328));
  XOR2_X1   g127(.A(G113gat), .B(G120gat), .Z(new_n329));
  INV_X1    g128(.A(KEYINPUT1), .ZN(new_n330));
  AOI22_X1  g129(.A1(new_n325), .A2(new_n328), .B1(new_n329), .B2(new_n330), .ZN(new_n331));
  INV_X1    g130(.A(G127gat), .ZN(new_n332));
  AND2_X1   g131(.A1(new_n332), .A2(G134gat), .ZN(new_n333));
  OAI21_X1  g132(.A(new_n330), .B1(new_n332), .B2(G134gat), .ZN(new_n334));
  NOR2_X1   g133(.A1(new_n333), .A2(new_n334), .ZN(new_n335));
  INV_X1    g134(.A(new_n335), .ZN(new_n336));
  OR2_X1    g135(.A1(KEYINPUT73), .A2(G120gat), .ZN(new_n337));
  INV_X1    g136(.A(KEYINPUT74), .ZN(new_n338));
  NAND2_X1  g137(.A1(KEYINPUT73), .A2(G120gat), .ZN(new_n339));
  NAND4_X1  g138(.A1(new_n337), .A2(new_n338), .A3(G113gat), .A4(new_n339), .ZN(new_n340));
  AND2_X1   g139(.A1(KEYINPUT73), .A2(G120gat), .ZN(new_n341));
  NOR2_X1   g140(.A1(KEYINPUT73), .A2(G120gat), .ZN(new_n342));
  INV_X1    g141(.A(G113gat), .ZN(new_n343));
  NOR3_X1   g142(.A1(new_n341), .A2(new_n342), .A3(new_n343), .ZN(new_n344));
  INV_X1    g143(.A(G120gat), .ZN(new_n345));
  OAI21_X1  g144(.A(KEYINPUT74), .B1(new_n345), .B2(G113gat), .ZN(new_n346));
  OAI21_X1  g145(.A(new_n340), .B1(new_n344), .B2(new_n346), .ZN(new_n347));
  INV_X1    g146(.A(KEYINPUT75), .ZN(new_n348));
  AOI21_X1  g147(.A(new_n336), .B1(new_n347), .B2(new_n348), .ZN(new_n349));
  OAI211_X1 g148(.A(KEYINPUT75), .B(new_n340), .C1(new_n344), .C2(new_n346), .ZN(new_n350));
  AOI21_X1  g149(.A(new_n331), .B1(new_n349), .B2(new_n350), .ZN(new_n351));
  NAND2_X1  g150(.A1(new_n323), .A2(new_n351), .ZN(new_n352));
  NAND2_X1  g151(.A1(new_n320), .A2(new_n306), .ZN(new_n353));
  INV_X1    g152(.A(KEYINPUT66), .ZN(new_n354));
  NAND2_X1  g153(.A1(new_n353), .A2(new_n354), .ZN(new_n355));
  NAND3_X1  g154(.A1(new_n355), .A2(new_n321), .A3(new_n305), .ZN(new_n356));
  NOR2_X1   g155(.A1(new_n341), .A2(new_n342), .ZN(new_n357));
  AOI21_X1  g156(.A(new_n346), .B1(new_n357), .B2(G113gat), .ZN(new_n358));
  NOR4_X1   g157(.A1(new_n341), .A2(new_n342), .A3(KEYINPUT74), .A4(new_n343), .ZN(new_n359));
  OAI21_X1  g158(.A(new_n348), .B1(new_n358), .B2(new_n359), .ZN(new_n360));
  NAND3_X1  g159(.A1(new_n360), .A2(new_n350), .A3(new_n335), .ZN(new_n361));
  INV_X1    g160(.A(new_n331), .ZN(new_n362));
  NAND2_X1  g161(.A1(new_n361), .A2(new_n362), .ZN(new_n363));
  NAND3_X1  g162(.A1(new_n356), .A2(new_n363), .A3(new_n292), .ZN(new_n364));
  NAND4_X1  g163(.A1(new_n352), .A2(G227gat), .A3(G233gat), .A4(new_n364), .ZN(new_n365));
  AOI21_X1  g164(.A(new_n270), .B1(new_n365), .B2(KEYINPUT32), .ZN(new_n366));
  INV_X1    g165(.A(KEYINPUT33), .ZN(new_n367));
  NAND2_X1  g166(.A1(new_n365), .A2(new_n367), .ZN(new_n368));
  NAND2_X1  g167(.A1(new_n366), .A2(new_n368), .ZN(new_n369));
  OR2_X1    g168(.A1(new_n270), .A2(KEYINPUT76), .ZN(new_n370));
  NAND2_X1  g169(.A1(new_n270), .A2(KEYINPUT76), .ZN(new_n371));
  NAND3_X1  g170(.A1(new_n370), .A2(KEYINPUT33), .A3(new_n371), .ZN(new_n372));
  NAND3_X1  g171(.A1(new_n365), .A2(KEYINPUT32), .A3(new_n372), .ZN(new_n373));
  NAND2_X1  g172(.A1(new_n369), .A2(new_n373), .ZN(new_n374));
  NAND2_X1  g173(.A1(new_n352), .A2(new_n364), .ZN(new_n375));
  NAND2_X1  g174(.A1(G227gat), .A2(G233gat), .ZN(new_n376));
  NAND2_X1  g175(.A1(new_n375), .A2(new_n376), .ZN(new_n377));
  INV_X1    g176(.A(KEYINPUT34), .ZN(new_n378));
  INV_X1    g177(.A(KEYINPUT77), .ZN(new_n379));
  AOI21_X1  g178(.A(new_n378), .B1(new_n376), .B2(new_n379), .ZN(new_n380));
  OR2_X1    g179(.A1(new_n377), .A2(new_n380), .ZN(new_n381));
  NAND2_X1  g180(.A1(new_n377), .A2(new_n380), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n381), .A2(new_n382), .ZN(new_n383));
  NAND2_X1  g182(.A1(new_n374), .A2(new_n383), .ZN(new_n384));
  INV_X1    g183(.A(new_n384), .ZN(new_n385));
  NAND4_X1  g184(.A1(new_n369), .A2(new_n381), .A3(new_n373), .A4(new_n382), .ZN(new_n386));
  INV_X1    g185(.A(new_n386), .ZN(new_n387));
  NOR2_X1   g186(.A1(new_n385), .A2(new_n387), .ZN(new_n388));
  XNOR2_X1  g187(.A(KEYINPUT31), .B(G50gat), .ZN(new_n389));
  INV_X1    g188(.A(G106gat), .ZN(new_n390));
  XNOR2_X1  g189(.A(new_n389), .B(new_n390), .ZN(new_n391));
  NAND2_X1  g190(.A1(G228gat), .A2(G233gat), .ZN(new_n392));
  INV_X1    g191(.A(new_n392), .ZN(new_n393));
  NAND2_X1  g192(.A1(G211gat), .A2(G218gat), .ZN(new_n394));
  INV_X1    g193(.A(KEYINPUT22), .ZN(new_n395));
  NAND2_X1  g194(.A1(new_n394), .A2(new_n395), .ZN(new_n396));
  NAND2_X1  g195(.A1(new_n396), .A2(KEYINPUT78), .ZN(new_n397));
  INV_X1    g196(.A(KEYINPUT78), .ZN(new_n398));
  NAND3_X1  g197(.A1(new_n394), .A2(new_n398), .A3(new_n395), .ZN(new_n399));
  XNOR2_X1  g198(.A(G197gat), .B(G204gat), .ZN(new_n400));
  NAND3_X1  g199(.A1(new_n397), .A2(new_n399), .A3(new_n400), .ZN(new_n401));
  INV_X1    g200(.A(G211gat), .ZN(new_n402));
  INV_X1    g201(.A(G218gat), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n402), .A2(new_n403), .ZN(new_n404));
  NAND3_X1  g203(.A1(new_n404), .A2(KEYINPUT79), .A3(new_n394), .ZN(new_n405));
  INV_X1    g204(.A(new_n405), .ZN(new_n406));
  NAND2_X1  g205(.A1(new_n401), .A2(new_n406), .ZN(new_n407));
  NAND4_X1  g206(.A1(new_n405), .A2(new_n397), .A3(new_n399), .A4(new_n400), .ZN(new_n408));
  NAND2_X1  g207(.A1(new_n407), .A2(new_n408), .ZN(new_n409));
  INV_X1    g208(.A(KEYINPUT3), .ZN(new_n410));
  NAND2_X1  g209(.A1(G155gat), .A2(G162gat), .ZN(new_n411));
  NAND2_X1  g210(.A1(new_n411), .A2(KEYINPUT2), .ZN(new_n412));
  OR2_X1    g211(.A1(G141gat), .A2(G148gat), .ZN(new_n413));
  NAND2_X1  g212(.A1(G141gat), .A2(G148gat), .ZN(new_n414));
  NAND3_X1  g213(.A1(new_n412), .A2(new_n413), .A3(new_n414), .ZN(new_n415));
  INV_X1    g214(.A(KEYINPUT81), .ZN(new_n416));
  XNOR2_X1  g215(.A(G155gat), .B(G162gat), .ZN(new_n417));
  AND3_X1   g216(.A1(new_n415), .A2(new_n416), .A3(new_n417), .ZN(new_n418));
  AOI21_X1  g217(.A(new_n417), .B1(new_n415), .B2(new_n416), .ZN(new_n419));
  OAI21_X1  g218(.A(new_n410), .B1(new_n418), .B2(new_n419), .ZN(new_n420));
  INV_X1    g219(.A(KEYINPUT83), .ZN(new_n421));
  NAND2_X1  g220(.A1(new_n420), .A2(new_n421), .ZN(new_n422));
  XNOR2_X1  g221(.A(G141gat), .B(G148gat), .ZN(new_n423));
  INV_X1    g222(.A(KEYINPUT2), .ZN(new_n424));
  AOI21_X1  g223(.A(new_n424), .B1(G155gat), .B2(G162gat), .ZN(new_n425));
  OAI21_X1  g224(.A(new_n416), .B1(new_n423), .B2(new_n425), .ZN(new_n426));
  INV_X1    g225(.A(new_n417), .ZN(new_n427));
  NAND2_X1  g226(.A1(new_n426), .A2(new_n427), .ZN(new_n428));
  NAND3_X1  g227(.A1(new_n415), .A2(new_n416), .A3(new_n417), .ZN(new_n429));
  NAND2_X1  g228(.A1(new_n428), .A2(new_n429), .ZN(new_n430));
  NAND3_X1  g229(.A1(new_n430), .A2(KEYINPUT83), .A3(new_n410), .ZN(new_n431));
  NAND2_X1  g230(.A1(new_n422), .A2(new_n431), .ZN(new_n432));
  INV_X1    g231(.A(KEYINPUT29), .ZN(new_n433));
  AOI21_X1  g232(.A(new_n409), .B1(new_n432), .B2(new_n433), .ZN(new_n434));
  NAND2_X1  g233(.A1(new_n409), .A2(new_n433), .ZN(new_n435));
  AOI21_X1  g234(.A(new_n430), .B1(new_n435), .B2(new_n410), .ZN(new_n436));
  OAI21_X1  g235(.A(new_n393), .B1(new_n434), .B2(new_n436), .ZN(new_n437));
  NAND2_X1  g236(.A1(new_n404), .A2(new_n394), .ZN(new_n438));
  NAND2_X1  g237(.A1(new_n401), .A2(new_n438), .ZN(new_n439));
  NAND2_X1  g238(.A1(new_n439), .A2(new_n433), .ZN(new_n440));
  NOR2_X1   g239(.A1(new_n401), .A2(new_n438), .ZN(new_n441));
  OAI21_X1  g240(.A(new_n410), .B1(new_n440), .B2(new_n441), .ZN(new_n442));
  INV_X1    g241(.A(new_n430), .ZN(new_n443));
  AOI21_X1  g242(.A(new_n393), .B1(new_n442), .B2(new_n443), .ZN(new_n444));
  AOI21_X1  g243(.A(KEYINPUT29), .B1(new_n422), .B2(new_n431), .ZN(new_n445));
  OAI21_X1  g244(.A(new_n444), .B1(new_n445), .B2(new_n409), .ZN(new_n446));
  NAND2_X1  g245(.A1(new_n437), .A2(new_n446), .ZN(new_n447));
  NAND2_X1  g246(.A1(new_n447), .A2(G22gat), .ZN(new_n448));
  INV_X1    g247(.A(KEYINPUT85), .ZN(new_n449));
  INV_X1    g248(.A(G78gat), .ZN(new_n450));
  INV_X1    g249(.A(G22gat), .ZN(new_n451));
  AOI21_X1  g250(.A(KEYINPUT83), .B1(new_n430), .B2(new_n410), .ZN(new_n452));
  AOI211_X1 g251(.A(new_n421), .B(KEYINPUT3), .C1(new_n428), .C2(new_n429), .ZN(new_n453));
  OAI21_X1  g252(.A(new_n433), .B1(new_n452), .B2(new_n453), .ZN(new_n454));
  INV_X1    g253(.A(new_n409), .ZN(new_n455));
  AOI21_X1  g254(.A(new_n436), .B1(new_n454), .B2(new_n455), .ZN(new_n456));
  OAI211_X1 g255(.A(new_n451), .B(new_n446), .C1(new_n456), .C2(new_n392), .ZN(new_n457));
  NAND4_X1  g256(.A1(new_n448), .A2(new_n449), .A3(new_n450), .A4(new_n457), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n457), .A2(new_n449), .ZN(new_n459));
  AOI21_X1  g258(.A(new_n451), .B1(new_n437), .B2(new_n446), .ZN(new_n460));
  OAI21_X1  g259(.A(G78gat), .B1(new_n459), .B2(new_n460), .ZN(new_n461));
  AOI21_X1  g260(.A(new_n391), .B1(new_n458), .B2(new_n461), .ZN(new_n462));
  INV_X1    g261(.A(new_n462), .ZN(new_n463));
  NAND3_X1  g262(.A1(new_n458), .A2(new_n461), .A3(new_n391), .ZN(new_n464));
  NAND2_X1  g263(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  NAND2_X1  g264(.A1(new_n388), .A2(new_n465), .ZN(new_n466));
  INV_X1    g265(.A(KEYINPUT5), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n363), .A2(KEYINPUT82), .ZN(new_n468));
  INV_X1    g267(.A(KEYINPUT82), .ZN(new_n469));
  NAND2_X1  g268(.A1(new_n351), .A2(new_n469), .ZN(new_n470));
  NAND3_X1  g269(.A1(new_n468), .A2(new_n470), .A3(new_n443), .ZN(new_n471));
  NAND3_X1  g270(.A1(new_n361), .A2(new_n430), .A3(new_n362), .ZN(new_n472));
  NAND2_X1  g271(.A1(new_n471), .A2(new_n472), .ZN(new_n473));
  NAND2_X1  g272(.A1(G225gat), .A2(G233gat), .ZN(new_n474));
  INV_X1    g273(.A(new_n474), .ZN(new_n475));
  AOI21_X1  g274(.A(new_n467), .B1(new_n473), .B2(new_n475), .ZN(new_n476));
  NOR3_X1   g275(.A1(new_n418), .A2(new_n419), .A3(new_n410), .ZN(new_n477));
  AOI21_X1  g276(.A(new_n477), .B1(new_n422), .B2(new_n431), .ZN(new_n478));
  NAND3_X1  g277(.A1(new_n478), .A2(new_n468), .A3(new_n470), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n472), .A2(KEYINPUT4), .ZN(new_n480));
  INV_X1    g279(.A(KEYINPUT4), .ZN(new_n481));
  NAND3_X1  g280(.A1(new_n351), .A2(new_n481), .A3(new_n430), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n480), .A2(new_n482), .ZN(new_n483));
  NAND3_X1  g282(.A1(new_n479), .A2(new_n483), .A3(new_n474), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n484), .A2(KEYINPUT84), .ZN(new_n485));
  NAND2_X1  g284(.A1(new_n476), .A2(new_n485), .ZN(new_n486));
  AOI21_X1  g285(.A(new_n474), .B1(new_n471), .B2(new_n472), .ZN(new_n487));
  OAI211_X1 g286(.A(KEYINPUT84), .B(new_n484), .C1(new_n487), .C2(new_n467), .ZN(new_n488));
  XNOR2_X1  g287(.A(G1gat), .B(G29gat), .ZN(new_n489));
  XNOR2_X1  g288(.A(new_n489), .B(KEYINPUT0), .ZN(new_n490));
  XNOR2_X1  g289(.A(G57gat), .B(G85gat), .ZN(new_n491));
  XOR2_X1   g290(.A(new_n490), .B(new_n491), .Z(new_n492));
  INV_X1    g291(.A(new_n492), .ZN(new_n493));
  NAND3_X1  g292(.A1(new_n486), .A2(new_n488), .A3(new_n493), .ZN(new_n494));
  INV_X1    g293(.A(KEYINPUT6), .ZN(new_n495));
  NOR2_X1   g294(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  INV_X1    g295(.A(KEYINPUT87), .ZN(new_n497));
  AND3_X1   g296(.A1(new_n486), .A2(new_n497), .A3(new_n488), .ZN(new_n498));
  AOI21_X1  g297(.A(new_n497), .B1(new_n486), .B2(new_n488), .ZN(new_n499));
  OAI21_X1  g298(.A(new_n493), .B1(new_n498), .B2(new_n499), .ZN(new_n500));
  NAND2_X1  g299(.A1(new_n486), .A2(new_n488), .ZN(new_n501));
  AOI21_X1  g300(.A(KEYINPUT6), .B1(new_n501), .B2(new_n492), .ZN(new_n502));
  AOI21_X1  g301(.A(new_n496), .B1(new_n500), .B2(new_n502), .ZN(new_n503));
  NOR2_X1   g302(.A1(new_n466), .A2(new_n503), .ZN(new_n504));
  XNOR2_X1  g303(.A(G8gat), .B(G36gat), .ZN(new_n505));
  XNOR2_X1  g304(.A(G64gat), .B(G92gat), .ZN(new_n506));
  XOR2_X1   g305(.A(new_n505), .B(new_n506), .Z(new_n507));
  INV_X1    g306(.A(new_n507), .ZN(new_n508));
  NAND2_X1  g307(.A1(new_n323), .A2(KEYINPUT80), .ZN(new_n509));
  AND2_X1   g308(.A1(G226gat), .A2(G233gat), .ZN(new_n510));
  INV_X1    g309(.A(KEYINPUT80), .ZN(new_n511));
  OAI211_X1 g310(.A(new_n511), .B(new_n292), .C1(new_n315), .C2(new_n322), .ZN(new_n512));
  NAND3_X1  g311(.A1(new_n509), .A2(new_n510), .A3(new_n512), .ZN(new_n513));
  NOR2_X1   g312(.A1(new_n510), .A2(KEYINPUT29), .ZN(new_n514));
  NAND2_X1  g313(.A1(new_n323), .A2(new_n514), .ZN(new_n515));
  NAND3_X1  g314(.A1(new_n513), .A2(new_n515), .A3(new_n455), .ZN(new_n516));
  INV_X1    g315(.A(new_n516), .ZN(new_n517));
  INV_X1    g316(.A(new_n512), .ZN(new_n518));
  AOI21_X1  g317(.A(new_n511), .B1(new_n356), .B2(new_n292), .ZN(new_n519));
  OAI21_X1  g318(.A(new_n514), .B1(new_n518), .B2(new_n519), .ZN(new_n520));
  NAND3_X1  g319(.A1(new_n356), .A2(new_n510), .A3(new_n292), .ZN(new_n521));
  AOI21_X1  g320(.A(new_n455), .B1(new_n520), .B2(new_n521), .ZN(new_n522));
  OAI21_X1  g321(.A(new_n508), .B1(new_n517), .B2(new_n522), .ZN(new_n523));
  INV_X1    g322(.A(new_n521), .ZN(new_n524));
  NAND2_X1  g323(.A1(new_n509), .A2(new_n512), .ZN(new_n525));
  AOI21_X1  g324(.A(new_n524), .B1(new_n525), .B2(new_n514), .ZN(new_n526));
  OAI211_X1 g325(.A(new_n516), .B(new_n507), .C1(new_n526), .C2(new_n455), .ZN(new_n527));
  NAND3_X1  g326(.A1(new_n523), .A2(KEYINPUT30), .A3(new_n527), .ZN(new_n528));
  INV_X1    g327(.A(new_n522), .ZN(new_n529));
  INV_X1    g328(.A(KEYINPUT30), .ZN(new_n530));
  NAND4_X1  g329(.A1(new_n529), .A2(new_n530), .A3(new_n516), .A4(new_n507), .ZN(new_n531));
  AND2_X1   g330(.A1(new_n528), .A2(new_n531), .ZN(new_n532));
  NOR2_X1   g331(.A1(new_n532), .A2(KEYINPUT35), .ZN(new_n533));
  NAND2_X1  g332(.A1(new_n504), .A2(new_n533), .ZN(new_n534));
  AND3_X1   g333(.A1(new_n458), .A2(new_n461), .A3(new_n391), .ZN(new_n535));
  NOR2_X1   g334(.A1(new_n535), .A2(new_n462), .ZN(new_n536));
  NOR3_X1   g335(.A1(new_n536), .A2(new_n387), .A3(new_n385), .ZN(new_n537));
  NAND2_X1  g336(.A1(new_n502), .A2(new_n494), .ZN(new_n538));
  INV_X1    g337(.A(new_n496), .ZN(new_n539));
  AOI22_X1  g338(.A1(new_n538), .A2(new_n539), .B1(new_n528), .B2(new_n531), .ZN(new_n540));
  NAND2_X1  g339(.A1(new_n537), .A2(new_n540), .ZN(new_n541));
  NAND2_X1  g340(.A1(new_n541), .A2(KEYINPUT35), .ZN(new_n542));
  NAND2_X1  g341(.A1(new_n534), .A2(new_n542), .ZN(new_n543));
  AND3_X1   g342(.A1(new_n384), .A2(KEYINPUT36), .A3(new_n386), .ZN(new_n544));
  AOI21_X1  g343(.A(KEYINPUT36), .B1(new_n384), .B2(new_n386), .ZN(new_n545));
  OR2_X1    g344(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  NAND2_X1  g345(.A1(new_n501), .A2(KEYINPUT87), .ZN(new_n547));
  NAND3_X1  g346(.A1(new_n486), .A2(new_n497), .A3(new_n488), .ZN(new_n548));
  AOI21_X1  g347(.A(new_n492), .B1(new_n547), .B2(new_n548), .ZN(new_n549));
  NAND2_X1  g348(.A1(new_n501), .A2(new_n492), .ZN(new_n550));
  NAND2_X1  g349(.A1(new_n550), .A2(new_n495), .ZN(new_n551));
  OAI211_X1 g350(.A(new_n539), .B(new_n527), .C1(new_n549), .C2(new_n551), .ZN(new_n552));
  INV_X1    g351(.A(KEYINPUT37), .ZN(new_n553));
  NOR2_X1   g352(.A1(new_n507), .A2(new_n553), .ZN(new_n554));
  INV_X1    g353(.A(new_n554), .ZN(new_n555));
  NAND2_X1  g354(.A1(new_n523), .A2(new_n555), .ZN(new_n556));
  INV_X1    g355(.A(KEYINPUT38), .ZN(new_n557));
  INV_X1    g356(.A(KEYINPUT88), .ZN(new_n558));
  NAND3_X1  g357(.A1(new_n526), .A2(new_n558), .A3(new_n455), .ZN(new_n559));
  NAND3_X1  g358(.A1(new_n520), .A2(new_n455), .A3(new_n521), .ZN(new_n560));
  NAND2_X1  g359(.A1(new_n560), .A2(KEYINPUT88), .ZN(new_n561));
  AOI21_X1  g360(.A(new_n455), .B1(new_n513), .B2(new_n515), .ZN(new_n562));
  OAI211_X1 g361(.A(KEYINPUT37), .B(new_n559), .C1(new_n561), .C2(new_n562), .ZN(new_n563));
  NAND3_X1  g362(.A1(new_n556), .A2(new_n557), .A3(new_n563), .ZN(new_n564));
  OAI21_X1  g363(.A(new_n516), .B1(new_n526), .B2(new_n455), .ZN(new_n565));
  AOI21_X1  g364(.A(new_n554), .B1(new_n565), .B2(new_n508), .ZN(new_n566));
  AOI21_X1  g365(.A(new_n553), .B1(new_n529), .B2(new_n516), .ZN(new_n567));
  OAI21_X1  g366(.A(KEYINPUT38), .B1(new_n566), .B2(new_n567), .ZN(new_n568));
  NAND2_X1  g367(.A1(new_n564), .A2(new_n568), .ZN(new_n569));
  NOR2_X1   g368(.A1(new_n552), .A2(new_n569), .ZN(new_n570));
  AOI21_X1  g369(.A(new_n474), .B1(new_n479), .B2(new_n483), .ZN(new_n571));
  INV_X1    g370(.A(KEYINPUT39), .ZN(new_n572));
  AOI21_X1  g371(.A(new_n493), .B1(new_n571), .B2(new_n572), .ZN(new_n573));
  NAND3_X1  g372(.A1(new_n471), .A2(new_n474), .A3(new_n472), .ZN(new_n574));
  AOI211_X1 g373(.A(KEYINPUT82), .B(new_n331), .C1(new_n349), .C2(new_n350), .ZN(new_n575));
  AOI21_X1  g374(.A(new_n469), .B1(new_n361), .B2(new_n362), .ZN(new_n576));
  NOR2_X1   g375(.A1(new_n575), .A2(new_n576), .ZN(new_n577));
  AOI22_X1  g376(.A1(new_n577), .A2(new_n478), .B1(new_n480), .B2(new_n482), .ZN(new_n578));
  OAI211_X1 g377(.A(KEYINPUT39), .B(new_n574), .C1(new_n578), .C2(new_n474), .ZN(new_n579));
  NAND2_X1  g378(.A1(new_n573), .A2(new_n579), .ZN(new_n580));
  INV_X1    g379(.A(KEYINPUT86), .ZN(new_n581));
  NAND2_X1  g380(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  INV_X1    g381(.A(KEYINPUT40), .ZN(new_n583));
  NAND2_X1  g382(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  NAND3_X1  g383(.A1(new_n580), .A2(new_n581), .A3(KEYINPUT40), .ZN(new_n585));
  NAND2_X1  g384(.A1(new_n584), .A2(new_n585), .ZN(new_n586));
  NAND2_X1  g385(.A1(new_n586), .A2(new_n500), .ZN(new_n587));
  NAND2_X1  g386(.A1(new_n528), .A2(new_n531), .ZN(new_n588));
  OAI21_X1  g387(.A(new_n465), .B1(new_n587), .B2(new_n588), .ZN(new_n589));
  OAI221_X1 g388(.A(new_n546), .B1(new_n540), .B2(new_n465), .C1(new_n570), .C2(new_n589), .ZN(new_n590));
  AOI21_X1  g389(.A(new_n267), .B1(new_n543), .B2(new_n590), .ZN(new_n591));
  INV_X1    g390(.A(G57gat), .ZN(new_n592));
  NAND2_X1  g391(.A1(new_n592), .A2(G64gat), .ZN(new_n593));
  INV_X1    g392(.A(G64gat), .ZN(new_n594));
  NAND2_X1  g393(.A1(new_n594), .A2(G57gat), .ZN(new_n595));
  INV_X1    g394(.A(KEYINPUT9), .ZN(new_n596));
  NAND2_X1  g395(.A1(G71gat), .A2(G78gat), .ZN(new_n597));
  AOI22_X1  g396(.A1(new_n593), .A2(new_n595), .B1(new_n596), .B2(new_n597), .ZN(new_n598));
  XNOR2_X1  g397(.A(G71gat), .B(G78gat), .ZN(new_n599));
  NAND2_X1  g398(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  INV_X1    g399(.A(KEYINPUT94), .ZN(new_n601));
  NAND2_X1  g400(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  NAND3_X1  g401(.A1(new_n598), .A2(KEYINPUT94), .A3(new_n599), .ZN(new_n603));
  NAND2_X1  g402(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  OR3_X1    g403(.A1(KEYINPUT93), .A2(G71gat), .A3(G78gat), .ZN(new_n605));
  OAI21_X1  g404(.A(KEYINPUT93), .B1(G71gat), .B2(G78gat), .ZN(new_n606));
  NAND2_X1  g405(.A1(new_n605), .A2(new_n606), .ZN(new_n607));
  AND2_X1   g406(.A1(new_n593), .A2(new_n595), .ZN(new_n608));
  OAI211_X1 g407(.A(new_n607), .B(new_n597), .C1(new_n608), .C2(new_n596), .ZN(new_n609));
  AOI21_X1  g408(.A(KEYINPUT21), .B1(new_n604), .B2(new_n609), .ZN(new_n610));
  XOR2_X1   g409(.A(new_n610), .B(KEYINPUT95), .Z(new_n611));
  NAND2_X1  g410(.A1(new_n611), .A2(KEYINPUT96), .ZN(new_n612));
  XNOR2_X1  g411(.A(new_n610), .B(KEYINPUT95), .ZN(new_n613));
  INV_X1    g412(.A(KEYINPUT96), .ZN(new_n614));
  NAND2_X1  g413(.A1(new_n613), .A2(new_n614), .ZN(new_n615));
  NAND2_X1  g414(.A1(new_n612), .A2(new_n615), .ZN(new_n616));
  XOR2_X1   g415(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n617));
  NAND2_X1  g416(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  INV_X1    g417(.A(new_n617), .ZN(new_n619));
  NAND3_X1  g418(.A1(new_n612), .A2(new_n615), .A3(new_n619), .ZN(new_n620));
  NAND2_X1  g419(.A1(new_n618), .A2(new_n620), .ZN(new_n621));
  XOR2_X1   g420(.A(G183gat), .B(G211gat), .Z(new_n622));
  NAND2_X1  g421(.A1(new_n621), .A2(new_n622), .ZN(new_n623));
  INV_X1    g422(.A(new_n622), .ZN(new_n624));
  NAND3_X1  g423(.A1(new_n618), .A2(new_n624), .A3(new_n620), .ZN(new_n625));
  NAND2_X1  g424(.A1(new_n623), .A2(new_n625), .ZN(new_n626));
  NAND3_X1  g425(.A1(new_n604), .A2(KEYINPUT21), .A3(new_n609), .ZN(new_n627));
  NAND2_X1  g426(.A1(new_n627), .A2(new_n237), .ZN(new_n628));
  XNOR2_X1  g427(.A(new_n628), .B(KEYINPUT97), .ZN(new_n629));
  XNOR2_X1  g428(.A(G127gat), .B(G155gat), .ZN(new_n630));
  NAND2_X1  g429(.A1(G231gat), .A2(G233gat), .ZN(new_n631));
  XNOR2_X1  g430(.A(new_n630), .B(new_n631), .ZN(new_n632));
  XNOR2_X1  g431(.A(new_n629), .B(new_n632), .ZN(new_n633));
  INV_X1    g432(.A(new_n633), .ZN(new_n634));
  NAND2_X1  g433(.A1(new_n626), .A2(new_n634), .ZN(new_n635));
  NAND3_X1  g434(.A1(new_n623), .A2(new_n625), .A3(new_n633), .ZN(new_n636));
  NAND2_X1  g435(.A1(new_n635), .A2(new_n636), .ZN(new_n637));
  NAND2_X1  g436(.A1(new_n225), .A2(new_n226), .ZN(new_n638));
  NAND2_X1  g437(.A1(G85gat), .A2(G92gat), .ZN(new_n639));
  NAND2_X1  g438(.A1(new_n639), .A2(KEYINPUT7), .ZN(new_n640));
  INV_X1    g439(.A(KEYINPUT7), .ZN(new_n641));
  NAND3_X1  g440(.A1(new_n641), .A2(G85gat), .A3(G92gat), .ZN(new_n642));
  NAND2_X1  g441(.A1(new_n640), .A2(new_n642), .ZN(new_n643));
  XNOR2_X1  g442(.A(G99gat), .B(G106gat), .ZN(new_n644));
  NAND2_X1  g443(.A1(G99gat), .A2(G106gat), .ZN(new_n645));
  INV_X1    g444(.A(G85gat), .ZN(new_n646));
  INV_X1    g445(.A(G92gat), .ZN(new_n647));
  AOI22_X1  g446(.A1(KEYINPUT8), .A2(new_n645), .B1(new_n646), .B2(new_n647), .ZN(new_n648));
  AND3_X1   g447(.A1(new_n643), .A2(new_n644), .A3(new_n648), .ZN(new_n649));
  AOI21_X1  g448(.A(new_n644), .B1(new_n643), .B2(new_n648), .ZN(new_n650));
  NOR2_X1   g449(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  AND2_X1   g450(.A1(G232gat), .A2(G233gat), .ZN(new_n652));
  AOI22_X1  g451(.A1(new_n638), .A2(new_n651), .B1(KEYINPUT41), .B2(new_n652), .ZN(new_n653));
  INV_X1    g452(.A(new_n651), .ZN(new_n654));
  NAND3_X1  g453(.A1(new_n254), .A2(new_n248), .A3(new_n654), .ZN(new_n655));
  XOR2_X1   g454(.A(G190gat), .B(G218gat), .Z(new_n656));
  INV_X1    g455(.A(new_n656), .ZN(new_n657));
  NAND3_X1  g456(.A1(new_n653), .A2(new_n655), .A3(new_n657), .ZN(new_n658));
  INV_X1    g457(.A(new_n658), .ZN(new_n659));
  AOI21_X1  g458(.A(new_n657), .B1(new_n653), .B2(new_n655), .ZN(new_n660));
  NOR2_X1   g459(.A1(new_n652), .A2(KEYINPUT41), .ZN(new_n661));
  XNOR2_X1  g460(.A(G134gat), .B(G162gat), .ZN(new_n662));
  XNOR2_X1  g461(.A(new_n661), .B(new_n662), .ZN(new_n663));
  INV_X1    g462(.A(new_n663), .ZN(new_n664));
  NOR3_X1   g463(.A1(new_n659), .A2(new_n660), .A3(new_n664), .ZN(new_n665));
  NAND2_X1  g464(.A1(new_n653), .A2(new_n655), .ZN(new_n666));
  NAND2_X1  g465(.A1(new_n666), .A2(new_n656), .ZN(new_n667));
  AOI21_X1  g466(.A(new_n663), .B1(new_n667), .B2(new_n658), .ZN(new_n668));
  NOR2_X1   g467(.A1(new_n665), .A2(new_n668), .ZN(new_n669));
  INV_X1    g468(.A(G230gat), .ZN(new_n670));
  INV_X1    g469(.A(G233gat), .ZN(new_n671));
  NOR2_X1   g470(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  OR2_X1    g471(.A1(new_n644), .A2(KEYINPUT98), .ZN(new_n673));
  AND3_X1   g472(.A1(new_n598), .A2(KEYINPUT94), .A3(new_n599), .ZN(new_n674));
  AOI21_X1  g473(.A(KEYINPUT94), .B1(new_n598), .B2(new_n599), .ZN(new_n675));
  OAI211_X1 g474(.A(new_n609), .B(new_n673), .C1(new_n674), .C2(new_n675), .ZN(new_n676));
  NAND2_X1  g475(.A1(new_n676), .A2(new_n654), .ZN(new_n677));
  NAND4_X1  g476(.A1(new_n604), .A2(new_n609), .A3(new_n651), .A4(new_n673), .ZN(new_n678));
  INV_X1    g477(.A(KEYINPUT10), .ZN(new_n679));
  NAND3_X1  g478(.A1(new_n677), .A2(new_n678), .A3(new_n679), .ZN(new_n680));
  NAND4_X1  g479(.A1(new_n604), .A2(KEYINPUT10), .A3(new_n651), .A4(new_n609), .ZN(new_n681));
  AOI21_X1  g480(.A(new_n672), .B1(new_n680), .B2(new_n681), .ZN(new_n682));
  INV_X1    g481(.A(new_n682), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n677), .A2(new_n678), .ZN(new_n684));
  NAND2_X1  g483(.A1(new_n684), .A2(new_n672), .ZN(new_n685));
  NAND2_X1  g484(.A1(new_n683), .A2(new_n685), .ZN(new_n686));
  XNOR2_X1  g485(.A(G120gat), .B(G148gat), .ZN(new_n687));
  XNOR2_X1  g486(.A(G176gat), .B(G204gat), .ZN(new_n688));
  XOR2_X1   g487(.A(new_n687), .B(new_n688), .Z(new_n689));
  INV_X1    g488(.A(new_n689), .ZN(new_n690));
  NAND2_X1  g489(.A1(new_n686), .A2(new_n690), .ZN(new_n691));
  NAND3_X1  g490(.A1(new_n683), .A2(new_n685), .A3(new_n689), .ZN(new_n692));
  NAND2_X1  g491(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  NOR3_X1   g492(.A1(new_n637), .A2(new_n669), .A3(new_n693), .ZN(new_n694));
  NAND2_X1  g493(.A1(new_n591), .A2(new_n694), .ZN(new_n695));
  AOI21_X1  g494(.A(new_n496), .B1(new_n494), .B2(new_n502), .ZN(new_n696));
  INV_X1    g495(.A(new_n696), .ZN(new_n697));
  NOR2_X1   g496(.A1(new_n695), .A2(new_n697), .ZN(new_n698));
  XOR2_X1   g497(.A(KEYINPUT99), .B(G1gat), .Z(new_n699));
  XNOR2_X1  g498(.A(new_n698), .B(new_n699), .ZN(G1324gat));
  INV_X1    g499(.A(new_n695), .ZN(new_n701));
  XOR2_X1   g500(.A(KEYINPUT16), .B(G8gat), .Z(new_n702));
  NAND3_X1  g501(.A1(new_n701), .A2(new_n532), .A3(new_n702), .ZN(new_n703));
  NAND2_X1  g502(.A1(new_n703), .A2(KEYINPUT100), .ZN(new_n704));
  OR2_X1    g503(.A1(new_n704), .A2(KEYINPUT42), .ZN(new_n705));
  OAI21_X1  g504(.A(G8gat), .B1(new_n695), .B2(new_n588), .ZN(new_n706));
  NAND2_X1  g505(.A1(new_n704), .A2(KEYINPUT42), .ZN(new_n707));
  NAND3_X1  g506(.A1(new_n705), .A2(new_n706), .A3(new_n707), .ZN(G1325gat));
  OAI21_X1  g507(.A(G15gat), .B1(new_n695), .B2(new_n546), .ZN(new_n709));
  INV_X1    g508(.A(G15gat), .ZN(new_n710));
  NAND2_X1  g509(.A1(new_n388), .A2(new_n710), .ZN(new_n711));
  OAI21_X1  g510(.A(new_n709), .B1(new_n695), .B2(new_n711), .ZN(G1326gat));
  NOR2_X1   g511(.A1(new_n695), .A2(new_n465), .ZN(new_n713));
  XOR2_X1   g512(.A(KEYINPUT43), .B(G22gat), .Z(new_n714));
  XNOR2_X1  g513(.A(new_n713), .B(new_n714), .ZN(G1327gat));
  INV_X1    g514(.A(new_n637), .ZN(new_n716));
  NOR2_X1   g515(.A1(new_n716), .A2(new_n693), .ZN(new_n717));
  INV_X1    g516(.A(new_n717), .ZN(new_n718));
  INV_X1    g517(.A(new_n669), .ZN(new_n719));
  NOR2_X1   g518(.A1(new_n718), .A2(new_n719), .ZN(new_n720));
  NAND4_X1  g519(.A1(new_n591), .A2(new_n210), .A3(new_n696), .A4(new_n720), .ZN(new_n721));
  OR2_X1    g520(.A1(new_n721), .A2(KEYINPUT101), .ZN(new_n722));
  NAND2_X1  g521(.A1(new_n721), .A2(KEYINPUT101), .ZN(new_n723));
  AND3_X1   g522(.A1(new_n722), .A2(KEYINPUT45), .A3(new_n723), .ZN(new_n724));
  AOI21_X1  g523(.A(KEYINPUT45), .B1(new_n722), .B2(new_n723), .ZN(new_n725));
  NOR2_X1   g524(.A1(new_n724), .A2(new_n725), .ZN(new_n726));
  OAI21_X1  g525(.A(new_n546), .B1(new_n570), .B2(new_n589), .ZN(new_n727));
  OAI21_X1  g526(.A(KEYINPUT103), .B1(new_n540), .B2(new_n465), .ZN(new_n728));
  INV_X1    g527(.A(KEYINPUT103), .ZN(new_n729));
  OAI211_X1 g528(.A(new_n729), .B(new_n536), .C1(new_n532), .C2(new_n696), .ZN(new_n730));
  NAND2_X1  g529(.A1(new_n728), .A2(new_n730), .ZN(new_n731));
  OAI21_X1  g530(.A(KEYINPUT104), .B1(new_n727), .B2(new_n731), .ZN(new_n732));
  NOR2_X1   g531(.A1(new_n544), .A2(new_n545), .ZN(new_n733));
  NAND4_X1  g532(.A1(new_n503), .A2(new_n527), .A3(new_n564), .A4(new_n568), .ZN(new_n734));
  NAND2_X1  g533(.A1(new_n547), .A2(new_n548), .ZN(new_n735));
  AOI22_X1  g534(.A1(new_n735), .A2(new_n493), .B1(new_n584), .B2(new_n585), .ZN(new_n736));
  AOI21_X1  g535(.A(new_n536), .B1(new_n736), .B2(new_n532), .ZN(new_n737));
  AOI21_X1  g536(.A(new_n733), .B1(new_n734), .B2(new_n737), .ZN(new_n738));
  INV_X1    g537(.A(KEYINPUT104), .ZN(new_n739));
  NAND4_X1  g538(.A1(new_n738), .A2(new_n739), .A3(new_n728), .A4(new_n730), .ZN(new_n740));
  NAND2_X1  g539(.A1(new_n732), .A2(new_n740), .ZN(new_n741));
  NAND2_X1  g540(.A1(new_n741), .A2(new_n543), .ZN(new_n742));
  INV_X1    g541(.A(KEYINPUT105), .ZN(new_n743));
  OAI21_X1  g542(.A(new_n743), .B1(new_n665), .B2(new_n668), .ZN(new_n744));
  OAI21_X1  g543(.A(new_n664), .B1(new_n659), .B2(new_n660), .ZN(new_n745));
  NAND3_X1  g544(.A1(new_n667), .A2(new_n663), .A3(new_n658), .ZN(new_n746));
  NAND3_X1  g545(.A1(new_n745), .A2(new_n746), .A3(KEYINPUT105), .ZN(new_n747));
  NAND2_X1  g546(.A1(new_n744), .A2(new_n747), .ZN(new_n748));
  NOR2_X1   g547(.A1(new_n748), .A2(KEYINPUT44), .ZN(new_n749));
  NAND2_X1  g548(.A1(new_n742), .A2(new_n749), .ZN(new_n750));
  INV_X1    g549(.A(KEYINPUT44), .ZN(new_n751));
  NAND2_X1  g550(.A1(new_n543), .A2(new_n590), .ZN(new_n752));
  AOI21_X1  g551(.A(new_n751), .B1(new_n752), .B2(new_n669), .ZN(new_n753));
  INV_X1    g552(.A(new_n753), .ZN(new_n754));
  NAND2_X1  g553(.A1(new_n750), .A2(new_n754), .ZN(new_n755));
  INV_X1    g554(.A(KEYINPUT102), .ZN(new_n756));
  NAND2_X1  g555(.A1(new_n266), .A2(new_n756), .ZN(new_n757));
  NAND3_X1  g556(.A1(new_n264), .A2(KEYINPUT102), .A3(new_n265), .ZN(new_n758));
  NAND2_X1  g557(.A1(new_n757), .A2(new_n758), .ZN(new_n759));
  NOR2_X1   g558(.A1(new_n718), .A2(new_n759), .ZN(new_n760));
  NAND2_X1  g559(.A1(new_n755), .A2(new_n760), .ZN(new_n761));
  OAI21_X1  g560(.A(G29gat), .B1(new_n761), .B2(new_n697), .ZN(new_n762));
  NAND2_X1  g561(.A1(new_n726), .A2(new_n762), .ZN(G1328gat));
  OAI21_X1  g562(.A(G36gat), .B1(new_n761), .B2(new_n588), .ZN(new_n764));
  NAND2_X1  g563(.A1(new_n591), .A2(new_n720), .ZN(new_n765));
  NOR3_X1   g564(.A1(new_n765), .A2(G36gat), .A3(new_n588), .ZN(new_n766));
  INV_X1    g565(.A(KEYINPUT46), .ZN(new_n767));
  OAI21_X1  g566(.A(new_n766), .B1(KEYINPUT106), .B2(new_n767), .ZN(new_n768));
  XNOR2_X1  g567(.A(KEYINPUT106), .B(KEYINPUT46), .ZN(new_n769));
  OAI211_X1 g568(.A(new_n764), .B(new_n768), .C1(new_n766), .C2(new_n769), .ZN(G1329gat));
  INV_X1    g569(.A(new_n749), .ZN(new_n771));
  AOI21_X1  g570(.A(new_n771), .B1(new_n741), .B2(new_n543), .ZN(new_n772));
  OAI211_X1 g571(.A(new_n733), .B(new_n760), .C1(new_n772), .C2(new_n753), .ZN(new_n773));
  NAND2_X1  g572(.A1(new_n773), .A2(G43gat), .ZN(new_n774));
  INV_X1    g573(.A(KEYINPUT107), .ZN(new_n775));
  NAND2_X1  g574(.A1(new_n774), .A2(new_n775), .ZN(new_n776));
  NAND4_X1  g575(.A1(new_n591), .A2(new_n213), .A3(new_n388), .A4(new_n720), .ZN(new_n777));
  NAND2_X1  g576(.A1(new_n774), .A2(new_n777), .ZN(new_n778));
  INV_X1    g577(.A(KEYINPUT47), .ZN(new_n779));
  NAND3_X1  g578(.A1(new_n776), .A2(new_n778), .A3(new_n779), .ZN(new_n780));
  OAI211_X1 g579(.A(new_n774), .B(new_n777), .C1(new_n775), .C2(KEYINPUT47), .ZN(new_n781));
  NAND2_X1  g580(.A1(new_n780), .A2(new_n781), .ZN(G1330gat));
  NAND4_X1  g581(.A1(new_n755), .A2(G50gat), .A3(new_n536), .A4(new_n760), .ZN(new_n783));
  OAI21_X1  g582(.A(new_n214), .B1(new_n765), .B2(new_n465), .ZN(new_n784));
  NAND2_X1  g583(.A1(new_n783), .A2(new_n784), .ZN(new_n785));
  NAND2_X1  g584(.A1(new_n785), .A2(KEYINPUT48), .ZN(new_n786));
  INV_X1    g585(.A(KEYINPUT48), .ZN(new_n787));
  NAND3_X1  g586(.A1(new_n783), .A2(new_n787), .A3(new_n784), .ZN(new_n788));
  NAND2_X1  g587(.A1(new_n786), .A2(new_n788), .ZN(G1331gat));
  INV_X1    g588(.A(new_n759), .ZN(new_n790));
  NAND3_X1  g589(.A1(new_n716), .A2(new_n719), .A3(new_n693), .ZN(new_n791));
  AOI211_X1 g590(.A(new_n790), .B(new_n791), .C1(new_n741), .C2(new_n543), .ZN(new_n792));
  NAND2_X1  g591(.A1(new_n792), .A2(new_n696), .ZN(new_n793));
  XNOR2_X1  g592(.A(new_n793), .B(G57gat), .ZN(G1332gat));
  NAND2_X1  g593(.A1(new_n792), .A2(new_n532), .ZN(new_n795));
  OAI21_X1  g594(.A(new_n795), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n796));
  XOR2_X1   g595(.A(KEYINPUT49), .B(G64gat), .Z(new_n797));
  OAI21_X1  g596(.A(new_n796), .B1(new_n795), .B2(new_n797), .ZN(G1333gat));
  INV_X1    g597(.A(G71gat), .ZN(new_n799));
  NAND3_X1  g598(.A1(new_n792), .A2(new_n799), .A3(new_n388), .ZN(new_n800));
  AND2_X1   g599(.A1(new_n792), .A2(new_n733), .ZN(new_n801));
  OAI21_X1  g600(.A(new_n800), .B1(new_n801), .B2(new_n799), .ZN(new_n802));
  INV_X1    g601(.A(KEYINPUT50), .ZN(new_n803));
  NAND2_X1  g602(.A1(new_n802), .A2(new_n803), .ZN(new_n804));
  OAI211_X1 g603(.A(KEYINPUT50), .B(new_n800), .C1(new_n801), .C2(new_n799), .ZN(new_n805));
  NAND2_X1  g604(.A1(new_n804), .A2(new_n805), .ZN(G1334gat));
  NAND2_X1  g605(.A1(new_n792), .A2(new_n536), .ZN(new_n807));
  XNOR2_X1  g606(.A(new_n807), .B(G78gat), .ZN(G1335gat));
  INV_X1    g607(.A(new_n693), .ZN(new_n809));
  NOR3_X1   g608(.A1(new_n716), .A2(new_n809), .A3(new_n790), .ZN(new_n810));
  NAND2_X1  g609(.A1(new_n755), .A2(new_n810), .ZN(new_n811));
  OAI21_X1  g610(.A(G85gat), .B1(new_n811), .B2(new_n697), .ZN(new_n812));
  NAND3_X1  g611(.A1(new_n637), .A2(new_n669), .A3(new_n759), .ZN(new_n813));
  INV_X1    g612(.A(new_n813), .ZN(new_n814));
  NAND2_X1  g613(.A1(new_n742), .A2(new_n814), .ZN(new_n815));
  INV_X1    g614(.A(KEYINPUT51), .ZN(new_n816));
  NAND2_X1  g615(.A1(new_n815), .A2(new_n816), .ZN(new_n817));
  NAND3_X1  g616(.A1(new_n742), .A2(KEYINPUT51), .A3(new_n814), .ZN(new_n818));
  NAND2_X1  g617(.A1(new_n817), .A2(new_n818), .ZN(new_n819));
  INV_X1    g618(.A(new_n819), .ZN(new_n820));
  NAND3_X1  g619(.A1(new_n696), .A2(new_n646), .A3(new_n693), .ZN(new_n821));
  OAI21_X1  g620(.A(new_n812), .B1(new_n820), .B2(new_n821), .ZN(G1336gat));
  INV_X1    g621(.A(KEYINPUT52), .ZN(new_n823));
  OAI211_X1 g622(.A(new_n532), .B(new_n810), .C1(new_n772), .C2(new_n753), .ZN(new_n824));
  NAND2_X1  g623(.A1(new_n824), .A2(G92gat), .ZN(new_n825));
  NAND3_X1  g624(.A1(new_n532), .A2(new_n647), .A3(new_n693), .ZN(new_n826));
  OAI211_X1 g625(.A(new_n823), .B(new_n825), .C1(new_n820), .C2(new_n826), .ZN(new_n827));
  INV_X1    g626(.A(new_n825), .ZN(new_n828));
  AOI21_X1  g627(.A(new_n826), .B1(new_n817), .B2(new_n818), .ZN(new_n829));
  OAI21_X1  g628(.A(KEYINPUT52), .B1(new_n828), .B2(new_n829), .ZN(new_n830));
  NAND2_X1  g629(.A1(new_n827), .A2(new_n830), .ZN(G1337gat));
  OAI21_X1  g630(.A(G99gat), .B1(new_n811), .B2(new_n546), .ZN(new_n832));
  INV_X1    g631(.A(G99gat), .ZN(new_n833));
  NAND3_X1  g632(.A1(new_n388), .A2(new_n833), .A3(new_n693), .ZN(new_n834));
  OAI21_X1  g633(.A(new_n832), .B1(new_n820), .B2(new_n834), .ZN(G1338gat));
  NOR3_X1   g634(.A1(new_n465), .A2(G106gat), .A3(new_n809), .ZN(new_n836));
  NAND2_X1  g635(.A1(new_n819), .A2(new_n836), .ZN(new_n837));
  OAI211_X1 g636(.A(new_n536), .B(new_n810), .C1(new_n772), .C2(new_n753), .ZN(new_n838));
  NAND2_X1  g637(.A1(new_n838), .A2(G106gat), .ZN(new_n839));
  INV_X1    g638(.A(KEYINPUT53), .ZN(new_n840));
  NAND3_X1  g639(.A1(new_n837), .A2(new_n839), .A3(new_n840), .ZN(new_n841));
  XNOR2_X1  g640(.A(new_n836), .B(KEYINPUT108), .ZN(new_n842));
  AOI22_X1  g641(.A1(new_n819), .A2(new_n842), .B1(new_n838), .B2(G106gat), .ZN(new_n843));
  OAI21_X1  g642(.A(new_n841), .B1(new_n843), .B2(new_n840), .ZN(G1339gat));
  INV_X1    g643(.A(new_n748), .ZN(new_n845));
  INV_X1    g644(.A(new_n692), .ZN(new_n846));
  AND3_X1   g645(.A1(new_n680), .A2(new_n672), .A3(new_n681), .ZN(new_n847));
  INV_X1    g646(.A(KEYINPUT54), .ZN(new_n848));
  NOR3_X1   g647(.A1(new_n847), .A2(new_n682), .A3(new_n848), .ZN(new_n849));
  INV_X1    g648(.A(KEYINPUT109), .ZN(new_n850));
  AOI211_X1 g649(.A(KEYINPUT54), .B(new_n672), .C1(new_n680), .C2(new_n681), .ZN(new_n851));
  OAI21_X1  g650(.A(new_n850), .B1(new_n851), .B2(new_n689), .ZN(new_n852));
  NAND2_X1  g651(.A1(new_n682), .A2(new_n848), .ZN(new_n853));
  NAND3_X1  g652(.A1(new_n853), .A2(KEYINPUT109), .A3(new_n690), .ZN(new_n854));
  AOI21_X1  g653(.A(new_n849), .B1(new_n852), .B2(new_n854), .ZN(new_n855));
  AOI21_X1  g654(.A(new_n846), .B1(new_n855), .B2(KEYINPUT55), .ZN(new_n856));
  INV_X1    g655(.A(new_n849), .ZN(new_n857));
  NOR3_X1   g656(.A1(new_n851), .A2(new_n850), .A3(new_n689), .ZN(new_n858));
  AOI21_X1  g657(.A(KEYINPUT109), .B1(new_n853), .B2(new_n690), .ZN(new_n859));
  OAI21_X1  g658(.A(new_n857), .B1(new_n858), .B2(new_n859), .ZN(new_n860));
  INV_X1    g659(.A(KEYINPUT55), .ZN(new_n861));
  NAND2_X1  g660(.A1(new_n860), .A2(new_n861), .ZN(new_n862));
  NAND4_X1  g661(.A1(new_n757), .A2(new_n758), .A3(new_n856), .A4(new_n862), .ZN(new_n863));
  OAI21_X1  g662(.A(new_n240), .B1(new_n243), .B2(new_n249), .ZN(new_n864));
  NAND2_X1  g663(.A1(new_n864), .A2(new_n203), .ZN(new_n865));
  INV_X1    g664(.A(KEYINPUT110), .ZN(new_n866));
  NAND4_X1  g665(.A1(new_n238), .A2(new_n240), .A3(new_n866), .A4(new_n205), .ZN(new_n867));
  NAND3_X1  g666(.A1(new_n238), .A2(new_n240), .A3(new_n205), .ZN(new_n868));
  NAND2_X1  g667(.A1(new_n868), .A2(KEYINPUT110), .ZN(new_n869));
  NAND3_X1  g668(.A1(new_n865), .A2(new_n867), .A3(new_n869), .ZN(new_n870));
  NAND2_X1  g669(.A1(new_n870), .A2(new_n261), .ZN(new_n871));
  NAND3_X1  g670(.A1(new_n871), .A2(new_n265), .A3(new_n693), .ZN(new_n872));
  AOI21_X1  g671(.A(new_n845), .B1(new_n863), .B2(new_n872), .ZN(new_n873));
  AND2_X1   g672(.A1(new_n871), .A2(new_n265), .ZN(new_n874));
  NAND3_X1  g673(.A1(new_n874), .A2(new_n856), .A3(new_n862), .ZN(new_n875));
  NOR2_X1   g674(.A1(new_n875), .A2(new_n748), .ZN(new_n876));
  OAI21_X1  g675(.A(new_n637), .B1(new_n873), .B2(new_n876), .ZN(new_n877));
  NAND2_X1  g676(.A1(new_n694), .A2(new_n759), .ZN(new_n878));
  NAND2_X1  g677(.A1(new_n877), .A2(new_n878), .ZN(new_n879));
  NOR2_X1   g678(.A1(new_n466), .A2(new_n697), .ZN(new_n880));
  AND2_X1   g679(.A1(new_n879), .A2(new_n880), .ZN(new_n881));
  NAND2_X1  g680(.A1(new_n881), .A2(KEYINPUT112), .ZN(new_n882));
  NAND2_X1  g681(.A1(new_n879), .A2(new_n880), .ZN(new_n883));
  INV_X1    g682(.A(KEYINPUT112), .ZN(new_n884));
  NAND2_X1  g683(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  AOI21_X1  g684(.A(new_n532), .B1(new_n882), .B2(new_n885), .ZN(new_n886));
  AOI21_X1  g685(.A(G113gat), .B1(new_n886), .B2(new_n790), .ZN(new_n887));
  NAND3_X1  g686(.A1(new_n881), .A2(KEYINPUT111), .A3(new_n588), .ZN(new_n888));
  INV_X1    g687(.A(KEYINPUT111), .ZN(new_n889));
  OAI21_X1  g688(.A(new_n889), .B1(new_n883), .B2(new_n532), .ZN(new_n890));
  NAND2_X1  g689(.A1(new_n888), .A2(new_n890), .ZN(new_n891));
  NOR3_X1   g690(.A1(new_n891), .A2(new_n343), .A3(new_n267), .ZN(new_n892));
  NOR2_X1   g691(.A1(new_n887), .A2(new_n892), .ZN(G1340gat));
  OAI21_X1  g692(.A(G120gat), .B1(new_n891), .B2(new_n809), .ZN(new_n894));
  NAND3_X1  g693(.A1(new_n886), .A2(new_n357), .A3(new_n693), .ZN(new_n895));
  NAND2_X1  g694(.A1(new_n894), .A2(new_n895), .ZN(G1341gat));
  NAND4_X1  g695(.A1(new_n886), .A2(new_n326), .A3(new_n327), .A4(new_n716), .ZN(new_n897));
  NAND2_X1  g696(.A1(new_n326), .A2(new_n327), .ZN(new_n898));
  OAI21_X1  g697(.A(new_n898), .B1(new_n891), .B2(new_n637), .ZN(new_n899));
  NAND2_X1  g698(.A1(new_n897), .A2(new_n899), .ZN(G1342gat));
  NOR2_X1   g699(.A1(new_n532), .A2(new_n719), .ZN(new_n901));
  NAND2_X1  g700(.A1(new_n901), .A2(new_n324), .ZN(new_n902));
  AOI21_X1  g701(.A(new_n902), .B1(new_n882), .B2(new_n885), .ZN(new_n903));
  INV_X1    g702(.A(KEYINPUT56), .ZN(new_n904));
  NAND2_X1  g703(.A1(new_n903), .A2(new_n904), .ZN(new_n905));
  NAND3_X1  g704(.A1(new_n888), .A2(new_n669), .A3(new_n890), .ZN(new_n906));
  AND3_X1   g705(.A1(new_n906), .A2(KEYINPUT113), .A3(G134gat), .ZN(new_n907));
  AOI21_X1  g706(.A(KEYINPUT113), .B1(new_n906), .B2(G134gat), .ZN(new_n908));
  NOR2_X1   g707(.A1(new_n903), .A2(new_n904), .ZN(new_n909));
  NOR2_X1   g708(.A1(new_n909), .A2(KEYINPUT114), .ZN(new_n910));
  INV_X1    g709(.A(KEYINPUT114), .ZN(new_n911));
  NOR3_X1   g710(.A1(new_n903), .A2(new_n911), .A3(new_n904), .ZN(new_n912));
  OAI221_X1 g711(.A(new_n905), .B1(new_n907), .B2(new_n908), .C1(new_n910), .C2(new_n912), .ZN(G1343gat));
  INV_X1    g712(.A(KEYINPUT118), .ZN(new_n914));
  INV_X1    g713(.A(KEYINPUT58), .ZN(new_n915));
  NAND2_X1  g714(.A1(new_n546), .A2(new_n696), .ZN(new_n916));
  INV_X1    g715(.A(new_n916), .ZN(new_n917));
  NAND2_X1  g716(.A1(new_n917), .A2(new_n588), .ZN(new_n918));
  INV_X1    g717(.A(new_n918), .ZN(new_n919));
  INV_X1    g718(.A(KEYINPUT57), .ZN(new_n920));
  NOR2_X1   g719(.A1(new_n465), .A2(new_n920), .ZN(new_n921));
  INV_X1    g720(.A(new_n921), .ZN(new_n922));
  NOR4_X1   g721(.A1(new_n637), .A2(new_n790), .A3(new_n669), .A4(new_n693), .ZN(new_n923));
  NAND2_X1  g722(.A1(new_n250), .A2(new_n251), .ZN(new_n924));
  INV_X1    g723(.A(new_n241), .ZN(new_n925));
  AND4_X1   g724(.A1(new_n262), .A2(new_n924), .A3(new_n256), .A4(new_n925), .ZN(new_n926));
  AOI21_X1  g725(.A(new_n262), .B1(new_n252), .B2(new_n256), .ZN(new_n927));
  OAI22_X1  g726(.A1(new_n926), .A2(new_n927), .B1(new_n855), .B2(KEYINPUT55), .ZN(new_n928));
  OAI211_X1 g727(.A(KEYINPUT55), .B(new_n857), .C1(new_n858), .C2(new_n859), .ZN(new_n929));
  NAND2_X1  g728(.A1(new_n929), .A2(new_n692), .ZN(new_n930));
  OAI21_X1  g729(.A(new_n872), .B1(new_n928), .B2(new_n930), .ZN(new_n931));
  NAND2_X1  g730(.A1(new_n931), .A2(new_n719), .ZN(new_n932));
  INV_X1    g731(.A(KEYINPUT115), .ZN(new_n933));
  AOI21_X1  g732(.A(new_n876), .B1(new_n932), .B2(new_n933), .ZN(new_n934));
  NAND3_X1  g733(.A1(new_n266), .A2(new_n856), .A3(new_n862), .ZN(new_n935));
  AOI21_X1  g734(.A(new_n669), .B1(new_n935), .B2(new_n872), .ZN(new_n936));
  NAND2_X1  g735(.A1(new_n936), .A2(KEYINPUT115), .ZN(new_n937));
  AOI21_X1  g736(.A(new_n716), .B1(new_n934), .B2(new_n937), .ZN(new_n938));
  AOI21_X1  g737(.A(new_n923), .B1(new_n938), .B2(KEYINPUT116), .ZN(new_n939));
  OAI22_X1  g738(.A1(new_n936), .A2(KEYINPUT115), .B1(new_n748), .B2(new_n875), .ZN(new_n940));
  NOR2_X1   g739(.A1(new_n932), .A2(new_n933), .ZN(new_n941));
  OAI21_X1  g740(.A(new_n637), .B1(new_n940), .B2(new_n941), .ZN(new_n942));
  INV_X1    g741(.A(KEYINPUT116), .ZN(new_n943));
  NAND2_X1  g742(.A1(new_n942), .A2(new_n943), .ZN(new_n944));
  AOI21_X1  g743(.A(new_n922), .B1(new_n939), .B2(new_n944), .ZN(new_n945));
  AOI21_X1  g744(.A(new_n465), .B1(new_n877), .B2(new_n878), .ZN(new_n946));
  NOR2_X1   g745(.A1(new_n946), .A2(KEYINPUT57), .ZN(new_n947));
  OAI211_X1 g746(.A(new_n790), .B(new_n919), .C1(new_n945), .C2(new_n947), .ZN(new_n948));
  NAND2_X1  g747(.A1(new_n948), .A2(G141gat), .ZN(new_n949));
  NOR2_X1   g748(.A1(new_n267), .A2(G141gat), .ZN(new_n950));
  NAND4_X1  g749(.A1(new_n946), .A2(new_n588), .A3(new_n917), .A4(new_n950), .ZN(new_n951));
  AOI21_X1  g750(.A(new_n915), .B1(new_n949), .B2(new_n951), .ZN(new_n952));
  AOI21_X1  g751(.A(KEYINPUT58), .B1(new_n951), .B2(KEYINPUT117), .ZN(new_n953));
  AOI211_X1 g752(.A(new_n465), .B(new_n916), .C1(new_n877), .C2(new_n878), .ZN(new_n954));
  INV_X1    g753(.A(KEYINPUT117), .ZN(new_n955));
  NAND4_X1  g754(.A1(new_n954), .A2(new_n955), .A3(new_n588), .A4(new_n950), .ZN(new_n956));
  NAND2_X1  g755(.A1(new_n953), .A2(new_n956), .ZN(new_n957));
  OAI211_X1 g756(.A(new_n266), .B(new_n919), .C1(new_n945), .C2(new_n947), .ZN(new_n958));
  AOI21_X1  g757(.A(new_n957), .B1(G141gat), .B2(new_n958), .ZN(new_n959));
  OAI21_X1  g758(.A(new_n914), .B1(new_n952), .B2(new_n959), .ZN(new_n960));
  NAND2_X1  g759(.A1(new_n958), .A2(G141gat), .ZN(new_n961));
  NAND3_X1  g760(.A1(new_n961), .A2(new_n956), .A3(new_n953), .ZN(new_n962));
  INV_X1    g761(.A(new_n954), .ZN(new_n963));
  NOR2_X1   g762(.A1(new_n963), .A2(new_n532), .ZN(new_n964));
  AOI22_X1  g763(.A1(new_n948), .A2(G141gat), .B1(new_n964), .B2(new_n950), .ZN(new_n965));
  OAI211_X1 g764(.A(new_n962), .B(KEYINPUT118), .C1(new_n915), .C2(new_n965), .ZN(new_n966));
  NAND2_X1  g765(.A1(new_n960), .A2(new_n966), .ZN(G1344gat));
  INV_X1    g766(.A(G148gat), .ZN(new_n968));
  NAND3_X1  g767(.A1(new_n964), .A2(new_n968), .A3(new_n693), .ZN(new_n969));
  INV_X1    g768(.A(KEYINPUT59), .ZN(new_n970));
  AOI21_X1  g769(.A(new_n922), .B1(new_n877), .B2(new_n878), .ZN(new_n971));
  INV_X1    g770(.A(KEYINPUT119), .ZN(new_n972));
  NAND2_X1  g771(.A1(new_n971), .A2(new_n972), .ZN(new_n973));
  OAI21_X1  g772(.A(new_n932), .B1(new_n719), .B2(new_n875), .ZN(new_n974));
  AOI22_X1  g773(.A1(new_n694), .A2(new_n267), .B1(new_n974), .B2(new_n637), .ZN(new_n975));
  OAI21_X1  g774(.A(new_n920), .B1(new_n975), .B2(new_n465), .ZN(new_n976));
  AND2_X1   g775(.A1(new_n976), .A2(new_n972), .ZN(new_n977));
  OAI21_X1  g776(.A(new_n973), .B1(new_n977), .B2(new_n971), .ZN(new_n978));
  NAND3_X1  g777(.A1(new_n978), .A2(new_n693), .A3(new_n919), .ZN(new_n979));
  AOI21_X1  g778(.A(new_n970), .B1(new_n979), .B2(G148gat), .ZN(new_n980));
  NAND2_X1  g779(.A1(new_n939), .A2(new_n944), .ZN(new_n981));
  NAND2_X1  g780(.A1(new_n981), .A2(new_n921), .ZN(new_n982));
  INV_X1    g781(.A(new_n947), .ZN(new_n983));
  AOI21_X1  g782(.A(new_n918), .B1(new_n982), .B2(new_n983), .ZN(new_n984));
  AOI211_X1 g783(.A(KEYINPUT59), .B(new_n968), .C1(new_n984), .C2(new_n693), .ZN(new_n985));
  OAI21_X1  g784(.A(new_n969), .B1(new_n980), .B2(new_n985), .ZN(G1345gat));
  NOR3_X1   g785(.A1(new_n963), .A2(new_n532), .A3(new_n637), .ZN(new_n987));
  INV_X1    g786(.A(KEYINPUT120), .ZN(new_n988));
  OR2_X1    g787(.A1(new_n987), .A2(new_n988), .ZN(new_n989));
  AOI21_X1  g788(.A(G155gat), .B1(new_n987), .B2(new_n988), .ZN(new_n990));
  AND2_X1   g789(.A1(new_n716), .A2(G155gat), .ZN(new_n991));
  AOI22_X1  g790(.A1(new_n989), .A2(new_n990), .B1(new_n984), .B2(new_n991), .ZN(G1346gat));
  INV_X1    g791(.A(G162gat), .ZN(new_n993));
  AOI21_X1  g792(.A(new_n993), .B1(new_n984), .B2(new_n845), .ZN(new_n994));
  AND3_X1   g793(.A1(new_n954), .A2(new_n993), .A3(new_n901), .ZN(new_n995));
  OR3_X1    g794(.A1(new_n994), .A2(KEYINPUT121), .A3(new_n995), .ZN(new_n996));
  OAI21_X1  g795(.A(KEYINPUT121), .B1(new_n994), .B2(new_n995), .ZN(new_n997));
  NAND2_X1  g796(.A1(new_n996), .A2(new_n997), .ZN(G1347gat));
  AOI21_X1  g797(.A(new_n696), .B1(new_n877), .B2(new_n878), .ZN(new_n999));
  XNOR2_X1  g798(.A(new_n999), .B(KEYINPUT122), .ZN(new_n1000));
  NOR2_X1   g799(.A1(new_n466), .A2(new_n588), .ZN(new_n1001));
  NOR2_X1   g800(.A1(new_n759), .A2(G169gat), .ZN(new_n1002));
  NAND3_X1  g801(.A1(new_n1000), .A2(new_n1001), .A3(new_n1002), .ZN(new_n1003));
  NOR2_X1   g802(.A1(new_n1003), .A2(KEYINPUT123), .ZN(new_n1004));
  INV_X1    g803(.A(KEYINPUT123), .ZN(new_n1005));
  NOR2_X1   g804(.A1(new_n696), .A2(new_n588), .ZN(new_n1006));
  XNOR2_X1  g805(.A(new_n1006), .B(KEYINPUT124), .ZN(new_n1007));
  AND2_X1   g806(.A1(new_n1007), .A2(new_n537), .ZN(new_n1008));
  NAND3_X1  g807(.A1(new_n1008), .A2(new_n266), .A3(new_n879), .ZN(new_n1009));
  AOI21_X1  g808(.A(new_n1005), .B1(new_n1009), .B2(G169gat), .ZN(new_n1010));
  AOI21_X1  g809(.A(new_n1004), .B1(new_n1003), .B2(new_n1010), .ZN(G1348gat));
  NAND2_X1  g810(.A1(new_n1008), .A2(new_n879), .ZN(new_n1012));
  INV_X1    g811(.A(G176gat), .ZN(new_n1013));
  NOR3_X1   g812(.A1(new_n1012), .A2(new_n1013), .A3(new_n809), .ZN(new_n1014));
  NAND2_X1  g813(.A1(new_n1000), .A2(new_n1001), .ZN(new_n1015));
  OAI21_X1  g814(.A(new_n1013), .B1(new_n1015), .B2(new_n809), .ZN(new_n1016));
  INV_X1    g815(.A(KEYINPUT125), .ZN(new_n1017));
  OR2_X1    g816(.A1(new_n1016), .A2(new_n1017), .ZN(new_n1018));
  NAND2_X1  g817(.A1(new_n1016), .A2(new_n1017), .ZN(new_n1019));
  AOI21_X1  g818(.A(new_n1014), .B1(new_n1018), .B2(new_n1019), .ZN(G1349gat));
  OAI21_X1  g819(.A(new_n303), .B1(new_n1012), .B2(new_n637), .ZN(new_n1021));
  NAND2_X1  g820(.A1(new_n716), .A2(new_n271), .ZN(new_n1022));
  OAI21_X1  g821(.A(new_n1021), .B1(new_n1015), .B2(new_n1022), .ZN(new_n1023));
  XNOR2_X1  g822(.A(new_n1023), .B(KEYINPUT60), .ZN(G1350gat));
  OAI21_X1  g823(.A(G190gat), .B1(new_n1012), .B2(new_n719), .ZN(new_n1025));
  XNOR2_X1  g824(.A(new_n1025), .B(KEYINPUT61), .ZN(new_n1026));
  NAND2_X1  g825(.A1(new_n845), .A2(new_n272), .ZN(new_n1027));
  OAI21_X1  g826(.A(new_n1026), .B1(new_n1015), .B2(new_n1027), .ZN(G1351gat));
  AND4_X1   g827(.A1(new_n532), .A2(new_n1000), .A3(new_n536), .A4(new_n546), .ZN(new_n1029));
  XOR2_X1   g828(.A(KEYINPUT126), .B(G197gat), .Z(new_n1030));
  NAND3_X1  g829(.A1(new_n1029), .A2(new_n790), .A3(new_n1030), .ZN(new_n1031));
  NAND2_X1  g830(.A1(new_n1007), .A2(new_n546), .ZN(new_n1032));
  XNOR2_X1  g831(.A(new_n1032), .B(KEYINPUT127), .ZN(new_n1033));
  NAND2_X1  g832(.A1(new_n978), .A2(new_n1033), .ZN(new_n1034));
  NOR2_X1   g833(.A1(new_n1034), .A2(new_n267), .ZN(new_n1035));
  OAI21_X1  g834(.A(new_n1031), .B1(new_n1035), .B2(new_n1030), .ZN(G1352gat));
  NOR2_X1   g835(.A1(new_n809), .A2(G204gat), .ZN(new_n1037));
  NAND2_X1  g836(.A1(new_n1029), .A2(new_n1037), .ZN(new_n1038));
  NAND2_X1  g837(.A1(new_n1038), .A2(KEYINPUT62), .ZN(new_n1039));
  NAND3_X1  g838(.A1(new_n978), .A2(new_n693), .A3(new_n1033), .ZN(new_n1040));
  NAND2_X1  g839(.A1(new_n1040), .A2(G204gat), .ZN(new_n1041));
  INV_X1    g840(.A(KEYINPUT62), .ZN(new_n1042));
  NAND3_X1  g841(.A1(new_n1029), .A2(new_n1042), .A3(new_n1037), .ZN(new_n1043));
  NAND3_X1  g842(.A1(new_n1039), .A2(new_n1041), .A3(new_n1043), .ZN(G1353gat));
  NAND3_X1  g843(.A1(new_n1029), .A2(new_n402), .A3(new_n716), .ZN(new_n1045));
  NAND3_X1  g844(.A1(new_n978), .A2(new_n716), .A3(new_n1033), .ZN(new_n1046));
  AND3_X1   g845(.A1(new_n1046), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n1047));
  AOI21_X1  g846(.A(KEYINPUT63), .B1(new_n1046), .B2(G211gat), .ZN(new_n1048));
  OAI21_X1  g847(.A(new_n1045), .B1(new_n1047), .B2(new_n1048), .ZN(G1354gat));
  OAI21_X1  g848(.A(G218gat), .B1(new_n1034), .B2(new_n719), .ZN(new_n1050));
  NAND3_X1  g849(.A1(new_n1029), .A2(new_n403), .A3(new_n845), .ZN(new_n1051));
  NAND2_X1  g850(.A1(new_n1050), .A2(new_n1051), .ZN(G1355gat));
endmodule


