

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301,
         n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312,
         n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323,
         n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334,
         n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
         n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
         n588, n589, n590, n591, n592;

  XNOR2_X1 U323 ( .A(n404), .B(n403), .ZN(n405) );
  XNOR2_X1 U324 ( .A(n347), .B(G50GAT), .ZN(n348) );
  INV_X1 U325 ( .A(KEYINPUT48), .ZN(n473) );
  XNOR2_X1 U326 ( .A(n349), .B(n348), .ZN(n350) );
  XNOR2_X1 U327 ( .A(n473), .B(KEYINPUT64), .ZN(n474) );
  INV_X1 U328 ( .A(KEYINPUT99), .ZN(n387) );
  XNOR2_X1 U329 ( .A(KEYINPUT98), .B(KEYINPUT36), .ZN(n408) );
  XNOR2_X1 U330 ( .A(n475), .B(n474), .ZN(n534) );
  XNOR2_X1 U331 ( .A(n548), .B(n408), .ZN(n465) );
  XOR2_X1 U332 ( .A(n355), .B(n354), .Z(n479) );
  XNOR2_X1 U333 ( .A(n406), .B(n405), .ZN(n407) );
  NOR2_X1 U334 ( .A1(n536), .A2(n481), .ZN(n573) );
  INV_X1 U335 ( .A(G50GAT), .ZN(n457) );
  INV_X1 U336 ( .A(G43GAT), .ZN(n454) );
  XNOR2_X1 U337 ( .A(n482), .B(G190GAT), .ZN(n483) );
  XNOR2_X1 U338 ( .A(n457), .B(KEYINPUT104), .ZN(n458) );
  XNOR2_X1 U339 ( .A(n454), .B(KEYINPUT40), .ZN(n455) );
  XNOR2_X1 U340 ( .A(n484), .B(n483), .ZN(G1351GAT) );
  XNOR2_X1 U341 ( .A(n459), .B(n458), .ZN(G1331GAT) );
  XOR2_X1 U342 ( .A(KEYINPUT84), .B(KEYINPUT20), .Z(n292) );
  XNOR2_X1 U343 ( .A(G43GAT), .B(G99GAT), .ZN(n291) );
  XNOR2_X1 U344 ( .A(n292), .B(n291), .ZN(n306) );
  XOR2_X1 U345 ( .A(KEYINPUT0), .B(G127GAT), .Z(n310) );
  XOR2_X1 U346 ( .A(G120GAT), .B(G71GAT), .Z(n434) );
  XOR2_X1 U347 ( .A(n310), .B(n434), .Z(n294) );
  XOR2_X1 U348 ( .A(G113GAT), .B(G15GAT), .Z(n424) );
  XOR2_X1 U349 ( .A(G190GAT), .B(G134GAT), .Z(n402) );
  XNOR2_X1 U350 ( .A(n424), .B(n402), .ZN(n293) );
  XNOR2_X1 U351 ( .A(n294), .B(n293), .ZN(n298) );
  XOR2_X1 U352 ( .A(KEYINPUT83), .B(KEYINPUT85), .Z(n296) );
  NAND2_X1 U353 ( .A1(G227GAT), .A2(G233GAT), .ZN(n295) );
  XNOR2_X1 U354 ( .A(n296), .B(n295), .ZN(n297) );
  XOR2_X1 U355 ( .A(n298), .B(n297), .Z(n304) );
  XNOR2_X1 U356 ( .A(G183GAT), .B(KEYINPUT18), .ZN(n299) );
  XNOR2_X1 U357 ( .A(n299), .B(KEYINPUT17), .ZN(n300) );
  XOR2_X1 U358 ( .A(n300), .B(KEYINPUT19), .Z(n302) );
  XNOR2_X1 U359 ( .A(G169GAT), .B(G176GAT), .ZN(n301) );
  XNOR2_X1 U360 ( .A(n302), .B(n301), .ZN(n330) );
  XNOR2_X1 U361 ( .A(n330), .B(KEYINPUT86), .ZN(n303) );
  XNOR2_X1 U362 ( .A(n304), .B(n303), .ZN(n305) );
  XNOR2_X1 U363 ( .A(n306), .B(n305), .ZN(n526) );
  INV_X1 U364 ( .A(n526), .ZN(n536) );
  XOR2_X1 U365 ( .A(KEYINPUT100), .B(KEYINPUT37), .Z(n411) );
  XOR2_X1 U366 ( .A(n526), .B(KEYINPUT87), .Z(n358) );
  XOR2_X1 U367 ( .A(G85GAT), .B(G120GAT), .Z(n308) );
  XNOR2_X1 U368 ( .A(G113GAT), .B(G134GAT), .ZN(n307) );
  XNOR2_X1 U369 ( .A(n308), .B(n307), .ZN(n309) );
  XOR2_X1 U370 ( .A(n309), .B(G162GAT), .Z(n312) );
  XNOR2_X1 U371 ( .A(G29GAT), .B(n310), .ZN(n311) );
  XNOR2_X1 U372 ( .A(n312), .B(n311), .ZN(n318) );
  XOR2_X1 U373 ( .A(KEYINPUT3), .B(KEYINPUT90), .Z(n314) );
  XNOR2_X1 U374 ( .A(G155GAT), .B(KEYINPUT2), .ZN(n313) );
  XNOR2_X1 U375 ( .A(n314), .B(n313), .ZN(n346) );
  XOR2_X1 U376 ( .A(n346), .B(KEYINPUT4), .Z(n316) );
  NAND2_X1 U377 ( .A1(G225GAT), .A2(G233GAT), .ZN(n315) );
  XNOR2_X1 U378 ( .A(n316), .B(n315), .ZN(n317) );
  XOR2_X1 U379 ( .A(n318), .B(n317), .Z(n326) );
  XOR2_X1 U380 ( .A(KEYINPUT6), .B(KEYINPUT93), .Z(n320) );
  XNOR2_X1 U381 ( .A(G141GAT), .B(G148GAT), .ZN(n319) );
  XNOR2_X1 U382 ( .A(n320), .B(n319), .ZN(n324) );
  XOR2_X1 U383 ( .A(G57GAT), .B(KEYINPUT1), .Z(n322) );
  XNOR2_X1 U384 ( .A(G1GAT), .B(KEYINPUT5), .ZN(n321) );
  XNOR2_X1 U385 ( .A(n322), .B(n321), .ZN(n323) );
  XNOR2_X1 U386 ( .A(n324), .B(n323), .ZN(n325) );
  XOR2_X1 U387 ( .A(n326), .B(n325), .Z(n522) );
  INV_X1 U388 ( .A(n522), .ZN(n500) );
  XOR2_X1 U389 ( .A(KEYINPUT21), .B(G211GAT), .Z(n328) );
  XNOR2_X1 U390 ( .A(KEYINPUT89), .B(G204GAT), .ZN(n327) );
  XNOR2_X1 U391 ( .A(n328), .B(n327), .ZN(n329) );
  XOR2_X1 U392 ( .A(G197GAT), .B(n329), .Z(n355) );
  XNOR2_X1 U393 ( .A(n330), .B(n355), .ZN(n340) );
  XOR2_X1 U394 ( .A(G92GAT), .B(G190GAT), .Z(n332) );
  XNOR2_X1 U395 ( .A(G36GAT), .B(G8GAT), .ZN(n331) );
  XNOR2_X1 U396 ( .A(n332), .B(n331), .ZN(n336) );
  XOR2_X1 U397 ( .A(KEYINPUT94), .B(KEYINPUT76), .Z(n334) );
  XOR2_X1 U398 ( .A(KEYINPUT72), .B(G64GAT), .Z(n436) );
  XNOR2_X1 U399 ( .A(G218GAT), .B(n436), .ZN(n333) );
  XNOR2_X1 U400 ( .A(n334), .B(n333), .ZN(n335) );
  XOR2_X1 U401 ( .A(n336), .B(n335), .Z(n338) );
  NAND2_X1 U402 ( .A1(G226GAT), .A2(G233GAT), .ZN(n337) );
  XNOR2_X1 U403 ( .A(n338), .B(n337), .ZN(n339) );
  XOR2_X1 U404 ( .A(n340), .B(n339), .Z(n505) );
  XNOR2_X1 U405 ( .A(n505), .B(KEYINPUT27), .ZN(n362) );
  NOR2_X1 U406 ( .A1(n500), .A2(n362), .ZN(n535) );
  XOR2_X1 U407 ( .A(KEYINPUT23), .B(KEYINPUT88), .Z(n342) );
  XNOR2_X1 U408 ( .A(KEYINPUT24), .B(KEYINPUT91), .ZN(n341) );
  XNOR2_X1 U409 ( .A(n342), .B(n341), .ZN(n353) );
  XOR2_X1 U410 ( .A(KEYINPUT92), .B(KEYINPUT22), .Z(n344) );
  XOR2_X1 U411 ( .A(G141GAT), .B(G22GAT), .Z(n423) );
  XOR2_X1 U412 ( .A(G148GAT), .B(G78GAT), .Z(n435) );
  XNOR2_X1 U413 ( .A(n423), .B(n435), .ZN(n343) );
  XNOR2_X1 U414 ( .A(n344), .B(n343), .ZN(n345) );
  XOR2_X1 U415 ( .A(n345), .B(G106GAT), .Z(n351) );
  XOR2_X1 U416 ( .A(G218GAT), .B(G162GAT), .Z(n401) );
  XOR2_X1 U417 ( .A(n401), .B(n346), .Z(n349) );
  NAND2_X1 U418 ( .A1(G228GAT), .A2(G233GAT), .ZN(n347) );
  XNOR2_X1 U419 ( .A(n351), .B(n350), .ZN(n352) );
  XOR2_X1 U420 ( .A(n353), .B(n352), .Z(n354) );
  XNOR2_X1 U421 ( .A(n479), .B(KEYINPUT28), .ZN(n539) );
  INV_X1 U422 ( .A(n539), .ZN(n497) );
  NAND2_X1 U423 ( .A1(n535), .A2(n497), .ZN(n356) );
  XOR2_X1 U424 ( .A(KEYINPUT95), .B(n356), .Z(n357) );
  NOR2_X1 U425 ( .A1(n358), .A2(n357), .ZN(n367) );
  NOR2_X1 U426 ( .A1(n536), .A2(n505), .ZN(n359) );
  NOR2_X1 U427 ( .A1(n479), .A2(n359), .ZN(n360) );
  XOR2_X1 U428 ( .A(KEYINPUT25), .B(n360), .Z(n364) );
  NAND2_X1 U429 ( .A1(n479), .A2(n536), .ZN(n361) );
  XNOR2_X1 U430 ( .A(n361), .B(KEYINPUT26), .ZN(n576) );
  NOR2_X1 U431 ( .A1(n362), .A2(n576), .ZN(n363) );
  NOR2_X1 U432 ( .A1(n364), .A2(n363), .ZN(n365) );
  NOR2_X1 U433 ( .A1(n522), .A2(n365), .ZN(n366) );
  NOR2_X1 U434 ( .A1(n367), .A2(n366), .ZN(n488) );
  XOR2_X1 U435 ( .A(KEYINPUT79), .B(KEYINPUT80), .Z(n369) );
  XNOR2_X1 U436 ( .A(G64GAT), .B(KEYINPUT81), .ZN(n368) );
  XNOR2_X1 U437 ( .A(n369), .B(n368), .ZN(n381) );
  XOR2_X1 U438 ( .A(G127GAT), .B(G71GAT), .Z(n371) );
  XNOR2_X1 U439 ( .A(G15GAT), .B(G183GAT), .ZN(n370) );
  XNOR2_X1 U440 ( .A(n371), .B(n370), .ZN(n379) );
  XOR2_X1 U441 ( .A(KEYINPUT82), .B(KEYINPUT14), .Z(n373) );
  XNOR2_X1 U442 ( .A(KEYINPUT12), .B(KEYINPUT15), .ZN(n372) );
  XNOR2_X1 U443 ( .A(n373), .B(n372), .ZN(n377) );
  XOR2_X1 U444 ( .A(G78GAT), .B(G155GAT), .Z(n375) );
  XNOR2_X1 U445 ( .A(G22GAT), .B(G211GAT), .ZN(n374) );
  XNOR2_X1 U446 ( .A(n375), .B(n374), .ZN(n376) );
  XOR2_X1 U447 ( .A(n377), .B(n376), .Z(n378) );
  XNOR2_X1 U448 ( .A(n379), .B(n378), .ZN(n380) );
  XNOR2_X1 U449 ( .A(n381), .B(n380), .ZN(n386) );
  XOR2_X1 U450 ( .A(G57GAT), .B(KEYINPUT13), .Z(n441) );
  XNOR2_X1 U451 ( .A(G1GAT), .B(KEYINPUT68), .ZN(n382) );
  XNOR2_X1 U452 ( .A(n382), .B(G8GAT), .ZN(n421) );
  XOR2_X1 U453 ( .A(n441), .B(n421), .Z(n384) );
  NAND2_X1 U454 ( .A1(G231GAT), .A2(G233GAT), .ZN(n383) );
  XNOR2_X1 U455 ( .A(n384), .B(n383), .ZN(n385) );
  XOR2_X1 U456 ( .A(n386), .B(n385), .Z(n485) );
  INV_X1 U457 ( .A(n485), .ZN(n587) );
  NOR2_X1 U458 ( .A1(n488), .A2(n587), .ZN(n388) );
  XNOR2_X1 U459 ( .A(n388), .B(n387), .ZN(n409) );
  XOR2_X1 U460 ( .A(G43GAT), .B(G29GAT), .Z(n390) );
  XNOR2_X1 U461 ( .A(G50GAT), .B(KEYINPUT7), .ZN(n389) );
  XNOR2_X1 U462 ( .A(n390), .B(n389), .ZN(n391) );
  XOR2_X1 U463 ( .A(n391), .B(KEYINPUT67), .Z(n393) );
  XNOR2_X1 U464 ( .A(G36GAT), .B(KEYINPUT8), .ZN(n392) );
  XNOR2_X1 U465 ( .A(n393), .B(n392), .ZN(n418) );
  INV_X1 U466 ( .A(KEYINPUT10), .ZN(n396) );
  XOR2_X1 U467 ( .A(G92GAT), .B(G85GAT), .Z(n395) );
  XNOR2_X1 U468 ( .A(G99GAT), .B(G106GAT), .ZN(n394) );
  XNOR2_X1 U469 ( .A(n395), .B(n394), .ZN(n447) );
  XNOR2_X1 U470 ( .A(n396), .B(n447), .ZN(n398) );
  NAND2_X1 U471 ( .A1(G232GAT), .A2(G233GAT), .ZN(n397) );
  XNOR2_X1 U472 ( .A(n398), .B(n397), .ZN(n406) );
  XOR2_X1 U473 ( .A(KEYINPUT76), .B(KEYINPUT11), .Z(n400) );
  XNOR2_X1 U474 ( .A(KEYINPUT77), .B(KEYINPUT9), .ZN(n399) );
  XOR2_X1 U475 ( .A(n400), .B(n399), .Z(n404) );
  XNOR2_X1 U476 ( .A(n402), .B(n401), .ZN(n403) );
  XNOR2_X1 U477 ( .A(n418), .B(n407), .ZN(n562) );
  INV_X1 U478 ( .A(n562), .ZN(n463) );
  XOR2_X1 U479 ( .A(KEYINPUT78), .B(n463), .Z(n548) );
  NAND2_X1 U480 ( .A1(n409), .A2(n465), .ZN(n410) );
  XNOR2_X1 U481 ( .A(n411), .B(n410), .ZN(n521) );
  XOR2_X1 U482 ( .A(KEYINPUT30), .B(KEYINPUT65), .Z(n413) );
  NAND2_X1 U483 ( .A1(G229GAT), .A2(G233GAT), .ZN(n412) );
  XNOR2_X1 U484 ( .A(n413), .B(n412), .ZN(n414) );
  XOR2_X1 U485 ( .A(n414), .B(KEYINPUT29), .Z(n420) );
  XOR2_X1 U486 ( .A(KEYINPUT66), .B(KEYINPUT69), .Z(n416) );
  XNOR2_X1 U487 ( .A(G169GAT), .B(G197GAT), .ZN(n415) );
  XNOR2_X1 U488 ( .A(n416), .B(n415), .ZN(n417) );
  XNOR2_X1 U489 ( .A(n418), .B(n417), .ZN(n419) );
  XNOR2_X1 U490 ( .A(n420), .B(n419), .ZN(n422) );
  XOR2_X1 U491 ( .A(n422), .B(n421), .Z(n426) );
  XNOR2_X1 U492 ( .A(n424), .B(n423), .ZN(n425) );
  XNOR2_X1 U493 ( .A(n426), .B(n425), .ZN(n578) );
  XNOR2_X1 U494 ( .A(n578), .B(KEYINPUT70), .ZN(n565) );
  INV_X1 U495 ( .A(KEYINPUT74), .ZN(n427) );
  NAND2_X1 U496 ( .A1(KEYINPUT31), .A2(n427), .ZN(n430) );
  INV_X1 U497 ( .A(KEYINPUT31), .ZN(n428) );
  NAND2_X1 U498 ( .A1(n428), .A2(KEYINPUT74), .ZN(n429) );
  NAND2_X1 U499 ( .A1(n430), .A2(n429), .ZN(n432) );
  XNOR2_X1 U500 ( .A(KEYINPUT32), .B(KEYINPUT73), .ZN(n431) );
  XNOR2_X1 U501 ( .A(n432), .B(n431), .ZN(n433) );
  XOR2_X1 U502 ( .A(n434), .B(n433), .Z(n440) );
  XNOR2_X1 U503 ( .A(n436), .B(n435), .ZN(n438) );
  AND2_X1 U504 ( .A1(G230GAT), .A2(G233GAT), .ZN(n437) );
  XNOR2_X1 U505 ( .A(n438), .B(n437), .ZN(n439) );
  XNOR2_X1 U506 ( .A(n440), .B(n439), .ZN(n442) );
  XNOR2_X1 U507 ( .A(n442), .B(n441), .ZN(n444) );
  XNOR2_X1 U508 ( .A(G176GAT), .B(G204GAT), .ZN(n443) );
  XNOR2_X1 U509 ( .A(n444), .B(n443), .ZN(n446) );
  INV_X1 U510 ( .A(KEYINPUT71), .ZN(n445) );
  XNOR2_X1 U511 ( .A(n446), .B(n445), .ZN(n449) );
  XNOR2_X1 U512 ( .A(n447), .B(KEYINPUT33), .ZN(n448) );
  XOR2_X1 U513 ( .A(n449), .B(n448), .Z(n583) );
  INV_X1 U514 ( .A(n583), .ZN(n468) );
  NAND2_X1 U515 ( .A1(n565), .A2(n468), .ZN(n450) );
  XOR2_X1 U516 ( .A(KEYINPUT75), .B(n450), .Z(n490) );
  NOR2_X1 U517 ( .A1(n521), .A2(n490), .ZN(n452) );
  XNOR2_X1 U518 ( .A(KEYINPUT102), .B(KEYINPUT38), .ZN(n451) );
  XNOR2_X1 U519 ( .A(n452), .B(n451), .ZN(n453) );
  XNOR2_X1 U520 ( .A(KEYINPUT101), .B(n453), .ZN(n504) );
  NOR2_X1 U521 ( .A1(n536), .A2(n504), .ZN(n456) );
  XNOR2_X1 U522 ( .A(n456), .B(n455), .ZN(G1330GAT) );
  NOR2_X1 U523 ( .A1(n497), .A2(n504), .ZN(n459) );
  INV_X1 U524 ( .A(n505), .ZN(n524) );
  XOR2_X1 U525 ( .A(n583), .B(KEYINPUT41), .Z(n507) );
  AND2_X1 U526 ( .A1(n578), .A2(n507), .ZN(n460) );
  XNOR2_X1 U527 ( .A(n460), .B(KEYINPUT46), .ZN(n461) );
  NOR2_X1 U528 ( .A1(n587), .A2(n461), .ZN(n462) );
  NAND2_X1 U529 ( .A1(n463), .A2(n462), .ZN(n464) );
  XNOR2_X1 U530 ( .A(n464), .B(KEYINPUT47), .ZN(n472) );
  NAND2_X1 U531 ( .A1(n465), .A2(n587), .ZN(n467) );
  XOR2_X1 U532 ( .A(KEYINPUT45), .B(KEYINPUT112), .Z(n466) );
  XNOR2_X1 U533 ( .A(n467), .B(n466), .ZN(n469) );
  NAND2_X1 U534 ( .A1(n469), .A2(n468), .ZN(n470) );
  NOR2_X1 U535 ( .A1(n565), .A2(n470), .ZN(n471) );
  NOR2_X1 U536 ( .A1(n472), .A2(n471), .ZN(n475) );
  NAND2_X1 U537 ( .A1(n524), .A2(n534), .ZN(n477) );
  XOR2_X1 U538 ( .A(KEYINPUT54), .B(KEYINPUT120), .Z(n476) );
  XNOR2_X1 U539 ( .A(n477), .B(n476), .ZN(n478) );
  NAND2_X1 U540 ( .A1(n500), .A2(n478), .ZN(n575) );
  NOR2_X1 U541 ( .A1(n575), .A2(n479), .ZN(n480) );
  XNOR2_X1 U542 ( .A(n480), .B(KEYINPUT55), .ZN(n481) );
  NAND2_X1 U543 ( .A1(n573), .A2(n548), .ZN(n484) );
  XOR2_X1 U544 ( .A(KEYINPUT123), .B(KEYINPUT58), .Z(n482) );
  XOR2_X1 U545 ( .A(KEYINPUT97), .B(KEYINPUT34), .Z(n492) );
  NOR2_X1 U546 ( .A1(n548), .A2(n485), .ZN(n486) );
  XOR2_X1 U547 ( .A(KEYINPUT16), .B(n486), .Z(n487) );
  NOR2_X1 U548 ( .A1(n488), .A2(n487), .ZN(n489) );
  XOR2_X1 U549 ( .A(KEYINPUT96), .B(n489), .Z(n509) );
  NOR2_X1 U550 ( .A1(n509), .A2(n490), .ZN(n498) );
  NAND2_X1 U551 ( .A1(n498), .A2(n522), .ZN(n491) );
  XNOR2_X1 U552 ( .A(n492), .B(n491), .ZN(n493) );
  XNOR2_X1 U553 ( .A(G1GAT), .B(n493), .ZN(G1324GAT) );
  NAND2_X1 U554 ( .A1(n498), .A2(n524), .ZN(n494) );
  XNOR2_X1 U555 ( .A(n494), .B(G8GAT), .ZN(G1325GAT) );
  XOR2_X1 U556 ( .A(G15GAT), .B(KEYINPUT35), .Z(n496) );
  NAND2_X1 U557 ( .A1(n498), .A2(n526), .ZN(n495) );
  XNOR2_X1 U558 ( .A(n496), .B(n495), .ZN(G1326GAT) );
  NAND2_X1 U559 ( .A1(n539), .A2(n498), .ZN(n499) );
  XNOR2_X1 U560 ( .A(n499), .B(G22GAT), .ZN(G1327GAT) );
  NOR2_X1 U561 ( .A1(n500), .A2(n504), .ZN(n502) );
  XNOR2_X1 U562 ( .A(KEYINPUT39), .B(KEYINPUT103), .ZN(n501) );
  XNOR2_X1 U563 ( .A(n502), .B(n501), .ZN(n503) );
  XOR2_X1 U564 ( .A(G29GAT), .B(n503), .Z(G1328GAT) );
  NOR2_X1 U565 ( .A1(n505), .A2(n504), .ZN(n506) );
  XOR2_X1 U566 ( .A(G36GAT), .B(n506), .Z(G1329GAT) );
  XOR2_X1 U567 ( .A(KEYINPUT42), .B(KEYINPUT106), .Z(n511) );
  INV_X1 U568 ( .A(n507), .ZN(n541) );
  NOR2_X1 U569 ( .A1(n541), .A2(n578), .ZN(n508) );
  XNOR2_X1 U570 ( .A(n508), .B(KEYINPUT105), .ZN(n520) );
  NOR2_X1 U571 ( .A1(n509), .A2(n520), .ZN(n517) );
  NAND2_X1 U572 ( .A1(n517), .A2(n522), .ZN(n510) );
  XNOR2_X1 U573 ( .A(n511), .B(n510), .ZN(n512) );
  XOR2_X1 U574 ( .A(G57GAT), .B(n512), .Z(G1332GAT) );
  XOR2_X1 U575 ( .A(G64GAT), .B(KEYINPUT107), .Z(n514) );
  NAND2_X1 U576 ( .A1(n517), .A2(n524), .ZN(n513) );
  XNOR2_X1 U577 ( .A(n514), .B(n513), .ZN(G1333GAT) );
  NAND2_X1 U578 ( .A1(n526), .A2(n517), .ZN(n515) );
  XNOR2_X1 U579 ( .A(n515), .B(KEYINPUT108), .ZN(n516) );
  XNOR2_X1 U580 ( .A(G71GAT), .B(n516), .ZN(G1334GAT) );
  XOR2_X1 U581 ( .A(G78GAT), .B(KEYINPUT43), .Z(n519) );
  NAND2_X1 U582 ( .A1(n517), .A2(n539), .ZN(n518) );
  XNOR2_X1 U583 ( .A(n519), .B(n518), .ZN(G1335GAT) );
  NOR2_X1 U584 ( .A1(n521), .A2(n520), .ZN(n531) );
  NAND2_X1 U585 ( .A1(n531), .A2(n522), .ZN(n523) );
  XNOR2_X1 U586 ( .A(G85GAT), .B(n523), .ZN(G1336GAT) );
  NAND2_X1 U587 ( .A1(n531), .A2(n524), .ZN(n525) );
  XNOR2_X1 U588 ( .A(n525), .B(G92GAT), .ZN(G1337GAT) );
  NAND2_X1 U589 ( .A1(n531), .A2(n526), .ZN(n527) );
  XNOR2_X1 U590 ( .A(G99GAT), .B(n527), .ZN(G1338GAT) );
  XOR2_X1 U591 ( .A(KEYINPUT111), .B(KEYINPUT44), .Z(n529) );
  XNOR2_X1 U592 ( .A(G106GAT), .B(KEYINPUT110), .ZN(n528) );
  XNOR2_X1 U593 ( .A(n529), .B(n528), .ZN(n530) );
  XOR2_X1 U594 ( .A(KEYINPUT109), .B(n530), .Z(n533) );
  NAND2_X1 U595 ( .A1(n531), .A2(n539), .ZN(n532) );
  XNOR2_X1 U596 ( .A(n533), .B(n532), .ZN(G1339GAT) );
  NAND2_X1 U597 ( .A1(n535), .A2(n534), .ZN(n552) );
  NOR2_X1 U598 ( .A1(n536), .A2(n552), .ZN(n537) );
  XNOR2_X1 U599 ( .A(n537), .B(KEYINPUT113), .ZN(n538) );
  NOR2_X1 U600 ( .A1(n539), .A2(n538), .ZN(n549) );
  NAND2_X1 U601 ( .A1(n549), .A2(n565), .ZN(n540) );
  XNOR2_X1 U602 ( .A(G113GAT), .B(n540), .ZN(G1340GAT) );
  XOR2_X1 U603 ( .A(KEYINPUT114), .B(KEYINPUT49), .Z(n543) );
  INV_X1 U604 ( .A(n541), .ZN(n568) );
  NAND2_X1 U605 ( .A1(n549), .A2(n568), .ZN(n542) );
  XNOR2_X1 U606 ( .A(n543), .B(n542), .ZN(n544) );
  XNOR2_X1 U607 ( .A(G120GAT), .B(n544), .ZN(G1341GAT) );
  XOR2_X1 U608 ( .A(KEYINPUT50), .B(KEYINPUT115), .Z(n546) );
  NAND2_X1 U609 ( .A1(n549), .A2(n587), .ZN(n545) );
  XNOR2_X1 U610 ( .A(n546), .B(n545), .ZN(n547) );
  XNOR2_X1 U611 ( .A(G127GAT), .B(n547), .ZN(G1342GAT) );
  XOR2_X1 U612 ( .A(G134GAT), .B(KEYINPUT51), .Z(n551) );
  NAND2_X1 U613 ( .A1(n549), .A2(n548), .ZN(n550) );
  XNOR2_X1 U614 ( .A(n551), .B(n550), .ZN(G1343GAT) );
  XOR2_X1 U615 ( .A(G141GAT), .B(KEYINPUT117), .Z(n555) );
  NOR2_X1 U616 ( .A1(n552), .A2(n576), .ZN(n553) );
  XNOR2_X1 U617 ( .A(n553), .B(KEYINPUT116), .ZN(n563) );
  NAND2_X1 U618 ( .A1(n578), .A2(n563), .ZN(n554) );
  XNOR2_X1 U619 ( .A(n555), .B(n554), .ZN(G1344GAT) );
  XOR2_X1 U620 ( .A(KEYINPUT53), .B(KEYINPUT119), .Z(n557) );
  XNOR2_X1 U621 ( .A(G148GAT), .B(KEYINPUT118), .ZN(n556) );
  XNOR2_X1 U622 ( .A(n557), .B(n556), .ZN(n558) );
  XOR2_X1 U623 ( .A(KEYINPUT52), .B(n558), .Z(n560) );
  NAND2_X1 U624 ( .A1(n563), .A2(n568), .ZN(n559) );
  XNOR2_X1 U625 ( .A(n560), .B(n559), .ZN(G1345GAT) );
  NAND2_X1 U626 ( .A1(n563), .A2(n587), .ZN(n561) );
  XNOR2_X1 U627 ( .A(n561), .B(G155GAT), .ZN(G1346GAT) );
  NAND2_X1 U628 ( .A1(n563), .A2(n562), .ZN(n564) );
  XNOR2_X1 U629 ( .A(n564), .B(G162GAT), .ZN(G1347GAT) );
  XOR2_X1 U630 ( .A(G169GAT), .B(KEYINPUT121), .Z(n567) );
  NAND2_X1 U631 ( .A1(n573), .A2(n565), .ZN(n566) );
  XNOR2_X1 U632 ( .A(n567), .B(n566), .ZN(G1348GAT) );
  XNOR2_X1 U633 ( .A(G176GAT), .B(KEYINPUT57), .ZN(n572) );
  NAND2_X1 U634 ( .A1(n573), .A2(n568), .ZN(n570) );
  XOR2_X1 U635 ( .A(KEYINPUT56), .B(KEYINPUT122), .Z(n569) );
  XNOR2_X1 U636 ( .A(n570), .B(n569), .ZN(n571) );
  XNOR2_X1 U637 ( .A(n572), .B(n571), .ZN(G1349GAT) );
  NAND2_X1 U638 ( .A1(n587), .A2(n573), .ZN(n574) );
  XNOR2_X1 U639 ( .A(n574), .B(G183GAT), .ZN(G1350GAT) );
  NOR2_X1 U640 ( .A1(n576), .A2(n575), .ZN(n577) );
  XNOR2_X1 U641 ( .A(n577), .B(KEYINPUT124), .ZN(n589) );
  NAND2_X1 U642 ( .A1(n578), .A2(n589), .ZN(n580) );
  XOR2_X1 U643 ( .A(G197GAT), .B(KEYINPUT125), .Z(n579) );
  XNOR2_X1 U644 ( .A(n580), .B(n579), .ZN(n582) );
  XOR2_X1 U645 ( .A(KEYINPUT59), .B(KEYINPUT60), .Z(n581) );
  XNOR2_X1 U646 ( .A(n582), .B(n581), .ZN(G1352GAT) );
  XOR2_X1 U647 ( .A(KEYINPUT61), .B(KEYINPUT126), .Z(n585) );
  NAND2_X1 U648 ( .A1(n589), .A2(n583), .ZN(n584) );
  XNOR2_X1 U649 ( .A(n585), .B(n584), .ZN(n586) );
  XNOR2_X1 U650 ( .A(G204GAT), .B(n586), .ZN(G1353GAT) );
  NAND2_X1 U651 ( .A1(n589), .A2(n587), .ZN(n588) );
  XNOR2_X1 U652 ( .A(n588), .B(G211GAT), .ZN(G1354GAT) );
  XOR2_X1 U653 ( .A(KEYINPUT62), .B(KEYINPUT127), .Z(n591) );
  NAND2_X1 U654 ( .A1(n465), .A2(n589), .ZN(n590) );
  XNOR2_X1 U655 ( .A(n591), .B(n590), .ZN(n592) );
  XNOR2_X1 U656 ( .A(n592), .B(G218GAT), .ZN(G1355GAT) );
endmodule

