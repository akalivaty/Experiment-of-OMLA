//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 0 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 0 0 1 1 1 0 0 0 1 1 1 1 1 0 0 1 0 0 1 0 1 0 1 0 0 1 1 1 0 1 0 1 0 0 0 1 0 0 0 0 1 0 0 0 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:23:32 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n679, new_n680, new_n681, new_n682, new_n683, new_n684, new_n685,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n692, new_n693,
    new_n694, new_n695, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n720, new_n721, new_n722, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n744, new_n745, new_n747, new_n748, new_n749,
    new_n750, new_n751, new_n752, new_n753, new_n755, new_n756, new_n757,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n772, new_n773,
    new_n774, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n796,
    new_n797, new_n798, new_n799, new_n800, new_n801, new_n802, new_n803,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n910,
    new_n911, new_n912, new_n913, new_n914, new_n915, new_n916, new_n917,
    new_n918, new_n919, new_n920, new_n921, new_n922, new_n923, new_n924,
    new_n925, new_n926, new_n927, new_n928, new_n929, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n951, new_n952, new_n953, new_n954,
    new_n956, new_n957, new_n958, new_n959, new_n960, new_n961, new_n962,
    new_n963, new_n964, new_n965, new_n966, new_n968, new_n969, new_n970,
    new_n971, new_n972, new_n973, new_n974, new_n975, new_n977, new_n978,
    new_n979, new_n980, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015;
  INV_X1    g000(.A(KEYINPUT68), .ZN(new_n187));
  INV_X1    g001(.A(KEYINPUT65), .ZN(new_n188));
  AND2_X1   g002(.A1(KEYINPUT0), .A2(G128), .ZN(new_n189));
  NOR2_X1   g003(.A1(KEYINPUT0), .A2(G128), .ZN(new_n190));
  NOR2_X1   g004(.A1(new_n189), .A2(new_n190), .ZN(new_n191));
  INV_X1    g005(.A(KEYINPUT64), .ZN(new_n192));
  INV_X1    g006(.A(G146), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n192), .A2(new_n193), .ZN(new_n194));
  NAND2_X1  g008(.A1(KEYINPUT64), .A2(G146), .ZN(new_n195));
  AOI21_X1  g009(.A(G143), .B1(new_n194), .B2(new_n195), .ZN(new_n196));
  INV_X1    g010(.A(G143), .ZN(new_n197));
  NOR2_X1   g011(.A1(new_n197), .A2(G146), .ZN(new_n198));
  OAI211_X1 g012(.A(new_n188), .B(new_n191), .C1(new_n196), .C2(new_n198), .ZN(new_n199));
  NAND3_X1  g013(.A1(new_n194), .A2(G143), .A3(new_n195), .ZN(new_n200));
  NOR2_X1   g014(.A1(new_n193), .A2(G143), .ZN(new_n201));
  INV_X1    g015(.A(new_n201), .ZN(new_n202));
  NAND3_X1  g016(.A1(new_n200), .A2(new_n189), .A3(new_n202), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n199), .A2(new_n203), .ZN(new_n204));
  AND2_X1   g018(.A1(KEYINPUT64), .A2(G146), .ZN(new_n205));
  NOR2_X1   g019(.A1(KEYINPUT64), .A2(G146), .ZN(new_n206));
  OAI21_X1  g020(.A(new_n197), .B1(new_n205), .B2(new_n206), .ZN(new_n207));
  INV_X1    g021(.A(new_n198), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  AOI21_X1  g023(.A(new_n188), .B1(new_n209), .B2(new_n191), .ZN(new_n210));
  OAI21_X1  g024(.A(new_n187), .B1(new_n204), .B2(new_n210), .ZN(new_n211));
  INV_X1    g025(.A(KEYINPUT11), .ZN(new_n212));
  INV_X1    g026(.A(G134), .ZN(new_n213));
  OAI21_X1  g027(.A(new_n212), .B1(new_n213), .B2(G137), .ZN(new_n214));
  INV_X1    g028(.A(G137), .ZN(new_n215));
  NAND3_X1  g029(.A1(new_n215), .A2(KEYINPUT11), .A3(G134), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n213), .A2(G137), .ZN(new_n217));
  NAND3_X1  g031(.A1(new_n214), .A2(new_n216), .A3(new_n217), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n218), .A2(G131), .ZN(new_n219));
  INV_X1    g033(.A(G131), .ZN(new_n220));
  NAND4_X1  g034(.A1(new_n214), .A2(new_n216), .A3(new_n220), .A4(new_n217), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n219), .A2(new_n221), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n194), .A2(new_n195), .ZN(new_n223));
  AOI21_X1  g037(.A(new_n198), .B1(new_n223), .B2(new_n197), .ZN(new_n224));
  XNOR2_X1  g038(.A(KEYINPUT0), .B(G128), .ZN(new_n225));
  OAI21_X1  g039(.A(KEYINPUT65), .B1(new_n224), .B2(new_n225), .ZN(new_n226));
  NAND4_X1  g040(.A1(new_n226), .A2(KEYINPUT68), .A3(new_n199), .A4(new_n203), .ZN(new_n227));
  NAND3_X1  g041(.A1(new_n211), .A2(new_n222), .A3(new_n227), .ZN(new_n228));
  OR2_X1    g042(.A1(KEYINPUT67), .A2(G119), .ZN(new_n229));
  NAND2_X1  g043(.A1(KEYINPUT67), .A2(G119), .ZN(new_n230));
  NAND3_X1  g044(.A1(new_n229), .A2(G116), .A3(new_n230), .ZN(new_n231));
  INV_X1    g045(.A(G119), .ZN(new_n232));
  OAI21_X1  g046(.A(new_n231), .B1(G116), .B2(new_n232), .ZN(new_n233));
  XNOR2_X1  g047(.A(KEYINPUT2), .B(G113), .ZN(new_n234));
  OR2_X1    g048(.A1(new_n233), .A2(new_n234), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n233), .A2(new_n234), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n235), .A2(new_n236), .ZN(new_n237));
  INV_X1    g051(.A(new_n237), .ZN(new_n238));
  XNOR2_X1  g052(.A(KEYINPUT66), .B(KEYINPUT1), .ZN(new_n239));
  NAND4_X1  g053(.A1(new_n200), .A2(G128), .A3(new_n239), .A4(new_n202), .ZN(new_n240));
  INV_X1    g054(.A(G128), .ZN(new_n241));
  INV_X1    g055(.A(KEYINPUT1), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n242), .A2(KEYINPUT66), .ZN(new_n243));
  INV_X1    g057(.A(KEYINPUT66), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n244), .A2(KEYINPUT1), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n243), .A2(new_n245), .ZN(new_n246));
  AOI21_X1  g060(.A(new_n241), .B1(new_n200), .B2(new_n246), .ZN(new_n247));
  OAI21_X1  g061(.A(new_n240), .B1(new_n247), .B2(new_n224), .ZN(new_n248));
  INV_X1    g062(.A(new_n217), .ZN(new_n249));
  NOR2_X1   g063(.A1(new_n213), .A2(G137), .ZN(new_n250));
  OAI21_X1  g064(.A(G131), .B1(new_n249), .B2(new_n250), .ZN(new_n251));
  NAND3_X1  g065(.A1(new_n248), .A2(new_n221), .A3(new_n251), .ZN(new_n252));
  NAND3_X1  g066(.A1(new_n228), .A2(new_n238), .A3(new_n252), .ZN(new_n253));
  INV_X1    g067(.A(KEYINPUT74), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n253), .A2(new_n254), .ZN(new_n255));
  NAND4_X1  g069(.A1(new_n228), .A2(KEYINPUT74), .A3(new_n238), .A4(new_n252), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n228), .A2(new_n252), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n257), .A2(new_n237), .ZN(new_n258));
  NAND3_X1  g072(.A1(new_n255), .A2(new_n256), .A3(new_n258), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n259), .A2(KEYINPUT28), .ZN(new_n260));
  INV_X1    g074(.A(KEYINPUT72), .ZN(new_n261));
  INV_X1    g075(.A(KEYINPUT28), .ZN(new_n262));
  AND3_X1   g076(.A1(new_n253), .A2(new_n261), .A3(new_n262), .ZN(new_n263));
  AOI21_X1  g077(.A(new_n261), .B1(new_n253), .B2(new_n262), .ZN(new_n264));
  NOR2_X1   g078(.A1(new_n263), .A2(new_n264), .ZN(new_n265));
  NOR2_X1   g079(.A1(G237), .A2(G953), .ZN(new_n266));
  NAND2_X1  g080(.A1(new_n266), .A2(G210), .ZN(new_n267));
  XOR2_X1   g081(.A(new_n267), .B(KEYINPUT71), .Z(new_n268));
  XNOR2_X1  g082(.A(KEYINPUT26), .B(G101), .ZN(new_n269));
  XNOR2_X1  g083(.A(KEYINPUT70), .B(KEYINPUT27), .ZN(new_n270));
  XNOR2_X1  g084(.A(new_n269), .B(new_n270), .ZN(new_n271));
  XNOR2_X1  g085(.A(new_n268), .B(new_n271), .ZN(new_n272));
  INV_X1    g086(.A(KEYINPUT29), .ZN(new_n273));
  NOR2_X1   g087(.A1(new_n272), .A2(new_n273), .ZN(new_n274));
  NAND3_X1  g088(.A1(new_n260), .A2(new_n265), .A3(new_n274), .ZN(new_n275));
  INV_X1    g089(.A(KEYINPUT75), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n275), .A2(new_n276), .ZN(new_n277));
  NAND4_X1  g091(.A1(new_n260), .A2(new_n265), .A3(KEYINPUT75), .A4(new_n274), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n277), .A2(new_n278), .ZN(new_n279));
  XOR2_X1   g093(.A(KEYINPUT76), .B(G902), .Z(new_n280));
  INV_X1    g094(.A(new_n253), .ZN(new_n281));
  NAND4_X1  g095(.A1(new_n226), .A2(new_n222), .A3(new_n199), .A4(new_n203), .ZN(new_n282));
  AOI21_X1  g096(.A(new_n238), .B1(new_n252), .B2(new_n282), .ZN(new_n283));
  OAI21_X1  g097(.A(KEYINPUT28), .B1(new_n281), .B2(new_n283), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n253), .A2(new_n262), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n285), .A2(KEYINPUT72), .ZN(new_n286));
  NAND3_X1  g100(.A1(new_n253), .A2(new_n261), .A3(new_n262), .ZN(new_n287));
  INV_X1    g101(.A(new_n272), .ZN(new_n288));
  NAND4_X1  g102(.A1(new_n284), .A2(new_n286), .A3(new_n287), .A4(new_n288), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n289), .A2(KEYINPUT73), .ZN(new_n290));
  INV_X1    g104(.A(KEYINPUT73), .ZN(new_n291));
  NAND4_X1  g105(.A1(new_n265), .A2(new_n291), .A3(new_n284), .A4(new_n288), .ZN(new_n292));
  NAND3_X1  g106(.A1(new_n228), .A2(KEYINPUT30), .A3(new_n252), .ZN(new_n293));
  INV_X1    g107(.A(KEYINPUT69), .ZN(new_n294));
  NAND2_X1  g108(.A1(new_n252), .A2(new_n282), .ZN(new_n295));
  INV_X1    g109(.A(KEYINPUT30), .ZN(new_n296));
  AOI21_X1  g110(.A(new_n294), .B1(new_n295), .B2(new_n296), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n293), .A2(new_n297), .ZN(new_n298));
  NAND4_X1  g112(.A1(new_n228), .A2(new_n294), .A3(KEYINPUT30), .A4(new_n252), .ZN(new_n299));
  AOI21_X1  g113(.A(new_n238), .B1(new_n298), .B2(new_n299), .ZN(new_n300));
  OAI21_X1  g114(.A(new_n272), .B1(new_n300), .B2(new_n281), .ZN(new_n301));
  NAND4_X1  g115(.A1(new_n290), .A2(new_n292), .A3(new_n273), .A4(new_n301), .ZN(new_n302));
  NAND3_X1  g116(.A1(new_n279), .A2(new_n280), .A3(new_n302), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n303), .A2(G472), .ZN(new_n304));
  INV_X1    g118(.A(KEYINPUT32), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n265), .A2(new_n284), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n306), .A2(new_n272), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n298), .A2(new_n299), .ZN(new_n308));
  AOI21_X1  g122(.A(new_n281), .B1(new_n308), .B2(new_n237), .ZN(new_n309));
  AOI21_X1  g123(.A(KEYINPUT31), .B1(new_n309), .B2(new_n288), .ZN(new_n310));
  INV_X1    g124(.A(KEYINPUT31), .ZN(new_n311));
  NOR4_X1   g125(.A1(new_n300), .A2(new_n311), .A3(new_n281), .A4(new_n272), .ZN(new_n312));
  OAI21_X1  g126(.A(new_n307), .B1(new_n310), .B2(new_n312), .ZN(new_n313));
  NOR2_X1   g127(.A1(G472), .A2(G902), .ZN(new_n314));
  AOI21_X1  g128(.A(new_n305), .B1(new_n313), .B2(new_n314), .ZN(new_n315));
  AND3_X1   g129(.A1(new_n313), .A2(new_n305), .A3(new_n314), .ZN(new_n316));
  OAI21_X1  g130(.A(new_n304), .B1(new_n315), .B2(new_n316), .ZN(new_n317));
  INV_X1    g131(.A(G104), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n318), .A2(G107), .ZN(new_n319));
  INV_X1    g133(.A(KEYINPUT86), .ZN(new_n320));
  NOR2_X1   g134(.A1(new_n318), .A2(G107), .ZN(new_n321));
  INV_X1    g135(.A(KEYINPUT3), .ZN(new_n322));
  AOI21_X1  g136(.A(new_n320), .B1(new_n321), .B2(new_n322), .ZN(new_n323));
  NOR4_X1   g137(.A1(new_n318), .A2(KEYINPUT86), .A3(KEYINPUT3), .A4(G107), .ZN(new_n324));
  OAI21_X1  g138(.A(new_n319), .B1(new_n323), .B2(new_n324), .ZN(new_n325));
  INV_X1    g139(.A(KEYINPUT85), .ZN(new_n326));
  OAI211_X1 g140(.A(new_n326), .B(KEYINPUT3), .C1(new_n318), .C2(G107), .ZN(new_n327));
  INV_X1    g141(.A(new_n327), .ZN(new_n328));
  INV_X1    g142(.A(G107), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n329), .A2(G104), .ZN(new_n330));
  AOI21_X1  g144(.A(new_n326), .B1(new_n330), .B2(KEYINPUT3), .ZN(new_n331));
  NOR2_X1   g145(.A1(new_n328), .A2(new_n331), .ZN(new_n332));
  OAI21_X1  g146(.A(G101), .B1(new_n325), .B2(new_n332), .ZN(new_n333));
  OAI21_X1  g147(.A(KEYINPUT3), .B1(new_n318), .B2(G107), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n334), .A2(KEYINPUT85), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n335), .A2(new_n327), .ZN(new_n336));
  NAND3_X1  g150(.A1(new_n322), .A2(new_n329), .A3(G104), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n337), .A2(KEYINPUT86), .ZN(new_n338));
  NAND4_X1  g152(.A1(new_n320), .A2(new_n322), .A3(new_n329), .A4(G104), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n338), .A2(new_n339), .ZN(new_n340));
  INV_X1    g154(.A(G101), .ZN(new_n341));
  NAND4_X1  g155(.A1(new_n336), .A2(new_n340), .A3(new_n341), .A4(new_n319), .ZN(new_n342));
  NAND3_X1  g156(.A1(new_n333), .A2(KEYINPUT4), .A3(new_n342), .ZN(new_n343));
  INV_X1    g157(.A(KEYINPUT4), .ZN(new_n344));
  OAI211_X1 g158(.A(new_n344), .B(G101), .C1(new_n325), .C2(new_n332), .ZN(new_n345));
  NAND3_X1  g159(.A1(new_n343), .A2(new_n237), .A3(new_n345), .ZN(new_n346));
  XOR2_X1   g160(.A(KEYINPUT67), .B(G119), .Z(new_n347));
  INV_X1    g161(.A(KEYINPUT5), .ZN(new_n348));
  NAND3_X1  g162(.A1(new_n347), .A2(new_n348), .A3(G116), .ZN(new_n349));
  OAI211_X1 g163(.A(new_n349), .B(G113), .C1(new_n233), .C2(new_n348), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n330), .A2(new_n319), .ZN(new_n351));
  NAND2_X1  g165(.A1(new_n351), .A2(G101), .ZN(new_n352));
  NAND4_X1  g166(.A1(new_n350), .A2(new_n235), .A3(new_n342), .A4(new_n352), .ZN(new_n353));
  NAND2_X1  g167(.A1(new_n346), .A2(new_n353), .ZN(new_n354));
  XOR2_X1   g168(.A(G110), .B(G122), .Z(new_n355));
  NAND2_X1  g169(.A1(new_n354), .A2(new_n355), .ZN(new_n356));
  INV_X1    g170(.A(new_n355), .ZN(new_n357));
  NAND3_X1  g171(.A1(new_n346), .A2(new_n357), .A3(new_n353), .ZN(new_n358));
  NAND3_X1  g172(.A1(new_n356), .A2(KEYINPUT6), .A3(new_n358), .ZN(new_n359));
  NOR3_X1   g173(.A1(new_n205), .A2(new_n206), .A3(new_n197), .ZN(new_n360));
  OAI21_X1  g174(.A(G128), .B1(new_n360), .B2(new_n239), .ZN(new_n361));
  NOR2_X1   g175(.A1(new_n205), .A2(new_n206), .ZN(new_n362));
  AOI21_X1  g176(.A(new_n201), .B1(new_n362), .B2(G143), .ZN(new_n363));
  NOR2_X1   g177(.A1(new_n246), .A2(new_n241), .ZN(new_n364));
  AOI22_X1  g178(.A1(new_n361), .A2(new_n209), .B1(new_n363), .B2(new_n364), .ZN(new_n365));
  XNOR2_X1  g179(.A(KEYINPUT80), .B(G125), .ZN(new_n366));
  INV_X1    g180(.A(new_n366), .ZN(new_n367));
  NAND3_X1  g181(.A1(new_n365), .A2(KEYINPUT88), .A3(new_n367), .ZN(new_n368));
  AOI21_X1  g182(.A(new_n225), .B1(new_n207), .B2(new_n208), .ZN(new_n369));
  AOI22_X1  g183(.A1(new_n369), .A2(new_n188), .B1(new_n363), .B2(new_n189), .ZN(new_n370));
  AOI21_X1  g184(.A(new_n367), .B1(new_n370), .B2(new_n226), .ZN(new_n371));
  INV_X1    g185(.A(KEYINPUT88), .ZN(new_n372));
  OAI21_X1  g186(.A(new_n372), .B1(new_n248), .B2(new_n366), .ZN(new_n373));
  OAI21_X1  g187(.A(new_n368), .B1(new_n371), .B2(new_n373), .ZN(new_n374));
  INV_X1    g188(.A(G953), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n375), .A2(G224), .ZN(new_n376));
  XNOR2_X1  g190(.A(new_n374), .B(new_n376), .ZN(new_n377));
  INV_X1    g191(.A(KEYINPUT6), .ZN(new_n378));
  NAND3_X1  g192(.A1(new_n354), .A2(new_n378), .A3(new_n355), .ZN(new_n379));
  NAND3_X1  g193(.A1(new_n359), .A2(new_n377), .A3(new_n379), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n380), .A2(KEYINPUT89), .ZN(new_n381));
  INV_X1    g195(.A(new_n358), .ZN(new_n382));
  XNOR2_X1  g196(.A(KEYINPUT90), .B(KEYINPUT8), .ZN(new_n383));
  XNOR2_X1  g197(.A(new_n355), .B(new_n383), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n350), .A2(new_n235), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n342), .A2(new_n352), .ZN(new_n386));
  NAND2_X1  g200(.A1(new_n385), .A2(new_n386), .ZN(new_n387));
  AOI21_X1  g201(.A(new_n384), .B1(new_n387), .B2(new_n353), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n376), .A2(KEYINPUT7), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n374), .A2(new_n389), .ZN(new_n390));
  INV_X1    g204(.A(new_n389), .ZN(new_n391));
  OAI211_X1 g205(.A(new_n368), .B(new_n391), .C1(new_n371), .C2(new_n373), .ZN(new_n392));
  AOI21_X1  g206(.A(new_n388), .B1(new_n390), .B2(new_n392), .ZN(new_n393));
  INV_X1    g207(.A(KEYINPUT91), .ZN(new_n394));
  AOI21_X1  g208(.A(new_n382), .B1(new_n393), .B2(new_n394), .ZN(new_n395));
  OAI21_X1  g209(.A(new_n366), .B1(new_n204), .B2(new_n210), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n365), .A2(new_n367), .ZN(new_n397));
  NAND3_X1  g211(.A1(new_n396), .A2(new_n397), .A3(new_n372), .ZN(new_n398));
  AOI21_X1  g212(.A(new_n391), .B1(new_n398), .B2(new_n368), .ZN(new_n399));
  INV_X1    g213(.A(new_n392), .ZN(new_n400));
  AND2_X1   g214(.A1(new_n387), .A2(new_n353), .ZN(new_n401));
  OAI22_X1  g215(.A1(new_n399), .A2(new_n400), .B1(new_n401), .B2(new_n384), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n402), .A2(KEYINPUT91), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n395), .A2(new_n403), .ZN(new_n404));
  INV_X1    g218(.A(G902), .ZN(new_n405));
  INV_X1    g219(.A(KEYINPUT89), .ZN(new_n406));
  NAND4_X1  g220(.A1(new_n359), .A2(new_n377), .A3(new_n406), .A4(new_n379), .ZN(new_n407));
  NAND4_X1  g221(.A1(new_n381), .A2(new_n404), .A3(new_n405), .A4(new_n407), .ZN(new_n408));
  OAI21_X1  g222(.A(G210), .B1(G237), .B2(G902), .ZN(new_n409));
  INV_X1    g223(.A(new_n409), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n408), .A2(new_n410), .ZN(new_n411));
  AOI21_X1  g225(.A(G902), .B1(new_n395), .B2(new_n403), .ZN(new_n412));
  NAND4_X1  g226(.A1(new_n412), .A2(new_n409), .A3(new_n381), .A4(new_n407), .ZN(new_n413));
  NAND3_X1  g227(.A1(new_n411), .A2(KEYINPUT92), .A3(new_n413), .ZN(new_n414));
  INV_X1    g228(.A(KEYINPUT92), .ZN(new_n415));
  NAND3_X1  g229(.A1(new_n408), .A2(new_n415), .A3(new_n410), .ZN(new_n416));
  NAND2_X1  g230(.A1(new_n414), .A2(new_n416), .ZN(new_n417));
  INV_X1    g231(.A(new_n417), .ZN(new_n418));
  INV_X1    g232(.A(G469), .ZN(new_n419));
  XNOR2_X1  g233(.A(G110), .B(G140), .ZN(new_n420));
  XNOR2_X1  g234(.A(new_n420), .B(KEYINPUT84), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n375), .A2(G227), .ZN(new_n422));
  XNOR2_X1  g236(.A(new_n421), .B(new_n422), .ZN(new_n423));
  AOI21_X1  g237(.A(new_n248), .B1(new_n342), .B2(new_n352), .ZN(new_n424));
  AOI21_X1  g238(.A(new_n241), .B1(new_n208), .B2(KEYINPUT1), .ZN(new_n425));
  OAI21_X1  g239(.A(new_n240), .B1(new_n363), .B2(new_n425), .ZN(new_n426));
  AND3_X1   g240(.A1(new_n426), .A2(new_n342), .A3(new_n352), .ZN(new_n427));
  OAI21_X1  g241(.A(new_n222), .B1(new_n424), .B2(new_n427), .ZN(new_n428));
  NAND2_X1  g242(.A1(KEYINPUT87), .A2(KEYINPUT12), .ZN(new_n429));
  INV_X1    g243(.A(KEYINPUT87), .ZN(new_n430));
  INV_X1    g244(.A(KEYINPUT12), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n430), .A2(new_n431), .ZN(new_n432));
  NAND3_X1  g246(.A1(new_n428), .A2(new_n429), .A3(new_n432), .ZN(new_n433));
  NAND4_X1  g247(.A1(new_n343), .A2(new_n211), .A3(new_n227), .A4(new_n345), .ZN(new_n434));
  INV_X1    g248(.A(new_n386), .ZN(new_n435));
  INV_X1    g249(.A(KEYINPUT10), .ZN(new_n436));
  NAND2_X1  g250(.A1(new_n361), .A2(new_n209), .ZN(new_n437));
  AOI21_X1  g251(.A(new_n436), .B1(new_n437), .B2(new_n240), .ZN(new_n438));
  NAND3_X1  g252(.A1(new_n426), .A2(new_n342), .A3(new_n352), .ZN(new_n439));
  AOI22_X1  g253(.A1(new_n435), .A2(new_n438), .B1(new_n439), .B2(new_n436), .ZN(new_n440));
  INV_X1    g254(.A(new_n222), .ZN(new_n441));
  NAND3_X1  g255(.A1(new_n434), .A2(new_n440), .A3(new_n441), .ZN(new_n442));
  OAI21_X1  g256(.A(new_n439), .B1(new_n435), .B2(new_n248), .ZN(new_n443));
  NAND4_X1  g257(.A1(new_n443), .A2(new_n430), .A3(new_n431), .A4(new_n222), .ZN(new_n444));
  AND4_X1   g258(.A1(new_n423), .A2(new_n433), .A3(new_n442), .A4(new_n444), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n434), .A2(new_n440), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n446), .A2(new_n222), .ZN(new_n447));
  AOI21_X1  g261(.A(new_n423), .B1(new_n447), .B2(new_n442), .ZN(new_n448));
  OAI211_X1 g262(.A(new_n419), .B(new_n280), .C1(new_n445), .C2(new_n448), .ZN(new_n449));
  INV_X1    g263(.A(new_n423), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n433), .A2(new_n444), .ZN(new_n451));
  INV_X1    g265(.A(new_n442), .ZN(new_n452));
  OAI21_X1  g266(.A(new_n450), .B1(new_n451), .B2(new_n452), .ZN(new_n453));
  NAND3_X1  g267(.A1(new_n447), .A2(new_n423), .A3(new_n442), .ZN(new_n454));
  NAND3_X1  g268(.A1(new_n453), .A2(G469), .A3(new_n454), .ZN(new_n455));
  NOR2_X1   g269(.A1(new_n419), .A2(new_n405), .ZN(new_n456));
  INV_X1    g270(.A(new_n456), .ZN(new_n457));
  NAND3_X1  g271(.A1(new_n449), .A2(new_n455), .A3(new_n457), .ZN(new_n458));
  OAI21_X1  g272(.A(G214), .B1(G237), .B2(G902), .ZN(new_n459));
  XNOR2_X1  g273(.A(KEYINPUT9), .B(G234), .ZN(new_n460));
  OAI21_X1  g274(.A(G221), .B1(new_n460), .B2(G902), .ZN(new_n461));
  NAND3_X1  g275(.A1(new_n458), .A2(new_n459), .A3(new_n461), .ZN(new_n462));
  XNOR2_X1  g276(.A(G113), .B(G122), .ZN(new_n463));
  XNOR2_X1  g277(.A(new_n463), .B(new_n318), .ZN(new_n464));
  INV_X1    g278(.A(G214), .ZN(new_n465));
  NOR3_X1   g279(.A1(new_n465), .A2(G237), .A3(G953), .ZN(new_n466));
  OAI21_X1  g280(.A(KEYINPUT93), .B1(new_n466), .B2(G143), .ZN(new_n467));
  NAND2_X1  g281(.A1(new_n266), .A2(G214), .ZN(new_n468));
  INV_X1    g282(.A(KEYINPUT93), .ZN(new_n469));
  NAND3_X1  g283(.A1(new_n468), .A2(new_n469), .A3(new_n197), .ZN(new_n470));
  INV_X1    g284(.A(G237), .ZN(new_n471));
  NAND4_X1  g285(.A1(new_n471), .A2(new_n375), .A3(G143), .A4(G214), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n472), .A2(KEYINPUT94), .ZN(new_n473));
  INV_X1    g287(.A(KEYINPUT94), .ZN(new_n474));
  NAND4_X1  g288(.A1(new_n266), .A2(new_n474), .A3(G143), .A4(G214), .ZN(new_n475));
  AOI22_X1  g289(.A1(new_n467), .A2(new_n470), .B1(new_n473), .B2(new_n475), .ZN(new_n476));
  NAND2_X1  g290(.A1(KEYINPUT18), .A2(G131), .ZN(new_n477));
  NOR2_X1   g291(.A1(G125), .A2(G140), .ZN(new_n478));
  AOI21_X1  g292(.A(new_n478), .B1(new_n366), .B2(G140), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n479), .A2(G146), .ZN(new_n480));
  XOR2_X1   g294(.A(G125), .B(G140), .Z(new_n481));
  OR2_X1    g295(.A1(new_n481), .A2(new_n223), .ZN(new_n482));
  AOI22_X1  g296(.A1(new_n476), .A2(new_n477), .B1(new_n480), .B2(new_n482), .ZN(new_n483));
  INV_X1    g297(.A(KEYINPUT18), .ZN(new_n484));
  NOR3_X1   g298(.A1(new_n466), .A2(KEYINPUT93), .A3(G143), .ZN(new_n485));
  AOI21_X1  g299(.A(new_n469), .B1(new_n468), .B2(new_n197), .ZN(new_n486));
  NOR2_X1   g300(.A1(new_n485), .A2(new_n486), .ZN(new_n487));
  AND2_X1   g301(.A1(new_n473), .A2(new_n475), .ZN(new_n488));
  OAI21_X1  g302(.A(G131), .B1(new_n487), .B2(new_n488), .ZN(new_n489));
  OAI21_X1  g303(.A(new_n483), .B1(new_n484), .B2(new_n489), .ZN(new_n490));
  INV_X1    g304(.A(KEYINPUT17), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n476), .A2(new_n220), .ZN(new_n492));
  AND3_X1   g306(.A1(new_n489), .A2(new_n491), .A3(new_n492), .ZN(new_n493));
  OAI211_X1 g307(.A(KEYINPUT17), .B(G131), .C1(new_n487), .C2(new_n488), .ZN(new_n494));
  INV_X1    g308(.A(KEYINPUT16), .ZN(new_n495));
  INV_X1    g309(.A(G140), .ZN(new_n496));
  NAND3_X1  g310(.A1(new_n366), .A2(new_n495), .A3(new_n496), .ZN(new_n497));
  OAI211_X1 g311(.A(G146), .B(new_n497), .C1(new_n479), .C2(new_n495), .ZN(new_n498));
  OAI21_X1  g312(.A(new_n497), .B1(new_n479), .B2(new_n495), .ZN(new_n499));
  NAND2_X1  g313(.A1(new_n499), .A2(new_n193), .ZN(new_n500));
  NAND3_X1  g314(.A1(new_n494), .A2(new_n498), .A3(new_n500), .ZN(new_n501));
  OAI211_X1 g315(.A(new_n464), .B(new_n490), .C1(new_n493), .C2(new_n501), .ZN(new_n502));
  INV_X1    g316(.A(new_n502), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n489), .A2(new_n492), .ZN(new_n504));
  INV_X1    g318(.A(KEYINPUT81), .ZN(new_n505));
  OR2_X1    g319(.A1(new_n498), .A2(new_n505), .ZN(new_n506));
  NAND2_X1  g320(.A1(new_n498), .A2(new_n505), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n479), .A2(KEYINPUT19), .ZN(new_n508));
  OR2_X1    g322(.A1(new_n481), .A2(KEYINPUT19), .ZN(new_n509));
  NAND3_X1  g323(.A1(new_n508), .A2(new_n362), .A3(new_n509), .ZN(new_n510));
  NAND4_X1  g324(.A1(new_n504), .A2(new_n506), .A3(new_n507), .A4(new_n510), .ZN(new_n511));
  AOI21_X1  g325(.A(new_n464), .B1(new_n511), .B2(new_n490), .ZN(new_n512));
  OAI21_X1  g326(.A(KEYINPUT95), .B1(new_n503), .B2(new_n512), .ZN(new_n513));
  NOR2_X1   g327(.A1(G475), .A2(G902), .ZN(new_n514));
  INV_X1    g328(.A(KEYINPUT95), .ZN(new_n515));
  AND2_X1   g329(.A1(new_n508), .A2(new_n509), .ZN(new_n516));
  AOI22_X1  g330(.A1(new_n362), .A2(new_n516), .B1(new_n489), .B2(new_n492), .ZN(new_n517));
  XNOR2_X1  g331(.A(new_n498), .B(KEYINPUT81), .ZN(new_n518));
  OR2_X1    g332(.A1(new_n489), .A2(new_n484), .ZN(new_n519));
  AOI22_X1  g333(.A1(new_n517), .A2(new_n518), .B1(new_n519), .B2(new_n483), .ZN(new_n520));
  OAI211_X1 g334(.A(new_n515), .B(new_n502), .C1(new_n520), .C2(new_n464), .ZN(new_n521));
  NAND3_X1  g335(.A1(new_n513), .A2(new_n514), .A3(new_n521), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n522), .A2(KEYINPUT20), .ZN(new_n523));
  NOR2_X1   g337(.A1(new_n503), .A2(new_n512), .ZN(new_n524));
  INV_X1    g338(.A(KEYINPUT20), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n514), .A2(new_n525), .ZN(new_n526));
  NOR2_X1   g340(.A1(new_n524), .A2(new_n526), .ZN(new_n527));
  INV_X1    g341(.A(new_n527), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n523), .A2(new_n528), .ZN(new_n529));
  INV_X1    g343(.A(G952), .ZN(new_n530));
  AND2_X1   g344(.A1(new_n530), .A2(KEYINPUT101), .ZN(new_n531));
  NOR2_X1   g345(.A1(new_n530), .A2(KEYINPUT101), .ZN(new_n532));
  OAI21_X1  g346(.A(new_n375), .B1(new_n531), .B2(new_n532), .ZN(new_n533));
  INV_X1    g347(.A(new_n533), .ZN(new_n534));
  NAND2_X1  g348(.A1(G234), .A2(G237), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n534), .A2(new_n535), .ZN(new_n536));
  INV_X1    g350(.A(new_n536), .ZN(new_n537));
  INV_X1    g351(.A(new_n280), .ZN(new_n538));
  NAND3_X1  g352(.A1(new_n538), .A2(G953), .A3(new_n535), .ZN(new_n539));
  INV_X1    g353(.A(new_n539), .ZN(new_n540));
  XNOR2_X1  g354(.A(KEYINPUT21), .B(G898), .ZN(new_n541));
  AOI21_X1  g355(.A(new_n537), .B1(new_n540), .B2(new_n541), .ZN(new_n542));
  INV_X1    g356(.A(new_n542), .ZN(new_n543));
  OAI21_X1  g357(.A(new_n490), .B1(new_n493), .B2(new_n501), .ZN(new_n544));
  INV_X1    g358(.A(new_n464), .ZN(new_n545));
  NAND2_X1  g359(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  AOI21_X1  g360(.A(G902), .B1(new_n546), .B2(new_n502), .ZN(new_n547));
  INV_X1    g361(.A(G475), .ZN(new_n548));
  NOR2_X1   g362(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  INV_X1    g363(.A(new_n549), .ZN(new_n550));
  INV_X1    g364(.A(G122), .ZN(new_n551));
  OAI21_X1  g365(.A(KEYINPUT97), .B1(new_n551), .B2(G116), .ZN(new_n552));
  INV_X1    g366(.A(KEYINPUT97), .ZN(new_n553));
  INV_X1    g367(.A(G116), .ZN(new_n554));
  NAND3_X1  g368(.A1(new_n553), .A2(new_n554), .A3(G122), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n552), .A2(new_n555), .ZN(new_n556));
  AND2_X1   g370(.A1(KEYINPUT96), .A2(G122), .ZN(new_n557));
  NOR2_X1   g371(.A1(KEYINPUT96), .A2(G122), .ZN(new_n558));
  OAI21_X1  g372(.A(G116), .B1(new_n557), .B2(new_n558), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n556), .A2(new_n559), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n560), .A2(G107), .ZN(new_n561));
  NAND3_X1  g375(.A1(new_n556), .A2(new_n559), .A3(new_n329), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n563), .A2(KEYINPUT98), .ZN(new_n564));
  INV_X1    g378(.A(KEYINPUT13), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n565), .A2(KEYINPUT99), .ZN(new_n566));
  OAI21_X1  g380(.A(new_n566), .B1(G128), .B2(new_n197), .ZN(new_n567));
  NOR2_X1   g381(.A1(new_n565), .A2(KEYINPUT99), .ZN(new_n568));
  OAI21_X1  g382(.A(G134), .B1(new_n567), .B2(new_n568), .ZN(new_n569));
  XNOR2_X1  g383(.A(G128), .B(G143), .ZN(new_n570));
  INV_X1    g384(.A(new_n570), .ZN(new_n571));
  XNOR2_X1  g385(.A(new_n569), .B(new_n571), .ZN(new_n572));
  INV_X1    g386(.A(KEYINPUT98), .ZN(new_n573));
  NAND3_X1  g387(.A1(new_n561), .A2(new_n573), .A3(new_n562), .ZN(new_n574));
  NAND3_X1  g388(.A1(new_n564), .A2(new_n572), .A3(new_n574), .ZN(new_n575));
  INV_X1    g389(.A(KEYINPUT100), .ZN(new_n576));
  OR2_X1    g390(.A1(new_n557), .A2(new_n558), .ZN(new_n577));
  AOI22_X1  g391(.A1(G116), .A2(new_n577), .B1(new_n556), .B2(KEYINPUT14), .ZN(new_n578));
  INV_X1    g392(.A(KEYINPUT14), .ZN(new_n579));
  NAND3_X1  g393(.A1(new_n552), .A2(new_n555), .A3(new_n579), .ZN(new_n580));
  AOI21_X1  g394(.A(new_n329), .B1(new_n578), .B2(new_n580), .ZN(new_n581));
  XNOR2_X1  g395(.A(new_n570), .B(new_n213), .ZN(new_n582));
  NAND2_X1  g396(.A1(new_n582), .A2(new_n562), .ZN(new_n583));
  OAI21_X1  g397(.A(new_n576), .B1(new_n581), .B2(new_n583), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n556), .A2(KEYINPUT14), .ZN(new_n585));
  NAND3_X1  g399(.A1(new_n585), .A2(new_n559), .A3(new_n580), .ZN(new_n586));
  NAND2_X1  g400(.A1(new_n586), .A2(G107), .ZN(new_n587));
  NAND4_X1  g401(.A1(new_n587), .A2(KEYINPUT100), .A3(new_n562), .A4(new_n582), .ZN(new_n588));
  NAND3_X1  g402(.A1(new_n575), .A2(new_n584), .A3(new_n588), .ZN(new_n589));
  INV_X1    g403(.A(new_n460), .ZN(new_n590));
  XOR2_X1   g404(.A(KEYINPUT77), .B(G217), .Z(new_n591));
  NAND3_X1  g405(.A1(new_n590), .A2(new_n375), .A3(new_n591), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n589), .A2(new_n592), .ZN(new_n593));
  INV_X1    g407(.A(new_n592), .ZN(new_n594));
  NAND4_X1  g408(.A1(new_n575), .A2(new_n584), .A3(new_n588), .A4(new_n594), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n593), .A2(new_n595), .ZN(new_n596));
  NAND2_X1  g410(.A1(new_n596), .A2(new_n280), .ZN(new_n597));
  INV_X1    g411(.A(G478), .ZN(new_n598));
  NOR2_X1   g412(.A1(new_n598), .A2(KEYINPUT15), .ZN(new_n599));
  INV_X1    g413(.A(new_n599), .ZN(new_n600));
  XNOR2_X1  g414(.A(new_n597), .B(new_n600), .ZN(new_n601));
  NAND4_X1  g415(.A1(new_n529), .A2(new_n543), .A3(new_n550), .A4(new_n601), .ZN(new_n602));
  INV_X1    g416(.A(KEYINPUT102), .ZN(new_n603));
  NAND2_X1  g417(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  AOI21_X1  g418(.A(new_n527), .B1(new_n522), .B2(KEYINPUT20), .ZN(new_n605));
  NOR2_X1   g419(.A1(new_n605), .A2(new_n549), .ZN(new_n606));
  NAND4_X1  g420(.A1(new_n606), .A2(KEYINPUT102), .A3(new_n543), .A4(new_n601), .ZN(new_n607));
  AOI21_X1  g421(.A(new_n462), .B1(new_n604), .B2(new_n607), .ZN(new_n608));
  NAND3_X1  g422(.A1(new_n375), .A2(G221), .A3(G234), .ZN(new_n609));
  XNOR2_X1  g423(.A(new_n609), .B(KEYINPUT82), .ZN(new_n610));
  XNOR2_X1  g424(.A(KEYINPUT22), .B(G137), .ZN(new_n611));
  XNOR2_X1  g425(.A(new_n610), .B(new_n611), .ZN(new_n612));
  OAI21_X1  g426(.A(KEYINPUT79), .B1(new_n347), .B2(G128), .ZN(new_n613));
  NAND2_X1  g427(.A1(new_n229), .A2(new_n230), .ZN(new_n614));
  OAI21_X1  g428(.A(KEYINPUT23), .B1(new_n614), .B2(new_n241), .ZN(new_n615));
  INV_X1    g429(.A(KEYINPUT79), .ZN(new_n616));
  NAND3_X1  g430(.A1(new_n614), .A2(new_n616), .A3(new_n241), .ZN(new_n617));
  NAND3_X1  g431(.A1(new_n613), .A2(new_n615), .A3(new_n617), .ZN(new_n618));
  INV_X1    g432(.A(G110), .ZN(new_n619));
  NAND3_X1  g433(.A1(new_n241), .A2(KEYINPUT23), .A3(G119), .ZN(new_n620));
  NAND3_X1  g434(.A1(new_n618), .A2(new_n619), .A3(new_n620), .ZN(new_n621));
  NAND2_X1  g435(.A1(new_n241), .A2(G119), .ZN(new_n622));
  OAI21_X1  g436(.A(new_n622), .B1(new_n614), .B2(new_n241), .ZN(new_n623));
  XNOR2_X1  g437(.A(KEYINPUT24), .B(G110), .ZN(new_n624));
  NAND2_X1  g438(.A1(new_n623), .A2(new_n624), .ZN(new_n625));
  NAND2_X1  g439(.A1(new_n621), .A2(new_n625), .ZN(new_n626));
  NAND3_X1  g440(.A1(new_n518), .A2(new_n626), .A3(new_n482), .ZN(new_n627));
  NAND2_X1  g441(.A1(new_n618), .A2(new_n620), .ZN(new_n628));
  NAND2_X1  g442(.A1(new_n628), .A2(G110), .ZN(new_n629));
  NAND2_X1  g443(.A1(new_n500), .A2(new_n498), .ZN(new_n630));
  OAI211_X1 g444(.A(new_n629), .B(new_n630), .C1(new_n623), .C2(new_n624), .ZN(new_n631));
  AND3_X1   g445(.A1(new_n627), .A2(new_n631), .A3(KEYINPUT83), .ZN(new_n632));
  AOI21_X1  g446(.A(KEYINPUT83), .B1(new_n627), .B2(new_n631), .ZN(new_n633));
  OAI21_X1  g447(.A(new_n612), .B1(new_n632), .B2(new_n633), .ZN(new_n634));
  INV_X1    g448(.A(new_n612), .ZN(new_n635));
  AND2_X1   g449(.A1(new_n627), .A2(new_n631), .ZN(new_n636));
  OAI21_X1  g450(.A(new_n635), .B1(new_n636), .B2(KEYINPUT83), .ZN(new_n637));
  NAND3_X1  g451(.A1(new_n634), .A2(new_n280), .A3(new_n637), .ZN(new_n638));
  NAND2_X1  g452(.A1(new_n638), .A2(KEYINPUT25), .ZN(new_n639));
  INV_X1    g453(.A(G234), .ZN(new_n640));
  OAI21_X1  g454(.A(new_n591), .B1(new_n538), .B2(new_n640), .ZN(new_n641));
  XNOR2_X1  g455(.A(new_n641), .B(KEYINPUT78), .ZN(new_n642));
  INV_X1    g456(.A(KEYINPUT25), .ZN(new_n643));
  NAND4_X1  g457(.A1(new_n634), .A2(new_n637), .A3(new_n643), .A4(new_n280), .ZN(new_n644));
  NAND3_X1  g458(.A1(new_n639), .A2(new_n642), .A3(new_n644), .ZN(new_n645));
  AND2_X1   g459(.A1(new_n634), .A2(new_n637), .ZN(new_n646));
  NOR2_X1   g460(.A1(new_n642), .A2(G902), .ZN(new_n647));
  NAND2_X1  g461(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  NAND2_X1  g462(.A1(new_n645), .A2(new_n648), .ZN(new_n649));
  INV_X1    g463(.A(new_n649), .ZN(new_n650));
  NAND4_X1  g464(.A1(new_n317), .A2(new_n418), .A3(new_n608), .A4(new_n650), .ZN(new_n651));
  XNOR2_X1  g465(.A(new_n651), .B(G101), .ZN(G3));
  AOI21_X1  g466(.A(new_n288), .B1(new_n265), .B2(new_n284), .ZN(new_n653));
  NAND2_X1  g467(.A1(new_n308), .A2(new_n237), .ZN(new_n654));
  NAND3_X1  g468(.A1(new_n654), .A2(new_n253), .A3(new_n288), .ZN(new_n655));
  NAND2_X1  g469(.A1(new_n655), .A2(new_n311), .ZN(new_n656));
  NAND3_X1  g470(.A1(new_n309), .A2(KEYINPUT31), .A3(new_n288), .ZN(new_n657));
  AOI21_X1  g471(.A(new_n653), .B1(new_n656), .B2(new_n657), .ZN(new_n658));
  OAI21_X1  g472(.A(G472), .B1(new_n658), .B2(new_n538), .ZN(new_n659));
  NAND2_X1  g473(.A1(new_n313), .A2(new_n314), .ZN(new_n660));
  AND2_X1   g474(.A1(new_n458), .A2(new_n461), .ZN(new_n661));
  AND4_X1   g475(.A1(new_n650), .A2(new_n659), .A3(new_n660), .A4(new_n661), .ZN(new_n662));
  INV_X1    g476(.A(new_n459), .ZN(new_n663));
  AOI21_X1  g477(.A(new_n663), .B1(new_n411), .B2(new_n413), .ZN(new_n664));
  NOR2_X1   g478(.A1(new_n538), .A2(new_n598), .ZN(new_n665));
  INV_X1    g479(.A(KEYINPUT103), .ZN(new_n666));
  AOI21_X1  g480(.A(KEYINPUT33), .B1(new_n596), .B2(new_n666), .ZN(new_n667));
  INV_X1    g481(.A(KEYINPUT33), .ZN(new_n668));
  AOI211_X1 g482(.A(KEYINPUT103), .B(new_n668), .C1(new_n593), .C2(new_n595), .ZN(new_n669));
  OAI21_X1  g483(.A(new_n665), .B1(new_n667), .B2(new_n669), .ZN(new_n670));
  NAND2_X1  g484(.A1(new_n597), .A2(new_n598), .ZN(new_n671));
  NAND2_X1  g485(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  INV_X1    g486(.A(new_n672), .ZN(new_n673));
  NOR2_X1   g487(.A1(new_n673), .A2(new_n606), .ZN(new_n674));
  AND3_X1   g488(.A1(new_n664), .A2(new_n543), .A3(new_n674), .ZN(new_n675));
  NAND2_X1  g489(.A1(new_n662), .A2(new_n675), .ZN(new_n676));
  XOR2_X1   g490(.A(KEYINPUT34), .B(G104), .Z(new_n677));
  XNOR2_X1  g491(.A(new_n676), .B(new_n677), .ZN(G6));
  XOR2_X1   g492(.A(new_n549), .B(KEYINPUT104), .Z(new_n679));
  INV_X1    g493(.A(new_n601), .ZN(new_n680));
  XNOR2_X1  g494(.A(new_n522), .B(KEYINPUT20), .ZN(new_n681));
  NAND3_X1  g495(.A1(new_n679), .A2(new_n680), .A3(new_n681), .ZN(new_n682));
  INV_X1    g496(.A(new_n682), .ZN(new_n683));
  NAND4_X1  g497(.A1(new_n662), .A2(new_n543), .A3(new_n664), .A4(new_n683), .ZN(new_n684));
  XOR2_X1   g498(.A(KEYINPUT35), .B(G107), .Z(new_n685));
  XNOR2_X1  g499(.A(new_n684), .B(new_n685), .ZN(G9));
  INV_X1    g500(.A(G472), .ZN(new_n687));
  AOI21_X1  g501(.A(new_n687), .B1(new_n313), .B2(new_n280), .ZN(new_n688));
  AOI21_X1  g502(.A(new_n688), .B1(new_n313), .B2(new_n314), .ZN(new_n689));
  NOR2_X1   g503(.A1(new_n612), .A2(KEYINPUT36), .ZN(new_n690));
  XOR2_X1   g504(.A(new_n636), .B(new_n690), .Z(new_n691));
  NAND2_X1  g505(.A1(new_n691), .A2(new_n647), .ZN(new_n692));
  NAND2_X1  g506(.A1(new_n645), .A2(new_n692), .ZN(new_n693));
  NAND4_X1  g507(.A1(new_n418), .A2(new_n608), .A3(new_n689), .A4(new_n693), .ZN(new_n694));
  XOR2_X1   g508(.A(KEYINPUT37), .B(G110), .Z(new_n695));
  XNOR2_X1  g509(.A(new_n694), .B(new_n695), .ZN(G12));
  NAND2_X1  g510(.A1(new_n411), .A2(new_n413), .ZN(new_n697));
  AND4_X1   g511(.A1(new_n697), .A2(new_n459), .A3(new_n661), .A4(new_n693), .ZN(new_n698));
  OAI21_X1  g512(.A(new_n536), .B1(new_n539), .B2(G900), .ZN(new_n699));
  NAND4_X1  g513(.A1(new_n679), .A2(new_n680), .A3(new_n681), .A4(new_n699), .ZN(new_n700));
  INV_X1    g514(.A(new_n700), .ZN(new_n701));
  NAND3_X1  g515(.A1(new_n317), .A2(new_n698), .A3(new_n701), .ZN(new_n702));
  XNOR2_X1  g516(.A(new_n702), .B(G128), .ZN(G30));
  XNOR2_X1  g517(.A(new_n417), .B(KEYINPUT38), .ZN(new_n704));
  XNOR2_X1  g518(.A(new_n699), .B(KEYINPUT39), .ZN(new_n705));
  NAND2_X1  g519(.A1(new_n661), .A2(new_n705), .ZN(new_n706));
  NAND2_X1  g520(.A1(new_n706), .A2(KEYINPUT40), .ZN(new_n707));
  AND2_X1   g521(.A1(new_n644), .A2(new_n642), .ZN(new_n708));
  AOI22_X1  g522(.A1(new_n708), .A2(new_n639), .B1(new_n647), .B2(new_n691), .ZN(new_n709));
  NOR2_X1   g523(.A1(new_n606), .A2(new_n601), .ZN(new_n710));
  NAND4_X1  g524(.A1(new_n707), .A2(new_n459), .A3(new_n709), .A4(new_n710), .ZN(new_n711));
  NOR2_X1   g525(.A1(new_n309), .A2(new_n272), .ZN(new_n712));
  OAI21_X1  g526(.A(new_n405), .B1(new_n259), .B2(new_n288), .ZN(new_n713));
  OAI21_X1  g527(.A(G472), .B1(new_n712), .B2(new_n713), .ZN(new_n714));
  OAI21_X1  g528(.A(new_n714), .B1(new_n316), .B2(new_n315), .ZN(new_n715));
  INV_X1    g529(.A(new_n715), .ZN(new_n716));
  NOR2_X1   g530(.A1(new_n706), .A2(KEYINPUT40), .ZN(new_n717));
  OR4_X1    g531(.A1(new_n704), .A2(new_n711), .A3(new_n716), .A4(new_n717), .ZN(new_n718));
  XNOR2_X1  g532(.A(new_n718), .B(G143), .ZN(G45));
  OAI211_X1 g533(.A(new_n672), .B(new_n699), .C1(new_n605), .C2(new_n549), .ZN(new_n720));
  INV_X1    g534(.A(new_n720), .ZN(new_n721));
  NAND3_X1  g535(.A1(new_n317), .A2(new_n698), .A3(new_n721), .ZN(new_n722));
  XNOR2_X1  g536(.A(new_n722), .B(G146), .ZN(G48));
  INV_X1    g537(.A(new_n314), .ZN(new_n724));
  OAI21_X1  g538(.A(KEYINPUT32), .B1(new_n658), .B2(new_n724), .ZN(new_n725));
  NAND3_X1  g539(.A1(new_n313), .A2(new_n305), .A3(new_n314), .ZN(new_n726));
  NAND2_X1  g540(.A1(new_n725), .A2(new_n726), .ZN(new_n727));
  AOI21_X1  g541(.A(new_n649), .B1(new_n727), .B2(new_n304), .ZN(new_n728));
  OR2_X1    g542(.A1(new_n445), .A2(new_n448), .ZN(new_n729));
  AOI21_X1  g543(.A(new_n419), .B1(new_n729), .B2(new_n280), .ZN(new_n730));
  INV_X1    g544(.A(new_n449), .ZN(new_n731));
  INV_X1    g545(.A(new_n461), .ZN(new_n732));
  NOR3_X1   g546(.A1(new_n730), .A2(new_n731), .A3(new_n732), .ZN(new_n733));
  NAND3_X1  g547(.A1(new_n728), .A2(new_n675), .A3(new_n733), .ZN(new_n734));
  XNOR2_X1  g548(.A(KEYINPUT41), .B(G113), .ZN(new_n735));
  XNOR2_X1  g549(.A(new_n734), .B(new_n735), .ZN(G15));
  AOI22_X1  g550(.A1(new_n725), .A2(new_n726), .B1(new_n303), .B2(G472), .ZN(new_n737));
  NAND2_X1  g551(.A1(new_n664), .A2(new_n733), .ZN(new_n738));
  NOR2_X1   g552(.A1(new_n737), .A2(new_n738), .ZN(new_n739));
  NOR3_X1   g553(.A1(new_n682), .A2(new_n649), .A3(new_n542), .ZN(new_n740));
  NAND2_X1  g554(.A1(new_n739), .A2(new_n740), .ZN(new_n741));
  XOR2_X1   g555(.A(KEYINPUT105), .B(G116), .Z(new_n742));
  XNOR2_X1  g556(.A(new_n741), .B(new_n742), .ZN(G18));
  AOI21_X1  g557(.A(new_n709), .B1(new_n604), .B2(new_n607), .ZN(new_n744));
  NAND2_X1  g558(.A1(new_n739), .A2(new_n744), .ZN(new_n745));
  XNOR2_X1  g559(.A(new_n745), .B(G119), .ZN(G21));
  NAND2_X1  g560(.A1(new_n656), .A2(new_n657), .ZN(new_n747));
  NAND2_X1  g561(.A1(new_n260), .A2(new_n265), .ZN(new_n748));
  NAND2_X1  g562(.A1(new_n748), .A2(new_n272), .ZN(new_n749));
  AOI21_X1  g563(.A(new_n724), .B1(new_n747), .B2(new_n749), .ZN(new_n750));
  NOR3_X1   g564(.A1(new_n688), .A2(new_n750), .A3(new_n649), .ZN(new_n751));
  AND3_X1   g565(.A1(new_n697), .A2(new_n710), .A3(new_n459), .ZN(new_n752));
  NAND4_X1  g566(.A1(new_n751), .A2(new_n752), .A3(new_n543), .A4(new_n733), .ZN(new_n753));
  XNOR2_X1  g567(.A(new_n753), .B(G122), .ZN(G24));
  NOR3_X1   g568(.A1(new_n688), .A2(new_n750), .A3(new_n709), .ZN(new_n755));
  AND3_X1   g569(.A1(new_n697), .A2(new_n733), .A3(new_n459), .ZN(new_n756));
  NAND3_X1  g570(.A1(new_n755), .A2(new_n756), .A3(new_n721), .ZN(new_n757));
  XNOR2_X1  g571(.A(new_n757), .B(G125), .ZN(G27));
  AOI21_X1  g572(.A(new_n462), .B1(new_n414), .B2(new_n416), .ZN(new_n759));
  NAND4_X1  g573(.A1(new_n317), .A2(new_n650), .A3(new_n721), .A4(new_n759), .ZN(new_n760));
  NAND2_X1  g574(.A1(new_n760), .A2(KEYINPUT106), .ZN(new_n761));
  INV_X1    g575(.A(KEYINPUT42), .ZN(new_n762));
  INV_X1    g576(.A(KEYINPUT106), .ZN(new_n763));
  NAND4_X1  g577(.A1(new_n728), .A2(new_n763), .A3(new_n721), .A4(new_n759), .ZN(new_n764));
  NAND4_X1  g578(.A1(new_n761), .A2(KEYINPUT107), .A3(new_n762), .A4(new_n764), .ZN(new_n765));
  OR2_X1    g579(.A1(new_n760), .A2(new_n762), .ZN(new_n766));
  NAND2_X1  g580(.A1(new_n765), .A2(new_n766), .ZN(new_n767));
  AOI21_X1  g581(.A(KEYINPUT42), .B1(new_n760), .B2(KEYINPUT106), .ZN(new_n768));
  AOI21_X1  g582(.A(KEYINPUT107), .B1(new_n768), .B2(new_n764), .ZN(new_n769));
  NOR2_X1   g583(.A1(new_n767), .A2(new_n769), .ZN(new_n770));
  XNOR2_X1  g584(.A(new_n770), .B(new_n220), .ZN(G33));
  INV_X1    g585(.A(new_n759), .ZN(new_n772));
  NOR2_X1   g586(.A1(new_n772), .A2(new_n700), .ZN(new_n773));
  NAND2_X1  g587(.A1(new_n773), .A2(new_n728), .ZN(new_n774));
  XNOR2_X1  g588(.A(new_n774), .B(G134), .ZN(G36));
  AND2_X1   g589(.A1(new_n453), .A2(new_n454), .ZN(new_n776));
  AND2_X1   g590(.A1(new_n776), .A2(KEYINPUT45), .ZN(new_n777));
  OAI21_X1  g591(.A(G469), .B1(new_n776), .B2(KEYINPUT45), .ZN(new_n778));
  OAI21_X1  g592(.A(new_n457), .B1(new_n777), .B2(new_n778), .ZN(new_n779));
  INV_X1    g593(.A(KEYINPUT46), .ZN(new_n780));
  AOI21_X1  g594(.A(new_n731), .B1(new_n779), .B2(new_n780), .ZN(new_n781));
  OAI21_X1  g595(.A(new_n781), .B1(new_n780), .B2(new_n779), .ZN(new_n782));
  NAND3_X1  g596(.A1(new_n782), .A2(new_n461), .A3(new_n705), .ZN(new_n783));
  XOR2_X1   g597(.A(new_n783), .B(KEYINPUT108), .Z(new_n784));
  NAND2_X1  g598(.A1(new_n417), .A2(new_n459), .ZN(new_n785));
  NAND2_X1  g599(.A1(KEYINPUT109), .A2(KEYINPUT43), .ZN(new_n786));
  XNOR2_X1  g600(.A(KEYINPUT109), .B(KEYINPUT43), .ZN(new_n787));
  NAND2_X1  g601(.A1(new_n529), .A2(new_n550), .ZN(new_n788));
  NOR2_X1   g602(.A1(new_n788), .A2(new_n673), .ZN(new_n789));
  MUX2_X1   g603(.A(new_n786), .B(new_n787), .S(new_n789), .Z(new_n790));
  NAND2_X1  g604(.A1(new_n790), .A2(new_n693), .ZN(new_n791));
  NOR2_X1   g605(.A1(new_n791), .A2(new_n689), .ZN(new_n792));
  AOI21_X1  g606(.A(new_n785), .B1(new_n792), .B2(KEYINPUT44), .ZN(new_n793));
  OAI211_X1 g607(.A(new_n784), .B(new_n793), .C1(KEYINPUT44), .C2(new_n792), .ZN(new_n794));
  XNOR2_X1  g608(.A(new_n794), .B(G137), .ZN(G39));
  INV_X1    g609(.A(KEYINPUT110), .ZN(new_n796));
  NAND2_X1  g610(.A1(new_n796), .A2(KEYINPUT47), .ZN(new_n797));
  XOR2_X1   g611(.A(KEYINPUT110), .B(KEYINPUT47), .Z(new_n798));
  NAND2_X1  g612(.A1(new_n782), .A2(new_n461), .ZN(new_n799));
  MUX2_X1   g613(.A(new_n797), .B(new_n798), .S(new_n799), .Z(new_n800));
  INV_X1    g614(.A(new_n785), .ZN(new_n801));
  NAND4_X1  g615(.A1(new_n801), .A2(new_n649), .A3(new_n737), .A4(new_n721), .ZN(new_n802));
  OR2_X1    g616(.A1(new_n800), .A2(new_n802), .ZN(new_n803));
  XNOR2_X1  g617(.A(new_n803), .B(G140), .ZN(G42));
  NOR2_X1   g618(.A1(new_n730), .A2(new_n731), .ZN(new_n805));
  XOR2_X1   g619(.A(new_n805), .B(KEYINPUT49), .Z(new_n806));
  NAND3_X1  g620(.A1(new_n789), .A2(new_n459), .A3(new_n461), .ZN(new_n807));
  NOR2_X1   g621(.A1(new_n806), .A2(new_n807), .ZN(new_n808));
  NAND4_X1  g622(.A1(new_n808), .A2(new_n704), .A3(new_n650), .A4(new_n716), .ZN(new_n809));
  INV_X1    g623(.A(KEYINPUT53), .ZN(new_n810));
  NAND4_X1  g624(.A1(new_n697), .A2(new_n661), .A3(new_n693), .A4(new_n459), .ZN(new_n811));
  NOR3_X1   g625(.A1(new_n737), .A2(new_n811), .A3(new_n700), .ZN(new_n812));
  NAND2_X1  g626(.A1(new_n747), .A2(new_n749), .ZN(new_n813));
  NAND2_X1  g627(.A1(new_n813), .A2(new_n314), .ZN(new_n814));
  NAND4_X1  g628(.A1(new_n659), .A2(new_n814), .A3(new_n721), .A4(new_n693), .ZN(new_n815));
  NOR2_X1   g629(.A1(new_n815), .A2(new_n738), .ZN(new_n816));
  NOR2_X1   g630(.A1(new_n812), .A2(new_n816), .ZN(new_n817));
  NOR2_X1   g631(.A1(new_n737), .A2(new_n811), .ZN(new_n818));
  NAND3_X1  g632(.A1(new_n458), .A2(new_n461), .A3(new_n699), .ZN(new_n819));
  NOR2_X1   g633(.A1(new_n693), .A2(new_n819), .ZN(new_n820));
  AND3_X1   g634(.A1(new_n820), .A2(new_n664), .A3(new_n710), .ZN(new_n821));
  AOI22_X1  g635(.A1(new_n818), .A2(new_n721), .B1(new_n821), .B2(new_n715), .ZN(new_n822));
  INV_X1    g636(.A(KEYINPUT113), .ZN(new_n823));
  NAND3_X1  g637(.A1(new_n817), .A2(new_n822), .A3(new_n823), .ZN(new_n824));
  NAND3_X1  g638(.A1(new_n715), .A2(new_n752), .A3(new_n820), .ZN(new_n825));
  NAND4_X1  g639(.A1(new_n702), .A2(new_n722), .A3(new_n757), .A4(new_n825), .ZN(new_n826));
  NAND2_X1  g640(.A1(new_n826), .A2(KEYINPUT113), .ZN(new_n827));
  NAND2_X1  g641(.A1(new_n824), .A2(new_n827), .ZN(new_n828));
  NAND2_X1  g642(.A1(new_n828), .A2(KEYINPUT52), .ZN(new_n829));
  INV_X1    g643(.A(KEYINPUT52), .ZN(new_n830));
  NAND3_X1  g644(.A1(new_n824), .A2(new_n827), .A3(new_n830), .ZN(new_n831));
  NAND2_X1  g645(.A1(new_n829), .A2(new_n831), .ZN(new_n832));
  AND2_X1   g646(.A1(new_n601), .A2(new_n699), .ZN(new_n833));
  NAND3_X1  g647(.A1(new_n679), .A2(new_n833), .A3(new_n681), .ZN(new_n834));
  NOR3_X1   g648(.A1(new_n737), .A2(new_n709), .A3(new_n834), .ZN(new_n835));
  AOI22_X1  g649(.A1(new_n773), .A2(new_n728), .B1(new_n835), .B2(new_n759), .ZN(new_n836));
  OAI21_X1  g650(.A(KEYINPUT111), .B1(new_n772), .B2(new_n815), .ZN(new_n837));
  INV_X1    g651(.A(KEYINPUT111), .ZN(new_n838));
  NAND4_X1  g652(.A1(new_n755), .A2(new_n759), .A3(new_n838), .A4(new_n721), .ZN(new_n839));
  NAND2_X1  g653(.A1(new_n837), .A2(new_n839), .ZN(new_n840));
  AND2_X1   g654(.A1(new_n836), .A2(new_n840), .ZN(new_n841));
  OAI211_X1 g655(.A(new_n317), .B(new_n756), .C1(new_n740), .C2(new_n744), .ZN(new_n842));
  NAND3_X1  g656(.A1(new_n734), .A2(new_n842), .A3(new_n651), .ZN(new_n843));
  NAND2_X1  g657(.A1(new_n788), .A2(new_n673), .ZN(new_n844));
  NAND2_X1  g658(.A1(new_n606), .A2(new_n601), .ZN(new_n845));
  AND4_X1   g659(.A1(new_n543), .A2(new_n844), .A3(new_n845), .A4(new_n459), .ZN(new_n846));
  NAND3_X1  g660(.A1(new_n662), .A2(new_n418), .A3(new_n846), .ZN(new_n847));
  NAND3_X1  g661(.A1(new_n847), .A2(new_n694), .A3(new_n753), .ZN(new_n848));
  NOR2_X1   g662(.A1(new_n843), .A2(new_n848), .ZN(new_n849));
  OAI211_X1 g663(.A(new_n841), .B(new_n849), .C1(new_n767), .C2(new_n769), .ZN(new_n850));
  OAI21_X1  g664(.A(new_n810), .B1(new_n832), .B2(new_n850), .ZN(new_n851));
  AND3_X1   g665(.A1(new_n734), .A2(new_n842), .A3(new_n651), .ZN(new_n852));
  INV_X1    g666(.A(new_n848), .ZN(new_n853));
  NAND4_X1  g667(.A1(new_n852), .A2(new_n853), .A3(new_n836), .A4(new_n840), .ZN(new_n854));
  AND2_X1   g668(.A1(new_n765), .A2(new_n766), .ZN(new_n855));
  INV_X1    g669(.A(new_n769), .ZN(new_n856));
  AOI21_X1  g670(.A(new_n854), .B1(new_n855), .B2(new_n856), .ZN(new_n857));
  INV_X1    g671(.A(KEYINPUT112), .ZN(new_n858));
  OAI21_X1  g672(.A(new_n858), .B1(new_n812), .B2(new_n816), .ZN(new_n859));
  NAND3_X1  g673(.A1(new_n702), .A2(new_n757), .A3(KEYINPUT112), .ZN(new_n860));
  NAND4_X1  g674(.A1(new_n859), .A2(new_n722), .A3(new_n825), .A4(new_n860), .ZN(new_n861));
  NAND2_X1  g675(.A1(new_n861), .A2(KEYINPUT52), .ZN(new_n862));
  AND2_X1   g676(.A1(new_n862), .A2(new_n831), .ZN(new_n863));
  NAND3_X1  g677(.A1(new_n857), .A2(new_n863), .A3(KEYINPUT53), .ZN(new_n864));
  INV_X1    g678(.A(KEYINPUT54), .ZN(new_n865));
  NAND3_X1  g679(.A1(new_n851), .A2(new_n864), .A3(new_n865), .ZN(new_n866));
  INV_X1    g680(.A(new_n866), .ZN(new_n867));
  AND3_X1   g681(.A1(new_n824), .A2(new_n827), .A3(new_n830), .ZN(new_n868));
  AOI21_X1  g682(.A(new_n830), .B1(new_n824), .B2(new_n827), .ZN(new_n869));
  NOR2_X1   g683(.A1(new_n868), .A2(new_n869), .ZN(new_n870));
  NAND3_X1  g684(.A1(new_n870), .A2(new_n857), .A3(KEYINPUT53), .ZN(new_n871));
  NAND2_X1  g685(.A1(new_n862), .A2(new_n831), .ZN(new_n872));
  NOR2_X1   g686(.A1(new_n850), .A2(new_n872), .ZN(new_n873));
  OAI21_X1  g687(.A(new_n871), .B1(KEYINPUT53), .B2(new_n873), .ZN(new_n874));
  AOI21_X1  g688(.A(new_n867), .B1(KEYINPUT54), .B2(new_n874), .ZN(new_n875));
  INV_X1    g689(.A(KEYINPUT51), .ZN(new_n876));
  NAND3_X1  g690(.A1(new_n704), .A2(new_n663), .A3(new_n733), .ZN(new_n877));
  NAND3_X1  g691(.A1(new_n790), .A2(new_n537), .A3(new_n751), .ZN(new_n878));
  NOR2_X1   g692(.A1(new_n877), .A2(new_n878), .ZN(new_n879));
  XNOR2_X1  g693(.A(new_n879), .B(KEYINPUT50), .ZN(new_n880));
  AND2_X1   g694(.A1(new_n733), .A2(new_n537), .ZN(new_n881));
  AND4_X1   g695(.A1(new_n650), .A2(new_n801), .A3(new_n716), .A4(new_n881), .ZN(new_n882));
  NOR2_X1   g696(.A1(new_n788), .A2(new_n672), .ZN(new_n883));
  AND3_X1   g697(.A1(new_n790), .A2(new_n801), .A3(new_n881), .ZN(new_n884));
  AOI22_X1  g698(.A1(new_n882), .A2(new_n883), .B1(new_n884), .B2(new_n755), .ZN(new_n885));
  NAND2_X1  g699(.A1(new_n880), .A2(new_n885), .ZN(new_n886));
  NAND2_X1  g700(.A1(new_n805), .A2(new_n732), .ZN(new_n887));
  NAND2_X1  g701(.A1(new_n800), .A2(new_n887), .ZN(new_n888));
  NOR2_X1   g702(.A1(new_n878), .A2(new_n785), .ZN(new_n889));
  AND2_X1   g703(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  OAI21_X1  g704(.A(new_n876), .B1(new_n886), .B2(new_n890), .ZN(new_n891));
  OR2_X1    g705(.A1(new_n891), .A2(KEYINPUT114), .ZN(new_n892));
  NAND2_X1  g706(.A1(new_n891), .A2(KEYINPUT114), .ZN(new_n893));
  NAND2_X1  g707(.A1(new_n884), .A2(new_n728), .ZN(new_n894));
  INV_X1    g708(.A(new_n894), .ZN(new_n895));
  OR2_X1    g709(.A1(new_n895), .A2(KEYINPUT116), .ZN(new_n896));
  NAND2_X1  g710(.A1(new_n895), .A2(KEYINPUT116), .ZN(new_n897));
  NAND3_X1  g711(.A1(new_n896), .A2(KEYINPUT48), .A3(new_n897), .ZN(new_n898));
  OAI21_X1  g712(.A(new_n534), .B1(new_n878), .B2(new_n738), .ZN(new_n899));
  AOI21_X1  g713(.A(new_n899), .B1(new_n674), .B2(new_n882), .ZN(new_n900));
  OAI211_X1 g714(.A(new_n898), .B(new_n900), .C1(KEYINPUT48), .C2(new_n896), .ZN(new_n901));
  NOR2_X1   g715(.A1(new_n886), .A2(new_n876), .ZN(new_n902));
  OR2_X1    g716(.A1(new_n888), .A2(KEYINPUT115), .ZN(new_n903));
  NAND2_X1  g717(.A1(new_n888), .A2(KEYINPUT115), .ZN(new_n904));
  NAND3_X1  g718(.A1(new_n903), .A2(new_n889), .A3(new_n904), .ZN(new_n905));
  AOI21_X1  g719(.A(new_n901), .B1(new_n902), .B2(new_n905), .ZN(new_n906));
  AND4_X1   g720(.A1(new_n875), .A2(new_n892), .A3(new_n893), .A4(new_n906), .ZN(new_n907));
  NOR2_X1   g721(.A1(G952), .A2(G953), .ZN(new_n908));
  OAI21_X1  g722(.A(new_n809), .B1(new_n907), .B2(new_n908), .ZN(G75));
  AND2_X1   g723(.A1(new_n359), .A2(new_n379), .ZN(new_n910));
  XOR2_X1   g724(.A(new_n910), .B(KEYINPUT117), .Z(new_n911));
  INV_X1    g725(.A(new_n911), .ZN(new_n912));
  AOI21_X1  g726(.A(new_n280), .B1(new_n851), .B2(new_n864), .ZN(new_n913));
  NAND2_X1  g727(.A1(new_n913), .A2(new_n410), .ZN(new_n914));
  INV_X1    g728(.A(new_n914), .ZN(new_n915));
  OAI21_X1  g729(.A(new_n912), .B1(new_n915), .B2(KEYINPUT56), .ZN(new_n916));
  INV_X1    g730(.A(KEYINPUT56), .ZN(new_n917));
  NAND3_X1  g731(.A1(new_n914), .A2(new_n917), .A3(new_n911), .ZN(new_n918));
  NAND2_X1  g732(.A1(new_n916), .A2(new_n918), .ZN(new_n919));
  XOR2_X1   g733(.A(new_n377), .B(KEYINPUT55), .Z(new_n920));
  INV_X1    g734(.A(new_n920), .ZN(new_n921));
  NAND2_X1  g735(.A1(new_n919), .A2(new_n921), .ZN(new_n922));
  NAND3_X1  g736(.A1(new_n916), .A2(new_n918), .A3(new_n920), .ZN(new_n923));
  NOR2_X1   g737(.A1(new_n375), .A2(G952), .ZN(new_n924));
  INV_X1    g738(.A(new_n924), .ZN(new_n925));
  NAND3_X1  g739(.A1(new_n922), .A2(new_n923), .A3(new_n925), .ZN(new_n926));
  NAND2_X1  g740(.A1(new_n926), .A2(KEYINPUT118), .ZN(new_n927));
  INV_X1    g741(.A(KEYINPUT118), .ZN(new_n928));
  NAND4_X1  g742(.A1(new_n922), .A2(new_n928), .A3(new_n923), .A4(new_n925), .ZN(new_n929));
  NAND2_X1  g743(.A1(new_n927), .A2(new_n929), .ZN(G51));
  XNOR2_X1  g744(.A(new_n456), .B(KEYINPUT57), .ZN(new_n931));
  AND2_X1   g745(.A1(new_n866), .A2(KEYINPUT119), .ZN(new_n932));
  AOI21_X1  g746(.A(KEYINPUT53), .B1(new_n870), .B2(new_n857), .ZN(new_n933));
  NOR3_X1   g747(.A1(new_n850), .A2(new_n872), .A3(new_n810), .ZN(new_n934));
  OAI21_X1  g748(.A(KEYINPUT54), .B1(new_n933), .B2(new_n934), .ZN(new_n935));
  INV_X1    g749(.A(KEYINPUT119), .ZN(new_n936));
  NAND4_X1  g750(.A1(new_n851), .A2(new_n864), .A3(new_n936), .A4(new_n865), .ZN(new_n937));
  NAND2_X1  g751(.A1(new_n935), .A2(new_n937), .ZN(new_n938));
  OAI21_X1  g752(.A(new_n931), .B1(new_n932), .B2(new_n938), .ZN(new_n939));
  INV_X1    g753(.A(KEYINPUT120), .ZN(new_n940));
  NAND3_X1  g754(.A1(new_n939), .A2(new_n940), .A3(new_n729), .ZN(new_n941));
  NOR2_X1   g755(.A1(new_n777), .A2(new_n778), .ZN(new_n942));
  NAND2_X1  g756(.A1(new_n913), .A2(new_n942), .ZN(new_n943));
  NAND2_X1  g757(.A1(new_n941), .A2(new_n943), .ZN(new_n944));
  AOI21_X1  g758(.A(new_n940), .B1(new_n939), .B2(new_n729), .ZN(new_n945));
  OAI21_X1  g759(.A(new_n925), .B1(new_n944), .B2(new_n945), .ZN(new_n946));
  NAND2_X1  g760(.A1(new_n946), .A2(KEYINPUT121), .ZN(new_n947));
  INV_X1    g761(.A(KEYINPUT121), .ZN(new_n948));
  OAI211_X1 g762(.A(new_n948), .B(new_n925), .C1(new_n944), .C2(new_n945), .ZN(new_n949));
  NAND2_X1  g763(.A1(new_n947), .A2(new_n949), .ZN(G54));
  NAND3_X1  g764(.A1(new_n913), .A2(KEYINPUT58), .A3(G475), .ZN(new_n951));
  NAND2_X1  g765(.A1(new_n513), .A2(new_n521), .ZN(new_n952));
  AND2_X1   g766(.A1(new_n951), .A2(new_n952), .ZN(new_n953));
  NOR2_X1   g767(.A1(new_n951), .A2(new_n952), .ZN(new_n954));
  NOR3_X1   g768(.A1(new_n953), .A2(new_n954), .A3(new_n924), .ZN(G60));
  OR2_X1    g769(.A1(new_n667), .A2(new_n669), .ZN(new_n956));
  INV_X1    g770(.A(new_n956), .ZN(new_n957));
  NAND2_X1  g771(.A1(G478), .A2(G902), .ZN(new_n958));
  XOR2_X1   g772(.A(new_n958), .B(KEYINPUT59), .Z(new_n959));
  OAI21_X1  g773(.A(new_n957), .B1(new_n875), .B2(new_n959), .ZN(new_n960));
  INV_X1    g774(.A(KEYINPUT122), .ZN(new_n961));
  OR2_X1    g775(.A1(new_n960), .A2(new_n961), .ZN(new_n962));
  OR2_X1    g776(.A1(new_n932), .A2(new_n938), .ZN(new_n963));
  NOR2_X1   g777(.A1(new_n957), .A2(new_n959), .ZN(new_n964));
  AOI21_X1  g778(.A(new_n924), .B1(new_n963), .B2(new_n964), .ZN(new_n965));
  NAND2_X1  g779(.A1(new_n960), .A2(new_n961), .ZN(new_n966));
  AND3_X1   g780(.A1(new_n962), .A2(new_n965), .A3(new_n966), .ZN(G63));
  NAND2_X1  g781(.A1(new_n851), .A2(new_n864), .ZN(new_n968));
  NAND2_X1  g782(.A1(G217), .A2(G902), .ZN(new_n969));
  XNOR2_X1  g783(.A(new_n969), .B(KEYINPUT123), .ZN(new_n970));
  XNOR2_X1  g784(.A(new_n970), .B(KEYINPUT60), .ZN(new_n971));
  NAND3_X1  g785(.A1(new_n968), .A2(new_n691), .A3(new_n971), .ZN(new_n972));
  XNOR2_X1  g786(.A(new_n972), .B(KEYINPUT124), .ZN(new_n973));
  AOI21_X1  g787(.A(new_n646), .B1(new_n968), .B2(new_n971), .ZN(new_n974));
  NOR3_X1   g788(.A1(new_n973), .A2(new_n924), .A3(new_n974), .ZN(new_n975));
  XNOR2_X1  g789(.A(new_n975), .B(KEYINPUT61), .ZN(G66));
  INV_X1    g790(.A(G224), .ZN(new_n977));
  OAI21_X1  g791(.A(G953), .B1(new_n541), .B2(new_n977), .ZN(new_n978));
  OAI21_X1  g792(.A(new_n978), .B1(new_n849), .B2(G953), .ZN(new_n979));
  OAI21_X1  g793(.A(new_n911), .B1(G898), .B2(new_n375), .ZN(new_n980));
  XNOR2_X1  g794(.A(new_n979), .B(new_n980), .ZN(G69));
  XOR2_X1   g795(.A(new_n308), .B(new_n516), .Z(new_n982));
  AND3_X1   g796(.A1(new_n859), .A2(new_n722), .A3(new_n860), .ZN(new_n983));
  NAND2_X1  g797(.A1(new_n983), .A2(new_n718), .ZN(new_n984));
  XOR2_X1   g798(.A(new_n984), .B(KEYINPUT62), .Z(new_n985));
  INV_X1    g799(.A(new_n728), .ZN(new_n986));
  NAND2_X1  g800(.A1(new_n844), .A2(new_n845), .ZN(new_n987));
  OR4_X1    g801(.A1(new_n986), .A2(new_n706), .A3(new_n785), .A4(new_n987), .ZN(new_n988));
  AND4_X1   g802(.A1(new_n794), .A2(new_n985), .A3(new_n803), .A4(new_n988), .ZN(new_n989));
  OAI21_X1  g803(.A(new_n982), .B1(new_n989), .B2(G953), .ZN(new_n990));
  OR2_X1    g804(.A1(new_n990), .A2(KEYINPUT125), .ZN(new_n991));
  NAND2_X1  g805(.A1(new_n990), .A2(KEYINPUT125), .ZN(new_n992));
  AOI21_X1  g806(.A(new_n982), .B1(G900), .B2(G953), .ZN(new_n993));
  NAND2_X1  g807(.A1(new_n803), .A2(new_n774), .ZN(new_n994));
  OAI21_X1  g808(.A(new_n793), .B1(KEYINPUT44), .B2(new_n792), .ZN(new_n995));
  INV_X1    g809(.A(new_n752), .ZN(new_n996));
  OAI21_X1  g810(.A(new_n995), .B1(new_n986), .B2(new_n996), .ZN(new_n997));
  AOI21_X1  g811(.A(new_n994), .B1(new_n784), .B2(new_n997), .ZN(new_n998));
  OAI211_X1 g812(.A(new_n998), .B(new_n983), .C1(new_n769), .C2(new_n767), .ZN(new_n999));
  OAI21_X1  g813(.A(new_n993), .B1(new_n999), .B2(G953), .ZN(new_n1000));
  NAND3_X1  g814(.A1(new_n991), .A2(new_n992), .A3(new_n1000), .ZN(new_n1001));
  AOI21_X1  g815(.A(new_n375), .B1(G227), .B2(G900), .ZN(new_n1002));
  XNOR2_X1  g816(.A(new_n1001), .B(new_n1002), .ZN(G72));
  NAND2_X1  g817(.A1(new_n309), .A2(new_n272), .ZN(new_n1004));
  INV_X1    g818(.A(new_n1004), .ZN(new_n1005));
  NOR3_X1   g819(.A1(new_n999), .A2(new_n848), .A3(new_n843), .ZN(new_n1006));
  XOR2_X1   g820(.A(KEYINPUT126), .B(KEYINPUT63), .Z(new_n1007));
  NOR2_X1   g821(.A1(new_n687), .A2(new_n405), .ZN(new_n1008));
  XNOR2_X1  g822(.A(new_n1007), .B(new_n1008), .ZN(new_n1009));
  OAI21_X1  g823(.A(new_n1005), .B1(new_n1006), .B2(new_n1009), .ZN(new_n1010));
  AND2_X1   g824(.A1(new_n989), .A2(new_n849), .ZN(new_n1011));
  OAI21_X1  g825(.A(new_n712), .B1(new_n1011), .B2(new_n1009), .ZN(new_n1012));
  NOR3_X1   g826(.A1(new_n1005), .A2(new_n712), .A3(new_n1009), .ZN(new_n1013));
  NAND2_X1  g827(.A1(new_n874), .A2(new_n1013), .ZN(new_n1014));
  NAND4_X1  g828(.A1(new_n1010), .A2(new_n1012), .A3(new_n925), .A4(new_n1014), .ZN(new_n1015));
  XNOR2_X1  g829(.A(new_n1015), .B(KEYINPUT127), .ZN(G57));
endmodule


