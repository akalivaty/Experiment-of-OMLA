//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 0 0 1 0 0 1 1 1 1 1 1 1 0 0 0 0 1 1 1 0 0 1 1 0 1 0 0 0 1 0 0 1 0 1 1 0 1 0 0 1 1 0 1 1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:28:46 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n442, new_n443, new_n444, new_n449, new_n453, new_n454, new_n455,
    new_n456, new_n457, new_n460, new_n461, new_n462, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n516, new_n517, new_n518, new_n519,
    new_n520, new_n521, new_n522, new_n523, new_n524, new_n525, new_n526,
    new_n527, new_n528, new_n529, new_n530, new_n531, new_n532, new_n533,
    new_n534, new_n535, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n544, new_n545, new_n546, new_n547, new_n548, new_n549,
    new_n550, new_n553, new_n554, new_n555, new_n557, new_n558, new_n559,
    new_n560, new_n561, new_n562, new_n563, new_n564, new_n565, new_n566,
    new_n567, new_n568, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n578, new_n579, new_n580, new_n581, new_n582, new_n583, new_n584,
    new_n585, new_n586, new_n587, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n614, new_n617, new_n619,
    new_n620, new_n622, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n837, new_n838, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1199, new_n1200, new_n1201, new_n1202,
    new_n1203, new_n1204;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  INV_X1    g016(.A(G2072), .ZN(new_n442));
  INV_X1    g017(.A(G2078), .ZN(new_n443));
  NOR2_X1   g018(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  NAND3_X1  g019(.A1(new_n444), .A2(G2084), .A3(G2090), .ZN(G158));
  NAND3_X1  g020(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g021(.A(G452), .Z(G391));
  AND2_X1   g022(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g023(.A1(G7), .A2(G661), .ZN(new_n449));
  XOR2_X1   g024(.A(new_n449), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g025(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g026(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g027(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n453));
  XNOR2_X1  g028(.A(new_n453), .B(KEYINPUT2), .ZN(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(new_n455));
  NOR4_X1   g030(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n456));
  INV_X1    g031(.A(new_n456), .ZN(new_n457));
  NOR2_X1   g032(.A1(new_n455), .A2(new_n457), .ZN(G325));
  INV_X1    g033(.A(G325), .ZN(G261));
  NAND2_X1  g034(.A1(new_n455), .A2(G2106), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n457), .A2(G567), .ZN(new_n461));
  NAND2_X1  g036(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  INV_X1    g037(.A(new_n462), .ZN(G319));
  INV_X1    g038(.A(G2104), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n464), .A2(KEYINPUT64), .ZN(new_n465));
  INV_X1    g040(.A(KEYINPUT64), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n466), .A2(G2104), .ZN(new_n467));
  NAND3_X1  g042(.A1(new_n465), .A2(new_n467), .A3(KEYINPUT3), .ZN(new_n468));
  OR2_X1    g043(.A1(new_n464), .A2(KEYINPUT3), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  NOR2_X1   g045(.A1(new_n470), .A2(G2105), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n471), .A2(G137), .ZN(new_n472));
  XNOR2_X1  g047(.A(KEYINPUT3), .B(G2104), .ZN(new_n473));
  AOI22_X1  g048(.A1(new_n473), .A2(G125), .B1(G113), .B2(G2104), .ZN(new_n474));
  INV_X1    g049(.A(G2105), .ZN(new_n475));
  OR2_X1    g050(.A1(new_n474), .A2(new_n475), .ZN(new_n476));
  AOI21_X1  g051(.A(G2105), .B1(new_n465), .B2(new_n467), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n477), .A2(G101), .ZN(new_n478));
  AND3_X1   g053(.A1(new_n472), .A2(new_n476), .A3(new_n478), .ZN(G160));
  NAND2_X1  g054(.A1(new_n471), .A2(G136), .ZN(new_n480));
  NOR2_X1   g055(.A1(new_n470), .A2(new_n475), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n481), .A2(G124), .ZN(new_n482));
  OR2_X1    g057(.A1(G100), .A2(G2105), .ZN(new_n483));
  OAI211_X1 g058(.A(new_n483), .B(G2104), .C1(G112), .C2(new_n475), .ZN(new_n484));
  NAND3_X1  g059(.A1(new_n480), .A2(new_n482), .A3(new_n484), .ZN(new_n485));
  INV_X1    g060(.A(new_n485), .ZN(G162));
  INV_X1    g061(.A(KEYINPUT4), .ZN(new_n487));
  AND2_X1   g062(.A1(new_n475), .A2(G138), .ZN(new_n488));
  NAND3_X1  g063(.A1(new_n473), .A2(new_n487), .A3(new_n488), .ZN(new_n489));
  NAND3_X1  g064(.A1(new_n468), .A2(new_n469), .A3(new_n488), .ZN(new_n490));
  AND3_X1   g065(.A1(new_n490), .A2(KEYINPUT65), .A3(KEYINPUT4), .ZN(new_n491));
  AOI21_X1  g066(.A(KEYINPUT65), .B1(new_n490), .B2(KEYINPUT4), .ZN(new_n492));
  OAI21_X1  g067(.A(new_n489), .B1(new_n491), .B2(new_n492), .ZN(new_n493));
  NAND4_X1  g068(.A1(new_n468), .A2(G126), .A3(G2105), .A4(new_n469), .ZN(new_n494));
  OR2_X1    g069(.A1(G102), .A2(G2105), .ZN(new_n495));
  OAI211_X1 g070(.A(new_n495), .B(G2104), .C1(G114), .C2(new_n475), .ZN(new_n496));
  NAND2_X1  g071(.A1(new_n494), .A2(new_n496), .ZN(new_n497));
  INV_X1    g072(.A(new_n497), .ZN(new_n498));
  NAND2_X1  g073(.A1(new_n493), .A2(new_n498), .ZN(new_n499));
  INV_X1    g074(.A(new_n499), .ZN(G164));
  XNOR2_X1  g075(.A(KEYINPUT5), .B(G543), .ZN(new_n501));
  AOI22_X1  g076(.A1(new_n501), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n502));
  INV_X1    g077(.A(G651), .ZN(new_n503));
  OR2_X1    g078(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  INV_X1    g079(.A(G50), .ZN(new_n505));
  XNOR2_X1  g080(.A(KEYINPUT6), .B(G651), .ZN(new_n506));
  NAND2_X1  g081(.A1(new_n506), .A2(G543), .ZN(new_n507));
  NAND2_X1  g082(.A1(new_n506), .A2(new_n501), .ZN(new_n508));
  INV_X1    g083(.A(KEYINPUT66), .ZN(new_n509));
  NAND2_X1  g084(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  NAND3_X1  g085(.A1(new_n506), .A2(new_n501), .A3(KEYINPUT66), .ZN(new_n511));
  NAND2_X1  g086(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  INV_X1    g087(.A(G88), .ZN(new_n513));
  OAI221_X1 g088(.A(new_n504), .B1(new_n505), .B2(new_n507), .C1(new_n512), .C2(new_n513), .ZN(G303));
  INV_X1    g089(.A(G303), .ZN(G166));
  INV_X1    g090(.A(KEYINPUT67), .ZN(new_n516));
  XNOR2_X1  g091(.A(new_n501), .B(new_n516), .ZN(new_n517));
  NAND3_X1  g092(.A1(new_n517), .A2(G63), .A3(G651), .ZN(new_n518));
  INV_X1    g093(.A(KEYINPUT68), .ZN(new_n519));
  XNOR2_X1  g094(.A(new_n518), .B(new_n519), .ZN(new_n520));
  INV_X1    g095(.A(new_n511), .ZN(new_n521));
  AOI21_X1  g096(.A(KEYINPUT66), .B1(new_n506), .B2(new_n501), .ZN(new_n522));
  NOR2_X1   g097(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  NAND2_X1  g098(.A1(new_n523), .A2(G89), .ZN(new_n524));
  INV_X1    g099(.A(new_n507), .ZN(new_n525));
  XOR2_X1   g100(.A(KEYINPUT69), .B(G51), .Z(new_n526));
  NAND3_X1  g101(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n527));
  NAND2_X1  g102(.A1(new_n527), .A2(KEYINPUT7), .ZN(new_n528));
  OR2_X1    g103(.A1(new_n527), .A2(KEYINPUT7), .ZN(new_n529));
  AOI22_X1  g104(.A1(new_n525), .A2(new_n526), .B1(new_n528), .B2(new_n529), .ZN(new_n530));
  NAND2_X1  g105(.A1(new_n524), .A2(new_n530), .ZN(new_n531));
  OAI21_X1  g106(.A(KEYINPUT70), .B1(new_n520), .B2(new_n531), .ZN(new_n532));
  XNOR2_X1  g107(.A(new_n518), .B(KEYINPUT68), .ZN(new_n533));
  INV_X1    g108(.A(KEYINPUT70), .ZN(new_n534));
  NAND4_X1  g109(.A1(new_n533), .A2(new_n534), .A3(new_n524), .A4(new_n530), .ZN(new_n535));
  NAND2_X1  g110(.A1(new_n532), .A2(new_n535), .ZN(G168));
  NAND2_X1  g111(.A1(new_n517), .A2(G64), .ZN(new_n537));
  NAND2_X1  g112(.A1(G77), .A2(G543), .ZN(new_n538));
  AOI21_X1  g113(.A(new_n503), .B1(new_n537), .B2(new_n538), .ZN(new_n539));
  NAND2_X1  g114(.A1(new_n525), .A2(G52), .ZN(new_n540));
  INV_X1    g115(.A(G90), .ZN(new_n541));
  OAI21_X1  g116(.A(new_n540), .B1(new_n512), .B2(new_n541), .ZN(new_n542));
  NOR2_X1   g117(.A1(new_n539), .A2(new_n542), .ZN(G171));
  NAND2_X1  g118(.A1(new_n517), .A2(G56), .ZN(new_n544));
  NAND2_X1  g119(.A1(G68), .A2(G543), .ZN(new_n545));
  AOI21_X1  g120(.A(new_n503), .B1(new_n544), .B2(new_n545), .ZN(new_n546));
  NAND2_X1  g121(.A1(new_n525), .A2(G43), .ZN(new_n547));
  INV_X1    g122(.A(G81), .ZN(new_n548));
  OAI21_X1  g123(.A(new_n547), .B1(new_n512), .B2(new_n548), .ZN(new_n549));
  NOR2_X1   g124(.A1(new_n546), .A2(new_n549), .ZN(new_n550));
  NAND2_X1  g125(.A1(new_n550), .A2(G860), .ZN(G153));
  NAND4_X1  g126(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g127(.A1(G1), .A2(G3), .ZN(new_n553));
  XNOR2_X1  g128(.A(new_n553), .B(KEYINPUT71), .ZN(new_n554));
  XNOR2_X1  g129(.A(new_n554), .B(KEYINPUT8), .ZN(new_n555));
  NAND4_X1  g130(.A1(G319), .A2(G483), .A3(G661), .A4(new_n555), .ZN(G188));
  OAI21_X1  g131(.A(KEYINPUT72), .B1(new_n521), .B2(new_n522), .ZN(new_n557));
  INV_X1    g132(.A(KEYINPUT72), .ZN(new_n558));
  NAND3_X1  g133(.A1(new_n510), .A2(new_n558), .A3(new_n511), .ZN(new_n559));
  NAND3_X1  g134(.A1(new_n557), .A2(new_n559), .A3(G91), .ZN(new_n560));
  NAND2_X1  g135(.A1(new_n501), .A2(G65), .ZN(new_n561));
  NAND2_X1  g136(.A1(G78), .A2(G543), .ZN(new_n562));
  XNOR2_X1  g137(.A(new_n562), .B(KEYINPUT73), .ZN(new_n563));
  AOI21_X1  g138(.A(new_n503), .B1(new_n561), .B2(new_n563), .ZN(new_n564));
  INV_X1    g139(.A(G53), .ZN(new_n565));
  OR3_X1    g140(.A1(new_n507), .A2(KEYINPUT9), .A3(new_n565), .ZN(new_n566));
  OAI21_X1  g141(.A(KEYINPUT9), .B1(new_n507), .B2(new_n565), .ZN(new_n567));
  AOI21_X1  g142(.A(new_n564), .B1(new_n566), .B2(new_n567), .ZN(new_n568));
  NAND2_X1  g143(.A1(new_n560), .A2(new_n568), .ZN(G299));
  INV_X1    g144(.A(G171), .ZN(G301));
  INV_X1    g145(.A(G168), .ZN(G286));
  XNOR2_X1  g146(.A(new_n501), .B(KEYINPUT67), .ZN(new_n572));
  INV_X1    g147(.A(G74), .ZN(new_n573));
  NAND2_X1  g148(.A1(new_n572), .A2(new_n573), .ZN(new_n574));
  AOI22_X1  g149(.A1(new_n574), .A2(G651), .B1(G49), .B2(new_n525), .ZN(new_n575));
  NAND3_X1  g150(.A1(new_n557), .A2(new_n559), .A3(G87), .ZN(new_n576));
  NAND2_X1  g151(.A1(new_n575), .A2(new_n576), .ZN(G288));
  NAND2_X1  g152(.A1(new_n557), .A2(new_n559), .ZN(new_n578));
  INV_X1    g153(.A(G86), .ZN(new_n579));
  OAI21_X1  g154(.A(KEYINPUT74), .B1(new_n578), .B2(new_n579), .ZN(new_n580));
  INV_X1    g155(.A(KEYINPUT74), .ZN(new_n581));
  NAND4_X1  g156(.A1(new_n557), .A2(new_n559), .A3(new_n581), .A4(G86), .ZN(new_n582));
  NAND2_X1  g157(.A1(new_n580), .A2(new_n582), .ZN(new_n583));
  AOI22_X1  g158(.A1(new_n501), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n584));
  INV_X1    g159(.A(G48), .ZN(new_n585));
  OAI22_X1  g160(.A1(new_n584), .A2(new_n503), .B1(new_n585), .B2(new_n507), .ZN(new_n586));
  INV_X1    g161(.A(new_n586), .ZN(new_n587));
  NAND2_X1  g162(.A1(new_n583), .A2(new_n587), .ZN(G305));
  AOI22_X1  g163(.A1(new_n523), .A2(G85), .B1(G47), .B2(new_n525), .ZN(new_n589));
  NAND2_X1  g164(.A1(G72), .A2(G543), .ZN(new_n590));
  INV_X1    g165(.A(G60), .ZN(new_n591));
  OAI21_X1  g166(.A(new_n590), .B1(new_n572), .B2(new_n591), .ZN(new_n592));
  NAND2_X1  g167(.A1(new_n592), .A2(G651), .ZN(new_n593));
  INV_X1    g168(.A(new_n593), .ZN(new_n594));
  OAI21_X1  g169(.A(new_n589), .B1(new_n594), .B2(KEYINPUT75), .ZN(new_n595));
  INV_X1    g170(.A(KEYINPUT75), .ZN(new_n596));
  NOR2_X1   g171(.A1(new_n593), .A2(new_n596), .ZN(new_n597));
  NOR2_X1   g172(.A1(new_n595), .A2(new_n597), .ZN(new_n598));
  INV_X1    g173(.A(new_n598), .ZN(G290));
  NAND2_X1  g174(.A1(G301), .A2(G868), .ZN(new_n600));
  INV_X1    g175(.A(KEYINPUT10), .ZN(new_n601));
  INV_X1    g176(.A(G92), .ZN(new_n602));
  OAI21_X1  g177(.A(new_n601), .B1(new_n578), .B2(new_n602), .ZN(new_n603));
  NAND4_X1  g178(.A1(new_n557), .A2(new_n559), .A3(KEYINPUT10), .A4(G92), .ZN(new_n604));
  NAND2_X1  g179(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  XNOR2_X1  g180(.A(KEYINPUT76), .B(G66), .ZN(new_n606));
  AOI22_X1  g181(.A1(new_n501), .A2(new_n606), .B1(G79), .B2(G543), .ZN(new_n607));
  INV_X1    g182(.A(new_n607), .ZN(new_n608));
  AOI22_X1  g183(.A1(new_n608), .A2(G651), .B1(G54), .B2(new_n525), .ZN(new_n609));
  NAND2_X1  g184(.A1(new_n605), .A2(new_n609), .ZN(new_n610));
  INV_X1    g185(.A(new_n610), .ZN(new_n611));
  OAI21_X1  g186(.A(new_n600), .B1(new_n611), .B2(G868), .ZN(G284));
  XNOR2_X1  g187(.A(G284), .B(KEYINPUT77), .ZN(G321));
  NOR2_X1   g188(.A1(G299), .A2(G868), .ZN(new_n614));
  AOI21_X1  g189(.A(new_n614), .B1(G168), .B2(G868), .ZN(G297));
  XOR2_X1   g190(.A(G297), .B(KEYINPUT78), .Z(G280));
  INV_X1    g191(.A(G559), .ZN(new_n617));
  OAI21_X1  g192(.A(new_n611), .B1(new_n617), .B2(G860), .ZN(G148));
  NAND2_X1  g193(.A1(new_n611), .A2(new_n617), .ZN(new_n619));
  NAND2_X1  g194(.A1(new_n619), .A2(G868), .ZN(new_n620));
  OAI21_X1  g195(.A(new_n620), .B1(G868), .B2(new_n550), .ZN(G323));
  XOR2_X1   g196(.A(KEYINPUT79), .B(KEYINPUT11), .Z(new_n622));
  XNOR2_X1  g197(.A(G323), .B(new_n622), .ZN(G282));
  NAND2_X1  g198(.A1(new_n477), .A2(new_n473), .ZN(new_n624));
  XOR2_X1   g199(.A(new_n624), .B(KEYINPUT12), .Z(new_n625));
  XNOR2_X1  g200(.A(new_n625), .B(KEYINPUT13), .ZN(new_n626));
  OR2_X1    g201(.A1(new_n626), .A2(G2100), .ZN(new_n627));
  NAND2_X1  g202(.A1(new_n481), .A2(G123), .ZN(new_n628));
  OR2_X1    g203(.A1(G99), .A2(G2105), .ZN(new_n629));
  OAI211_X1 g204(.A(new_n629), .B(G2104), .C1(G111), .C2(new_n475), .ZN(new_n630));
  NAND2_X1  g205(.A1(new_n628), .A2(new_n630), .ZN(new_n631));
  AOI21_X1  g206(.A(new_n631), .B1(G135), .B2(new_n471), .ZN(new_n632));
  XNOR2_X1  g207(.A(new_n632), .B(G2096), .ZN(new_n633));
  NAND2_X1  g208(.A1(new_n626), .A2(G2100), .ZN(new_n634));
  NAND3_X1  g209(.A1(new_n627), .A2(new_n633), .A3(new_n634), .ZN(new_n635));
  XOR2_X1   g210(.A(new_n635), .B(KEYINPUT80), .Z(G156));
  XNOR2_X1  g211(.A(G2427), .B(G2438), .ZN(new_n637));
  XNOR2_X1  g212(.A(new_n637), .B(G2430), .ZN(new_n638));
  XNOR2_X1  g213(.A(KEYINPUT15), .B(G2435), .ZN(new_n639));
  OR2_X1    g214(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  NAND2_X1  g215(.A1(new_n638), .A2(new_n639), .ZN(new_n641));
  NAND3_X1  g216(.A1(new_n640), .A2(KEYINPUT14), .A3(new_n641), .ZN(new_n642));
  XOR2_X1   g217(.A(G2443), .B(G2446), .Z(new_n643));
  XNOR2_X1  g218(.A(new_n642), .B(new_n643), .ZN(new_n644));
  XOR2_X1   g219(.A(KEYINPUT81), .B(KEYINPUT16), .Z(new_n645));
  XNOR2_X1  g220(.A(new_n645), .B(KEYINPUT82), .ZN(new_n646));
  XOR2_X1   g221(.A(G2451), .B(G2454), .Z(new_n647));
  XNOR2_X1  g222(.A(new_n646), .B(new_n647), .ZN(new_n648));
  XNOR2_X1  g223(.A(new_n644), .B(new_n648), .ZN(new_n649));
  XNOR2_X1  g224(.A(G1341), .B(G1348), .ZN(new_n650));
  XNOR2_X1  g225(.A(new_n650), .B(KEYINPUT83), .ZN(new_n651));
  OAI21_X1  g226(.A(G14), .B1(new_n649), .B2(new_n651), .ZN(new_n652));
  NAND2_X1  g227(.A1(new_n649), .A2(new_n651), .ZN(new_n653));
  NAND2_X1  g228(.A1(new_n653), .A2(KEYINPUT84), .ZN(new_n654));
  INV_X1    g229(.A(KEYINPUT84), .ZN(new_n655));
  NAND3_X1  g230(.A1(new_n649), .A2(new_n655), .A3(new_n651), .ZN(new_n656));
  AOI21_X1  g231(.A(new_n652), .B1(new_n654), .B2(new_n656), .ZN(G401));
  XOR2_X1   g232(.A(G2084), .B(G2090), .Z(new_n658));
  XNOR2_X1  g233(.A(G2067), .B(G2678), .ZN(new_n659));
  XNOR2_X1  g234(.A(new_n659), .B(KEYINPUT85), .ZN(new_n660));
  NOR2_X1   g235(.A1(G2072), .A2(G2078), .ZN(new_n661));
  NOR2_X1   g236(.A1(new_n444), .A2(new_n661), .ZN(new_n662));
  AOI21_X1  g237(.A(new_n658), .B1(new_n660), .B2(new_n662), .ZN(new_n663));
  XNOR2_X1  g238(.A(new_n662), .B(KEYINPUT17), .ZN(new_n664));
  OAI21_X1  g239(.A(new_n663), .B1(new_n660), .B2(new_n664), .ZN(new_n665));
  OAI211_X1 g240(.A(new_n658), .B(new_n659), .C1(new_n444), .C2(new_n661), .ZN(new_n666));
  XOR2_X1   g241(.A(new_n666), .B(KEYINPUT18), .Z(new_n667));
  NAND3_X1  g242(.A1(new_n664), .A2(new_n660), .A3(new_n658), .ZN(new_n668));
  NAND3_X1  g243(.A1(new_n665), .A2(new_n667), .A3(new_n668), .ZN(new_n669));
  XOR2_X1   g244(.A(G2096), .B(G2100), .Z(new_n670));
  XNOR2_X1  g245(.A(new_n669), .B(new_n670), .ZN(G227));
  XOR2_X1   g246(.A(G1971), .B(G1976), .Z(new_n672));
  XNOR2_X1  g247(.A(KEYINPUT86), .B(KEYINPUT19), .ZN(new_n673));
  XNOR2_X1  g248(.A(new_n672), .B(new_n673), .ZN(new_n674));
  XNOR2_X1  g249(.A(G1956), .B(G2474), .ZN(new_n675));
  XNOR2_X1  g250(.A(G1961), .B(G1966), .ZN(new_n676));
  NOR2_X1   g251(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  INV_X1    g252(.A(new_n677), .ZN(new_n678));
  NOR2_X1   g253(.A1(new_n674), .A2(new_n678), .ZN(new_n679));
  XOR2_X1   g254(.A(new_n679), .B(KEYINPUT20), .Z(new_n680));
  NAND2_X1  g255(.A1(new_n675), .A2(new_n676), .ZN(new_n681));
  NAND3_X1  g256(.A1(new_n674), .A2(new_n678), .A3(new_n681), .ZN(new_n682));
  OR2_X1    g257(.A1(new_n674), .A2(new_n681), .ZN(new_n683));
  NAND3_X1  g258(.A1(new_n680), .A2(new_n682), .A3(new_n683), .ZN(new_n684));
  XNOR2_X1  g259(.A(new_n684), .B(G1981), .ZN(new_n685));
  XNOR2_X1  g260(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n686));
  XNOR2_X1  g261(.A(new_n686), .B(KEYINPUT87), .ZN(new_n687));
  XOR2_X1   g262(.A(G1991), .B(G1996), .Z(new_n688));
  XNOR2_X1  g263(.A(new_n687), .B(new_n688), .ZN(new_n689));
  XNOR2_X1  g264(.A(new_n685), .B(new_n689), .ZN(new_n690));
  XNOR2_X1  g265(.A(KEYINPUT88), .B(G1986), .ZN(new_n691));
  XNOR2_X1  g266(.A(new_n690), .B(new_n691), .ZN(new_n692));
  INV_X1    g267(.A(new_n692), .ZN(G229));
  NOR2_X1   g268(.A1(G16), .A2(G23), .ZN(new_n694));
  NAND2_X1  g269(.A1(G288), .A2(KEYINPUT90), .ZN(new_n695));
  INV_X1    g270(.A(KEYINPUT90), .ZN(new_n696));
  NAND3_X1  g271(.A1(new_n575), .A2(new_n696), .A3(new_n576), .ZN(new_n697));
  AND2_X1   g272(.A1(new_n695), .A2(new_n697), .ZN(new_n698));
  AOI21_X1  g273(.A(new_n694), .B1(new_n698), .B2(G16), .ZN(new_n699));
  XOR2_X1   g274(.A(KEYINPUT33), .B(G1976), .Z(new_n700));
  OR2_X1    g275(.A1(new_n699), .A2(new_n700), .ZN(new_n701));
  NAND2_X1  g276(.A1(new_n699), .A2(new_n700), .ZN(new_n702));
  INV_X1    g277(.A(G16), .ZN(new_n703));
  OR2_X1    g278(.A1(new_n703), .A2(KEYINPUT89), .ZN(new_n704));
  NAND2_X1  g279(.A1(new_n703), .A2(KEYINPUT89), .ZN(new_n705));
  NAND2_X1  g280(.A1(new_n704), .A2(new_n705), .ZN(new_n706));
  NOR2_X1   g281(.A1(new_n706), .A2(G22), .ZN(new_n707));
  AOI21_X1  g282(.A(new_n707), .B1(G166), .B2(new_n706), .ZN(new_n708));
  XNOR2_X1  g283(.A(KEYINPUT91), .B(G1971), .ZN(new_n709));
  XNOR2_X1  g284(.A(new_n708), .B(new_n709), .ZN(new_n710));
  NAND3_X1  g285(.A1(new_n701), .A2(new_n702), .A3(new_n710), .ZN(new_n711));
  NAND2_X1  g286(.A1(new_n703), .A2(G6), .ZN(new_n712));
  AOI21_X1  g287(.A(new_n586), .B1(new_n580), .B2(new_n582), .ZN(new_n713));
  OAI21_X1  g288(.A(new_n712), .B1(new_n713), .B2(new_n703), .ZN(new_n714));
  XNOR2_X1  g289(.A(KEYINPUT32), .B(G1981), .ZN(new_n715));
  XNOR2_X1  g290(.A(new_n714), .B(new_n715), .ZN(new_n716));
  OAI21_X1  g291(.A(KEYINPUT92), .B1(new_n711), .B2(new_n716), .ZN(new_n717));
  AND2_X1   g292(.A1(new_n702), .A2(new_n710), .ZN(new_n718));
  INV_X1    g293(.A(KEYINPUT92), .ZN(new_n719));
  INV_X1    g294(.A(new_n716), .ZN(new_n720));
  NAND4_X1  g295(.A1(new_n718), .A2(new_n719), .A3(new_n720), .A4(new_n701), .ZN(new_n721));
  NAND2_X1  g296(.A1(new_n717), .A2(new_n721), .ZN(new_n722));
  INV_X1    g297(.A(KEYINPUT34), .ZN(new_n723));
  NAND2_X1  g298(.A1(new_n722), .A2(new_n723), .ZN(new_n724));
  NAND3_X1  g299(.A1(new_n717), .A2(KEYINPUT34), .A3(new_n721), .ZN(new_n725));
  NOR2_X1   g300(.A1(new_n706), .A2(G24), .ZN(new_n726));
  AOI21_X1  g301(.A(new_n726), .B1(new_n598), .B2(new_n706), .ZN(new_n727));
  XNOR2_X1  g302(.A(new_n727), .B(G1986), .ZN(new_n728));
  NAND2_X1  g303(.A1(new_n471), .A2(G131), .ZN(new_n729));
  NAND2_X1  g304(.A1(new_n481), .A2(G119), .ZN(new_n730));
  NOR2_X1   g305(.A1(new_n475), .A2(G107), .ZN(new_n731));
  OAI21_X1  g306(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n732));
  OAI211_X1 g307(.A(new_n729), .B(new_n730), .C1(new_n731), .C2(new_n732), .ZN(new_n733));
  MUX2_X1   g308(.A(G25), .B(new_n733), .S(G29), .Z(new_n734));
  XOR2_X1   g309(.A(KEYINPUT35), .B(G1991), .Z(new_n735));
  INV_X1    g310(.A(new_n735), .ZN(new_n736));
  XNOR2_X1  g311(.A(new_n734), .B(new_n736), .ZN(new_n737));
  NOR3_X1   g312(.A1(new_n728), .A2(KEYINPUT93), .A3(new_n737), .ZN(new_n738));
  NAND3_X1  g313(.A1(new_n724), .A2(new_n725), .A3(new_n738), .ZN(new_n739));
  NAND2_X1  g314(.A1(new_n739), .A2(KEYINPUT36), .ZN(new_n740));
  INV_X1    g315(.A(KEYINPUT36), .ZN(new_n741));
  NAND4_X1  g316(.A1(new_n724), .A2(new_n741), .A3(new_n725), .A4(new_n738), .ZN(new_n742));
  NAND3_X1  g317(.A1(new_n704), .A2(G20), .A3(new_n705), .ZN(new_n743));
  XOR2_X1   g318(.A(new_n743), .B(KEYINPUT23), .Z(new_n744));
  AOI21_X1  g319(.A(new_n744), .B1(G299), .B2(G16), .ZN(new_n745));
  XNOR2_X1  g320(.A(new_n745), .B(G1956), .ZN(new_n746));
  INV_X1    g321(.A(G29), .ZN(new_n747));
  NAND2_X1  g322(.A1(new_n747), .A2(G35), .ZN(new_n748));
  OAI21_X1  g323(.A(new_n748), .B1(G162), .B2(new_n747), .ZN(new_n749));
  XOR2_X1   g324(.A(new_n749), .B(KEYINPUT29), .Z(new_n750));
  INV_X1    g325(.A(G2090), .ZN(new_n751));
  OAI21_X1  g326(.A(new_n746), .B1(new_n750), .B2(new_n751), .ZN(new_n752));
  XOR2_X1   g327(.A(new_n752), .B(KEYINPUT100), .Z(new_n753));
  NAND2_X1  g328(.A1(new_n611), .A2(G16), .ZN(new_n754));
  OAI21_X1  g329(.A(new_n754), .B1(G4), .B2(G16), .ZN(new_n755));
  INV_X1    g330(.A(G1348), .ZN(new_n756));
  NAND2_X1  g331(.A1(new_n755), .A2(new_n756), .ZN(new_n757));
  NAND2_X1  g332(.A1(new_n750), .A2(new_n751), .ZN(new_n758));
  NOR2_X1   g333(.A1(new_n706), .A2(G19), .ZN(new_n759));
  AOI21_X1  g334(.A(new_n759), .B1(new_n550), .B2(new_n706), .ZN(new_n760));
  XNOR2_X1  g335(.A(KEYINPUT94), .B(G1341), .ZN(new_n761));
  XNOR2_X1  g336(.A(new_n760), .B(new_n761), .ZN(new_n762));
  NAND2_X1  g337(.A1(new_n747), .A2(G26), .ZN(new_n763));
  XNOR2_X1  g338(.A(new_n763), .B(KEYINPUT28), .ZN(new_n764));
  NAND2_X1  g339(.A1(new_n471), .A2(G140), .ZN(new_n765));
  NAND2_X1  g340(.A1(new_n481), .A2(G128), .ZN(new_n766));
  INV_X1    g341(.A(G104), .ZN(new_n767));
  AND3_X1   g342(.A1(new_n767), .A2(new_n475), .A3(KEYINPUT95), .ZN(new_n768));
  AOI21_X1  g343(.A(KEYINPUT95), .B1(new_n767), .B2(new_n475), .ZN(new_n769));
  OAI221_X1 g344(.A(G2104), .B1(G116), .B2(new_n475), .C1(new_n768), .C2(new_n769), .ZN(new_n770));
  NAND3_X1  g345(.A1(new_n765), .A2(new_n766), .A3(new_n770), .ZN(new_n771));
  INV_X1    g346(.A(new_n771), .ZN(new_n772));
  OAI21_X1  g347(.A(new_n764), .B1(new_n772), .B2(new_n747), .ZN(new_n773));
  XNOR2_X1  g348(.A(new_n773), .B(G2067), .ZN(new_n774));
  NOR2_X1   g349(.A1(new_n762), .A2(new_n774), .ZN(new_n775));
  NAND3_X1  g350(.A1(new_n757), .A2(new_n758), .A3(new_n775), .ZN(new_n776));
  NOR2_X1   g351(.A1(new_n755), .A2(new_n756), .ZN(new_n777));
  NOR2_X1   g352(.A1(new_n776), .A2(new_n777), .ZN(new_n778));
  AND2_X1   g353(.A1(new_n747), .A2(G33), .ZN(new_n779));
  NAND3_X1  g354(.A1(new_n475), .A2(G103), .A3(G2104), .ZN(new_n780));
  XOR2_X1   g355(.A(new_n780), .B(KEYINPUT25), .Z(new_n781));
  AOI22_X1  g356(.A1(new_n473), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n782));
  INV_X1    g357(.A(new_n471), .ZN(new_n783));
  INV_X1    g358(.A(G139), .ZN(new_n784));
  OAI221_X1 g359(.A(new_n781), .B1(new_n475), .B2(new_n782), .C1(new_n783), .C2(new_n784), .ZN(new_n785));
  AOI21_X1  g360(.A(new_n779), .B1(new_n785), .B2(G29), .ZN(new_n786));
  INV_X1    g361(.A(G34), .ZN(new_n787));
  OR2_X1    g362(.A1(new_n787), .A2(KEYINPUT24), .ZN(new_n788));
  AOI21_X1  g363(.A(G29), .B1(new_n787), .B2(KEYINPUT24), .ZN(new_n789));
  AOI22_X1  g364(.A1(G160), .A2(G29), .B1(new_n788), .B2(new_n789), .ZN(new_n790));
  AOI22_X1  g365(.A1(new_n442), .A2(new_n786), .B1(new_n790), .B2(G2084), .ZN(new_n791));
  OR2_X1    g366(.A1(new_n786), .A2(new_n442), .ZN(new_n792));
  NAND2_X1  g367(.A1(new_n471), .A2(G141), .ZN(new_n793));
  NAND2_X1  g368(.A1(new_n481), .A2(G129), .ZN(new_n794));
  NAND3_X1  g369(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n795));
  INV_X1    g370(.A(KEYINPUT26), .ZN(new_n796));
  OR2_X1    g371(.A1(new_n795), .A2(new_n796), .ZN(new_n797));
  NAND2_X1  g372(.A1(new_n795), .A2(new_n796), .ZN(new_n798));
  AOI22_X1  g373(.A1(G105), .A2(new_n477), .B1(new_n797), .B2(new_n798), .ZN(new_n799));
  NAND3_X1  g374(.A1(new_n793), .A2(new_n794), .A3(new_n799), .ZN(new_n800));
  MUX2_X1   g375(.A(G32), .B(new_n800), .S(G29), .Z(new_n801));
  XOR2_X1   g376(.A(KEYINPUT27), .B(G1996), .Z(new_n802));
  OAI211_X1 g377(.A(new_n791), .B(new_n792), .C1(new_n801), .C2(new_n802), .ZN(new_n803));
  XNOR2_X1  g378(.A(new_n803), .B(KEYINPUT96), .ZN(new_n804));
  NOR2_X1   g379(.A1(G16), .A2(G21), .ZN(new_n805));
  AOI21_X1  g380(.A(new_n805), .B1(G168), .B2(G16), .ZN(new_n806));
  INV_X1    g381(.A(G1966), .ZN(new_n807));
  XNOR2_X1  g382(.A(new_n806), .B(new_n807), .ZN(new_n808));
  NAND2_X1  g383(.A1(new_n703), .A2(G5), .ZN(new_n809));
  OAI21_X1  g384(.A(new_n809), .B1(G171), .B2(new_n703), .ZN(new_n810));
  INV_X1    g385(.A(G1961), .ZN(new_n811));
  XNOR2_X1  g386(.A(new_n810), .B(new_n811), .ZN(new_n812));
  NAND2_X1  g387(.A1(new_n801), .A2(new_n802), .ZN(new_n813));
  NAND2_X1  g388(.A1(new_n812), .A2(new_n813), .ZN(new_n814));
  NAND2_X1  g389(.A1(new_n632), .A2(G29), .ZN(new_n815));
  INV_X1    g390(.A(KEYINPUT97), .ZN(new_n816));
  NAND2_X1  g391(.A1(new_n815), .A2(new_n816), .ZN(new_n817));
  XOR2_X1   g392(.A(KEYINPUT31), .B(G11), .Z(new_n818));
  INV_X1    g393(.A(KEYINPUT30), .ZN(new_n819));
  OAI21_X1  g394(.A(new_n747), .B1(new_n819), .B2(G28), .ZN(new_n820));
  INV_X1    g395(.A(KEYINPUT98), .ZN(new_n821));
  OR2_X1    g396(.A1(new_n820), .A2(new_n821), .ZN(new_n822));
  AOI22_X1  g397(.A1(new_n820), .A2(new_n821), .B1(new_n819), .B2(G28), .ZN(new_n823));
  AOI21_X1  g398(.A(new_n818), .B1(new_n822), .B2(new_n823), .ZN(new_n824));
  NAND2_X1  g399(.A1(new_n817), .A2(new_n824), .ZN(new_n825));
  OAI22_X1  g400(.A1(new_n815), .A2(new_n816), .B1(new_n790), .B2(G2084), .ZN(new_n826));
  NOR3_X1   g401(.A1(new_n814), .A2(new_n825), .A3(new_n826), .ZN(new_n827));
  NAND2_X1  g402(.A1(new_n747), .A2(G27), .ZN(new_n828));
  OAI21_X1  g403(.A(new_n828), .B1(G164), .B2(new_n747), .ZN(new_n829));
  XNOR2_X1  g404(.A(new_n829), .B(new_n443), .ZN(new_n830));
  NAND4_X1  g405(.A1(new_n804), .A2(new_n808), .A3(new_n827), .A4(new_n830), .ZN(new_n831));
  OAI211_X1 g406(.A(new_n753), .B(new_n778), .C1(new_n831), .C2(KEYINPUT99), .ZN(new_n832));
  AND2_X1   g407(.A1(new_n831), .A2(KEYINPUT99), .ZN(new_n833));
  OR3_X1    g408(.A1(new_n832), .A2(new_n833), .A3(KEYINPUT101), .ZN(new_n834));
  OAI21_X1  g409(.A(KEYINPUT101), .B1(new_n832), .B2(new_n833), .ZN(new_n835));
  AOI22_X1  g410(.A1(new_n740), .A2(new_n742), .B1(new_n834), .B2(new_n835), .ZN(G311));
  NAND2_X1  g411(.A1(new_n740), .A2(new_n742), .ZN(new_n837));
  NAND2_X1  g412(.A1(new_n834), .A2(new_n835), .ZN(new_n838));
  NAND2_X1  g413(.A1(new_n837), .A2(new_n838), .ZN(G150));
  NAND2_X1  g414(.A1(G80), .A2(G543), .ZN(new_n840));
  INV_X1    g415(.A(G67), .ZN(new_n841));
  OAI21_X1  g416(.A(new_n840), .B1(new_n572), .B2(new_n841), .ZN(new_n842));
  NAND2_X1  g417(.A1(new_n842), .A2(G651), .ZN(new_n843));
  INV_X1    g418(.A(KEYINPUT102), .ZN(new_n844));
  NAND2_X1  g419(.A1(new_n843), .A2(new_n844), .ZN(new_n845));
  NAND3_X1  g420(.A1(new_n842), .A2(KEYINPUT102), .A3(G651), .ZN(new_n846));
  NAND2_X1  g421(.A1(new_n525), .A2(G55), .ZN(new_n847));
  INV_X1    g422(.A(G93), .ZN(new_n848));
  OAI21_X1  g423(.A(new_n847), .B1(new_n512), .B2(new_n848), .ZN(new_n849));
  INV_X1    g424(.A(new_n849), .ZN(new_n850));
  NAND3_X1  g425(.A1(new_n845), .A2(new_n846), .A3(new_n850), .ZN(new_n851));
  NAND2_X1  g426(.A1(new_n851), .A2(new_n550), .ZN(new_n852));
  INV_X1    g427(.A(KEYINPUT103), .ZN(new_n853));
  NAND2_X1  g428(.A1(new_n852), .A2(new_n853), .ZN(new_n854));
  NAND3_X1  g429(.A1(new_n851), .A2(KEYINPUT103), .A3(new_n550), .ZN(new_n855));
  NAND2_X1  g430(.A1(new_n854), .A2(new_n855), .ZN(new_n856));
  INV_X1    g431(.A(KEYINPUT104), .ZN(new_n857));
  OAI21_X1  g432(.A(new_n857), .B1(new_n851), .B2(new_n550), .ZN(new_n858));
  INV_X1    g433(.A(new_n550), .ZN(new_n859));
  AOI21_X1  g434(.A(new_n849), .B1(new_n843), .B2(new_n844), .ZN(new_n860));
  NAND4_X1  g435(.A1(new_n859), .A2(new_n860), .A3(KEYINPUT104), .A4(new_n846), .ZN(new_n861));
  NAND2_X1  g436(.A1(new_n858), .A2(new_n861), .ZN(new_n862));
  NAND2_X1  g437(.A1(new_n856), .A2(new_n862), .ZN(new_n863));
  INV_X1    g438(.A(KEYINPUT38), .ZN(new_n864));
  NAND3_X1  g439(.A1(new_n611), .A2(new_n864), .A3(G559), .ZN(new_n865));
  OAI21_X1  g440(.A(KEYINPUT38), .B1(new_n610), .B2(new_n617), .ZN(new_n866));
  NAND2_X1  g441(.A1(new_n865), .A2(new_n866), .ZN(new_n867));
  XNOR2_X1  g442(.A(new_n863), .B(new_n867), .ZN(new_n868));
  NAND2_X1  g443(.A1(new_n868), .A2(KEYINPUT39), .ZN(new_n869));
  INV_X1    g444(.A(G860), .ZN(new_n870));
  NAND2_X1  g445(.A1(new_n869), .A2(new_n870), .ZN(new_n871));
  OR3_X1    g446(.A1(new_n868), .A2(KEYINPUT105), .A3(KEYINPUT39), .ZN(new_n872));
  OAI21_X1  g447(.A(KEYINPUT105), .B1(new_n868), .B2(KEYINPUT39), .ZN(new_n873));
  AOI21_X1  g448(.A(new_n871), .B1(new_n872), .B2(new_n873), .ZN(new_n874));
  INV_X1    g449(.A(KEYINPUT107), .ZN(new_n875));
  NAND2_X1  g450(.A1(new_n851), .A2(G860), .ZN(new_n876));
  XOR2_X1   g451(.A(KEYINPUT106), .B(KEYINPUT37), .Z(new_n877));
  XNOR2_X1  g452(.A(new_n876), .B(new_n877), .ZN(new_n878));
  INV_X1    g453(.A(new_n878), .ZN(new_n879));
  OR3_X1    g454(.A1(new_n874), .A2(new_n875), .A3(new_n879), .ZN(new_n880));
  OAI21_X1  g455(.A(new_n875), .B1(new_n874), .B2(new_n879), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n880), .A2(new_n881), .ZN(G145));
  INV_X1    g457(.A(G37), .ZN(new_n883));
  INV_X1    g458(.A(KEYINPUT108), .ZN(new_n884));
  AND3_X1   g459(.A1(new_n494), .A2(new_n884), .A3(new_n496), .ZN(new_n885));
  AOI21_X1  g460(.A(new_n884), .B1(new_n494), .B2(new_n496), .ZN(new_n886));
  NOR2_X1   g461(.A1(new_n885), .A2(new_n886), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n493), .A2(new_n887), .ZN(new_n888));
  XNOR2_X1  g463(.A(new_n888), .B(new_n771), .ZN(new_n889));
  XNOR2_X1  g464(.A(new_n889), .B(new_n800), .ZN(new_n890));
  XNOR2_X1  g465(.A(new_n890), .B(new_n785), .ZN(new_n891));
  XNOR2_X1  g466(.A(new_n733), .B(KEYINPUT109), .ZN(new_n892));
  INV_X1    g467(.A(new_n625), .ZN(new_n893));
  NAND2_X1  g468(.A1(new_n892), .A2(new_n893), .ZN(new_n894));
  INV_X1    g469(.A(new_n894), .ZN(new_n895));
  NAND2_X1  g470(.A1(new_n471), .A2(G142), .ZN(new_n896));
  NAND2_X1  g471(.A1(new_n481), .A2(G130), .ZN(new_n897));
  OR2_X1    g472(.A1(G106), .A2(G2105), .ZN(new_n898));
  OAI211_X1 g473(.A(new_n898), .B(G2104), .C1(G118), .C2(new_n475), .ZN(new_n899));
  NAND3_X1  g474(.A1(new_n896), .A2(new_n897), .A3(new_n899), .ZN(new_n900));
  NOR2_X1   g475(.A1(new_n892), .A2(new_n893), .ZN(new_n901));
  NOR3_X1   g476(.A1(new_n895), .A2(new_n900), .A3(new_n901), .ZN(new_n902));
  INV_X1    g477(.A(new_n900), .ZN(new_n903));
  INV_X1    g478(.A(new_n892), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n904), .A2(new_n625), .ZN(new_n905));
  AOI21_X1  g480(.A(new_n903), .B1(new_n905), .B2(new_n894), .ZN(new_n906));
  OAI21_X1  g481(.A(new_n891), .B1(new_n902), .B2(new_n906), .ZN(new_n907));
  INV_X1    g482(.A(KEYINPUT110), .ZN(new_n908));
  OAI21_X1  g483(.A(new_n908), .B1(new_n902), .B2(new_n906), .ZN(new_n909));
  OAI21_X1  g484(.A(new_n900), .B1(new_n895), .B2(new_n901), .ZN(new_n910));
  NAND3_X1  g485(.A1(new_n905), .A2(new_n894), .A3(new_n903), .ZN(new_n911));
  NAND3_X1  g486(.A1(new_n910), .A2(KEYINPUT110), .A3(new_n911), .ZN(new_n912));
  INV_X1    g487(.A(new_n785), .ZN(new_n913));
  AND2_X1   g488(.A1(new_n890), .A2(new_n913), .ZN(new_n914));
  NOR2_X1   g489(.A1(new_n890), .A2(new_n913), .ZN(new_n915));
  OAI211_X1 g490(.A(new_n909), .B(new_n912), .C1(new_n914), .C2(new_n915), .ZN(new_n916));
  XNOR2_X1  g491(.A(new_n632), .B(G160), .ZN(new_n917));
  XNOR2_X1  g492(.A(new_n917), .B(new_n485), .ZN(new_n918));
  INV_X1    g493(.A(new_n918), .ZN(new_n919));
  NAND3_X1  g494(.A1(new_n907), .A2(new_n916), .A3(new_n919), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n909), .A2(new_n912), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n921), .A2(new_n891), .ZN(new_n922));
  AND2_X1   g497(.A1(new_n922), .A2(new_n916), .ZN(new_n923));
  OAI211_X1 g498(.A(new_n883), .B(new_n920), .C1(new_n923), .C2(new_n919), .ZN(new_n924));
  XNOR2_X1  g499(.A(new_n924), .B(KEYINPUT40), .ZN(G395));
  OR2_X1    g500(.A1(new_n698), .A2(G303), .ZN(new_n926));
  NAND2_X1  g501(.A1(new_n698), .A2(G303), .ZN(new_n927));
  NAND2_X1  g502(.A1(new_n926), .A2(new_n927), .ZN(new_n928));
  NAND2_X1  g503(.A1(G290), .A2(new_n713), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n598), .A2(G305), .ZN(new_n930));
  NAND2_X1  g505(.A1(new_n929), .A2(new_n930), .ZN(new_n931));
  NAND2_X1  g506(.A1(new_n928), .A2(new_n931), .ZN(new_n932));
  NAND4_X1  g507(.A1(new_n926), .A2(new_n929), .A3(new_n927), .A4(new_n930), .ZN(new_n933));
  AND3_X1   g508(.A1(new_n932), .A2(KEYINPUT112), .A3(new_n933), .ZN(new_n934));
  AOI21_X1  g509(.A(KEYINPUT112), .B1(new_n932), .B2(new_n933), .ZN(new_n935));
  OAI21_X1  g510(.A(KEYINPUT42), .B1(new_n934), .B2(new_n935), .ZN(new_n936));
  INV_X1    g511(.A(KEYINPUT42), .ZN(new_n937));
  NAND3_X1  g512(.A1(new_n932), .A2(new_n937), .A3(new_n933), .ZN(new_n938));
  XNOR2_X1  g513(.A(new_n938), .B(KEYINPUT113), .ZN(new_n939));
  NAND2_X1  g514(.A1(new_n619), .A2(KEYINPUT111), .ZN(new_n940));
  INV_X1    g515(.A(new_n940), .ZN(new_n941));
  NOR2_X1   g516(.A1(new_n619), .A2(KEYINPUT111), .ZN(new_n942));
  OR3_X1    g517(.A1(new_n941), .A2(new_n863), .A3(new_n942), .ZN(new_n943));
  OAI21_X1  g518(.A(new_n863), .B1(new_n941), .B2(new_n942), .ZN(new_n944));
  NAND2_X1  g519(.A1(new_n943), .A2(new_n944), .ZN(new_n945));
  NAND2_X1  g520(.A1(new_n610), .A2(G299), .ZN(new_n946));
  INV_X1    g521(.A(new_n946), .ZN(new_n947));
  NOR2_X1   g522(.A1(new_n610), .A2(G299), .ZN(new_n948));
  NOR2_X1   g523(.A1(new_n947), .A2(new_n948), .ZN(new_n949));
  NAND2_X1  g524(.A1(new_n949), .A2(KEYINPUT41), .ZN(new_n950));
  INV_X1    g525(.A(new_n948), .ZN(new_n951));
  NAND2_X1  g526(.A1(new_n951), .A2(new_n946), .ZN(new_n952));
  INV_X1    g527(.A(KEYINPUT41), .ZN(new_n953));
  NAND2_X1  g528(.A1(new_n952), .A2(new_n953), .ZN(new_n954));
  NAND2_X1  g529(.A1(new_n950), .A2(new_n954), .ZN(new_n955));
  NAND2_X1  g530(.A1(new_n945), .A2(new_n955), .ZN(new_n956));
  NAND3_X1  g531(.A1(new_n943), .A2(new_n952), .A3(new_n944), .ZN(new_n957));
  AND4_X1   g532(.A1(new_n936), .A2(new_n939), .A3(new_n956), .A4(new_n957), .ZN(new_n958));
  AOI22_X1  g533(.A1(new_n939), .A2(new_n936), .B1(new_n956), .B2(new_n957), .ZN(new_n959));
  OAI21_X1  g534(.A(G868), .B1(new_n958), .B2(new_n959), .ZN(new_n960));
  INV_X1    g535(.A(G868), .ZN(new_n961));
  NAND2_X1  g536(.A1(new_n851), .A2(new_n961), .ZN(new_n962));
  NAND2_X1  g537(.A1(new_n960), .A2(new_n962), .ZN(G295));
  NAND2_X1  g538(.A1(new_n960), .A2(new_n962), .ZN(G331));
  INV_X1    g539(.A(KEYINPUT44), .ZN(new_n965));
  INV_X1    g540(.A(KEYINPUT43), .ZN(new_n966));
  NOR2_X1   g541(.A1(new_n934), .A2(new_n935), .ZN(new_n967));
  NAND2_X1  g542(.A1(G168), .A2(G171), .ZN(new_n968));
  NAND3_X1  g543(.A1(new_n532), .A2(new_n535), .A3(G301), .ZN(new_n969));
  NAND2_X1  g544(.A1(new_n968), .A2(new_n969), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n863), .A2(new_n970), .ZN(new_n971));
  NAND4_X1  g546(.A1(new_n856), .A2(new_n862), .A3(new_n968), .A4(new_n969), .ZN(new_n972));
  NAND2_X1  g547(.A1(new_n971), .A2(new_n972), .ZN(new_n973));
  NAND2_X1  g548(.A1(new_n973), .A2(new_n949), .ZN(new_n974));
  NAND4_X1  g549(.A1(new_n971), .A2(new_n950), .A3(new_n954), .A4(new_n972), .ZN(new_n975));
  NAND2_X1  g550(.A1(new_n974), .A2(new_n975), .ZN(new_n976));
  NAND2_X1  g551(.A1(new_n967), .A2(new_n976), .ZN(new_n977));
  OAI211_X1 g552(.A(new_n974), .B(new_n975), .C1(new_n934), .C2(new_n935), .ZN(new_n978));
  AND4_X1   g553(.A1(new_n966), .A2(new_n977), .A3(new_n883), .A4(new_n978), .ZN(new_n979));
  AOI21_X1  g554(.A(G37), .B1(new_n967), .B2(new_n976), .ZN(new_n980));
  AOI21_X1  g555(.A(new_n966), .B1(new_n980), .B2(new_n978), .ZN(new_n981));
  OAI21_X1  g556(.A(new_n965), .B1(new_n979), .B2(new_n981), .ZN(new_n982));
  NAND3_X1  g557(.A1(new_n977), .A2(new_n883), .A3(new_n978), .ZN(new_n983));
  NAND2_X1  g558(.A1(new_n983), .A2(KEYINPUT43), .ZN(new_n984));
  NAND3_X1  g559(.A1(new_n980), .A2(new_n966), .A3(new_n978), .ZN(new_n985));
  NAND3_X1  g560(.A1(new_n984), .A2(KEYINPUT44), .A3(new_n985), .ZN(new_n986));
  NAND2_X1  g561(.A1(new_n982), .A2(new_n986), .ZN(G397));
  AOI21_X1  g562(.A(G1384), .B1(new_n493), .B2(new_n887), .ZN(new_n988));
  NAND4_X1  g563(.A1(new_n472), .A2(new_n476), .A3(G40), .A4(new_n478), .ZN(new_n989));
  NOR3_X1   g564(.A1(new_n988), .A2(KEYINPUT45), .A3(new_n989), .ZN(new_n990));
  INV_X1    g565(.A(new_n990), .ZN(new_n991));
  NOR3_X1   g566(.A1(G290), .A2(new_n991), .A3(G1986), .ZN(new_n992));
  XOR2_X1   g567(.A(new_n992), .B(KEYINPUT48), .Z(new_n993));
  XNOR2_X1  g568(.A(new_n771), .B(G2067), .ZN(new_n994));
  XNOR2_X1  g569(.A(new_n800), .B(G1996), .ZN(new_n995));
  OAI21_X1  g570(.A(new_n990), .B1(new_n994), .B2(new_n995), .ZN(new_n996));
  INV_X1    g571(.A(KEYINPUT114), .ZN(new_n997));
  OR2_X1    g572(.A1(new_n996), .A2(new_n997), .ZN(new_n998));
  NAND2_X1  g573(.A1(new_n996), .A2(new_n997), .ZN(new_n999));
  NAND2_X1  g574(.A1(new_n998), .A2(new_n999), .ZN(new_n1000));
  XNOR2_X1  g575(.A(new_n733), .B(new_n736), .ZN(new_n1001));
  XNOR2_X1  g576(.A(new_n1001), .B(KEYINPUT115), .ZN(new_n1002));
  AOI21_X1  g577(.A(new_n1000), .B1(new_n990), .B2(new_n1002), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n993), .A2(new_n1003), .ZN(new_n1004));
  INV_X1    g579(.A(KEYINPUT46), .ZN(new_n1005));
  OR3_X1    g580(.A1(new_n991), .A2(new_n1005), .A3(G1996), .ZN(new_n1006));
  OAI21_X1  g581(.A(new_n990), .B1(new_n800), .B2(new_n994), .ZN(new_n1007));
  OAI21_X1  g582(.A(new_n1005), .B1(new_n991), .B2(G1996), .ZN(new_n1008));
  NAND3_X1  g583(.A1(new_n1006), .A2(new_n1007), .A3(new_n1008), .ZN(new_n1009));
  XNOR2_X1  g584(.A(new_n1009), .B(KEYINPUT47), .ZN(new_n1010));
  NAND2_X1  g585(.A1(new_n1004), .A2(new_n1010), .ZN(new_n1011));
  NOR2_X1   g586(.A1(new_n733), .A2(new_n736), .ZN(new_n1012));
  NAND3_X1  g587(.A1(new_n998), .A2(new_n999), .A3(new_n1012), .ZN(new_n1013));
  INV_X1    g588(.A(G2067), .ZN(new_n1014));
  NAND2_X1  g589(.A1(new_n772), .A2(new_n1014), .ZN(new_n1015));
  AND3_X1   g590(.A1(new_n1013), .A2(KEYINPUT125), .A3(new_n1015), .ZN(new_n1016));
  AOI21_X1  g591(.A(KEYINPUT125), .B1(new_n1013), .B2(new_n1015), .ZN(new_n1017));
  NOR3_X1   g592(.A1(new_n1016), .A2(new_n1017), .A3(new_n991), .ZN(new_n1018));
  OR3_X1    g593(.A1(new_n1011), .A2(new_n1018), .A3(KEYINPUT126), .ZN(new_n1019));
  OAI21_X1  g594(.A(KEYINPUT126), .B1(new_n1011), .B2(new_n1018), .ZN(new_n1020));
  NAND2_X1  g595(.A1(new_n1019), .A2(new_n1020), .ZN(new_n1021));
  INV_X1    g596(.A(new_n989), .ZN(new_n1022));
  INV_X1    g597(.A(G1384), .ZN(new_n1023));
  NAND3_X1  g598(.A1(new_n888), .A2(new_n1022), .A3(new_n1023), .ZN(new_n1024));
  AND2_X1   g599(.A1(new_n1024), .A2(G8), .ZN(new_n1025));
  NOR2_X1   g600(.A1(G288), .A2(G1976), .ZN(new_n1026));
  XNOR2_X1  g601(.A(new_n1026), .B(KEYINPUT118), .ZN(new_n1027));
  INV_X1    g602(.A(KEYINPUT117), .ZN(new_n1028));
  INV_X1    g603(.A(KEYINPUT49), .ZN(new_n1029));
  NOR2_X1   g604(.A1(G305), .A2(G1981), .ZN(new_n1030));
  NOR2_X1   g605(.A1(new_n512), .A2(new_n579), .ZN(new_n1031));
  OAI21_X1  g606(.A(G1981), .B1(new_n1031), .B2(new_n586), .ZN(new_n1032));
  INV_X1    g607(.A(KEYINPUT116), .ZN(new_n1033));
  NAND2_X1  g608(.A1(new_n1032), .A2(new_n1033), .ZN(new_n1034));
  OAI211_X1 g609(.A(KEYINPUT116), .B(G1981), .C1(new_n1031), .C2(new_n586), .ZN(new_n1035));
  NAND2_X1  g610(.A1(new_n1034), .A2(new_n1035), .ZN(new_n1036));
  OAI211_X1 g611(.A(new_n1028), .B(new_n1029), .C1(new_n1030), .C2(new_n1036), .ZN(new_n1037));
  INV_X1    g612(.A(G1981), .ZN(new_n1038));
  AOI21_X1  g613(.A(new_n1036), .B1(new_n1038), .B2(new_n713), .ZN(new_n1039));
  OAI21_X1  g614(.A(KEYINPUT49), .B1(new_n1039), .B2(KEYINPUT117), .ZN(new_n1040));
  AOI21_X1  g615(.A(new_n1027), .B1(new_n1037), .B2(new_n1040), .ZN(new_n1041));
  OAI21_X1  g616(.A(new_n1025), .B1(new_n1041), .B2(new_n1030), .ZN(new_n1042));
  NAND3_X1  g617(.A1(new_n1037), .A2(new_n1040), .A3(new_n1025), .ZN(new_n1043));
  INV_X1    g618(.A(new_n489), .ZN(new_n1044));
  NAND2_X1  g619(.A1(new_n490), .A2(KEYINPUT4), .ZN(new_n1045));
  INV_X1    g620(.A(KEYINPUT65), .ZN(new_n1046));
  NAND2_X1  g621(.A1(new_n1045), .A2(new_n1046), .ZN(new_n1047));
  NAND3_X1  g622(.A1(new_n490), .A2(KEYINPUT65), .A3(KEYINPUT4), .ZN(new_n1048));
  AOI21_X1  g623(.A(new_n1044), .B1(new_n1047), .B2(new_n1048), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n497), .A2(KEYINPUT108), .ZN(new_n1050));
  NAND3_X1  g625(.A1(new_n494), .A2(new_n884), .A3(new_n496), .ZN(new_n1051));
  NAND2_X1  g626(.A1(new_n1050), .A2(new_n1051), .ZN(new_n1052));
  OAI211_X1 g627(.A(KEYINPUT45), .B(new_n1023), .C1(new_n1049), .C2(new_n1052), .ZN(new_n1053));
  AOI21_X1  g628(.A(G1384), .B1(new_n493), .B2(new_n498), .ZN(new_n1054));
  OAI211_X1 g629(.A(new_n1053), .B(new_n1022), .C1(KEYINPUT45), .C2(new_n1054), .ZN(new_n1055));
  INV_X1    g630(.A(G1971), .ZN(new_n1056));
  NAND2_X1  g631(.A1(new_n1055), .A2(new_n1056), .ZN(new_n1057));
  INV_X1    g632(.A(KEYINPUT50), .ZN(new_n1058));
  OAI211_X1 g633(.A(new_n1058), .B(new_n1023), .C1(new_n1049), .C2(new_n1052), .ZN(new_n1059));
  OAI211_X1 g634(.A(new_n1059), .B(new_n1022), .C1(new_n1058), .C2(new_n1054), .ZN(new_n1060));
  OAI21_X1  g635(.A(new_n1057), .B1(G2090), .B2(new_n1060), .ZN(new_n1061));
  AND2_X1   g636(.A1(new_n1061), .A2(G8), .ZN(new_n1062));
  NAND2_X1  g637(.A1(G303), .A2(G8), .ZN(new_n1063));
  XOR2_X1   g638(.A(new_n1063), .B(KEYINPUT55), .Z(new_n1064));
  INV_X1    g639(.A(KEYINPUT52), .ZN(new_n1065));
  NAND3_X1  g640(.A1(new_n695), .A2(G1976), .A3(new_n697), .ZN(new_n1066));
  AOI21_X1  g641(.A(new_n1065), .B1(new_n1025), .B2(new_n1066), .ZN(new_n1067));
  AND2_X1   g642(.A1(new_n1025), .A2(new_n1066), .ZN(new_n1068));
  INV_X1    g643(.A(G1976), .ZN(new_n1069));
  AOI21_X1  g644(.A(KEYINPUT52), .B1(G288), .B2(new_n1069), .ZN(new_n1070));
  AOI21_X1  g645(.A(new_n1067), .B1(new_n1068), .B2(new_n1070), .ZN(new_n1071));
  NAND4_X1  g646(.A1(new_n1043), .A2(new_n1062), .A3(new_n1064), .A4(new_n1071), .ZN(new_n1072));
  AND2_X1   g647(.A1(new_n1042), .A2(new_n1072), .ZN(new_n1073));
  NAND3_X1  g648(.A1(new_n1061), .A2(G8), .A3(new_n1064), .ZN(new_n1074));
  NAND3_X1  g649(.A1(new_n1043), .A2(new_n1074), .A3(new_n1071), .ZN(new_n1075));
  NOR2_X1   g650(.A1(KEYINPUT50), .A2(G1384), .ZN(new_n1076));
  OAI21_X1  g651(.A(new_n1076), .B1(new_n1049), .B2(new_n497), .ZN(new_n1077));
  OAI211_X1 g652(.A(new_n1077), .B(new_n1022), .C1(new_n988), .C2(new_n1058), .ZN(new_n1078));
  NAND2_X1  g653(.A1(new_n1078), .A2(KEYINPUT119), .ZN(new_n1079));
  NAND2_X1  g654(.A1(new_n1079), .A2(new_n751), .ZN(new_n1080));
  NOR2_X1   g655(.A1(new_n1078), .A2(KEYINPUT119), .ZN(new_n1081));
  OAI21_X1  g656(.A(new_n1057), .B1(new_n1080), .B2(new_n1081), .ZN(new_n1082));
  AOI21_X1  g657(.A(new_n1064), .B1(new_n1082), .B2(G8), .ZN(new_n1083));
  NOR2_X1   g658(.A1(new_n1075), .A2(new_n1083), .ZN(new_n1084));
  INV_X1    g659(.A(KEYINPUT120), .ZN(new_n1085));
  NOR2_X1   g660(.A1(new_n989), .A2(G2084), .ZN(new_n1086));
  OAI211_X1 g661(.A(new_n1059), .B(new_n1086), .C1(new_n1058), .C2(new_n1054), .ZN(new_n1087));
  OAI211_X1 g662(.A(KEYINPUT45), .B(new_n1023), .C1(new_n1049), .C2(new_n497), .ZN(new_n1088));
  OAI211_X1 g663(.A(new_n1088), .B(new_n1022), .C1(new_n988), .C2(KEYINPUT45), .ZN(new_n1089));
  AOI22_X1  g664(.A1(new_n1085), .A2(new_n1087), .B1(new_n1089), .B2(new_n807), .ZN(new_n1090));
  OR2_X1    g665(.A1(new_n1087), .A2(new_n1085), .ZN(new_n1091));
  NAND2_X1  g666(.A1(new_n1090), .A2(new_n1091), .ZN(new_n1092));
  AND3_X1   g667(.A1(new_n1092), .A2(G8), .A3(G168), .ZN(new_n1093));
  AOI21_X1  g668(.A(KEYINPUT63), .B1(new_n1084), .B2(new_n1093), .ZN(new_n1094));
  OAI211_X1 g669(.A(new_n1093), .B(KEYINPUT63), .C1(new_n1064), .C2(new_n1062), .ZN(new_n1095));
  NOR2_X1   g670(.A1(new_n1095), .A2(new_n1075), .ZN(new_n1096));
  OAI21_X1  g671(.A(new_n1073), .B1(new_n1094), .B2(new_n1096), .ZN(new_n1097));
  INV_X1    g672(.A(KEYINPUT53), .ZN(new_n1098));
  OAI21_X1  g673(.A(new_n1098), .B1(new_n1055), .B2(G2078), .ZN(new_n1099));
  NOR2_X1   g674(.A1(new_n1098), .A2(G2078), .ZN(new_n1100));
  AND2_X1   g675(.A1(new_n1053), .A2(new_n1100), .ZN(new_n1101));
  OAI21_X1  g676(.A(new_n1023), .B1(new_n1049), .B2(new_n1052), .ZN(new_n1102));
  INV_X1    g677(.A(KEYINPUT45), .ZN(new_n1103));
  AOI21_X1  g678(.A(new_n989), .B1(new_n1102), .B2(new_n1103), .ZN(new_n1104));
  AOI21_X1  g679(.A(G171), .B1(new_n1101), .B2(new_n1104), .ZN(new_n1105));
  NAND2_X1  g680(.A1(new_n1060), .A2(new_n811), .ZN(new_n1106));
  NAND3_X1  g681(.A1(new_n1099), .A2(new_n1105), .A3(new_n1106), .ZN(new_n1107));
  INV_X1    g682(.A(KEYINPUT122), .ZN(new_n1108));
  NAND2_X1  g683(.A1(new_n1107), .A2(new_n1108), .ZN(new_n1109));
  INV_X1    g684(.A(new_n1099), .ZN(new_n1110));
  NAND3_X1  g685(.A1(new_n1104), .A2(new_n1088), .A3(new_n1100), .ZN(new_n1111));
  NAND2_X1  g686(.A1(new_n1106), .A2(new_n1111), .ZN(new_n1112));
  OAI21_X1  g687(.A(G171), .B1(new_n1110), .B2(new_n1112), .ZN(new_n1113));
  NAND4_X1  g688(.A1(new_n1099), .A2(new_n1105), .A3(KEYINPUT122), .A4(new_n1106), .ZN(new_n1114));
  NAND3_X1  g689(.A1(new_n1109), .A2(new_n1113), .A3(new_n1114), .ZN(new_n1115));
  INV_X1    g690(.A(KEYINPUT54), .ZN(new_n1116));
  NAND2_X1  g691(.A1(new_n1115), .A2(new_n1116), .ZN(new_n1117));
  NAND2_X1  g692(.A1(new_n1117), .A2(KEYINPUT123), .ZN(new_n1118));
  NAND3_X1  g693(.A1(new_n1090), .A2(G168), .A3(new_n1091), .ZN(new_n1119));
  NAND2_X1  g694(.A1(new_n1119), .A2(G8), .ZN(new_n1120));
  NAND2_X1  g695(.A1(new_n1120), .A2(KEYINPUT51), .ZN(new_n1121));
  AOI21_X1  g696(.A(G168), .B1(new_n1090), .B2(new_n1091), .ZN(new_n1122));
  INV_X1    g697(.A(KEYINPUT51), .ZN(new_n1123));
  OAI211_X1 g698(.A(G8), .B(new_n1119), .C1(new_n1122), .C2(new_n1123), .ZN(new_n1124));
  NAND2_X1  g699(.A1(new_n1101), .A2(new_n1104), .ZN(new_n1125));
  NAND3_X1  g700(.A1(new_n1099), .A2(new_n1106), .A3(new_n1125), .ZN(new_n1126));
  INV_X1    g701(.A(KEYINPUT124), .ZN(new_n1127));
  NAND2_X1  g702(.A1(new_n1126), .A2(new_n1127), .ZN(new_n1128));
  NAND4_X1  g703(.A1(new_n1099), .A2(new_n1125), .A3(KEYINPUT124), .A4(new_n1106), .ZN(new_n1129));
  NAND3_X1  g704(.A1(new_n1128), .A2(G171), .A3(new_n1129), .ZN(new_n1130));
  NAND4_X1  g705(.A1(new_n1099), .A2(G301), .A3(new_n1111), .A4(new_n1106), .ZN(new_n1131));
  AND2_X1   g706(.A1(new_n1131), .A2(KEYINPUT54), .ZN(new_n1132));
  AOI22_X1  g707(.A1(new_n1121), .A2(new_n1124), .B1(new_n1130), .B2(new_n1132), .ZN(new_n1133));
  INV_X1    g708(.A(G1956), .ZN(new_n1134));
  NAND2_X1  g709(.A1(new_n1078), .A2(new_n1134), .ZN(new_n1135));
  OAI21_X1  g710(.A(new_n1023), .B1(new_n1049), .B2(new_n497), .ZN(new_n1136));
  NAND2_X1  g711(.A1(new_n1136), .A2(new_n1103), .ZN(new_n1137));
  XNOR2_X1  g712(.A(KEYINPUT56), .B(G2072), .ZN(new_n1138));
  NAND4_X1  g713(.A1(new_n1137), .A2(new_n1053), .A3(new_n1022), .A4(new_n1138), .ZN(new_n1139));
  NAND2_X1  g714(.A1(G299), .A2(KEYINPUT57), .ZN(new_n1140));
  INV_X1    g715(.A(KEYINPUT57), .ZN(new_n1141));
  NAND3_X1  g716(.A1(new_n560), .A2(new_n1141), .A3(new_n568), .ZN(new_n1142));
  NAND2_X1  g717(.A1(new_n1140), .A2(new_n1142), .ZN(new_n1143));
  INV_X1    g718(.A(new_n1143), .ZN(new_n1144));
  AND3_X1   g719(.A1(new_n1135), .A2(new_n1139), .A3(new_n1144), .ZN(new_n1145));
  INV_X1    g720(.A(new_n1145), .ZN(new_n1146));
  OAI21_X1  g721(.A(KEYINPUT121), .B1(new_n1024), .B2(G2067), .ZN(new_n1147));
  INV_X1    g722(.A(KEYINPUT121), .ZN(new_n1148));
  NAND4_X1  g723(.A1(new_n988), .A2(new_n1148), .A3(new_n1014), .A4(new_n1022), .ZN(new_n1149));
  AND2_X1   g724(.A1(new_n1147), .A2(new_n1149), .ZN(new_n1150));
  NAND2_X1  g725(.A1(new_n1060), .A2(new_n756), .ZN(new_n1151));
  AOI21_X1  g726(.A(new_n610), .B1(new_n1150), .B2(new_n1151), .ZN(new_n1152));
  AOI21_X1  g727(.A(new_n1144), .B1(new_n1135), .B2(new_n1139), .ZN(new_n1153));
  OAI21_X1  g728(.A(new_n1146), .B1(new_n1152), .B2(new_n1153), .ZN(new_n1154));
  INV_X1    g729(.A(KEYINPUT61), .ZN(new_n1155));
  OAI21_X1  g730(.A(new_n1155), .B1(new_n1145), .B2(new_n1153), .ZN(new_n1156));
  AOI21_X1  g731(.A(KEYINPUT60), .B1(new_n1150), .B2(new_n1151), .ZN(new_n1157));
  NAND4_X1  g732(.A1(new_n1151), .A2(KEYINPUT60), .A3(new_n1147), .A4(new_n1149), .ZN(new_n1158));
  NAND2_X1  g733(.A1(new_n1158), .A2(new_n611), .ZN(new_n1159));
  OAI21_X1  g734(.A(new_n1156), .B1(new_n1157), .B2(new_n1159), .ZN(new_n1160));
  NOR2_X1   g735(.A1(new_n989), .A2(G1996), .ZN(new_n1161));
  OAI211_X1 g736(.A(new_n1053), .B(new_n1161), .C1(KEYINPUT45), .C2(new_n1054), .ZN(new_n1162));
  XOR2_X1   g737(.A(KEYINPUT58), .B(G1341), .Z(new_n1163));
  NAND2_X1  g738(.A1(new_n1024), .A2(new_n1163), .ZN(new_n1164));
  NAND2_X1  g739(.A1(new_n1162), .A2(new_n1164), .ZN(new_n1165));
  NAND2_X1  g740(.A1(new_n1165), .A2(new_n550), .ZN(new_n1166));
  NAND2_X1  g741(.A1(new_n1166), .A2(KEYINPUT59), .ZN(new_n1167));
  INV_X1    g742(.A(KEYINPUT59), .ZN(new_n1168));
  NAND3_X1  g743(.A1(new_n1165), .A2(new_n1168), .A3(new_n550), .ZN(new_n1169));
  NAND2_X1  g744(.A1(new_n1167), .A2(new_n1169), .ZN(new_n1170));
  NAND4_X1  g745(.A1(new_n1150), .A2(KEYINPUT60), .A3(new_n610), .A4(new_n1151), .ZN(new_n1171));
  AOI21_X1  g746(.A(new_n1143), .B1(new_n1078), .B2(new_n1134), .ZN(new_n1172));
  AOI21_X1  g747(.A(new_n1155), .B1(new_n1172), .B2(new_n1139), .ZN(new_n1173));
  AND4_X1   g748(.A1(new_n1137), .A2(new_n1053), .A3(new_n1022), .A4(new_n1138), .ZN(new_n1174));
  NAND2_X1  g749(.A1(new_n1102), .A2(KEYINPUT50), .ZN(new_n1175));
  AOI21_X1  g750(.A(new_n989), .B1(new_n499), .B2(new_n1076), .ZN(new_n1176));
  AOI21_X1  g751(.A(G1956), .B1(new_n1175), .B2(new_n1176), .ZN(new_n1177));
  OAI21_X1  g752(.A(new_n1143), .B1(new_n1174), .B2(new_n1177), .ZN(new_n1178));
  NAND2_X1  g753(.A1(new_n1173), .A2(new_n1178), .ZN(new_n1179));
  NAND3_X1  g754(.A1(new_n1170), .A2(new_n1171), .A3(new_n1179), .ZN(new_n1180));
  OAI21_X1  g755(.A(new_n1154), .B1(new_n1160), .B2(new_n1180), .ZN(new_n1181));
  INV_X1    g756(.A(KEYINPUT123), .ZN(new_n1182));
  NAND3_X1  g757(.A1(new_n1115), .A2(new_n1182), .A3(new_n1116), .ZN(new_n1183));
  NAND4_X1  g758(.A1(new_n1118), .A2(new_n1133), .A3(new_n1181), .A4(new_n1183), .ZN(new_n1184));
  AOI21_X1  g759(.A(new_n1123), .B1(new_n1092), .B2(G286), .ZN(new_n1185));
  NOR2_X1   g760(.A1(new_n1185), .A2(new_n1120), .ZN(new_n1186));
  AOI21_X1  g761(.A(new_n1123), .B1(new_n1119), .B2(G8), .ZN(new_n1187));
  OAI21_X1  g762(.A(KEYINPUT62), .B1(new_n1186), .B2(new_n1187), .ZN(new_n1188));
  INV_X1    g763(.A(new_n1113), .ZN(new_n1189));
  INV_X1    g764(.A(KEYINPUT62), .ZN(new_n1190));
  NAND3_X1  g765(.A1(new_n1121), .A2(new_n1124), .A3(new_n1190), .ZN(new_n1191));
  NAND3_X1  g766(.A1(new_n1188), .A2(new_n1189), .A3(new_n1191), .ZN(new_n1192));
  NAND2_X1  g767(.A1(new_n1184), .A2(new_n1192), .ZN(new_n1193));
  AOI21_X1  g768(.A(new_n1097), .B1(new_n1193), .B2(new_n1084), .ZN(new_n1194));
  XNOR2_X1  g769(.A(new_n598), .B(G1986), .ZN(new_n1195));
  OAI21_X1  g770(.A(new_n1003), .B1(new_n991), .B2(new_n1195), .ZN(new_n1196));
  OAI21_X1  g771(.A(new_n1021), .B1(new_n1194), .B2(new_n1196), .ZN(G329));
  assign    G231 = 1'b0;
  NOR2_X1   g772(.A1(G227), .A2(new_n462), .ZN(new_n1199));
  INV_X1    g773(.A(new_n1199), .ZN(new_n1200));
  OR3_X1    g774(.A1(G401), .A2(KEYINPUT127), .A3(new_n1200), .ZN(new_n1201));
  OAI21_X1  g775(.A(KEYINPUT127), .B1(G401), .B2(new_n1200), .ZN(new_n1202));
  AND3_X1   g776(.A1(new_n692), .A2(new_n1201), .A3(new_n1202), .ZN(new_n1203));
  NAND2_X1  g777(.A1(new_n1203), .A2(new_n924), .ZN(new_n1204));
  AOI21_X1  g778(.A(new_n1204), .B1(new_n984), .B2(new_n985), .ZN(G308));
  OAI211_X1 g779(.A(new_n924), .B(new_n1203), .C1(new_n979), .C2(new_n981), .ZN(G225));
endmodule


