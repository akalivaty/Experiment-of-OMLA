//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 0 0 1 1 1 0 1 1 0 0 1 1 1 0 0 0 1 1 1 1 1 0 0 0 1 0 0 1 0 0 1 0 1 0 1 0 1 0 0 1 0 0 0 0 0 0 1 1 0 1 1 0 0 1 0 1 0 1 0 0 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:32:16 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n437, new_n444, new_n445, new_n446, new_n451, new_n452,
    new_n454, new_n457, new_n458, new_n459, new_n460, new_n463, new_n464,
    new_n465, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n524, new_n525, new_n526,
    new_n527, new_n528, new_n529, new_n530, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n550, new_n552,
    new_n553, new_n555, new_n556, new_n557, new_n558, new_n559, new_n560,
    new_n561, new_n562, new_n563, new_n564, new_n565, new_n566, new_n567,
    new_n568, new_n569, new_n570, new_n573, new_n574, new_n575, new_n577,
    new_n578, new_n579, new_n580, new_n581, new_n582, new_n583, new_n585,
    new_n586, new_n587, new_n588, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n602,
    new_n605, new_n607, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1149, new_n1150, new_n1151, new_n1152, new_n1153, new_n1154,
    new_n1155, new_n1156;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(new_n436));
  INV_X1    g011(.A(KEYINPUT64), .ZN(new_n437));
  XNOR2_X1  g012(.A(new_n436), .B(new_n437), .ZN(G220));
  INV_X1    g013(.A(G96), .ZN(G221));
  INV_X1    g014(.A(G69), .ZN(G235));
  INV_X1    g015(.A(G120), .ZN(G236));
  XOR2_X1   g016(.A(KEYINPUT65), .B(G57), .Z(G237));
  INV_X1    g017(.A(G108), .ZN(G238));
  INV_X1    g018(.A(G2072), .ZN(new_n444));
  INV_X1    g019(.A(G2078), .ZN(new_n445));
  NOR2_X1   g020(.A1(new_n444), .A2(new_n445), .ZN(new_n446));
  NAND3_X1  g021(.A1(new_n446), .A2(G2084), .A3(G2090), .ZN(G158));
  NAND3_X1  g022(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g023(.A(G452), .Z(G391));
  AND2_X1   g024(.A1(G94), .A2(G452), .ZN(G173));
  XNOR2_X1  g025(.A(KEYINPUT66), .B(KEYINPUT1), .ZN(new_n451));
  NAND2_X1  g026(.A1(G7), .A2(G661), .ZN(new_n452));
  XNOR2_X1  g027(.A(new_n451), .B(new_n452), .ZN(G223));
  INV_X1    g028(.A(new_n452), .ZN(new_n454));
  NAND2_X1  g029(.A1(new_n454), .A2(G567), .ZN(G234));
  NAND2_X1  g030(.A1(new_n454), .A2(G2106), .ZN(G217));
  NOR4_X1   g031(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n457));
  XOR2_X1   g032(.A(new_n457), .B(KEYINPUT2), .Z(new_n458));
  NOR4_X1   g033(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n459));
  XNOR2_X1  g034(.A(new_n459), .B(KEYINPUT67), .ZN(new_n460));
  NOR2_X1   g035(.A1(new_n458), .A2(new_n460), .ZN(G325));
  INV_X1    g036(.A(G325), .ZN(G261));
  NAND2_X1  g037(.A1(new_n458), .A2(G2106), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n460), .A2(G567), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  INV_X1    g040(.A(new_n465), .ZN(G319));
  INV_X1    g041(.A(G125), .ZN(new_n467));
  INV_X1    g042(.A(KEYINPUT3), .ZN(new_n468));
  INV_X1    g043(.A(G2104), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  NAND2_X1  g045(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n471));
  AOI21_X1  g046(.A(new_n467), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  AND2_X1   g047(.A1(G113), .A2(G2104), .ZN(new_n473));
  OAI21_X1  g048(.A(G2105), .B1(new_n472), .B2(new_n473), .ZN(new_n474));
  INV_X1    g049(.A(G101), .ZN(new_n475));
  NOR3_X1   g050(.A1(new_n475), .A2(new_n469), .A3(G2105), .ZN(new_n476));
  AOI21_X1  g051(.A(G2105), .B1(new_n470), .B2(new_n471), .ZN(new_n477));
  AOI21_X1  g052(.A(new_n476), .B1(new_n477), .B2(G137), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n474), .A2(new_n478), .ZN(new_n479));
  INV_X1    g054(.A(new_n479), .ZN(G160));
  AND2_X1   g055(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n481));
  NOR2_X1   g056(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n482));
  NOR2_X1   g057(.A1(new_n481), .A2(new_n482), .ZN(new_n483));
  INV_X1    g058(.A(G2105), .ZN(new_n484));
  NOR2_X1   g059(.A1(new_n483), .A2(new_n484), .ZN(new_n485));
  NAND2_X1  g060(.A1(new_n485), .A2(G124), .ZN(new_n486));
  MUX2_X1   g061(.A(G100), .B(G112), .S(G2105), .Z(new_n487));
  NAND2_X1  g062(.A1(new_n487), .A2(G2104), .ZN(new_n488));
  NAND2_X1  g063(.A1(new_n486), .A2(new_n488), .ZN(new_n489));
  AOI21_X1  g064(.A(new_n489), .B1(G136), .B2(new_n477), .ZN(G162));
  INV_X1    g065(.A(G126), .ZN(new_n491));
  AOI21_X1  g066(.A(new_n491), .B1(new_n470), .B2(new_n471), .ZN(new_n492));
  AND2_X1   g067(.A1(G114), .A2(G2104), .ZN(new_n493));
  OAI21_X1  g068(.A(G2105), .B1(new_n492), .B2(new_n493), .ZN(new_n494));
  NAND2_X1  g069(.A1(KEYINPUT4), .A2(G138), .ZN(new_n495));
  AOI21_X1  g070(.A(new_n495), .B1(new_n470), .B2(new_n471), .ZN(new_n496));
  NAND2_X1  g071(.A1(G102), .A2(G2104), .ZN(new_n497));
  INV_X1    g072(.A(new_n497), .ZN(new_n498));
  OAI21_X1  g073(.A(new_n484), .B1(new_n496), .B2(new_n498), .ZN(new_n499));
  OAI211_X1 g074(.A(G138), .B(new_n484), .C1(new_n481), .C2(new_n482), .ZN(new_n500));
  INV_X1    g075(.A(KEYINPUT4), .ZN(new_n501));
  NAND2_X1  g076(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  NAND3_X1  g077(.A1(new_n494), .A2(new_n499), .A3(new_n502), .ZN(new_n503));
  INV_X1    g078(.A(new_n503), .ZN(G164));
  INV_X1    g079(.A(G543), .ZN(new_n505));
  INV_X1    g080(.A(KEYINPUT6), .ZN(new_n506));
  INV_X1    g081(.A(KEYINPUT68), .ZN(new_n507));
  INV_X1    g082(.A(G651), .ZN(new_n508));
  OAI21_X1  g083(.A(new_n506), .B1(new_n507), .B2(new_n508), .ZN(new_n509));
  NAND3_X1  g084(.A1(KEYINPUT68), .A2(KEYINPUT6), .A3(G651), .ZN(new_n510));
  AOI21_X1  g085(.A(new_n505), .B1(new_n509), .B2(new_n510), .ZN(new_n511));
  NAND2_X1  g086(.A1(new_n511), .A2(G50), .ZN(new_n512));
  INV_X1    g087(.A(G88), .ZN(new_n513));
  NAND2_X1  g088(.A1(new_n509), .A2(new_n510), .ZN(new_n514));
  OR2_X1    g089(.A1(KEYINPUT5), .A2(G543), .ZN(new_n515));
  NAND2_X1  g090(.A1(KEYINPUT5), .A2(G543), .ZN(new_n516));
  NAND2_X1  g091(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  NAND2_X1  g092(.A1(new_n514), .A2(new_n517), .ZN(new_n518));
  OAI21_X1  g093(.A(new_n512), .B1(new_n513), .B2(new_n518), .ZN(new_n519));
  AOI22_X1  g094(.A1(new_n517), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n520));
  NOR2_X1   g095(.A1(new_n520), .A2(new_n508), .ZN(new_n521));
  OR2_X1    g096(.A1(new_n519), .A2(new_n521), .ZN(G303));
  INV_X1    g097(.A(G303), .ZN(G166));
  AND2_X1   g098(.A1(new_n514), .A2(new_n517), .ZN(new_n524));
  AND2_X1   g099(.A1(new_n524), .A2(G89), .ZN(new_n525));
  NAND2_X1  g100(.A1(new_n511), .A2(G51), .ZN(new_n526));
  NAND3_X1  g101(.A1(new_n517), .A2(G63), .A3(G651), .ZN(new_n527));
  NAND3_X1  g102(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n528));
  XNOR2_X1  g103(.A(new_n528), .B(KEYINPUT7), .ZN(new_n529));
  NAND3_X1  g104(.A1(new_n526), .A2(new_n527), .A3(new_n529), .ZN(new_n530));
  NOR2_X1   g105(.A1(new_n525), .A2(new_n530), .ZN(G168));
  NAND2_X1  g106(.A1(new_n511), .A2(G52), .ZN(new_n532));
  INV_X1    g107(.A(G90), .ZN(new_n533));
  OAI21_X1  g108(.A(new_n532), .B1(new_n533), .B2(new_n518), .ZN(new_n534));
  AOI22_X1  g109(.A1(new_n517), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n535));
  NOR2_X1   g110(.A1(new_n535), .A2(new_n508), .ZN(new_n536));
  OR2_X1    g111(.A1(new_n534), .A2(new_n536), .ZN(G301));
  INV_X1    g112(.A(G301), .ZN(G171));
  AOI22_X1  g113(.A1(new_n517), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n539));
  OR2_X1    g114(.A1(new_n539), .A2(new_n508), .ZN(new_n540));
  NAND2_X1  g115(.A1(new_n524), .A2(G81), .ZN(new_n541));
  NAND2_X1  g116(.A1(new_n511), .A2(G43), .ZN(new_n542));
  AOI21_X1  g117(.A(KEYINPUT69), .B1(new_n541), .B2(new_n542), .ZN(new_n543));
  INV_X1    g118(.A(G81), .ZN(new_n544));
  OAI211_X1 g119(.A(new_n542), .B(KEYINPUT69), .C1(new_n544), .C2(new_n518), .ZN(new_n545));
  INV_X1    g120(.A(new_n545), .ZN(new_n546));
  OAI21_X1  g121(.A(new_n540), .B1(new_n543), .B2(new_n546), .ZN(new_n547));
  INV_X1    g122(.A(G860), .ZN(new_n548));
  OR2_X1    g123(.A1(new_n547), .A2(new_n548), .ZN(G153));
  AND3_X1   g124(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n550));
  NAND2_X1  g125(.A1(new_n550), .A2(G36), .ZN(G176));
  NAND2_X1  g126(.A1(G1), .A2(G3), .ZN(new_n552));
  XNOR2_X1  g127(.A(new_n552), .B(KEYINPUT8), .ZN(new_n553));
  NAND2_X1  g128(.A1(new_n550), .A2(new_n553), .ZN(G188));
  NAND3_X1  g129(.A1(new_n511), .A2(KEYINPUT70), .A3(G53), .ZN(new_n555));
  INV_X1    g130(.A(KEYINPUT9), .ZN(new_n556));
  NAND2_X1  g131(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  NAND4_X1  g132(.A1(new_n511), .A2(KEYINPUT70), .A3(KEYINPUT9), .A4(G53), .ZN(new_n558));
  INV_X1    g133(.A(KEYINPUT71), .ZN(new_n559));
  INV_X1    g134(.A(G65), .ZN(new_n560));
  AOI21_X1  g135(.A(new_n560), .B1(new_n515), .B2(new_n516), .ZN(new_n561));
  NAND2_X1  g136(.A1(G78), .A2(G543), .ZN(new_n562));
  INV_X1    g137(.A(new_n562), .ZN(new_n563));
  OAI211_X1 g138(.A(new_n559), .B(G651), .C1(new_n561), .C2(new_n563), .ZN(new_n564));
  NAND3_X1  g139(.A1(new_n557), .A2(new_n558), .A3(new_n564), .ZN(new_n565));
  OAI21_X1  g140(.A(G651), .B1(new_n561), .B2(new_n563), .ZN(new_n566));
  INV_X1    g141(.A(new_n566), .ZN(new_n567));
  INV_X1    g142(.A(G91), .ZN(new_n568));
  OAI22_X1  g143(.A1(new_n567), .A2(new_n559), .B1(new_n568), .B2(new_n518), .ZN(new_n569));
  NOR2_X1   g144(.A1(new_n565), .A2(new_n569), .ZN(new_n570));
  INV_X1    g145(.A(new_n570), .ZN(G299));
  INV_X1    g146(.A(G168), .ZN(G286));
  NAND2_X1  g147(.A1(new_n524), .A2(G87), .ZN(new_n573));
  NAND2_X1  g148(.A1(new_n511), .A2(G49), .ZN(new_n574));
  OAI21_X1  g149(.A(G651), .B1(new_n517), .B2(G74), .ZN(new_n575));
  NAND3_X1  g150(.A1(new_n573), .A2(new_n574), .A3(new_n575), .ZN(G288));
  NAND2_X1  g151(.A1(new_n511), .A2(G48), .ZN(new_n577));
  INV_X1    g152(.A(G61), .ZN(new_n578));
  AOI21_X1  g153(.A(new_n578), .B1(new_n515), .B2(new_n516), .ZN(new_n579));
  AND2_X1   g154(.A1(G73), .A2(G543), .ZN(new_n580));
  OAI21_X1  g155(.A(G651), .B1(new_n579), .B2(new_n580), .ZN(new_n581));
  NAND3_X1  g156(.A1(new_n514), .A2(G86), .A3(new_n517), .ZN(new_n582));
  AND3_X1   g157(.A1(new_n577), .A2(new_n581), .A3(new_n582), .ZN(new_n583));
  INV_X1    g158(.A(new_n583), .ZN(G305));
  NAND2_X1  g159(.A1(new_n524), .A2(G85), .ZN(new_n585));
  AOI22_X1  g160(.A1(new_n517), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n586));
  INV_X1    g161(.A(new_n511), .ZN(new_n587));
  XOR2_X1   g162(.A(KEYINPUT72), .B(G47), .Z(new_n588));
  OAI221_X1 g163(.A(new_n585), .B1(new_n508), .B2(new_n586), .C1(new_n587), .C2(new_n588), .ZN(G290));
  INV_X1    g164(.A(G868), .ZN(new_n590));
  NOR2_X1   g165(.A1(G301), .A2(new_n590), .ZN(new_n591));
  AND3_X1   g166(.A1(new_n514), .A2(G92), .A3(new_n517), .ZN(new_n592));
  XNOR2_X1  g167(.A(new_n592), .B(KEYINPUT10), .ZN(new_n593));
  AND2_X1   g168(.A1(new_n511), .A2(KEYINPUT73), .ZN(new_n594));
  NOR2_X1   g169(.A1(new_n511), .A2(KEYINPUT73), .ZN(new_n595));
  OAI21_X1  g170(.A(G54), .B1(new_n594), .B2(new_n595), .ZN(new_n596));
  AOI22_X1  g171(.A1(new_n517), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n597));
  OR2_X1    g172(.A1(new_n597), .A2(new_n508), .ZN(new_n598));
  AND3_X1   g173(.A1(new_n593), .A2(new_n596), .A3(new_n598), .ZN(new_n599));
  AOI21_X1  g174(.A(new_n591), .B1(new_n599), .B2(new_n590), .ZN(G284));
  AOI21_X1  g175(.A(new_n591), .B1(new_n599), .B2(new_n590), .ZN(G321));
  NOR2_X1   g176(.A1(G286), .A2(new_n590), .ZN(new_n602));
  AOI21_X1  g177(.A(new_n602), .B1(new_n590), .B2(new_n570), .ZN(G297));
  AOI21_X1  g178(.A(new_n602), .B1(new_n590), .B2(new_n570), .ZN(G280));
  XNOR2_X1  g179(.A(KEYINPUT74), .B(G559), .ZN(new_n605));
  OAI21_X1  g180(.A(new_n599), .B1(G860), .B2(new_n605), .ZN(G148));
  NAND2_X1  g181(.A1(new_n599), .A2(new_n605), .ZN(new_n607));
  MUX2_X1   g182(.A(new_n547), .B(new_n607), .S(G868), .Z(G323));
  XNOR2_X1  g183(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g184(.A1(new_n477), .A2(G2104), .ZN(new_n610));
  XNOR2_X1  g185(.A(new_n610), .B(KEYINPUT12), .ZN(new_n611));
  INV_X1    g186(.A(G2100), .ZN(new_n612));
  AOI22_X1  g187(.A1(new_n611), .A2(KEYINPUT13), .B1(KEYINPUT75), .B2(new_n612), .ZN(new_n613));
  OAI21_X1  g188(.A(new_n613), .B1(KEYINPUT13), .B2(new_n611), .ZN(new_n614));
  OR3_X1    g189(.A1(new_n614), .A2(KEYINPUT75), .A3(new_n612), .ZN(new_n615));
  OAI21_X1  g190(.A(new_n614), .B1(KEYINPUT75), .B2(new_n612), .ZN(new_n616));
  NAND2_X1  g191(.A1(new_n485), .A2(G123), .ZN(new_n617));
  NAND2_X1  g192(.A1(new_n477), .A2(G135), .ZN(new_n618));
  AND2_X1   g193(.A1(G111), .A2(G2105), .ZN(new_n619));
  AOI21_X1  g194(.A(new_n619), .B1(G99), .B2(new_n484), .ZN(new_n620));
  OAI211_X1 g195(.A(new_n617), .B(new_n618), .C1(new_n469), .C2(new_n620), .ZN(new_n621));
  XOR2_X1   g196(.A(new_n621), .B(G2096), .Z(new_n622));
  NAND3_X1  g197(.A1(new_n615), .A2(new_n616), .A3(new_n622), .ZN(G156));
  XNOR2_X1  g198(.A(KEYINPUT15), .B(G2435), .ZN(new_n624));
  INV_X1    g199(.A(G2438), .ZN(new_n625));
  XNOR2_X1  g200(.A(new_n624), .B(new_n625), .ZN(new_n626));
  XNOR2_X1  g201(.A(new_n626), .B(G2427), .ZN(new_n627));
  INV_X1    g202(.A(G2430), .ZN(new_n628));
  OR2_X1    g203(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  NAND2_X1  g204(.A1(new_n627), .A2(new_n628), .ZN(new_n630));
  NAND3_X1  g205(.A1(new_n629), .A2(KEYINPUT14), .A3(new_n630), .ZN(new_n631));
  XNOR2_X1  g206(.A(G2451), .B(G2454), .ZN(new_n632));
  XNOR2_X1  g207(.A(G2443), .B(G2446), .ZN(new_n633));
  XNOR2_X1  g208(.A(new_n632), .B(new_n633), .ZN(new_n634));
  XOR2_X1   g209(.A(KEYINPUT76), .B(KEYINPUT16), .Z(new_n635));
  XNOR2_X1  g210(.A(new_n634), .B(new_n635), .ZN(new_n636));
  XNOR2_X1  g211(.A(new_n631), .B(new_n636), .ZN(new_n637));
  XNOR2_X1  g212(.A(G1341), .B(G1348), .ZN(new_n638));
  INV_X1    g213(.A(new_n638), .ZN(new_n639));
  NAND2_X1  g214(.A1(new_n637), .A2(new_n639), .ZN(new_n640));
  NAND2_X1  g215(.A1(new_n640), .A2(G14), .ZN(new_n641));
  OAI21_X1  g216(.A(KEYINPUT77), .B1(new_n637), .B2(new_n639), .ZN(new_n642));
  INV_X1    g217(.A(new_n637), .ZN(new_n643));
  INV_X1    g218(.A(KEYINPUT77), .ZN(new_n644));
  NAND3_X1  g219(.A1(new_n643), .A2(new_n644), .A3(new_n638), .ZN(new_n645));
  AOI21_X1  g220(.A(new_n641), .B1(new_n642), .B2(new_n645), .ZN(G401));
  XNOR2_X1  g221(.A(G2084), .B(G2090), .ZN(new_n647));
  INV_X1    g222(.A(KEYINPUT78), .ZN(new_n648));
  XNOR2_X1  g223(.A(new_n647), .B(new_n648), .ZN(new_n649));
  NOR2_X1   g224(.A1(G2072), .A2(G2078), .ZN(new_n650));
  NOR2_X1   g225(.A1(new_n446), .A2(new_n650), .ZN(new_n651));
  INV_X1    g226(.A(new_n651), .ZN(new_n652));
  XNOR2_X1  g227(.A(G2067), .B(G2678), .ZN(new_n653));
  NAND3_X1  g228(.A1(new_n649), .A2(new_n652), .A3(new_n653), .ZN(new_n654));
  XOR2_X1   g229(.A(new_n654), .B(KEYINPUT18), .Z(new_n655));
  INV_X1    g230(.A(new_n649), .ZN(new_n656));
  NAND2_X1  g231(.A1(new_n652), .A2(KEYINPUT17), .ZN(new_n657));
  NAND2_X1  g232(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  NAND2_X1  g233(.A1(new_n658), .A2(new_n653), .ZN(new_n659));
  OAI21_X1  g234(.A(KEYINPUT17), .B1(new_n649), .B2(new_n653), .ZN(new_n660));
  NAND2_X1  g235(.A1(new_n660), .A2(new_n651), .ZN(new_n661));
  OAI211_X1 g236(.A(new_n659), .B(new_n661), .C1(new_n656), .C2(new_n657), .ZN(new_n662));
  NAND2_X1  g237(.A1(new_n655), .A2(new_n662), .ZN(new_n663));
  XNOR2_X1  g238(.A(new_n663), .B(G2096), .ZN(new_n664));
  XNOR2_X1  g239(.A(KEYINPUT79), .B(G2100), .ZN(new_n665));
  XNOR2_X1  g240(.A(new_n664), .B(new_n665), .ZN(G227));
  XNOR2_X1  g241(.A(G1961), .B(G1966), .ZN(new_n667));
  XNOR2_X1  g242(.A(new_n667), .B(KEYINPUT80), .ZN(new_n668));
  XNOR2_X1  g243(.A(G1956), .B(G2474), .ZN(new_n669));
  INV_X1    g244(.A(new_n669), .ZN(new_n670));
  NAND2_X1  g245(.A1(new_n668), .A2(new_n670), .ZN(new_n671));
  XNOR2_X1  g246(.A(G1971), .B(G1976), .ZN(new_n672));
  XNOR2_X1  g247(.A(new_n672), .B(KEYINPUT19), .ZN(new_n673));
  NOR2_X1   g248(.A1(new_n671), .A2(new_n673), .ZN(new_n674));
  XOR2_X1   g249(.A(new_n674), .B(KEYINPUT20), .Z(new_n675));
  NOR2_X1   g250(.A1(new_n668), .A2(new_n670), .ZN(new_n676));
  INV_X1    g251(.A(new_n676), .ZN(new_n677));
  NAND3_X1  g252(.A1(new_n677), .A2(new_n673), .A3(new_n671), .ZN(new_n678));
  OAI211_X1 g253(.A(new_n675), .B(new_n678), .C1(new_n673), .C2(new_n677), .ZN(new_n679));
  XOR2_X1   g254(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n680));
  XNOR2_X1  g255(.A(new_n679), .B(new_n680), .ZN(new_n681));
  XNOR2_X1  g256(.A(G1991), .B(G1996), .ZN(new_n682));
  XNOR2_X1  g257(.A(G1981), .B(G1986), .ZN(new_n683));
  XNOR2_X1  g258(.A(new_n682), .B(new_n683), .ZN(new_n684));
  XNOR2_X1  g259(.A(new_n681), .B(new_n684), .ZN(new_n685));
  INV_X1    g260(.A(new_n685), .ZN(G229));
  NOR2_X1   g261(.A1(G6), .A2(G16), .ZN(new_n687));
  AOI21_X1  g262(.A(new_n687), .B1(new_n583), .B2(G16), .ZN(new_n688));
  XNOR2_X1  g263(.A(new_n688), .B(KEYINPUT83), .ZN(new_n689));
  XNOR2_X1  g264(.A(KEYINPUT32), .B(G1981), .ZN(new_n690));
  XNOR2_X1  g265(.A(new_n689), .B(new_n690), .ZN(new_n691));
  NOR2_X1   g266(.A1(G16), .A2(G23), .ZN(new_n692));
  XOR2_X1   g267(.A(new_n692), .B(KEYINPUT84), .Z(new_n693));
  INV_X1    g268(.A(G16), .ZN(new_n694));
  OAI21_X1  g269(.A(new_n693), .B1(G288), .B2(new_n694), .ZN(new_n695));
  XNOR2_X1  g270(.A(KEYINPUT33), .B(G1976), .ZN(new_n696));
  XNOR2_X1  g271(.A(new_n696), .B(KEYINPUT85), .ZN(new_n697));
  XNOR2_X1  g272(.A(new_n695), .B(new_n697), .ZN(new_n698));
  NOR2_X1   g273(.A1(G16), .A2(G22), .ZN(new_n699));
  AOI21_X1  g274(.A(new_n699), .B1(G166), .B2(G16), .ZN(new_n700));
  XNOR2_X1  g275(.A(new_n700), .B(G1971), .ZN(new_n701));
  NOR3_X1   g276(.A1(new_n691), .A2(new_n698), .A3(new_n701), .ZN(new_n702));
  INV_X1    g277(.A(KEYINPUT34), .ZN(new_n703));
  AND2_X1   g278(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  NOR2_X1   g279(.A1(new_n702), .A2(new_n703), .ZN(new_n705));
  MUX2_X1   g280(.A(G95), .B(G107), .S(G2105), .Z(new_n706));
  AOI22_X1  g281(.A1(new_n485), .A2(G119), .B1(G2104), .B2(new_n706), .ZN(new_n707));
  INV_X1    g282(.A(G131), .ZN(new_n708));
  INV_X1    g283(.A(new_n477), .ZN(new_n709));
  OAI21_X1  g284(.A(new_n707), .B1(new_n708), .B2(new_n709), .ZN(new_n710));
  INV_X1    g285(.A(G29), .ZN(new_n711));
  OR2_X1    g286(.A1(new_n711), .A2(KEYINPUT81), .ZN(new_n712));
  NAND2_X1  g287(.A1(new_n711), .A2(KEYINPUT81), .ZN(new_n713));
  NAND2_X1  g288(.A1(new_n712), .A2(new_n713), .ZN(new_n714));
  MUX2_X1   g289(.A(G25), .B(new_n710), .S(new_n714), .Z(new_n715));
  XNOR2_X1  g290(.A(KEYINPUT35), .B(G1991), .ZN(new_n716));
  XNOR2_X1  g291(.A(new_n715), .B(new_n716), .ZN(new_n717));
  MUX2_X1   g292(.A(G24), .B(G290), .S(G16), .Z(new_n718));
  XOR2_X1   g293(.A(KEYINPUT82), .B(G1986), .Z(new_n719));
  XOR2_X1   g294(.A(new_n718), .B(new_n719), .Z(new_n720));
  NOR4_X1   g295(.A1(new_n704), .A2(new_n705), .A3(new_n717), .A4(new_n720), .ZN(new_n721));
  XNOR2_X1  g296(.A(new_n721), .B(KEYINPUT36), .ZN(new_n722));
  XOR2_X1   g297(.A(KEYINPUT93), .B(KEYINPUT26), .Z(new_n723));
  NAND3_X1  g298(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n724));
  XNOR2_X1  g299(.A(new_n723), .B(new_n724), .ZN(new_n725));
  NAND2_X1  g300(.A1(new_n485), .A2(G129), .ZN(new_n726));
  NAND3_X1  g301(.A1(new_n484), .A2(G105), .A3(G2104), .ZN(new_n727));
  XOR2_X1   g302(.A(new_n727), .B(KEYINPUT92), .Z(new_n728));
  NAND2_X1  g303(.A1(new_n477), .A2(G141), .ZN(new_n729));
  NAND4_X1  g304(.A1(new_n725), .A2(new_n726), .A3(new_n728), .A4(new_n729), .ZN(new_n730));
  MUX2_X1   g305(.A(G32), .B(new_n730), .S(G29), .Z(new_n731));
  XOR2_X1   g306(.A(new_n731), .B(KEYINPUT94), .Z(new_n732));
  XNOR2_X1  g307(.A(KEYINPUT27), .B(G1996), .ZN(new_n733));
  INV_X1    g308(.A(new_n733), .ZN(new_n734));
  NAND2_X1  g309(.A1(new_n732), .A2(new_n734), .ZN(new_n735));
  INV_X1    g310(.A(G34), .ZN(new_n736));
  AOI21_X1  g311(.A(new_n714), .B1(KEYINPUT24), .B2(new_n736), .ZN(new_n737));
  NAND2_X1  g312(.A1(new_n737), .A2(KEYINPUT91), .ZN(new_n738));
  OAI21_X1  g313(.A(new_n738), .B1(KEYINPUT24), .B2(new_n736), .ZN(new_n739));
  NOR2_X1   g314(.A1(new_n737), .A2(KEYINPUT91), .ZN(new_n740));
  OAI22_X1  g315(.A1(new_n739), .A2(new_n740), .B1(new_n711), .B2(new_n479), .ZN(new_n741));
  INV_X1    g316(.A(G2084), .ZN(new_n742));
  AND2_X1   g317(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  XNOR2_X1  g318(.A(KEYINPUT31), .B(G11), .ZN(new_n744));
  OR2_X1    g319(.A1(KEYINPUT30), .A2(G28), .ZN(new_n745));
  NAND2_X1  g320(.A1(KEYINPUT30), .A2(G28), .ZN(new_n746));
  AND2_X1   g321(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  INV_X1    g322(.A(new_n714), .ZN(new_n748));
  OAI221_X1 g323(.A(new_n744), .B1(G29), .B2(new_n747), .C1(new_n621), .C2(new_n748), .ZN(new_n749));
  NOR2_X1   g324(.A1(new_n743), .A2(new_n749), .ZN(new_n750));
  OAI211_X1 g325(.A(new_n735), .B(new_n750), .C1(new_n742), .C2(new_n741), .ZN(new_n751));
  NAND2_X1  g326(.A1(new_n694), .A2(G5), .ZN(new_n752));
  OAI21_X1  g327(.A(new_n752), .B1(G171), .B2(new_n694), .ZN(new_n753));
  INV_X1    g328(.A(G1961), .ZN(new_n754));
  XNOR2_X1  g329(.A(new_n753), .B(new_n754), .ZN(new_n755));
  INV_X1    g330(.A(G1966), .ZN(new_n756));
  NOR2_X1   g331(.A1(G168), .A2(new_n694), .ZN(new_n757));
  AOI21_X1  g332(.A(new_n757), .B1(new_n694), .B2(G21), .ZN(new_n758));
  NAND2_X1  g333(.A1(new_n748), .A2(G26), .ZN(new_n759));
  XNOR2_X1  g334(.A(new_n759), .B(KEYINPUT28), .ZN(new_n760));
  NAND2_X1  g335(.A1(new_n485), .A2(G128), .ZN(new_n761));
  INV_X1    g336(.A(KEYINPUT87), .ZN(new_n762));
  XNOR2_X1  g337(.A(new_n761), .B(new_n762), .ZN(new_n763));
  MUX2_X1   g338(.A(G104), .B(G116), .S(G2105), .Z(new_n764));
  AOI22_X1  g339(.A1(G140), .A2(new_n477), .B1(new_n764), .B2(G2104), .ZN(new_n765));
  NAND2_X1  g340(.A1(new_n763), .A2(new_n765), .ZN(new_n766));
  INV_X1    g341(.A(new_n766), .ZN(new_n767));
  OAI21_X1  g342(.A(new_n760), .B1(new_n767), .B2(new_n711), .ZN(new_n768));
  OAI221_X1 g343(.A(new_n755), .B1(new_n756), .B2(new_n758), .C1(G2067), .C2(new_n768), .ZN(new_n769));
  NOR2_X1   g344(.A1(new_n732), .A2(new_n734), .ZN(new_n770));
  AOI22_X1  g345(.A1(new_n768), .A2(G2067), .B1(new_n758), .B2(new_n756), .ZN(new_n771));
  NOR2_X1   g346(.A1(new_n714), .A2(G27), .ZN(new_n772));
  AOI21_X1  g347(.A(new_n772), .B1(G164), .B2(new_n714), .ZN(new_n773));
  XNOR2_X1  g348(.A(new_n773), .B(new_n445), .ZN(new_n774));
  NAND2_X1  g349(.A1(new_n771), .A2(new_n774), .ZN(new_n775));
  NOR4_X1   g350(.A1(new_n751), .A2(new_n769), .A3(new_n770), .A4(new_n775), .ZN(new_n776));
  MUX2_X1   g351(.A(G19), .B(new_n547), .S(G16), .Z(new_n777));
  XNOR2_X1  g352(.A(KEYINPUT86), .B(G1341), .ZN(new_n778));
  XOR2_X1   g353(.A(new_n777), .B(new_n778), .Z(new_n779));
  NAND2_X1  g354(.A1(new_n694), .A2(G20), .ZN(new_n780));
  XNOR2_X1  g355(.A(new_n780), .B(KEYINPUT23), .ZN(new_n781));
  OAI21_X1  g356(.A(new_n781), .B1(new_n570), .B2(new_n694), .ZN(new_n782));
  INV_X1    g357(.A(G1956), .ZN(new_n783));
  NOR2_X1   g358(.A1(new_n782), .A2(new_n783), .ZN(new_n784));
  AND2_X1   g359(.A1(new_n782), .A2(new_n783), .ZN(new_n785));
  OAI211_X1 g360(.A(new_n776), .B(new_n779), .C1(new_n784), .C2(new_n785), .ZN(new_n786));
  NAND3_X1  g361(.A1(new_n484), .A2(G103), .A3(G2104), .ZN(new_n787));
  XNOR2_X1  g362(.A(new_n787), .B(KEYINPUT88), .ZN(new_n788));
  INV_X1    g363(.A(KEYINPUT25), .ZN(new_n789));
  AOI22_X1  g364(.A1(new_n788), .A2(new_n789), .B1(G139), .B2(new_n477), .ZN(new_n790));
  OAI21_X1  g365(.A(new_n790), .B1(new_n789), .B2(new_n788), .ZN(new_n791));
  XNOR2_X1  g366(.A(new_n791), .B(KEYINPUT89), .ZN(new_n792));
  NAND2_X1  g367(.A1(G115), .A2(G2104), .ZN(new_n793));
  INV_X1    g368(.A(G127), .ZN(new_n794));
  OAI21_X1  g369(.A(new_n793), .B1(new_n483), .B2(new_n794), .ZN(new_n795));
  INV_X1    g370(.A(KEYINPUT90), .ZN(new_n796));
  AOI21_X1  g371(.A(new_n484), .B1(new_n795), .B2(new_n796), .ZN(new_n797));
  OAI21_X1  g372(.A(new_n797), .B1(new_n796), .B2(new_n795), .ZN(new_n798));
  NAND2_X1  g373(.A1(new_n792), .A2(new_n798), .ZN(new_n799));
  MUX2_X1   g374(.A(G33), .B(new_n799), .S(G29), .Z(new_n800));
  XNOR2_X1  g375(.A(new_n800), .B(new_n444), .ZN(new_n801));
  NOR2_X1   g376(.A1(new_n714), .A2(G35), .ZN(new_n802));
  AOI21_X1  g377(.A(new_n802), .B1(G162), .B2(new_n714), .ZN(new_n803));
  XNOR2_X1  g378(.A(new_n803), .B(KEYINPUT29), .ZN(new_n804));
  INV_X1    g379(.A(G2090), .ZN(new_n805));
  XNOR2_X1  g380(.A(new_n804), .B(new_n805), .ZN(new_n806));
  NAND2_X1  g381(.A1(new_n599), .A2(G16), .ZN(new_n807));
  OAI21_X1  g382(.A(new_n807), .B1(G4), .B2(G16), .ZN(new_n808));
  INV_X1    g383(.A(G1348), .ZN(new_n809));
  OR2_X1    g384(.A1(new_n808), .A2(new_n809), .ZN(new_n810));
  NAND2_X1  g385(.A1(new_n808), .A2(new_n809), .ZN(new_n811));
  NAND4_X1  g386(.A1(new_n801), .A2(new_n806), .A3(new_n810), .A4(new_n811), .ZN(new_n812));
  NOR3_X1   g387(.A1(new_n722), .A2(new_n786), .A3(new_n812), .ZN(G311));
  INV_X1    g388(.A(G311), .ZN(G150));
  NAND2_X1  g389(.A1(new_n511), .A2(G55), .ZN(new_n815));
  XNOR2_X1  g390(.A(KEYINPUT95), .B(G93), .ZN(new_n816));
  OAI21_X1  g391(.A(new_n815), .B1(new_n518), .B2(new_n816), .ZN(new_n817));
  AOI22_X1  g392(.A1(new_n517), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n818));
  NOR2_X1   g393(.A1(new_n818), .A2(new_n508), .ZN(new_n819));
  NOR2_X1   g394(.A1(new_n817), .A2(new_n819), .ZN(new_n820));
  NOR2_X1   g395(.A1(new_n820), .A2(new_n548), .ZN(new_n821));
  XNOR2_X1  g396(.A(new_n821), .B(KEYINPUT37), .ZN(new_n822));
  INV_X1    g397(.A(new_n820), .ZN(new_n823));
  NAND2_X1  g398(.A1(new_n547), .A2(new_n823), .ZN(new_n824));
  OAI211_X1 g399(.A(new_n540), .B(new_n820), .C1(new_n543), .C2(new_n546), .ZN(new_n825));
  NAND2_X1  g400(.A1(new_n824), .A2(new_n825), .ZN(new_n826));
  XNOR2_X1  g401(.A(new_n826), .B(KEYINPUT38), .ZN(new_n827));
  NAND2_X1  g402(.A1(new_n599), .A2(G559), .ZN(new_n828));
  XNOR2_X1  g403(.A(new_n827), .B(new_n828), .ZN(new_n829));
  INV_X1    g404(.A(new_n829), .ZN(new_n830));
  OR2_X1    g405(.A1(new_n830), .A2(KEYINPUT39), .ZN(new_n831));
  INV_X1    g406(.A(KEYINPUT96), .ZN(new_n832));
  AND2_X1   g407(.A1(new_n831), .A2(new_n832), .ZN(new_n833));
  AOI21_X1  g408(.A(G860), .B1(new_n830), .B2(KEYINPUT39), .ZN(new_n834));
  OAI21_X1  g409(.A(new_n834), .B1(new_n831), .B2(new_n832), .ZN(new_n835));
  OAI21_X1  g410(.A(new_n822), .B1(new_n833), .B2(new_n835), .ZN(G145));
  NAND2_X1  g411(.A1(new_n799), .A2(KEYINPUT98), .ZN(new_n837));
  XNOR2_X1  g412(.A(new_n766), .B(new_n503), .ZN(new_n838));
  XNOR2_X1  g413(.A(new_n838), .B(new_n730), .ZN(new_n839));
  XNOR2_X1  g414(.A(new_n710), .B(new_n611), .ZN(new_n840));
  MUX2_X1   g415(.A(G106), .B(G118), .S(G2105), .Z(new_n841));
  AOI22_X1  g416(.A1(new_n485), .A2(G130), .B1(G2104), .B2(new_n841), .ZN(new_n842));
  INV_X1    g417(.A(G142), .ZN(new_n843));
  OAI21_X1  g418(.A(new_n842), .B1(new_n843), .B2(new_n709), .ZN(new_n844));
  XNOR2_X1  g419(.A(new_n840), .B(new_n844), .ZN(new_n845));
  INV_X1    g420(.A(new_n845), .ZN(new_n846));
  OR2_X1    g421(.A1(new_n799), .A2(KEYINPUT98), .ZN(new_n847));
  NAND3_X1  g422(.A1(new_n839), .A2(new_n846), .A3(new_n847), .ZN(new_n848));
  INV_X1    g423(.A(new_n848), .ZN(new_n849));
  AOI21_X1  g424(.A(new_n846), .B1(new_n839), .B2(new_n847), .ZN(new_n850));
  OAI21_X1  g425(.A(new_n837), .B1(new_n849), .B2(new_n850), .ZN(new_n851));
  INV_X1    g426(.A(new_n850), .ZN(new_n852));
  INV_X1    g427(.A(new_n837), .ZN(new_n853));
  NAND3_X1  g428(.A1(new_n852), .A2(new_n853), .A3(new_n848), .ZN(new_n854));
  NAND2_X1  g429(.A1(new_n851), .A2(new_n854), .ZN(new_n855));
  XNOR2_X1  g430(.A(G162), .B(new_n479), .ZN(new_n856));
  XOR2_X1   g431(.A(new_n621), .B(KEYINPUT97), .Z(new_n857));
  XNOR2_X1  g432(.A(new_n856), .B(new_n857), .ZN(new_n858));
  INV_X1    g433(.A(new_n858), .ZN(new_n859));
  NAND2_X1  g434(.A1(new_n855), .A2(new_n859), .ZN(new_n860));
  INV_X1    g435(.A(G37), .ZN(new_n861));
  NAND3_X1  g436(.A1(new_n851), .A2(new_n854), .A3(new_n858), .ZN(new_n862));
  NAND3_X1  g437(.A1(new_n860), .A2(new_n861), .A3(new_n862), .ZN(new_n863));
  XNOR2_X1  g438(.A(new_n863), .B(KEYINPUT40), .ZN(G395));
  XNOR2_X1  g439(.A(new_n826), .B(new_n607), .ZN(new_n865));
  NAND2_X1  g440(.A1(new_n599), .A2(G299), .ZN(new_n866));
  NAND2_X1  g441(.A1(new_n866), .A2(KEYINPUT99), .ZN(new_n867));
  NAND3_X1  g442(.A1(new_n593), .A2(new_n596), .A3(new_n598), .ZN(new_n868));
  OR3_X1    g443(.A1(new_n868), .A2(new_n570), .A3(KEYINPUT99), .ZN(new_n869));
  NAND2_X1  g444(.A1(new_n868), .A2(new_n570), .ZN(new_n870));
  NAND3_X1  g445(.A1(new_n867), .A2(new_n869), .A3(new_n870), .ZN(new_n871));
  NAND2_X1  g446(.A1(new_n865), .A2(new_n871), .ZN(new_n872));
  XNOR2_X1  g447(.A(new_n872), .B(KEYINPUT100), .ZN(new_n873));
  NAND2_X1  g448(.A1(new_n866), .A2(new_n870), .ZN(new_n874));
  INV_X1    g449(.A(KEYINPUT41), .ZN(new_n875));
  NAND2_X1  g450(.A1(new_n874), .A2(new_n875), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n876), .A2(KEYINPUT101), .ZN(new_n877));
  NAND4_X1  g452(.A1(new_n867), .A2(KEYINPUT41), .A3(new_n869), .A4(new_n870), .ZN(new_n878));
  INV_X1    g453(.A(KEYINPUT101), .ZN(new_n879));
  NAND3_X1  g454(.A1(new_n874), .A2(new_n879), .A3(new_n875), .ZN(new_n880));
  NAND3_X1  g455(.A1(new_n877), .A2(new_n878), .A3(new_n880), .ZN(new_n881));
  INV_X1    g456(.A(new_n881), .ZN(new_n882));
  OAI21_X1  g457(.A(new_n873), .B1(new_n882), .B2(new_n865), .ZN(new_n883));
  XNOR2_X1  g458(.A(G290), .B(G288), .ZN(new_n884));
  XNOR2_X1  g459(.A(G303), .B(G305), .ZN(new_n885));
  XOR2_X1   g460(.A(new_n884), .B(new_n885), .Z(new_n886));
  XNOR2_X1  g461(.A(KEYINPUT102), .B(KEYINPUT42), .ZN(new_n887));
  XOR2_X1   g462(.A(new_n886), .B(new_n887), .Z(new_n888));
  INV_X1    g463(.A(new_n888), .ZN(new_n889));
  OAI21_X1  g464(.A(KEYINPUT103), .B1(new_n883), .B2(new_n889), .ZN(new_n890));
  INV_X1    g465(.A(KEYINPUT100), .ZN(new_n891));
  XNOR2_X1  g466(.A(new_n872), .B(new_n891), .ZN(new_n892));
  NOR2_X1   g467(.A1(new_n882), .A2(new_n865), .ZN(new_n893));
  NOR2_X1   g468(.A1(new_n892), .A2(new_n893), .ZN(new_n894));
  OAI21_X1  g469(.A(KEYINPUT104), .B1(new_n894), .B2(new_n888), .ZN(new_n895));
  INV_X1    g470(.A(KEYINPUT104), .ZN(new_n896));
  NAND3_X1  g471(.A1(new_n883), .A2(new_n896), .A3(new_n889), .ZN(new_n897));
  INV_X1    g472(.A(KEYINPUT103), .ZN(new_n898));
  NAND3_X1  g473(.A1(new_n894), .A2(new_n898), .A3(new_n888), .ZN(new_n899));
  NAND4_X1  g474(.A1(new_n890), .A2(new_n895), .A3(new_n897), .A4(new_n899), .ZN(new_n900));
  MUX2_X1   g475(.A(new_n823), .B(new_n900), .S(G868), .Z(G295));
  MUX2_X1   g476(.A(new_n823), .B(new_n900), .S(G868), .Z(G331));
  XNOR2_X1  g477(.A(G301), .B(G168), .ZN(new_n903));
  INV_X1    g478(.A(new_n903), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n904), .A2(new_n826), .ZN(new_n905));
  NAND3_X1  g480(.A1(new_n903), .A2(new_n824), .A3(new_n825), .ZN(new_n906));
  NAND2_X1  g481(.A1(new_n905), .A2(new_n906), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n881), .A2(new_n907), .ZN(new_n908));
  INV_X1    g483(.A(KEYINPUT105), .ZN(new_n909));
  INV_X1    g484(.A(new_n871), .ZN(new_n910));
  NOR2_X1   g485(.A1(new_n910), .A2(new_n907), .ZN(new_n911));
  INV_X1    g486(.A(new_n911), .ZN(new_n912));
  AND3_X1   g487(.A1(new_n908), .A2(new_n909), .A3(new_n912), .ZN(new_n913));
  AOI21_X1  g488(.A(new_n909), .B1(new_n908), .B2(new_n912), .ZN(new_n914));
  OAI21_X1  g489(.A(new_n886), .B1(new_n913), .B2(new_n914), .ZN(new_n915));
  INV_X1    g490(.A(new_n886), .ZN(new_n916));
  NAND3_X1  g491(.A1(new_n908), .A2(new_n916), .A3(new_n912), .ZN(new_n917));
  AND2_X1   g492(.A1(new_n917), .A2(new_n861), .ZN(new_n918));
  NAND3_X1  g493(.A1(new_n915), .A2(new_n918), .A3(KEYINPUT43), .ZN(new_n919));
  INV_X1    g494(.A(KEYINPUT44), .ZN(new_n920));
  INV_X1    g495(.A(KEYINPUT106), .ZN(new_n921));
  OAI21_X1  g496(.A(new_n886), .B1(new_n912), .B2(new_n921), .ZN(new_n922));
  INV_X1    g497(.A(new_n907), .ZN(new_n923));
  OAI21_X1  g498(.A(new_n910), .B1(new_n923), .B2(new_n875), .ZN(new_n924));
  NAND3_X1  g499(.A1(new_n907), .A2(KEYINPUT41), .A3(new_n874), .ZN(new_n925));
  AOI21_X1  g500(.A(KEYINPUT106), .B1(new_n924), .B2(new_n925), .ZN(new_n926));
  OAI211_X1 g501(.A(new_n861), .B(new_n917), .C1(new_n922), .C2(new_n926), .ZN(new_n927));
  INV_X1    g502(.A(KEYINPUT43), .ZN(new_n928));
  NAND2_X1  g503(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  NAND3_X1  g504(.A1(new_n919), .A2(new_n920), .A3(new_n929), .ZN(new_n930));
  AOI21_X1  g505(.A(new_n920), .B1(new_n927), .B2(KEYINPUT43), .ZN(new_n931));
  NAND3_X1  g506(.A1(new_n915), .A2(new_n918), .A3(new_n928), .ZN(new_n932));
  AND3_X1   g507(.A1(new_n931), .A2(new_n932), .A3(KEYINPUT107), .ZN(new_n933));
  AOI21_X1  g508(.A(KEYINPUT107), .B1(new_n931), .B2(new_n932), .ZN(new_n934));
  OAI21_X1  g509(.A(new_n930), .B1(new_n933), .B2(new_n934), .ZN(G397));
  XNOR2_X1  g510(.A(new_n766), .B(G2067), .ZN(new_n936));
  XNOR2_X1  g511(.A(new_n730), .B(G1996), .ZN(new_n937));
  OR2_X1    g512(.A1(new_n936), .A2(new_n937), .ZN(new_n938));
  AND2_X1   g513(.A1(new_n710), .A2(new_n716), .ZN(new_n939));
  NOR2_X1   g514(.A1(new_n710), .A2(new_n716), .ZN(new_n940));
  NOR3_X1   g515(.A1(new_n938), .A2(new_n939), .A3(new_n940), .ZN(new_n941));
  INV_X1    g516(.A(G1384), .ZN(new_n942));
  NAND2_X1  g517(.A1(new_n503), .A2(new_n942), .ZN(new_n943));
  INV_X1    g518(.A(KEYINPUT45), .ZN(new_n944));
  NAND2_X1  g519(.A1(new_n943), .A2(new_n944), .ZN(new_n945));
  NAND3_X1  g520(.A1(new_n474), .A2(new_n478), .A3(G40), .ZN(new_n946));
  INV_X1    g521(.A(KEYINPUT108), .ZN(new_n947));
  NAND2_X1  g522(.A1(new_n946), .A2(new_n947), .ZN(new_n948));
  NAND4_X1  g523(.A1(new_n474), .A2(new_n478), .A3(KEYINPUT108), .A4(G40), .ZN(new_n949));
  NAND2_X1  g524(.A1(new_n948), .A2(new_n949), .ZN(new_n950));
  NOR2_X1   g525(.A1(new_n945), .A2(new_n950), .ZN(new_n951));
  INV_X1    g526(.A(new_n951), .ZN(new_n952));
  OR3_X1    g527(.A1(new_n952), .A2(G1986), .A3(G290), .ZN(new_n953));
  XNOR2_X1  g528(.A(KEYINPUT126), .B(KEYINPUT48), .ZN(new_n954));
  OAI22_X1  g529(.A1(new_n941), .A2(new_n952), .B1(new_n953), .B2(new_n954), .ZN(new_n955));
  AOI21_X1  g530(.A(new_n955), .B1(new_n953), .B2(new_n954), .ZN(new_n956));
  NOR2_X1   g531(.A1(new_n952), .A2(G1996), .ZN(new_n957));
  XOR2_X1   g532(.A(new_n957), .B(KEYINPUT46), .Z(new_n958));
  OAI21_X1  g533(.A(new_n951), .B1(new_n936), .B2(new_n730), .ZN(new_n959));
  NAND2_X1  g534(.A1(new_n958), .A2(new_n959), .ZN(new_n960));
  XOR2_X1   g535(.A(new_n960), .B(KEYINPUT47), .Z(new_n961));
  XNOR2_X1  g536(.A(new_n940), .B(KEYINPUT125), .ZN(new_n962));
  OAI22_X1  g537(.A1(new_n938), .A2(new_n962), .B1(G2067), .B2(new_n766), .ZN(new_n963));
  AOI211_X1 g538(.A(new_n956), .B(new_n961), .C1(new_n951), .C2(new_n963), .ZN(new_n964));
  OAI21_X1  g539(.A(KEYINPUT57), .B1(new_n565), .B2(new_n569), .ZN(new_n965));
  AOI22_X1  g540(.A1(new_n567), .A2(new_n559), .B1(new_n555), .B2(new_n556), .ZN(new_n966));
  AOI22_X1  g541(.A1(G91), .A2(new_n524), .B1(new_n566), .B2(KEYINPUT71), .ZN(new_n967));
  INV_X1    g542(.A(KEYINPUT57), .ZN(new_n968));
  NAND4_X1  g543(.A1(new_n966), .A2(new_n967), .A3(new_n968), .A4(new_n558), .ZN(new_n969));
  AND2_X1   g544(.A1(new_n965), .A2(new_n969), .ZN(new_n970));
  AND3_X1   g545(.A1(new_n503), .A2(KEYINPUT50), .A3(new_n942), .ZN(new_n971));
  AOI21_X1  g546(.A(KEYINPUT50), .B1(new_n503), .B2(new_n942), .ZN(new_n972));
  OAI211_X1 g547(.A(new_n948), .B(new_n949), .C1(new_n971), .C2(new_n972), .ZN(new_n973));
  NAND2_X1  g548(.A1(new_n973), .A2(new_n783), .ZN(new_n974));
  AND3_X1   g549(.A1(new_n503), .A2(KEYINPUT45), .A3(new_n942), .ZN(new_n975));
  AOI21_X1  g550(.A(KEYINPUT45), .B1(new_n503), .B2(new_n942), .ZN(new_n976));
  NOR2_X1   g551(.A1(new_n975), .A2(new_n976), .ZN(new_n977));
  AND2_X1   g552(.A1(new_n948), .A2(new_n949), .ZN(new_n978));
  XOR2_X1   g553(.A(KEYINPUT56), .B(G2072), .Z(new_n979));
  INV_X1    g554(.A(new_n979), .ZN(new_n980));
  NAND3_X1  g555(.A1(new_n977), .A2(new_n978), .A3(new_n980), .ZN(new_n981));
  AOI21_X1  g556(.A(new_n970), .B1(new_n974), .B2(new_n981), .ZN(new_n982));
  INV_X1    g557(.A(G2067), .ZN(new_n983));
  INV_X1    g558(.A(new_n495), .ZN(new_n984));
  OAI21_X1  g559(.A(new_n984), .B1(new_n481), .B2(new_n482), .ZN(new_n985));
  NAND2_X1  g560(.A1(new_n985), .A2(new_n497), .ZN(new_n986));
  AOI22_X1  g561(.A1(new_n986), .A2(new_n484), .B1(new_n501), .B2(new_n500), .ZN(new_n987));
  AOI21_X1  g562(.A(G1384), .B1(new_n987), .B2(new_n494), .ZN(new_n988));
  AND4_X1   g563(.A1(new_n983), .A2(new_n988), .A3(new_n948), .A4(new_n949), .ZN(new_n989));
  AOI21_X1  g564(.A(new_n989), .B1(new_n973), .B2(new_n809), .ZN(new_n990));
  NOR2_X1   g565(.A1(new_n990), .A2(new_n868), .ZN(new_n991));
  NAND3_X1  g566(.A1(new_n974), .A2(new_n981), .A3(new_n970), .ZN(new_n992));
  AOI21_X1  g567(.A(new_n982), .B1(new_n991), .B2(new_n992), .ZN(new_n993));
  NAND2_X1  g568(.A1(new_n965), .A2(new_n969), .ZN(new_n994));
  NAND2_X1  g569(.A1(new_n988), .A2(KEYINPUT50), .ZN(new_n995));
  INV_X1    g570(.A(KEYINPUT50), .ZN(new_n996));
  NAND2_X1  g571(.A1(new_n943), .A2(new_n996), .ZN(new_n997));
  NAND2_X1  g572(.A1(new_n995), .A2(new_n997), .ZN(new_n998));
  AOI21_X1  g573(.A(G1956), .B1(new_n998), .B2(new_n978), .ZN(new_n999));
  NOR4_X1   g574(.A1(new_n950), .A2(new_n975), .A3(new_n976), .A4(new_n979), .ZN(new_n1000));
  OAI21_X1  g575(.A(new_n994), .B1(new_n999), .B2(new_n1000), .ZN(new_n1001));
  NAND3_X1  g576(.A1(new_n1001), .A2(KEYINPUT61), .A3(new_n992), .ZN(new_n1002));
  INV_X1    g577(.A(KEYINPUT119), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n1002), .A2(new_n1003), .ZN(new_n1004));
  NAND2_X1  g579(.A1(KEYINPUT118), .A2(KEYINPUT59), .ZN(new_n1005));
  NAND3_X1  g580(.A1(new_n503), .A2(KEYINPUT45), .A3(new_n942), .ZN(new_n1006));
  XNOR2_X1  g581(.A(KEYINPUT117), .B(G1996), .ZN(new_n1007));
  NAND4_X1  g582(.A1(new_n978), .A2(new_n945), .A3(new_n1006), .A4(new_n1007), .ZN(new_n1008));
  NAND3_X1  g583(.A1(new_n988), .A2(new_n948), .A3(new_n949), .ZN(new_n1009));
  XOR2_X1   g584(.A(KEYINPUT58), .B(G1341), .Z(new_n1010));
  NAND2_X1  g585(.A1(new_n1009), .A2(new_n1010), .ZN(new_n1011));
  AOI21_X1  g586(.A(new_n547), .B1(new_n1008), .B2(new_n1011), .ZN(new_n1012));
  NOR2_X1   g587(.A1(KEYINPUT118), .A2(KEYINPUT59), .ZN(new_n1013));
  INV_X1    g588(.A(new_n1013), .ZN(new_n1014));
  NOR2_X1   g589(.A1(new_n1012), .A2(new_n1014), .ZN(new_n1015));
  AOI211_X1 g590(.A(new_n1013), .B(new_n547), .C1(new_n1008), .C2(new_n1011), .ZN(new_n1016));
  OAI21_X1  g591(.A(new_n1005), .B1(new_n1015), .B2(new_n1016), .ZN(new_n1017));
  INV_X1    g592(.A(KEYINPUT61), .ZN(new_n1018));
  INV_X1    g593(.A(new_n992), .ZN(new_n1019));
  OAI21_X1  g594(.A(new_n1018), .B1(new_n1019), .B2(new_n982), .ZN(new_n1020));
  NAND4_X1  g595(.A1(new_n1001), .A2(KEYINPUT119), .A3(KEYINPUT61), .A4(new_n992), .ZN(new_n1021));
  NAND4_X1  g596(.A1(new_n1004), .A2(new_n1017), .A3(new_n1020), .A4(new_n1021), .ZN(new_n1022));
  NOR2_X1   g597(.A1(new_n990), .A2(KEYINPUT60), .ZN(new_n1023));
  INV_X1    g598(.A(KEYINPUT120), .ZN(new_n1024));
  NAND4_X1  g599(.A1(new_n990), .A2(new_n1024), .A3(KEYINPUT60), .A4(new_n868), .ZN(new_n1025));
  NAND3_X1  g600(.A1(new_n978), .A2(new_n983), .A3(new_n988), .ZN(new_n1026));
  AOI21_X1  g601(.A(new_n950), .B1(new_n997), .B2(new_n995), .ZN(new_n1027));
  OAI211_X1 g602(.A(new_n1026), .B(KEYINPUT60), .C1(new_n1027), .C2(G1348), .ZN(new_n1028));
  NAND2_X1  g603(.A1(new_n1028), .A2(new_n599), .ZN(new_n1029));
  AND2_X1   g604(.A1(new_n1025), .A2(new_n1029), .ZN(new_n1030));
  OAI21_X1  g605(.A(KEYINPUT120), .B1(new_n1028), .B2(new_n599), .ZN(new_n1031));
  AOI21_X1  g606(.A(new_n1023), .B1(new_n1030), .B2(new_n1031), .ZN(new_n1032));
  OAI21_X1  g607(.A(new_n993), .B1(new_n1022), .B2(new_n1032), .ZN(new_n1033));
  INV_X1    g608(.A(KEYINPUT116), .ZN(new_n1034));
  OAI21_X1  g609(.A(new_n1034), .B1(new_n973), .B2(G2084), .ZN(new_n1035));
  NAND4_X1  g610(.A1(new_n998), .A2(KEYINPUT116), .A3(new_n742), .A4(new_n978), .ZN(new_n1036));
  NAND4_X1  g611(.A1(new_n945), .A2(new_n948), .A3(new_n949), .A4(new_n1006), .ZN(new_n1037));
  NAND2_X1  g612(.A1(new_n1037), .A2(new_n756), .ZN(new_n1038));
  NAND3_X1  g613(.A1(new_n1035), .A2(new_n1036), .A3(new_n1038), .ZN(new_n1039));
  XNOR2_X1  g614(.A(KEYINPUT111), .B(G8), .ZN(new_n1040));
  INV_X1    g615(.A(new_n1040), .ZN(new_n1041));
  NAND3_X1  g616(.A1(new_n1039), .A2(G286), .A3(new_n1041), .ZN(new_n1042));
  INV_X1    g617(.A(KEYINPUT51), .ZN(new_n1043));
  NAND2_X1  g618(.A1(new_n1039), .A2(G8), .ZN(new_n1044));
  NAND2_X1  g619(.A1(G286), .A2(new_n1041), .ZN(new_n1045));
  AOI21_X1  g620(.A(new_n1043), .B1(new_n1044), .B2(new_n1045), .ZN(new_n1046));
  NAND2_X1  g621(.A1(new_n1045), .A2(new_n1043), .ZN(new_n1047));
  AOI21_X1  g622(.A(new_n1047), .B1(new_n1039), .B2(new_n1041), .ZN(new_n1048));
  OAI21_X1  g623(.A(new_n1042), .B1(new_n1046), .B2(new_n1048), .ZN(new_n1049));
  INV_X1    g624(.A(KEYINPUT122), .ZN(new_n1050));
  NAND3_X1  g625(.A1(new_n977), .A2(new_n445), .A3(new_n978), .ZN(new_n1051));
  INV_X1    g626(.A(KEYINPUT53), .ZN(new_n1052));
  OR2_X1    g627(.A1(new_n1051), .A2(new_n1052), .ZN(new_n1053));
  AOI22_X1  g628(.A1(new_n1051), .A2(new_n1052), .B1(new_n754), .B2(new_n973), .ZN(new_n1054));
  NAND3_X1  g629(.A1(new_n1053), .A2(new_n1054), .A3(G301), .ZN(new_n1055));
  NAND2_X1  g630(.A1(new_n1055), .A2(KEYINPUT54), .ZN(new_n1056));
  NOR3_X1   g631(.A1(new_n946), .A2(new_n1052), .A3(G2078), .ZN(new_n1057));
  NAND2_X1  g632(.A1(new_n977), .A2(new_n1057), .ZN(new_n1058));
  AOI21_X1  g633(.A(G301), .B1(new_n1054), .B2(new_n1058), .ZN(new_n1059));
  OAI21_X1  g634(.A(new_n1050), .B1(new_n1056), .B2(new_n1059), .ZN(new_n1060));
  INV_X1    g635(.A(new_n1059), .ZN(new_n1061));
  NAND4_X1  g636(.A1(new_n1061), .A2(KEYINPUT122), .A3(KEYINPUT54), .A4(new_n1055), .ZN(new_n1062));
  NAND2_X1  g637(.A1(new_n1060), .A2(new_n1062), .ZN(new_n1063));
  NAND2_X1  g638(.A1(new_n1009), .A2(new_n1041), .ZN(new_n1064));
  INV_X1    g639(.A(new_n1064), .ZN(new_n1065));
  INV_X1    g640(.A(G288), .ZN(new_n1066));
  NAND2_X1  g641(.A1(new_n1066), .A2(G1976), .ZN(new_n1067));
  INV_X1    g642(.A(G1976), .ZN(new_n1068));
  AOI21_X1  g643(.A(KEYINPUT52), .B1(G288), .B2(new_n1068), .ZN(new_n1069));
  NAND3_X1  g644(.A1(new_n1065), .A2(new_n1067), .A3(new_n1069), .ZN(new_n1070));
  AOI21_X1  g645(.A(new_n1064), .B1(G1976), .B2(new_n1066), .ZN(new_n1071));
  INV_X1    g646(.A(KEYINPUT52), .ZN(new_n1072));
  OAI21_X1  g647(.A(new_n1070), .B1(new_n1071), .B2(new_n1072), .ZN(new_n1073));
  INV_X1    g648(.A(G1981), .ZN(new_n1074));
  NAND4_X1  g649(.A1(new_n577), .A2(new_n581), .A3(new_n582), .A4(new_n1074), .ZN(new_n1075));
  XNOR2_X1  g650(.A(new_n1075), .B(KEYINPUT112), .ZN(new_n1076));
  NAND2_X1  g651(.A1(G305), .A2(G1981), .ZN(new_n1077));
  AND3_X1   g652(.A1(new_n1076), .A2(KEYINPUT49), .A3(new_n1077), .ZN(new_n1078));
  AOI21_X1  g653(.A(KEYINPUT49), .B1(new_n1076), .B2(new_n1077), .ZN(new_n1079));
  NOR3_X1   g654(.A1(new_n1078), .A2(new_n1079), .A3(new_n1064), .ZN(new_n1080));
  NOR2_X1   g655(.A1(new_n1073), .A2(new_n1080), .ZN(new_n1081));
  NOR2_X1   g656(.A1(new_n973), .A2(G2090), .ZN(new_n1082));
  XOR2_X1   g657(.A(KEYINPUT109), .B(G1971), .Z(new_n1083));
  AOI21_X1  g658(.A(new_n1083), .B1(new_n977), .B2(new_n978), .ZN(new_n1084));
  OAI21_X1  g659(.A(KEYINPUT110), .B1(new_n1082), .B2(new_n1084), .ZN(new_n1085));
  INV_X1    g660(.A(new_n1083), .ZN(new_n1086));
  NAND2_X1  g661(.A1(new_n1037), .A2(new_n1086), .ZN(new_n1087));
  INV_X1    g662(.A(KEYINPUT110), .ZN(new_n1088));
  OAI211_X1 g663(.A(new_n1087), .B(new_n1088), .C1(G2090), .C2(new_n973), .ZN(new_n1089));
  NAND2_X1  g664(.A1(G303), .A2(G8), .ZN(new_n1090));
  XNOR2_X1  g665(.A(new_n1090), .B(KEYINPUT55), .ZN(new_n1091));
  INV_X1    g666(.A(new_n1091), .ZN(new_n1092));
  NAND4_X1  g667(.A1(new_n1085), .A2(new_n1089), .A3(new_n1092), .A4(G8), .ZN(new_n1093));
  INV_X1    g668(.A(KEYINPUT115), .ZN(new_n1094));
  NOR2_X1   g669(.A1(new_n973), .A2(new_n1094), .ZN(new_n1095));
  AOI21_X1  g670(.A(KEYINPUT115), .B1(new_n998), .B2(new_n978), .ZN(new_n1096));
  OAI21_X1  g671(.A(new_n805), .B1(new_n1095), .B2(new_n1096), .ZN(new_n1097));
  AOI21_X1  g672(.A(new_n1040), .B1(new_n1097), .B2(new_n1087), .ZN(new_n1098));
  OAI211_X1 g673(.A(new_n1081), .B(new_n1093), .C1(new_n1098), .C2(new_n1092), .ZN(new_n1099));
  XNOR2_X1  g674(.A(KEYINPUT121), .B(KEYINPUT54), .ZN(new_n1100));
  NAND2_X1  g675(.A1(new_n1053), .A2(new_n1054), .ZN(new_n1101));
  NAND2_X1  g676(.A1(new_n1101), .A2(G171), .ZN(new_n1102));
  NAND3_X1  g677(.A1(new_n1054), .A2(G301), .A3(new_n1058), .ZN(new_n1103));
  AOI21_X1  g678(.A(new_n1100), .B1(new_n1102), .B2(new_n1103), .ZN(new_n1104));
  NOR2_X1   g679(.A1(new_n1099), .A2(new_n1104), .ZN(new_n1105));
  NAND4_X1  g680(.A1(new_n1033), .A2(new_n1049), .A3(new_n1063), .A4(new_n1105), .ZN(new_n1106));
  INV_X1    g681(.A(KEYINPUT123), .ZN(new_n1107));
  XOR2_X1   g682(.A(new_n1064), .B(KEYINPUT113), .Z(new_n1108));
  NAND2_X1  g683(.A1(new_n1066), .A2(new_n1068), .ZN(new_n1109));
  OAI21_X1  g684(.A(new_n1076), .B1(new_n1080), .B2(new_n1109), .ZN(new_n1110));
  OAI21_X1  g685(.A(new_n1108), .B1(new_n1110), .B2(KEYINPUT114), .ZN(new_n1111));
  INV_X1    g686(.A(KEYINPUT114), .ZN(new_n1112));
  NAND2_X1  g687(.A1(new_n1076), .A2(new_n1077), .ZN(new_n1113));
  INV_X1    g688(.A(KEYINPUT49), .ZN(new_n1114));
  NAND2_X1  g689(.A1(new_n1113), .A2(new_n1114), .ZN(new_n1115));
  NAND2_X1  g690(.A1(new_n1115), .A2(new_n1065), .ZN(new_n1116));
  OAI211_X1 g691(.A(new_n1068), .B(new_n1066), .C1(new_n1116), .C2(new_n1078), .ZN(new_n1117));
  AOI21_X1  g692(.A(new_n1112), .B1(new_n1117), .B2(new_n1076), .ZN(new_n1118));
  INV_X1    g693(.A(new_n1081), .ZN(new_n1119));
  OAI22_X1  g694(.A1(new_n1111), .A2(new_n1118), .B1(new_n1093), .B2(new_n1119), .ZN(new_n1120));
  INV_X1    g695(.A(KEYINPUT63), .ZN(new_n1121));
  NAND3_X1  g696(.A1(new_n1039), .A2(G168), .A3(new_n1041), .ZN(new_n1122));
  OAI21_X1  g697(.A(new_n1121), .B1(new_n1099), .B2(new_n1122), .ZN(new_n1123));
  NOR2_X1   g698(.A1(new_n1122), .A2(new_n1121), .ZN(new_n1124));
  NAND3_X1  g699(.A1(new_n1085), .A2(new_n1089), .A3(G8), .ZN(new_n1125));
  NAND2_X1  g700(.A1(new_n1125), .A2(new_n1091), .ZN(new_n1126));
  NAND4_X1  g701(.A1(new_n1124), .A2(new_n1126), .A3(new_n1093), .A4(new_n1081), .ZN(new_n1127));
  AOI21_X1  g702(.A(new_n1120), .B1(new_n1123), .B2(new_n1127), .ZN(new_n1128));
  AND3_X1   g703(.A1(new_n1106), .A2(new_n1107), .A3(new_n1128), .ZN(new_n1129));
  AOI21_X1  g704(.A(new_n1107), .B1(new_n1106), .B2(new_n1128), .ZN(new_n1130));
  INV_X1    g705(.A(KEYINPUT62), .ZN(new_n1131));
  OAI211_X1 g706(.A(new_n1131), .B(new_n1042), .C1(new_n1046), .C2(new_n1048), .ZN(new_n1132));
  NAND2_X1  g707(.A1(new_n1081), .A2(new_n1093), .ZN(new_n1133));
  NAND2_X1  g708(.A1(new_n1097), .A2(new_n1087), .ZN(new_n1134));
  AOI21_X1  g709(.A(new_n1092), .B1(new_n1134), .B2(new_n1041), .ZN(new_n1135));
  NOR2_X1   g710(.A1(new_n1133), .A2(new_n1135), .ZN(new_n1136));
  INV_X1    g711(.A(new_n1102), .ZN(new_n1137));
  NAND4_X1  g712(.A1(new_n1132), .A2(new_n1136), .A3(KEYINPUT124), .A4(new_n1137), .ZN(new_n1138));
  NAND2_X1  g713(.A1(new_n1049), .A2(KEYINPUT62), .ZN(new_n1139));
  NAND2_X1  g714(.A1(new_n1138), .A2(new_n1139), .ZN(new_n1140));
  NOR2_X1   g715(.A1(new_n1099), .A2(new_n1102), .ZN(new_n1141));
  AOI21_X1  g716(.A(KEYINPUT124), .B1(new_n1141), .B2(new_n1132), .ZN(new_n1142));
  NOR2_X1   g717(.A1(new_n1140), .A2(new_n1142), .ZN(new_n1143));
  NOR3_X1   g718(.A1(new_n1129), .A2(new_n1130), .A3(new_n1143), .ZN(new_n1144));
  XOR2_X1   g719(.A(G290), .B(G1986), .Z(new_n1145));
  AOI21_X1  g720(.A(new_n952), .B1(new_n941), .B2(new_n1145), .ZN(new_n1146));
  OAI21_X1  g721(.A(new_n964), .B1(new_n1144), .B2(new_n1146), .ZN(G329));
  assign    G231 = 1'b0;
  OR2_X1    g722(.A1(G227), .A2(new_n465), .ZN(new_n1149));
  OAI21_X1  g723(.A(KEYINPUT127), .B1(new_n1149), .B2(G401), .ZN(new_n1150));
  NOR2_X1   g724(.A1(G227), .A2(new_n465), .ZN(new_n1151));
  INV_X1    g725(.A(KEYINPUT127), .ZN(new_n1152));
  AND2_X1   g726(.A1(new_n645), .A2(new_n642), .ZN(new_n1153));
  OAI211_X1 g727(.A(new_n1151), .B(new_n1152), .C1(new_n1153), .C2(new_n641), .ZN(new_n1154));
  AOI21_X1  g728(.A(G229), .B1(new_n1150), .B2(new_n1154), .ZN(new_n1155));
  AND2_X1   g729(.A1(new_n1155), .A2(new_n863), .ZN(new_n1156));
  AND3_X1   g730(.A1(new_n1156), .A2(new_n929), .A3(new_n919), .ZN(G308));
  NAND3_X1  g731(.A1(new_n1156), .A2(new_n929), .A3(new_n919), .ZN(G225));
endmodule


