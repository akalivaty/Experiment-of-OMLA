

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301,
         n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312,
         n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323,
         n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334,
         n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
         n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582;

  XOR2_X1 U323 ( .A(n572), .B(KEYINPUT41), .Z(n553) );
  XOR2_X1 U324 ( .A(n390), .B(n389), .Z(n291) );
  XNOR2_X1 U325 ( .A(n391), .B(n291), .ZN(n392) );
  XNOR2_X1 U326 ( .A(n393), .B(n392), .ZN(n397) );
  NOR2_X1 U327 ( .A1(n530), .A2(n451), .ZN(n562) );
  XNOR2_X1 U328 ( .A(n453), .B(n452), .ZN(n454) );
  XNOR2_X1 U329 ( .A(n455), .B(n454), .ZN(G1349GAT) );
  XNOR2_X1 U330 ( .A(G169GAT), .B(G176GAT), .ZN(n298) );
  XOR2_X1 U331 ( .A(KEYINPUT18), .B(KEYINPUT19), .Z(n293) );
  XNOR2_X1 U332 ( .A(KEYINPUT17), .B(KEYINPUT80), .ZN(n292) );
  XNOR2_X1 U333 ( .A(n293), .B(n292), .ZN(n294) );
  XOR2_X1 U334 ( .A(n294), .B(KEYINPUT81), .Z(n296) );
  XNOR2_X1 U335 ( .A(G190GAT), .B(G183GAT), .ZN(n295) );
  XNOR2_X1 U336 ( .A(n296), .B(n295), .ZN(n297) );
  XOR2_X1 U337 ( .A(n298), .B(n297), .Z(n342) );
  XOR2_X1 U338 ( .A(KEYINPUT84), .B(KEYINPUT83), .Z(n300) );
  XNOR2_X1 U339 ( .A(G15GAT), .B(KEYINPUT79), .ZN(n299) );
  XNOR2_X1 U340 ( .A(n300), .B(n299), .ZN(n301) );
  XOR2_X1 U341 ( .A(n342), .B(n301), .Z(n311) );
  XOR2_X1 U342 ( .A(G127GAT), .B(KEYINPUT0), .Z(n303) );
  XNOR2_X1 U343 ( .A(G113GAT), .B(KEYINPUT78), .ZN(n302) );
  XNOR2_X1 U344 ( .A(n303), .B(n302), .ZN(n441) );
  XOR2_X1 U345 ( .A(G43GAT), .B(G134GAT), .Z(n356) );
  XOR2_X1 U346 ( .A(n441), .B(n356), .Z(n305) );
  NAND2_X1 U347 ( .A1(G227GAT), .A2(G233GAT), .ZN(n304) );
  XNOR2_X1 U348 ( .A(n305), .B(n304), .ZN(n306) );
  XOR2_X1 U349 ( .A(n306), .B(KEYINPUT82), .Z(n309) );
  XNOR2_X1 U350 ( .A(G99GAT), .B(G71GAT), .ZN(n307) );
  XNOR2_X1 U351 ( .A(n307), .B(G120GAT), .ZN(n395) );
  XNOR2_X1 U352 ( .A(n395), .B(KEYINPUT20), .ZN(n308) );
  XNOR2_X1 U353 ( .A(n309), .B(n308), .ZN(n310) );
  XNOR2_X1 U354 ( .A(n311), .B(n310), .ZN(n530) );
  XOR2_X1 U355 ( .A(KEYINPUT22), .B(KEYINPUT86), .Z(n313) );
  XNOR2_X1 U356 ( .A(KEYINPUT24), .B(KEYINPUT91), .ZN(n312) );
  XNOR2_X1 U357 ( .A(n313), .B(n312), .ZN(n317) );
  XOR2_X1 U358 ( .A(KEYINPUT90), .B(KEYINPUT23), .Z(n315) );
  XOR2_X1 U359 ( .A(G141GAT), .B(G22GAT), .Z(n407) );
  XOR2_X1 U360 ( .A(G50GAT), .B(G162GAT), .Z(n355) );
  XNOR2_X1 U361 ( .A(n407), .B(n355), .ZN(n314) );
  XNOR2_X1 U362 ( .A(n315), .B(n314), .ZN(n316) );
  XOR2_X1 U363 ( .A(n317), .B(n316), .Z(n319) );
  NAND2_X1 U364 ( .A1(G228GAT), .A2(G233GAT), .ZN(n318) );
  XNOR2_X1 U365 ( .A(n319), .B(n318), .ZN(n321) );
  XNOR2_X1 U366 ( .A(G155GAT), .B(KEYINPUT3), .ZN(n320) );
  XNOR2_X1 U367 ( .A(n320), .B(KEYINPUT2), .ZN(n430) );
  XOR2_X1 U368 ( .A(n321), .B(n430), .Z(n330) );
  XOR2_X1 U369 ( .A(KEYINPUT21), .B(KEYINPUT87), .Z(n323) );
  XNOR2_X1 U370 ( .A(G218GAT), .B(KEYINPUT89), .ZN(n322) );
  XNOR2_X1 U371 ( .A(n323), .B(n322), .ZN(n324) );
  XOR2_X1 U372 ( .A(n324), .B(KEYINPUT88), .Z(n326) );
  XNOR2_X1 U373 ( .A(G197GAT), .B(G211GAT), .ZN(n325) );
  XNOR2_X1 U374 ( .A(n326), .B(n325), .ZN(n341) );
  XOR2_X1 U375 ( .A(G78GAT), .B(G148GAT), .Z(n328) );
  XNOR2_X1 U376 ( .A(G106GAT), .B(G204GAT), .ZN(n327) );
  XNOR2_X1 U377 ( .A(n328), .B(n327), .ZN(n394) );
  XNOR2_X1 U378 ( .A(n341), .B(n394), .ZN(n329) );
  XNOR2_X1 U379 ( .A(n330), .B(n329), .ZN(n465) );
  XOR2_X1 U380 ( .A(G204GAT), .B(KEYINPUT96), .Z(n332) );
  NAND2_X1 U381 ( .A1(G226GAT), .A2(G233GAT), .ZN(n331) );
  XNOR2_X1 U382 ( .A(n332), .B(n331), .ZN(n333) );
  XOR2_X1 U383 ( .A(G8GAT), .B(KEYINPUT74), .Z(n363) );
  XOR2_X1 U384 ( .A(n333), .B(n363), .Z(n339) );
  INV_X1 U385 ( .A(G64GAT), .ZN(n334) );
  NAND2_X1 U386 ( .A1(G92GAT), .A2(n334), .ZN(n337) );
  INV_X1 U387 ( .A(G92GAT), .ZN(n335) );
  NAND2_X1 U388 ( .A1(n335), .A2(G64GAT), .ZN(n336) );
  NAND2_X1 U389 ( .A1(n337), .A2(n336), .ZN(n380) );
  XNOR2_X1 U390 ( .A(G36GAT), .B(n380), .ZN(n338) );
  XNOR2_X1 U391 ( .A(n339), .B(n338), .ZN(n340) );
  XNOR2_X1 U392 ( .A(n341), .B(n340), .ZN(n344) );
  INV_X1 U393 ( .A(n342), .ZN(n343) );
  XOR2_X1 U394 ( .A(n344), .B(n343), .Z(n457) );
  XNOR2_X1 U395 ( .A(KEYINPUT48), .B(KEYINPUT64), .ZN(n425) );
  XOR2_X1 U396 ( .A(KEYINPUT9), .B(KEYINPUT10), .Z(n346) );
  XNOR2_X1 U397 ( .A(G218GAT), .B(KEYINPUT11), .ZN(n345) );
  XNOR2_X1 U398 ( .A(n346), .B(n345), .ZN(n360) );
  XOR2_X1 U399 ( .A(KEYINPUT68), .B(G85GAT), .Z(n384) );
  XOR2_X1 U400 ( .A(G29GAT), .B(G36GAT), .Z(n348) );
  XNOR2_X1 U401 ( .A(KEYINPUT8), .B(KEYINPUT7), .ZN(n347) );
  XNOR2_X1 U402 ( .A(n348), .B(n347), .ZN(n404) );
  XOR2_X1 U403 ( .A(n384), .B(n404), .Z(n350) );
  NAND2_X1 U404 ( .A1(G232GAT), .A2(G233GAT), .ZN(n349) );
  XNOR2_X1 U405 ( .A(n350), .B(n349), .ZN(n354) );
  XOR2_X1 U406 ( .A(G92GAT), .B(G106GAT), .Z(n352) );
  XNOR2_X1 U407 ( .A(G190GAT), .B(G99GAT), .ZN(n351) );
  XNOR2_X1 U408 ( .A(n352), .B(n351), .ZN(n353) );
  XOR2_X1 U409 ( .A(n354), .B(n353), .Z(n358) );
  XNOR2_X1 U410 ( .A(n356), .B(n355), .ZN(n357) );
  XNOR2_X1 U411 ( .A(n358), .B(n357), .ZN(n359) );
  XNOR2_X1 U412 ( .A(n360), .B(n359), .ZN(n563) );
  XOR2_X1 U413 ( .A(G155GAT), .B(G78GAT), .Z(n362) );
  XNOR2_X1 U414 ( .A(G71GAT), .B(G127GAT), .ZN(n361) );
  XNOR2_X1 U415 ( .A(n362), .B(n361), .ZN(n364) );
  XOR2_X1 U416 ( .A(n364), .B(n363), .Z(n366) );
  XNOR2_X1 U417 ( .A(G22GAT), .B(G211GAT), .ZN(n365) );
  XNOR2_X1 U418 ( .A(n366), .B(n365), .ZN(n371) );
  XOR2_X1 U419 ( .A(KEYINPUT13), .B(G57GAT), .Z(n381) );
  XNOR2_X1 U420 ( .A(G15GAT), .B(G1GAT), .ZN(n367) );
  XNOR2_X1 U421 ( .A(n367), .B(KEYINPUT66), .ZN(n403) );
  XOR2_X1 U422 ( .A(n381), .B(n403), .Z(n369) );
  NAND2_X1 U423 ( .A1(G231GAT), .A2(G233GAT), .ZN(n368) );
  XNOR2_X1 U424 ( .A(n369), .B(n368), .ZN(n370) );
  XOR2_X1 U425 ( .A(n371), .B(n370), .Z(n379) );
  XOR2_X1 U426 ( .A(KEYINPUT76), .B(KEYINPUT77), .Z(n373) );
  XNOR2_X1 U427 ( .A(G183GAT), .B(G64GAT), .ZN(n372) );
  XNOR2_X1 U428 ( .A(n373), .B(n372), .ZN(n377) );
  XOR2_X1 U429 ( .A(KEYINPUT14), .B(KEYINPUT12), .Z(n375) );
  XNOR2_X1 U430 ( .A(KEYINPUT75), .B(KEYINPUT15), .ZN(n374) );
  XNOR2_X1 U431 ( .A(n375), .B(n374), .ZN(n376) );
  XNOR2_X1 U432 ( .A(n377), .B(n376), .ZN(n378) );
  XOR2_X1 U433 ( .A(n379), .B(n378), .Z(n576) );
  INV_X1 U434 ( .A(n576), .ZN(n488) );
  XOR2_X1 U435 ( .A(KEYINPUT113), .B(KEYINPUT46), .Z(n414) );
  XOR2_X1 U436 ( .A(KEYINPUT32), .B(n380), .Z(n383) );
  XNOR2_X1 U437 ( .A(G176GAT), .B(n381), .ZN(n382) );
  XOR2_X1 U438 ( .A(n383), .B(n382), .Z(n385) );
  XNOR2_X1 U439 ( .A(n385), .B(n384), .ZN(n393) );
  XOR2_X1 U440 ( .A(KEYINPUT33), .B(KEYINPUT31), .Z(n387) );
  NAND2_X1 U441 ( .A1(G230GAT), .A2(G233GAT), .ZN(n386) );
  XNOR2_X1 U442 ( .A(n387), .B(n386), .ZN(n388) );
  XNOR2_X1 U443 ( .A(KEYINPUT71), .B(n388), .ZN(n391) );
  XOR2_X1 U444 ( .A(KEYINPUT67), .B(KEYINPUT70), .Z(n390) );
  XNOR2_X1 U445 ( .A(KEYINPUT69), .B(KEYINPUT72), .ZN(n389) );
  XNOR2_X1 U446 ( .A(n395), .B(n394), .ZN(n396) );
  XNOR2_X1 U447 ( .A(n397), .B(n396), .ZN(n572) );
  XOR2_X1 U448 ( .A(KEYINPUT29), .B(G113GAT), .Z(n399) );
  XNOR2_X1 U449 ( .A(G169GAT), .B(G197GAT), .ZN(n398) );
  XNOR2_X1 U450 ( .A(n399), .B(n398), .ZN(n412) );
  XOR2_X1 U451 ( .A(G8GAT), .B(KEYINPUT65), .Z(n401) );
  NAND2_X1 U452 ( .A1(G229GAT), .A2(G233GAT), .ZN(n400) );
  XNOR2_X1 U453 ( .A(n401), .B(n400), .ZN(n402) );
  XOR2_X1 U454 ( .A(n402), .B(KEYINPUT30), .Z(n406) );
  XNOR2_X1 U455 ( .A(n404), .B(n403), .ZN(n405) );
  XNOR2_X1 U456 ( .A(n406), .B(n405), .ZN(n408) );
  XOR2_X1 U457 ( .A(n408), .B(n407), .Z(n410) );
  XNOR2_X1 U458 ( .A(G50GAT), .B(G43GAT), .ZN(n409) );
  XNOR2_X1 U459 ( .A(n410), .B(n409), .ZN(n411) );
  XOR2_X1 U460 ( .A(n412), .B(n411), .Z(n502) );
  INV_X1 U461 ( .A(n502), .ZN(n568) );
  NAND2_X1 U462 ( .A1(n553), .A2(n568), .ZN(n413) );
  XNOR2_X1 U463 ( .A(n414), .B(n413), .ZN(n415) );
  NAND2_X1 U464 ( .A1(n488), .A2(n415), .ZN(n416) );
  NOR2_X1 U465 ( .A1(n563), .A2(n416), .ZN(n417) );
  XNOR2_X1 U466 ( .A(n417), .B(KEYINPUT47), .ZN(n423) );
  XNOR2_X1 U467 ( .A(KEYINPUT36), .B(KEYINPUT103), .ZN(n418) );
  XNOR2_X1 U468 ( .A(n418), .B(n563), .ZN(n580) );
  NOR2_X1 U469 ( .A1(n488), .A2(n580), .ZN(n419) );
  XOR2_X1 U470 ( .A(KEYINPUT45), .B(n419), .Z(n420) );
  NOR2_X1 U471 ( .A1(n572), .A2(n420), .ZN(n421) );
  NAND2_X1 U472 ( .A1(n421), .A2(n502), .ZN(n422) );
  NAND2_X1 U473 ( .A1(n423), .A2(n422), .ZN(n424) );
  XNOR2_X1 U474 ( .A(n425), .B(n424), .ZN(n528) );
  NAND2_X1 U475 ( .A1(n457), .A2(n528), .ZN(n426) );
  XNOR2_X1 U476 ( .A(n426), .B(KEYINPUT54), .ZN(n427) );
  XNOR2_X1 U477 ( .A(n427), .B(KEYINPUT125), .ZN(n449) );
  XOR2_X1 U478 ( .A(KEYINPUT4), .B(KEYINPUT5), .Z(n429) );
  XNOR2_X1 U479 ( .A(KEYINPUT94), .B(KEYINPUT93), .ZN(n428) );
  XNOR2_X1 U480 ( .A(n429), .B(n428), .ZN(n434) );
  XOR2_X1 U481 ( .A(n430), .B(KEYINPUT95), .Z(n432) );
  NAND2_X1 U482 ( .A1(G225GAT), .A2(G233GAT), .ZN(n431) );
  XNOR2_X1 U483 ( .A(n432), .B(n431), .ZN(n433) );
  XNOR2_X1 U484 ( .A(n434), .B(n433), .ZN(n448) );
  XOR2_X1 U485 ( .A(G148GAT), .B(G120GAT), .Z(n436) );
  XNOR2_X1 U486 ( .A(G1GAT), .B(G141GAT), .ZN(n435) );
  XNOR2_X1 U487 ( .A(n436), .B(n435), .ZN(n440) );
  XOR2_X1 U488 ( .A(KEYINPUT1), .B(KEYINPUT6), .Z(n438) );
  XNOR2_X1 U489 ( .A(G57GAT), .B(KEYINPUT92), .ZN(n437) );
  XNOR2_X1 U490 ( .A(n438), .B(n437), .ZN(n439) );
  XOR2_X1 U491 ( .A(n440), .B(n439), .Z(n446) );
  XOR2_X1 U492 ( .A(G85GAT), .B(G162GAT), .Z(n443) );
  XNOR2_X1 U493 ( .A(G29GAT), .B(n441), .ZN(n442) );
  XNOR2_X1 U494 ( .A(n443), .B(n442), .ZN(n444) );
  XNOR2_X1 U495 ( .A(G134GAT), .B(n444), .ZN(n445) );
  XNOR2_X1 U496 ( .A(n446), .B(n445), .ZN(n447) );
  XOR2_X1 U497 ( .A(n448), .B(n447), .Z(n471) );
  INV_X1 U498 ( .A(n471), .ZN(n515) );
  NAND2_X1 U499 ( .A1(n449), .A2(n515), .ZN(n567) );
  NOR2_X1 U500 ( .A1(n465), .A2(n567), .ZN(n450) );
  XNOR2_X1 U501 ( .A(n450), .B(KEYINPUT55), .ZN(n451) );
  NAND2_X1 U502 ( .A1(n562), .A2(n553), .ZN(n455) );
  XOR2_X1 U503 ( .A(KEYINPUT57), .B(KEYINPUT126), .Z(n453) );
  XNOR2_X1 U504 ( .A(G176GAT), .B(KEYINPUT56), .ZN(n452) );
  NOR2_X1 U505 ( .A1(n502), .A2(n572), .ZN(n456) );
  XOR2_X1 U506 ( .A(KEYINPUT73), .B(n456), .Z(n491) );
  INV_X1 U507 ( .A(n457), .ZN(n519) );
  XNOR2_X1 U508 ( .A(KEYINPUT27), .B(n519), .ZN(n468) );
  NOR2_X1 U509 ( .A1(n515), .A2(n468), .ZN(n458) );
  XOR2_X1 U510 ( .A(KEYINPUT97), .B(n458), .Z(n527) );
  XOR2_X1 U511 ( .A(n465), .B(KEYINPUT28), .Z(n532) );
  NAND2_X1 U512 ( .A1(n527), .A2(n532), .ZN(n460) );
  XNOR2_X1 U513 ( .A(KEYINPUT85), .B(n530), .ZN(n459) );
  NOR2_X1 U514 ( .A1(n460), .A2(n459), .ZN(n474) );
  XNOR2_X1 U515 ( .A(KEYINPUT25), .B(KEYINPUT100), .ZN(n461) );
  XNOR2_X1 U516 ( .A(n461), .B(KEYINPUT99), .ZN(n464) );
  NOR2_X1 U517 ( .A1(n530), .A2(n519), .ZN(n462) );
  NOR2_X1 U518 ( .A1(n465), .A2(n462), .ZN(n463) );
  XNOR2_X1 U519 ( .A(n464), .B(n463), .ZN(n470) );
  NAND2_X1 U520 ( .A1(n465), .A2(n530), .ZN(n466) );
  XNOR2_X1 U521 ( .A(n466), .B(KEYINPUT26), .ZN(n467) );
  XNOR2_X1 U522 ( .A(KEYINPUT98), .B(n467), .ZN(n566) );
  NOR2_X1 U523 ( .A1(n468), .A2(n566), .ZN(n469) );
  NOR2_X1 U524 ( .A1(n470), .A2(n469), .ZN(n472) );
  NOR2_X1 U525 ( .A1(n472), .A2(n471), .ZN(n473) );
  NOR2_X1 U526 ( .A1(n474), .A2(n473), .ZN(n486) );
  NOR2_X1 U527 ( .A1(n488), .A2(n563), .ZN(n475) );
  XOR2_X1 U528 ( .A(KEYINPUT16), .B(n475), .Z(n476) );
  NOR2_X1 U529 ( .A1(n486), .A2(n476), .ZN(n477) );
  XOR2_X1 U530 ( .A(KEYINPUT101), .B(n477), .Z(n503) );
  NAND2_X1 U531 ( .A1(n491), .A2(n503), .ZN(n484) );
  NOR2_X1 U532 ( .A1(n515), .A2(n484), .ZN(n479) );
  XNOR2_X1 U533 ( .A(KEYINPUT34), .B(KEYINPUT102), .ZN(n478) );
  XNOR2_X1 U534 ( .A(n479), .B(n478), .ZN(n480) );
  XOR2_X1 U535 ( .A(G1GAT), .B(n480), .Z(G1324GAT) );
  NOR2_X1 U536 ( .A1(n519), .A2(n484), .ZN(n481) );
  XOR2_X1 U537 ( .A(G8GAT), .B(n481), .Z(G1325GAT) );
  NOR2_X1 U538 ( .A1(n530), .A2(n484), .ZN(n483) );
  XNOR2_X1 U539 ( .A(G15GAT), .B(KEYINPUT35), .ZN(n482) );
  XNOR2_X1 U540 ( .A(n483), .B(n482), .ZN(G1326GAT) );
  NOR2_X1 U541 ( .A1(n532), .A2(n484), .ZN(n485) );
  XOR2_X1 U542 ( .A(G22GAT), .B(n485), .Z(G1327GAT) );
  XNOR2_X1 U543 ( .A(G29GAT), .B(KEYINPUT39), .ZN(n494) );
  XNOR2_X1 U544 ( .A(KEYINPUT37), .B(KEYINPUT104), .ZN(n490) );
  NOR2_X1 U545 ( .A1(n486), .A2(n580), .ZN(n487) );
  NAND2_X1 U546 ( .A1(n488), .A2(n487), .ZN(n489) );
  XNOR2_X1 U547 ( .A(n490), .B(n489), .ZN(n513) );
  NAND2_X1 U548 ( .A1(n491), .A2(n513), .ZN(n492) );
  XNOR2_X1 U549 ( .A(KEYINPUT38), .B(n492), .ZN(n500) );
  NOR2_X1 U550 ( .A1(n515), .A2(n500), .ZN(n493) );
  XNOR2_X1 U551 ( .A(n494), .B(n493), .ZN(G1328GAT) );
  NOR2_X1 U552 ( .A1(n519), .A2(n500), .ZN(n495) );
  XOR2_X1 U553 ( .A(G36GAT), .B(n495), .Z(G1329GAT) );
  XOR2_X1 U554 ( .A(KEYINPUT40), .B(KEYINPUT105), .Z(n497) );
  XNOR2_X1 U555 ( .A(G43GAT), .B(KEYINPUT106), .ZN(n496) );
  XNOR2_X1 U556 ( .A(n497), .B(n496), .ZN(n499) );
  NOR2_X1 U557 ( .A1(n530), .A2(n500), .ZN(n498) );
  XOR2_X1 U558 ( .A(n499), .B(n498), .Z(G1330GAT) );
  NOR2_X1 U559 ( .A1(n532), .A2(n500), .ZN(n501) );
  XOR2_X1 U560 ( .A(G50GAT), .B(n501), .Z(G1331GAT) );
  AND2_X1 U561 ( .A1(n502), .A2(n553), .ZN(n514) );
  NAND2_X1 U562 ( .A1(n503), .A2(n514), .ZN(n509) );
  NOR2_X1 U563 ( .A1(n515), .A2(n509), .ZN(n505) );
  XNOR2_X1 U564 ( .A(KEYINPUT107), .B(KEYINPUT42), .ZN(n504) );
  XNOR2_X1 U565 ( .A(n505), .B(n504), .ZN(n506) );
  XNOR2_X1 U566 ( .A(G57GAT), .B(n506), .ZN(G1332GAT) );
  NOR2_X1 U567 ( .A1(n519), .A2(n509), .ZN(n507) );
  XOR2_X1 U568 ( .A(G64GAT), .B(n507), .Z(G1333GAT) );
  NOR2_X1 U569 ( .A1(n530), .A2(n509), .ZN(n508) );
  XOR2_X1 U570 ( .A(G71GAT), .B(n508), .Z(G1334GAT) );
  NOR2_X1 U571 ( .A1(n532), .A2(n509), .ZN(n511) );
  XNOR2_X1 U572 ( .A(KEYINPUT108), .B(KEYINPUT43), .ZN(n510) );
  XNOR2_X1 U573 ( .A(n511), .B(n510), .ZN(n512) );
  XNOR2_X1 U574 ( .A(G78GAT), .B(n512), .ZN(G1335GAT) );
  NAND2_X1 U575 ( .A1(n514), .A2(n513), .ZN(n523) );
  NOR2_X1 U576 ( .A1(n515), .A2(n523), .ZN(n517) );
  XNOR2_X1 U577 ( .A(KEYINPUT109), .B(KEYINPUT110), .ZN(n516) );
  XNOR2_X1 U578 ( .A(n517), .B(n516), .ZN(n518) );
  XNOR2_X1 U579 ( .A(G85GAT), .B(n518), .ZN(G1336GAT) );
  NOR2_X1 U580 ( .A1(n519), .A2(n523), .ZN(n520) );
  XOR2_X1 U581 ( .A(G92GAT), .B(n520), .Z(G1337GAT) );
  NOR2_X1 U582 ( .A1(n530), .A2(n523), .ZN(n522) );
  XNOR2_X1 U583 ( .A(G99GAT), .B(KEYINPUT111), .ZN(n521) );
  XNOR2_X1 U584 ( .A(n522), .B(n521), .ZN(G1338GAT) );
  NOR2_X1 U585 ( .A1(n532), .A2(n523), .ZN(n525) );
  XNOR2_X1 U586 ( .A(KEYINPUT44), .B(KEYINPUT112), .ZN(n524) );
  XNOR2_X1 U587 ( .A(n525), .B(n524), .ZN(n526) );
  XOR2_X1 U588 ( .A(G106GAT), .B(n526), .Z(G1339GAT) );
  NAND2_X1 U589 ( .A1(n528), .A2(n527), .ZN(n529) );
  XNOR2_X1 U590 ( .A(n529), .B(KEYINPUT114), .ZN(n545) );
  NOR2_X1 U591 ( .A1(n530), .A2(n545), .ZN(n531) );
  NAND2_X1 U592 ( .A1(n532), .A2(n531), .ZN(n533) );
  XNOR2_X1 U593 ( .A(KEYINPUT115), .B(n533), .ZN(n541) );
  NAND2_X1 U594 ( .A1(n568), .A2(n541), .ZN(n534) );
  XNOR2_X1 U595 ( .A(n534), .B(KEYINPUT116), .ZN(n535) );
  XNOR2_X1 U596 ( .A(G113GAT), .B(n535), .ZN(G1340GAT) );
  XOR2_X1 U597 ( .A(KEYINPUT117), .B(KEYINPUT49), .Z(n537) );
  NAND2_X1 U598 ( .A1(n541), .A2(n553), .ZN(n536) );
  XNOR2_X1 U599 ( .A(n537), .B(n536), .ZN(n538) );
  XOR2_X1 U600 ( .A(G120GAT), .B(n538), .Z(G1341GAT) );
  NAND2_X1 U601 ( .A1(n576), .A2(n541), .ZN(n539) );
  XNOR2_X1 U602 ( .A(n539), .B(KEYINPUT50), .ZN(n540) );
  XNOR2_X1 U603 ( .A(G127GAT), .B(n540), .ZN(G1342GAT) );
  XOR2_X1 U604 ( .A(KEYINPUT51), .B(KEYINPUT118), .Z(n543) );
  NAND2_X1 U605 ( .A1(n541), .A2(n563), .ZN(n542) );
  XNOR2_X1 U606 ( .A(n543), .B(n542), .ZN(n544) );
  XNOR2_X1 U607 ( .A(G134GAT), .B(n544), .ZN(G1343GAT) );
  NOR2_X1 U608 ( .A1(n545), .A2(n566), .ZN(n546) );
  XOR2_X1 U609 ( .A(KEYINPUT119), .B(n546), .Z(n558) );
  NAND2_X1 U610 ( .A1(n558), .A2(n568), .ZN(n547) );
  XNOR2_X1 U611 ( .A(G141GAT), .B(n547), .ZN(G1344GAT) );
  XOR2_X1 U612 ( .A(KEYINPUT120), .B(KEYINPUT122), .Z(n549) );
  XNOR2_X1 U613 ( .A(KEYINPUT52), .B(KEYINPUT53), .ZN(n548) );
  XNOR2_X1 U614 ( .A(n549), .B(n548), .ZN(n550) );
  XOR2_X1 U615 ( .A(n550), .B(KEYINPUT123), .Z(n552) );
  XNOR2_X1 U616 ( .A(G148GAT), .B(KEYINPUT121), .ZN(n551) );
  XNOR2_X1 U617 ( .A(n552), .B(n551), .ZN(n555) );
  NAND2_X1 U618 ( .A1(n558), .A2(n553), .ZN(n554) );
  XOR2_X1 U619 ( .A(n555), .B(n554), .Z(G1345GAT) );
  NAND2_X1 U620 ( .A1(n576), .A2(n558), .ZN(n556) );
  XNOR2_X1 U621 ( .A(n556), .B(KEYINPUT124), .ZN(n557) );
  XNOR2_X1 U622 ( .A(G155GAT), .B(n557), .ZN(G1346GAT) );
  NAND2_X1 U623 ( .A1(n563), .A2(n558), .ZN(n559) );
  XNOR2_X1 U624 ( .A(n559), .B(G162GAT), .ZN(G1347GAT) );
  NAND2_X1 U625 ( .A1(n568), .A2(n562), .ZN(n560) );
  XNOR2_X1 U626 ( .A(n560), .B(G169GAT), .ZN(G1348GAT) );
  NAND2_X1 U627 ( .A1(n576), .A2(n562), .ZN(n561) );
  XNOR2_X1 U628 ( .A(n561), .B(G183GAT), .ZN(G1350GAT) );
  NAND2_X1 U629 ( .A1(n563), .A2(n562), .ZN(n564) );
  XNOR2_X1 U630 ( .A(n564), .B(KEYINPUT58), .ZN(n565) );
  XNOR2_X1 U631 ( .A(G190GAT), .B(n565), .ZN(G1351GAT) );
  XOR2_X1 U632 ( .A(KEYINPUT60), .B(KEYINPUT59), .Z(n570) );
  NOR2_X1 U633 ( .A1(n567), .A2(n566), .ZN(n578) );
  NAND2_X1 U634 ( .A1(n578), .A2(n568), .ZN(n569) );
  XNOR2_X1 U635 ( .A(n570), .B(n569), .ZN(n571) );
  XNOR2_X1 U636 ( .A(G197GAT), .B(n571), .ZN(G1352GAT) );
  XOR2_X1 U637 ( .A(KEYINPUT61), .B(KEYINPUT127), .Z(n574) );
  NAND2_X1 U638 ( .A1(n578), .A2(n572), .ZN(n573) );
  XNOR2_X1 U639 ( .A(n574), .B(n573), .ZN(n575) );
  XOR2_X1 U640 ( .A(G204GAT), .B(n575), .Z(G1353GAT) );
  NAND2_X1 U641 ( .A1(n576), .A2(n578), .ZN(n577) );
  XNOR2_X1 U642 ( .A(n577), .B(G211GAT), .ZN(G1354GAT) );
  INV_X1 U643 ( .A(n578), .ZN(n579) );
  NOR2_X1 U644 ( .A1(n580), .A2(n579), .ZN(n581) );
  XOR2_X1 U645 ( .A(KEYINPUT62), .B(n581), .Z(n582) );
  XNOR2_X1 U646 ( .A(G218GAT), .B(n582), .ZN(G1355GAT) );
endmodule

