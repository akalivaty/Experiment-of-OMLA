//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 0 1 1 1 1 1 0 0 1 0 0 1 1 0 1 1 1 0 1 0 0 0 1 0 0 0 1 1 1 0 1 0 1 1 0 0 0 0 1 0 1 0 0 1 0 1 1 1 1 1 0 0 0 0 0 1 0 1 0 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:23:13 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n620, new_n621, new_n622,
    new_n623, new_n624, new_n625, new_n626, new_n628, new_n629, new_n630,
    new_n631, new_n632, new_n633, new_n634, new_n635, new_n636, new_n637,
    new_n638, new_n639, new_n640, new_n641, new_n643, new_n644, new_n645,
    new_n646, new_n647, new_n648, new_n649, new_n650, new_n651, new_n652,
    new_n653, new_n654, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n692, new_n693, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n718, new_n719, new_n720, new_n721,
    new_n722, new_n723, new_n724, new_n725, new_n726, new_n727, new_n728,
    new_n729, new_n730, new_n731, new_n732, new_n733, new_n734, new_n735,
    new_n736, new_n737, new_n738, new_n740, new_n741, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n764, new_n765, new_n766,
    new_n767, new_n768, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n788, new_n789,
    new_n790, new_n791, new_n792, new_n793, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n921, new_n922, new_n923, new_n924, new_n926, new_n927,
    new_n928, new_n929, new_n930, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n939, new_n940, new_n942, new_n943,
    new_n944, new_n945, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n973,
    new_n974, new_n975, new_n976, new_n977, new_n978, new_n979, new_n980,
    new_n981, new_n982, new_n983;
  INV_X1    g000(.A(G952), .ZN(new_n187));
  AOI211_X1 g001(.A(G953), .B(new_n187), .C1(G234), .C2(G237), .ZN(new_n188));
  INV_X1    g002(.A(G902), .ZN(new_n189));
  INV_X1    g003(.A(G953), .ZN(new_n190));
  AOI211_X1 g004(.A(new_n189), .B(new_n190), .C1(G234), .C2(G237), .ZN(new_n191));
  XNOR2_X1  g005(.A(KEYINPUT21), .B(G898), .ZN(new_n192));
  AOI21_X1  g006(.A(new_n188), .B1(new_n191), .B2(new_n192), .ZN(new_n193));
  INV_X1    g007(.A(new_n193), .ZN(new_n194));
  OAI21_X1  g008(.A(G214), .B1(G237), .B2(G902), .ZN(new_n195));
  XOR2_X1   g009(.A(new_n195), .B(KEYINPUT82), .Z(new_n196));
  INV_X1    g010(.A(new_n196), .ZN(new_n197));
  OAI21_X1  g011(.A(G210), .B1(G237), .B2(G902), .ZN(new_n198));
  INV_X1    g012(.A(G104), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n199), .A2(G107), .ZN(new_n200));
  OR2_X1    g014(.A1(KEYINPUT75), .A2(KEYINPUT3), .ZN(new_n201));
  INV_X1    g015(.A(G107), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n202), .A2(G104), .ZN(new_n203));
  OAI21_X1  g017(.A(new_n200), .B1(new_n201), .B2(new_n203), .ZN(new_n204));
  NOR2_X1   g018(.A1(KEYINPUT75), .A2(KEYINPUT3), .ZN(new_n205));
  NOR2_X1   g019(.A1(new_n199), .A2(G107), .ZN(new_n206));
  NAND2_X1  g020(.A1(KEYINPUT75), .A2(KEYINPUT3), .ZN(new_n207));
  AOI21_X1  g021(.A(new_n205), .B1(new_n206), .B2(new_n207), .ZN(new_n208));
  OAI21_X1  g022(.A(G101), .B1(new_n204), .B2(new_n208), .ZN(new_n209));
  AND2_X1   g023(.A1(KEYINPUT75), .A2(KEYINPUT3), .ZN(new_n210));
  OAI21_X1  g024(.A(new_n201), .B1(new_n203), .B2(new_n210), .ZN(new_n211));
  INV_X1    g025(.A(G101), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n206), .A2(new_n205), .ZN(new_n213));
  NAND4_X1  g027(.A1(new_n211), .A2(new_n212), .A3(new_n200), .A4(new_n213), .ZN(new_n214));
  NAND3_X1  g028(.A1(new_n209), .A2(KEYINPUT4), .A3(new_n214), .ZN(new_n215));
  INV_X1    g029(.A(G119), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n216), .A2(G116), .ZN(new_n217));
  INV_X1    g031(.A(G116), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n218), .A2(G119), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n217), .A2(new_n219), .ZN(new_n220));
  NAND2_X1  g034(.A1(KEYINPUT2), .A2(G113), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n221), .A2(KEYINPUT67), .ZN(new_n222));
  INV_X1    g036(.A(KEYINPUT67), .ZN(new_n223));
  NAND3_X1  g037(.A1(new_n223), .A2(KEYINPUT2), .A3(G113), .ZN(new_n224));
  AND2_X1   g038(.A1(new_n222), .A2(new_n224), .ZN(new_n225));
  NOR2_X1   g039(.A1(KEYINPUT2), .A2(G113), .ZN(new_n226));
  OAI21_X1  g040(.A(new_n220), .B1(new_n225), .B2(new_n226), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n222), .A2(new_n224), .ZN(new_n228));
  OR2_X1    g042(.A1(KEYINPUT2), .A2(G113), .ZN(new_n229));
  NAND4_X1  g043(.A1(new_n228), .A2(new_n229), .A3(new_n217), .A4(new_n219), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n227), .A2(new_n230), .ZN(new_n231));
  INV_X1    g045(.A(KEYINPUT83), .ZN(new_n232));
  INV_X1    g046(.A(KEYINPUT4), .ZN(new_n233));
  OAI211_X1 g047(.A(new_n233), .B(G101), .C1(new_n204), .C2(new_n208), .ZN(new_n234));
  NAND4_X1  g048(.A1(new_n215), .A2(new_n231), .A3(new_n232), .A4(new_n234), .ZN(new_n235));
  NOR2_X1   g049(.A1(new_n202), .A2(G104), .ZN(new_n236));
  OAI21_X1  g050(.A(G101), .B1(new_n206), .B2(new_n236), .ZN(new_n237));
  AND2_X1   g051(.A1(new_n214), .A2(new_n237), .ZN(new_n238));
  OR2_X1    g052(.A1(new_n217), .A2(KEYINPUT5), .ZN(new_n239));
  NAND3_X1  g053(.A1(new_n217), .A2(new_n219), .A3(KEYINPUT5), .ZN(new_n240));
  NAND4_X1  g054(.A1(new_n239), .A2(KEYINPUT84), .A3(new_n240), .A4(G113), .ZN(new_n241));
  NAND3_X1  g055(.A1(new_n239), .A2(G113), .A3(new_n240), .ZN(new_n242));
  INV_X1    g056(.A(KEYINPUT84), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n242), .A2(new_n243), .ZN(new_n244));
  NAND4_X1  g058(.A1(new_n238), .A2(new_n230), .A3(new_n241), .A4(new_n244), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n235), .A2(new_n245), .ZN(new_n246));
  AOI21_X1  g060(.A(new_n236), .B1(new_n205), .B2(new_n206), .ZN(new_n247));
  AOI21_X1  g061(.A(new_n212), .B1(new_n247), .B2(new_n211), .ZN(new_n248));
  AOI22_X1  g062(.A1(new_n233), .A2(new_n248), .B1(new_n227), .B2(new_n230), .ZN(new_n249));
  AOI21_X1  g063(.A(new_n232), .B1(new_n249), .B2(new_n215), .ZN(new_n250));
  OAI21_X1  g064(.A(KEYINPUT85), .B1(new_n246), .B2(new_n250), .ZN(new_n251));
  NAND3_X1  g065(.A1(new_n215), .A2(new_n231), .A3(new_n234), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n252), .A2(KEYINPUT83), .ZN(new_n253));
  INV_X1    g067(.A(KEYINPUT85), .ZN(new_n254));
  NAND4_X1  g068(.A1(new_n253), .A2(new_n254), .A3(new_n245), .A4(new_n235), .ZN(new_n255));
  XNOR2_X1  g069(.A(G110), .B(G122), .ZN(new_n256));
  INV_X1    g070(.A(new_n256), .ZN(new_n257));
  NAND3_X1  g071(.A1(new_n251), .A2(new_n255), .A3(new_n257), .ZN(new_n258));
  NAND4_X1  g072(.A1(new_n253), .A2(new_n245), .A3(new_n235), .A4(new_n256), .ZN(new_n259));
  AND2_X1   g073(.A1(new_n259), .A2(KEYINPUT6), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n258), .A2(new_n260), .ZN(new_n261));
  INV_X1    g075(.A(G143), .ZN(new_n262));
  OAI21_X1  g076(.A(KEYINPUT1), .B1(new_n262), .B2(G146), .ZN(new_n263));
  NOR2_X1   g077(.A1(new_n262), .A2(G146), .ZN(new_n264));
  INV_X1    g078(.A(G146), .ZN(new_n265));
  NOR2_X1   g079(.A1(new_n265), .A2(G143), .ZN(new_n266));
  OAI211_X1 g080(.A(G128), .B(new_n263), .C1(new_n264), .C2(new_n266), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n265), .A2(G143), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n262), .A2(G146), .ZN(new_n269));
  INV_X1    g083(.A(G128), .ZN(new_n270));
  OAI211_X1 g084(.A(new_n268), .B(new_n269), .C1(KEYINPUT1), .C2(new_n270), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n267), .A2(new_n271), .ZN(new_n272));
  INV_X1    g086(.A(G125), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n272), .A2(new_n273), .ZN(new_n274));
  NAND4_X1  g088(.A1(new_n268), .A2(new_n269), .A3(KEYINPUT0), .A4(G128), .ZN(new_n275));
  NOR2_X1   g089(.A1(new_n264), .A2(new_n266), .ZN(new_n276));
  XNOR2_X1  g090(.A(KEYINPUT0), .B(G128), .ZN(new_n277));
  OAI21_X1  g091(.A(new_n275), .B1(new_n276), .B2(new_n277), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n278), .A2(G125), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n274), .A2(new_n279), .ZN(new_n280));
  INV_X1    g094(.A(G224), .ZN(new_n281));
  NOR2_X1   g095(.A1(new_n281), .A2(G953), .ZN(new_n282));
  NOR2_X1   g096(.A1(new_n280), .A2(new_n282), .ZN(new_n283));
  INV_X1    g097(.A(new_n282), .ZN(new_n284));
  AOI21_X1  g098(.A(new_n284), .B1(new_n274), .B2(new_n279), .ZN(new_n285));
  NOR2_X1   g099(.A1(new_n283), .A2(new_n285), .ZN(new_n286));
  INV_X1    g100(.A(new_n286), .ZN(new_n287));
  INV_X1    g101(.A(KEYINPUT6), .ZN(new_n288));
  NAND4_X1  g102(.A1(new_n251), .A2(new_n288), .A3(new_n255), .A4(new_n257), .ZN(new_n289));
  NAND3_X1  g103(.A1(new_n261), .A2(new_n287), .A3(new_n289), .ZN(new_n290));
  INV_X1    g104(.A(KEYINPUT86), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n290), .A2(new_n291), .ZN(new_n292));
  NAND4_X1  g106(.A1(new_n261), .A2(KEYINPUT86), .A3(new_n287), .A4(new_n289), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n292), .A2(new_n293), .ZN(new_n294));
  OAI22_X1  g108(.A1(new_n283), .A2(new_n285), .B1(KEYINPUT7), .B2(new_n282), .ZN(new_n295));
  XOR2_X1   g109(.A(new_n256), .B(KEYINPUT8), .Z(new_n296));
  NAND2_X1  g110(.A1(new_n242), .A2(new_n230), .ZN(new_n297));
  AOI21_X1  g111(.A(new_n296), .B1(new_n238), .B2(new_n297), .ZN(new_n298));
  NAND2_X1  g112(.A1(new_n214), .A2(new_n237), .ZN(new_n299));
  NAND4_X1  g113(.A1(new_n299), .A2(new_n244), .A3(new_n230), .A4(new_n241), .ZN(new_n300));
  NOR2_X1   g114(.A1(new_n282), .A2(KEYINPUT7), .ZN(new_n301));
  AOI22_X1  g115(.A1(new_n298), .A2(new_n300), .B1(new_n280), .B2(new_n301), .ZN(new_n302));
  NAND3_X1  g116(.A1(new_n259), .A2(new_n295), .A3(new_n302), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n303), .A2(new_n189), .ZN(new_n304));
  INV_X1    g118(.A(KEYINPUT87), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n304), .A2(new_n305), .ZN(new_n306));
  NAND3_X1  g120(.A1(new_n303), .A2(KEYINPUT87), .A3(new_n189), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n306), .A2(new_n307), .ZN(new_n308));
  INV_X1    g122(.A(new_n308), .ZN(new_n309));
  AOI21_X1  g123(.A(new_n198), .B1(new_n294), .B2(new_n309), .ZN(new_n310));
  INV_X1    g124(.A(new_n198), .ZN(new_n311));
  AOI211_X1 g125(.A(new_n311), .B(new_n308), .C1(new_n292), .C2(new_n293), .ZN(new_n312));
  OAI211_X1 g126(.A(new_n194), .B(new_n197), .C1(new_n310), .C2(new_n312), .ZN(new_n313));
  INV_X1    g127(.A(G237), .ZN(new_n314));
  NAND3_X1  g128(.A1(new_n314), .A2(new_n190), .A3(G214), .ZN(new_n315));
  XNOR2_X1  g129(.A(new_n315), .B(new_n262), .ZN(new_n316));
  INV_X1    g130(.A(KEYINPUT18), .ZN(new_n317));
  INV_X1    g131(.A(G131), .ZN(new_n318));
  NOR2_X1   g132(.A1(new_n317), .A2(new_n318), .ZN(new_n319));
  XNOR2_X1  g133(.A(G125), .B(G140), .ZN(new_n320));
  OR2_X1    g134(.A1(new_n320), .A2(new_n265), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n320), .A2(new_n265), .ZN(new_n322));
  AOI22_X1  g136(.A1(new_n316), .A2(new_n319), .B1(new_n321), .B2(new_n322), .ZN(new_n323));
  XNOR2_X1  g137(.A(new_n315), .B(G143), .ZN(new_n324));
  OAI21_X1  g138(.A(new_n324), .B1(new_n317), .B2(new_n318), .ZN(new_n325));
  AND2_X1   g139(.A1(new_n325), .A2(KEYINPUT88), .ZN(new_n326));
  NOR2_X1   g140(.A1(new_n325), .A2(KEYINPUT88), .ZN(new_n327));
  OAI21_X1  g141(.A(new_n323), .B1(new_n326), .B2(new_n327), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n320), .A2(KEYINPUT16), .ZN(new_n329));
  OR3_X1    g143(.A1(new_n273), .A2(KEYINPUT16), .A3(G140), .ZN(new_n330));
  NAND3_X1  g144(.A1(new_n329), .A2(G146), .A3(new_n330), .ZN(new_n331));
  INV_X1    g145(.A(new_n331), .ZN(new_n332));
  AOI21_X1  g146(.A(G146), .B1(new_n329), .B2(new_n330), .ZN(new_n333));
  OR3_X1    g147(.A1(new_n332), .A2(KEYINPUT92), .A3(new_n333), .ZN(new_n334));
  OAI21_X1  g148(.A(KEYINPUT92), .B1(new_n332), .B2(new_n333), .ZN(new_n335));
  NAND3_X1  g149(.A1(new_n316), .A2(KEYINPUT17), .A3(G131), .ZN(new_n336));
  NAND3_X1  g150(.A1(new_n334), .A2(new_n335), .A3(new_n336), .ZN(new_n337));
  OAI21_X1  g151(.A(KEYINPUT89), .B1(new_n316), .B2(G131), .ZN(new_n338));
  INV_X1    g152(.A(KEYINPUT89), .ZN(new_n339));
  NAND3_X1  g153(.A1(new_n324), .A2(new_n339), .A3(new_n318), .ZN(new_n340));
  OAI211_X1 g154(.A(new_n338), .B(new_n340), .C1(new_n318), .C2(new_n324), .ZN(new_n341));
  NOR2_X1   g155(.A1(new_n341), .A2(KEYINPUT17), .ZN(new_n342));
  OAI21_X1  g156(.A(new_n328), .B1(new_n337), .B2(new_n342), .ZN(new_n343));
  XNOR2_X1  g157(.A(G113), .B(G122), .ZN(new_n344));
  XNOR2_X1  g158(.A(new_n344), .B(KEYINPUT91), .ZN(new_n345));
  XNOR2_X1  g159(.A(KEYINPUT90), .B(G104), .ZN(new_n346));
  XNOR2_X1  g160(.A(new_n345), .B(new_n346), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n347), .A2(KEYINPUT93), .ZN(new_n348));
  AND2_X1   g162(.A1(new_n343), .A2(new_n348), .ZN(new_n349));
  OAI21_X1  g163(.A(new_n189), .B1(new_n343), .B2(new_n348), .ZN(new_n350));
  OAI21_X1  g164(.A(G475), .B1(new_n349), .B2(new_n350), .ZN(new_n351));
  INV_X1    g165(.A(KEYINPUT20), .ZN(new_n352));
  XOR2_X1   g166(.A(new_n320), .B(KEYINPUT19), .Z(new_n353));
  OR2_X1    g167(.A1(new_n353), .A2(G146), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n331), .A2(KEYINPUT73), .ZN(new_n355));
  INV_X1    g169(.A(KEYINPUT73), .ZN(new_n356));
  NAND4_X1  g170(.A1(new_n329), .A2(new_n356), .A3(G146), .A4(new_n330), .ZN(new_n357));
  NAND4_X1  g171(.A1(new_n341), .A2(new_n354), .A3(new_n355), .A4(new_n357), .ZN(new_n358));
  NAND2_X1  g172(.A1(new_n358), .A2(new_n328), .ZN(new_n359));
  NAND2_X1  g173(.A1(new_n359), .A2(new_n347), .ZN(new_n360));
  INV_X1    g174(.A(new_n347), .ZN(new_n361));
  OAI211_X1 g175(.A(new_n328), .B(new_n361), .C1(new_n337), .C2(new_n342), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n360), .A2(new_n362), .ZN(new_n363));
  NOR2_X1   g177(.A1(G475), .A2(G902), .ZN(new_n364));
  AOI21_X1  g178(.A(new_n352), .B1(new_n363), .B2(new_n364), .ZN(new_n365));
  INV_X1    g179(.A(new_n364), .ZN(new_n366));
  AOI211_X1 g180(.A(KEYINPUT20), .B(new_n366), .C1(new_n360), .C2(new_n362), .ZN(new_n367));
  OAI21_X1  g181(.A(new_n351), .B1(new_n365), .B2(new_n367), .ZN(new_n368));
  INV_X1    g182(.A(new_n368), .ZN(new_n369));
  NOR2_X1   g183(.A1(new_n270), .A2(G143), .ZN(new_n370));
  NOR2_X1   g184(.A1(new_n262), .A2(G128), .ZN(new_n371));
  NOR2_X1   g185(.A1(new_n370), .A2(new_n371), .ZN(new_n372));
  INV_X1    g186(.A(G134), .ZN(new_n373));
  XNOR2_X1  g187(.A(new_n372), .B(new_n373), .ZN(new_n374));
  XNOR2_X1  g188(.A(G116), .B(G122), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n375), .A2(new_n202), .ZN(new_n376));
  NAND3_X1  g190(.A1(new_n218), .A2(KEYINPUT14), .A3(G122), .ZN(new_n377));
  INV_X1    g191(.A(new_n375), .ZN(new_n378));
  OAI211_X1 g192(.A(G107), .B(new_n377), .C1(new_n378), .C2(KEYINPUT14), .ZN(new_n379));
  NAND3_X1  g193(.A1(new_n374), .A2(new_n376), .A3(new_n379), .ZN(new_n380));
  NOR2_X1   g194(.A1(new_n370), .A2(KEYINPUT13), .ZN(new_n381));
  NOR2_X1   g195(.A1(new_n381), .A2(new_n371), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n370), .A2(KEYINPUT13), .ZN(new_n383));
  AOI21_X1  g197(.A(new_n373), .B1(new_n382), .B2(new_n383), .ZN(new_n384));
  XNOR2_X1  g198(.A(new_n375), .B(new_n202), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n372), .A2(new_n373), .ZN(new_n386));
  NAND2_X1  g200(.A1(new_n385), .A2(new_n386), .ZN(new_n387));
  OAI21_X1  g201(.A(new_n380), .B1(new_n384), .B2(new_n387), .ZN(new_n388));
  XNOR2_X1  g202(.A(KEYINPUT9), .B(G234), .ZN(new_n389));
  INV_X1    g203(.A(G217), .ZN(new_n390));
  NOR3_X1   g204(.A1(new_n389), .A2(new_n390), .A3(G953), .ZN(new_n391));
  INV_X1    g205(.A(new_n391), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n388), .A2(new_n392), .ZN(new_n393));
  OAI211_X1 g207(.A(new_n380), .B(new_n391), .C1(new_n384), .C2(new_n387), .ZN(new_n394));
  NAND3_X1  g208(.A1(new_n393), .A2(KEYINPUT94), .A3(new_n394), .ZN(new_n395));
  INV_X1    g209(.A(KEYINPUT94), .ZN(new_n396));
  NAND3_X1  g210(.A1(new_n388), .A2(new_n396), .A3(new_n392), .ZN(new_n397));
  NAND3_X1  g211(.A1(new_n395), .A2(new_n189), .A3(new_n397), .ZN(new_n398));
  INV_X1    g212(.A(G478), .ZN(new_n399));
  NOR2_X1   g213(.A1(new_n399), .A2(KEYINPUT15), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n398), .A2(new_n400), .ZN(new_n401));
  INV_X1    g215(.A(new_n400), .ZN(new_n402));
  NAND4_X1  g216(.A1(new_n395), .A2(new_n189), .A3(new_n397), .A4(new_n402), .ZN(new_n403));
  AND3_X1   g217(.A1(new_n401), .A2(KEYINPUT95), .A3(new_n403), .ZN(new_n404));
  AOI21_X1  g218(.A(KEYINPUT95), .B1(new_n401), .B2(new_n403), .ZN(new_n405));
  NOR2_X1   g219(.A1(new_n404), .A2(new_n405), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n369), .A2(new_n406), .ZN(new_n407));
  NOR2_X1   g221(.A1(new_n313), .A2(new_n407), .ZN(new_n408));
  INV_X1    g222(.A(KEYINPUT25), .ZN(new_n409));
  XNOR2_X1  g223(.A(KEYINPUT24), .B(G110), .ZN(new_n410));
  INV_X1    g224(.A(KEYINPUT72), .ZN(new_n411));
  OR2_X1    g225(.A1(new_n410), .A2(new_n411), .ZN(new_n412));
  XNOR2_X1  g226(.A(G119), .B(G128), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n410), .A2(new_n411), .ZN(new_n414));
  NAND3_X1  g228(.A1(new_n412), .A2(new_n413), .A3(new_n414), .ZN(new_n415));
  INV_X1    g229(.A(KEYINPUT23), .ZN(new_n416));
  OAI21_X1  g230(.A(new_n416), .B1(new_n216), .B2(G128), .ZN(new_n417));
  NAND3_X1  g231(.A1(new_n270), .A2(KEYINPUT23), .A3(G119), .ZN(new_n418));
  OAI211_X1 g232(.A(new_n417), .B(new_n418), .C1(G119), .C2(new_n270), .ZN(new_n419));
  NAND2_X1  g233(.A1(new_n419), .A2(G110), .ZN(new_n420));
  OAI211_X1 g234(.A(new_n415), .B(new_n420), .C1(new_n332), .C2(new_n333), .ZN(new_n421));
  AOI21_X1  g235(.A(new_n413), .B1(new_n412), .B2(new_n414), .ZN(new_n422));
  NOR2_X1   g236(.A1(new_n419), .A2(G110), .ZN(new_n423));
  OAI21_X1  g237(.A(new_n322), .B1(new_n422), .B2(new_n423), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n355), .A2(new_n357), .ZN(new_n425));
  OAI21_X1  g239(.A(new_n421), .B1(new_n424), .B2(new_n425), .ZN(new_n426));
  XNOR2_X1  g240(.A(KEYINPUT22), .B(G137), .ZN(new_n427));
  NAND3_X1  g241(.A1(new_n190), .A2(G221), .A3(G234), .ZN(new_n428));
  XNOR2_X1  g242(.A(new_n427), .B(new_n428), .ZN(new_n429));
  INV_X1    g243(.A(new_n429), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n426), .A2(new_n430), .ZN(new_n431));
  OAI211_X1 g245(.A(new_n421), .B(new_n429), .C1(new_n424), .C2(new_n425), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n431), .A2(new_n432), .ZN(new_n433));
  OAI21_X1  g247(.A(new_n409), .B1(new_n433), .B2(G902), .ZN(new_n434));
  NAND4_X1  g248(.A1(new_n431), .A2(KEYINPUT25), .A3(new_n189), .A4(new_n432), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n434), .A2(new_n435), .ZN(new_n436));
  AOI21_X1  g250(.A(new_n390), .B1(G234), .B2(new_n189), .ZN(new_n437));
  NAND3_X1  g251(.A1(new_n436), .A2(KEYINPUT74), .A3(new_n437), .ZN(new_n438));
  INV_X1    g252(.A(new_n438), .ZN(new_n439));
  AOI21_X1  g253(.A(KEYINPUT74), .B1(new_n436), .B2(new_n437), .ZN(new_n440));
  NOR3_X1   g254(.A1(new_n433), .A2(G902), .A3(new_n437), .ZN(new_n441));
  NOR3_X1   g255(.A1(new_n439), .A2(new_n440), .A3(new_n441), .ZN(new_n442));
  INV_X1    g256(.A(new_n442), .ZN(new_n443));
  NOR2_X1   g257(.A1(G472), .A2(G902), .ZN(new_n444));
  INV_X1    g258(.A(KEYINPUT30), .ZN(new_n445));
  INV_X1    g259(.A(G137), .ZN(new_n446));
  NAND3_X1  g260(.A1(new_n446), .A2(KEYINPUT11), .A3(G134), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n373), .A2(G137), .ZN(new_n448));
  AND2_X1   g262(.A1(new_n447), .A2(new_n448), .ZN(new_n449));
  INV_X1    g263(.A(KEYINPUT64), .ZN(new_n450));
  INV_X1    g264(.A(KEYINPUT11), .ZN(new_n451));
  OAI21_X1  g265(.A(new_n451), .B1(new_n373), .B2(G137), .ZN(new_n452));
  NAND4_X1  g266(.A1(new_n449), .A2(new_n450), .A3(new_n318), .A4(new_n452), .ZN(new_n453));
  NAND4_X1  g267(.A1(new_n452), .A2(new_n447), .A3(new_n318), .A4(new_n448), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n454), .A2(KEYINPUT64), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n453), .A2(new_n455), .ZN(new_n456));
  INV_X1    g270(.A(KEYINPUT66), .ZN(new_n457));
  NOR2_X1   g271(.A1(new_n373), .A2(G137), .ZN(new_n458));
  NOR2_X1   g272(.A1(new_n446), .A2(G134), .ZN(new_n459));
  OAI21_X1  g273(.A(G131), .B1(new_n458), .B2(new_n459), .ZN(new_n460));
  AND3_X1   g274(.A1(new_n267), .A2(new_n460), .A3(new_n271), .ZN(new_n461));
  NAND3_X1  g275(.A1(new_n456), .A2(new_n457), .A3(new_n461), .ZN(new_n462));
  NAND3_X1  g276(.A1(new_n452), .A2(new_n447), .A3(new_n448), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n463), .A2(KEYINPUT65), .ZN(new_n464));
  INV_X1    g278(.A(KEYINPUT65), .ZN(new_n465));
  NAND4_X1  g279(.A1(new_n452), .A2(new_n447), .A3(new_n465), .A4(new_n448), .ZN(new_n466));
  AND2_X1   g280(.A1(new_n466), .A2(G131), .ZN(new_n467));
  AOI22_X1  g281(.A1(new_n464), .A2(new_n467), .B1(new_n453), .B2(new_n455), .ZN(new_n468));
  OAI21_X1  g282(.A(new_n462), .B1(new_n468), .B2(new_n278), .ZN(new_n469));
  NAND3_X1  g283(.A1(new_n267), .A2(new_n460), .A3(new_n271), .ZN(new_n470));
  AOI21_X1  g284(.A(new_n470), .B1(new_n453), .B2(new_n455), .ZN(new_n471));
  NOR2_X1   g285(.A1(new_n471), .A2(new_n457), .ZN(new_n472));
  OAI21_X1  g286(.A(new_n445), .B1(new_n469), .B2(new_n472), .ZN(new_n473));
  NAND3_X1  g287(.A1(new_n464), .A2(G131), .A3(new_n466), .ZN(new_n474));
  AOI21_X1  g288(.A(new_n278), .B1(new_n456), .B2(new_n474), .ZN(new_n475));
  NOR2_X1   g289(.A1(new_n475), .A2(new_n471), .ZN(new_n476));
  NAND2_X1  g290(.A1(new_n476), .A2(KEYINPUT30), .ZN(new_n477));
  NAND3_X1  g291(.A1(new_n473), .A2(new_n231), .A3(new_n477), .ZN(new_n478));
  XOR2_X1   g292(.A(KEYINPUT26), .B(G101), .Z(new_n479));
  NAND3_X1  g293(.A1(new_n314), .A2(new_n190), .A3(G210), .ZN(new_n480));
  XNOR2_X1  g294(.A(new_n479), .B(new_n480), .ZN(new_n481));
  XNOR2_X1  g295(.A(KEYINPUT69), .B(KEYINPUT27), .ZN(new_n482));
  XNOR2_X1  g296(.A(new_n481), .B(new_n482), .ZN(new_n483));
  INV_X1    g297(.A(KEYINPUT68), .ZN(new_n484));
  NAND2_X1  g298(.A1(new_n231), .A2(new_n484), .ZN(new_n485));
  NAND3_X1  g299(.A1(new_n227), .A2(new_n230), .A3(KEYINPUT68), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n485), .A2(new_n486), .ZN(new_n487));
  AOI21_X1  g301(.A(new_n483), .B1(new_n476), .B2(new_n487), .ZN(new_n488));
  AND3_X1   g302(.A1(new_n478), .A2(KEYINPUT70), .A3(new_n488), .ZN(new_n489));
  AOI21_X1  g303(.A(KEYINPUT70), .B1(new_n478), .B2(new_n488), .ZN(new_n490));
  INV_X1    g304(.A(KEYINPUT31), .ZN(new_n491));
  NOR3_X1   g305(.A1(new_n489), .A2(new_n490), .A3(new_n491), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n476), .A2(new_n487), .ZN(new_n493));
  INV_X1    g307(.A(new_n483), .ZN(new_n494));
  NAND2_X1  g308(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  NOR3_X1   g309(.A1(new_n475), .A2(new_n445), .A3(new_n471), .ZN(new_n496));
  AND2_X1   g310(.A1(new_n454), .A2(KEYINPUT64), .ZN(new_n497));
  NOR2_X1   g311(.A1(new_n454), .A2(KEYINPUT64), .ZN(new_n498));
  AOI21_X1  g312(.A(new_n465), .B1(new_n449), .B2(new_n452), .ZN(new_n499));
  NAND2_X1  g313(.A1(new_n466), .A2(G131), .ZN(new_n500));
  OAI22_X1  g314(.A1(new_n497), .A2(new_n498), .B1(new_n499), .B2(new_n500), .ZN(new_n501));
  INV_X1    g315(.A(new_n278), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  XNOR2_X1  g317(.A(new_n454), .B(new_n450), .ZN(new_n504));
  OAI21_X1  g318(.A(KEYINPUT66), .B1(new_n504), .B2(new_n470), .ZN(new_n505));
  NAND3_X1  g319(.A1(new_n503), .A2(new_n505), .A3(new_n462), .ZN(new_n506));
  AOI21_X1  g320(.A(new_n496), .B1(new_n445), .B2(new_n506), .ZN(new_n507));
  AOI21_X1  g321(.A(new_n495), .B1(new_n507), .B2(new_n231), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n508), .A2(new_n491), .ZN(new_n509));
  INV_X1    g323(.A(KEYINPUT28), .ZN(new_n510));
  NAND2_X1  g324(.A1(new_n493), .A2(new_n510), .ZN(new_n511));
  AOI22_X1  g325(.A1(new_n506), .A2(new_n231), .B1(new_n476), .B2(new_n487), .ZN(new_n512));
  OAI21_X1  g326(.A(new_n511), .B1(new_n512), .B2(new_n510), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n513), .A2(new_n483), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n509), .A2(new_n514), .ZN(new_n515));
  OAI21_X1  g329(.A(new_n444), .B1(new_n492), .B2(new_n515), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n516), .A2(KEYINPUT32), .ZN(new_n517));
  INV_X1    g331(.A(new_n444), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n478), .A2(new_n488), .ZN(new_n519));
  INV_X1    g333(.A(KEYINPUT70), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  NAND3_X1  g335(.A1(new_n478), .A2(KEYINPUT70), .A3(new_n488), .ZN(new_n522));
  NAND3_X1  g336(.A1(new_n521), .A2(KEYINPUT31), .A3(new_n522), .ZN(new_n523));
  AOI22_X1  g337(.A1(new_n491), .A2(new_n508), .B1(new_n513), .B2(new_n483), .ZN(new_n524));
  AOI21_X1  g338(.A(new_n518), .B1(new_n523), .B2(new_n524), .ZN(new_n525));
  INV_X1    g339(.A(KEYINPUT32), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n517), .A2(new_n527), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n478), .A2(new_n493), .ZN(new_n529));
  NAND2_X1  g343(.A1(new_n529), .A2(new_n483), .ZN(new_n530));
  INV_X1    g344(.A(KEYINPUT29), .ZN(new_n531));
  OAI211_X1 g345(.A(new_n530), .B(new_n531), .C1(new_n483), .C2(new_n513), .ZN(new_n532));
  INV_X1    g346(.A(new_n487), .ZN(new_n533));
  OAI22_X1  g347(.A1(new_n468), .A2(new_n278), .B1(new_n504), .B2(new_n470), .ZN(new_n534));
  NAND2_X1  g348(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  AOI21_X1  g349(.A(new_n510), .B1(new_n535), .B2(new_n493), .ZN(new_n536));
  NOR2_X1   g350(.A1(new_n533), .A2(new_n534), .ZN(new_n537));
  NOR2_X1   g351(.A1(new_n537), .A2(KEYINPUT28), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n494), .A2(KEYINPUT29), .ZN(new_n539));
  NOR3_X1   g353(.A1(new_n536), .A2(new_n538), .A3(new_n539), .ZN(new_n540));
  OAI21_X1  g354(.A(KEYINPUT71), .B1(new_n540), .B2(G902), .ZN(new_n541));
  INV_X1    g355(.A(KEYINPUT71), .ZN(new_n542));
  NOR2_X1   g356(.A1(new_n476), .A2(new_n487), .ZN(new_n543));
  OAI21_X1  g357(.A(KEYINPUT28), .B1(new_n537), .B2(new_n543), .ZN(new_n544));
  NAND2_X1  g358(.A1(new_n544), .A2(new_n511), .ZN(new_n545));
  OAI211_X1 g359(.A(new_n542), .B(new_n189), .C1(new_n545), .C2(new_n539), .ZN(new_n546));
  NAND3_X1  g360(.A1(new_n532), .A2(new_n541), .A3(new_n546), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n547), .A2(G472), .ZN(new_n548));
  AOI21_X1  g362(.A(new_n443), .B1(new_n528), .B2(new_n548), .ZN(new_n549));
  OAI21_X1  g363(.A(G221), .B1(new_n389), .B2(G902), .ZN(new_n550));
  INV_X1    g364(.A(new_n550), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n214), .A2(KEYINPUT4), .ZN(new_n552));
  OAI211_X1 g366(.A(new_n502), .B(new_n234), .C1(new_n552), .C2(new_n248), .ZN(new_n553));
  XNOR2_X1  g367(.A(KEYINPUT76), .B(KEYINPUT10), .ZN(new_n554));
  OAI21_X1  g368(.A(new_n554), .B1(new_n299), .B2(new_n272), .ZN(new_n555));
  INV_X1    g369(.A(new_n272), .ZN(new_n556));
  NAND4_X1  g370(.A1(new_n556), .A2(KEYINPUT10), .A3(new_n214), .A4(new_n237), .ZN(new_n557));
  AND3_X1   g371(.A1(new_n553), .A2(new_n555), .A3(new_n557), .ZN(new_n558));
  INV_X1    g372(.A(KEYINPUT12), .ZN(new_n559));
  OAI21_X1  g373(.A(new_n559), .B1(new_n468), .B2(KEYINPUT77), .ZN(new_n560));
  NOR2_X1   g374(.A1(new_n299), .A2(new_n272), .ZN(new_n561));
  AOI22_X1  g375(.A1(new_n214), .A2(new_n237), .B1(new_n271), .B2(new_n267), .ZN(new_n562));
  OAI21_X1  g376(.A(new_n501), .B1(new_n561), .B2(new_n562), .ZN(new_n563));
  AOI22_X1  g377(.A1(new_n558), .A2(new_n468), .B1(new_n560), .B2(new_n563), .ZN(new_n564));
  XNOR2_X1  g378(.A(G110), .B(G140), .ZN(new_n565));
  INV_X1    g379(.A(G227), .ZN(new_n566));
  NOR2_X1   g380(.A1(new_n566), .A2(G953), .ZN(new_n567));
  XNOR2_X1  g381(.A(new_n565), .B(new_n567), .ZN(new_n568));
  INV_X1    g382(.A(new_n568), .ZN(new_n569));
  NAND3_X1  g383(.A1(new_n556), .A2(new_n214), .A3(new_n237), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n299), .A2(new_n272), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n570), .A2(new_n571), .ZN(new_n572));
  NAND4_X1  g386(.A1(new_n572), .A2(KEYINPUT77), .A3(new_n559), .A4(new_n501), .ZN(new_n573));
  NAND4_X1  g387(.A1(new_n564), .A2(KEYINPUT79), .A3(new_n569), .A4(new_n573), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n560), .A2(new_n563), .ZN(new_n575));
  NAND4_X1  g389(.A1(new_n553), .A2(new_n555), .A3(new_n468), .A4(new_n557), .ZN(new_n576));
  NAND4_X1  g390(.A1(new_n575), .A2(new_n573), .A3(new_n569), .A4(new_n576), .ZN(new_n577));
  INV_X1    g391(.A(KEYINPUT79), .ZN(new_n578));
  NAND2_X1  g392(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n574), .A2(new_n579), .ZN(new_n580));
  NAND3_X1  g394(.A1(new_n553), .A2(new_n555), .A3(new_n557), .ZN(new_n581));
  NAND2_X1  g395(.A1(new_n581), .A2(new_n501), .ZN(new_n582));
  NAND3_X1  g396(.A1(new_n582), .A2(KEYINPUT78), .A3(new_n576), .ZN(new_n583));
  INV_X1    g397(.A(KEYINPUT78), .ZN(new_n584));
  NAND3_X1  g398(.A1(new_n581), .A2(new_n584), .A3(new_n501), .ZN(new_n585));
  NAND3_X1  g399(.A1(new_n583), .A2(new_n568), .A3(new_n585), .ZN(new_n586));
  INV_X1    g400(.A(KEYINPUT80), .ZN(new_n587));
  NAND2_X1  g401(.A1(new_n586), .A2(new_n587), .ZN(new_n588));
  NAND4_X1  g402(.A1(new_n583), .A2(KEYINPUT80), .A3(new_n568), .A4(new_n585), .ZN(new_n589));
  NAND3_X1  g403(.A1(new_n580), .A2(new_n588), .A3(new_n589), .ZN(new_n590));
  INV_X1    g404(.A(G469), .ZN(new_n591));
  NAND3_X1  g405(.A1(new_n590), .A2(new_n591), .A3(new_n189), .ZN(new_n592));
  NAND3_X1  g406(.A1(new_n575), .A2(new_n573), .A3(new_n576), .ZN(new_n593));
  NAND2_X1  g407(.A1(new_n593), .A2(new_n568), .ZN(new_n594));
  INV_X1    g408(.A(new_n594), .ZN(new_n595));
  AOI21_X1  g409(.A(new_n568), .B1(new_n583), .B2(new_n585), .ZN(new_n596));
  NOR2_X1   g410(.A1(new_n595), .A2(new_n596), .ZN(new_n597));
  OAI21_X1  g411(.A(G469), .B1(new_n597), .B2(G902), .ZN(new_n598));
  AOI21_X1  g412(.A(new_n551), .B1(new_n592), .B2(new_n598), .ZN(new_n599));
  XNOR2_X1  g413(.A(new_n599), .B(KEYINPUT81), .ZN(new_n600));
  NAND3_X1  g414(.A1(new_n408), .A2(new_n549), .A3(new_n600), .ZN(new_n601));
  XNOR2_X1  g415(.A(new_n601), .B(G101), .ZN(G3));
  AOI21_X1  g416(.A(G902), .B1(new_n523), .B2(new_n524), .ZN(new_n603));
  INV_X1    g417(.A(G472), .ZN(new_n604));
  NOR2_X1   g418(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  NOR2_X1   g419(.A1(new_n605), .A2(new_n525), .ZN(new_n606));
  AND3_X1   g420(.A1(new_n600), .A2(new_n442), .A3(new_n606), .ZN(new_n607));
  INV_X1    g421(.A(KEYINPUT33), .ZN(new_n608));
  NAND3_X1  g422(.A1(new_n395), .A2(new_n608), .A3(new_n397), .ZN(new_n609));
  NAND3_X1  g423(.A1(new_n393), .A2(KEYINPUT33), .A3(new_n394), .ZN(new_n610));
  AND2_X1   g424(.A1(new_n609), .A2(new_n610), .ZN(new_n611));
  NAND3_X1  g425(.A1(new_n611), .A2(G478), .A3(new_n189), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n398), .A2(new_n399), .ZN(new_n613));
  NAND2_X1  g427(.A1(new_n612), .A2(new_n613), .ZN(new_n614));
  INV_X1    g428(.A(new_n614), .ZN(new_n615));
  NOR3_X1   g429(.A1(new_n313), .A2(new_n369), .A3(new_n615), .ZN(new_n616));
  NAND2_X1  g430(.A1(new_n607), .A2(new_n616), .ZN(new_n617));
  XOR2_X1   g431(.A(KEYINPUT34), .B(G104), .Z(new_n618));
  XNOR2_X1  g432(.A(new_n617), .B(new_n618), .ZN(G6));
  NOR2_X1   g433(.A1(new_n406), .A2(new_n368), .ZN(new_n620));
  INV_X1    g434(.A(new_n620), .ZN(new_n621));
  NOR2_X1   g435(.A1(new_n313), .A2(new_n621), .ZN(new_n622));
  NAND2_X1  g436(.A1(new_n607), .A2(new_n622), .ZN(new_n623));
  XNOR2_X1  g437(.A(KEYINPUT97), .B(G107), .ZN(new_n624));
  XNOR2_X1  g438(.A(new_n623), .B(new_n624), .ZN(new_n625));
  XNOR2_X1  g439(.A(KEYINPUT96), .B(KEYINPUT35), .ZN(new_n626));
  XNOR2_X1  g440(.A(new_n625), .B(new_n626), .ZN(G9));
  NAND2_X1  g441(.A1(new_n436), .A2(new_n437), .ZN(new_n628));
  INV_X1    g442(.A(KEYINPUT74), .ZN(new_n629));
  NAND2_X1  g443(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  NOR2_X1   g444(.A1(new_n430), .A2(KEYINPUT36), .ZN(new_n631));
  XOR2_X1   g445(.A(new_n631), .B(KEYINPUT98), .Z(new_n632));
  XNOR2_X1  g446(.A(new_n632), .B(new_n426), .ZN(new_n633));
  OR3_X1    g447(.A1(new_n633), .A2(G902), .A3(new_n437), .ZN(new_n634));
  NAND3_X1  g448(.A1(new_n630), .A2(new_n634), .A3(new_n438), .ZN(new_n635));
  OAI211_X1 g449(.A(new_n635), .B(new_n516), .C1(new_n604), .C2(new_n603), .ZN(new_n636));
  INV_X1    g450(.A(KEYINPUT99), .ZN(new_n637));
  XNOR2_X1  g451(.A(new_n636), .B(new_n637), .ZN(new_n638));
  NAND3_X1  g452(.A1(new_n638), .A2(new_n408), .A3(new_n600), .ZN(new_n639));
  XNOR2_X1  g453(.A(KEYINPUT37), .B(G110), .ZN(new_n640));
  XNOR2_X1  g454(.A(new_n640), .B(KEYINPUT100), .ZN(new_n641));
  XNOR2_X1  g455(.A(new_n639), .B(new_n641), .ZN(G12));
  INV_X1    g456(.A(KEYINPUT101), .ZN(new_n643));
  NAND2_X1  g457(.A1(new_n523), .A2(new_n524), .ZN(new_n644));
  AOI21_X1  g458(.A(new_n526), .B1(new_n644), .B2(new_n444), .ZN(new_n645));
  AOI211_X1 g459(.A(KEYINPUT32), .B(new_n518), .C1(new_n523), .C2(new_n524), .ZN(new_n646));
  OAI21_X1  g460(.A(new_n548), .B1(new_n645), .B2(new_n646), .ZN(new_n647));
  NAND2_X1  g461(.A1(new_n592), .A2(new_n598), .ZN(new_n648));
  AOI21_X1  g462(.A(KEYINPUT81), .B1(new_n648), .B2(new_n550), .ZN(new_n649));
  INV_X1    g463(.A(KEYINPUT81), .ZN(new_n650));
  AOI211_X1 g464(.A(new_n650), .B(new_n551), .C1(new_n592), .C2(new_n598), .ZN(new_n651));
  OAI211_X1 g465(.A(new_n647), .B(new_n635), .C1(new_n649), .C2(new_n651), .ZN(new_n652));
  INV_X1    g466(.A(G900), .ZN(new_n653));
  NAND2_X1  g467(.A1(new_n191), .A2(new_n653), .ZN(new_n654));
  INV_X1    g468(.A(new_n188), .ZN(new_n655));
  NAND2_X1  g469(.A1(new_n654), .A2(new_n655), .ZN(new_n656));
  INV_X1    g470(.A(new_n656), .ZN(new_n657));
  NOR3_X1   g471(.A1(new_n406), .A2(new_n368), .A3(new_n657), .ZN(new_n658));
  OAI211_X1 g472(.A(new_n658), .B(new_n197), .C1(new_n310), .C2(new_n312), .ZN(new_n659));
  OAI21_X1  g473(.A(new_n643), .B1(new_n652), .B2(new_n659), .ZN(new_n660));
  INV_X1    g474(.A(new_n659), .ZN(new_n661));
  INV_X1    g475(.A(new_n635), .ZN(new_n662));
  AOI21_X1  g476(.A(new_n662), .B1(new_n528), .B2(new_n548), .ZN(new_n663));
  NAND4_X1  g477(.A1(new_n661), .A2(new_n600), .A3(new_n663), .A4(KEYINPUT101), .ZN(new_n664));
  NAND2_X1  g478(.A1(new_n660), .A2(new_n664), .ZN(new_n665));
  XNOR2_X1  g479(.A(new_n665), .B(G128), .ZN(G30));
  NAND2_X1  g480(.A1(new_n294), .A2(new_n309), .ZN(new_n667));
  NAND2_X1  g481(.A1(new_n667), .A2(new_n311), .ZN(new_n668));
  NAND3_X1  g482(.A1(new_n294), .A2(new_n198), .A3(new_n309), .ZN(new_n669));
  NAND2_X1  g483(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  XOR2_X1   g484(.A(new_n670), .B(KEYINPUT38), .Z(new_n671));
  NOR2_X1   g485(.A1(new_n489), .A2(new_n490), .ZN(new_n672));
  OAI21_X1  g486(.A(new_n483), .B1(new_n537), .B2(new_n543), .ZN(new_n673));
  NAND2_X1  g487(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  AOI21_X1  g488(.A(new_n604), .B1(new_n674), .B2(new_n189), .ZN(new_n675));
  AOI21_X1  g489(.A(new_n675), .B1(new_n517), .B2(new_n527), .ZN(new_n676));
  NOR2_X1   g490(.A1(new_n369), .A2(new_n406), .ZN(new_n677));
  NAND3_X1  g491(.A1(new_n677), .A2(new_n662), .A3(new_n197), .ZN(new_n678));
  NOR3_X1   g492(.A1(new_n671), .A2(new_n676), .A3(new_n678), .ZN(new_n679));
  XNOR2_X1  g493(.A(new_n656), .B(KEYINPUT39), .ZN(new_n680));
  NAND2_X1  g494(.A1(new_n600), .A2(new_n680), .ZN(new_n681));
  OR2_X1    g495(.A1(new_n681), .A2(KEYINPUT40), .ZN(new_n682));
  NAND2_X1  g496(.A1(new_n681), .A2(KEYINPUT40), .ZN(new_n683));
  NAND3_X1  g497(.A1(new_n679), .A2(new_n682), .A3(new_n683), .ZN(new_n684));
  XNOR2_X1  g498(.A(new_n684), .B(G143), .ZN(G45));
  INV_X1    g499(.A(new_n652), .ZN(new_n686));
  AND3_X1   g500(.A1(new_n614), .A2(new_n368), .A3(new_n656), .ZN(new_n687));
  OAI211_X1 g501(.A(new_n197), .B(new_n687), .C1(new_n310), .C2(new_n312), .ZN(new_n688));
  INV_X1    g502(.A(KEYINPUT102), .ZN(new_n689));
  NAND2_X1  g503(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  AOI21_X1  g504(.A(new_n196), .B1(new_n668), .B2(new_n669), .ZN(new_n691));
  NAND3_X1  g505(.A1(new_n691), .A2(KEYINPUT102), .A3(new_n687), .ZN(new_n692));
  NAND3_X1  g506(.A1(new_n686), .A2(new_n690), .A3(new_n692), .ZN(new_n693));
  XNOR2_X1  g507(.A(new_n693), .B(G146), .ZN(G48));
  NAND2_X1  g508(.A1(new_n590), .A2(new_n189), .ZN(new_n695));
  NAND2_X1  g509(.A1(new_n695), .A2(G469), .ZN(new_n696));
  AND3_X1   g510(.A1(new_n696), .A2(new_n550), .A3(new_n592), .ZN(new_n697));
  AND3_X1   g511(.A1(new_n647), .A2(new_n697), .A3(new_n442), .ZN(new_n698));
  NAND2_X1  g512(.A1(new_n616), .A2(new_n698), .ZN(new_n699));
  XNOR2_X1  g513(.A(KEYINPUT41), .B(G113), .ZN(new_n700));
  XNOR2_X1  g514(.A(new_n699), .B(new_n700), .ZN(G15));
  INV_X1    g515(.A(KEYINPUT103), .ZN(new_n702));
  NAND4_X1  g516(.A1(new_n670), .A2(new_n194), .A3(new_n197), .A4(new_n620), .ZN(new_n703));
  NAND3_X1  g517(.A1(new_n647), .A2(new_n697), .A3(new_n442), .ZN(new_n704));
  OAI21_X1  g518(.A(new_n702), .B1(new_n703), .B2(new_n704), .ZN(new_n705));
  NAND3_X1  g519(.A1(new_n622), .A2(new_n698), .A3(KEYINPUT103), .ZN(new_n706));
  NAND2_X1  g520(.A1(new_n705), .A2(new_n706), .ZN(new_n707));
  XNOR2_X1  g521(.A(KEYINPUT104), .B(G116), .ZN(new_n708));
  XNOR2_X1  g522(.A(new_n707), .B(new_n708), .ZN(G18));
  NOR2_X1   g523(.A1(new_n407), .A2(new_n193), .ZN(new_n710));
  AND3_X1   g524(.A1(new_n647), .A2(new_n635), .A3(new_n710), .ZN(new_n711));
  OAI21_X1  g525(.A(new_n197), .B1(new_n310), .B2(new_n312), .ZN(new_n712));
  NAND3_X1  g526(.A1(new_n696), .A2(new_n550), .A3(new_n592), .ZN(new_n713));
  NOR2_X1   g527(.A1(new_n712), .A2(new_n713), .ZN(new_n714));
  NAND2_X1  g528(.A1(new_n711), .A2(new_n714), .ZN(new_n715));
  XOR2_X1   g529(.A(KEYINPUT105), .B(G119), .Z(new_n716));
  XNOR2_X1  g530(.A(new_n715), .B(new_n716), .ZN(G21));
  INV_X1    g531(.A(KEYINPUT106), .ZN(new_n718));
  OAI21_X1  g532(.A(new_n718), .B1(new_n536), .B2(new_n538), .ZN(new_n719));
  NAND3_X1  g533(.A1(new_n544), .A2(KEYINPUT106), .A3(new_n511), .ZN(new_n720));
  NAND3_X1  g534(.A1(new_n719), .A2(new_n720), .A3(new_n483), .ZN(new_n721));
  NAND3_X1  g535(.A1(new_n523), .A2(new_n721), .A3(KEYINPUT107), .ZN(new_n722));
  NAND2_X1  g536(.A1(new_n722), .A2(new_n509), .ZN(new_n723));
  AOI21_X1  g537(.A(KEYINPUT107), .B1(new_n523), .B2(new_n721), .ZN(new_n724));
  OAI21_X1  g538(.A(new_n444), .B1(new_n723), .B2(new_n724), .ZN(new_n725));
  INV_X1    g539(.A(new_n605), .ZN(new_n726));
  NAND3_X1  g540(.A1(new_n725), .A2(new_n442), .A3(new_n726), .ZN(new_n727));
  NAND2_X1  g541(.A1(new_n727), .A2(KEYINPUT108), .ZN(new_n728));
  INV_X1    g542(.A(KEYINPUT108), .ZN(new_n729));
  NAND4_X1  g543(.A1(new_n725), .A2(new_n726), .A3(new_n729), .A4(new_n442), .ZN(new_n730));
  NAND2_X1  g544(.A1(new_n728), .A2(new_n730), .ZN(new_n731));
  OAI211_X1 g545(.A(new_n677), .B(new_n197), .C1(new_n310), .C2(new_n312), .ZN(new_n732));
  NOR3_X1   g546(.A1(new_n732), .A2(new_n193), .A3(new_n713), .ZN(new_n733));
  NAND2_X1  g547(.A1(new_n731), .A2(new_n733), .ZN(new_n734));
  NAND2_X1  g548(.A1(new_n734), .A2(KEYINPUT109), .ZN(new_n735));
  INV_X1    g549(.A(KEYINPUT109), .ZN(new_n736));
  NAND3_X1  g550(.A1(new_n731), .A2(new_n736), .A3(new_n733), .ZN(new_n737));
  NAND2_X1  g551(.A1(new_n735), .A2(new_n737), .ZN(new_n738));
  XNOR2_X1  g552(.A(new_n738), .B(G122), .ZN(G24));
  NAND4_X1  g553(.A1(new_n725), .A2(new_n726), .A3(new_n635), .A4(new_n687), .ZN(new_n740));
  NOR3_X1   g554(.A1(new_n740), .A2(new_n712), .A3(new_n713), .ZN(new_n741));
  XNOR2_X1  g555(.A(new_n741), .B(new_n273), .ZN(G27));
  INV_X1    g556(.A(KEYINPUT42), .ZN(new_n743));
  NOR2_X1   g557(.A1(new_n594), .A2(KEYINPUT110), .ZN(new_n744));
  INV_X1    g558(.A(KEYINPUT110), .ZN(new_n745));
  AOI21_X1  g559(.A(new_n745), .B1(new_n593), .B2(new_n568), .ZN(new_n746));
  NOR3_X1   g560(.A1(new_n744), .A2(new_n596), .A3(new_n746), .ZN(new_n747));
  OAI21_X1  g561(.A(G469), .B1(new_n747), .B2(G902), .ZN(new_n748));
  AOI211_X1 g562(.A(KEYINPUT111), .B(new_n551), .C1(new_n748), .C2(new_n592), .ZN(new_n749));
  INV_X1    g563(.A(new_n749), .ZN(new_n750));
  AOI21_X1  g564(.A(new_n551), .B1(new_n748), .B2(new_n592), .ZN(new_n751));
  INV_X1    g565(.A(KEYINPUT111), .ZN(new_n752));
  OR2_X1    g566(.A1(new_n751), .A2(new_n752), .ZN(new_n753));
  NOR3_X1   g567(.A1(new_n310), .A2(new_n312), .A3(new_n196), .ZN(new_n754));
  NAND4_X1  g568(.A1(new_n549), .A2(new_n750), .A3(new_n753), .A4(new_n754), .ZN(new_n755));
  INV_X1    g569(.A(new_n687), .ZN(new_n756));
  OAI21_X1  g570(.A(new_n743), .B1(new_n755), .B2(new_n756), .ZN(new_n757));
  NAND3_X1  g571(.A1(new_n668), .A2(new_n197), .A3(new_n669), .ZN(new_n758));
  NOR2_X1   g572(.A1(new_n751), .A2(new_n752), .ZN(new_n759));
  NOR3_X1   g573(.A1(new_n758), .A2(new_n759), .A3(new_n749), .ZN(new_n760));
  NAND4_X1  g574(.A1(new_n760), .A2(KEYINPUT42), .A3(new_n549), .A4(new_n687), .ZN(new_n761));
  NAND2_X1  g575(.A1(new_n757), .A2(new_n761), .ZN(new_n762));
  XNOR2_X1  g576(.A(new_n762), .B(G131), .ZN(G33));
  INV_X1    g577(.A(new_n658), .ZN(new_n764));
  OAI21_X1  g578(.A(KEYINPUT112), .B1(new_n755), .B2(new_n764), .ZN(new_n765));
  INV_X1    g579(.A(KEYINPUT112), .ZN(new_n766));
  NAND4_X1  g580(.A1(new_n760), .A2(new_n766), .A3(new_n549), .A4(new_n658), .ZN(new_n767));
  NAND2_X1  g581(.A1(new_n765), .A2(new_n767), .ZN(new_n768));
  XNOR2_X1  g582(.A(new_n768), .B(G134), .ZN(G36));
  NAND2_X1  g583(.A1(new_n747), .A2(KEYINPUT45), .ZN(new_n770));
  OAI211_X1 g584(.A(new_n770), .B(G469), .C1(KEYINPUT45), .C2(new_n597), .ZN(new_n771));
  NAND2_X1  g585(.A1(G469), .A2(G902), .ZN(new_n772));
  NAND2_X1  g586(.A1(new_n771), .A2(new_n772), .ZN(new_n773));
  INV_X1    g587(.A(KEYINPUT46), .ZN(new_n774));
  NAND3_X1  g588(.A1(new_n773), .A2(KEYINPUT113), .A3(new_n774), .ZN(new_n775));
  OAI211_X1 g589(.A(new_n775), .B(new_n592), .C1(new_n774), .C2(new_n773), .ZN(new_n776));
  AOI21_X1  g590(.A(KEYINPUT113), .B1(new_n773), .B2(new_n774), .ZN(new_n777));
  NOR2_X1   g591(.A1(new_n776), .A2(new_n777), .ZN(new_n778));
  NOR2_X1   g592(.A1(new_n778), .A2(new_n551), .ZN(new_n779));
  NAND2_X1  g593(.A1(new_n779), .A2(new_n680), .ZN(new_n780));
  NAND2_X1  g594(.A1(new_n369), .A2(new_n614), .ZN(new_n781));
  XNOR2_X1  g595(.A(new_n781), .B(KEYINPUT43), .ZN(new_n782));
  NOR3_X1   g596(.A1(new_n782), .A2(new_n606), .A3(new_n662), .ZN(new_n783));
  AOI21_X1  g597(.A(new_n758), .B1(new_n783), .B2(KEYINPUT44), .ZN(new_n784));
  OAI21_X1  g598(.A(new_n784), .B1(KEYINPUT44), .B2(new_n783), .ZN(new_n785));
  NOR2_X1   g599(.A1(new_n780), .A2(new_n785), .ZN(new_n786));
  XNOR2_X1  g600(.A(new_n786), .B(new_n446), .ZN(G39));
  NOR2_X1   g601(.A1(new_n779), .A2(KEYINPUT47), .ZN(new_n788));
  INV_X1    g602(.A(new_n788), .ZN(new_n789));
  NAND2_X1  g603(.A1(new_n779), .A2(KEYINPUT47), .ZN(new_n790));
  NAND2_X1  g604(.A1(new_n789), .A2(new_n790), .ZN(new_n791));
  NOR4_X1   g605(.A1(new_n758), .A2(new_n647), .A3(new_n756), .A4(new_n442), .ZN(new_n792));
  NAND2_X1  g606(.A1(new_n791), .A2(new_n792), .ZN(new_n793));
  XNOR2_X1  g607(.A(new_n793), .B(G140), .ZN(G42));
  NOR2_X1   g608(.A1(new_n758), .A2(new_n713), .ZN(new_n795));
  INV_X1    g609(.A(new_n795), .ZN(new_n796));
  NAND3_X1  g610(.A1(new_n676), .A2(new_n442), .A3(new_n188), .ZN(new_n797));
  NOR2_X1   g611(.A1(new_n796), .A2(new_n797), .ZN(new_n798));
  NOR2_X1   g612(.A1(new_n615), .A2(new_n369), .ZN(new_n799));
  NAND2_X1  g613(.A1(new_n798), .A2(new_n799), .ZN(new_n800));
  NAND3_X1  g614(.A1(new_n800), .A2(G952), .A3(new_n190), .ZN(new_n801));
  NOR2_X1   g615(.A1(new_n782), .A2(new_n655), .ZN(new_n802));
  NAND2_X1  g616(.A1(new_n802), .A2(new_n795), .ZN(new_n803));
  INV_X1    g617(.A(new_n549), .ZN(new_n804));
  NOR2_X1   g618(.A1(new_n803), .A2(new_n804), .ZN(new_n805));
  XNOR2_X1  g619(.A(new_n805), .B(KEYINPUT48), .ZN(new_n806));
  AND2_X1   g620(.A1(new_n731), .A2(new_n802), .ZN(new_n807));
  AOI211_X1 g621(.A(new_n801), .B(new_n806), .C1(new_n714), .C2(new_n807), .ZN(new_n808));
  NAND3_X1  g622(.A1(new_n697), .A2(KEYINPUT118), .A3(new_n196), .ZN(new_n809));
  INV_X1    g623(.A(KEYINPUT118), .ZN(new_n810));
  OAI21_X1  g624(.A(new_n810), .B1(new_n713), .B2(new_n197), .ZN(new_n811));
  NAND4_X1  g625(.A1(new_n807), .A2(new_n671), .A3(new_n809), .A4(new_n811), .ZN(new_n812));
  XNOR2_X1  g626(.A(new_n812), .B(KEYINPUT50), .ZN(new_n813));
  NAND3_X1  g627(.A1(new_n798), .A2(new_n369), .A3(new_n615), .ZN(new_n814));
  NAND3_X1  g628(.A1(new_n725), .A2(new_n726), .A3(new_n635), .ZN(new_n815));
  OAI21_X1  g629(.A(new_n814), .B1(new_n815), .B2(new_n803), .ZN(new_n816));
  NOR2_X1   g630(.A1(new_n813), .A2(new_n816), .ZN(new_n817));
  INV_X1    g631(.A(new_n817), .ZN(new_n818));
  NAND2_X1  g632(.A1(new_n696), .A2(new_n592), .ZN(new_n819));
  INV_X1    g633(.A(new_n819), .ZN(new_n820));
  AOI21_X1  g634(.A(new_n791), .B1(new_n551), .B2(new_n820), .ZN(new_n821));
  NAND2_X1  g635(.A1(new_n807), .A2(new_n754), .ZN(new_n822));
  OAI21_X1  g636(.A(KEYINPUT51), .B1(new_n821), .B2(new_n822), .ZN(new_n823));
  NAND2_X1  g637(.A1(new_n820), .A2(new_n551), .ZN(new_n824));
  INV_X1    g638(.A(KEYINPUT117), .ZN(new_n825));
  OAI21_X1  g639(.A(new_n824), .B1(new_n791), .B2(new_n825), .ZN(new_n826));
  AOI21_X1  g640(.A(KEYINPUT117), .B1(new_n789), .B2(new_n790), .ZN(new_n827));
  OAI211_X1 g641(.A(new_n754), .B(new_n807), .C1(new_n826), .C2(new_n827), .ZN(new_n828));
  AND2_X1   g642(.A1(new_n828), .A2(new_n817), .ZN(new_n829));
  OAI221_X1 g643(.A(new_n808), .B1(new_n818), .B2(new_n823), .C1(new_n829), .C2(KEYINPUT51), .ZN(new_n830));
  NAND2_X1  g644(.A1(new_n401), .A2(new_n403), .ZN(new_n831));
  NOR4_X1   g645(.A1(new_n758), .A2(new_n368), .A3(new_n831), .A4(new_n657), .ZN(new_n832));
  INV_X1    g646(.A(new_n740), .ZN(new_n833));
  AOI22_X1  g647(.A1(new_n832), .A2(new_n686), .B1(new_n760), .B2(new_n833), .ZN(new_n834));
  NAND3_X1  g648(.A1(new_n762), .A2(new_n768), .A3(new_n834), .ZN(new_n835));
  INV_X1    g649(.A(new_n737), .ZN(new_n836));
  AOI21_X1  g650(.A(new_n736), .B1(new_n731), .B2(new_n733), .ZN(new_n837));
  NOR2_X1   g651(.A1(new_n836), .A2(new_n837), .ZN(new_n838));
  AOI21_X1  g652(.A(new_n799), .B1(new_n369), .B2(new_n831), .ZN(new_n839));
  NOR2_X1   g653(.A1(new_n839), .A2(new_n313), .ZN(new_n840));
  NAND2_X1  g654(.A1(new_n607), .A2(new_n840), .ZN(new_n841));
  AOI22_X1  g655(.A1(new_n616), .A2(new_n698), .B1(new_n711), .B2(new_n714), .ZN(new_n842));
  OAI211_X1 g656(.A(new_n408), .B(new_n600), .C1(new_n638), .C2(new_n549), .ZN(new_n843));
  NAND4_X1  g657(.A1(new_n707), .A2(new_n841), .A3(new_n842), .A4(new_n843), .ZN(new_n844));
  NOR3_X1   g658(.A1(new_n835), .A2(new_n838), .A3(new_n844), .ZN(new_n845));
  INV_X1    g659(.A(KEYINPUT52), .ZN(new_n846));
  NAND3_X1  g660(.A1(new_n751), .A2(new_n662), .A3(new_n656), .ZN(new_n847));
  NOR3_X1   g661(.A1(new_n732), .A2(new_n847), .A3(new_n676), .ZN(new_n848));
  INV_X1    g662(.A(new_n688), .ZN(new_n849));
  AOI21_X1  g663(.A(new_n652), .B1(KEYINPUT102), .B2(new_n849), .ZN(new_n850));
  AOI21_X1  g664(.A(new_n848), .B1(new_n850), .B2(new_n690), .ZN(new_n851));
  AOI21_X1  g665(.A(new_n741), .B1(new_n660), .B2(new_n664), .ZN(new_n852));
  AND3_X1   g666(.A1(new_n851), .A2(new_n852), .A3(KEYINPUT115), .ZN(new_n853));
  AOI21_X1  g667(.A(KEYINPUT115), .B1(new_n851), .B2(new_n852), .ZN(new_n854));
  OAI21_X1  g668(.A(new_n846), .B1(new_n853), .B2(new_n854), .ZN(new_n855));
  INV_X1    g669(.A(new_n741), .ZN(new_n856));
  INV_X1    g670(.A(new_n848), .ZN(new_n857));
  NAND4_X1  g671(.A1(new_n665), .A2(new_n693), .A3(new_n856), .A4(new_n857), .ZN(new_n858));
  INV_X1    g672(.A(KEYINPUT115), .ZN(new_n859));
  NAND2_X1  g673(.A1(new_n858), .A2(new_n859), .ZN(new_n860));
  NAND3_X1  g674(.A1(new_n851), .A2(KEYINPUT115), .A3(new_n852), .ZN(new_n861));
  NAND3_X1  g675(.A1(new_n860), .A2(KEYINPUT52), .A3(new_n861), .ZN(new_n862));
  NAND3_X1  g676(.A1(new_n845), .A2(new_n855), .A3(new_n862), .ZN(new_n863));
  INV_X1    g677(.A(KEYINPUT53), .ZN(new_n864));
  NAND2_X1  g678(.A1(new_n863), .A2(new_n864), .ZN(new_n865));
  AOI21_X1  g679(.A(KEYINPUT52), .B1(new_n860), .B2(new_n861), .ZN(new_n866));
  AND4_X1   g680(.A1(new_n707), .A2(new_n841), .A3(new_n842), .A4(new_n843), .ZN(new_n867));
  AOI22_X1  g681(.A1(new_n757), .A2(new_n761), .B1(new_n765), .B2(new_n767), .ZN(new_n868));
  NAND4_X1  g682(.A1(new_n867), .A2(new_n868), .A3(new_n738), .A4(new_n834), .ZN(new_n869));
  NOR2_X1   g683(.A1(new_n866), .A2(new_n869), .ZN(new_n870));
  NAND2_X1  g684(.A1(new_n858), .A2(KEYINPUT52), .ZN(new_n871));
  NAND3_X1  g685(.A1(new_n870), .A2(KEYINPUT53), .A3(new_n871), .ZN(new_n872));
  INV_X1    g686(.A(KEYINPUT54), .ZN(new_n873));
  NAND3_X1  g687(.A1(new_n865), .A2(new_n872), .A3(new_n873), .ZN(new_n874));
  OR2_X1    g688(.A1(new_n874), .A2(KEYINPUT116), .ZN(new_n875));
  NAND2_X1  g689(.A1(new_n870), .A2(new_n871), .ZN(new_n876));
  NAND2_X1  g690(.A1(new_n876), .A2(new_n864), .ZN(new_n877));
  OAI21_X1  g691(.A(new_n877), .B1(new_n864), .B2(new_n863), .ZN(new_n878));
  NAND2_X1  g692(.A1(new_n878), .A2(KEYINPUT54), .ZN(new_n879));
  NAND2_X1  g693(.A1(new_n874), .A2(KEYINPUT116), .ZN(new_n880));
  NAND3_X1  g694(.A1(new_n875), .A2(new_n879), .A3(new_n880), .ZN(new_n881));
  OAI22_X1  g695(.A1(new_n830), .A2(new_n881), .B1(G952), .B2(G953), .ZN(new_n882));
  NOR4_X1   g696(.A1(new_n443), .A2(new_n781), .A3(new_n551), .A4(new_n196), .ZN(new_n883));
  INV_X1    g697(.A(KEYINPUT49), .ZN(new_n884));
  OAI21_X1  g698(.A(new_n883), .B1(new_n884), .B2(new_n820), .ZN(new_n885));
  XNOR2_X1  g699(.A(new_n885), .B(KEYINPUT114), .ZN(new_n886));
  NAND2_X1  g700(.A1(new_n820), .A2(new_n884), .ZN(new_n887));
  NAND3_X1  g701(.A1(new_n671), .A2(new_n676), .A3(new_n887), .ZN(new_n888));
  OAI21_X1  g702(.A(new_n882), .B1(new_n886), .B2(new_n888), .ZN(G75));
  NOR2_X1   g703(.A1(new_n190), .A2(G952), .ZN(new_n890));
  INV_X1    g704(.A(new_n890), .ZN(new_n891));
  AOI21_X1  g705(.A(new_n189), .B1(new_n865), .B2(new_n872), .ZN(new_n892));
  AOI21_X1  g706(.A(KEYINPUT56), .B1(new_n892), .B2(G210), .ZN(new_n893));
  NAND2_X1  g707(.A1(new_n261), .A2(new_n289), .ZN(new_n894));
  NAND2_X1  g708(.A1(new_n894), .A2(new_n286), .ZN(new_n895));
  NAND2_X1  g709(.A1(new_n895), .A2(new_n290), .ZN(new_n896));
  XOR2_X1   g710(.A(new_n896), .B(KEYINPUT55), .Z(new_n897));
  OAI21_X1  g711(.A(new_n891), .B1(new_n893), .B2(new_n897), .ZN(new_n898));
  AOI21_X1  g712(.A(new_n898), .B1(new_n893), .B2(new_n897), .ZN(G51));
  AOI211_X1 g713(.A(new_n189), .B(new_n771), .C1(new_n865), .C2(new_n872), .ZN(new_n900));
  INV_X1    g714(.A(new_n590), .ZN(new_n901));
  AOI21_X1  g715(.A(KEYINPUT53), .B1(new_n870), .B2(new_n862), .ZN(new_n902));
  AND4_X1   g716(.A1(KEYINPUT53), .A2(new_n845), .A3(new_n855), .A4(new_n871), .ZN(new_n903));
  OAI21_X1  g717(.A(KEYINPUT54), .B1(new_n902), .B2(new_n903), .ZN(new_n904));
  NAND2_X1  g718(.A1(new_n904), .A2(KEYINPUT119), .ZN(new_n905));
  NAND2_X1  g719(.A1(new_n865), .A2(new_n872), .ZN(new_n906));
  INV_X1    g720(.A(KEYINPUT119), .ZN(new_n907));
  NAND3_X1  g721(.A1(new_n906), .A2(new_n907), .A3(KEYINPUT54), .ZN(new_n908));
  NAND3_X1  g722(.A1(new_n905), .A2(new_n874), .A3(new_n908), .ZN(new_n909));
  XOR2_X1   g723(.A(new_n772), .B(KEYINPUT57), .Z(new_n910));
  AOI21_X1  g724(.A(new_n901), .B1(new_n909), .B2(new_n910), .ZN(new_n911));
  INV_X1    g725(.A(KEYINPUT120), .ZN(new_n912));
  AOI21_X1  g726(.A(new_n900), .B1(new_n911), .B2(new_n912), .ZN(new_n913));
  AOI21_X1  g727(.A(new_n873), .B1(new_n865), .B2(new_n872), .ZN(new_n914));
  OAI21_X1  g728(.A(new_n874), .B1(new_n914), .B2(new_n907), .ZN(new_n915));
  NOR2_X1   g729(.A1(new_n904), .A2(KEYINPUT119), .ZN(new_n916));
  OAI21_X1  g730(.A(new_n910), .B1(new_n915), .B2(new_n916), .ZN(new_n917));
  NAND2_X1  g731(.A1(new_n917), .A2(new_n590), .ZN(new_n918));
  NAND2_X1  g732(.A1(new_n918), .A2(KEYINPUT120), .ZN(new_n919));
  AOI21_X1  g733(.A(new_n890), .B1(new_n913), .B2(new_n919), .ZN(G54));
  NAND3_X1  g734(.A1(new_n892), .A2(KEYINPUT58), .A3(G475), .ZN(new_n921));
  INV_X1    g735(.A(new_n363), .ZN(new_n922));
  AND2_X1   g736(.A1(new_n921), .A2(new_n922), .ZN(new_n923));
  NOR2_X1   g737(.A1(new_n921), .A2(new_n922), .ZN(new_n924));
  NOR3_X1   g738(.A1(new_n923), .A2(new_n924), .A3(new_n890), .ZN(G60));
  NAND2_X1  g739(.A1(G478), .A2(G902), .ZN(new_n926));
  XOR2_X1   g740(.A(new_n926), .B(KEYINPUT59), .Z(new_n927));
  INV_X1    g741(.A(new_n927), .ZN(new_n928));
  AOI21_X1  g742(.A(new_n611), .B1(new_n881), .B2(new_n928), .ZN(new_n929));
  AND3_X1   g743(.A1(new_n909), .A2(new_n611), .A3(new_n928), .ZN(new_n930));
  NOR3_X1   g744(.A1(new_n929), .A2(new_n930), .A3(new_n890), .ZN(G63));
  NAND2_X1  g745(.A1(G217), .A2(G902), .ZN(new_n932));
  XOR2_X1   g746(.A(new_n932), .B(KEYINPUT60), .Z(new_n933));
  NAND2_X1  g747(.A1(new_n906), .A2(new_n933), .ZN(new_n934));
  NAND2_X1  g748(.A1(new_n934), .A2(new_n433), .ZN(new_n935));
  NAND2_X1  g749(.A1(new_n935), .A2(new_n891), .ZN(new_n936));
  NOR2_X1   g750(.A1(new_n934), .A2(new_n633), .ZN(new_n937));
  INV_X1    g751(.A(KEYINPUT61), .ZN(new_n938));
  OAI22_X1  g752(.A1(new_n936), .A2(new_n937), .B1(KEYINPUT121), .B2(new_n938), .ZN(new_n939));
  NAND2_X1  g753(.A1(new_n938), .A2(KEYINPUT121), .ZN(new_n940));
  XNOR2_X1  g754(.A(new_n939), .B(new_n940), .ZN(G66));
  OAI21_X1  g755(.A(G953), .B1(new_n192), .B2(new_n281), .ZN(new_n942));
  NOR2_X1   g756(.A1(new_n838), .A2(new_n844), .ZN(new_n943));
  OAI21_X1  g757(.A(new_n942), .B1(new_n943), .B2(G953), .ZN(new_n944));
  OAI21_X1  g758(.A(new_n894), .B1(G898), .B2(new_n190), .ZN(new_n945));
  XNOR2_X1  g759(.A(new_n944), .B(new_n945), .ZN(G69));
  XOR2_X1   g760(.A(new_n507), .B(new_n353), .Z(new_n947));
  INV_X1    g761(.A(new_n681), .ZN(new_n948));
  NOR3_X1   g762(.A1(new_n804), .A2(new_n758), .A3(new_n839), .ZN(new_n949));
  AOI21_X1  g763(.A(new_n786), .B1(new_n948), .B2(new_n949), .ZN(new_n950));
  NAND2_X1  g764(.A1(new_n950), .A2(new_n793), .ZN(new_n951));
  NAND2_X1  g765(.A1(new_n852), .A2(new_n693), .ZN(new_n952));
  XNOR2_X1  g766(.A(new_n952), .B(KEYINPUT122), .ZN(new_n953));
  NAND2_X1  g767(.A1(new_n953), .A2(new_n684), .ZN(new_n954));
  AOI21_X1  g768(.A(new_n951), .B1(new_n954), .B2(KEYINPUT62), .ZN(new_n955));
  OR2_X1    g769(.A1(new_n954), .A2(KEYINPUT62), .ZN(new_n956));
  AOI211_X1 g770(.A(G953), .B(new_n947), .C1(new_n955), .C2(new_n956), .ZN(new_n957));
  NAND2_X1  g771(.A1(new_n653), .A2(G953), .ZN(new_n958));
  XNOR2_X1  g772(.A(new_n958), .B(KEYINPUT123), .ZN(new_n959));
  NAND2_X1  g773(.A1(new_n947), .A2(new_n959), .ZN(new_n960));
  NOR2_X1   g774(.A1(new_n868), .A2(KEYINPUT124), .ZN(new_n961));
  NAND3_X1  g775(.A1(new_n549), .A2(new_n691), .A3(new_n677), .ZN(new_n962));
  AOI21_X1  g776(.A(new_n780), .B1(new_n785), .B2(new_n962), .ZN(new_n963));
  AOI211_X1 g777(.A(new_n961), .B(new_n963), .C1(new_n791), .C2(new_n792), .ZN(new_n964));
  NAND2_X1  g778(.A1(new_n868), .A2(KEYINPUT124), .ZN(new_n965));
  NAND3_X1  g779(.A1(new_n964), .A2(new_n953), .A3(new_n965), .ZN(new_n966));
  AOI21_X1  g780(.A(new_n960), .B1(new_n966), .B2(new_n190), .ZN(new_n967));
  INV_X1    g781(.A(KEYINPUT125), .ZN(new_n968));
  OAI21_X1  g782(.A(G953), .B1(new_n566), .B2(new_n653), .ZN(new_n969));
  OAI22_X1  g783(.A1(new_n957), .A2(new_n967), .B1(new_n968), .B2(new_n969), .ZN(new_n970));
  NAND2_X1  g784(.A1(new_n969), .A2(new_n968), .ZN(new_n971));
  XNOR2_X1  g785(.A(new_n970), .B(new_n971), .ZN(G72));
  INV_X1    g786(.A(new_n529), .ZN(new_n973));
  NAND3_X1  g787(.A1(new_n955), .A2(new_n943), .A3(new_n956), .ZN(new_n974));
  NAND2_X1  g788(.A1(G472), .A2(G902), .ZN(new_n975));
  XOR2_X1   g789(.A(new_n975), .B(KEYINPUT63), .Z(new_n976));
  XNOR2_X1  g790(.A(new_n976), .B(KEYINPUT126), .ZN(new_n977));
  AOI211_X1 g791(.A(new_n483), .B(new_n973), .C1(new_n974), .C2(new_n977), .ZN(new_n978));
  INV_X1    g792(.A(new_n943), .ZN(new_n979));
  OAI21_X1  g793(.A(new_n977), .B1(new_n966), .B2(new_n979), .ZN(new_n980));
  AND3_X1   g794(.A1(new_n980), .A2(new_n483), .A3(new_n973), .ZN(new_n981));
  NAND2_X1  g795(.A1(new_n672), .A2(new_n530), .ZN(new_n982));
  AND3_X1   g796(.A1(new_n878), .A2(new_n976), .A3(new_n982), .ZN(new_n983));
  NOR4_X1   g797(.A1(new_n978), .A2(new_n981), .A3(new_n890), .A4(new_n983), .ZN(G57));
endmodule


