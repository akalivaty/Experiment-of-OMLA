//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 0 0 1 0 0 1 0 0 0 1 1 1 0 1 1 1 0 1 1 1 0 0 1 0 1 1 1 0 1 1 1 0 0 0 0 1 0 0 1 1 0 0 0 1 1 0 0 1 0 1 0 1 0 0 1 0 1 0 0 0 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:25:13 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n697, new_n698, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n716, new_n718, new_n720, new_n721,
    new_n722, new_n723, new_n724, new_n725, new_n726, new_n727, new_n729,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n742, new_n743, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n774, new_n775,
    new_n776, new_n777, new_n778, new_n779, new_n780, new_n781, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n898, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n906, new_n907, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n925, new_n926,
    new_n927, new_n928, new_n930, new_n931, new_n932, new_n933, new_n934,
    new_n935, new_n936, new_n938, new_n939, new_n940, new_n941, new_n942,
    new_n943, new_n944, new_n945, new_n946, new_n948, new_n949, new_n950,
    new_n951, new_n952, new_n953, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n982, new_n983, new_n984, new_n985, new_n986, new_n987,
    new_n988, new_n989, new_n990, new_n991, new_n992, new_n993, new_n994,
    new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001;
  OAI21_X1  g000(.A(G214), .B1(G237), .B2(G902), .ZN(new_n187));
  INV_X1    g001(.A(new_n187), .ZN(new_n188));
  OAI21_X1  g002(.A(G210), .B1(G237), .B2(G902), .ZN(new_n189));
  XOR2_X1   g003(.A(new_n189), .B(KEYINPUT82), .Z(new_n190));
  INV_X1    g004(.A(new_n190), .ZN(new_n191));
  AND2_X1   g005(.A1(KEYINPUT64), .A2(G146), .ZN(new_n192));
  NOR2_X1   g006(.A1(KEYINPUT64), .A2(G146), .ZN(new_n193));
  OAI21_X1  g007(.A(G143), .B1(new_n192), .B2(new_n193), .ZN(new_n194));
  INV_X1    g008(.A(KEYINPUT1), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n195), .A2(KEYINPUT68), .ZN(new_n196));
  INV_X1    g010(.A(KEYINPUT68), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n197), .A2(KEYINPUT1), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n196), .A2(new_n198), .ZN(new_n199));
  INV_X1    g013(.A(G146), .ZN(new_n200));
  NOR2_X1   g014(.A1(new_n200), .A2(G143), .ZN(new_n201));
  INV_X1    g015(.A(new_n201), .ZN(new_n202));
  NAND4_X1  g016(.A1(new_n194), .A2(new_n199), .A3(G128), .A4(new_n202), .ZN(new_n203));
  XNOR2_X1  g017(.A(KEYINPUT69), .B(G128), .ZN(new_n204));
  XNOR2_X1  g018(.A(KEYINPUT68), .B(KEYINPUT1), .ZN(new_n205));
  AOI21_X1  g019(.A(new_n204), .B1(new_n194), .B2(new_n205), .ZN(new_n206));
  INV_X1    g020(.A(G143), .ZN(new_n207));
  NOR2_X1   g021(.A1(new_n207), .A2(G146), .ZN(new_n208));
  NOR2_X1   g022(.A1(new_n192), .A2(new_n193), .ZN(new_n209));
  AOI21_X1  g023(.A(new_n208), .B1(new_n209), .B2(new_n207), .ZN(new_n210));
  OAI21_X1  g024(.A(new_n203), .B1(new_n206), .B2(new_n210), .ZN(new_n211));
  OR2_X1    g025(.A1(new_n211), .A2(G125), .ZN(new_n212));
  NAND3_X1  g026(.A1(new_n194), .A2(G128), .A3(new_n202), .ZN(new_n213));
  INV_X1    g027(.A(KEYINPUT0), .ZN(new_n214));
  XOR2_X1   g028(.A(KEYINPUT0), .B(G128), .Z(new_n215));
  INV_X1    g029(.A(new_n215), .ZN(new_n216));
  OAI22_X1  g030(.A1(new_n213), .A2(new_n214), .B1(new_n210), .B2(new_n216), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n217), .A2(G125), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n212), .A2(new_n218), .ZN(new_n219));
  INV_X1    g033(.A(KEYINPUT80), .ZN(new_n220));
  INV_X1    g034(.A(G224), .ZN(new_n221));
  OAI21_X1  g035(.A(new_n220), .B1(new_n221), .B2(G953), .ZN(new_n222));
  INV_X1    g036(.A(G953), .ZN(new_n223));
  NAND3_X1  g037(.A1(new_n223), .A2(KEYINPUT80), .A3(G224), .ZN(new_n224));
  NAND2_X1  g038(.A1(new_n222), .A2(new_n224), .ZN(new_n225));
  XOR2_X1   g039(.A(new_n225), .B(KEYINPUT81), .Z(new_n226));
  XNOR2_X1  g040(.A(new_n219), .B(new_n226), .ZN(new_n227));
  XOR2_X1   g041(.A(G110), .B(G122), .Z(new_n228));
  INV_X1    g042(.A(G104), .ZN(new_n229));
  OAI21_X1  g043(.A(KEYINPUT3), .B1(new_n229), .B2(G107), .ZN(new_n230));
  INV_X1    g044(.A(KEYINPUT77), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n230), .A2(new_n231), .ZN(new_n232));
  NOR2_X1   g046(.A1(new_n229), .A2(G107), .ZN(new_n233));
  INV_X1    g047(.A(KEYINPUT3), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n233), .A2(new_n234), .ZN(new_n235));
  INV_X1    g049(.A(G107), .ZN(new_n236));
  NOR2_X1   g050(.A1(new_n236), .A2(G104), .ZN(new_n237));
  INV_X1    g051(.A(new_n237), .ZN(new_n238));
  OAI211_X1 g052(.A(KEYINPUT77), .B(KEYINPUT3), .C1(new_n229), .C2(G107), .ZN(new_n239));
  NAND4_X1  g053(.A1(new_n232), .A2(new_n235), .A3(new_n238), .A4(new_n239), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n240), .A2(G101), .ZN(new_n241));
  AOI21_X1  g055(.A(new_n237), .B1(new_n234), .B2(new_n233), .ZN(new_n242));
  INV_X1    g056(.A(G101), .ZN(new_n243));
  NAND4_X1  g057(.A1(new_n242), .A2(new_n243), .A3(new_n232), .A4(new_n239), .ZN(new_n244));
  NAND3_X1  g058(.A1(new_n241), .A2(KEYINPUT4), .A3(new_n244), .ZN(new_n245));
  XOR2_X1   g059(.A(KEYINPUT2), .B(G113), .Z(new_n246));
  XNOR2_X1  g060(.A(G116), .B(G119), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n246), .A2(new_n247), .ZN(new_n248));
  INV_X1    g062(.A(KEYINPUT70), .ZN(new_n249));
  XNOR2_X1  g063(.A(new_n247), .B(new_n249), .ZN(new_n250));
  OAI21_X1  g064(.A(new_n248), .B1(new_n250), .B2(new_n246), .ZN(new_n251));
  INV_X1    g065(.A(KEYINPUT4), .ZN(new_n252));
  NAND3_X1  g066(.A1(new_n240), .A2(new_n252), .A3(G101), .ZN(new_n253));
  NAND3_X1  g067(.A1(new_n245), .A2(new_n251), .A3(new_n253), .ZN(new_n254));
  INV_X1    g068(.A(G113), .ZN(new_n255));
  INV_X1    g069(.A(G116), .ZN(new_n256));
  NOR2_X1   g070(.A1(new_n256), .A2(G119), .ZN(new_n257));
  INV_X1    g071(.A(KEYINPUT5), .ZN(new_n258));
  AOI21_X1  g072(.A(new_n255), .B1(new_n257), .B2(new_n258), .ZN(new_n259));
  XNOR2_X1  g073(.A(new_n247), .B(KEYINPUT70), .ZN(new_n260));
  OAI21_X1  g074(.A(new_n259), .B1(new_n260), .B2(new_n258), .ZN(new_n261));
  OAI21_X1  g075(.A(G101), .B1(new_n233), .B2(new_n237), .ZN(new_n262));
  AND2_X1   g076(.A1(new_n244), .A2(new_n262), .ZN(new_n263));
  NAND3_X1  g077(.A1(new_n261), .A2(new_n263), .A3(new_n248), .ZN(new_n264));
  INV_X1    g078(.A(KEYINPUT79), .ZN(new_n265));
  AND3_X1   g079(.A1(new_n254), .A2(new_n264), .A3(new_n265), .ZN(new_n266));
  AOI21_X1  g080(.A(new_n265), .B1(new_n254), .B2(new_n264), .ZN(new_n267));
  OAI21_X1  g081(.A(new_n228), .B1(new_n266), .B2(new_n267), .ZN(new_n268));
  INV_X1    g082(.A(KEYINPUT6), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n254), .A2(new_n264), .ZN(new_n270));
  NOR2_X1   g084(.A1(new_n270), .A2(new_n228), .ZN(new_n271));
  OAI21_X1  g085(.A(new_n268), .B1(new_n269), .B2(new_n271), .ZN(new_n272));
  OAI211_X1 g086(.A(KEYINPUT6), .B(new_n228), .C1(new_n266), .C2(new_n267), .ZN(new_n273));
  AOI21_X1  g087(.A(new_n227), .B1(new_n272), .B2(new_n273), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n244), .A2(new_n262), .ZN(new_n275));
  NAND3_X1  g089(.A1(new_n261), .A2(new_n248), .A3(new_n275), .ZN(new_n276));
  XOR2_X1   g090(.A(new_n228), .B(KEYINPUT8), .Z(new_n277));
  NAND2_X1  g091(.A1(new_n247), .A2(KEYINPUT5), .ZN(new_n278));
  AOI22_X1  g092(.A1(new_n278), .A2(new_n259), .B1(new_n246), .B2(new_n247), .ZN(new_n279));
  OAI211_X1 g093(.A(new_n276), .B(new_n277), .C1(new_n275), .C2(new_n279), .ZN(new_n280));
  NAND3_X1  g094(.A1(new_n222), .A2(KEYINPUT7), .A3(new_n224), .ZN(new_n281));
  AND3_X1   g095(.A1(new_n212), .A2(new_n218), .A3(new_n281), .ZN(new_n282));
  AOI21_X1  g096(.A(new_n281), .B1(new_n212), .B2(new_n218), .ZN(new_n283));
  OAI221_X1 g097(.A(new_n280), .B1(new_n270), .B2(new_n228), .C1(new_n282), .C2(new_n283), .ZN(new_n284));
  INV_X1    g098(.A(G902), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n284), .A2(new_n285), .ZN(new_n286));
  OAI21_X1  g100(.A(new_n191), .B1(new_n274), .B2(new_n286), .ZN(new_n287));
  INV_X1    g101(.A(new_n228), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n270), .A2(KEYINPUT79), .ZN(new_n289));
  NAND3_X1  g103(.A1(new_n254), .A2(new_n264), .A3(new_n265), .ZN(new_n290));
  AOI21_X1  g104(.A(new_n288), .B1(new_n289), .B2(new_n290), .ZN(new_n291));
  NOR2_X1   g105(.A1(new_n271), .A2(new_n269), .ZN(new_n292));
  OAI21_X1  g106(.A(new_n273), .B1(new_n291), .B2(new_n292), .ZN(new_n293));
  INV_X1    g107(.A(new_n227), .ZN(new_n294));
  NAND2_X1  g108(.A1(new_n293), .A2(new_n294), .ZN(new_n295));
  INV_X1    g109(.A(new_n286), .ZN(new_n296));
  NAND3_X1  g110(.A1(new_n295), .A2(new_n296), .A3(new_n189), .ZN(new_n297));
  AOI21_X1  g111(.A(new_n188), .B1(new_n287), .B2(new_n297), .ZN(new_n298));
  NAND3_X1  g112(.A1(new_n256), .A2(KEYINPUT14), .A3(G122), .ZN(new_n299));
  XNOR2_X1  g113(.A(G116), .B(G122), .ZN(new_n300));
  INV_X1    g114(.A(new_n300), .ZN(new_n301));
  OAI211_X1 g115(.A(G107), .B(new_n299), .C1(new_n301), .C2(KEYINPUT14), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n300), .A2(new_n236), .ZN(new_n303));
  NAND2_X1  g117(.A1(KEYINPUT69), .A2(G128), .ZN(new_n304));
  INV_X1    g118(.A(new_n304), .ZN(new_n305));
  NOR2_X1   g119(.A1(KEYINPUT69), .A2(G128), .ZN(new_n306));
  OAI21_X1  g120(.A(G143), .B1(new_n305), .B2(new_n306), .ZN(new_n307));
  INV_X1    g121(.A(G134), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n207), .A2(G128), .ZN(new_n309));
  AND3_X1   g123(.A1(new_n307), .A2(new_n308), .A3(new_n309), .ZN(new_n310));
  AOI21_X1  g124(.A(new_n308), .B1(new_n307), .B2(new_n309), .ZN(new_n311));
  OAI211_X1 g125(.A(new_n302), .B(new_n303), .C1(new_n310), .C2(new_n311), .ZN(new_n312));
  NAND3_X1  g126(.A1(new_n207), .A2(KEYINPUT13), .A3(G128), .ZN(new_n313));
  XOR2_X1   g127(.A(new_n313), .B(KEYINPUT86), .Z(new_n314));
  INV_X1    g128(.A(new_n306), .ZN(new_n315));
  AOI21_X1  g129(.A(new_n207), .B1(new_n315), .B2(new_n304), .ZN(new_n316));
  INV_X1    g130(.A(KEYINPUT13), .ZN(new_n317));
  OAI21_X1  g131(.A(new_n309), .B1(new_n316), .B2(new_n317), .ZN(new_n318));
  AOI21_X1  g132(.A(new_n308), .B1(new_n314), .B2(new_n318), .ZN(new_n319));
  XNOR2_X1  g133(.A(new_n300), .B(new_n236), .ZN(new_n320));
  NAND3_X1  g134(.A1(new_n307), .A2(new_n308), .A3(new_n309), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n320), .A2(new_n321), .ZN(new_n322));
  OAI21_X1  g136(.A(new_n312), .B1(new_n319), .B2(new_n322), .ZN(new_n323));
  XNOR2_X1  g137(.A(KEYINPUT9), .B(G234), .ZN(new_n324));
  INV_X1    g138(.A(G217), .ZN(new_n325));
  NOR3_X1   g139(.A1(new_n324), .A2(new_n325), .A3(G953), .ZN(new_n326));
  INV_X1    g140(.A(new_n326), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n323), .A2(new_n327), .ZN(new_n328));
  INV_X1    g142(.A(KEYINPUT87), .ZN(new_n329));
  OAI211_X1 g143(.A(new_n312), .B(new_n326), .C1(new_n319), .C2(new_n322), .ZN(new_n330));
  NAND3_X1  g144(.A1(new_n328), .A2(new_n329), .A3(new_n330), .ZN(new_n331));
  INV_X1    g145(.A(KEYINPUT89), .ZN(new_n332));
  NAND3_X1  g146(.A1(new_n323), .A2(KEYINPUT87), .A3(new_n327), .ZN(new_n333));
  NAND4_X1  g147(.A1(new_n331), .A2(new_n332), .A3(new_n285), .A4(new_n333), .ZN(new_n334));
  INV_X1    g148(.A(KEYINPUT15), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n335), .A2(G478), .ZN(new_n336));
  AND3_X1   g150(.A1(new_n334), .A2(KEYINPUT88), .A3(new_n336), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n334), .A2(KEYINPUT88), .ZN(new_n338));
  INV_X1    g152(.A(KEYINPUT88), .ZN(new_n339));
  NAND4_X1  g153(.A1(new_n331), .A2(new_n339), .A3(new_n285), .A4(new_n333), .ZN(new_n340));
  AND3_X1   g154(.A1(new_n340), .A2(new_n335), .A3(G478), .ZN(new_n341));
  AOI21_X1  g155(.A(new_n337), .B1(new_n338), .B2(new_n341), .ZN(new_n342));
  NOR2_X1   g156(.A1(G237), .A2(G953), .ZN(new_n343));
  NAND3_X1  g157(.A1(new_n343), .A2(G143), .A3(G214), .ZN(new_n344));
  INV_X1    g158(.A(new_n344), .ZN(new_n345));
  AOI21_X1  g159(.A(G143), .B1(new_n343), .B2(G214), .ZN(new_n346));
  OAI21_X1  g160(.A(G131), .B1(new_n345), .B2(new_n346), .ZN(new_n347));
  INV_X1    g161(.A(KEYINPUT17), .ZN(new_n348));
  INV_X1    g162(.A(G237), .ZN(new_n349));
  NAND3_X1  g163(.A1(new_n349), .A2(new_n223), .A3(G214), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n350), .A2(new_n207), .ZN(new_n351));
  INV_X1    g165(.A(G131), .ZN(new_n352));
  NAND3_X1  g166(.A1(new_n351), .A2(new_n352), .A3(new_n344), .ZN(new_n353));
  NAND3_X1  g167(.A1(new_n347), .A2(new_n348), .A3(new_n353), .ZN(new_n354));
  INV_X1    g168(.A(KEYINPUT16), .ZN(new_n355));
  INV_X1    g169(.A(G140), .ZN(new_n356));
  NAND3_X1  g170(.A1(new_n355), .A2(new_n356), .A3(G125), .ZN(new_n357));
  NAND2_X1  g171(.A1(G125), .A2(G140), .ZN(new_n358));
  INV_X1    g172(.A(new_n358), .ZN(new_n359));
  NOR2_X1   g173(.A1(G125), .A2(G140), .ZN(new_n360));
  NOR2_X1   g174(.A1(new_n359), .A2(new_n360), .ZN(new_n361));
  OAI21_X1  g175(.A(new_n357), .B1(new_n361), .B2(new_n355), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n362), .A2(new_n200), .ZN(new_n363));
  OAI211_X1 g177(.A(G146), .B(new_n357), .C1(new_n361), .C2(new_n355), .ZN(new_n364));
  AOI21_X1  g178(.A(new_n352), .B1(new_n351), .B2(new_n344), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n365), .A2(KEYINPUT17), .ZN(new_n366));
  NAND4_X1  g180(.A1(new_n354), .A2(new_n363), .A3(new_n364), .A4(new_n366), .ZN(new_n367));
  XNOR2_X1  g181(.A(G113), .B(G122), .ZN(new_n368));
  XNOR2_X1  g182(.A(new_n368), .B(new_n229), .ZN(new_n369));
  NAND2_X1  g183(.A1(KEYINPUT18), .A2(G131), .ZN(new_n370));
  NAND3_X1  g184(.A1(new_n351), .A2(new_n344), .A3(new_n370), .ZN(new_n371));
  INV_X1    g185(.A(new_n370), .ZN(new_n372));
  OAI21_X1  g186(.A(new_n372), .B1(new_n345), .B2(new_n346), .ZN(new_n373));
  OR2_X1    g187(.A1(G125), .A2(G140), .ZN(new_n374));
  NAND3_X1  g188(.A1(new_n374), .A2(G146), .A3(new_n358), .ZN(new_n375));
  INV_X1    g189(.A(KEYINPUT83), .ZN(new_n376));
  XNOR2_X1  g190(.A(new_n375), .B(new_n376), .ZN(new_n377));
  INV_X1    g191(.A(KEYINPUT74), .ZN(new_n378));
  OAI21_X1  g192(.A(new_n378), .B1(new_n359), .B2(new_n360), .ZN(new_n379));
  NAND3_X1  g193(.A1(new_n374), .A2(KEYINPUT74), .A3(new_n358), .ZN(new_n380));
  AOI21_X1  g194(.A(new_n209), .B1(new_n379), .B2(new_n380), .ZN(new_n381));
  OAI211_X1 g195(.A(new_n371), .B(new_n373), .C1(new_n377), .C2(new_n381), .ZN(new_n382));
  AND3_X1   g196(.A1(new_n367), .A2(new_n369), .A3(new_n382), .ZN(new_n383));
  NAND2_X1  g197(.A1(new_n367), .A2(new_n382), .ZN(new_n384));
  INV_X1    g198(.A(new_n369), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n384), .A2(new_n385), .ZN(new_n386));
  NAND2_X1  g200(.A1(new_n386), .A2(KEYINPUT85), .ZN(new_n387));
  INV_X1    g201(.A(KEYINPUT85), .ZN(new_n388));
  NAND3_X1  g202(.A1(new_n384), .A2(new_n388), .A3(new_n385), .ZN(new_n389));
  AOI21_X1  g203(.A(new_n383), .B1(new_n387), .B2(new_n389), .ZN(new_n390));
  OAI21_X1  g204(.A(G475), .B1(new_n390), .B2(G902), .ZN(new_n391));
  INV_X1    g205(.A(G475), .ZN(new_n392));
  INV_X1    g206(.A(KEYINPUT84), .ZN(new_n393));
  INV_X1    g207(.A(new_n353), .ZN(new_n394));
  OAI21_X1  g208(.A(new_n393), .B1(new_n394), .B2(new_n365), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n379), .A2(new_n380), .ZN(new_n396));
  INV_X1    g210(.A(KEYINPUT19), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n396), .A2(new_n397), .ZN(new_n398));
  OR2_X1    g212(.A1(KEYINPUT64), .A2(G146), .ZN(new_n399));
  NAND2_X1  g213(.A1(KEYINPUT64), .A2(G146), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n399), .A2(new_n400), .ZN(new_n401));
  NOR3_X1   g215(.A1(new_n359), .A2(new_n360), .A3(new_n397), .ZN(new_n402));
  INV_X1    g216(.A(new_n402), .ZN(new_n403));
  NAND3_X1  g217(.A1(new_n398), .A2(new_n401), .A3(new_n403), .ZN(new_n404));
  NAND3_X1  g218(.A1(new_n347), .A2(KEYINPUT84), .A3(new_n353), .ZN(new_n405));
  NAND4_X1  g219(.A1(new_n395), .A2(new_n404), .A3(new_n364), .A4(new_n405), .ZN(new_n406));
  AOI21_X1  g220(.A(new_n369), .B1(new_n406), .B2(new_n382), .ZN(new_n407));
  OAI211_X1 g221(.A(new_n392), .B(new_n285), .C1(new_n407), .C2(new_n383), .ZN(new_n408));
  NAND2_X1  g222(.A1(new_n408), .A2(KEYINPUT20), .ZN(new_n409));
  NAND3_X1  g223(.A1(new_n367), .A2(new_n382), .A3(new_n369), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n373), .A2(new_n371), .ZN(new_n411));
  INV_X1    g225(.A(new_n381), .ZN(new_n412));
  XNOR2_X1  g226(.A(new_n375), .B(KEYINPUT83), .ZN(new_n413));
  AOI21_X1  g227(.A(new_n411), .B1(new_n412), .B2(new_n413), .ZN(new_n414));
  AND3_X1   g228(.A1(new_n347), .A2(KEYINPUT84), .A3(new_n353), .ZN(new_n415));
  AOI21_X1  g229(.A(KEYINPUT84), .B1(new_n347), .B2(new_n353), .ZN(new_n416));
  NOR2_X1   g230(.A1(new_n415), .A2(new_n416), .ZN(new_n417));
  INV_X1    g231(.A(new_n364), .ZN(new_n418));
  AOI21_X1  g232(.A(new_n402), .B1(new_n396), .B2(new_n397), .ZN(new_n419));
  AOI21_X1  g233(.A(new_n418), .B1(new_n419), .B2(new_n401), .ZN(new_n420));
  AOI21_X1  g234(.A(new_n414), .B1(new_n417), .B2(new_n420), .ZN(new_n421));
  OAI21_X1  g235(.A(new_n410), .B1(new_n421), .B2(new_n369), .ZN(new_n422));
  INV_X1    g236(.A(KEYINPUT20), .ZN(new_n423));
  NAND4_X1  g237(.A1(new_n422), .A2(new_n423), .A3(new_n392), .A4(new_n285), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n409), .A2(new_n424), .ZN(new_n425));
  INV_X1    g239(.A(G952), .ZN(new_n426));
  NOR2_X1   g240(.A1(new_n426), .A2(G953), .ZN(new_n427));
  NAND2_X1  g241(.A1(G234), .A2(G237), .ZN(new_n428));
  NAND2_X1  g242(.A1(new_n427), .A2(new_n428), .ZN(new_n429));
  XOR2_X1   g243(.A(KEYINPUT21), .B(G898), .Z(new_n430));
  NAND3_X1  g244(.A1(new_n428), .A2(G902), .A3(G953), .ZN(new_n431));
  OAI21_X1  g245(.A(new_n429), .B1(new_n430), .B2(new_n431), .ZN(new_n432));
  NAND3_X1  g246(.A1(new_n391), .A2(new_n425), .A3(new_n432), .ZN(new_n433));
  INV_X1    g247(.A(KEYINPUT90), .ZN(new_n434));
  NOR3_X1   g248(.A1(new_n342), .A2(new_n433), .A3(new_n434), .ZN(new_n435));
  AND3_X1   g249(.A1(new_n391), .A2(new_n425), .A3(new_n432), .ZN(new_n436));
  NAND3_X1  g250(.A1(new_n334), .A2(KEYINPUT88), .A3(new_n336), .ZN(new_n437));
  INV_X1    g251(.A(new_n338), .ZN(new_n438));
  NAND3_X1  g252(.A1(new_n340), .A2(new_n335), .A3(G478), .ZN(new_n439));
  OAI21_X1  g253(.A(new_n437), .B1(new_n438), .B2(new_n439), .ZN(new_n440));
  AOI21_X1  g254(.A(KEYINPUT90), .B1(new_n436), .B2(new_n440), .ZN(new_n441));
  OAI21_X1  g255(.A(new_n298), .B1(new_n435), .B2(new_n441), .ZN(new_n442));
  INV_X1    g256(.A(G469), .ZN(new_n443));
  INV_X1    g257(.A(new_n213), .ZN(new_n444));
  INV_X1    g258(.A(new_n208), .ZN(new_n445));
  OAI21_X1  g259(.A(new_n445), .B1(new_n401), .B2(G143), .ZN(new_n446));
  AOI22_X1  g260(.A1(new_n444), .A2(KEYINPUT0), .B1(new_n446), .B2(new_n215), .ZN(new_n447));
  NAND3_X1  g261(.A1(new_n245), .A2(new_n447), .A3(new_n253), .ZN(new_n448));
  INV_X1    g262(.A(KEYINPUT10), .ZN(new_n449));
  OAI21_X1  g263(.A(G128), .B1(new_n208), .B2(new_n195), .ZN(new_n450));
  AOI21_X1  g264(.A(new_n207), .B1(new_n399), .B2(new_n400), .ZN(new_n451));
  OAI21_X1  g265(.A(new_n450), .B1(new_n451), .B2(new_n201), .ZN(new_n452));
  AND2_X1   g266(.A1(new_n452), .A2(new_n203), .ZN(new_n453));
  OAI21_X1  g267(.A(new_n449), .B1(new_n453), .B2(new_n275), .ZN(new_n454));
  INV_X1    g268(.A(KEYINPUT11), .ZN(new_n455));
  OAI21_X1  g269(.A(new_n455), .B1(new_n308), .B2(G137), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n456), .A2(KEYINPUT65), .ZN(new_n457));
  INV_X1    g271(.A(KEYINPUT65), .ZN(new_n458));
  OAI211_X1 g272(.A(new_n458), .B(new_n455), .C1(new_n308), .C2(G137), .ZN(new_n459));
  INV_X1    g273(.A(G137), .ZN(new_n460));
  NAND3_X1  g274(.A1(new_n460), .A2(KEYINPUT11), .A3(G134), .ZN(new_n461));
  INV_X1    g275(.A(KEYINPUT66), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  NAND4_X1  g277(.A1(new_n460), .A2(KEYINPUT66), .A3(KEYINPUT11), .A4(G134), .ZN(new_n464));
  AOI22_X1  g278(.A1(new_n457), .A2(new_n459), .B1(new_n463), .B2(new_n464), .ZN(new_n465));
  NOR2_X1   g279(.A1(new_n460), .A2(G134), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n466), .A2(KEYINPUT67), .ZN(new_n467));
  INV_X1    g281(.A(KEYINPUT67), .ZN(new_n468));
  OAI21_X1  g282(.A(new_n468), .B1(new_n460), .B2(G134), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n467), .A2(new_n469), .ZN(new_n470));
  AOI21_X1  g284(.A(new_n352), .B1(new_n465), .B2(new_n470), .ZN(new_n471));
  NAND2_X1  g285(.A1(new_n457), .A2(new_n459), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n463), .A2(new_n464), .ZN(new_n473));
  NAND4_X1  g287(.A1(new_n472), .A2(new_n473), .A3(new_n470), .A4(new_n352), .ZN(new_n474));
  INV_X1    g288(.A(new_n474), .ZN(new_n475));
  NOR2_X1   g289(.A1(new_n471), .A2(new_n475), .ZN(new_n476));
  NAND4_X1  g290(.A1(new_n211), .A2(KEYINPUT10), .A3(new_n244), .A4(new_n262), .ZN(new_n477));
  NAND4_X1  g291(.A1(new_n448), .A2(new_n454), .A3(new_n476), .A4(new_n477), .ZN(new_n478));
  XNOR2_X1  g292(.A(G110), .B(G140), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n223), .A2(G227), .ZN(new_n480));
  XNOR2_X1  g294(.A(new_n479), .B(new_n480), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n478), .A2(new_n481), .ZN(new_n482));
  NAND2_X1  g296(.A1(new_n452), .A2(new_n203), .ZN(new_n483));
  NAND3_X1  g297(.A1(new_n483), .A2(new_n244), .A3(new_n262), .ZN(new_n484));
  OAI21_X1  g298(.A(new_n484), .B1(new_n263), .B2(new_n211), .ZN(new_n485));
  NAND3_X1  g299(.A1(new_n472), .A2(new_n470), .A3(new_n473), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n486), .A2(G131), .ZN(new_n487));
  NAND2_X1  g301(.A1(new_n487), .A2(new_n474), .ZN(new_n488));
  NAND3_X1  g302(.A1(new_n485), .A2(KEYINPUT12), .A3(new_n488), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n485), .A2(new_n488), .ZN(new_n490));
  INV_X1    g304(.A(KEYINPUT12), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  AOI21_X1  g306(.A(new_n482), .B1(new_n489), .B2(new_n492), .ZN(new_n493));
  NAND3_X1  g307(.A1(new_n448), .A2(new_n454), .A3(new_n477), .ZN(new_n494));
  NAND2_X1  g308(.A1(new_n494), .A2(new_n488), .ZN(new_n495));
  AOI21_X1  g309(.A(new_n481), .B1(new_n495), .B2(new_n478), .ZN(new_n496));
  OAI211_X1 g310(.A(new_n443), .B(new_n285), .C1(new_n493), .C2(new_n496), .ZN(new_n497));
  AND3_X1   g311(.A1(new_n485), .A2(KEYINPUT12), .A3(new_n488), .ZN(new_n498));
  AOI21_X1  g312(.A(KEYINPUT12), .B1(new_n485), .B2(new_n488), .ZN(new_n499));
  OAI21_X1  g313(.A(new_n478), .B1(new_n498), .B2(new_n499), .ZN(new_n500));
  INV_X1    g314(.A(new_n481), .ZN(new_n501));
  NAND2_X1  g315(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  AND2_X1   g316(.A1(new_n478), .A2(new_n481), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n503), .A2(new_n495), .ZN(new_n504));
  NAND3_X1  g318(.A1(new_n502), .A2(G469), .A3(new_n504), .ZN(new_n505));
  NAND2_X1  g319(.A1(G469), .A2(G902), .ZN(new_n506));
  NAND3_X1  g320(.A1(new_n497), .A2(new_n505), .A3(new_n506), .ZN(new_n507));
  INV_X1    g321(.A(G221), .ZN(new_n508));
  INV_X1    g322(.A(new_n324), .ZN(new_n509));
  AOI21_X1  g323(.A(new_n508), .B1(new_n509), .B2(new_n285), .ZN(new_n510));
  INV_X1    g324(.A(new_n510), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n507), .A2(new_n511), .ZN(new_n512));
  INV_X1    g326(.A(KEYINPUT78), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  NAND3_X1  g328(.A1(new_n507), .A2(KEYINPUT78), .A3(new_n511), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  OAI21_X1  g330(.A(KEYINPUT91), .B1(new_n442), .B2(new_n516), .ZN(new_n517));
  AND3_X1   g331(.A1(new_n507), .A2(KEYINPUT78), .A3(new_n511), .ZN(new_n518));
  AOI21_X1  g332(.A(KEYINPUT78), .B1(new_n507), .B2(new_n511), .ZN(new_n519));
  NOR2_X1   g333(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  INV_X1    g334(.A(KEYINPUT91), .ZN(new_n521));
  OAI21_X1  g335(.A(new_n434), .B1(new_n342), .B2(new_n433), .ZN(new_n522));
  NAND3_X1  g336(.A1(new_n436), .A2(new_n440), .A3(KEYINPUT90), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  NAND4_X1  g338(.A1(new_n520), .A2(new_n521), .A3(new_n298), .A4(new_n524), .ZN(new_n525));
  AOI21_X1  g339(.A(new_n217), .B1(new_n487), .B2(new_n474), .ZN(new_n526));
  NOR2_X1   g340(.A1(new_n308), .A2(G137), .ZN(new_n527));
  OAI21_X1  g341(.A(G131), .B1(new_n466), .B2(new_n527), .ZN(new_n528));
  AND3_X1   g342(.A1(new_n211), .A2(new_n474), .A3(new_n528), .ZN(new_n529));
  NOR3_X1   g343(.A1(new_n526), .A2(new_n529), .A3(new_n251), .ZN(new_n530));
  INV_X1    g344(.A(new_n251), .ZN(new_n531));
  OAI21_X1  g345(.A(new_n447), .B1(new_n471), .B2(new_n475), .ZN(new_n532));
  NAND3_X1  g346(.A1(new_n211), .A2(new_n474), .A3(new_n528), .ZN(new_n533));
  AOI21_X1  g347(.A(new_n531), .B1(new_n532), .B2(new_n533), .ZN(new_n534));
  OAI21_X1  g348(.A(KEYINPUT28), .B1(new_n530), .B2(new_n534), .ZN(new_n535));
  NAND3_X1  g349(.A1(new_n532), .A2(new_n531), .A3(new_n533), .ZN(new_n536));
  INV_X1    g350(.A(KEYINPUT28), .ZN(new_n537));
  NAND2_X1  g351(.A1(new_n536), .A2(new_n537), .ZN(new_n538));
  XNOR2_X1  g352(.A(KEYINPUT26), .B(KEYINPUT27), .ZN(new_n539));
  XNOR2_X1  g353(.A(new_n539), .B(G101), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n343), .A2(G210), .ZN(new_n541));
  XNOR2_X1  g355(.A(new_n540), .B(new_n541), .ZN(new_n542));
  NAND3_X1  g356(.A1(new_n535), .A2(new_n538), .A3(new_n542), .ZN(new_n543));
  INV_X1    g357(.A(KEYINPUT29), .ZN(new_n544));
  OAI21_X1  g358(.A(KEYINPUT30), .B1(new_n526), .B2(new_n529), .ZN(new_n545));
  INV_X1    g359(.A(KEYINPUT30), .ZN(new_n546));
  NAND3_X1  g360(.A1(new_n532), .A2(new_n546), .A3(new_n533), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n545), .A2(new_n547), .ZN(new_n548));
  AOI21_X1  g362(.A(new_n530), .B1(new_n548), .B2(new_n251), .ZN(new_n549));
  OAI211_X1 g363(.A(new_n543), .B(new_n544), .C1(new_n542), .C2(new_n549), .ZN(new_n550));
  OAI211_X1 g364(.A(new_n550), .B(new_n285), .C1(new_n544), .C2(new_n543), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n551), .A2(G472), .ZN(new_n552));
  NOR2_X1   g366(.A1(G472), .A2(G902), .ZN(new_n553));
  XOR2_X1   g367(.A(new_n553), .B(KEYINPUT71), .Z(new_n554));
  INV_X1    g368(.A(new_n554), .ZN(new_n555));
  INV_X1    g369(.A(new_n542), .ZN(new_n556));
  INV_X1    g370(.A(new_n538), .ZN(new_n557));
  OAI21_X1  g371(.A(new_n251), .B1(new_n526), .B2(new_n529), .ZN(new_n558));
  AOI21_X1  g372(.A(new_n537), .B1(new_n558), .B2(new_n536), .ZN(new_n559));
  OAI21_X1  g373(.A(new_n556), .B1(new_n557), .B2(new_n559), .ZN(new_n560));
  AOI21_X1  g374(.A(new_n531), .B1(new_n545), .B2(new_n547), .ZN(new_n561));
  NOR3_X1   g375(.A1(new_n561), .A2(new_n530), .A3(new_n556), .ZN(new_n562));
  INV_X1    g376(.A(KEYINPUT31), .ZN(new_n563));
  OAI21_X1  g377(.A(new_n560), .B1(new_n562), .B2(new_n563), .ZN(new_n564));
  NOR4_X1   g378(.A1(new_n561), .A2(KEYINPUT31), .A3(new_n530), .A4(new_n556), .ZN(new_n565));
  OAI211_X1 g379(.A(KEYINPUT32), .B(new_n555), .C1(new_n564), .C2(new_n565), .ZN(new_n566));
  INV_X1    g380(.A(KEYINPUT72), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n549), .A2(new_n542), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n569), .A2(KEYINPUT31), .ZN(new_n570));
  INV_X1    g384(.A(new_n565), .ZN(new_n571));
  NAND3_X1  g385(.A1(new_n570), .A2(new_n571), .A3(new_n560), .ZN(new_n572));
  AOI21_X1  g386(.A(KEYINPUT32), .B1(new_n572), .B2(new_n555), .ZN(new_n573));
  NOR2_X1   g387(.A1(new_n568), .A2(new_n573), .ZN(new_n574));
  INV_X1    g388(.A(KEYINPUT32), .ZN(new_n575));
  AOI21_X1  g389(.A(new_n563), .B1(new_n549), .B2(new_n542), .ZN(new_n576));
  AOI21_X1  g390(.A(new_n542), .B1(new_n535), .B2(new_n538), .ZN(new_n577));
  NOR3_X1   g391(.A1(new_n576), .A2(new_n565), .A3(new_n577), .ZN(new_n578));
  OAI211_X1 g392(.A(KEYINPUT72), .B(new_n575), .C1(new_n578), .C2(new_n554), .ZN(new_n579));
  INV_X1    g393(.A(new_n579), .ZN(new_n580));
  OAI21_X1  g394(.A(new_n552), .B1(new_n574), .B2(new_n580), .ZN(new_n581));
  INV_X1    g395(.A(KEYINPUT25), .ZN(new_n582));
  INV_X1    g396(.A(G128), .ZN(new_n583));
  NOR2_X1   g397(.A1(new_n583), .A2(G119), .ZN(new_n584));
  AOI21_X1  g398(.A(new_n584), .B1(new_n204), .B2(G119), .ZN(new_n585));
  XOR2_X1   g399(.A(KEYINPUT24), .B(G110), .Z(new_n586));
  NOR2_X1   g400(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  XOR2_X1   g401(.A(new_n587), .B(KEYINPUT73), .Z(new_n588));
  AOI21_X1  g402(.A(KEYINPUT23), .B1(new_n583), .B2(G119), .ZN(new_n589));
  INV_X1    g403(.A(new_n589), .ZN(new_n590));
  INV_X1    g404(.A(KEYINPUT23), .ZN(new_n591));
  OAI21_X1  g405(.A(new_n590), .B1(new_n585), .B2(new_n591), .ZN(new_n592));
  NOR2_X1   g406(.A1(new_n592), .A2(G110), .ZN(new_n593));
  OAI211_X1 g407(.A(new_n364), .B(new_n412), .C1(new_n588), .C2(new_n593), .ZN(new_n594));
  AOI22_X1  g408(.A1(new_n363), .A2(new_n364), .B1(new_n585), .B2(new_n586), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n592), .A2(G110), .ZN(new_n596));
  NAND2_X1  g410(.A1(new_n595), .A2(new_n596), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n594), .A2(new_n597), .ZN(new_n598));
  XNOR2_X1  g412(.A(KEYINPUT22), .B(G137), .ZN(new_n599));
  XNOR2_X1  g413(.A(new_n599), .B(KEYINPUT75), .ZN(new_n600));
  NAND3_X1  g414(.A1(new_n223), .A2(G221), .A3(G234), .ZN(new_n601));
  XOR2_X1   g415(.A(new_n600), .B(new_n601), .Z(new_n602));
  NAND2_X1  g416(.A1(new_n602), .A2(KEYINPUT76), .ZN(new_n603));
  OR2_X1    g417(.A1(new_n602), .A2(KEYINPUT76), .ZN(new_n604));
  NAND3_X1  g418(.A1(new_n598), .A2(new_n603), .A3(new_n604), .ZN(new_n605));
  NAND4_X1  g419(.A1(new_n594), .A2(new_n597), .A3(KEYINPUT76), .A4(new_n602), .ZN(new_n606));
  NAND2_X1  g420(.A1(new_n605), .A2(new_n606), .ZN(new_n607));
  AOI21_X1  g421(.A(new_n582), .B1(new_n607), .B2(new_n285), .ZN(new_n608));
  INV_X1    g422(.A(new_n608), .ZN(new_n609));
  AOI21_X1  g423(.A(new_n325), .B1(G234), .B2(new_n285), .ZN(new_n610));
  NAND3_X1  g424(.A1(new_n607), .A2(new_n582), .A3(new_n285), .ZN(new_n611));
  NAND3_X1  g425(.A1(new_n609), .A2(new_n610), .A3(new_n611), .ZN(new_n612));
  NOR2_X1   g426(.A1(new_n610), .A2(G902), .ZN(new_n613));
  NAND2_X1  g427(.A1(new_n607), .A2(new_n613), .ZN(new_n614));
  NAND2_X1  g428(.A1(new_n612), .A2(new_n614), .ZN(new_n615));
  INV_X1    g429(.A(new_n615), .ZN(new_n616));
  NAND4_X1  g430(.A1(new_n517), .A2(new_n525), .A3(new_n581), .A4(new_n616), .ZN(new_n617));
  XNOR2_X1  g431(.A(new_n617), .B(G101), .ZN(G3));
  INV_X1    g432(.A(G472), .ZN(new_n619));
  AOI21_X1  g433(.A(new_n619), .B1(new_n572), .B2(new_n285), .ZN(new_n620));
  NOR2_X1   g434(.A1(new_n578), .A2(new_n554), .ZN(new_n621));
  OR2_X1    g435(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  NOR3_X1   g436(.A1(new_n622), .A2(new_n516), .A3(new_n615), .ZN(new_n623));
  INV_X1    g437(.A(new_n189), .ZN(new_n624));
  OAI21_X1  g438(.A(new_n624), .B1(new_n274), .B2(new_n286), .ZN(new_n625));
  AOI21_X1  g439(.A(new_n188), .B1(new_n625), .B2(new_n297), .ZN(new_n626));
  NAND2_X1  g440(.A1(new_n626), .A2(new_n432), .ZN(new_n627));
  NAND3_X1  g441(.A1(new_n331), .A2(new_n285), .A3(new_n333), .ZN(new_n628));
  INV_X1    g442(.A(G478), .ZN(new_n629));
  NAND2_X1  g443(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  XNOR2_X1  g444(.A(new_n630), .B(KEYINPUT92), .ZN(new_n631));
  INV_X1    g445(.A(KEYINPUT33), .ZN(new_n632));
  NAND3_X1  g446(.A1(new_n331), .A2(new_n632), .A3(new_n333), .ZN(new_n633));
  NAND3_X1  g447(.A1(new_n328), .A2(KEYINPUT33), .A3(new_n330), .ZN(new_n634));
  AND2_X1   g448(.A1(new_n633), .A2(new_n634), .ZN(new_n635));
  NAND3_X1  g449(.A1(new_n635), .A2(G478), .A3(new_n285), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n631), .A2(new_n636), .ZN(new_n637));
  NAND2_X1  g451(.A1(new_n391), .A2(new_n425), .ZN(new_n638));
  NAND2_X1  g452(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  NOR2_X1   g453(.A1(new_n627), .A2(new_n639), .ZN(new_n640));
  NAND2_X1  g454(.A1(new_n623), .A2(new_n640), .ZN(new_n641));
  XOR2_X1   g455(.A(KEYINPUT34), .B(G104), .Z(new_n642));
  XNOR2_X1  g456(.A(new_n641), .B(new_n642), .ZN(G6));
  INV_X1    g457(.A(KEYINPUT93), .ZN(new_n644));
  AOI21_X1  g458(.A(new_n644), .B1(new_n408), .B2(KEYINPUT20), .ZN(new_n645));
  AOI21_X1  g459(.A(new_n645), .B1(new_n425), .B2(new_n644), .ZN(new_n646));
  OR2_X1    g460(.A1(new_n646), .A2(KEYINPUT94), .ZN(new_n647));
  NAND2_X1  g461(.A1(new_n646), .A2(KEYINPUT94), .ZN(new_n648));
  NAND4_X1  g462(.A1(new_n647), .A2(new_n648), .A3(new_n391), .A4(new_n342), .ZN(new_n649));
  NOR2_X1   g463(.A1(new_n627), .A2(new_n649), .ZN(new_n650));
  NAND2_X1  g464(.A1(new_n623), .A2(new_n650), .ZN(new_n651));
  XOR2_X1   g465(.A(KEYINPUT35), .B(G107), .Z(new_n652));
  XNOR2_X1  g466(.A(new_n651), .B(new_n652), .ZN(G9));
  AOI211_X1 g467(.A(KEYINPUT25), .B(G902), .C1(new_n605), .C2(new_n606), .ZN(new_n654));
  NOR2_X1   g468(.A1(new_n608), .A2(new_n654), .ZN(new_n655));
  NOR2_X1   g469(.A1(new_n602), .A2(KEYINPUT36), .ZN(new_n656));
  XNOR2_X1  g470(.A(new_n598), .B(new_n656), .ZN(new_n657));
  AOI22_X1  g471(.A1(new_n655), .A2(new_n610), .B1(new_n613), .B2(new_n657), .ZN(new_n658));
  NOR3_X1   g472(.A1(new_n658), .A2(new_n621), .A3(new_n620), .ZN(new_n659));
  NAND3_X1  g473(.A1(new_n517), .A2(new_n525), .A3(new_n659), .ZN(new_n660));
  XNOR2_X1  g474(.A(new_n660), .B(G110), .ZN(new_n661));
  XOR2_X1   g475(.A(KEYINPUT95), .B(KEYINPUT37), .Z(new_n662));
  XNOR2_X1  g476(.A(new_n661), .B(new_n662), .ZN(G12));
  NAND2_X1  g477(.A1(new_n657), .A2(new_n613), .ZN(new_n664));
  NAND2_X1  g478(.A1(new_n612), .A2(new_n664), .ZN(new_n665));
  AND2_X1   g479(.A1(new_n665), .A2(new_n626), .ZN(new_n666));
  OR2_X1    g480(.A1(new_n431), .A2(G900), .ZN(new_n667));
  NAND2_X1  g481(.A1(new_n667), .A2(new_n429), .ZN(new_n668));
  INV_X1    g482(.A(new_n668), .ZN(new_n669));
  NOR2_X1   g483(.A1(new_n649), .A2(new_n669), .ZN(new_n670));
  NAND4_X1  g484(.A1(new_n581), .A2(new_n666), .A3(new_n520), .A4(new_n670), .ZN(new_n671));
  XNOR2_X1  g485(.A(new_n671), .B(G128), .ZN(G30));
  AOI21_X1  g486(.A(new_n542), .B1(new_n558), .B2(new_n536), .ZN(new_n673));
  AOI21_X1  g487(.A(new_n562), .B1(KEYINPUT96), .B2(new_n673), .ZN(new_n674));
  OAI21_X1  g488(.A(new_n674), .B1(KEYINPUT96), .B2(new_n673), .ZN(new_n675));
  AOI21_X1  g489(.A(new_n619), .B1(new_n675), .B2(new_n285), .ZN(new_n676));
  INV_X1    g490(.A(new_n676), .ZN(new_n677));
  OAI21_X1  g491(.A(new_n677), .B1(new_n574), .B2(new_n580), .ZN(new_n678));
  INV_X1    g492(.A(KEYINPUT97), .ZN(new_n679));
  NAND2_X1  g493(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  OAI21_X1  g494(.A(new_n575), .B1(new_n578), .B2(new_n554), .ZN(new_n681));
  NAND3_X1  g495(.A1(new_n681), .A2(new_n567), .A3(new_n566), .ZN(new_n682));
  NAND2_X1  g496(.A1(new_n682), .A2(new_n579), .ZN(new_n683));
  NAND3_X1  g497(.A1(new_n683), .A2(KEYINPUT97), .A3(new_n677), .ZN(new_n684));
  NAND2_X1  g498(.A1(new_n680), .A2(new_n684), .ZN(new_n685));
  AND2_X1   g499(.A1(new_n287), .A2(new_n297), .ZN(new_n686));
  XNOR2_X1  g500(.A(new_n686), .B(KEYINPUT38), .ZN(new_n687));
  NOR3_X1   g501(.A1(new_n687), .A2(new_n188), .A3(new_n665), .ZN(new_n688));
  XOR2_X1   g502(.A(new_n668), .B(KEYINPUT39), .Z(new_n689));
  OAI21_X1  g503(.A(KEYINPUT40), .B1(new_n516), .B2(new_n689), .ZN(new_n690));
  NOR3_X1   g504(.A1(new_n516), .A2(KEYINPUT40), .A3(new_n689), .ZN(new_n691));
  NAND2_X1  g505(.A1(new_n342), .A2(new_n638), .ZN(new_n692));
  NOR2_X1   g506(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  NAND4_X1  g507(.A1(new_n685), .A2(new_n688), .A3(new_n690), .A4(new_n693), .ZN(new_n694));
  XNOR2_X1  g508(.A(new_n694), .B(KEYINPUT98), .ZN(new_n695));
  XNOR2_X1  g509(.A(new_n695), .B(new_n207), .ZN(G45));
  NOR2_X1   g510(.A1(new_n639), .A2(new_n669), .ZN(new_n697));
  NAND4_X1  g511(.A1(new_n581), .A2(new_n666), .A3(new_n520), .A4(new_n697), .ZN(new_n698));
  XNOR2_X1  g512(.A(new_n698), .B(G146), .ZN(G48));
  NAND2_X1  g513(.A1(new_n581), .A2(new_n616), .ZN(new_n700));
  INV_X1    g514(.A(KEYINPUT99), .ZN(new_n701));
  OAI21_X1  g515(.A(new_n503), .B1(new_n498), .B2(new_n499), .ZN(new_n702));
  AND2_X1   g516(.A1(new_n495), .A2(new_n478), .ZN(new_n703));
  OAI21_X1  g517(.A(new_n702), .B1(new_n703), .B2(new_n481), .ZN(new_n704));
  NAND2_X1  g518(.A1(new_n704), .A2(new_n285), .ZN(new_n705));
  NAND2_X1  g519(.A1(new_n705), .A2(G469), .ZN(new_n706));
  NAND2_X1  g520(.A1(new_n706), .A2(new_n497), .ZN(new_n707));
  OAI21_X1  g521(.A(new_n701), .B1(new_n707), .B2(new_n510), .ZN(new_n708));
  NAND4_X1  g522(.A1(new_n706), .A2(KEYINPUT99), .A3(new_n511), .A4(new_n497), .ZN(new_n709));
  AND2_X1   g523(.A1(new_n708), .A2(new_n709), .ZN(new_n710));
  INV_X1    g524(.A(new_n710), .ZN(new_n711));
  NOR2_X1   g525(.A1(new_n700), .A2(new_n711), .ZN(new_n712));
  NAND2_X1  g526(.A1(new_n712), .A2(new_n640), .ZN(new_n713));
  XNOR2_X1  g527(.A(KEYINPUT41), .B(G113), .ZN(new_n714));
  XNOR2_X1  g528(.A(new_n713), .B(new_n714), .ZN(G15));
  NAND2_X1  g529(.A1(new_n712), .A2(new_n650), .ZN(new_n716));
  XNOR2_X1  g530(.A(new_n716), .B(G116), .ZN(G18));
  NAND4_X1  g531(.A1(new_n710), .A2(new_n581), .A3(new_n666), .A4(new_n524), .ZN(new_n718));
  XNOR2_X1  g532(.A(new_n718), .B(G119), .ZN(G21));
  NOR2_X1   g533(.A1(new_n622), .A2(new_n615), .ZN(new_n720));
  INV_X1    g534(.A(KEYINPUT100), .ZN(new_n721));
  INV_X1    g535(.A(new_n638), .ZN(new_n722));
  OAI21_X1  g536(.A(new_n721), .B1(new_n722), .B2(new_n440), .ZN(new_n723));
  NAND3_X1  g537(.A1(new_n342), .A2(KEYINPUT100), .A3(new_n638), .ZN(new_n724));
  NAND2_X1  g538(.A1(new_n723), .A2(new_n724), .ZN(new_n725));
  NOR2_X1   g539(.A1(new_n627), .A2(new_n725), .ZN(new_n726));
  NAND3_X1  g540(.A1(new_n710), .A2(new_n720), .A3(new_n726), .ZN(new_n727));
  XNOR2_X1  g541(.A(new_n727), .B(G122), .ZN(G24));
  NAND4_X1  g542(.A1(new_n710), .A2(new_n659), .A3(new_n626), .A4(new_n697), .ZN(new_n729));
  XNOR2_X1  g543(.A(new_n729), .B(G125), .ZN(G27));
  NAND3_X1  g544(.A1(new_n287), .A2(new_n297), .A3(new_n187), .ZN(new_n731));
  NOR2_X1   g545(.A1(new_n731), .A2(new_n512), .ZN(new_n732));
  NAND3_X1  g546(.A1(new_n552), .A2(new_n681), .A3(new_n566), .ZN(new_n733));
  NAND4_X1  g547(.A1(new_n616), .A2(new_n697), .A3(new_n732), .A4(new_n733), .ZN(new_n734));
  NAND2_X1  g548(.A1(new_n734), .A2(KEYINPUT42), .ZN(new_n735));
  NOR3_X1   g549(.A1(new_n639), .A2(KEYINPUT42), .A3(new_n669), .ZN(new_n736));
  NAND4_X1  g550(.A1(new_n581), .A2(new_n616), .A3(new_n732), .A4(new_n736), .ZN(new_n737));
  AND3_X1   g551(.A1(new_n735), .A2(new_n737), .A3(KEYINPUT101), .ZN(new_n738));
  AOI21_X1  g552(.A(KEYINPUT101), .B1(new_n735), .B2(new_n737), .ZN(new_n739));
  NOR2_X1   g553(.A1(new_n738), .A2(new_n739), .ZN(new_n740));
  XNOR2_X1  g554(.A(new_n740), .B(new_n352), .ZN(G33));
  INV_X1    g555(.A(new_n700), .ZN(new_n742));
  NAND3_X1  g556(.A1(new_n742), .A2(new_n670), .A3(new_n732), .ZN(new_n743));
  XNOR2_X1  g557(.A(new_n743), .B(G134), .ZN(G36));
  AOI22_X1  g558(.A1(new_n500), .A2(new_n501), .B1(new_n503), .B2(new_n495), .ZN(new_n745));
  OAI21_X1  g559(.A(G469), .B1(new_n745), .B2(KEYINPUT45), .ZN(new_n746));
  INV_X1    g560(.A(KEYINPUT102), .ZN(new_n747));
  NAND2_X1  g561(.A1(new_n746), .A2(new_n747), .ZN(new_n748));
  NAND2_X1  g562(.A1(new_n745), .A2(KEYINPUT45), .ZN(new_n749));
  OAI211_X1 g563(.A(KEYINPUT102), .B(G469), .C1(new_n745), .C2(KEYINPUT45), .ZN(new_n750));
  NAND3_X1  g564(.A1(new_n748), .A2(new_n749), .A3(new_n750), .ZN(new_n751));
  NAND2_X1  g565(.A1(new_n751), .A2(new_n506), .ZN(new_n752));
  INV_X1    g566(.A(KEYINPUT46), .ZN(new_n753));
  NAND2_X1  g567(.A1(new_n752), .A2(new_n753), .ZN(new_n754));
  NAND3_X1  g568(.A1(new_n751), .A2(KEYINPUT46), .A3(new_n506), .ZN(new_n755));
  NAND3_X1  g569(.A1(new_n754), .A2(new_n497), .A3(new_n755), .ZN(new_n756));
  NAND2_X1  g570(.A1(new_n756), .A2(new_n511), .ZN(new_n757));
  INV_X1    g571(.A(KEYINPUT103), .ZN(new_n758));
  OR3_X1    g572(.A1(new_n757), .A2(new_n758), .A3(new_n689), .ZN(new_n759));
  AOI21_X1  g573(.A(new_n638), .B1(new_n631), .B2(new_n636), .ZN(new_n760));
  INV_X1    g574(.A(new_n760), .ZN(new_n761));
  INV_X1    g575(.A(KEYINPUT104), .ZN(new_n762));
  NOR2_X1   g576(.A1(new_n762), .A2(KEYINPUT43), .ZN(new_n763));
  NAND2_X1  g577(.A1(new_n761), .A2(new_n763), .ZN(new_n764));
  AOI21_X1  g578(.A(new_n760), .B1(new_n762), .B2(KEYINPUT43), .ZN(new_n765));
  OAI21_X1  g579(.A(new_n764), .B1(new_n765), .B2(new_n763), .ZN(new_n766));
  NAND3_X1  g580(.A1(new_n766), .A2(new_n622), .A3(new_n665), .ZN(new_n767));
  INV_X1    g581(.A(KEYINPUT44), .ZN(new_n768));
  AOI21_X1  g582(.A(new_n731), .B1(new_n767), .B2(new_n768), .ZN(new_n769));
  OR2_X1    g583(.A1(new_n767), .A2(new_n768), .ZN(new_n770));
  OAI21_X1  g584(.A(new_n758), .B1(new_n757), .B2(new_n689), .ZN(new_n771));
  NAND4_X1  g585(.A1(new_n759), .A2(new_n769), .A3(new_n770), .A4(new_n771), .ZN(new_n772));
  XNOR2_X1  g586(.A(new_n772), .B(G137), .ZN(G39));
  INV_X1    g587(.A(KEYINPUT105), .ZN(new_n774));
  OAI21_X1  g588(.A(new_n757), .B1(new_n774), .B2(KEYINPUT47), .ZN(new_n775));
  INV_X1    g589(.A(new_n731), .ZN(new_n776));
  XOR2_X1   g590(.A(KEYINPUT105), .B(KEYINPUT47), .Z(new_n777));
  NAND3_X1  g591(.A1(new_n756), .A2(new_n511), .A3(new_n777), .ZN(new_n778));
  NAND4_X1  g592(.A1(new_n775), .A2(new_n697), .A3(new_n776), .A4(new_n778), .ZN(new_n779));
  NAND3_X1  g593(.A1(new_n683), .A2(new_n552), .A3(new_n615), .ZN(new_n780));
  NOR2_X1   g594(.A1(new_n779), .A2(new_n780), .ZN(new_n781));
  XNOR2_X1  g595(.A(new_n781), .B(new_n356), .ZN(G42));
  NAND2_X1  g596(.A1(new_n426), .A2(new_n223), .ZN(new_n783));
  AND3_X1   g597(.A1(new_n647), .A2(new_n648), .A3(new_n391), .ZN(new_n784));
  NAND4_X1  g598(.A1(new_n581), .A2(new_n520), .A3(new_n440), .A4(new_n784), .ZN(new_n785));
  OR3_X1    g599(.A1(new_n622), .A2(new_n512), .A3(new_n639), .ZN(new_n786));
  NAND2_X1  g600(.A1(new_n785), .A2(new_n786), .ZN(new_n787));
  NAND4_X1  g601(.A1(new_n787), .A2(new_n665), .A3(new_n668), .A4(new_n776), .ZN(new_n788));
  NAND2_X1  g602(.A1(new_n788), .A2(new_n743), .ZN(new_n789));
  NAND4_X1  g603(.A1(new_n713), .A2(new_n716), .A3(new_n718), .A4(new_n727), .ZN(new_n790));
  NOR3_X1   g604(.A1(new_n686), .A2(new_n639), .A3(new_n188), .ZN(new_n791));
  NAND4_X1  g605(.A1(new_n720), .A2(new_n791), .A3(new_n520), .A4(new_n432), .ZN(new_n792));
  NAND2_X1  g606(.A1(new_n617), .A2(new_n792), .ZN(new_n793));
  INV_X1    g607(.A(KEYINPUT106), .ZN(new_n794));
  NAND2_X1  g608(.A1(new_n793), .A2(new_n794), .ZN(new_n795));
  NOR2_X1   g609(.A1(new_n440), .A2(new_n638), .ZN(new_n796));
  INV_X1    g610(.A(KEYINPUT107), .ZN(new_n797));
  XNOR2_X1  g611(.A(new_n796), .B(new_n797), .ZN(new_n798));
  NAND4_X1  g612(.A1(new_n623), .A2(new_n298), .A3(new_n432), .A4(new_n798), .ZN(new_n799));
  AND2_X1   g613(.A1(new_n799), .A2(new_n660), .ZN(new_n800));
  NAND3_X1  g614(.A1(new_n617), .A2(KEYINPUT106), .A3(new_n792), .ZN(new_n801));
  NAND3_X1  g615(.A1(new_n795), .A2(new_n800), .A3(new_n801), .ZN(new_n802));
  NAND2_X1  g616(.A1(new_n802), .A2(KEYINPUT108), .ZN(new_n803));
  INV_X1    g617(.A(KEYINPUT108), .ZN(new_n804));
  NAND4_X1  g618(.A1(new_n795), .A2(new_n800), .A3(new_n804), .A4(new_n801), .ZN(new_n805));
  AOI211_X1 g619(.A(new_n789), .B(new_n790), .C1(new_n803), .C2(new_n805), .ZN(new_n806));
  AND3_X1   g620(.A1(new_n729), .A2(new_n671), .A3(new_n698), .ZN(new_n807));
  INV_X1    g621(.A(KEYINPUT109), .ZN(new_n808));
  NAND3_X1  g622(.A1(new_n626), .A2(new_n723), .A3(new_n724), .ZN(new_n809));
  NOR4_X1   g623(.A1(new_n809), .A2(new_n665), .A3(new_n512), .A4(new_n669), .ZN(new_n810));
  AOI21_X1  g624(.A(new_n808), .B1(new_n685), .B2(new_n810), .ZN(new_n811));
  AOI21_X1  g625(.A(KEYINPUT97), .B1(new_n683), .B2(new_n677), .ZN(new_n812));
  AOI211_X1 g626(.A(new_n679), .B(new_n676), .C1(new_n682), .C2(new_n579), .ZN(new_n813));
  OAI211_X1 g627(.A(new_n810), .B(new_n808), .C1(new_n812), .C2(new_n813), .ZN(new_n814));
  INV_X1    g628(.A(new_n814), .ZN(new_n815));
  OAI21_X1  g629(.A(new_n807), .B1(new_n811), .B2(new_n815), .ZN(new_n816));
  INV_X1    g630(.A(KEYINPUT110), .ZN(new_n817));
  NAND2_X1  g631(.A1(new_n816), .A2(new_n817), .ZN(new_n818));
  INV_X1    g632(.A(KEYINPUT52), .ZN(new_n819));
  OAI21_X1  g633(.A(new_n810), .B1(new_n812), .B2(new_n813), .ZN(new_n820));
  NAND2_X1  g634(.A1(new_n820), .A2(KEYINPUT109), .ZN(new_n821));
  NAND2_X1  g635(.A1(new_n821), .A2(new_n814), .ZN(new_n822));
  NAND3_X1  g636(.A1(new_n822), .A2(KEYINPUT110), .A3(new_n807), .ZN(new_n823));
  NAND3_X1  g637(.A1(new_n818), .A2(new_n819), .A3(new_n823), .ZN(new_n824));
  NAND3_X1  g638(.A1(new_n822), .A2(KEYINPUT52), .A3(new_n807), .ZN(new_n825));
  NAND2_X1  g639(.A1(new_n824), .A2(new_n825), .ZN(new_n826));
  AND3_X1   g640(.A1(new_n735), .A2(new_n737), .A3(KEYINPUT53), .ZN(new_n827));
  AND3_X1   g641(.A1(new_n806), .A2(new_n826), .A3(new_n827), .ZN(new_n828));
  OAI211_X1 g642(.A(new_n788), .B(new_n743), .C1(new_n739), .C2(new_n738), .ZN(new_n829));
  AOI211_X1 g643(.A(new_n790), .B(new_n829), .C1(new_n803), .C2(new_n805), .ZN(new_n830));
  NAND3_X1  g644(.A1(new_n729), .A2(new_n671), .A3(new_n698), .ZN(new_n831));
  AOI211_X1 g645(.A(new_n817), .B(new_n831), .C1(new_n821), .C2(new_n814), .ZN(new_n832));
  AOI21_X1  g646(.A(KEYINPUT110), .B1(new_n822), .B2(new_n807), .ZN(new_n833));
  OAI21_X1  g647(.A(KEYINPUT52), .B1(new_n832), .B2(new_n833), .ZN(new_n834));
  NAND2_X1  g648(.A1(new_n834), .A2(new_n824), .ZN(new_n835));
  AOI21_X1  g649(.A(KEYINPUT53), .B1(new_n830), .B2(new_n835), .ZN(new_n836));
  XOR2_X1   g650(.A(KEYINPUT112), .B(KEYINPUT54), .Z(new_n837));
  NOR3_X1   g651(.A1(new_n828), .A2(new_n836), .A3(new_n837), .ZN(new_n838));
  INV_X1    g652(.A(KEYINPUT53), .ZN(new_n839));
  AND2_X1   g653(.A1(new_n824), .A2(new_n825), .ZN(new_n840));
  INV_X1    g654(.A(new_n829), .ZN(new_n841));
  INV_X1    g655(.A(new_n790), .ZN(new_n842));
  AND3_X1   g656(.A1(new_n617), .A2(KEYINPUT106), .A3(new_n792), .ZN(new_n843));
  AOI21_X1  g657(.A(KEYINPUT106), .B1(new_n617), .B2(new_n792), .ZN(new_n844));
  NOR2_X1   g658(.A1(new_n843), .A2(new_n844), .ZN(new_n845));
  AOI21_X1  g659(.A(new_n804), .B1(new_n845), .B2(new_n800), .ZN(new_n846));
  INV_X1    g660(.A(new_n805), .ZN(new_n847));
  OAI211_X1 g661(.A(new_n841), .B(new_n842), .C1(new_n846), .C2(new_n847), .ZN(new_n848));
  OAI21_X1  g662(.A(new_n839), .B1(new_n840), .B2(new_n848), .ZN(new_n849));
  NAND2_X1  g663(.A1(new_n849), .A2(KEYINPUT111), .ZN(new_n850));
  AOI21_X1  g664(.A(new_n848), .B1(new_n824), .B2(new_n834), .ZN(new_n851));
  NAND2_X1  g665(.A1(new_n851), .A2(KEYINPUT53), .ZN(new_n852));
  INV_X1    g666(.A(KEYINPUT111), .ZN(new_n853));
  OAI211_X1 g667(.A(new_n853), .B(new_n839), .C1(new_n840), .C2(new_n848), .ZN(new_n854));
  NAND3_X1  g668(.A1(new_n850), .A2(new_n852), .A3(new_n854), .ZN(new_n855));
  AOI21_X1  g669(.A(new_n838), .B1(new_n855), .B2(KEYINPUT54), .ZN(new_n856));
  INV_X1    g670(.A(new_n685), .ZN(new_n857));
  INV_X1    g671(.A(new_n429), .ZN(new_n858));
  NOR2_X1   g672(.A1(new_n711), .A2(new_n731), .ZN(new_n859));
  NAND4_X1  g673(.A1(new_n857), .A2(new_n616), .A3(new_n858), .A4(new_n859), .ZN(new_n860));
  OR2_X1    g674(.A1(new_n860), .A2(new_n639), .ZN(new_n861));
  NAND2_X1  g675(.A1(new_n766), .A2(new_n858), .ZN(new_n862));
  XOR2_X1   g676(.A(new_n862), .B(KEYINPUT113), .Z(new_n863));
  AND2_X1   g677(.A1(new_n863), .A2(new_n720), .ZN(new_n864));
  NAND3_X1  g678(.A1(new_n864), .A2(new_n626), .A3(new_n710), .ZN(new_n865));
  INV_X1    g679(.A(KEYINPUT51), .ZN(new_n866));
  NOR2_X1   g680(.A1(new_n711), .A2(new_n187), .ZN(new_n867));
  OAI211_X1 g681(.A(new_n863), .B(new_n720), .C1(KEYINPUT114), .C2(new_n867), .ZN(new_n868));
  NAND2_X1  g682(.A1(new_n867), .A2(KEYINPUT114), .ZN(new_n869));
  NAND2_X1  g683(.A1(new_n869), .A2(new_n687), .ZN(new_n870));
  OR3_X1    g684(.A1(new_n868), .A2(KEYINPUT50), .A3(new_n870), .ZN(new_n871));
  AND3_X1   g685(.A1(new_n863), .A2(KEYINPUT115), .A3(new_n859), .ZN(new_n872));
  AOI21_X1  g686(.A(KEYINPUT115), .B1(new_n863), .B2(new_n859), .ZN(new_n873));
  OAI21_X1  g687(.A(new_n659), .B1(new_n872), .B2(new_n873), .ZN(new_n874));
  OAI21_X1  g688(.A(KEYINPUT50), .B1(new_n868), .B2(new_n870), .ZN(new_n875));
  OR3_X1    g689(.A1(new_n860), .A2(new_n638), .A3(new_n637), .ZN(new_n876));
  NAND4_X1  g690(.A1(new_n871), .A2(new_n874), .A3(new_n875), .A4(new_n876), .ZN(new_n877));
  NAND2_X1  g691(.A1(new_n775), .A2(new_n778), .ZN(new_n878));
  OAI21_X1  g692(.A(new_n878), .B1(new_n511), .B2(new_n707), .ZN(new_n879));
  AND3_X1   g693(.A1(new_n864), .A2(new_n776), .A3(new_n879), .ZN(new_n880));
  OAI21_X1  g694(.A(new_n866), .B1(new_n877), .B2(new_n880), .ZN(new_n881));
  NAND2_X1  g695(.A1(new_n881), .A2(new_n427), .ZN(new_n882));
  OR2_X1    g696(.A1(new_n879), .A2(KEYINPUT116), .ZN(new_n883));
  NAND2_X1  g697(.A1(new_n879), .A2(KEYINPUT116), .ZN(new_n884));
  AND4_X1   g698(.A1(new_n776), .A2(new_n883), .A3(new_n864), .A4(new_n884), .ZN(new_n885));
  NOR3_X1   g699(.A1(new_n877), .A2(new_n885), .A3(new_n866), .ZN(new_n886));
  NOR2_X1   g700(.A1(new_n882), .A2(new_n886), .ZN(new_n887));
  NAND4_X1  g701(.A1(new_n856), .A2(new_n861), .A3(new_n865), .A4(new_n887), .ZN(new_n888));
  AND2_X1   g702(.A1(new_n616), .A2(new_n733), .ZN(new_n889));
  OAI21_X1  g703(.A(new_n889), .B1(new_n872), .B2(new_n873), .ZN(new_n890));
  XOR2_X1   g704(.A(new_n890), .B(KEYINPUT48), .Z(new_n891));
  OAI21_X1  g705(.A(new_n783), .B1(new_n888), .B2(new_n891), .ZN(new_n892));
  XNOR2_X1  g706(.A(new_n707), .B(KEYINPUT49), .ZN(new_n893));
  NOR3_X1   g707(.A1(new_n893), .A2(new_n615), .A3(new_n188), .ZN(new_n894));
  AND3_X1   g708(.A1(new_n687), .A2(new_n511), .A3(new_n760), .ZN(new_n895));
  NAND3_X1  g709(.A1(new_n857), .A2(new_n894), .A3(new_n895), .ZN(new_n896));
  NAND2_X1  g710(.A1(new_n892), .A2(new_n896), .ZN(G75));
  XNOR2_X1  g711(.A(new_n293), .B(new_n227), .ZN(new_n898));
  XNOR2_X1  g712(.A(new_n898), .B(KEYINPUT55), .ZN(new_n899));
  NOR2_X1   g713(.A1(new_n828), .A2(new_n836), .ZN(new_n900));
  NOR2_X1   g714(.A1(new_n900), .A2(new_n285), .ZN(new_n901));
  NAND2_X1  g715(.A1(new_n901), .A2(G210), .ZN(new_n902));
  INV_X1    g716(.A(KEYINPUT56), .ZN(new_n903));
  AOI21_X1  g717(.A(new_n899), .B1(new_n902), .B2(new_n903), .ZN(new_n904));
  NOR2_X1   g718(.A1(new_n223), .A2(G952), .ZN(new_n905));
  NAND2_X1  g719(.A1(new_n899), .A2(new_n903), .ZN(new_n906));
  AOI21_X1  g720(.A(new_n906), .B1(new_n901), .B2(new_n191), .ZN(new_n907));
  NOR3_X1   g721(.A1(new_n904), .A2(new_n905), .A3(new_n907), .ZN(G51));
  OAI21_X1  g722(.A(new_n837), .B1(new_n828), .B2(new_n836), .ZN(new_n909));
  INV_X1    g723(.A(new_n837), .ZN(new_n910));
  NAND3_X1  g724(.A1(new_n806), .A2(new_n826), .A3(new_n827), .ZN(new_n911));
  OAI211_X1 g725(.A(new_n910), .B(new_n911), .C1(new_n851), .C2(KEYINPUT53), .ZN(new_n912));
  NAND3_X1  g726(.A1(new_n909), .A2(KEYINPUT117), .A3(new_n912), .ZN(new_n913));
  INV_X1    g727(.A(KEYINPUT117), .ZN(new_n914));
  OAI211_X1 g728(.A(new_n914), .B(new_n837), .C1(new_n828), .C2(new_n836), .ZN(new_n915));
  XOR2_X1   g729(.A(new_n506), .B(KEYINPUT57), .Z(new_n916));
  NAND3_X1  g730(.A1(new_n913), .A2(new_n915), .A3(new_n916), .ZN(new_n917));
  NAND2_X1  g731(.A1(new_n917), .A2(KEYINPUT118), .ZN(new_n918));
  INV_X1    g732(.A(KEYINPUT118), .ZN(new_n919));
  NAND4_X1  g733(.A1(new_n913), .A2(new_n919), .A3(new_n915), .A4(new_n916), .ZN(new_n920));
  XOR2_X1   g734(.A(new_n704), .B(KEYINPUT119), .Z(new_n921));
  NAND3_X1  g735(.A1(new_n918), .A2(new_n920), .A3(new_n921), .ZN(new_n922));
  OR3_X1    g736(.A1(new_n900), .A2(new_n285), .A3(new_n751), .ZN(new_n923));
  AOI21_X1  g737(.A(new_n905), .B1(new_n922), .B2(new_n923), .ZN(G54));
  NAND3_X1  g738(.A1(new_n901), .A2(KEYINPUT58), .A3(G475), .ZN(new_n925));
  INV_X1    g739(.A(new_n422), .ZN(new_n926));
  AND2_X1   g740(.A1(new_n925), .A2(new_n926), .ZN(new_n927));
  NOR2_X1   g741(.A1(new_n925), .A2(new_n926), .ZN(new_n928));
  NOR3_X1   g742(.A1(new_n927), .A2(new_n928), .A3(new_n905), .ZN(G60));
  INV_X1    g743(.A(new_n635), .ZN(new_n930));
  NAND2_X1  g744(.A1(G478), .A2(G902), .ZN(new_n931));
  XOR2_X1   g745(.A(new_n931), .B(KEYINPUT59), .Z(new_n932));
  OAI21_X1  g746(.A(new_n930), .B1(new_n856), .B2(new_n932), .ZN(new_n933));
  INV_X1    g747(.A(new_n905), .ZN(new_n934));
  INV_X1    g748(.A(new_n932), .ZN(new_n935));
  NAND4_X1  g749(.A1(new_n913), .A2(new_n635), .A3(new_n915), .A4(new_n935), .ZN(new_n936));
  AND3_X1   g750(.A1(new_n933), .A2(new_n934), .A3(new_n936), .ZN(G63));
  XNOR2_X1  g751(.A(KEYINPUT120), .B(KEYINPUT60), .ZN(new_n938));
  NAND2_X1  g752(.A1(G217), .A2(G902), .ZN(new_n939));
  XNOR2_X1  g753(.A(new_n938), .B(new_n939), .ZN(new_n940));
  NOR2_X1   g754(.A1(new_n900), .A2(new_n940), .ZN(new_n941));
  NAND2_X1  g755(.A1(new_n941), .A2(new_n657), .ZN(new_n942));
  XNOR2_X1  g756(.A(new_n607), .B(KEYINPUT121), .ZN(new_n943));
  INV_X1    g757(.A(new_n943), .ZN(new_n944));
  OAI211_X1 g758(.A(new_n942), .B(new_n934), .C1(new_n941), .C2(new_n944), .ZN(new_n945));
  INV_X1    g759(.A(KEYINPUT61), .ZN(new_n946));
  XNOR2_X1  g760(.A(new_n945), .B(new_n946), .ZN(G66));
  INV_X1    g761(.A(new_n430), .ZN(new_n948));
  OAI21_X1  g762(.A(G953), .B1(new_n948), .B2(new_n221), .ZN(new_n949));
  AOI21_X1  g763(.A(new_n790), .B1(new_n803), .B2(new_n805), .ZN(new_n950));
  OAI21_X1  g764(.A(new_n949), .B1(new_n950), .B2(G953), .ZN(new_n951));
  XNOR2_X1  g765(.A(new_n951), .B(KEYINPUT122), .ZN(new_n952));
  OAI211_X1 g766(.A(new_n272), .B(new_n273), .C1(G898), .C2(new_n223), .ZN(new_n953));
  XNOR2_X1  g767(.A(new_n952), .B(new_n953), .ZN(G69));
  XNOR2_X1  g768(.A(new_n548), .B(new_n419), .ZN(new_n955));
  OAI211_X1 g769(.A(new_n772), .B(new_n743), .C1(new_n780), .C2(new_n779), .ZN(new_n956));
  INV_X1    g770(.A(new_n956), .ZN(new_n957));
  NAND2_X1  g771(.A1(new_n807), .A2(KEYINPUT123), .ZN(new_n958));
  INV_X1    g772(.A(KEYINPUT123), .ZN(new_n959));
  NAND2_X1  g773(.A1(new_n831), .A2(new_n959), .ZN(new_n960));
  NAND2_X1  g774(.A1(new_n958), .A2(new_n960), .ZN(new_n961));
  NOR2_X1   g775(.A1(new_n961), .A2(new_n740), .ZN(new_n962));
  NAND3_X1  g776(.A1(new_n759), .A2(new_n889), .A3(new_n771), .ZN(new_n963));
  OAI211_X1 g777(.A(new_n957), .B(new_n962), .C1(new_n809), .C2(new_n963), .ZN(new_n964));
  OAI21_X1  g778(.A(new_n955), .B1(new_n964), .B2(G953), .ZN(new_n965));
  AOI21_X1  g779(.A(new_n965), .B1(G900), .B2(G953), .ZN(new_n966));
  INV_X1    g780(.A(new_n798), .ZN(new_n967));
  NAND2_X1  g781(.A1(new_n967), .A2(new_n639), .ZN(new_n968));
  NOR3_X1   g782(.A1(new_n516), .A2(new_n689), .A3(new_n731), .ZN(new_n969));
  NAND3_X1  g783(.A1(new_n742), .A2(new_n968), .A3(new_n969), .ZN(new_n970));
  OAI211_X1 g784(.A(new_n772), .B(new_n970), .C1(new_n780), .C2(new_n779), .ZN(new_n971));
  NAND3_X1  g785(.A1(new_n958), .A2(new_n694), .A3(new_n960), .ZN(new_n972));
  INV_X1    g786(.A(KEYINPUT62), .ZN(new_n973));
  OR2_X1    g787(.A1(new_n972), .A2(new_n973), .ZN(new_n974));
  NAND2_X1  g788(.A1(new_n972), .A2(new_n973), .ZN(new_n975));
  AOI21_X1  g789(.A(new_n971), .B1(new_n974), .B2(new_n975), .ZN(new_n976));
  INV_X1    g790(.A(new_n976), .ZN(new_n977));
  AOI21_X1  g791(.A(new_n955), .B1(new_n977), .B2(new_n223), .ZN(new_n978));
  NOR3_X1   g792(.A1(new_n966), .A2(KEYINPUT124), .A3(new_n978), .ZN(new_n979));
  AOI21_X1  g793(.A(new_n223), .B1(G227), .B2(G900), .ZN(new_n980));
  XOR2_X1   g794(.A(new_n979), .B(new_n980), .Z(G72));
  NAND2_X1  g795(.A1(G472), .A2(G902), .ZN(new_n982));
  XOR2_X1   g796(.A(new_n982), .B(KEYINPUT63), .Z(new_n983));
  INV_X1    g797(.A(new_n950), .ZN(new_n984));
  OAI21_X1  g798(.A(new_n983), .B1(new_n964), .B2(new_n984), .ZN(new_n985));
  NAND3_X1  g799(.A1(new_n985), .A2(new_n556), .A3(new_n549), .ZN(new_n986));
  INV_X1    g800(.A(new_n983), .ZN(new_n987));
  AOI21_X1  g801(.A(new_n987), .B1(new_n976), .B2(new_n950), .ZN(new_n988));
  INV_X1    g802(.A(KEYINPUT125), .ZN(new_n989));
  NAND2_X1  g803(.A1(new_n988), .A2(new_n989), .ZN(new_n990));
  NAND2_X1  g804(.A1(new_n990), .A2(new_n542), .ZN(new_n991));
  OAI22_X1  g805(.A1(new_n988), .A2(new_n989), .B1(new_n530), .B2(new_n561), .ZN(new_n992));
  OAI211_X1 g806(.A(new_n934), .B(new_n986), .C1(new_n991), .C2(new_n992), .ZN(new_n993));
  INV_X1    g807(.A(new_n993), .ZN(new_n994));
  NOR2_X1   g808(.A1(new_n549), .A2(new_n542), .ZN(new_n995));
  XNOR2_X1  g809(.A(new_n995), .B(KEYINPUT126), .ZN(new_n996));
  OAI211_X1 g810(.A(new_n855), .B(new_n983), .C1(new_n562), .C2(new_n996), .ZN(new_n997));
  NAND2_X1  g811(.A1(new_n994), .A2(new_n997), .ZN(new_n998));
  NAND2_X1  g812(.A1(new_n998), .A2(KEYINPUT127), .ZN(new_n999));
  INV_X1    g813(.A(KEYINPUT127), .ZN(new_n1000));
  NAND3_X1  g814(.A1(new_n994), .A2(new_n1000), .A3(new_n997), .ZN(new_n1001));
  NAND2_X1  g815(.A1(new_n999), .A2(new_n1001), .ZN(G57));
endmodule


