//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 1 0 1 1 0 1 1 1 1 1 1 1 0 1 1 1 1 1 1 1 1 0 0 0 0 0 0 0 0 1 1 1 1 1 0 0 1 1 1 1 0 1 1 1 1 1 0 1 0 0 0 1 1 0 0 1 0 0 0 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:20:56 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n682, new_n683, new_n684, new_n685, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n710,
    new_n711, new_n712, new_n713, new_n714, new_n715, new_n716, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n750, new_n751, new_n752, new_n753, new_n755, new_n756, new_n757,
    new_n758, new_n759, new_n760, new_n761, new_n762, new_n763, new_n764,
    new_n766, new_n768, new_n769, new_n770, new_n771, new_n772, new_n773,
    new_n774, new_n775, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n786, new_n787, new_n788, new_n789,
    new_n790, new_n791, new_n792, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n850, new_n851, new_n852, new_n854, new_n855, new_n856,
    new_n858, new_n859, new_n860, new_n861, new_n862, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n902,
    new_n903, new_n904, new_n906, new_n907, new_n908, new_n909, new_n910,
    new_n911, new_n912, new_n913, new_n914, new_n915, new_n916, new_n917,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n930, new_n931, new_n932, new_n933,
    new_n935, new_n936, new_n937, new_n939, new_n940, new_n941, new_n942,
    new_n943, new_n945, new_n946, new_n947, new_n948, new_n949, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n957, new_n958, new_n959,
    new_n960, new_n961, new_n962, new_n963, new_n964, new_n965, new_n966,
    new_n967, new_n968, new_n969, new_n970, new_n971, new_n972, new_n974,
    new_n975, new_n976;
  INV_X1    g000(.A(G64gat), .ZN(new_n202));
  NAND3_X1  g001(.A1(new_n202), .A2(KEYINPUT100), .A3(G57gat), .ZN(new_n203));
  INV_X1    g002(.A(KEYINPUT9), .ZN(new_n204));
  NOR3_X1   g003(.A1(new_n204), .A2(G71gat), .A3(G78gat), .ZN(new_n205));
  NAND2_X1  g004(.A1(G71gat), .A2(G78gat), .ZN(new_n206));
  INV_X1    g005(.A(new_n206), .ZN(new_n207));
  OAI21_X1  g006(.A(new_n203), .B1(new_n205), .B2(new_n207), .ZN(new_n208));
  NAND2_X1  g007(.A1(new_n202), .A2(G57gat), .ZN(new_n209));
  INV_X1    g008(.A(G57gat), .ZN(new_n210));
  NAND2_X1  g009(.A1(new_n210), .A2(G64gat), .ZN(new_n211));
  INV_X1    g010(.A(KEYINPUT100), .ZN(new_n212));
  AND3_X1   g011(.A1(new_n209), .A2(new_n211), .A3(new_n212), .ZN(new_n213));
  AOI21_X1  g012(.A(new_n204), .B1(new_n209), .B2(new_n211), .ZN(new_n214));
  OR2_X1    g013(.A1(G71gat), .A2(G78gat), .ZN(new_n215));
  NAND2_X1  g014(.A1(new_n215), .A2(new_n206), .ZN(new_n216));
  OAI22_X1  g015(.A1(new_n208), .A2(new_n213), .B1(new_n214), .B2(new_n216), .ZN(new_n217));
  INV_X1    g016(.A(KEYINPUT21), .ZN(new_n218));
  NAND2_X1  g017(.A1(new_n217), .A2(new_n218), .ZN(new_n219));
  NAND2_X1  g018(.A1(G231gat), .A2(G233gat), .ZN(new_n220));
  XNOR2_X1  g019(.A(new_n219), .B(new_n220), .ZN(new_n221));
  XNOR2_X1  g020(.A(new_n221), .B(G127gat), .ZN(new_n222));
  XNOR2_X1  g021(.A(G15gat), .B(G22gat), .ZN(new_n223));
  INV_X1    g022(.A(G1gat), .ZN(new_n224));
  NAND2_X1  g023(.A1(new_n224), .A2(KEYINPUT16), .ZN(new_n225));
  AND2_X1   g024(.A1(new_n223), .A2(new_n225), .ZN(new_n226));
  NOR2_X1   g025(.A1(new_n223), .A2(G1gat), .ZN(new_n227));
  OAI21_X1  g026(.A(G8gat), .B1(new_n226), .B2(new_n227), .ZN(new_n228));
  OR2_X1    g027(.A1(new_n223), .A2(G1gat), .ZN(new_n229));
  INV_X1    g028(.A(G8gat), .ZN(new_n230));
  NAND2_X1  g029(.A1(new_n223), .A2(new_n225), .ZN(new_n231));
  NAND3_X1  g030(.A1(new_n229), .A2(new_n230), .A3(new_n231), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n228), .A2(new_n232), .ZN(new_n233));
  INV_X1    g032(.A(new_n233), .ZN(new_n234));
  OAI21_X1  g033(.A(new_n234), .B1(new_n218), .B2(new_n217), .ZN(new_n235));
  XNOR2_X1  g034(.A(new_n222), .B(new_n235), .ZN(new_n236));
  XNOR2_X1  g035(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n237));
  XNOR2_X1  g036(.A(new_n237), .B(KEYINPUT101), .ZN(new_n238));
  XNOR2_X1  g037(.A(new_n238), .B(G155gat), .ZN(new_n239));
  XNOR2_X1  g038(.A(G183gat), .B(G211gat), .ZN(new_n240));
  XNOR2_X1  g039(.A(new_n240), .B(KEYINPUT102), .ZN(new_n241));
  XNOR2_X1  g040(.A(new_n239), .B(new_n241), .ZN(new_n242));
  XNOR2_X1  g041(.A(new_n236), .B(new_n242), .ZN(new_n243));
  INV_X1    g042(.A(new_n243), .ZN(new_n244));
  INV_X1    g043(.A(KEYINPUT17), .ZN(new_n245));
  XNOR2_X1  g044(.A(G43gat), .B(G50gat), .ZN(new_n246));
  NAND2_X1  g045(.A1(new_n246), .A2(KEYINPUT15), .ZN(new_n247));
  NAND2_X1  g046(.A1(G29gat), .A2(G36gat), .ZN(new_n248));
  XNOR2_X1  g047(.A(new_n248), .B(KEYINPUT95), .ZN(new_n249));
  NAND2_X1  g048(.A1(new_n247), .A2(new_n249), .ZN(new_n250));
  INV_X1    g049(.A(KEYINPUT14), .ZN(new_n251));
  INV_X1    g050(.A(G29gat), .ZN(new_n252));
  INV_X1    g051(.A(G36gat), .ZN(new_n253));
  NAND3_X1  g052(.A1(new_n251), .A2(new_n252), .A3(new_n253), .ZN(new_n254));
  OAI21_X1  g053(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n255));
  NAND2_X1  g054(.A1(new_n254), .A2(new_n255), .ZN(new_n256));
  OAI21_X1  g055(.A(new_n256), .B1(KEYINPUT15), .B2(new_n246), .ZN(new_n257));
  NOR2_X1   g056(.A1(new_n250), .A2(new_n257), .ZN(new_n258));
  NAND2_X1  g057(.A1(new_n255), .A2(KEYINPUT94), .ZN(new_n259));
  INV_X1    g058(.A(KEYINPUT94), .ZN(new_n260));
  OAI211_X1 g059(.A(new_n260), .B(KEYINPUT14), .C1(G29gat), .C2(G36gat), .ZN(new_n261));
  NAND3_X1  g060(.A1(new_n259), .A2(new_n261), .A3(new_n254), .ZN(new_n262));
  AOI21_X1  g061(.A(new_n247), .B1(new_n262), .B2(new_n248), .ZN(new_n263));
  OAI21_X1  g062(.A(new_n245), .B1(new_n258), .B2(new_n263), .ZN(new_n264));
  NAND2_X1  g063(.A1(new_n262), .A2(new_n248), .ZN(new_n265));
  NAND3_X1  g064(.A1(new_n265), .A2(KEYINPUT15), .A3(new_n246), .ZN(new_n266));
  OR2_X1    g065(.A1(new_n246), .A2(KEYINPUT15), .ZN(new_n267));
  NAND4_X1  g066(.A1(new_n267), .A2(new_n247), .A3(new_n249), .A4(new_n256), .ZN(new_n268));
  NAND3_X1  g067(.A1(new_n266), .A2(KEYINPUT17), .A3(new_n268), .ZN(new_n269));
  NAND2_X1  g068(.A1(G99gat), .A2(G106gat), .ZN(new_n270));
  NAND2_X1  g069(.A1(new_n270), .A2(KEYINPUT8), .ZN(new_n271));
  NAND2_X1  g070(.A1(G85gat), .A2(G92gat), .ZN(new_n272));
  INV_X1    g071(.A(KEYINPUT7), .ZN(new_n273));
  NAND2_X1  g072(.A1(new_n272), .A2(new_n273), .ZN(new_n274));
  INV_X1    g073(.A(G85gat), .ZN(new_n275));
  INV_X1    g074(.A(G92gat), .ZN(new_n276));
  NAND2_X1  g075(.A1(new_n275), .A2(new_n276), .ZN(new_n277));
  NAND3_X1  g076(.A1(KEYINPUT7), .A2(G85gat), .A3(G92gat), .ZN(new_n278));
  NAND4_X1  g077(.A1(new_n271), .A2(new_n274), .A3(new_n277), .A4(new_n278), .ZN(new_n279));
  XNOR2_X1  g078(.A(G99gat), .B(G106gat), .ZN(new_n280));
  INV_X1    g079(.A(new_n280), .ZN(new_n281));
  NAND2_X1  g080(.A1(new_n279), .A2(new_n281), .ZN(new_n282));
  AOI22_X1  g081(.A1(KEYINPUT8), .A2(new_n270), .B1(new_n275), .B2(new_n276), .ZN(new_n283));
  NAND4_X1  g082(.A1(new_n283), .A2(new_n280), .A3(new_n274), .A4(new_n278), .ZN(new_n284));
  NAND2_X1  g083(.A1(new_n282), .A2(new_n284), .ZN(new_n285));
  NAND3_X1  g084(.A1(new_n264), .A2(new_n269), .A3(new_n285), .ZN(new_n286));
  NAND2_X1  g085(.A1(new_n266), .A2(new_n268), .ZN(new_n287));
  AND2_X1   g086(.A1(new_n282), .A2(new_n284), .ZN(new_n288));
  NAND2_X1  g087(.A1(new_n287), .A2(new_n288), .ZN(new_n289));
  AND2_X1   g088(.A1(G232gat), .A2(G233gat), .ZN(new_n290));
  NAND2_X1  g089(.A1(new_n290), .A2(KEYINPUT41), .ZN(new_n291));
  AOI21_X1  g090(.A(KEYINPUT103), .B1(new_n289), .B2(new_n291), .ZN(new_n292));
  INV_X1    g091(.A(KEYINPUT103), .ZN(new_n293));
  INV_X1    g092(.A(new_n291), .ZN(new_n294));
  AOI211_X1 g093(.A(new_n293), .B(new_n294), .C1(new_n287), .C2(new_n288), .ZN(new_n295));
  OAI21_X1  g094(.A(new_n286), .B1(new_n292), .B2(new_n295), .ZN(new_n296));
  XOR2_X1   g095(.A(G190gat), .B(G218gat), .Z(new_n297));
  NAND2_X1  g096(.A1(new_n296), .A2(new_n297), .ZN(new_n298));
  NOR2_X1   g097(.A1(new_n290), .A2(KEYINPUT41), .ZN(new_n299));
  XNOR2_X1  g098(.A(G134gat), .B(G162gat), .ZN(new_n300));
  XNOR2_X1  g099(.A(new_n299), .B(new_n300), .ZN(new_n301));
  INV_X1    g100(.A(new_n297), .ZN(new_n302));
  OAI211_X1 g101(.A(new_n302), .B(new_n286), .C1(new_n292), .C2(new_n295), .ZN(new_n303));
  AND3_X1   g102(.A1(new_n298), .A2(new_n301), .A3(new_n303), .ZN(new_n304));
  AOI21_X1  g103(.A(new_n301), .B1(new_n298), .B2(new_n303), .ZN(new_n305));
  NOR2_X1   g104(.A1(new_n304), .A2(new_n305), .ZN(new_n306));
  NOR2_X1   g105(.A1(new_n244), .A2(new_n306), .ZN(new_n307));
  NAND2_X1  g106(.A1(new_n287), .A2(new_n233), .ZN(new_n308));
  NAND4_X1  g107(.A1(new_n266), .A2(new_n268), .A3(new_n228), .A4(new_n232), .ZN(new_n309));
  NAND3_X1  g108(.A1(new_n308), .A2(new_n309), .A3(KEYINPUT97), .ZN(new_n310));
  NAND2_X1  g109(.A1(G229gat), .A2(G233gat), .ZN(new_n311));
  XOR2_X1   g110(.A(new_n311), .B(KEYINPUT13), .Z(new_n312));
  INV_X1    g111(.A(KEYINPUT97), .ZN(new_n313));
  NAND3_X1  g112(.A1(new_n287), .A2(new_n313), .A3(new_n233), .ZN(new_n314));
  NAND3_X1  g113(.A1(new_n310), .A2(new_n312), .A3(new_n314), .ZN(new_n315));
  NAND2_X1  g114(.A1(new_n315), .A2(KEYINPUT98), .ZN(new_n316));
  INV_X1    g115(.A(KEYINPUT98), .ZN(new_n317));
  NAND4_X1  g116(.A1(new_n310), .A2(new_n317), .A3(new_n312), .A4(new_n314), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n316), .A2(new_n318), .ZN(new_n319));
  AOI22_X1  g118(.A1(new_n266), .A2(new_n268), .B1(new_n228), .B2(new_n232), .ZN(new_n320));
  AOI21_X1  g119(.A(new_n233), .B1(new_n287), .B2(new_n245), .ZN(new_n321));
  AOI21_X1  g120(.A(new_n320), .B1(new_n321), .B2(new_n269), .ZN(new_n322));
  INV_X1    g121(.A(KEYINPUT96), .ZN(new_n323));
  NAND4_X1  g122(.A1(new_n322), .A2(new_n323), .A3(KEYINPUT18), .A4(new_n311), .ZN(new_n324));
  NAND3_X1  g123(.A1(new_n234), .A2(new_n264), .A3(new_n269), .ZN(new_n325));
  NAND4_X1  g124(.A1(new_n325), .A2(KEYINPUT18), .A3(new_n311), .A4(new_n308), .ZN(new_n326));
  NAND2_X1  g125(.A1(new_n326), .A2(KEYINPUT96), .ZN(new_n327));
  NAND2_X1  g126(.A1(new_n324), .A2(new_n327), .ZN(new_n328));
  AOI21_X1  g127(.A(KEYINPUT18), .B1(new_n322), .B2(new_n311), .ZN(new_n329));
  INV_X1    g128(.A(new_n329), .ZN(new_n330));
  NAND3_X1  g129(.A1(new_n319), .A2(new_n328), .A3(new_n330), .ZN(new_n331));
  XNOR2_X1  g130(.A(G113gat), .B(G141gat), .ZN(new_n332));
  XNOR2_X1  g131(.A(G169gat), .B(G197gat), .ZN(new_n333));
  XNOR2_X1  g132(.A(new_n332), .B(new_n333), .ZN(new_n334));
  XNOR2_X1  g133(.A(KEYINPUT93), .B(KEYINPUT11), .ZN(new_n335));
  XNOR2_X1  g134(.A(new_n334), .B(new_n335), .ZN(new_n336));
  XOR2_X1   g135(.A(new_n336), .B(KEYINPUT12), .Z(new_n337));
  OAI21_X1  g136(.A(new_n337), .B1(new_n329), .B2(KEYINPUT99), .ZN(new_n338));
  INV_X1    g137(.A(new_n338), .ZN(new_n339));
  NAND2_X1  g138(.A1(new_n331), .A2(new_n339), .ZN(new_n340));
  AOI21_X1  g139(.A(new_n329), .B1(new_n316), .B2(new_n318), .ZN(new_n341));
  NAND3_X1  g140(.A1(new_n341), .A2(new_n338), .A3(new_n328), .ZN(new_n342));
  NAND2_X1  g141(.A1(new_n340), .A2(new_n342), .ZN(new_n343));
  NAND2_X1  g142(.A1(new_n285), .A2(new_n217), .ZN(new_n344));
  INV_X1    g143(.A(KEYINPUT10), .ZN(new_n345));
  NAND3_X1  g144(.A1(new_n209), .A2(new_n211), .A3(new_n212), .ZN(new_n346));
  OAI211_X1 g145(.A(new_n346), .B(new_n203), .C1(new_n207), .C2(new_n205), .ZN(new_n347));
  XNOR2_X1  g146(.A(G57gat), .B(G64gat), .ZN(new_n348));
  OAI211_X1 g147(.A(new_n206), .B(new_n215), .C1(new_n348), .C2(new_n204), .ZN(new_n349));
  NAND4_X1  g148(.A1(new_n347), .A2(new_n282), .A3(new_n349), .A4(new_n284), .ZN(new_n350));
  NAND3_X1  g149(.A1(new_n344), .A2(new_n345), .A3(new_n350), .ZN(new_n351));
  NAND4_X1  g150(.A1(new_n288), .A2(KEYINPUT10), .A3(new_n347), .A4(new_n349), .ZN(new_n352));
  NAND2_X1  g151(.A1(new_n351), .A2(new_n352), .ZN(new_n353));
  NAND2_X1  g152(.A1(G230gat), .A2(G233gat), .ZN(new_n354));
  NAND2_X1  g153(.A1(new_n353), .A2(new_n354), .ZN(new_n355));
  AND2_X1   g154(.A1(new_n344), .A2(new_n350), .ZN(new_n356));
  OAI21_X1  g155(.A(new_n355), .B1(new_n356), .B2(new_n354), .ZN(new_n357));
  XNOR2_X1  g156(.A(G120gat), .B(G148gat), .ZN(new_n358));
  XNOR2_X1  g157(.A(G176gat), .B(G204gat), .ZN(new_n359));
  XOR2_X1   g158(.A(new_n358), .B(new_n359), .Z(new_n360));
  INV_X1    g159(.A(new_n360), .ZN(new_n361));
  NOR2_X1   g160(.A1(new_n357), .A2(new_n361), .ZN(new_n362));
  INV_X1    g161(.A(new_n362), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n357), .A2(new_n361), .ZN(new_n364));
  NAND2_X1  g163(.A1(new_n363), .A2(new_n364), .ZN(new_n365));
  INV_X1    g164(.A(new_n365), .ZN(new_n366));
  NAND3_X1  g165(.A1(new_n307), .A2(new_n343), .A3(new_n366), .ZN(new_n367));
  XNOR2_X1  g166(.A(G155gat), .B(G162gat), .ZN(new_n368));
  INV_X1    g167(.A(KEYINPUT2), .ZN(new_n369));
  INV_X1    g168(.A(G148gat), .ZN(new_n370));
  NAND2_X1  g169(.A1(new_n370), .A2(G141gat), .ZN(new_n371));
  INV_X1    g170(.A(G141gat), .ZN(new_n372));
  NAND2_X1  g171(.A1(new_n372), .A2(G148gat), .ZN(new_n373));
  NAND2_X1  g172(.A1(new_n371), .A2(new_n373), .ZN(new_n374));
  AOI21_X1  g173(.A(new_n368), .B1(new_n369), .B2(new_n374), .ZN(new_n375));
  INV_X1    g174(.A(new_n375), .ZN(new_n376));
  XOR2_X1   g175(.A(KEYINPUT83), .B(KEYINPUT3), .Z(new_n377));
  NAND2_X1  g176(.A1(KEYINPUT82), .A2(G162gat), .ZN(new_n378));
  NAND2_X1  g177(.A1(new_n378), .A2(KEYINPUT2), .ZN(new_n379));
  NAND2_X1  g178(.A1(new_n368), .A2(new_n379), .ZN(new_n380));
  INV_X1    g179(.A(new_n380), .ZN(new_n381));
  INV_X1    g180(.A(KEYINPUT80), .ZN(new_n382));
  XNOR2_X1  g181(.A(new_n371), .B(new_n382), .ZN(new_n383));
  INV_X1    g182(.A(new_n383), .ZN(new_n384));
  XNOR2_X1  g183(.A(KEYINPUT78), .B(G141gat), .ZN(new_n385));
  INV_X1    g184(.A(KEYINPUT79), .ZN(new_n386));
  NAND3_X1  g185(.A1(new_n385), .A2(new_n386), .A3(G148gat), .ZN(new_n387));
  INV_X1    g186(.A(new_n387), .ZN(new_n388));
  AOI21_X1  g187(.A(new_n386), .B1(new_n385), .B2(G148gat), .ZN(new_n389));
  OAI21_X1  g188(.A(new_n384), .B1(new_n388), .B2(new_n389), .ZN(new_n390));
  INV_X1    g189(.A(KEYINPUT81), .ZN(new_n391));
  OAI21_X1  g190(.A(new_n381), .B1(new_n390), .B2(new_n391), .ZN(new_n392));
  XOR2_X1   g191(.A(KEYINPUT78), .B(G141gat), .Z(new_n393));
  OAI21_X1  g192(.A(KEYINPUT79), .B1(new_n393), .B2(new_n370), .ZN(new_n394));
  AOI21_X1  g193(.A(new_n383), .B1(new_n394), .B2(new_n387), .ZN(new_n395));
  NOR2_X1   g194(.A1(new_n395), .A2(KEYINPUT81), .ZN(new_n396));
  OAI211_X1 g195(.A(new_n376), .B(new_n377), .C1(new_n392), .C2(new_n396), .ZN(new_n397));
  XNOR2_X1  g196(.A(G113gat), .B(G120gat), .ZN(new_n398));
  NOR2_X1   g197(.A1(new_n398), .A2(KEYINPUT71), .ZN(new_n399));
  AND2_X1   g198(.A1(G127gat), .A2(G134gat), .ZN(new_n400));
  NOR2_X1   g199(.A1(G127gat), .A2(G134gat), .ZN(new_n401));
  NOR2_X1   g200(.A1(new_n400), .A2(new_n401), .ZN(new_n402));
  XNOR2_X1  g201(.A(KEYINPUT72), .B(KEYINPUT1), .ZN(new_n403));
  NOR3_X1   g202(.A1(new_n399), .A2(new_n402), .A3(new_n403), .ZN(new_n404));
  NAND2_X1  g203(.A1(new_n398), .A2(KEYINPUT71), .ZN(new_n405));
  OR2_X1    g204(.A1(new_n398), .A2(KEYINPUT1), .ZN(new_n406));
  XOR2_X1   g205(.A(KEYINPUT70), .B(G127gat), .Z(new_n407));
  AOI21_X1  g206(.A(new_n401), .B1(new_n407), .B2(G134gat), .ZN(new_n408));
  AOI22_X1  g207(.A1(new_n404), .A2(new_n405), .B1(new_n406), .B2(new_n408), .ZN(new_n409));
  INV_X1    g208(.A(new_n409), .ZN(new_n410));
  INV_X1    g209(.A(KEYINPUT3), .ZN(new_n411));
  AOI21_X1  g210(.A(new_n380), .B1(new_n395), .B2(KEYINPUT81), .ZN(new_n412));
  NAND2_X1  g211(.A1(new_n390), .A2(new_n391), .ZN(new_n413));
  AOI21_X1  g212(.A(new_n375), .B1(new_n412), .B2(new_n413), .ZN(new_n414));
  OAI211_X1 g213(.A(new_n397), .B(new_n410), .C1(new_n411), .C2(new_n414), .ZN(new_n415));
  NAND2_X1  g214(.A1(G225gat), .A2(G233gat), .ZN(new_n416));
  OAI211_X1 g215(.A(new_n409), .B(new_n376), .C1(new_n392), .C2(new_n396), .ZN(new_n417));
  INV_X1    g216(.A(KEYINPUT4), .ZN(new_n418));
  NAND2_X1  g217(.A1(new_n417), .A2(new_n418), .ZN(new_n419));
  NAND3_X1  g218(.A1(new_n414), .A2(KEYINPUT4), .A3(new_n409), .ZN(new_n420));
  NAND4_X1  g219(.A1(new_n415), .A2(new_n416), .A3(new_n419), .A4(new_n420), .ZN(new_n421));
  XOR2_X1   g220(.A(KEYINPUT86), .B(KEYINPUT5), .Z(new_n422));
  INV_X1    g221(.A(new_n422), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n423), .A2(KEYINPUT84), .ZN(new_n424));
  NAND2_X1  g223(.A1(new_n421), .A2(new_n424), .ZN(new_n425));
  AND2_X1   g224(.A1(new_n419), .A2(new_n420), .ZN(new_n426));
  INV_X1    g225(.A(new_n424), .ZN(new_n427));
  NAND4_X1  g226(.A1(new_n426), .A2(new_n416), .A3(new_n415), .A4(new_n427), .ZN(new_n428));
  OAI21_X1  g227(.A(new_n376), .B1(new_n392), .B2(new_n396), .ZN(new_n429));
  NAND2_X1  g228(.A1(new_n429), .A2(new_n410), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n430), .A2(new_n417), .ZN(new_n431));
  INV_X1    g230(.A(KEYINPUT85), .ZN(new_n432));
  INV_X1    g231(.A(new_n416), .ZN(new_n433));
  NAND3_X1  g232(.A1(new_n431), .A2(new_n432), .A3(new_n433), .ZN(new_n434));
  NAND2_X1  g233(.A1(new_n434), .A2(new_n423), .ZN(new_n435));
  AOI21_X1  g234(.A(new_n416), .B1(new_n430), .B2(new_n417), .ZN(new_n436));
  NOR2_X1   g235(.A1(new_n436), .A2(new_n432), .ZN(new_n437));
  OAI211_X1 g236(.A(new_n425), .B(new_n428), .C1(new_n435), .C2(new_n437), .ZN(new_n438));
  XOR2_X1   g237(.A(G1gat), .B(G29gat), .Z(new_n439));
  XNOR2_X1  g238(.A(G57gat), .B(G85gat), .ZN(new_n440));
  XNOR2_X1  g239(.A(new_n439), .B(new_n440), .ZN(new_n441));
  XNOR2_X1  g240(.A(KEYINPUT87), .B(KEYINPUT0), .ZN(new_n442));
  XNOR2_X1  g241(.A(new_n441), .B(new_n442), .ZN(new_n443));
  INV_X1    g242(.A(new_n443), .ZN(new_n444));
  NAND2_X1  g243(.A1(new_n438), .A2(new_n444), .ZN(new_n445));
  INV_X1    g244(.A(KEYINPUT6), .ZN(new_n446));
  AOI21_X1  g245(.A(new_n422), .B1(new_n436), .B2(new_n432), .ZN(new_n447));
  OAI21_X1  g246(.A(new_n447), .B1(new_n432), .B2(new_n436), .ZN(new_n448));
  NAND4_X1  g247(.A1(new_n448), .A2(new_n443), .A3(new_n428), .A4(new_n425), .ZN(new_n449));
  NAND3_X1  g248(.A1(new_n445), .A2(new_n446), .A3(new_n449), .ZN(new_n450));
  OR3_X1    g249(.A1(new_n438), .A2(new_n446), .A3(new_n444), .ZN(new_n451));
  NAND2_X1  g250(.A1(G226gat), .A2(G233gat), .ZN(new_n452));
  INV_X1    g251(.A(new_n452), .ZN(new_n453));
  NAND2_X1  g252(.A1(G169gat), .A2(G176gat), .ZN(new_n454));
  XNOR2_X1  g253(.A(new_n454), .B(KEYINPUT66), .ZN(new_n455));
  NOR2_X1   g254(.A1(G169gat), .A2(G176gat), .ZN(new_n456));
  NAND2_X1  g255(.A1(new_n456), .A2(KEYINPUT23), .ZN(new_n457));
  NAND2_X1  g256(.A1(new_n455), .A2(new_n457), .ZN(new_n458));
  XNOR2_X1  g257(.A(new_n458), .B(KEYINPUT67), .ZN(new_n459));
  XNOR2_X1  g258(.A(KEYINPUT65), .B(KEYINPUT23), .ZN(new_n460));
  OAI21_X1  g259(.A(new_n460), .B1(G169gat), .B2(G176gat), .ZN(new_n461));
  AND2_X1   g260(.A1(new_n461), .A2(KEYINPUT25), .ZN(new_n462));
  NAND2_X1  g261(.A1(G183gat), .A2(G190gat), .ZN(new_n463));
  NOR2_X1   g262(.A1(new_n463), .A2(KEYINPUT24), .ZN(new_n464));
  XOR2_X1   g263(.A(G183gat), .B(G190gat), .Z(new_n465));
  AOI21_X1  g264(.A(new_n464), .B1(new_n465), .B2(KEYINPUT24), .ZN(new_n466));
  AND2_X1   g265(.A1(new_n462), .A2(new_n466), .ZN(new_n467));
  NAND3_X1  g266(.A1(new_n456), .A2(KEYINPUT64), .A3(KEYINPUT23), .ZN(new_n468));
  AND2_X1   g267(.A1(new_n455), .A2(new_n468), .ZN(new_n469));
  INV_X1    g268(.A(KEYINPUT64), .ZN(new_n470));
  NAND2_X1  g269(.A1(new_n457), .A2(new_n470), .ZN(new_n471));
  NAND4_X1  g270(.A1(new_n469), .A2(new_n466), .A3(new_n461), .A4(new_n471), .ZN(new_n472));
  INV_X1    g271(.A(KEYINPUT25), .ZN(new_n473));
  AOI22_X1  g272(.A1(new_n459), .A2(new_n467), .B1(new_n472), .B2(new_n473), .ZN(new_n474));
  INV_X1    g273(.A(KEYINPUT77), .ZN(new_n475));
  XNOR2_X1  g274(.A(new_n456), .B(KEYINPUT26), .ZN(new_n476));
  NAND2_X1  g275(.A1(new_n476), .A2(new_n455), .ZN(new_n477));
  NAND2_X1  g276(.A1(new_n477), .A2(new_n463), .ZN(new_n478));
  XNOR2_X1  g277(.A(KEYINPUT27), .B(G183gat), .ZN(new_n479));
  XNOR2_X1  g278(.A(new_n479), .B(KEYINPUT69), .ZN(new_n480));
  INV_X1    g279(.A(G190gat), .ZN(new_n481));
  NAND3_X1  g280(.A1(new_n480), .A2(KEYINPUT28), .A3(new_n481), .ZN(new_n482));
  AOI21_X1  g281(.A(KEYINPUT28), .B1(new_n479), .B2(new_n481), .ZN(new_n483));
  INV_X1    g282(.A(new_n483), .ZN(new_n484));
  AOI21_X1  g283(.A(new_n478), .B1(new_n482), .B2(new_n484), .ZN(new_n485));
  NOR3_X1   g284(.A1(new_n474), .A2(new_n475), .A3(new_n485), .ZN(new_n486));
  NOR2_X1   g285(.A1(new_n458), .A2(KEYINPUT67), .ZN(new_n487));
  INV_X1    g286(.A(KEYINPUT67), .ZN(new_n488));
  AOI21_X1  g287(.A(new_n488), .B1(new_n455), .B2(new_n457), .ZN(new_n489));
  OAI211_X1 g288(.A(new_n466), .B(new_n462), .C1(new_n487), .C2(new_n489), .ZN(new_n490));
  NAND4_X1  g289(.A1(new_n461), .A2(new_n468), .A3(new_n455), .A4(new_n471), .ZN(new_n491));
  INV_X1    g290(.A(new_n466), .ZN(new_n492));
  OAI21_X1  g291(.A(new_n473), .B1(new_n491), .B2(new_n492), .ZN(new_n493));
  NAND2_X1  g292(.A1(new_n490), .A2(new_n493), .ZN(new_n494));
  NAND2_X1  g293(.A1(new_n482), .A2(new_n484), .ZN(new_n495));
  INV_X1    g294(.A(new_n478), .ZN(new_n496));
  NAND2_X1  g295(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  AOI21_X1  g296(.A(KEYINPUT77), .B1(new_n494), .B2(new_n497), .ZN(new_n498));
  OAI21_X1  g297(.A(new_n453), .B1(new_n486), .B2(new_n498), .ZN(new_n499));
  INV_X1    g298(.A(KEYINPUT68), .ZN(new_n500));
  AND3_X1   g299(.A1(new_n490), .A2(new_n500), .A3(new_n493), .ZN(new_n501));
  AOI21_X1  g300(.A(new_n500), .B1(new_n490), .B2(new_n493), .ZN(new_n502));
  OAI21_X1  g301(.A(new_n497), .B1(new_n501), .B2(new_n502), .ZN(new_n503));
  NOR2_X1   g302(.A1(new_n453), .A2(KEYINPUT29), .ZN(new_n504));
  NAND2_X1  g303(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  AOI21_X1  g304(.A(KEYINPUT22), .B1(G211gat), .B2(G218gat), .ZN(new_n506));
  XNOR2_X1  g305(.A(KEYINPUT75), .B(G197gat), .ZN(new_n507));
  OR2_X1    g306(.A1(new_n507), .A2(G204gat), .ZN(new_n508));
  NAND2_X1  g307(.A1(new_n507), .A2(G204gat), .ZN(new_n509));
  AOI21_X1  g308(.A(new_n506), .B1(new_n508), .B2(new_n509), .ZN(new_n510));
  INV_X1    g309(.A(KEYINPUT76), .ZN(new_n511));
  XOR2_X1   g310(.A(G211gat), .B(G218gat), .Z(new_n512));
  OR3_X1    g311(.A1(new_n510), .A2(new_n511), .A3(new_n512), .ZN(new_n513));
  OAI21_X1  g312(.A(new_n512), .B1(new_n510), .B2(new_n511), .ZN(new_n514));
  NAND2_X1  g313(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  AND3_X1   g314(.A1(new_n499), .A2(new_n505), .A3(new_n515), .ZN(new_n516));
  OAI21_X1  g315(.A(new_n475), .B1(new_n474), .B2(new_n485), .ZN(new_n517));
  NAND3_X1  g316(.A1(new_n494), .A2(new_n497), .A3(KEYINPUT77), .ZN(new_n518));
  NAND3_X1  g317(.A1(new_n517), .A2(new_n518), .A3(new_n504), .ZN(new_n519));
  OAI211_X1 g318(.A(new_n497), .B(new_n453), .C1(new_n501), .C2(new_n502), .ZN(new_n520));
  AOI21_X1  g319(.A(new_n515), .B1(new_n519), .B2(new_n520), .ZN(new_n521));
  NOR2_X1   g320(.A1(new_n516), .A2(new_n521), .ZN(new_n522));
  INV_X1    g321(.A(KEYINPUT30), .ZN(new_n523));
  XNOR2_X1  g322(.A(G8gat), .B(G36gat), .ZN(new_n524));
  XNOR2_X1  g323(.A(G64gat), .B(G92gat), .ZN(new_n525));
  XOR2_X1   g324(.A(new_n524), .B(new_n525), .Z(new_n526));
  NAND3_X1  g325(.A1(new_n522), .A2(new_n523), .A3(new_n526), .ZN(new_n527));
  INV_X1    g326(.A(new_n526), .ZN(new_n528));
  OAI21_X1  g327(.A(new_n528), .B1(new_n516), .B2(new_n521), .ZN(new_n529));
  NAND2_X1  g328(.A1(new_n519), .A2(new_n520), .ZN(new_n530));
  INV_X1    g329(.A(new_n515), .ZN(new_n531));
  NAND2_X1  g330(.A1(new_n530), .A2(new_n531), .ZN(new_n532));
  NAND3_X1  g331(.A1(new_n499), .A2(new_n505), .A3(new_n515), .ZN(new_n533));
  NAND3_X1  g332(.A1(new_n532), .A2(new_n533), .A3(new_n526), .ZN(new_n534));
  NAND3_X1  g333(.A1(new_n529), .A2(KEYINPUT30), .A3(new_n534), .ZN(new_n535));
  AOI22_X1  g334(.A1(new_n450), .A2(new_n451), .B1(new_n527), .B2(new_n535), .ZN(new_n536));
  INV_X1    g335(.A(KEYINPUT35), .ZN(new_n537));
  XNOR2_X1  g336(.A(G78gat), .B(G106gat), .ZN(new_n538));
  XNOR2_X1  g337(.A(new_n538), .B(G22gat), .ZN(new_n539));
  INV_X1    g338(.A(new_n539), .ZN(new_n540));
  AND2_X1   g339(.A1(G228gat), .A2(G233gat), .ZN(new_n541));
  INV_X1    g340(.A(KEYINPUT29), .ZN(new_n542));
  NAND2_X1  g341(.A1(new_n531), .A2(new_n542), .ZN(new_n543));
  AOI21_X1  g342(.A(new_n414), .B1(new_n543), .B2(new_n411), .ZN(new_n544));
  AOI21_X1  g343(.A(KEYINPUT29), .B1(new_n414), .B2(new_n377), .ZN(new_n545));
  NOR2_X1   g344(.A1(new_n545), .A2(new_n531), .ZN(new_n546));
  OAI21_X1  g345(.A(new_n541), .B1(new_n544), .B2(new_n546), .ZN(new_n547));
  AND2_X1   g346(.A1(new_n510), .A2(KEYINPUT88), .ZN(new_n548));
  NOR2_X1   g347(.A1(new_n510), .A2(KEYINPUT88), .ZN(new_n549));
  INV_X1    g348(.A(new_n512), .ZN(new_n550));
  NOR3_X1   g349(.A1(new_n548), .A2(new_n549), .A3(new_n550), .ZN(new_n551));
  NAND2_X1  g350(.A1(new_n549), .A2(new_n550), .ZN(new_n552));
  NAND2_X1  g351(.A1(new_n552), .A2(new_n542), .ZN(new_n553));
  OAI21_X1  g352(.A(new_n377), .B1(new_n551), .B2(new_n553), .ZN(new_n554));
  AOI21_X1  g353(.A(new_n541), .B1(new_n554), .B2(new_n429), .ZN(new_n555));
  OAI21_X1  g354(.A(KEYINPUT89), .B1(new_n545), .B2(new_n531), .ZN(new_n556));
  NAND2_X1  g355(.A1(new_n397), .A2(new_n542), .ZN(new_n557));
  INV_X1    g356(.A(KEYINPUT89), .ZN(new_n558));
  NAND3_X1  g357(.A1(new_n557), .A2(new_n558), .A3(new_n515), .ZN(new_n559));
  NAND3_X1  g358(.A1(new_n555), .A2(new_n556), .A3(new_n559), .ZN(new_n560));
  XNOR2_X1  g359(.A(KEYINPUT31), .B(G50gat), .ZN(new_n561));
  INV_X1    g360(.A(new_n561), .ZN(new_n562));
  NAND3_X1  g361(.A1(new_n547), .A2(new_n560), .A3(new_n562), .ZN(new_n563));
  INV_X1    g362(.A(new_n563), .ZN(new_n564));
  AOI21_X1  g363(.A(new_n562), .B1(new_n547), .B2(new_n560), .ZN(new_n565));
  OAI21_X1  g364(.A(new_n540), .B1(new_n564), .B2(new_n565), .ZN(new_n566));
  INV_X1    g365(.A(new_n565), .ZN(new_n567));
  NAND3_X1  g366(.A1(new_n567), .A2(new_n539), .A3(new_n563), .ZN(new_n568));
  AND2_X1   g367(.A1(new_n566), .A2(new_n568), .ZN(new_n569));
  NAND3_X1  g368(.A1(new_n536), .A2(new_n537), .A3(new_n569), .ZN(new_n570));
  INV_X1    g369(.A(new_n570), .ZN(new_n571));
  INV_X1    g370(.A(KEYINPUT74), .ZN(new_n572));
  NAND2_X1  g371(.A1(new_n503), .A2(new_n409), .ZN(new_n573));
  INV_X1    g372(.A(G227gat), .ZN(new_n574));
  INV_X1    g373(.A(G233gat), .ZN(new_n575));
  NOR2_X1   g374(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  OAI211_X1 g375(.A(new_n410), .B(new_n497), .C1(new_n501), .C2(new_n502), .ZN(new_n577));
  NAND3_X1  g376(.A1(new_n573), .A2(new_n576), .A3(new_n577), .ZN(new_n578));
  XNOR2_X1  g377(.A(G15gat), .B(G43gat), .ZN(new_n579));
  XNOR2_X1  g378(.A(G71gat), .B(G99gat), .ZN(new_n580));
  XNOR2_X1  g379(.A(new_n579), .B(new_n580), .ZN(new_n581));
  INV_X1    g380(.A(KEYINPUT33), .ZN(new_n582));
  OR2_X1    g381(.A1(new_n581), .A2(new_n582), .ZN(new_n583));
  NAND3_X1  g382(.A1(new_n578), .A2(KEYINPUT32), .A3(new_n583), .ZN(new_n584));
  NAND2_X1  g383(.A1(new_n584), .A2(KEYINPUT73), .ZN(new_n585));
  INV_X1    g384(.A(KEYINPUT73), .ZN(new_n586));
  NAND4_X1  g385(.A1(new_n578), .A2(new_n586), .A3(KEYINPUT32), .A4(new_n583), .ZN(new_n587));
  NAND2_X1  g386(.A1(new_n585), .A2(new_n587), .ZN(new_n588));
  AOI21_X1  g387(.A(new_n581), .B1(new_n578), .B2(KEYINPUT32), .ZN(new_n589));
  NAND2_X1  g388(.A1(new_n578), .A2(new_n582), .ZN(new_n590));
  NAND2_X1  g389(.A1(new_n589), .A2(new_n590), .ZN(new_n591));
  NAND2_X1  g390(.A1(new_n588), .A2(new_n591), .ZN(new_n592));
  AOI21_X1  g391(.A(new_n576), .B1(new_n573), .B2(new_n577), .ZN(new_n593));
  INV_X1    g392(.A(KEYINPUT34), .ZN(new_n594));
  NOR2_X1   g393(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  AOI211_X1 g394(.A(KEYINPUT34), .B(new_n576), .C1(new_n573), .C2(new_n577), .ZN(new_n596));
  NOR2_X1   g395(.A1(new_n595), .A2(new_n596), .ZN(new_n597));
  INV_X1    g396(.A(new_n597), .ZN(new_n598));
  NAND2_X1  g397(.A1(new_n592), .A2(new_n598), .ZN(new_n599));
  AOI22_X1  g398(.A1(new_n585), .A2(new_n587), .B1(new_n590), .B2(new_n589), .ZN(new_n600));
  NAND2_X1  g399(.A1(new_n600), .A2(new_n597), .ZN(new_n601));
  AOI21_X1  g400(.A(new_n572), .B1(new_n599), .B2(new_n601), .ZN(new_n602));
  AOI21_X1  g401(.A(KEYINPUT74), .B1(new_n600), .B2(new_n597), .ZN(new_n603));
  NOR3_X1   g402(.A1(new_n602), .A2(KEYINPUT92), .A3(new_n603), .ZN(new_n604));
  INV_X1    g403(.A(KEYINPUT92), .ZN(new_n605));
  AND3_X1   g404(.A1(new_n588), .A2(new_n597), .A3(new_n591), .ZN(new_n606));
  AOI21_X1  g405(.A(new_n597), .B1(new_n588), .B2(new_n591), .ZN(new_n607));
  OAI21_X1  g406(.A(KEYINPUT74), .B1(new_n606), .B2(new_n607), .ZN(new_n608));
  INV_X1    g407(.A(new_n603), .ZN(new_n609));
  AOI21_X1  g408(.A(new_n605), .B1(new_n608), .B2(new_n609), .ZN(new_n610));
  OAI21_X1  g409(.A(new_n571), .B1(new_n604), .B2(new_n610), .ZN(new_n611));
  NAND2_X1  g410(.A1(new_n599), .A2(new_n601), .ZN(new_n612));
  NAND2_X1  g411(.A1(new_n566), .A2(new_n568), .ZN(new_n613));
  NOR2_X1   g412(.A1(new_n612), .A2(new_n613), .ZN(new_n614));
  AOI21_X1  g413(.A(new_n537), .B1(new_n614), .B2(new_n536), .ZN(new_n615));
  INV_X1    g414(.A(new_n615), .ZN(new_n616));
  NAND2_X1  g415(.A1(new_n611), .A2(new_n616), .ZN(new_n617));
  AND2_X1   g416(.A1(new_n450), .A2(new_n451), .ZN(new_n618));
  INV_X1    g417(.A(KEYINPUT37), .ZN(new_n619));
  OAI211_X1 g418(.A(KEYINPUT91), .B(new_n528), .C1(new_n522), .C2(new_n619), .ZN(new_n620));
  INV_X1    g419(.A(KEYINPUT91), .ZN(new_n621));
  AOI21_X1  g420(.A(new_n619), .B1(new_n532), .B2(new_n533), .ZN(new_n622));
  OAI21_X1  g421(.A(new_n621), .B1(new_n622), .B2(new_n526), .ZN(new_n623));
  NAND2_X1  g422(.A1(new_n522), .A2(new_n619), .ZN(new_n624));
  NAND3_X1  g423(.A1(new_n620), .A2(new_n623), .A3(new_n624), .ZN(new_n625));
  NAND2_X1  g424(.A1(new_n625), .A2(KEYINPUT38), .ZN(new_n626));
  AOI211_X1 g425(.A(KEYINPUT38), .B(new_n526), .C1(new_n522), .C2(new_n619), .ZN(new_n627));
  NAND2_X1  g426(.A1(new_n530), .A2(new_n515), .ZN(new_n628));
  NAND3_X1  g427(.A1(new_n499), .A2(new_n505), .A3(new_n531), .ZN(new_n629));
  NAND3_X1  g428(.A1(new_n628), .A2(KEYINPUT37), .A3(new_n629), .ZN(new_n630));
  AOI22_X1  g429(.A1(new_n627), .A2(new_n630), .B1(new_n522), .B2(new_n526), .ZN(new_n631));
  NAND3_X1  g430(.A1(new_n618), .A2(new_n626), .A3(new_n631), .ZN(new_n632));
  NOR2_X1   g431(.A1(KEYINPUT90), .A2(KEYINPUT40), .ZN(new_n633));
  AOI21_X1  g432(.A(new_n416), .B1(new_n426), .B2(new_n415), .ZN(new_n634));
  INV_X1    g433(.A(KEYINPUT39), .ZN(new_n635));
  NAND2_X1  g434(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  NAND2_X1  g435(.A1(new_n636), .A2(new_n444), .ZN(new_n637));
  OAI21_X1  g436(.A(KEYINPUT39), .B1(new_n431), .B2(new_n433), .ZN(new_n638));
  NOR2_X1   g437(.A1(new_n634), .A2(new_n638), .ZN(new_n639));
  OAI21_X1  g438(.A(new_n633), .B1(new_n637), .B2(new_n639), .ZN(new_n640));
  INV_X1    g439(.A(new_n639), .ZN(new_n641));
  INV_X1    g440(.A(new_n633), .ZN(new_n642));
  NAND4_X1  g441(.A1(new_n641), .A2(new_n444), .A3(new_n642), .A4(new_n636), .ZN(new_n643));
  AND2_X1   g442(.A1(new_n640), .A2(new_n643), .ZN(new_n644));
  AND3_X1   g443(.A1(new_n535), .A2(new_n449), .A3(new_n527), .ZN(new_n645));
  AOI21_X1  g444(.A(new_n613), .B1(new_n644), .B2(new_n645), .ZN(new_n646));
  NAND2_X1  g445(.A1(new_n632), .A2(new_n646), .ZN(new_n647));
  NAND2_X1  g446(.A1(new_n450), .A2(new_n451), .ZN(new_n648));
  NAND2_X1  g447(.A1(new_n535), .A2(new_n527), .ZN(new_n649));
  NAND2_X1  g448(.A1(new_n648), .A2(new_n649), .ZN(new_n650));
  NAND2_X1  g449(.A1(new_n650), .A2(new_n613), .ZN(new_n651));
  AOI21_X1  g450(.A(KEYINPUT36), .B1(new_n608), .B2(new_n609), .ZN(new_n652));
  NAND3_X1  g451(.A1(new_n599), .A2(KEYINPUT36), .A3(new_n601), .ZN(new_n653));
  INV_X1    g452(.A(new_n653), .ZN(new_n654));
  OAI211_X1 g453(.A(new_n647), .B(new_n651), .C1(new_n652), .C2(new_n654), .ZN(new_n655));
  AOI21_X1  g454(.A(new_n367), .B1(new_n617), .B2(new_n655), .ZN(new_n656));
  NAND2_X1  g455(.A1(new_n656), .A2(new_n618), .ZN(new_n657));
  XNOR2_X1  g456(.A(new_n657), .B(G1gat), .ZN(G1324gat));
  INV_X1    g457(.A(new_n649), .ZN(new_n659));
  AND2_X1   g458(.A1(new_n656), .A2(new_n659), .ZN(new_n660));
  OR2_X1    g459(.A1(new_n660), .A2(new_n230), .ZN(new_n661));
  INV_X1    g460(.A(KEYINPUT42), .ZN(new_n662));
  XOR2_X1   g461(.A(KEYINPUT16), .B(G8gat), .Z(new_n663));
  AOI21_X1  g462(.A(new_n662), .B1(new_n660), .B2(new_n663), .ZN(new_n664));
  INV_X1    g463(.A(KEYINPUT104), .ZN(new_n665));
  NOR2_X1   g464(.A1(new_n663), .A2(new_n665), .ZN(new_n666));
  NAND2_X1  g465(.A1(new_n662), .A2(KEYINPUT104), .ZN(new_n667));
  AOI21_X1  g466(.A(new_n666), .B1(new_n663), .B2(new_n667), .ZN(new_n668));
  AOI22_X1  g467(.A1(new_n661), .A2(new_n664), .B1(new_n660), .B2(new_n668), .ZN(G1325gat));
  INV_X1    g468(.A(KEYINPUT36), .ZN(new_n670));
  OAI21_X1  g469(.A(new_n670), .B1(new_n602), .B2(new_n603), .ZN(new_n671));
  NAND2_X1  g470(.A1(new_n671), .A2(new_n653), .ZN(new_n672));
  INV_X1    g471(.A(new_n672), .ZN(new_n673));
  NAND2_X1  g472(.A1(new_n656), .A2(new_n673), .ZN(new_n674));
  OAI21_X1  g473(.A(KEYINPUT92), .B1(new_n602), .B2(new_n603), .ZN(new_n675));
  NAND3_X1  g474(.A1(new_n608), .A2(new_n605), .A3(new_n609), .ZN(new_n676));
  NAND2_X1  g475(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  INV_X1    g476(.A(new_n677), .ZN(new_n678));
  NOR2_X1   g477(.A1(new_n678), .A2(G15gat), .ZN(new_n679));
  AOI22_X1  g478(.A1(new_n674), .A2(G15gat), .B1(new_n656), .B2(new_n679), .ZN(new_n680));
  XOR2_X1   g479(.A(new_n680), .B(KEYINPUT105), .Z(G1326gat));
  NAND2_X1  g480(.A1(new_n656), .A2(new_n613), .ZN(new_n682));
  XNOR2_X1  g481(.A(new_n682), .B(KEYINPUT106), .ZN(new_n683));
  XNOR2_X1  g482(.A(KEYINPUT43), .B(G22gat), .ZN(new_n684));
  INV_X1    g483(.A(new_n684), .ZN(new_n685));
  XNOR2_X1  g484(.A(new_n683), .B(new_n685), .ZN(G1327gat));
  AOI21_X1  g485(.A(new_n570), .B1(new_n675), .B2(new_n676), .ZN(new_n687));
  OAI21_X1  g486(.A(new_n655), .B1(new_n687), .B2(new_n615), .ZN(new_n688));
  INV_X1    g487(.A(new_n343), .ZN(new_n689));
  NOR3_X1   g488(.A1(new_n689), .A2(new_n243), .A3(new_n365), .ZN(new_n690));
  NAND3_X1  g489(.A1(new_n688), .A2(new_n306), .A3(new_n690), .ZN(new_n691));
  INV_X1    g490(.A(new_n691), .ZN(new_n692));
  NAND3_X1  g491(.A1(new_n692), .A2(new_n252), .A3(new_n618), .ZN(new_n693));
  XNOR2_X1  g492(.A(new_n693), .B(KEYINPUT45), .ZN(new_n694));
  NAND2_X1  g493(.A1(new_n688), .A2(new_n306), .ZN(new_n695));
  NAND2_X1  g494(.A1(new_n695), .A2(KEYINPUT44), .ZN(new_n696));
  INV_X1    g495(.A(new_n306), .ZN(new_n697));
  AOI21_X1  g496(.A(KEYINPUT107), .B1(new_n650), .B2(new_n613), .ZN(new_n698));
  INV_X1    g497(.A(KEYINPUT107), .ZN(new_n699));
  NOR3_X1   g498(.A1(new_n536), .A2(new_n569), .A3(new_n699), .ZN(new_n700));
  NOR2_X1   g499(.A1(new_n698), .A2(new_n700), .ZN(new_n701));
  NAND3_X1  g500(.A1(new_n701), .A2(new_n672), .A3(new_n647), .ZN(new_n702));
  AOI21_X1  g501(.A(new_n697), .B1(new_n617), .B2(new_n702), .ZN(new_n703));
  XOR2_X1   g502(.A(KEYINPUT108), .B(KEYINPUT44), .Z(new_n704));
  NAND2_X1  g503(.A1(new_n703), .A2(new_n704), .ZN(new_n705));
  NAND2_X1  g504(.A1(new_n696), .A2(new_n705), .ZN(new_n706));
  NAND2_X1  g505(.A1(new_n706), .A2(new_n690), .ZN(new_n707));
  OAI21_X1  g506(.A(G29gat), .B1(new_n707), .B2(new_n648), .ZN(new_n708));
  NAND2_X1  g507(.A1(new_n694), .A2(new_n708), .ZN(G1328gat));
  NAND3_X1  g508(.A1(new_n706), .A2(new_n659), .A3(new_n690), .ZN(new_n710));
  INV_X1    g509(.A(KEYINPUT109), .ZN(new_n711));
  NAND2_X1  g510(.A1(new_n710), .A2(new_n711), .ZN(new_n712));
  NAND4_X1  g511(.A1(new_n706), .A2(KEYINPUT109), .A3(new_n659), .A4(new_n690), .ZN(new_n713));
  NAND3_X1  g512(.A1(new_n712), .A2(G36gat), .A3(new_n713), .ZN(new_n714));
  NOR3_X1   g513(.A1(new_n691), .A2(G36gat), .A3(new_n649), .ZN(new_n715));
  XNOR2_X1  g514(.A(new_n715), .B(KEYINPUT46), .ZN(new_n716));
  NAND2_X1  g515(.A1(new_n714), .A2(new_n716), .ZN(G1329gat));
  INV_X1    g516(.A(G43gat), .ZN(new_n718));
  OAI21_X1  g517(.A(new_n718), .B1(new_n691), .B2(new_n678), .ZN(new_n719));
  NAND2_X1  g518(.A1(new_n673), .A2(G43gat), .ZN(new_n720));
  OAI21_X1  g519(.A(new_n719), .B1(new_n707), .B2(new_n720), .ZN(new_n721));
  NAND2_X1  g520(.A1(new_n721), .A2(KEYINPUT47), .ZN(new_n722));
  INV_X1    g521(.A(KEYINPUT47), .ZN(new_n723));
  OAI211_X1 g522(.A(new_n719), .B(new_n723), .C1(new_n707), .C2(new_n720), .ZN(new_n724));
  NAND2_X1  g523(.A1(new_n722), .A2(new_n724), .ZN(G1330gat));
  INV_X1    g524(.A(new_n704), .ZN(new_n726));
  AOI211_X1 g525(.A(new_n697), .B(new_n726), .C1(new_n617), .C2(new_n702), .ZN(new_n727));
  INV_X1    g526(.A(KEYINPUT44), .ZN(new_n728));
  AOI21_X1  g527(.A(new_n728), .B1(new_n688), .B2(new_n306), .ZN(new_n729));
  OAI211_X1 g528(.A(new_n613), .B(new_n690), .C1(new_n727), .C2(new_n729), .ZN(new_n730));
  NAND2_X1  g529(.A1(new_n730), .A2(G50gat), .ZN(new_n731));
  NOR2_X1   g530(.A1(new_n569), .A2(G50gat), .ZN(new_n732));
  XNOR2_X1  g531(.A(new_n732), .B(KEYINPUT110), .ZN(new_n733));
  NAND2_X1  g532(.A1(new_n692), .A2(new_n733), .ZN(new_n734));
  NAND2_X1  g533(.A1(new_n731), .A2(new_n734), .ZN(new_n735));
  INV_X1    g534(.A(KEYINPUT48), .ZN(new_n736));
  NAND2_X1  g535(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  NAND3_X1  g536(.A1(new_n731), .A2(KEYINPUT48), .A3(new_n734), .ZN(new_n738));
  NAND2_X1  g537(.A1(new_n737), .A2(new_n738), .ZN(G1331gat));
  NAND2_X1  g538(.A1(new_n617), .A2(new_n702), .ZN(new_n740));
  INV_X1    g539(.A(new_n740), .ZN(new_n741));
  NAND3_X1  g540(.A1(new_n307), .A2(new_n689), .A3(new_n365), .ZN(new_n742));
  NOR2_X1   g541(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  INV_X1    g542(.A(KEYINPUT111), .ZN(new_n744));
  NAND2_X1  g543(.A1(new_n648), .A2(new_n744), .ZN(new_n745));
  NAND3_X1  g544(.A1(new_n450), .A2(new_n451), .A3(KEYINPUT111), .ZN(new_n746));
  NAND2_X1  g545(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  NAND2_X1  g546(.A1(new_n743), .A2(new_n747), .ZN(new_n748));
  XNOR2_X1  g547(.A(new_n748), .B(G57gat), .ZN(G1332gat));
  NOR3_X1   g548(.A1(new_n741), .A2(new_n649), .A3(new_n742), .ZN(new_n750));
  NOR2_X1   g549(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n751));
  AND2_X1   g550(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n752));
  OAI21_X1  g551(.A(new_n750), .B1(new_n751), .B2(new_n752), .ZN(new_n753));
  OAI21_X1  g552(.A(new_n753), .B1(new_n750), .B2(new_n751), .ZN(G1333gat));
  INV_X1    g553(.A(KEYINPUT112), .ZN(new_n755));
  XNOR2_X1  g554(.A(new_n677), .B(new_n755), .ZN(new_n756));
  NAND2_X1  g555(.A1(new_n743), .A2(new_n756), .ZN(new_n757));
  INV_X1    g556(.A(G71gat), .ZN(new_n758));
  NAND2_X1  g557(.A1(new_n757), .A2(new_n758), .ZN(new_n759));
  NAND3_X1  g558(.A1(new_n743), .A2(G71gat), .A3(new_n673), .ZN(new_n760));
  NAND2_X1  g559(.A1(new_n759), .A2(new_n760), .ZN(new_n761));
  NAND2_X1  g560(.A1(new_n761), .A2(KEYINPUT50), .ZN(new_n762));
  INV_X1    g561(.A(KEYINPUT50), .ZN(new_n763));
  NAND3_X1  g562(.A1(new_n759), .A2(new_n763), .A3(new_n760), .ZN(new_n764));
  NAND2_X1  g563(.A1(new_n762), .A2(new_n764), .ZN(G1334gat));
  NAND2_X1  g564(.A1(new_n743), .A2(new_n613), .ZN(new_n766));
  XNOR2_X1  g565(.A(new_n766), .B(G78gat), .ZN(G1335gat));
  NOR3_X1   g566(.A1(new_n648), .A2(G85gat), .A3(new_n366), .ZN(new_n768));
  NOR2_X1   g567(.A1(new_n243), .A2(new_n343), .ZN(new_n769));
  AND4_X1   g568(.A1(KEYINPUT51), .A2(new_n740), .A3(new_n306), .A4(new_n769), .ZN(new_n770));
  AOI21_X1  g569(.A(KEYINPUT51), .B1(new_n703), .B2(new_n769), .ZN(new_n771));
  OAI21_X1  g570(.A(new_n768), .B1(new_n770), .B2(new_n771), .ZN(new_n772));
  NAND2_X1  g571(.A1(new_n769), .A2(new_n365), .ZN(new_n773));
  AOI21_X1  g572(.A(new_n773), .B1(new_n696), .B2(new_n705), .ZN(new_n774));
  AND2_X1   g573(.A1(new_n774), .A2(new_n618), .ZN(new_n775));
  OAI21_X1  g574(.A(new_n772), .B1(new_n775), .B2(new_n275), .ZN(G1336gat));
  INV_X1    g575(.A(new_n773), .ZN(new_n777));
  OAI211_X1 g576(.A(new_n659), .B(new_n777), .C1(new_n727), .C2(new_n729), .ZN(new_n778));
  NAND2_X1  g577(.A1(new_n778), .A2(G92gat), .ZN(new_n779));
  NOR3_X1   g578(.A1(new_n649), .A2(G92gat), .A3(new_n366), .ZN(new_n780));
  OAI21_X1  g579(.A(new_n780), .B1(new_n770), .B2(new_n771), .ZN(new_n781));
  XNOR2_X1  g580(.A(KEYINPUT113), .B(KEYINPUT52), .ZN(new_n782));
  AND3_X1   g581(.A1(new_n779), .A2(new_n781), .A3(new_n782), .ZN(new_n783));
  AOI21_X1  g582(.A(new_n782), .B1(new_n779), .B2(new_n781), .ZN(new_n784));
  NOR2_X1   g583(.A1(new_n783), .A2(new_n784), .ZN(G1337gat));
  NAND3_X1  g584(.A1(new_n706), .A2(new_n673), .A3(new_n777), .ZN(new_n786));
  NAND2_X1  g585(.A1(new_n786), .A2(KEYINPUT114), .ZN(new_n787));
  INV_X1    g586(.A(KEYINPUT114), .ZN(new_n788));
  NAND3_X1  g587(.A1(new_n774), .A2(new_n788), .A3(new_n673), .ZN(new_n789));
  NAND3_X1  g588(.A1(new_n787), .A2(G99gat), .A3(new_n789), .ZN(new_n790));
  NOR3_X1   g589(.A1(new_n678), .A2(G99gat), .A3(new_n366), .ZN(new_n791));
  OAI21_X1  g590(.A(new_n791), .B1(new_n770), .B2(new_n771), .ZN(new_n792));
  NAND2_X1  g591(.A1(new_n790), .A2(new_n792), .ZN(G1338gat));
  OAI211_X1 g592(.A(new_n613), .B(new_n777), .C1(new_n727), .C2(new_n729), .ZN(new_n794));
  NAND2_X1  g593(.A1(new_n794), .A2(G106gat), .ZN(new_n795));
  NOR2_X1   g594(.A1(new_n366), .A2(G106gat), .ZN(new_n796));
  OAI211_X1 g595(.A(new_n613), .B(new_n796), .C1(new_n770), .C2(new_n771), .ZN(new_n797));
  NAND2_X1  g596(.A1(new_n795), .A2(new_n797), .ZN(new_n798));
  NAND2_X1  g597(.A1(new_n798), .A2(KEYINPUT53), .ZN(new_n799));
  INV_X1    g598(.A(KEYINPUT53), .ZN(new_n800));
  NAND3_X1  g599(.A1(new_n795), .A2(new_n797), .A3(new_n800), .ZN(new_n801));
  NAND2_X1  g600(.A1(new_n799), .A2(new_n801), .ZN(G1339gat));
  INV_X1    g601(.A(KEYINPUT54), .ZN(new_n803));
  NAND3_X1  g602(.A1(new_n353), .A2(new_n803), .A3(new_n354), .ZN(new_n804));
  NAND2_X1  g603(.A1(new_n804), .A2(new_n361), .ZN(new_n805));
  INV_X1    g604(.A(KEYINPUT115), .ZN(new_n806));
  AND3_X1   g605(.A1(new_n344), .A2(new_n345), .A3(new_n350), .ZN(new_n807));
  INV_X1    g606(.A(new_n354), .ZN(new_n808));
  OAI21_X1  g607(.A(new_n808), .B1(new_n350), .B2(new_n345), .ZN(new_n809));
  OAI21_X1  g608(.A(KEYINPUT54), .B1(new_n807), .B2(new_n809), .ZN(new_n810));
  AOI21_X1  g609(.A(new_n808), .B1(new_n351), .B2(new_n352), .ZN(new_n811));
  OAI21_X1  g610(.A(new_n806), .B1(new_n810), .B2(new_n811), .ZN(new_n812));
  AND4_X1   g611(.A1(new_n347), .A2(new_n282), .A3(new_n349), .A4(new_n284), .ZN(new_n813));
  AOI21_X1  g612(.A(new_n354), .B1(new_n813), .B2(KEYINPUT10), .ZN(new_n814));
  AOI21_X1  g613(.A(new_n803), .B1(new_n814), .B2(new_n351), .ZN(new_n815));
  NAND3_X1  g614(.A1(new_n355), .A2(new_n815), .A3(KEYINPUT115), .ZN(new_n816));
  AOI21_X1  g615(.A(new_n805), .B1(new_n812), .B2(new_n816), .ZN(new_n817));
  AOI21_X1  g616(.A(new_n362), .B1(new_n817), .B2(KEYINPUT55), .ZN(new_n818));
  AOI21_X1  g617(.A(new_n360), .B1(new_n811), .B2(new_n803), .ZN(new_n819));
  NOR3_X1   g618(.A1(new_n810), .A2(new_n806), .A3(new_n811), .ZN(new_n820));
  AOI21_X1  g619(.A(KEYINPUT115), .B1(new_n355), .B2(new_n815), .ZN(new_n821));
  OAI21_X1  g620(.A(new_n819), .B1(new_n820), .B2(new_n821), .ZN(new_n822));
  INV_X1    g621(.A(KEYINPUT55), .ZN(new_n823));
  NAND2_X1  g622(.A1(new_n822), .A2(new_n823), .ZN(new_n824));
  NAND3_X1  g623(.A1(new_n343), .A2(new_n818), .A3(new_n824), .ZN(new_n825));
  INV_X1    g624(.A(new_n337), .ZN(new_n826));
  NAND3_X1  g625(.A1(new_n341), .A2(new_n826), .A3(new_n328), .ZN(new_n827));
  NOR2_X1   g626(.A1(new_n322), .A2(new_n311), .ZN(new_n828));
  AOI21_X1  g627(.A(new_n312), .B1(new_n310), .B2(new_n314), .ZN(new_n829));
  OAI21_X1  g628(.A(new_n336), .B1(new_n828), .B2(new_n829), .ZN(new_n830));
  NAND3_X1  g629(.A1(new_n827), .A2(new_n365), .A3(new_n830), .ZN(new_n831));
  AOI21_X1  g630(.A(new_n306), .B1(new_n825), .B2(new_n831), .ZN(new_n832));
  NAND3_X1  g631(.A1(new_n306), .A2(new_n818), .A3(new_n824), .ZN(new_n833));
  AND3_X1   g632(.A1(new_n827), .A2(KEYINPUT116), .A3(new_n830), .ZN(new_n834));
  AOI21_X1  g633(.A(KEYINPUT116), .B1(new_n827), .B2(new_n830), .ZN(new_n835));
  NOR3_X1   g634(.A1(new_n833), .A2(new_n834), .A3(new_n835), .ZN(new_n836));
  OAI21_X1  g635(.A(new_n244), .B1(new_n832), .B2(new_n836), .ZN(new_n837));
  NAND3_X1  g636(.A1(new_n307), .A2(new_n689), .A3(new_n366), .ZN(new_n838));
  NAND2_X1  g637(.A1(new_n837), .A2(new_n838), .ZN(new_n839));
  NAND2_X1  g638(.A1(new_n839), .A2(new_n747), .ZN(new_n840));
  NOR3_X1   g639(.A1(new_n840), .A2(new_n613), .A3(new_n612), .ZN(new_n841));
  AND2_X1   g640(.A1(new_n841), .A2(new_n649), .ZN(new_n842));
  NOR2_X1   g641(.A1(new_n689), .A2(G113gat), .ZN(new_n843));
  XNOR2_X1  g642(.A(new_n843), .B(KEYINPUT117), .ZN(new_n844));
  NAND2_X1  g643(.A1(new_n842), .A2(new_n844), .ZN(new_n845));
  NOR2_X1   g644(.A1(new_n648), .A2(new_n659), .ZN(new_n846));
  NAND4_X1  g645(.A1(new_n677), .A2(new_n569), .A3(new_n839), .A4(new_n846), .ZN(new_n847));
  OAI21_X1  g646(.A(G113gat), .B1(new_n847), .B2(new_n689), .ZN(new_n848));
  NAND2_X1  g647(.A1(new_n845), .A2(new_n848), .ZN(G1340gat));
  INV_X1    g648(.A(G120gat), .ZN(new_n850));
  NOR3_X1   g649(.A1(new_n847), .A2(new_n850), .A3(new_n366), .ZN(new_n851));
  NAND2_X1  g650(.A1(new_n842), .A2(new_n365), .ZN(new_n852));
  AOI21_X1  g651(.A(new_n851), .B1(new_n852), .B2(new_n850), .ZN(G1341gat));
  NOR2_X1   g652(.A1(new_n244), .A2(new_n407), .ZN(new_n854));
  NAND2_X1  g653(.A1(new_n842), .A2(new_n854), .ZN(new_n855));
  OAI21_X1  g654(.A(new_n407), .B1(new_n847), .B2(new_n244), .ZN(new_n856));
  NAND2_X1  g655(.A1(new_n855), .A2(new_n856), .ZN(G1342gat));
  NOR3_X1   g656(.A1(new_n659), .A2(G134gat), .A3(new_n697), .ZN(new_n858));
  NAND2_X1  g657(.A1(new_n841), .A2(new_n858), .ZN(new_n859));
  NAND2_X1  g658(.A1(new_n859), .A2(KEYINPUT56), .ZN(new_n860));
  XNOR2_X1  g659(.A(new_n860), .B(KEYINPUT118), .ZN(new_n861));
  OAI21_X1  g660(.A(G134gat), .B1(new_n847), .B2(new_n697), .ZN(new_n862));
  OAI211_X1 g661(.A(new_n861), .B(new_n862), .C1(KEYINPUT56), .C2(new_n859), .ZN(G1343gat));
  INV_X1    g662(.A(KEYINPUT119), .ZN(new_n864));
  OAI21_X1  g663(.A(new_n823), .B1(new_n817), .B2(new_n864), .ZN(new_n865));
  AOI211_X1 g664(.A(KEYINPUT119), .B(new_n805), .C1(new_n812), .C2(new_n816), .ZN(new_n866));
  OAI211_X1 g665(.A(KEYINPUT120), .B(new_n818), .C1(new_n865), .C2(new_n866), .ZN(new_n867));
  NAND2_X1  g666(.A1(new_n867), .A2(new_n343), .ZN(new_n868));
  NAND2_X1  g667(.A1(new_n822), .A2(KEYINPUT119), .ZN(new_n869));
  NAND2_X1  g668(.A1(new_n817), .A2(new_n864), .ZN(new_n870));
  NAND3_X1  g669(.A1(new_n869), .A2(new_n823), .A3(new_n870), .ZN(new_n871));
  AOI21_X1  g670(.A(KEYINPUT120), .B1(new_n871), .B2(new_n818), .ZN(new_n872));
  OAI21_X1  g671(.A(new_n831), .B1(new_n868), .B2(new_n872), .ZN(new_n873));
  AOI21_X1  g672(.A(new_n836), .B1(new_n873), .B2(new_n697), .ZN(new_n874));
  OAI21_X1  g673(.A(new_n838), .B1(new_n874), .B2(new_n243), .ZN(new_n875));
  AND2_X1   g674(.A1(new_n875), .A2(new_n613), .ZN(new_n876));
  NAND2_X1  g675(.A1(new_n876), .A2(KEYINPUT57), .ZN(new_n877));
  INV_X1    g676(.A(KEYINPUT121), .ZN(new_n878));
  NAND2_X1  g677(.A1(new_n839), .A2(new_n613), .ZN(new_n879));
  INV_X1    g678(.A(KEYINPUT57), .ZN(new_n880));
  AOI21_X1  g679(.A(new_n878), .B1(new_n879), .B2(new_n880), .ZN(new_n881));
  NAND2_X1  g680(.A1(new_n877), .A2(new_n881), .ZN(new_n882));
  NAND3_X1  g681(.A1(new_n876), .A2(new_n878), .A3(KEYINPUT57), .ZN(new_n883));
  AND2_X1   g682(.A1(new_n672), .A2(new_n846), .ZN(new_n884));
  NAND4_X1  g683(.A1(new_n882), .A2(new_n343), .A3(new_n883), .A4(new_n884), .ZN(new_n885));
  NAND2_X1  g684(.A1(new_n885), .A2(new_n393), .ZN(new_n886));
  NOR4_X1   g685(.A1(new_n673), .A2(new_n840), .A3(new_n659), .A4(new_n569), .ZN(new_n887));
  NAND3_X1  g686(.A1(new_n887), .A2(new_n372), .A3(new_n343), .ZN(new_n888));
  AND2_X1   g687(.A1(new_n886), .A2(new_n888), .ZN(new_n889));
  AOI21_X1  g688(.A(KEYINPUT58), .B1(new_n886), .B2(KEYINPUT122), .ZN(new_n890));
  XNOR2_X1  g689(.A(new_n889), .B(new_n890), .ZN(G1344gat));
  NAND3_X1  g690(.A1(new_n887), .A2(new_n370), .A3(new_n365), .ZN(new_n892));
  AND3_X1   g691(.A1(new_n882), .A2(new_n883), .A3(new_n884), .ZN(new_n893));
  AOI211_X1 g692(.A(KEYINPUT59), .B(new_n370), .C1(new_n893), .C2(new_n365), .ZN(new_n894));
  INV_X1    g693(.A(KEYINPUT59), .ZN(new_n895));
  AOI21_X1  g694(.A(KEYINPUT57), .B1(new_n875), .B2(new_n613), .ZN(new_n896));
  AOI211_X1 g695(.A(new_n880), .B(new_n569), .C1(new_n837), .C2(new_n838), .ZN(new_n897));
  OR2_X1    g696(.A1(new_n896), .A2(new_n897), .ZN(new_n898));
  NAND3_X1  g697(.A1(new_n898), .A2(new_n365), .A3(new_n884), .ZN(new_n899));
  AOI21_X1  g698(.A(new_n895), .B1(new_n899), .B2(G148gat), .ZN(new_n900));
  OAI21_X1  g699(.A(new_n892), .B1(new_n894), .B2(new_n900), .ZN(G1345gat));
  INV_X1    g700(.A(G155gat), .ZN(new_n902));
  NAND3_X1  g701(.A1(new_n887), .A2(new_n902), .A3(new_n243), .ZN(new_n903));
  AND2_X1   g702(.A1(new_n893), .A2(new_n243), .ZN(new_n904));
  OAI21_X1  g703(.A(new_n903), .B1(new_n904), .B2(new_n902), .ZN(G1346gat));
  XNOR2_X1  g704(.A(KEYINPUT82), .B(G162gat), .ZN(new_n906));
  NOR2_X1   g705(.A1(new_n697), .A2(new_n906), .ZN(new_n907));
  NAND2_X1  g706(.A1(new_n887), .A2(new_n907), .ZN(new_n908));
  INV_X1    g707(.A(KEYINPUT123), .ZN(new_n909));
  XNOR2_X1  g708(.A(new_n908), .B(new_n909), .ZN(new_n910));
  NAND4_X1  g709(.A1(new_n882), .A2(new_n306), .A3(new_n883), .A4(new_n884), .ZN(new_n911));
  AND2_X1   g710(.A1(new_n911), .A2(KEYINPUT124), .ZN(new_n912));
  OAI21_X1  g711(.A(new_n906), .B1(new_n911), .B2(KEYINPUT124), .ZN(new_n913));
  OAI21_X1  g712(.A(new_n910), .B1(new_n912), .B2(new_n913), .ZN(new_n914));
  INV_X1    g713(.A(KEYINPUT125), .ZN(new_n915));
  NAND2_X1  g714(.A1(new_n914), .A2(new_n915), .ZN(new_n916));
  OAI211_X1 g715(.A(new_n910), .B(KEYINPUT125), .C1(new_n912), .C2(new_n913), .ZN(new_n917));
  NAND2_X1  g716(.A1(new_n916), .A2(new_n917), .ZN(G1347gat));
  NAND2_X1  g717(.A1(new_n839), .A2(new_n648), .ZN(new_n919));
  INV_X1    g718(.A(new_n919), .ZN(new_n920));
  NOR3_X1   g719(.A1(new_n612), .A2(new_n649), .A3(new_n613), .ZN(new_n921));
  NAND2_X1  g720(.A1(new_n920), .A2(new_n921), .ZN(new_n922));
  INV_X1    g721(.A(new_n922), .ZN(new_n923));
  AOI21_X1  g722(.A(G169gat), .B1(new_n923), .B2(new_n343), .ZN(new_n924));
  NAND3_X1  g723(.A1(new_n745), .A2(new_n659), .A3(new_n746), .ZN(new_n925));
  AOI211_X1 g724(.A(new_n613), .B(new_n925), .C1(new_n837), .C2(new_n838), .ZN(new_n926));
  AND2_X1   g725(.A1(new_n756), .A2(new_n926), .ZN(new_n927));
  AND2_X1   g726(.A1(new_n343), .A2(G169gat), .ZN(new_n928));
  AOI21_X1  g727(.A(new_n924), .B1(new_n927), .B2(new_n928), .ZN(G1348gat));
  INV_X1    g728(.A(G176gat), .ZN(new_n930));
  NAND3_X1  g729(.A1(new_n923), .A2(new_n930), .A3(new_n365), .ZN(new_n931));
  NAND2_X1  g730(.A1(new_n927), .A2(new_n365), .ZN(new_n932));
  INV_X1    g731(.A(new_n932), .ZN(new_n933));
  OAI21_X1  g732(.A(new_n931), .B1(new_n933), .B2(new_n930), .ZN(G1349gat));
  AND3_X1   g733(.A1(new_n923), .A2(new_n480), .A3(new_n243), .ZN(new_n935));
  NAND2_X1  g734(.A1(new_n927), .A2(new_n243), .ZN(new_n936));
  AOI21_X1  g735(.A(new_n935), .B1(new_n936), .B2(G183gat), .ZN(new_n937));
  XOR2_X1   g736(.A(new_n937), .B(KEYINPUT60), .Z(G1350gat));
  NAND3_X1  g737(.A1(new_n923), .A2(new_n481), .A3(new_n306), .ZN(new_n939));
  NAND2_X1  g738(.A1(new_n927), .A2(new_n306), .ZN(new_n940));
  NAND2_X1  g739(.A1(new_n940), .A2(G190gat), .ZN(new_n941));
  AND2_X1   g740(.A1(new_n941), .A2(KEYINPUT61), .ZN(new_n942));
  NOR2_X1   g741(.A1(new_n941), .A2(KEYINPUT61), .ZN(new_n943));
  OAI21_X1  g742(.A(new_n939), .B1(new_n942), .B2(new_n943), .ZN(G1351gat));
  NOR4_X1   g743(.A1(new_n673), .A2(new_n919), .A3(new_n649), .A4(new_n569), .ZN(new_n945));
  AOI21_X1  g744(.A(G197gat), .B1(new_n945), .B2(new_n343), .ZN(new_n946));
  AOI21_X1  g745(.A(new_n925), .B1(new_n671), .B2(new_n653), .ZN(new_n947));
  AND2_X1   g746(.A1(new_n898), .A2(new_n947), .ZN(new_n948));
  AND2_X1   g747(.A1(new_n343), .A2(G197gat), .ZN(new_n949));
  AOI21_X1  g748(.A(new_n946), .B1(new_n948), .B2(new_n949), .ZN(G1352gat));
  INV_X1    g749(.A(G204gat), .ZN(new_n951));
  NAND3_X1  g750(.A1(new_n945), .A2(new_n951), .A3(new_n365), .ZN(new_n952));
  XOR2_X1   g751(.A(new_n952), .B(KEYINPUT62), .Z(new_n953));
  NAND2_X1  g752(.A1(new_n948), .A2(new_n365), .ZN(new_n954));
  INV_X1    g753(.A(new_n954), .ZN(new_n955));
  OAI21_X1  g754(.A(new_n953), .B1(new_n951), .B2(new_n955), .ZN(G1353gat));
  INV_X1    g755(.A(KEYINPUT63), .ZN(new_n957));
  OAI211_X1 g756(.A(new_n243), .B(new_n947), .C1(new_n896), .C2(new_n897), .ZN(new_n958));
  AND2_X1   g757(.A1(new_n958), .A2(KEYINPUT126), .ZN(new_n959));
  OAI21_X1  g758(.A(G211gat), .B1(new_n958), .B2(KEYINPUT126), .ZN(new_n960));
  OAI21_X1  g759(.A(new_n957), .B1(new_n959), .B2(new_n960), .ZN(new_n961));
  INV_X1    g760(.A(KEYINPUT126), .ZN(new_n962));
  NAND4_X1  g761(.A1(new_n898), .A2(new_n962), .A3(new_n243), .A4(new_n947), .ZN(new_n963));
  NAND2_X1  g762(.A1(new_n958), .A2(KEYINPUT126), .ZN(new_n964));
  NAND4_X1  g763(.A1(new_n963), .A2(KEYINPUT63), .A3(new_n964), .A4(G211gat), .ZN(new_n965));
  NAND2_X1  g764(.A1(new_n961), .A2(new_n965), .ZN(new_n966));
  INV_X1    g765(.A(G211gat), .ZN(new_n967));
  NAND3_X1  g766(.A1(new_n945), .A2(new_n967), .A3(new_n243), .ZN(new_n968));
  NAND2_X1  g767(.A1(new_n966), .A2(new_n968), .ZN(new_n969));
  INV_X1    g768(.A(KEYINPUT127), .ZN(new_n970));
  NAND2_X1  g769(.A1(new_n969), .A2(new_n970), .ZN(new_n971));
  NAND3_X1  g770(.A1(new_n966), .A2(KEYINPUT127), .A3(new_n968), .ZN(new_n972));
  NAND2_X1  g771(.A1(new_n971), .A2(new_n972), .ZN(G1354gat));
  INV_X1    g772(.A(G218gat), .ZN(new_n974));
  AOI21_X1  g773(.A(new_n974), .B1(new_n948), .B2(new_n306), .ZN(new_n975));
  AND3_X1   g774(.A1(new_n945), .A2(new_n974), .A3(new_n306), .ZN(new_n976));
  OR2_X1    g775(.A1(new_n975), .A2(new_n976), .ZN(G1355gat));
endmodule


