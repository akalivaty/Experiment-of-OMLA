

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n359, n360, n361, n362, n363, n364, n365, n366, n367, n369, n370,
         n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381,
         n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392,
         n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403,
         n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414,
         n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425,
         n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436,
         n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447,
         n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458,
         n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469,
         n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480,
         n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491,
         n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502,
         n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n513,
         n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
         n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
         n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590,
         n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601,
         n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612,
         n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623,
         n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634,
         n635, n636, n637, n638, n639, n640, n641, n642, n643, n644, n645,
         n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, n656,
         n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n667,
         n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678,
         n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689,
         n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700,
         n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711,
         n712, n713, n714, n715, n716, n717, n718, n719, n720, n721, n722,
         n723, n724, n725, n726, n727, n728, n729, n730, n731, n732, n733,
         n734, n735, n736, n737, n738, n739, n740, n741, n742, n743, n744,
         n745, n746, n747, n748, n749, n750, n751, n752, n753, n754, n755,
         n756, n757, n758, n759, n760, n761, n762, n763, n764, n765, n766,
         n767, n768, n769, n770, n771, n772, n773, n774, n775, n776, n777,
         n778, n779, n780, n781, n782, n783, n784, n785, n786, n787, n788,
         n789, n790, n791, n792, n793, n794, n795, n796;

  BUF_X1 U380 ( .A(n701), .Z(n787) );
  NOR2_X1 U381 ( .A1(n556), .A2(n619), .ZN(n755) );
  NOR2_X1 U382 ( .A1(G953), .A2(G237), .ZN(n511) );
  XNOR2_X1 U383 ( .A(n649), .B(n640), .ZN(n701) );
  AND2_X2 U384 ( .A1(n711), .A2(n710), .ZN(n758) );
  INV_X1 U385 ( .A(G953), .ZN(n788) );
  XOR2_X1 U386 ( .A(KEYINPUT69), .B(n461), .Z(n359) );
  XNOR2_X2 U387 ( .A(n633), .B(n584), .ZN(n681) );
  XNOR2_X2 U388 ( .A(n552), .B(n425), .ZN(n756) );
  XNOR2_X2 U389 ( .A(n597), .B(KEYINPUT108), .ZN(n753) );
  AND2_X2 U390 ( .A1(n599), .A2(n598), .ZN(n600) );
  XNOR2_X2 U391 ( .A(n589), .B(n528), .ZN(n599) );
  AND2_X1 U392 ( .A1(n551), .A2(n673), .ZN(n552) );
  INV_X2 U393 ( .A(G125), .ZN(n404) );
  NOR2_X1 U394 ( .A1(n740), .A2(n769), .ZN(n741) );
  NOR2_X1 U395 ( .A1(n697), .A2(n696), .ZN(n698) );
  NOR2_X1 U396 ( .A1(n733), .A2(n769), .ZN(n735) );
  NAND2_X1 U397 ( .A1(n709), .A2(n371), .ZN(n711) );
  OR2_X1 U398 ( .A1(n787), .A2(n651), .ZN(n642) );
  AND2_X1 U399 ( .A1(n701), .A2(n700), .ZN(n702) );
  BUF_X1 U400 ( .A(n703), .Z(n770) );
  NOR2_X1 U401 ( .A1(n567), .A2(n569), .ZN(n570) );
  AND2_X1 U402 ( .A1(n562), .A2(n561), .ZN(n563) );
  AND2_X1 U403 ( .A1(n725), .A2(n629), .ZN(n374) );
  NOR2_X1 U404 ( .A1(n721), .A2(n796), .ZN(n596) );
  NAND2_X1 U405 ( .A1(n409), .A2(n407), .ZN(n721) );
  NAND2_X1 U406 ( .A1(n408), .A2(n367), .ZN(n407) );
  NAND2_X1 U407 ( .A1(n383), .A2(n387), .ZN(n604) );
  XNOR2_X1 U408 ( .A(n555), .B(n554), .ZN(n744) );
  AND2_X1 U409 ( .A1(n386), .A2(n384), .ZN(n383) );
  NAND2_X1 U410 ( .A1(n582), .A2(n360), .ZN(n623) );
  NAND2_X1 U411 ( .A1(n410), .A2(KEYINPUT40), .ZN(n405) );
  XNOR2_X1 U412 ( .A(n400), .B(n510), .ZN(n535) );
  BUF_X2 U413 ( .A(n575), .Z(n589) );
  XNOR2_X1 U414 ( .A(n442), .B(n441), .ZN(n583) );
  XNOR2_X1 U415 ( .A(n479), .B(n478), .ZN(n620) );
  XNOR2_X1 U416 ( .A(n403), .B(n468), .ZN(n784) );
  XNOR2_X1 U417 ( .A(n516), .B(KEYINPUT16), .ZN(n429) );
  XNOR2_X1 U418 ( .A(n459), .B(KEYINPUT4), .ZN(n494) );
  NOR2_X1 U419 ( .A1(n381), .A2(G953), .ZN(n380) );
  INV_X1 U420 ( .A(KEYINPUT31), .ZN(n425) );
  NAND2_X1 U421 ( .A1(n376), .A2(n639), .ZN(n649) );
  AND2_X1 U422 ( .A1(n422), .A2(n421), .ZN(n420) );
  NOR2_X1 U423 ( .A1(n606), .A2(n419), .ZN(n418) );
  XNOR2_X1 U424 ( .A(n382), .B(n380), .ZN(n461) );
  XNOR2_X1 U425 ( .A(KEYINPUT8), .B(KEYINPUT68), .ZN(n382) );
  AND2_X1 U426 ( .A1(n662), .A2(n661), .ZN(n433) );
  NAND2_X1 U427 ( .A1(n413), .A2(n412), .ZN(n411) );
  INV_X1 U428 ( .A(n623), .ZN(n413) );
  AND2_X1 U429 ( .A1(n416), .A2(n415), .ZN(n414) );
  NAND2_X1 U430 ( .A1(n623), .A2(n417), .ZN(n416) );
  XNOR2_X1 U431 ( .A(n458), .B(n457), .ZN(n460) );
  XNOR2_X1 U432 ( .A(G122), .B(G134), .ZN(n457) );
  OR2_X1 U433 ( .A1(n753), .A2(n389), .ZN(n386) );
  AND2_X1 U434 ( .A1(n600), .A2(n389), .ZN(n385) );
  AND2_X1 U435 ( .A1(n388), .A2(n602), .ZN(n387) );
  NAND2_X1 U436 ( .A1(n730), .A2(n507), .ZN(n479) );
  XNOR2_X1 U437 ( .A(n466), .B(n378), .ZN(n377) );
  OR2_X1 U438 ( .A1(n766), .A2(G902), .ZN(n379) );
  NOR2_X1 U439 ( .A1(n756), .A2(KEYINPUT99), .ZN(n423) );
  AND2_X1 U440 ( .A1(n560), .A2(n430), .ZN(n561) );
  INV_X1 U441 ( .A(G234), .ZN(n381) );
  NOR2_X1 U442 ( .A1(n597), .A2(n755), .ZN(n390) );
  INV_X1 U443 ( .A(KEYINPUT39), .ZN(n417) );
  XNOR2_X1 U444 ( .A(G104), .B(G143), .ZN(n471) );
  XNOR2_X1 U445 ( .A(n494), .B(n493), .ZN(n785) );
  XNOR2_X1 U446 ( .A(G134), .B(G131), .ZN(n492) );
  OR2_X1 U447 ( .A1(G902), .A2(G237), .ZN(n431) );
  NOR2_X1 U448 ( .A1(n681), .A2(n680), .ZN(n685) );
  INV_X1 U449 ( .A(KEYINPUT110), .ZN(n389) );
  INV_X1 U450 ( .A(G478), .ZN(n378) );
  INV_X1 U451 ( .A(KEYINPUT67), .ZN(n398) );
  NOR2_X2 U452 ( .A1(n535), .A2(n665), .ZN(n399) );
  XNOR2_X1 U453 ( .A(G116), .B(G113), .ZN(n512) );
  XNOR2_X1 U454 ( .A(G137), .B(G119), .ZN(n501) );
  XNOR2_X1 U455 ( .A(n467), .B(G140), .ZN(n403) );
  XNOR2_X1 U456 ( .A(n477), .B(n391), .ZN(n730) );
  XNOR2_X1 U457 ( .A(n784), .B(n392), .ZN(n391) );
  XNOR2_X1 U458 ( .A(n476), .B(n475), .ZN(n477) );
  XNOR2_X1 U459 ( .A(n470), .B(n471), .ZN(n392) );
  XNOR2_X1 U460 ( .A(n785), .B(G146), .ZN(n521) );
  XNOR2_X1 U461 ( .A(n427), .B(KEYINPUT90), .ZN(n426) );
  XNOR2_X1 U462 ( .A(n396), .B(KEYINPUT41), .ZN(n677) );
  NAND2_X1 U463 ( .A1(n682), .A2(n685), .ZN(n396) );
  NAND2_X1 U464 ( .A1(n414), .A2(n411), .ZN(n636) );
  NAND2_X1 U465 ( .A1(n361), .A2(n414), .ZN(n406) );
  BUF_X1 U466 ( .A(n535), .Z(n666) );
  XNOR2_X1 U467 ( .A(G110), .B(G104), .ZN(n434) );
  XNOR2_X1 U468 ( .A(n465), .B(n464), .ZN(n766) );
  BUF_X1 U469 ( .A(n758), .Z(n765) );
  XNOR2_X1 U470 ( .A(n544), .B(n543), .ZN(n728) );
  NOR2_X1 U471 ( .A1(n581), .A2(n587), .ZN(n360) );
  INV_X1 U472 ( .A(n606), .ZN(n684) );
  XNOR2_X1 U473 ( .A(n390), .B(KEYINPUT104), .ZN(n606) );
  AND2_X1 U474 ( .A1(n411), .A2(n410), .ZN(n361) );
  XOR2_X1 U475 ( .A(n459), .B(KEYINPUT9), .Z(n362) );
  AND2_X1 U476 ( .A1(n508), .A2(G217), .ZN(n363) );
  XOR2_X1 U477 ( .A(n531), .B(KEYINPUT80), .Z(n364) );
  AND2_X1 U478 ( .A1(n753), .A2(n600), .ZN(n365) );
  AND2_X1 U479 ( .A1(n619), .A2(n556), .ZN(n597) );
  NOR2_X1 U480 ( .A1(n661), .A2(n526), .ZN(n366) );
  AND2_X1 U481 ( .A1(n597), .A2(KEYINPUT40), .ZN(n367) );
  XOR2_X1 U482 ( .A(KEYINPUT53), .B(n699), .Z(G75) );
  NOR2_X1 U483 ( .A1(n557), .A2(n599), .ZN(n369) );
  XNOR2_X1 U484 ( .A(n485), .B(KEYINPUT22), .ZN(n370) );
  XOR2_X1 U485 ( .A(n708), .B(KEYINPUT65), .Z(n371) );
  XOR2_X1 U486 ( .A(n712), .B(KEYINPUT62), .Z(n372) );
  XNOR2_X1 U487 ( .A(n596), .B(KEYINPUT46), .ZN(n375) );
  XNOR2_X1 U488 ( .A(n373), .B(n630), .ZN(n376) );
  NAND2_X1 U489 ( .A1(n375), .A2(n374), .ZN(n373) );
  XNOR2_X2 U490 ( .A(n379), .B(n377), .ZN(n619) );
  NAND2_X1 U491 ( .A1(n753), .A2(n385), .ZN(n384) );
  OR2_X1 U492 ( .A1(n600), .A2(n389), .ZN(n388) );
  INV_X2 U493 ( .A(G116), .ZN(n395) );
  XNOR2_X2 U494 ( .A(n393), .B(n429), .ZN(n776) );
  XNOR2_X2 U495 ( .A(n458), .B(n469), .ZN(n393) );
  XNOR2_X2 U496 ( .A(n394), .B(G122), .ZN(n469) );
  XNOR2_X2 U497 ( .A(n395), .B(G107), .ZN(n458) );
  INV_X2 U498 ( .A(G113), .ZN(n394) );
  NAND2_X1 U499 ( .A1(n397), .A2(n366), .ZN(n527) );
  NAND2_X1 U500 ( .A1(n397), .A2(n364), .ZN(n534) );
  AND2_X1 U501 ( .A1(n397), .A2(n369), .ZN(n742) );
  XNOR2_X2 U502 ( .A(n486), .B(n370), .ZN(n397) );
  XNOR2_X2 U503 ( .A(n538), .B(n537), .ZN(n688) );
  XNOR2_X2 U504 ( .A(n496), .B(G469), .ZN(n592) );
  XNOR2_X2 U505 ( .A(n399), .B(n398), .ZN(n662) );
  NAND2_X1 U506 ( .A1(n717), .A2(n507), .ZN(n400) );
  XNOR2_X1 U507 ( .A(n401), .B(KEYINPUT63), .ZN(G57) );
  NAND2_X1 U508 ( .A1(n402), .A2(n715), .ZN(n401) );
  XNOR2_X1 U509 ( .A(n713), .B(n372), .ZN(n402) );
  XNOR2_X2 U510 ( .A(n404), .B(G146), .ZN(n467) );
  NAND2_X1 U511 ( .A1(n406), .A2(n405), .ZN(n409) );
  INV_X1 U512 ( .A(n636), .ZN(n408) );
  NAND2_X1 U513 ( .A1(n585), .A2(n586), .ZN(n410) );
  NOR2_X1 U514 ( .A1(n681), .A2(n417), .ZN(n412) );
  NAND2_X1 U515 ( .A1(n681), .A2(n417), .ZN(n415) );
  NAND2_X1 U516 ( .A1(n420), .A2(n418), .ZN(n560) );
  AND2_X1 U517 ( .A1(n756), .A2(KEYINPUT99), .ZN(n419) );
  NAND2_X1 U518 ( .A1(n744), .A2(KEYINPUT99), .ZN(n421) );
  NAND2_X1 U519 ( .A1(n424), .A2(n423), .ZN(n422) );
  INV_X1 U520 ( .A(n744), .ZN(n424) );
  XNOR2_X1 U521 ( .A(n428), .B(n426), .ZN(n437) );
  NAND2_X1 U522 ( .A1(n788), .A2(G224), .ZN(n427) );
  XNOR2_X1 U523 ( .A(n467), .B(n436), .ZN(n428) );
  XNOR2_X2 U524 ( .A(KEYINPUT3), .B(G119), .ZN(n516) );
  NAND2_X1 U525 ( .A1(n718), .A2(n715), .ZN(n719) );
  XNOR2_X1 U526 ( .A(n717), .B(n716), .ZN(n718) );
  NAND2_X1 U527 ( .A1(n758), .A2(G217), .ZN(n716) );
  XNOR2_X1 U528 ( .A(n601), .B(n447), .ZN(n607) );
  NAND2_X1 U529 ( .A1(n446), .A2(n445), .ZN(n601) );
  INV_X1 U530 ( .A(n583), .ZN(n446) );
  AND2_X1 U531 ( .A1(n559), .A2(n558), .ZN(n430) );
  XOR2_X1 U532 ( .A(n588), .B(KEYINPUT71), .Z(n432) );
  INV_X1 U533 ( .A(n769), .ZN(n715) );
  INV_X1 U534 ( .A(n469), .ZN(n470) );
  INV_X1 U535 ( .A(KEYINPUT85), .ZN(n704) );
  INV_X1 U536 ( .A(n680), .ZN(n445) );
  INV_X1 U537 ( .A(KEYINPUT103), .ZN(n466) );
  XNOR2_X1 U538 ( .A(n460), .B(n362), .ZN(n463) );
  XNOR2_X1 U539 ( .A(n463), .B(n462), .ZN(n465) );
  XNOR2_X1 U540 ( .A(n434), .B(KEYINPUT89), .ZN(n778) );
  XNOR2_X2 U541 ( .A(KEYINPUT66), .B(G101), .ZN(n514) );
  XNOR2_X1 U542 ( .A(n514), .B(KEYINPUT73), .ZN(n435) );
  XNOR2_X1 U543 ( .A(n778), .B(n435), .ZN(n490) );
  XNOR2_X1 U544 ( .A(n776), .B(n490), .ZN(n439) );
  XNOR2_X1 U545 ( .A(KEYINPUT17), .B(KEYINPUT18), .ZN(n436) );
  XNOR2_X2 U546 ( .A(G143), .B(G128), .ZN(n459) );
  XNOR2_X1 U547 ( .A(n437), .B(n494), .ZN(n438) );
  XNOR2_X1 U548 ( .A(n439), .B(n438), .ZN(n736) );
  XNOR2_X1 U549 ( .A(G902), .B(KEYINPUT88), .ZN(n440) );
  XNOR2_X1 U550 ( .A(n440), .B(KEYINPUT15), .ZN(n707) );
  NAND2_X1 U551 ( .A1(n736), .A2(n707), .ZN(n442) );
  XNOR2_X1 U552 ( .A(KEYINPUT76), .B(n431), .ZN(n443) );
  NAND2_X1 U553 ( .A1(n443), .A2(G210), .ZN(n441) );
  NAND2_X1 U554 ( .A1(n443), .A2(G214), .ZN(n444) );
  XNOR2_X1 U555 ( .A(n444), .B(KEYINPUT91), .ZN(n680) );
  INV_X1 U556 ( .A(KEYINPUT19), .ZN(n447) );
  XOR2_X1 U557 ( .A(KEYINPUT92), .B(KEYINPUT14), .Z(n449) );
  NAND2_X1 U558 ( .A1(G237), .A2(G234), .ZN(n448) );
  XNOR2_X1 U559 ( .A(n449), .B(n448), .ZN(n450) );
  XNOR2_X1 U560 ( .A(KEYINPUT75), .B(n450), .ZN(n453) );
  NAND2_X1 U561 ( .A1(n453), .A2(G902), .ZN(n451) );
  XNOR2_X1 U562 ( .A(n451), .B(KEYINPUT93), .ZN(n577) );
  NOR2_X1 U563 ( .A1(G898), .A2(n788), .ZN(n781) );
  NAND2_X1 U564 ( .A1(n577), .A2(n781), .ZN(n452) );
  XNOR2_X1 U565 ( .A(n452), .B(KEYINPUT94), .ZN(n454) );
  NAND2_X1 U566 ( .A1(G952), .A2(n453), .ZN(n694) );
  OR2_X1 U567 ( .A1(n694), .A2(G953), .ZN(n579) );
  AND2_X1 U568 ( .A1(n454), .A2(n579), .ZN(n455) );
  NOR2_X2 U569 ( .A1(n607), .A2(n455), .ZN(n456) );
  XNOR2_X2 U570 ( .A(n456), .B(KEYINPUT0), .ZN(n551) );
  NAND2_X1 U571 ( .A1(G217), .A2(n359), .ZN(n462) );
  XNOR2_X1 U572 ( .A(KEYINPUT102), .B(KEYINPUT7), .ZN(n464) );
  XOR2_X1 U573 ( .A(KEYINPUT70), .B(KEYINPUT10), .Z(n468) );
  XOR2_X1 U574 ( .A(KEYINPUT101), .B(KEYINPUT100), .Z(n473) );
  NAND2_X1 U575 ( .A1(n511), .A2(G214), .ZN(n472) );
  XNOR2_X1 U576 ( .A(n473), .B(n472), .ZN(n474) );
  XOR2_X1 U577 ( .A(n474), .B(KEYINPUT12), .Z(n476) );
  XOR2_X1 U578 ( .A(KEYINPUT11), .B(G131), .Z(n475) );
  INV_X1 U579 ( .A(G902), .ZN(n507) );
  XNOR2_X1 U580 ( .A(KEYINPUT13), .B(G475), .ZN(n478) );
  AND2_X1 U581 ( .A1(n619), .A2(n620), .ZN(n682) );
  NAND2_X1 U582 ( .A1(n707), .A2(G234), .ZN(n480) );
  XNOR2_X1 U583 ( .A(n480), .B(KEYINPUT20), .ZN(n508) );
  AND2_X1 U584 ( .A1(n508), .A2(G221), .ZN(n482) );
  INV_X1 U585 ( .A(KEYINPUT21), .ZN(n481) );
  XNOR2_X1 U586 ( .A(n482), .B(n481), .ZN(n665) );
  INV_X1 U587 ( .A(n665), .ZN(n483) );
  AND2_X1 U588 ( .A1(n682), .A2(n483), .ZN(n484) );
  NAND2_X1 U589 ( .A1(n551), .A2(n484), .ZN(n486) );
  INV_X1 U590 ( .A(KEYINPUT74), .ZN(n485) );
  XOR2_X1 U591 ( .A(G140), .B(G107), .Z(n488) );
  NAND2_X1 U592 ( .A1(G227), .A2(n788), .ZN(n487) );
  XNOR2_X1 U593 ( .A(n488), .B(n487), .ZN(n489) );
  XNOR2_X1 U594 ( .A(n490), .B(n489), .ZN(n495) );
  INV_X1 U595 ( .A(G137), .ZN(n491) );
  XNOR2_X1 U596 ( .A(n492), .B(n491), .ZN(n493) );
  XNOR2_X1 U597 ( .A(n495), .B(n521), .ZN(n761) );
  NAND2_X1 U598 ( .A1(n761), .A2(n507), .ZN(n496) );
  XNOR2_X2 U599 ( .A(n592), .B(KEYINPUT1), .ZN(n661) );
  XOR2_X1 U600 ( .A(G128), .B(G110), .Z(n498) );
  XNOR2_X1 U601 ( .A(KEYINPUT72), .B(KEYINPUT23), .ZN(n497) );
  XNOR2_X1 U602 ( .A(n498), .B(n497), .ZN(n499) );
  XNOR2_X1 U603 ( .A(KEYINPUT24), .B(n499), .ZN(n500) );
  XNOR2_X1 U604 ( .A(n784), .B(n500), .ZN(n506) );
  NAND2_X1 U605 ( .A1(G221), .A2(n359), .ZN(n504) );
  XOR2_X1 U606 ( .A(KEYINPUT95), .B(KEYINPUT78), .Z(n502) );
  XNOR2_X1 U607 ( .A(n502), .B(n501), .ZN(n503) );
  XNOR2_X1 U608 ( .A(n504), .B(n503), .ZN(n505) );
  XNOR2_X1 U609 ( .A(n506), .B(n505), .ZN(n717) );
  XOR2_X1 U610 ( .A(KEYINPUT96), .B(KEYINPUT25), .Z(n509) );
  XNOR2_X1 U611 ( .A(n509), .B(n363), .ZN(n510) );
  NAND2_X1 U612 ( .A1(n511), .A2(G210), .ZN(n513) );
  XNOR2_X1 U613 ( .A(n513), .B(n512), .ZN(n515) );
  XNOR2_X1 U614 ( .A(n515), .B(n514), .ZN(n519) );
  XNOR2_X1 U615 ( .A(KEYINPUT77), .B(KEYINPUT5), .ZN(n517) );
  XNOR2_X1 U616 ( .A(n516), .B(n517), .ZN(n518) );
  XNOR2_X1 U617 ( .A(n519), .B(n518), .ZN(n520) );
  XNOR2_X1 U618 ( .A(n521), .B(n520), .ZN(n712) );
  OR2_X1 U619 ( .A1(n712), .A2(G902), .ZN(n524) );
  INV_X1 U620 ( .A(KEYINPUT97), .ZN(n522) );
  XNOR2_X1 U621 ( .A(n522), .B(G472), .ZN(n523) );
  XNOR2_X1 U622 ( .A(n524), .B(n523), .ZN(n575) );
  INV_X1 U623 ( .A(n589), .ZN(n525) );
  NAND2_X1 U624 ( .A1(n666), .A2(n525), .ZN(n526) );
  XNOR2_X2 U625 ( .A(n527), .B(KEYINPUT106), .ZN(n729) );
  AND2_X1 U626 ( .A1(n661), .A2(n666), .ZN(n530) );
  XNOR2_X1 U627 ( .A(KEYINPUT105), .B(KEYINPUT6), .ZN(n528) );
  INV_X1 U628 ( .A(n599), .ZN(n529) );
  NAND2_X1 U629 ( .A1(n530), .A2(n529), .ZN(n531) );
  INV_X1 U630 ( .A(KEYINPUT79), .ZN(n532) );
  XNOR2_X1 U631 ( .A(n532), .B(KEYINPUT32), .ZN(n533) );
  XNOR2_X2 U632 ( .A(n534), .B(n533), .ZN(n727) );
  NAND2_X1 U633 ( .A1(n729), .A2(n727), .ZN(n567) );
  NAND2_X1 U634 ( .A1(n567), .A2(KEYINPUT64), .ZN(n545) );
  NAND2_X1 U635 ( .A1(n433), .A2(n599), .ZN(n538) );
  INV_X1 U636 ( .A(KEYINPUT107), .ZN(n536) );
  XNOR2_X1 U637 ( .A(n536), .B(KEYINPUT33), .ZN(n537) );
  NAND2_X1 U638 ( .A1(n688), .A2(n551), .ZN(n540) );
  INV_X1 U639 ( .A(KEYINPUT34), .ZN(n539) );
  XNOR2_X1 U640 ( .A(n540), .B(n539), .ZN(n542) );
  NOR2_X1 U641 ( .A1(n619), .A2(n620), .ZN(n541) );
  NAND2_X1 U642 ( .A1(n542), .A2(n541), .ZN(n544) );
  INV_X1 U643 ( .A(KEYINPUT35), .ZN(n543) );
  NAND2_X1 U644 ( .A1(n545), .A2(n728), .ZN(n546) );
  NAND2_X1 U645 ( .A1(n546), .A2(KEYINPUT44), .ZN(n564) );
  INV_X1 U646 ( .A(KEYINPUT64), .ZN(n547) );
  AND2_X1 U647 ( .A1(n727), .A2(n547), .ZN(n548) );
  NAND2_X1 U648 ( .A1(n729), .A2(n548), .ZN(n562) );
  NAND2_X1 U649 ( .A1(n662), .A2(n589), .ZN(n550) );
  INV_X1 U650 ( .A(n661), .ZN(n549) );
  NOR2_X1 U651 ( .A1(n550), .A2(n549), .ZN(n673) );
  NAND2_X1 U652 ( .A1(n662), .A2(n592), .ZN(n574) );
  NOR2_X1 U653 ( .A1(n574), .A2(n589), .ZN(n553) );
  NAND2_X1 U654 ( .A1(n551), .A2(n553), .ZN(n555) );
  INV_X1 U655 ( .A(KEYINPUT98), .ZN(n554) );
  INV_X1 U656 ( .A(n620), .ZN(n556) );
  OR2_X1 U657 ( .A1(n661), .A2(n666), .ZN(n557) );
  INV_X1 U658 ( .A(n742), .ZN(n559) );
  OR2_X1 U659 ( .A1(KEYINPUT64), .A2(KEYINPUT44), .ZN(n558) );
  NAND2_X1 U660 ( .A1(n564), .A2(n563), .ZN(n566) );
  INV_X1 U661 ( .A(KEYINPUT87), .ZN(n565) );
  XNOR2_X1 U662 ( .A(n566), .B(n565), .ZN(n571) );
  INV_X1 U663 ( .A(n728), .ZN(n568) );
  OR2_X1 U664 ( .A1(n568), .A2(KEYINPUT44), .ZN(n569) );
  NOR2_X2 U665 ( .A1(n571), .A2(n570), .ZN(n573) );
  INV_X1 U666 ( .A(KEYINPUT45), .ZN(n572) );
  XNOR2_X1 U667 ( .A(n573), .B(n572), .ZN(n703) );
  NOR2_X1 U668 ( .A1(n770), .A2(KEYINPUT83), .ZN(n644) );
  INV_X1 U669 ( .A(n574), .ZN(n582) );
  NAND2_X1 U670 ( .A1(n575), .A2(n445), .ZN(n576) );
  XNOR2_X1 U671 ( .A(n576), .B(KEYINPUT30), .ZN(n581) );
  NAND2_X1 U672 ( .A1(G953), .A2(n577), .ZN(n578) );
  OR2_X1 U673 ( .A1(n578), .A2(G900), .ZN(n580) );
  AND2_X1 U674 ( .A1(n580), .A2(n579), .ZN(n587) );
  BUF_X2 U675 ( .A(n583), .Z(n633) );
  INV_X1 U676 ( .A(KEYINPUT38), .ZN(n584) );
  INV_X1 U677 ( .A(n597), .ZN(n585) );
  INV_X1 U678 ( .A(KEYINPUT40), .ZN(n586) );
  NOR2_X1 U679 ( .A1(n587), .A2(n665), .ZN(n588) );
  AND2_X1 U680 ( .A1(n666), .A2(n432), .ZN(n598) );
  NAND2_X1 U681 ( .A1(n598), .A2(n589), .ZN(n591) );
  INV_X1 U682 ( .A(KEYINPUT28), .ZN(n590) );
  XNOR2_X1 U683 ( .A(n591), .B(n590), .ZN(n593) );
  AND2_X1 U684 ( .A1(n593), .A2(n592), .ZN(n609) );
  NAND2_X1 U685 ( .A1(n677), .A2(n609), .ZN(n595) );
  XNOR2_X1 U686 ( .A(KEYINPUT109), .B(KEYINPUT42), .ZN(n594) );
  XNOR2_X1 U687 ( .A(n595), .B(n594), .ZN(n796) );
  INV_X1 U688 ( .A(n601), .ZN(n602) );
  INV_X1 U689 ( .A(KEYINPUT36), .ZN(n603) );
  XNOR2_X1 U690 ( .A(n604), .B(n603), .ZN(n605) );
  NAND2_X1 U691 ( .A1(n605), .A2(n661), .ZN(n725) );
  NAND2_X1 U692 ( .A1(n606), .A2(KEYINPUT82), .ZN(n611) );
  INV_X1 U693 ( .A(n607), .ZN(n608) );
  NAND2_X1 U694 ( .A1(n609), .A2(n608), .ZN(n612) );
  INV_X1 U695 ( .A(KEYINPUT47), .ZN(n613) );
  NOR2_X1 U696 ( .A1(n612), .A2(n613), .ZN(n610) );
  NAND2_X1 U697 ( .A1(n611), .A2(n610), .ZN(n617) );
  INV_X1 U698 ( .A(n612), .ZN(n751) );
  NAND2_X1 U699 ( .A1(n684), .A2(n751), .ZN(n615) );
  AND2_X1 U700 ( .A1(n613), .A2(KEYINPUT82), .ZN(n614) );
  NAND2_X1 U701 ( .A1(n615), .A2(n614), .ZN(n616) );
  NAND2_X1 U702 ( .A1(n617), .A2(n616), .ZN(n628) );
  INV_X1 U703 ( .A(KEYINPUT82), .ZN(n618) );
  NAND2_X1 U704 ( .A1(n684), .A2(n618), .ZN(n626) );
  INV_X1 U705 ( .A(n619), .ZN(n622) );
  NOR2_X1 U706 ( .A1(n633), .A2(n620), .ZN(n621) );
  NAND2_X1 U707 ( .A1(n622), .A2(n621), .ZN(n624) );
  NOR2_X1 U708 ( .A1(n624), .A2(n623), .ZN(n750) );
  INV_X1 U709 ( .A(n750), .ZN(n625) );
  AND2_X1 U710 ( .A1(n626), .A2(n625), .ZN(n627) );
  AND2_X1 U711 ( .A1(n628), .A2(n627), .ZN(n629) );
  INV_X1 U712 ( .A(KEYINPUT48), .ZN(n630) );
  NOR2_X1 U713 ( .A1(n661), .A2(n680), .ZN(n631) );
  NAND2_X1 U714 ( .A1(n365), .A2(n631), .ZN(n632) );
  XNOR2_X1 U715 ( .A(n632), .B(KEYINPUT43), .ZN(n634) );
  NAND2_X1 U716 ( .A1(n634), .A2(n633), .ZN(n722) );
  INV_X1 U717 ( .A(n755), .ZN(n635) );
  OR2_X1 U718 ( .A1(n636), .A2(n635), .ZN(n638) );
  INV_X1 U719 ( .A(KEYINPUT111), .ZN(n637) );
  XNOR2_X1 U720 ( .A(n638), .B(n637), .ZN(n795) );
  AND2_X1 U721 ( .A1(n722), .A2(n795), .ZN(n639) );
  INV_X1 U722 ( .A(KEYINPUT86), .ZN(n640) );
  INV_X1 U723 ( .A(KEYINPUT84), .ZN(n651) );
  XOR2_X1 U724 ( .A(KEYINPUT2), .B(KEYINPUT81), .Z(n646) );
  INV_X1 U725 ( .A(n646), .ZN(n641) );
  NAND2_X1 U726 ( .A1(n642), .A2(n641), .ZN(n643) );
  OR2_X1 U727 ( .A1(n644), .A2(n643), .ZN(n648) );
  NOR2_X1 U728 ( .A1(n651), .A2(KEYINPUT83), .ZN(n645) );
  NAND2_X1 U729 ( .A1(n646), .A2(n645), .ZN(n647) );
  NAND2_X1 U730 ( .A1(n648), .A2(n647), .ZN(n657) );
  INV_X1 U731 ( .A(KEYINPUT2), .ZN(n706) );
  NOR2_X1 U732 ( .A1(n649), .A2(n706), .ZN(n650) );
  NAND2_X1 U733 ( .A1(n770), .A2(n650), .ZN(n710) );
  INV_X1 U734 ( .A(n710), .ZN(n655) );
  NAND2_X1 U735 ( .A1(n770), .A2(KEYINPUT83), .ZN(n653) );
  NAND2_X1 U736 ( .A1(n787), .A2(n651), .ZN(n652) );
  NAND2_X1 U737 ( .A1(n653), .A2(n652), .ZN(n654) );
  NOR2_X1 U738 ( .A1(n655), .A2(n654), .ZN(n656) );
  NAND2_X1 U739 ( .A1(n657), .A2(n656), .ZN(n660) );
  NAND2_X1 U740 ( .A1(n677), .A2(n688), .ZN(n658) );
  XNOR2_X1 U741 ( .A(n658), .B(KEYINPUT120), .ZN(n659) );
  NAND2_X1 U742 ( .A1(n660), .A2(n659), .ZN(n697) );
  XOR2_X1 U743 ( .A(KEYINPUT50), .B(KEYINPUT116), .Z(n664) );
  NOR2_X1 U744 ( .A1(n662), .A2(n661), .ZN(n663) );
  XOR2_X1 U745 ( .A(n664), .B(n663), .Z(n672) );
  NAND2_X1 U746 ( .A1(n666), .A2(n665), .ZN(n667) );
  XNOR2_X1 U747 ( .A(n667), .B(KEYINPUT114), .ZN(n668) );
  XNOR2_X1 U748 ( .A(n668), .B(KEYINPUT49), .ZN(n669) );
  NOR2_X1 U749 ( .A1(n669), .A2(n589), .ZN(n670) );
  XNOR2_X1 U750 ( .A(n670), .B(KEYINPUT115), .ZN(n671) );
  NOR2_X1 U751 ( .A1(n672), .A2(n671), .ZN(n674) );
  NOR2_X1 U752 ( .A1(n674), .A2(n673), .ZN(n676) );
  XOR2_X1 U753 ( .A(KEYINPUT117), .B(KEYINPUT51), .Z(n675) );
  XNOR2_X1 U754 ( .A(n676), .B(n675), .ZN(n678) );
  NAND2_X1 U755 ( .A1(n678), .A2(n677), .ZN(n679) );
  XNOR2_X1 U756 ( .A(n679), .B(KEYINPUT118), .ZN(n691) );
  NAND2_X1 U757 ( .A1(n681), .A2(n680), .ZN(n683) );
  NAND2_X1 U758 ( .A1(n683), .A2(n682), .ZN(n687) );
  NAND2_X1 U759 ( .A1(n685), .A2(n684), .ZN(n686) );
  NAND2_X1 U760 ( .A1(n687), .A2(n686), .ZN(n689) );
  NAND2_X1 U761 ( .A1(n689), .A2(n688), .ZN(n690) );
  NAND2_X1 U762 ( .A1(n691), .A2(n690), .ZN(n692) );
  XOR2_X1 U763 ( .A(KEYINPUT52), .B(n692), .Z(n693) );
  NOR2_X1 U764 ( .A1(n694), .A2(n693), .ZN(n695) );
  XOR2_X1 U765 ( .A(KEYINPUT119), .B(n695), .Z(n696) );
  NAND2_X1 U766 ( .A1(n788), .A2(n698), .ZN(n699) );
  INV_X1 U767 ( .A(n707), .ZN(n700) );
  NAND2_X1 U768 ( .A1(n703), .A2(n702), .ZN(n705) );
  XNOR2_X1 U769 ( .A(n705), .B(n704), .ZN(n709) );
  OR2_X1 U770 ( .A1(n707), .A2(n706), .ZN(n708) );
  NAND2_X1 U771 ( .A1(n758), .A2(G472), .ZN(n713) );
  INV_X1 U772 ( .A(G952), .ZN(n714) );
  AND2_X1 U773 ( .A1(n714), .A2(G953), .ZN(n769) );
  XNOR2_X1 U774 ( .A(n719), .B(KEYINPUT123), .ZN(G66) );
  XNOR2_X1 U775 ( .A(G131), .B(KEYINPUT127), .ZN(n720) );
  XNOR2_X1 U776 ( .A(n721), .B(n720), .ZN(G33) );
  XNOR2_X1 U777 ( .A(n722), .B(G140), .ZN(G42) );
  XOR2_X1 U778 ( .A(KEYINPUT112), .B(KEYINPUT113), .Z(n724) );
  XNOR2_X1 U779 ( .A(G125), .B(KEYINPUT37), .ZN(n723) );
  XNOR2_X1 U780 ( .A(n724), .B(n723), .ZN(n726) );
  XOR2_X1 U781 ( .A(n726), .B(n725), .Z(G27) );
  XNOR2_X1 U782 ( .A(n727), .B(G119), .ZN(G21) );
  XNOR2_X1 U783 ( .A(n728), .B(G122), .ZN(G24) );
  XNOR2_X1 U784 ( .A(n729), .B(G110), .ZN(G12) );
  NAND2_X1 U785 ( .A1(n758), .A2(G475), .ZN(n732) );
  XNOR2_X1 U786 ( .A(n730), .B(KEYINPUT59), .ZN(n731) );
  XNOR2_X1 U787 ( .A(n732), .B(n731), .ZN(n733) );
  XNOR2_X1 U788 ( .A(KEYINPUT122), .B(KEYINPUT60), .ZN(n734) );
  XNOR2_X1 U789 ( .A(n735), .B(n734), .ZN(G60) );
  NAND2_X1 U790 ( .A1(n758), .A2(G210), .ZN(n739) );
  XNOR2_X1 U791 ( .A(KEYINPUT54), .B(KEYINPUT55), .ZN(n737) );
  XNOR2_X1 U792 ( .A(n736), .B(n737), .ZN(n738) );
  XNOR2_X1 U793 ( .A(n739), .B(n738), .ZN(n740) );
  XNOR2_X1 U794 ( .A(n741), .B(KEYINPUT56), .ZN(G51) );
  XOR2_X1 U795 ( .A(G101), .B(n742), .Z(G3) );
  NAND2_X1 U796 ( .A1(n744), .A2(n753), .ZN(n743) );
  XNOR2_X1 U797 ( .A(n743), .B(G104), .ZN(G6) );
  XOR2_X1 U798 ( .A(KEYINPUT27), .B(KEYINPUT26), .Z(n746) );
  NAND2_X1 U799 ( .A1(n755), .A2(n744), .ZN(n745) );
  XNOR2_X1 U800 ( .A(n746), .B(n745), .ZN(n747) );
  XNOR2_X1 U801 ( .A(G107), .B(n747), .ZN(G9) );
  XOR2_X1 U802 ( .A(G128), .B(KEYINPUT29), .Z(n749) );
  NAND2_X1 U803 ( .A1(n751), .A2(n755), .ZN(n748) );
  XNOR2_X1 U804 ( .A(n749), .B(n748), .ZN(G30) );
  XOR2_X1 U805 ( .A(G143), .B(n750), .Z(G45) );
  NAND2_X1 U806 ( .A1(n753), .A2(n751), .ZN(n752) );
  XNOR2_X1 U807 ( .A(n752), .B(G146), .ZN(G48) );
  NAND2_X1 U808 ( .A1(n753), .A2(n756), .ZN(n754) );
  XNOR2_X1 U809 ( .A(n754), .B(G113), .ZN(G15) );
  NAND2_X1 U810 ( .A1(n756), .A2(n755), .ZN(n757) );
  XNOR2_X1 U811 ( .A(n757), .B(G116), .ZN(G18) );
  NAND2_X1 U812 ( .A1(n765), .A2(G469), .ZN(n763) );
  XNOR2_X1 U813 ( .A(KEYINPUT58), .B(KEYINPUT121), .ZN(n759) );
  XOR2_X1 U814 ( .A(n759), .B(KEYINPUT57), .Z(n760) );
  XNOR2_X1 U815 ( .A(n761), .B(n760), .ZN(n762) );
  XNOR2_X1 U816 ( .A(n763), .B(n762), .ZN(n764) );
  NOR2_X1 U817 ( .A1(n769), .A2(n764), .ZN(G54) );
  NAND2_X1 U818 ( .A1(n765), .A2(G478), .ZN(n767) );
  XNOR2_X1 U819 ( .A(n767), .B(n766), .ZN(n768) );
  NOR2_X1 U820 ( .A1(n769), .A2(n768), .ZN(G63) );
  NAND2_X1 U821 ( .A1(n770), .A2(n788), .ZN(n775) );
  NAND2_X1 U822 ( .A1(G224), .A2(G953), .ZN(n771) );
  XNOR2_X1 U823 ( .A(n771), .B(KEYINPUT124), .ZN(n772) );
  XNOR2_X1 U824 ( .A(KEYINPUT61), .B(n772), .ZN(n773) );
  NAND2_X1 U825 ( .A1(n773), .A2(G898), .ZN(n774) );
  NAND2_X1 U826 ( .A1(n775), .A2(n774), .ZN(n783) );
  XNOR2_X1 U827 ( .A(G101), .B(n776), .ZN(n777) );
  XNOR2_X1 U828 ( .A(n777), .B(KEYINPUT125), .ZN(n779) );
  XNOR2_X1 U829 ( .A(n779), .B(n778), .ZN(n780) );
  NOR2_X1 U830 ( .A1(n781), .A2(n780), .ZN(n782) );
  XNOR2_X1 U831 ( .A(n783), .B(n782), .ZN(G69) );
  XNOR2_X1 U832 ( .A(n784), .B(KEYINPUT126), .ZN(n786) );
  XNOR2_X1 U833 ( .A(n786), .B(n785), .ZN(n790) );
  XOR2_X1 U834 ( .A(n790), .B(n787), .Z(n789) );
  NAND2_X1 U835 ( .A1(n789), .A2(n788), .ZN(n794) );
  XNOR2_X1 U836 ( .A(G227), .B(n790), .ZN(n791) );
  NAND2_X1 U837 ( .A1(n791), .A2(G900), .ZN(n792) );
  NAND2_X1 U838 ( .A1(n792), .A2(G953), .ZN(n793) );
  NAND2_X1 U839 ( .A1(n794), .A2(n793), .ZN(G72) );
  XNOR2_X1 U840 ( .A(G134), .B(n795), .ZN(G36) );
  XOR2_X1 U841 ( .A(G137), .B(n796), .Z(G39) );
endmodule

