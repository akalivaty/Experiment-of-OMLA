//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 1 1 1 1 1 1 1 1 1 0 1 0 0 1 1 0 0 1 1 1 0 1 0 1 0 1 0 0 1 1 1 0 1 1 0 1 0 0 0 1 0 1 1 1 1 0 1 0 0 1 1 0 0 0 0 0 0 0 0 1 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:42:23 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n205, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n236, new_n237,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n244, new_n245,
    new_n246, new_n248, new_n249, new_n250, new_n251, new_n252, new_n253,
    new_n254, new_n255, new_n256, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1108, new_n1109, new_n1110, new_n1111, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1186, new_n1187, new_n1188, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1251, new_n1252,
    new_n1253, new_n1254, new_n1255, new_n1256, new_n1257, new_n1258,
    new_n1259, new_n1260, new_n1261, new_n1262, new_n1263, new_n1264,
    new_n1265, new_n1266, new_n1268, new_n1269, new_n1270, new_n1271,
    new_n1272, new_n1273, new_n1274, new_n1275, new_n1276, new_n1277,
    new_n1278, new_n1279, new_n1280, new_n1281, new_n1282, new_n1283,
    new_n1284, new_n1285, new_n1286, new_n1287, new_n1288, new_n1289,
    new_n1290, new_n1291, new_n1292, new_n1293, new_n1295, new_n1296,
    new_n1297, new_n1298, new_n1299, new_n1300, new_n1301, new_n1303,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1346,
    new_n1347, new_n1348, new_n1349, new_n1350, new_n1351, new_n1352,
    new_n1353, new_n1354, new_n1355, new_n1357, new_n1358, new_n1359,
    new_n1360, new_n1361, new_n1362, new_n1363, new_n1364;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND3_X1  g0002(.A1(new_n201), .A2(KEYINPUT64), .A3(new_n202), .ZN(new_n203));
  INV_X1    g0003(.A(new_n203), .ZN(new_n204));
  AOI21_X1  g0004(.A(KEYINPUT64), .B1(new_n201), .B2(new_n202), .ZN(new_n205));
  NOR3_X1   g0005(.A1(new_n204), .A2(new_n205), .A3(G77), .ZN(G353));
  OAI21_X1  g0006(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0007(.A(G1), .ZN(new_n208));
  INV_X1    g0008(.A(G20), .ZN(new_n209));
  NOR2_X1   g0009(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  INV_X1    g0010(.A(new_n210), .ZN(new_n211));
  NOR2_X1   g0011(.A1(new_n211), .A2(G13), .ZN(new_n212));
  OAI211_X1 g0012(.A(new_n212), .B(G250), .C1(G257), .C2(G264), .ZN(new_n213));
  XOR2_X1   g0013(.A(new_n213), .B(KEYINPUT0), .Z(new_n214));
  AND2_X1   g0014(.A1(G107), .A2(G264), .ZN(new_n215));
  INV_X1    g0015(.A(G87), .ZN(new_n216));
  INV_X1    g0016(.A(G250), .ZN(new_n217));
  INV_X1    g0017(.A(G97), .ZN(new_n218));
  INV_X1    g0018(.A(G257), .ZN(new_n219));
  OAI22_X1  g0019(.A1(new_n216), .A2(new_n217), .B1(new_n218), .B2(new_n219), .ZN(new_n220));
  AOI211_X1 g0020(.A(new_n215), .B(new_n220), .C1(G68), .C2(G238), .ZN(new_n221));
  NAND2_X1  g0021(.A1(G116), .A2(G270), .ZN(new_n222));
  AND2_X1   g0022(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  INV_X1    g0023(.A(G226), .ZN(new_n224));
  INV_X1    g0024(.A(G77), .ZN(new_n225));
  INV_X1    g0025(.A(G244), .ZN(new_n226));
  OAI221_X1 g0026(.A(new_n223), .B1(new_n202), .B2(new_n224), .C1(new_n225), .C2(new_n226), .ZN(new_n227));
  INV_X1    g0027(.A(G58), .ZN(new_n228));
  INV_X1    g0028(.A(G232), .ZN(new_n229));
  NOR2_X1   g0029(.A1(new_n228), .A2(new_n229), .ZN(new_n230));
  OAI21_X1  g0030(.A(new_n211), .B1(new_n227), .B2(new_n230), .ZN(new_n231));
  XNOR2_X1  g0031(.A(new_n231), .B(KEYINPUT1), .ZN(new_n232));
  NAND2_X1  g0032(.A1(G1), .A2(G13), .ZN(new_n233));
  NOR2_X1   g0033(.A1(new_n233), .A2(new_n209), .ZN(new_n234));
  XOR2_X1   g0034(.A(new_n234), .B(KEYINPUT65), .Z(new_n235));
  OAI21_X1  g0035(.A(G50), .B1(G58), .B2(G68), .ZN(new_n236));
  INV_X1    g0036(.A(new_n236), .ZN(new_n237));
  AOI211_X1 g0037(.A(new_n214), .B(new_n232), .C1(new_n235), .C2(new_n237), .ZN(G361));
  XNOR2_X1  g0038(.A(G250), .B(G257), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n239), .B(G264), .ZN(new_n240));
  XOR2_X1   g0040(.A(new_n240), .B(G270), .Z(new_n241));
  XNOR2_X1  g0041(.A(G238), .B(G244), .ZN(new_n242));
  XNOR2_X1  g0042(.A(KEYINPUT66), .B(KEYINPUT2), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XOR2_X1   g0044(.A(G226), .B(G232), .Z(new_n245));
  XNOR2_X1  g0045(.A(new_n244), .B(new_n245), .ZN(new_n246));
  XOR2_X1   g0046(.A(new_n241), .B(new_n246), .Z(G358));
  XNOR2_X1  g0047(.A(G87), .B(G97), .ZN(new_n248));
  INV_X1    g0048(.A(G107), .ZN(new_n249));
  XNOR2_X1  g0049(.A(new_n248), .B(new_n249), .ZN(new_n250));
  INV_X1    g0050(.A(G116), .ZN(new_n251));
  XNOR2_X1  g0051(.A(new_n250), .B(new_n251), .ZN(new_n252));
  XNOR2_X1  g0052(.A(new_n252), .B(KEYINPUT67), .ZN(new_n253));
  XNOR2_X1  g0053(.A(G68), .B(G77), .ZN(new_n254));
  XNOR2_X1  g0054(.A(new_n254), .B(new_n202), .ZN(new_n255));
  XNOR2_X1  g0055(.A(new_n255), .B(new_n228), .ZN(new_n256));
  XNOR2_X1  g0056(.A(new_n253), .B(new_n256), .ZN(G351));
  INV_X1    g0057(.A(KEYINPUT70), .ZN(new_n258));
  NAND3_X1  g0058(.A1(new_n208), .A2(G13), .A3(G20), .ZN(new_n259));
  INV_X1    g0059(.A(new_n259), .ZN(new_n260));
  NAND3_X1  g0060(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n261), .A2(new_n233), .ZN(new_n262));
  OAI21_X1  g0062(.A(new_n258), .B1(new_n260), .B2(new_n262), .ZN(new_n263));
  NAND4_X1  g0063(.A1(new_n259), .A2(KEYINPUT70), .A3(new_n233), .A4(new_n261), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n263), .A2(new_n264), .ZN(new_n265));
  AND3_X1   g0065(.A1(new_n208), .A2(KEYINPUT77), .A3(G33), .ZN(new_n266));
  AOI21_X1  g0066(.A(KEYINPUT77), .B1(new_n208), .B2(G33), .ZN(new_n267));
  NOR2_X1   g0067(.A1(new_n266), .A2(new_n267), .ZN(new_n268));
  INV_X1    g0068(.A(new_n268), .ZN(new_n269));
  NAND3_X1  g0069(.A1(new_n265), .A2(G116), .A3(new_n269), .ZN(new_n270));
  INV_X1    g0070(.A(G13), .ZN(new_n271));
  NOR2_X1   g0071(.A1(new_n271), .A2(G1), .ZN(new_n272));
  NAND3_X1  g0072(.A1(new_n272), .A2(G20), .A3(new_n251), .ZN(new_n273));
  NAND2_X1  g0073(.A1(G33), .A2(G283), .ZN(new_n274));
  OAI211_X1 g0074(.A(new_n274), .B(new_n209), .C1(G33), .C2(new_n218), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n251), .A2(G20), .ZN(new_n276));
  NAND3_X1  g0076(.A1(new_n275), .A2(new_n276), .A3(new_n262), .ZN(new_n277));
  INV_X1    g0077(.A(KEYINPUT20), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n277), .A2(new_n278), .ZN(new_n279));
  NAND4_X1  g0079(.A1(new_n275), .A2(KEYINPUT20), .A3(new_n262), .A4(new_n276), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n279), .A2(new_n280), .ZN(new_n281));
  AND3_X1   g0081(.A1(new_n270), .A2(new_n273), .A3(new_n281), .ZN(new_n282));
  INV_X1    g0082(.A(G1698), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n283), .A2(G257), .ZN(new_n284));
  NAND2_X1  g0084(.A1(G264), .A2(G1698), .ZN(new_n285));
  AND2_X1   g0085(.A1(KEYINPUT3), .A2(G33), .ZN(new_n286));
  NOR2_X1   g0086(.A1(KEYINPUT3), .A2(G33), .ZN(new_n287));
  OAI211_X1 g0087(.A(new_n284), .B(new_n285), .C1(new_n286), .C2(new_n287), .ZN(new_n288));
  AOI21_X1  g0088(.A(new_n233), .B1(G33), .B2(G41), .ZN(new_n289));
  INV_X1    g0089(.A(KEYINPUT3), .ZN(new_n290));
  INV_X1    g0090(.A(G33), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n290), .A2(new_n291), .ZN(new_n292));
  INV_X1    g0092(.A(G303), .ZN(new_n293));
  NAND2_X1  g0093(.A1(KEYINPUT3), .A2(G33), .ZN(new_n294));
  NAND3_X1  g0094(.A1(new_n292), .A2(new_n293), .A3(new_n294), .ZN(new_n295));
  NAND3_X1  g0095(.A1(new_n288), .A2(new_n289), .A3(new_n295), .ZN(new_n296));
  INV_X1    g0096(.A(G45), .ZN(new_n297));
  NOR2_X1   g0097(.A1(new_n297), .A2(G1), .ZN(new_n298));
  NAND2_X1  g0098(.A1(KEYINPUT5), .A2(G41), .ZN(new_n299));
  INV_X1    g0099(.A(new_n299), .ZN(new_n300));
  NOR2_X1   g0100(.A1(KEYINPUT5), .A2(G41), .ZN(new_n301));
  OAI21_X1  g0101(.A(new_n298), .B1(new_n300), .B2(new_n301), .ZN(new_n302));
  INV_X1    g0102(.A(G41), .ZN(new_n303));
  OAI211_X1 g0103(.A(G1), .B(G13), .C1(new_n291), .C2(new_n303), .ZN(new_n304));
  NAND3_X1  g0104(.A1(new_n302), .A2(G270), .A3(new_n304), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n208), .A2(G45), .ZN(new_n306));
  OR2_X1    g0106(.A1(KEYINPUT5), .A2(G41), .ZN(new_n307));
  AOI21_X1  g0107(.A(new_n306), .B1(new_n307), .B2(new_n299), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n308), .A2(G274), .ZN(new_n309));
  NAND3_X1  g0109(.A1(new_n296), .A2(new_n305), .A3(new_n309), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n310), .A2(G200), .ZN(new_n311));
  NAND4_X1  g0111(.A1(new_n296), .A2(new_n305), .A3(new_n309), .A4(G190), .ZN(new_n312));
  NAND4_X1  g0112(.A1(new_n282), .A2(KEYINPUT81), .A3(new_n311), .A4(new_n312), .ZN(new_n313));
  INV_X1    g0113(.A(KEYINPUT81), .ZN(new_n314));
  NAND4_X1  g0114(.A1(new_n270), .A2(new_n312), .A3(new_n273), .A4(new_n281), .ZN(new_n315));
  INV_X1    g0115(.A(new_n311), .ZN(new_n316));
  OAI21_X1  g0116(.A(new_n314), .B1(new_n315), .B2(new_n316), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n313), .A2(new_n317), .ZN(new_n318));
  NAND3_X1  g0118(.A1(new_n270), .A2(new_n273), .A3(new_n281), .ZN(new_n319));
  INV_X1    g0119(.A(G179), .ZN(new_n320));
  NOR2_X1   g0120(.A1(new_n310), .A2(new_n320), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n319), .A2(new_n321), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n310), .A2(G169), .ZN(new_n323));
  AOI21_X1  g0123(.A(new_n268), .B1(new_n263), .B2(new_n264), .ZN(new_n324));
  AOI22_X1  g0124(.A1(new_n324), .A2(G116), .B1(new_n279), .B2(new_n280), .ZN(new_n325));
  AOI21_X1  g0125(.A(new_n323), .B1(new_n325), .B2(new_n273), .ZN(new_n326));
  INV_X1    g0126(.A(KEYINPUT80), .ZN(new_n327));
  OAI21_X1  g0127(.A(KEYINPUT21), .B1(new_n326), .B2(new_n327), .ZN(new_n328));
  AND2_X1   g0128(.A1(new_n310), .A2(G169), .ZN(new_n329));
  AOI21_X1  g0129(.A(new_n327), .B1(new_n319), .B2(new_n329), .ZN(new_n330));
  INV_X1    g0130(.A(KEYINPUT21), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n330), .A2(new_n331), .ZN(new_n332));
  NAND4_X1  g0132(.A1(new_n318), .A2(new_n322), .A3(new_n328), .A4(new_n332), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n333), .A2(KEYINPUT82), .ZN(new_n334));
  NOR2_X1   g0134(.A1(new_n330), .A2(new_n331), .ZN(new_n335));
  AOI211_X1 g0135(.A(new_n327), .B(KEYINPUT21), .C1(new_n319), .C2(new_n329), .ZN(new_n336));
  NOR2_X1   g0136(.A1(new_n335), .A2(new_n336), .ZN(new_n337));
  INV_X1    g0137(.A(KEYINPUT82), .ZN(new_n338));
  NAND4_X1  g0138(.A1(new_n337), .A2(new_n338), .A3(new_n322), .A4(new_n318), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n334), .A2(new_n339), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n292), .A2(new_n294), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n283), .A2(G222), .ZN(new_n342));
  INV_X1    g0142(.A(G223), .ZN(new_n343));
  OAI211_X1 g0143(.A(new_n341), .B(new_n342), .C1(new_n343), .C2(new_n283), .ZN(new_n344));
  OAI211_X1 g0144(.A(new_n344), .B(new_n289), .C1(G77), .C2(new_n341), .ZN(new_n345));
  OAI21_X1  g0145(.A(new_n208), .B1(G41), .B2(G45), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n304), .A2(new_n346), .ZN(new_n347));
  INV_X1    g0147(.A(new_n347), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n348), .A2(G226), .ZN(new_n349));
  AOI21_X1  g0149(.A(G1), .B1(new_n303), .B2(new_n297), .ZN(new_n350));
  INV_X1    g0150(.A(KEYINPUT68), .ZN(new_n351));
  NAND3_X1  g0151(.A1(new_n350), .A2(new_n351), .A3(G274), .ZN(new_n352));
  INV_X1    g0152(.A(G274), .ZN(new_n353));
  OAI21_X1  g0153(.A(KEYINPUT68), .B1(new_n346), .B2(new_n353), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n352), .A2(new_n354), .ZN(new_n355));
  NAND3_X1  g0155(.A1(new_n345), .A2(new_n349), .A3(new_n355), .ZN(new_n356));
  INV_X1    g0156(.A(G169), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n356), .A2(new_n357), .ZN(new_n358));
  OAI21_X1  g0158(.A(new_n358), .B1(G179), .B2(new_n356), .ZN(new_n359));
  INV_X1    g0159(.A(new_n205), .ZN(new_n360));
  AOI21_X1  g0160(.A(new_n209), .B1(new_n360), .B2(new_n203), .ZN(new_n361));
  XNOR2_X1  g0161(.A(KEYINPUT8), .B(G58), .ZN(new_n362));
  NOR2_X1   g0162(.A1(new_n291), .A2(G20), .ZN(new_n363));
  INV_X1    g0163(.A(new_n363), .ZN(new_n364));
  INV_X1    g0164(.A(G150), .ZN(new_n365));
  NOR2_X1   g0165(.A1(G20), .A2(G33), .ZN(new_n366));
  INV_X1    g0166(.A(new_n366), .ZN(new_n367));
  OAI22_X1  g0167(.A1(new_n362), .A2(new_n364), .B1(new_n365), .B2(new_n367), .ZN(new_n368));
  OAI21_X1  g0168(.A(new_n262), .B1(new_n361), .B2(new_n368), .ZN(new_n369));
  NOR2_X1   g0169(.A1(new_n260), .A2(new_n262), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n208), .A2(G20), .ZN(new_n371));
  NAND3_X1  g0171(.A1(new_n370), .A2(G50), .A3(new_n371), .ZN(new_n372));
  OAI211_X1 g0172(.A(new_n369), .B(new_n372), .C1(G50), .C2(new_n259), .ZN(new_n373));
  INV_X1    g0173(.A(new_n373), .ZN(new_n374));
  NOR2_X1   g0174(.A1(new_n359), .A2(new_n374), .ZN(new_n375));
  INV_X1    g0175(.A(KEYINPUT71), .ZN(new_n376));
  NOR2_X1   g0176(.A1(new_n373), .A2(new_n376), .ZN(new_n377));
  INV_X1    g0177(.A(new_n362), .ZN(new_n378));
  AOI22_X1  g0178(.A1(new_n378), .A2(new_n363), .B1(G150), .B2(new_n366), .ZN(new_n379));
  OAI21_X1  g0179(.A(G20), .B1(new_n204), .B2(new_n205), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n379), .A2(new_n380), .ZN(new_n381));
  AOI22_X1  g0181(.A1(new_n381), .A2(new_n262), .B1(new_n202), .B2(new_n260), .ZN(new_n382));
  AOI21_X1  g0182(.A(KEYINPUT71), .B1(new_n382), .B2(new_n372), .ZN(new_n383));
  OAI21_X1  g0183(.A(KEYINPUT9), .B1(new_n377), .B2(new_n383), .ZN(new_n384));
  NAND2_X1  g0184(.A1(new_n373), .A2(new_n376), .ZN(new_n385));
  NAND3_X1  g0185(.A1(new_n382), .A2(KEYINPUT71), .A3(new_n372), .ZN(new_n386));
  INV_X1    g0186(.A(KEYINPUT9), .ZN(new_n387));
  NAND3_X1  g0187(.A1(new_n385), .A2(new_n386), .A3(new_n387), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n356), .A2(G200), .ZN(new_n389));
  INV_X1    g0189(.A(new_n356), .ZN(new_n390));
  NAND2_X1  g0190(.A1(new_n390), .A2(G190), .ZN(new_n391));
  NAND4_X1  g0191(.A1(new_n384), .A2(new_n388), .A3(new_n389), .A4(new_n391), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n392), .A2(KEYINPUT10), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n385), .A2(new_n386), .ZN(new_n394));
  AOI22_X1  g0194(.A1(new_n394), .A2(KEYINPUT9), .B1(G190), .B2(new_n390), .ZN(new_n395));
  INV_X1    g0195(.A(KEYINPUT10), .ZN(new_n396));
  NAND4_X1  g0196(.A1(new_n395), .A2(new_n396), .A3(new_n388), .A4(new_n389), .ZN(new_n397));
  AOI21_X1  g0197(.A(new_n375), .B1(new_n393), .B2(new_n397), .ZN(new_n398));
  AOI22_X1  g0198(.A1(new_n348), .A2(G232), .B1(new_n352), .B2(new_n354), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n343), .A2(new_n283), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n224), .A2(G1698), .ZN(new_n401));
  OAI211_X1 g0201(.A(new_n400), .B(new_n401), .C1(new_n286), .C2(new_n287), .ZN(new_n402));
  NAND2_X1  g0202(.A1(G33), .A2(G87), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n402), .A2(new_n403), .ZN(new_n404));
  AOI21_X1  g0204(.A(KEYINPUT75), .B1(new_n404), .B2(new_n289), .ZN(new_n405));
  INV_X1    g0205(.A(KEYINPUT75), .ZN(new_n406));
  AOI211_X1 g0206(.A(new_n406), .B(new_n304), .C1(new_n402), .C2(new_n403), .ZN(new_n407));
  OAI211_X1 g0207(.A(new_n320), .B(new_n399), .C1(new_n405), .C2(new_n407), .ZN(new_n408));
  OAI21_X1  g0208(.A(new_n355), .B1(new_n229), .B2(new_n347), .ZN(new_n409));
  AOI21_X1  g0209(.A(new_n304), .B1(new_n402), .B2(new_n403), .ZN(new_n410));
  OAI21_X1  g0210(.A(new_n357), .B1(new_n409), .B2(new_n410), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n408), .A2(new_n411), .ZN(new_n412));
  INV_X1    g0212(.A(new_n412), .ZN(new_n413));
  INV_X1    g0213(.A(KEYINPUT16), .ZN(new_n414));
  INV_X1    g0214(.A(G68), .ZN(new_n415));
  NAND3_X1  g0215(.A1(new_n292), .A2(new_n209), .A3(new_n294), .ZN(new_n416));
  INV_X1    g0216(.A(KEYINPUT7), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n416), .A2(new_n417), .ZN(new_n418));
  NOR2_X1   g0218(.A1(new_n286), .A2(new_n287), .ZN(new_n419));
  NAND3_X1  g0219(.A1(new_n419), .A2(KEYINPUT7), .A3(new_n209), .ZN(new_n420));
  AOI21_X1  g0220(.A(new_n415), .B1(new_n418), .B2(new_n420), .ZN(new_n421));
  NOR2_X1   g0221(.A1(new_n228), .A2(new_n415), .ZN(new_n422));
  OAI21_X1  g0222(.A(G20), .B1(new_n422), .B2(new_n201), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n366), .A2(G159), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n423), .A2(new_n424), .ZN(new_n425));
  OAI21_X1  g0225(.A(new_n414), .B1(new_n421), .B2(new_n425), .ZN(new_n426));
  AOI21_X1  g0226(.A(KEYINPUT7), .B1(new_n419), .B2(new_n209), .ZN(new_n427));
  NOR4_X1   g0227(.A1(new_n286), .A2(new_n287), .A3(new_n417), .A4(G20), .ZN(new_n428));
  OAI21_X1  g0228(.A(G68), .B1(new_n427), .B2(new_n428), .ZN(new_n429));
  INV_X1    g0229(.A(new_n425), .ZN(new_n430));
  NAND3_X1  g0230(.A1(new_n429), .A2(KEYINPUT16), .A3(new_n430), .ZN(new_n431));
  NAND3_X1  g0231(.A1(new_n426), .A2(new_n431), .A3(new_n262), .ZN(new_n432));
  INV_X1    g0232(.A(KEYINPUT74), .ZN(new_n433));
  AOI21_X1  g0233(.A(new_n362), .B1(new_n208), .B2(G20), .ZN(new_n434));
  AOI22_X1  g0234(.A1(new_n434), .A2(new_n370), .B1(new_n260), .B2(new_n362), .ZN(new_n435));
  AND3_X1   g0235(.A1(new_n432), .A2(new_n433), .A3(new_n435), .ZN(new_n436));
  AOI21_X1  g0236(.A(new_n433), .B1(new_n432), .B2(new_n435), .ZN(new_n437));
  OAI21_X1  g0237(.A(new_n413), .B1(new_n436), .B2(new_n437), .ZN(new_n438));
  INV_X1    g0238(.A(KEYINPUT18), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n438), .A2(new_n439), .ZN(new_n440));
  NAND2_X1  g0240(.A1(new_n432), .A2(new_n435), .ZN(new_n441));
  NAND2_X1  g0241(.A1(new_n441), .A2(KEYINPUT74), .ZN(new_n442));
  NAND3_X1  g0242(.A1(new_n432), .A2(new_n433), .A3(new_n435), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  NAND3_X1  g0244(.A1(new_n444), .A2(KEYINPUT18), .A3(new_n413), .ZN(new_n445));
  INV_X1    g0245(.A(G190), .ZN(new_n446));
  OAI211_X1 g0246(.A(new_n446), .B(new_n399), .C1(new_n405), .C2(new_n407), .ZN(new_n447));
  INV_X1    g0247(.A(G200), .ZN(new_n448));
  OAI21_X1  g0248(.A(new_n448), .B1(new_n409), .B2(new_n410), .ZN(new_n449));
  NAND2_X1  g0249(.A1(new_n447), .A2(new_n449), .ZN(new_n450));
  XNOR2_X1  g0250(.A(KEYINPUT76), .B(KEYINPUT17), .ZN(new_n451));
  INV_X1    g0251(.A(new_n451), .ZN(new_n452));
  NAND4_X1  g0252(.A1(new_n450), .A2(new_n432), .A3(new_n435), .A4(new_n452), .ZN(new_n453));
  NAND3_X1  g0253(.A1(new_n450), .A2(new_n432), .A3(new_n435), .ZN(new_n454));
  INV_X1    g0254(.A(KEYINPUT17), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n455), .A2(KEYINPUT76), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n454), .A2(new_n456), .ZN(new_n457));
  AOI22_X1  g0257(.A1(new_n440), .A2(new_n445), .B1(new_n453), .B2(new_n457), .ZN(new_n458));
  NAND2_X1  g0258(.A1(G238), .A2(G1698), .ZN(new_n459));
  OAI211_X1 g0259(.A(new_n341), .B(new_n459), .C1(new_n229), .C2(G1698), .ZN(new_n460));
  OAI21_X1  g0260(.A(new_n460), .B1(G107), .B2(new_n341), .ZN(new_n461));
  NAND2_X1  g0261(.A1(new_n461), .A2(KEYINPUT69), .ZN(new_n462));
  INV_X1    g0262(.A(KEYINPUT69), .ZN(new_n463));
  OAI211_X1 g0263(.A(new_n460), .B(new_n463), .C1(G107), .C2(new_n341), .ZN(new_n464));
  NAND3_X1  g0264(.A1(new_n462), .A2(new_n289), .A3(new_n464), .ZN(new_n465));
  AOI22_X1  g0265(.A1(new_n348), .A2(G244), .B1(new_n352), .B2(new_n354), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  NOR2_X1   g0267(.A1(new_n467), .A2(new_n446), .ZN(new_n468));
  AOI21_X1  g0268(.A(new_n448), .B1(new_n465), .B2(new_n466), .ZN(new_n469));
  XOR2_X1   g0269(.A(KEYINPUT15), .B(G87), .Z(new_n470));
  INV_X1    g0270(.A(new_n470), .ZN(new_n471));
  NOR2_X1   g0271(.A1(new_n471), .A2(new_n364), .ZN(new_n472));
  OAI22_X1  g0272(.A1(new_n362), .A2(new_n367), .B1(new_n209), .B2(new_n225), .ZN(new_n473));
  OAI21_X1  g0273(.A(new_n262), .B1(new_n472), .B2(new_n473), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n260), .A2(new_n225), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n265), .A2(new_n371), .ZN(new_n476));
  OAI211_X1 g0276(.A(new_n474), .B(new_n475), .C1(new_n225), .C2(new_n476), .ZN(new_n477));
  NOR3_X1   g0277(.A1(new_n468), .A2(new_n469), .A3(new_n477), .ZN(new_n478));
  INV_X1    g0278(.A(new_n478), .ZN(new_n479));
  NAND3_X1  g0279(.A1(new_n398), .A2(new_n458), .A3(new_n479), .ZN(new_n480));
  INV_X1    g0280(.A(KEYINPUT14), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n224), .A2(new_n283), .ZN(new_n482));
  OAI211_X1 g0282(.A(new_n341), .B(new_n482), .C1(G232), .C2(new_n283), .ZN(new_n483));
  NOR2_X1   g0283(.A1(new_n291), .A2(new_n218), .ZN(new_n484));
  INV_X1    g0284(.A(new_n484), .ZN(new_n485));
  AOI21_X1  g0285(.A(new_n304), .B1(new_n483), .B2(new_n485), .ZN(new_n486));
  INV_X1    g0286(.A(new_n486), .ZN(new_n487));
  NAND3_X1  g0287(.A1(new_n304), .A2(G238), .A3(new_n346), .ZN(new_n488));
  NAND3_X1  g0288(.A1(new_n355), .A2(KEYINPUT72), .A3(new_n488), .ZN(new_n489));
  INV_X1    g0289(.A(new_n489), .ZN(new_n490));
  AOI21_X1  g0290(.A(KEYINPUT72), .B1(new_n355), .B2(new_n488), .ZN(new_n491));
  OAI21_X1  g0291(.A(new_n487), .B1(new_n490), .B2(new_n491), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n492), .A2(KEYINPUT13), .ZN(new_n493));
  INV_X1    g0293(.A(KEYINPUT13), .ZN(new_n494));
  OAI211_X1 g0294(.A(new_n487), .B(new_n494), .C1(new_n490), .C2(new_n491), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n493), .A2(new_n495), .ZN(new_n496));
  AOI21_X1  g0296(.A(new_n481), .B1(new_n496), .B2(G169), .ZN(new_n497));
  INV_X1    g0297(.A(new_n497), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n495), .A2(KEYINPUT73), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n355), .A2(new_n488), .ZN(new_n500));
  INV_X1    g0300(.A(KEYINPUT72), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  AOI21_X1  g0302(.A(new_n486), .B1(new_n502), .B2(new_n489), .ZN(new_n503));
  NOR2_X1   g0303(.A1(new_n503), .A2(new_n494), .ZN(new_n504));
  NOR2_X1   g0304(.A1(new_n499), .A2(new_n504), .ZN(new_n505));
  NOR3_X1   g0305(.A1(new_n503), .A2(KEYINPUT73), .A3(new_n494), .ZN(new_n506));
  OAI21_X1  g0306(.A(G179), .B1(new_n505), .B2(new_n506), .ZN(new_n507));
  AOI211_X1 g0307(.A(KEYINPUT14), .B(new_n357), .C1(new_n493), .C2(new_n495), .ZN(new_n508));
  INV_X1    g0308(.A(new_n508), .ZN(new_n509));
  NAND3_X1  g0309(.A1(new_n498), .A2(new_n507), .A3(new_n509), .ZN(new_n510));
  AOI22_X1  g0310(.A1(new_n366), .A2(G50), .B1(G20), .B2(new_n415), .ZN(new_n511));
  OAI21_X1  g0311(.A(new_n511), .B1(new_n364), .B2(new_n225), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n512), .A2(new_n262), .ZN(new_n513));
  XNOR2_X1  g0313(.A(new_n513), .B(KEYINPUT11), .ZN(new_n514));
  NAND3_X1  g0314(.A1(new_n265), .A2(G68), .A3(new_n371), .ZN(new_n515));
  NAND3_X1  g0315(.A1(new_n272), .A2(G20), .A3(new_n415), .ZN(new_n516));
  XNOR2_X1  g0316(.A(new_n516), .B(KEYINPUT12), .ZN(new_n517));
  NAND3_X1  g0317(.A1(new_n514), .A2(new_n515), .A3(new_n517), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n510), .A2(new_n518), .ZN(new_n519));
  OAI21_X1  g0319(.A(G190), .B1(new_n505), .B2(new_n506), .ZN(new_n520));
  INV_X1    g0320(.A(new_n518), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n496), .A2(G200), .ZN(new_n522));
  NAND3_X1  g0322(.A1(new_n520), .A2(new_n521), .A3(new_n522), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n467), .A2(new_n357), .ZN(new_n524));
  NAND3_X1  g0324(.A1(new_n465), .A2(new_n320), .A3(new_n466), .ZN(new_n525));
  NAND3_X1  g0325(.A1(new_n524), .A2(new_n477), .A3(new_n525), .ZN(new_n526));
  NAND3_X1  g0326(.A1(new_n519), .A2(new_n523), .A3(new_n526), .ZN(new_n527));
  NOR2_X1   g0327(.A1(new_n480), .A2(new_n527), .ZN(new_n528));
  NOR2_X1   g0328(.A1(new_n209), .A2(G107), .ZN(new_n529));
  XNOR2_X1  g0329(.A(new_n529), .B(KEYINPUT23), .ZN(new_n530));
  NAND3_X1  g0330(.A1(new_n209), .A2(G33), .A3(G116), .ZN(new_n531));
  XNOR2_X1  g0331(.A(new_n531), .B(KEYINPUT83), .ZN(new_n532));
  INV_X1    g0332(.A(KEYINPUT22), .ZN(new_n533));
  AOI21_X1  g0333(.A(G20), .B1(new_n292), .B2(new_n294), .ZN(new_n534));
  AOI21_X1  g0334(.A(new_n533), .B1(new_n534), .B2(G87), .ZN(new_n535));
  OAI211_X1 g0335(.A(new_n209), .B(G87), .C1(new_n286), .C2(new_n287), .ZN(new_n536));
  NOR2_X1   g0336(.A1(new_n536), .A2(KEYINPUT22), .ZN(new_n537));
  OAI211_X1 g0337(.A(new_n530), .B(new_n532), .C1(new_n535), .C2(new_n537), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n538), .A2(KEYINPUT84), .ZN(new_n539));
  XNOR2_X1  g0339(.A(new_n536), .B(KEYINPUT22), .ZN(new_n540));
  INV_X1    g0340(.A(KEYINPUT84), .ZN(new_n541));
  NAND4_X1  g0341(.A1(new_n540), .A2(new_n541), .A3(new_n530), .A4(new_n532), .ZN(new_n542));
  NAND3_X1  g0342(.A1(new_n539), .A2(new_n542), .A3(KEYINPUT24), .ZN(new_n543));
  INV_X1    g0343(.A(KEYINPUT24), .ZN(new_n544));
  NAND3_X1  g0344(.A1(new_n538), .A2(KEYINPUT84), .A3(new_n544), .ZN(new_n545));
  NAND3_X1  g0345(.A1(new_n543), .A2(new_n262), .A3(new_n545), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n217), .A2(new_n283), .ZN(new_n547));
  OAI211_X1 g0347(.A(new_n341), .B(new_n547), .C1(G257), .C2(new_n283), .ZN(new_n548));
  INV_X1    g0348(.A(new_n548), .ZN(new_n549));
  INV_X1    g0349(.A(G294), .ZN(new_n550));
  NOR2_X1   g0350(.A1(new_n291), .A2(new_n550), .ZN(new_n551));
  OAI21_X1  g0351(.A(new_n289), .B1(new_n549), .B2(new_n551), .ZN(new_n552));
  NAND3_X1  g0352(.A1(new_n302), .A2(G264), .A3(new_n304), .ZN(new_n553));
  NAND3_X1  g0353(.A1(new_n552), .A2(new_n309), .A3(new_n553), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n554), .A2(new_n448), .ZN(new_n555));
  NAND4_X1  g0355(.A1(new_n552), .A2(new_n446), .A3(new_n309), .A4(new_n553), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n272), .A2(new_n529), .ZN(new_n558));
  XNOR2_X1  g0358(.A(new_n558), .B(KEYINPUT25), .ZN(new_n559));
  NOR3_X1   g0359(.A1(new_n268), .A2(new_n262), .A3(new_n260), .ZN(new_n560));
  AOI21_X1  g0360(.A(new_n559), .B1(G107), .B2(new_n560), .ZN(new_n561));
  NAND3_X1  g0361(.A1(new_n546), .A2(new_n557), .A3(new_n561), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n562), .A2(KEYINPUT85), .ZN(new_n563));
  INV_X1    g0363(.A(KEYINPUT85), .ZN(new_n564));
  NAND4_X1  g0364(.A1(new_n546), .A2(new_n557), .A3(new_n564), .A4(new_n561), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n563), .A2(new_n565), .ZN(new_n566));
  OAI21_X1  g0366(.A(G244), .B1(new_n286), .B2(new_n287), .ZN(new_n567));
  INV_X1    g0367(.A(KEYINPUT4), .ZN(new_n568));
  AOI22_X1  g0368(.A1(new_n567), .A2(new_n568), .B1(G33), .B2(G283), .ZN(new_n569));
  NAND4_X1  g0369(.A1(new_n341), .A2(KEYINPUT4), .A3(G244), .A4(new_n283), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n569), .A2(new_n570), .ZN(new_n571));
  AOI21_X1  g0371(.A(new_n568), .B1(new_n341), .B2(G250), .ZN(new_n572));
  NOR2_X1   g0372(.A1(new_n572), .A2(new_n283), .ZN(new_n573));
  OAI21_X1  g0373(.A(new_n289), .B1(new_n571), .B2(new_n573), .ZN(new_n574));
  NOR3_X1   g0374(.A1(new_n308), .A2(new_n219), .A3(new_n289), .ZN(new_n575));
  INV_X1    g0375(.A(new_n575), .ZN(new_n576));
  NAND3_X1  g0376(.A1(new_n574), .A2(new_n309), .A3(new_n576), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n577), .A2(G169), .ZN(new_n578));
  NAND4_X1  g0378(.A1(new_n574), .A2(G179), .A3(new_n309), .A4(new_n576), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n260), .A2(new_n218), .ZN(new_n580));
  OAI21_X1  g0380(.A(G107), .B1(new_n427), .B2(new_n428), .ZN(new_n581));
  INV_X1    g0381(.A(KEYINPUT6), .ZN(new_n582));
  NOR2_X1   g0382(.A1(new_n218), .A2(new_n249), .ZN(new_n583));
  NOR2_X1   g0383(.A1(G97), .A2(G107), .ZN(new_n584));
  OAI21_X1  g0384(.A(new_n582), .B1(new_n583), .B2(new_n584), .ZN(new_n585));
  NAND3_X1  g0385(.A1(new_n249), .A2(KEYINPUT6), .A3(G97), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n587), .A2(G20), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n366), .A2(G77), .ZN(new_n589));
  NAND3_X1  g0389(.A1(new_n581), .A2(new_n588), .A3(new_n589), .ZN(new_n590));
  AOI22_X1  g0390(.A1(new_n590), .A2(new_n262), .B1(G97), .B2(new_n560), .ZN(new_n591));
  AOI22_X1  g0391(.A1(new_n578), .A2(new_n579), .B1(new_n580), .B2(new_n591), .ZN(new_n592));
  INV_X1    g0392(.A(new_n592), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n560), .A2(G97), .ZN(new_n594));
  AOI21_X1  g0394(.A(new_n249), .B1(new_n418), .B2(new_n420), .ZN(new_n595));
  INV_X1    g0395(.A(new_n589), .ZN(new_n596));
  AOI21_X1  g0396(.A(new_n209), .B1(new_n585), .B2(new_n586), .ZN(new_n597));
  NOR3_X1   g0397(.A1(new_n595), .A2(new_n596), .A3(new_n597), .ZN(new_n598));
  INV_X1    g0398(.A(new_n262), .ZN(new_n599));
  OAI211_X1 g0399(.A(new_n580), .B(new_n594), .C1(new_n598), .C2(new_n599), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n600), .A2(KEYINPUT78), .ZN(new_n601));
  INV_X1    g0401(.A(KEYINPUT78), .ZN(new_n602));
  NAND3_X1  g0402(.A1(new_n591), .A2(new_n602), .A3(new_n580), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n601), .A2(new_n603), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n577), .A2(new_n448), .ZN(new_n605));
  OAI211_X1 g0405(.A(new_n569), .B(new_n570), .C1(new_n283), .C2(new_n572), .ZN(new_n606));
  AOI21_X1  g0406(.A(new_n575), .B1(new_n606), .B2(new_n289), .ZN(new_n607));
  NAND3_X1  g0407(.A1(new_n607), .A2(new_n446), .A3(new_n309), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n605), .A2(new_n608), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n604), .A2(new_n609), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n546), .A2(new_n561), .ZN(new_n611));
  NOR2_X1   g0411(.A1(new_n554), .A2(G179), .ZN(new_n612));
  AOI21_X1  g0412(.A(new_n612), .B1(new_n357), .B2(new_n554), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n611), .A2(new_n613), .ZN(new_n614));
  INV_X1    g0414(.A(KEYINPUT19), .ZN(new_n615));
  OAI21_X1  g0415(.A(new_n615), .B1(new_n364), .B2(new_n218), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n534), .A2(G68), .ZN(new_n617));
  NOR3_X1   g0417(.A1(G87), .A2(G97), .A3(G107), .ZN(new_n618));
  XNOR2_X1  g0418(.A(new_n618), .B(KEYINPUT79), .ZN(new_n619));
  AOI21_X1  g0419(.A(G20), .B1(new_n484), .B2(KEYINPUT19), .ZN(new_n620));
  OAI211_X1 g0420(.A(new_n616), .B(new_n617), .C1(new_n619), .C2(new_n620), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n621), .A2(new_n262), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n560), .A2(new_n470), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n471), .A2(new_n260), .ZN(new_n624));
  NAND3_X1  g0424(.A1(new_n622), .A2(new_n623), .A3(new_n624), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n226), .A2(G1698), .ZN(new_n626));
  OAI221_X1 g0426(.A(new_n626), .B1(G238), .B2(G1698), .C1(new_n286), .C2(new_n287), .ZN(new_n627));
  NAND2_X1  g0427(.A1(G33), .A2(G116), .ZN(new_n628));
  AOI21_X1  g0428(.A(new_n304), .B1(new_n627), .B2(new_n628), .ZN(new_n629));
  NOR2_X1   g0429(.A1(new_n298), .A2(G250), .ZN(new_n630));
  NOR2_X1   g0430(.A1(new_n306), .A2(G274), .ZN(new_n631));
  NOR3_X1   g0431(.A1(new_n630), .A2(new_n631), .A3(new_n289), .ZN(new_n632));
  NOR2_X1   g0432(.A1(new_n629), .A2(new_n632), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n633), .A2(new_n320), .ZN(new_n634));
  INV_X1    g0434(.A(new_n633), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n635), .A2(new_n357), .ZN(new_n636));
  NAND3_X1  g0436(.A1(new_n625), .A2(new_n634), .A3(new_n636), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n635), .A2(G200), .ZN(new_n638));
  AOI22_X1  g0438(.A1(new_n621), .A2(new_n262), .B1(new_n260), .B2(new_n471), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n633), .A2(G190), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n560), .A2(G87), .ZN(new_n641));
  NAND4_X1  g0441(.A1(new_n638), .A2(new_n639), .A3(new_n640), .A4(new_n641), .ZN(new_n642));
  AND2_X1   g0442(.A1(new_n637), .A2(new_n642), .ZN(new_n643));
  AND4_X1   g0443(.A1(new_n593), .A2(new_n610), .A3(new_n614), .A4(new_n643), .ZN(new_n644));
  AND4_X1   g0444(.A1(new_n340), .A2(new_n528), .A3(new_n566), .A4(new_n644), .ZN(G372));
  INV_X1    g0445(.A(new_n435), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n429), .A2(new_n430), .ZN(new_n647));
  AOI21_X1  g0447(.A(new_n599), .B1(new_n647), .B2(new_n414), .ZN(new_n648));
  AOI21_X1  g0448(.A(new_n646), .B1(new_n648), .B2(new_n431), .ZN(new_n649));
  OAI21_X1  g0449(.A(new_n439), .B1(new_n649), .B2(new_n412), .ZN(new_n650));
  NAND3_X1  g0450(.A1(new_n413), .A2(new_n441), .A3(KEYINPUT18), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  INV_X1    g0452(.A(new_n652), .ZN(new_n653));
  INV_X1    g0453(.A(new_n506), .ZN(new_n654));
  NAND3_X1  g0454(.A1(new_n493), .A2(KEYINPUT73), .A3(new_n495), .ZN(new_n655));
  AOI21_X1  g0455(.A(new_n446), .B1(new_n654), .B2(new_n655), .ZN(new_n656));
  INV_X1    g0456(.A(new_n522), .ZN(new_n657));
  NOR3_X1   g0457(.A1(new_n656), .A2(new_n657), .A3(new_n518), .ZN(new_n658));
  OAI21_X1  g0458(.A(new_n519), .B1(new_n658), .B2(new_n526), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n457), .A2(new_n453), .ZN(new_n660));
  AOI21_X1  g0460(.A(new_n653), .B1(new_n659), .B2(new_n660), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n393), .A2(new_n397), .ZN(new_n662));
  INV_X1    g0462(.A(new_n662), .ZN(new_n663));
  OAI22_X1  g0463(.A1(new_n661), .A2(new_n663), .B1(new_n374), .B2(new_n359), .ZN(new_n664));
  INV_X1    g0464(.A(new_n664), .ZN(new_n665));
  AOI22_X1  g0465(.A1(new_n601), .A2(new_n603), .B1(new_n608), .B2(new_n605), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n637), .A2(new_n642), .ZN(new_n667));
  NOR3_X1   g0467(.A1(new_n666), .A2(new_n592), .A3(new_n667), .ZN(new_n668));
  NAND3_X1  g0468(.A1(new_n614), .A2(new_n322), .A3(new_n337), .ZN(new_n669));
  NAND3_X1  g0469(.A1(new_n668), .A2(new_n566), .A3(new_n669), .ZN(new_n670));
  INV_X1    g0470(.A(new_n309), .ZN(new_n671));
  AOI211_X1 g0471(.A(new_n671), .B(new_n575), .C1(new_n606), .C2(new_n289), .ZN(new_n672));
  OAI21_X1  g0472(.A(new_n579), .B1(new_n672), .B2(new_n357), .ZN(new_n673));
  NAND4_X1  g0473(.A1(new_n673), .A2(new_n637), .A3(new_n642), .A4(new_n600), .ZN(new_n674));
  INV_X1    g0474(.A(KEYINPUT26), .ZN(new_n675));
  OAI21_X1  g0475(.A(KEYINPUT86), .B1(new_n674), .B2(new_n675), .ZN(new_n676));
  NAND3_X1  g0476(.A1(new_n673), .A2(new_n601), .A3(new_n603), .ZN(new_n677));
  OAI21_X1  g0477(.A(new_n675), .B1(new_n677), .B2(new_n667), .ZN(new_n678));
  INV_X1    g0478(.A(KEYINPUT86), .ZN(new_n679));
  NAND4_X1  g0479(.A1(new_n643), .A2(new_n679), .A3(new_n592), .A4(KEYINPUT26), .ZN(new_n680));
  NAND3_X1  g0480(.A1(new_n676), .A2(new_n678), .A3(new_n680), .ZN(new_n681));
  NAND3_X1  g0481(.A1(new_n670), .A2(new_n637), .A3(new_n681), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n528), .A2(new_n682), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n665), .A2(new_n683), .ZN(G369));
  NAND2_X1  g0484(.A1(new_n337), .A2(new_n322), .ZN(new_n685));
  INV_X1    g0485(.A(KEYINPUT87), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n272), .A2(new_n209), .ZN(new_n687));
  INV_X1    g0487(.A(new_n687), .ZN(new_n688));
  INV_X1    g0488(.A(KEYINPUT27), .ZN(new_n689));
  OAI21_X1  g0489(.A(new_n686), .B1(new_n688), .B2(new_n689), .ZN(new_n690));
  INV_X1    g0490(.A(G213), .ZN(new_n691));
  AOI21_X1  g0491(.A(new_n691), .B1(new_n688), .B2(new_n689), .ZN(new_n692));
  NAND3_X1  g0492(.A1(new_n687), .A2(KEYINPUT87), .A3(KEYINPUT27), .ZN(new_n693));
  NAND3_X1  g0493(.A1(new_n690), .A2(new_n692), .A3(new_n693), .ZN(new_n694));
  INV_X1    g0494(.A(G343), .ZN(new_n695));
  NOR2_X1   g0495(.A1(new_n694), .A2(new_n695), .ZN(new_n696));
  INV_X1    g0496(.A(new_n696), .ZN(new_n697));
  NOR2_X1   g0497(.A1(new_n697), .A2(new_n282), .ZN(new_n698));
  INV_X1    g0498(.A(new_n698), .ZN(new_n699));
  MUX2_X1   g0499(.A(new_n685), .B(new_n340), .S(new_n699), .Z(new_n700));
  NAND2_X1  g0500(.A1(new_n700), .A2(G330), .ZN(new_n701));
  INV_X1    g0501(.A(new_n614), .ZN(new_n702));
  NAND2_X1  g0502(.A1(new_n702), .A2(new_n697), .ZN(new_n703));
  AOI22_X1  g0503(.A1(new_n563), .A2(new_n565), .B1(new_n611), .B2(new_n696), .ZN(new_n704));
  OAI21_X1  g0504(.A(new_n703), .B1(new_n704), .B2(new_n702), .ZN(new_n705));
  NOR2_X1   g0505(.A1(new_n701), .A2(new_n705), .ZN(new_n706));
  INV_X1    g0506(.A(new_n706), .ZN(new_n707));
  NAND4_X1  g0507(.A1(new_n704), .A2(new_n685), .A3(new_n614), .A4(new_n697), .ZN(new_n708));
  INV_X1    g0508(.A(KEYINPUT88), .ZN(new_n709));
  NAND3_X1  g0509(.A1(new_n708), .A2(new_n709), .A3(new_n703), .ZN(new_n710));
  INV_X1    g0510(.A(new_n710), .ZN(new_n711));
  AOI21_X1  g0511(.A(new_n709), .B1(new_n708), .B2(new_n703), .ZN(new_n712));
  OAI21_X1  g0512(.A(new_n707), .B1(new_n711), .B2(new_n712), .ZN(G399));
  INV_X1    g0513(.A(new_n212), .ZN(new_n714));
  NOR2_X1   g0514(.A1(new_n714), .A2(G41), .ZN(new_n715));
  INV_X1    g0515(.A(new_n715), .ZN(new_n716));
  NAND2_X1  g0516(.A1(new_n619), .A2(new_n251), .ZN(new_n717));
  INV_X1    g0517(.A(new_n717), .ZN(new_n718));
  NAND3_X1  g0518(.A1(new_n716), .A2(G1), .A3(new_n718), .ZN(new_n719));
  OAI21_X1  g0519(.A(new_n719), .B1(new_n236), .B2(new_n716), .ZN(new_n720));
  XNOR2_X1  g0520(.A(new_n720), .B(KEYINPUT28), .ZN(new_n721));
  NOR2_X1   g0521(.A1(new_n666), .A2(new_n592), .ZN(new_n722));
  NAND4_X1  g0522(.A1(new_n566), .A2(new_n669), .A3(new_n722), .A4(new_n642), .ZN(new_n723));
  OAI21_X1  g0523(.A(KEYINPUT26), .B1(new_n677), .B2(new_n667), .ZN(new_n724));
  NAND3_X1  g0524(.A1(new_n643), .A2(new_n675), .A3(new_n592), .ZN(new_n725));
  AND3_X1   g0525(.A1(new_n724), .A2(new_n637), .A3(new_n725), .ZN(new_n726));
  AND2_X1   g0526(.A1(new_n723), .A2(new_n726), .ZN(new_n727));
  OAI21_X1  g0527(.A(KEYINPUT29), .B1(new_n727), .B2(new_n696), .ZN(new_n728));
  INV_X1    g0528(.A(KEYINPUT29), .ZN(new_n729));
  NAND3_X1  g0529(.A1(new_n682), .A2(new_n729), .A3(new_n697), .ZN(new_n730));
  NAND2_X1  g0530(.A1(new_n728), .A2(new_n730), .ZN(new_n731));
  NAND4_X1  g0531(.A1(new_n644), .A2(new_n340), .A3(new_n566), .A4(new_n697), .ZN(new_n732));
  INV_X1    g0532(.A(KEYINPUT31), .ZN(new_n733));
  NOR2_X1   g0533(.A1(new_n554), .A2(new_n635), .ZN(new_n734));
  NAND2_X1  g0534(.A1(new_n321), .A2(KEYINPUT89), .ZN(new_n735));
  INV_X1    g0535(.A(KEYINPUT89), .ZN(new_n736));
  OAI21_X1  g0536(.A(new_n736), .B1(new_n310), .B2(new_n320), .ZN(new_n737));
  NAND2_X1  g0537(.A1(new_n735), .A2(new_n737), .ZN(new_n738));
  NAND3_X1  g0538(.A1(new_n734), .A2(new_n738), .A3(new_n607), .ZN(new_n739));
  INV_X1    g0539(.A(KEYINPUT90), .ZN(new_n740));
  INV_X1    g0540(.A(KEYINPUT30), .ZN(new_n741));
  NAND3_X1  g0541(.A1(new_n739), .A2(new_n740), .A3(new_n741), .ZN(new_n742));
  INV_X1    g0542(.A(new_n742), .ZN(new_n743));
  AOI21_X1  g0543(.A(new_n740), .B1(new_n739), .B2(new_n741), .ZN(new_n744));
  NAND4_X1  g0544(.A1(new_n734), .A2(new_n738), .A3(KEYINPUT30), .A4(new_n607), .ZN(new_n745));
  AND2_X1   g0545(.A1(new_n635), .A2(new_n310), .ZN(new_n746));
  NAND4_X1  g0546(.A1(new_n746), .A2(new_n320), .A3(new_n554), .A4(new_n577), .ZN(new_n747));
  NAND2_X1  g0547(.A1(new_n745), .A2(new_n747), .ZN(new_n748));
  NOR3_X1   g0548(.A1(new_n743), .A2(new_n744), .A3(new_n748), .ZN(new_n749));
  OAI21_X1  g0549(.A(new_n733), .B1(new_n749), .B2(new_n697), .ZN(new_n750));
  AND2_X1   g0550(.A1(new_n739), .A2(new_n741), .ZN(new_n751));
  OAI211_X1 g0551(.A(KEYINPUT31), .B(new_n696), .C1(new_n751), .C2(new_n748), .ZN(new_n752));
  NAND3_X1  g0552(.A1(new_n732), .A2(new_n750), .A3(new_n752), .ZN(new_n753));
  AND2_X1   g0553(.A1(new_n753), .A2(G330), .ZN(new_n754));
  NOR2_X1   g0554(.A1(new_n731), .A2(new_n754), .ZN(new_n755));
  NAND2_X1  g0555(.A1(new_n755), .A2(KEYINPUT91), .ZN(new_n756));
  INV_X1    g0556(.A(KEYINPUT91), .ZN(new_n757));
  OAI21_X1  g0557(.A(new_n757), .B1(new_n731), .B2(new_n754), .ZN(new_n758));
  NAND2_X1  g0558(.A1(new_n756), .A2(new_n758), .ZN(new_n759));
  OAI21_X1  g0559(.A(new_n721), .B1(new_n759), .B2(G1), .ZN(new_n760));
  XOR2_X1   g0560(.A(new_n760), .B(KEYINPUT92), .Z(G364));
  INV_X1    g0561(.A(new_n701), .ZN(new_n762));
  NOR2_X1   g0562(.A1(new_n271), .A2(G20), .ZN(new_n763));
  NAND2_X1  g0563(.A1(new_n763), .A2(G45), .ZN(new_n764));
  NAND3_X1  g0564(.A1(new_n716), .A2(G1), .A3(new_n764), .ZN(new_n765));
  INV_X1    g0565(.A(new_n765), .ZN(new_n766));
  NOR2_X1   g0566(.A1(new_n762), .A2(new_n766), .ZN(new_n767));
  OAI21_X1  g0567(.A(new_n767), .B1(G330), .B2(new_n700), .ZN(new_n768));
  AOI21_X1  g0568(.A(new_n233), .B1(G20), .B2(new_n357), .ZN(new_n769));
  NOR3_X1   g0569(.A1(G13), .A2(G20), .A3(G33), .ZN(new_n770));
  NOR2_X1   g0570(.A1(new_n769), .A2(new_n770), .ZN(new_n771));
  INV_X1    g0571(.A(new_n771), .ZN(new_n772));
  NAND2_X1  g0572(.A1(new_n256), .A2(G45), .ZN(new_n773));
  NAND2_X1  g0573(.A1(new_n212), .A2(new_n419), .ZN(new_n774));
  AOI21_X1  g0574(.A(new_n774), .B1(new_n297), .B2(new_n237), .ZN(new_n775));
  AOI22_X1  g0575(.A1(new_n773), .A2(new_n775), .B1(new_n251), .B2(new_n714), .ZN(new_n776));
  XOR2_X1   g0576(.A(G355), .B(KEYINPUT93), .Z(new_n777));
  NAND3_X1  g0577(.A1(new_n777), .A2(new_n212), .A3(new_n341), .ZN(new_n778));
  AOI21_X1  g0578(.A(new_n772), .B1(new_n776), .B2(new_n778), .ZN(new_n779));
  NAND2_X1  g0579(.A1(new_n446), .A2(G20), .ZN(new_n780));
  XNOR2_X1  g0580(.A(new_n780), .B(KEYINPUT95), .ZN(new_n781));
  NOR2_X1   g0581(.A1(G179), .A2(G200), .ZN(new_n782));
  INV_X1    g0582(.A(new_n782), .ZN(new_n783));
  NOR2_X1   g0583(.A1(new_n781), .A2(new_n783), .ZN(new_n784));
  NAND2_X1  g0584(.A1(G20), .A2(G179), .ZN(new_n785));
  NOR3_X1   g0585(.A1(new_n785), .A2(new_n446), .A3(G200), .ZN(new_n786));
  AOI22_X1  g0586(.A1(new_n784), .A2(G329), .B1(G322), .B2(new_n786), .ZN(new_n787));
  INV_X1    g0587(.A(new_n785), .ZN(new_n788));
  NAND3_X1  g0588(.A1(new_n788), .A2(G190), .A3(G200), .ZN(new_n789));
  INV_X1    g0589(.A(new_n789), .ZN(new_n790));
  NAND2_X1  g0590(.A1(new_n790), .A2(G326), .ZN(new_n791));
  NAND3_X1  g0591(.A1(new_n787), .A2(new_n419), .A3(new_n791), .ZN(new_n792));
  NOR2_X1   g0592(.A1(new_n448), .A2(G179), .ZN(new_n793));
  INV_X1    g0593(.A(new_n793), .ZN(new_n794));
  NOR3_X1   g0594(.A1(new_n794), .A2(new_n209), .A3(new_n446), .ZN(new_n795));
  INV_X1    g0595(.A(new_n795), .ZN(new_n796));
  NOR2_X1   g0596(.A1(new_n796), .A2(new_n293), .ZN(new_n797));
  NOR3_X1   g0597(.A1(new_n785), .A2(new_n448), .A3(G190), .ZN(new_n798));
  INV_X1    g0598(.A(new_n798), .ZN(new_n799));
  OR2_X1    g0599(.A1(KEYINPUT33), .A2(G317), .ZN(new_n800));
  NAND2_X1  g0600(.A1(KEYINPUT33), .A2(G317), .ZN(new_n801));
  AOI21_X1  g0601(.A(new_n799), .B1(new_n800), .B2(new_n801), .ZN(new_n802));
  AOI21_X1  g0602(.A(new_n209), .B1(new_n782), .B2(G190), .ZN(new_n803));
  NOR2_X1   g0603(.A1(new_n803), .A2(new_n550), .ZN(new_n804));
  NOR4_X1   g0604(.A1(new_n792), .A2(new_n797), .A3(new_n802), .A4(new_n804), .ZN(new_n805));
  INV_X1    g0605(.A(G283), .ZN(new_n806));
  NOR2_X1   g0606(.A1(new_n781), .A2(new_n794), .ZN(new_n807));
  INV_X1    g0607(.A(new_n807), .ZN(new_n808));
  OAI21_X1  g0608(.A(new_n805), .B1(new_n806), .B2(new_n808), .ZN(new_n809));
  NOR3_X1   g0609(.A1(new_n785), .A2(G190), .A3(G200), .ZN(new_n810));
  AOI21_X1  g0610(.A(new_n809), .B1(G311), .B2(new_n810), .ZN(new_n811));
  XNOR2_X1  g0611(.A(new_n811), .B(KEYINPUT97), .ZN(new_n812));
  NAND2_X1  g0612(.A1(new_n784), .A2(G159), .ZN(new_n813));
  XNOR2_X1  g0613(.A(new_n813), .B(KEYINPUT32), .ZN(new_n814));
  AOI211_X1 g0614(.A(new_n419), .B(new_n814), .C1(G50), .C2(new_n790), .ZN(new_n815));
  NAND2_X1  g0615(.A1(new_n798), .A2(G68), .ZN(new_n816));
  NAND2_X1  g0616(.A1(new_n795), .A2(G87), .ZN(new_n817));
  INV_X1    g0617(.A(KEYINPUT96), .ZN(new_n818));
  AND2_X1   g0618(.A1(new_n803), .A2(new_n818), .ZN(new_n819));
  NOR2_X1   g0619(.A1(new_n803), .A2(new_n818), .ZN(new_n820));
  NOR2_X1   g0620(.A1(new_n819), .A2(new_n820), .ZN(new_n821));
  INV_X1    g0621(.A(new_n821), .ZN(new_n822));
  NAND2_X1  g0622(.A1(new_n822), .A2(G97), .ZN(new_n823));
  INV_X1    g0623(.A(new_n810), .ZN(new_n824));
  INV_X1    g0624(.A(new_n786), .ZN(new_n825));
  OAI22_X1  g0625(.A1(new_n824), .A2(new_n225), .B1(new_n825), .B2(new_n228), .ZN(new_n826));
  NAND2_X1  g0626(.A1(new_n826), .A2(KEYINPUT94), .ZN(new_n827));
  NAND2_X1  g0627(.A1(new_n823), .A2(new_n827), .ZN(new_n828));
  NOR2_X1   g0628(.A1(new_n826), .A2(KEYINPUT94), .ZN(new_n829));
  NOR2_X1   g0629(.A1(new_n808), .A2(new_n249), .ZN(new_n830));
  NOR3_X1   g0630(.A1(new_n828), .A2(new_n829), .A3(new_n830), .ZN(new_n831));
  NAND4_X1  g0631(.A1(new_n815), .A2(new_n816), .A3(new_n817), .A4(new_n831), .ZN(new_n832));
  NAND2_X1  g0632(.A1(new_n812), .A2(new_n832), .ZN(new_n833));
  AOI211_X1 g0633(.A(new_n779), .B(new_n765), .C1(new_n833), .C2(new_n769), .ZN(new_n834));
  XOR2_X1   g0634(.A(new_n770), .B(KEYINPUT98), .Z(new_n835));
  OAI21_X1  g0635(.A(new_n834), .B1(new_n700), .B2(new_n835), .ZN(new_n836));
  AND2_X1   g0636(.A1(new_n768), .A2(new_n836), .ZN(new_n837));
  INV_X1    g0637(.A(new_n837), .ZN(G396));
  INV_X1    g0638(.A(KEYINPUT100), .ZN(new_n839));
  NAND2_X1  g0639(.A1(new_n526), .A2(new_n839), .ZN(new_n840));
  NAND4_X1  g0640(.A1(new_n524), .A2(KEYINPUT100), .A3(new_n477), .A4(new_n525), .ZN(new_n841));
  AOI21_X1  g0641(.A(new_n478), .B1(new_n840), .B2(new_n841), .ZN(new_n842));
  NAND3_X1  g0642(.A1(new_n682), .A2(new_n697), .A3(new_n842), .ZN(new_n843));
  AND2_X1   g0643(.A1(new_n682), .A2(new_n697), .ZN(new_n844));
  NOR2_X1   g0644(.A1(new_n526), .A2(new_n697), .ZN(new_n845));
  NAND2_X1  g0645(.A1(new_n477), .A2(new_n696), .ZN(new_n846));
  AOI21_X1  g0646(.A(new_n845), .B1(new_n842), .B2(new_n846), .ZN(new_n847));
  INV_X1    g0647(.A(new_n847), .ZN(new_n848));
  OAI21_X1  g0648(.A(new_n843), .B1(new_n844), .B2(new_n848), .ZN(new_n849));
  XNOR2_X1  g0649(.A(new_n849), .B(new_n754), .ZN(new_n850));
  NAND2_X1  g0650(.A1(new_n850), .A2(new_n765), .ZN(new_n851));
  NOR2_X1   g0651(.A1(G13), .A2(G33), .ZN(new_n852));
  NAND2_X1  g0652(.A1(new_n847), .A2(new_n852), .ZN(new_n853));
  NOR2_X1   g0653(.A1(new_n769), .A2(new_n852), .ZN(new_n854));
  XNOR2_X1  g0654(.A(new_n854), .B(KEYINPUT99), .ZN(new_n855));
  NAND2_X1  g0655(.A1(new_n855), .A2(new_n225), .ZN(new_n856));
  AOI22_X1  g0656(.A1(G116), .A2(new_n810), .B1(new_n786), .B2(G294), .ZN(new_n857));
  NAND2_X1  g0657(.A1(new_n784), .A2(G311), .ZN(new_n858));
  NAND2_X1  g0658(.A1(new_n798), .A2(G283), .ZN(new_n859));
  NAND4_X1  g0659(.A1(new_n823), .A2(new_n857), .A3(new_n858), .A4(new_n859), .ZN(new_n860));
  NOR2_X1   g0660(.A1(new_n796), .A2(new_n249), .ZN(new_n861));
  NOR2_X1   g0661(.A1(new_n789), .A2(new_n293), .ZN(new_n862));
  OAI21_X1  g0662(.A(new_n419), .B1(new_n808), .B2(new_n216), .ZN(new_n863));
  NOR4_X1   g0663(.A1(new_n860), .A2(new_n861), .A3(new_n862), .A4(new_n863), .ZN(new_n864));
  NAND2_X1  g0664(.A1(new_n790), .A2(G137), .ZN(new_n865));
  AOI22_X1  g0665(.A1(G143), .A2(new_n786), .B1(new_n810), .B2(G159), .ZN(new_n866));
  OAI211_X1 g0666(.A(new_n865), .B(new_n866), .C1(new_n365), .C2(new_n799), .ZN(new_n867));
  INV_X1    g0667(.A(KEYINPUT34), .ZN(new_n868));
  OAI221_X1 g0668(.A(new_n341), .B1(new_n202), .B2(new_n796), .C1(new_n867), .C2(new_n868), .ZN(new_n869));
  AND2_X1   g0669(.A1(new_n867), .A2(new_n868), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n807), .A2(G68), .ZN(new_n871));
  OAI21_X1  g0671(.A(new_n871), .B1(new_n228), .B2(new_n803), .ZN(new_n872));
  INV_X1    g0672(.A(new_n784), .ZN(new_n873));
  INV_X1    g0673(.A(G132), .ZN(new_n874));
  NOR2_X1   g0674(.A1(new_n873), .A2(new_n874), .ZN(new_n875));
  NOR4_X1   g0675(.A1(new_n869), .A2(new_n870), .A3(new_n872), .A4(new_n875), .ZN(new_n876));
  OAI21_X1  g0676(.A(new_n769), .B1(new_n864), .B2(new_n876), .ZN(new_n877));
  NAND4_X1  g0677(.A1(new_n853), .A2(new_n766), .A3(new_n856), .A4(new_n877), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n851), .A2(new_n878), .ZN(G384));
  INV_X1    g0679(.A(new_n694), .ZN(new_n880));
  OAI21_X1  g0680(.A(new_n880), .B1(new_n436), .B2(new_n437), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n413), .A2(new_n441), .ZN(new_n882));
  NAND3_X1  g0682(.A1(new_n881), .A2(new_n454), .A3(new_n882), .ZN(new_n883));
  AOI22_X1  g0683(.A1(new_n650), .A2(new_n651), .B1(new_n457), .B2(new_n453), .ZN(new_n884));
  OAI211_X1 g0684(.A(KEYINPUT37), .B(new_n883), .C1(new_n884), .C2(new_n881), .ZN(new_n885));
  INV_X1    g0685(.A(KEYINPUT103), .ZN(new_n886));
  INV_X1    g0686(.A(new_n454), .ZN(new_n887));
  AOI21_X1  g0687(.A(new_n887), .B1(new_n444), .B2(new_n413), .ZN(new_n888));
  AOI21_X1  g0688(.A(KEYINPUT37), .B1(new_n444), .B2(new_n880), .ZN(new_n889));
  AOI21_X1  g0689(.A(KEYINPUT38), .B1(new_n888), .B2(new_n889), .ZN(new_n890));
  AND3_X1   g0690(.A1(new_n885), .A2(new_n886), .A3(new_n890), .ZN(new_n891));
  AOI21_X1  g0691(.A(new_n886), .B1(new_n885), .B2(new_n890), .ZN(new_n892));
  NOR2_X1   g0692(.A1(new_n891), .A2(new_n892), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n440), .A2(new_n445), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n894), .A2(new_n660), .ZN(new_n895));
  AOI21_X1  g0695(.A(KEYINPUT16), .B1(new_n429), .B2(new_n430), .ZN(new_n896));
  OAI21_X1  g0696(.A(KEYINPUT101), .B1(new_n896), .B2(new_n599), .ZN(new_n897));
  INV_X1    g0697(.A(KEYINPUT101), .ZN(new_n898));
  NAND3_X1  g0698(.A1(new_n426), .A2(new_n898), .A3(new_n262), .ZN(new_n899));
  NAND3_X1  g0699(.A1(new_n897), .A2(new_n431), .A3(new_n899), .ZN(new_n900));
  INV_X1    g0700(.A(KEYINPUT102), .ZN(new_n901));
  AND3_X1   g0701(.A1(new_n900), .A2(new_n901), .A3(new_n435), .ZN(new_n902));
  AOI21_X1  g0702(.A(new_n901), .B1(new_n900), .B2(new_n435), .ZN(new_n903));
  NOR2_X1   g0703(.A1(new_n902), .A2(new_n903), .ZN(new_n904));
  NAND3_X1  g0704(.A1(new_n895), .A2(new_n880), .A3(new_n904), .ZN(new_n905));
  INV_X1    g0705(.A(KEYINPUT37), .ZN(new_n906));
  AOI21_X1  g0706(.A(new_n887), .B1(new_n904), .B2(new_n413), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n900), .A2(new_n435), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n908), .A2(KEYINPUT102), .ZN(new_n909));
  NAND3_X1  g0709(.A1(new_n900), .A2(new_n901), .A3(new_n435), .ZN(new_n910));
  NAND3_X1  g0710(.A1(new_n909), .A2(new_n880), .A3(new_n910), .ZN(new_n911));
  AOI21_X1  g0711(.A(new_n906), .B1(new_n907), .B2(new_n911), .ZN(new_n912));
  AND4_X1   g0712(.A1(new_n906), .A2(new_n438), .A3(new_n881), .A4(new_n454), .ZN(new_n913));
  OAI211_X1 g0713(.A(KEYINPUT38), .B(new_n905), .C1(new_n912), .C2(new_n913), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n893), .A2(new_n914), .ZN(new_n915));
  OAI211_X1 g0715(.A(new_n518), .B(new_n696), .C1(new_n658), .C2(new_n510), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n518), .A2(new_n696), .ZN(new_n917));
  AOI21_X1  g0717(.A(new_n320), .B1(new_n654), .B2(new_n655), .ZN(new_n918));
  NOR3_X1   g0718(.A1(new_n918), .A2(new_n497), .A3(new_n508), .ZN(new_n919));
  OAI211_X1 g0719(.A(new_n523), .B(new_n917), .C1(new_n919), .C2(new_n521), .ZN(new_n920));
  AOI21_X1  g0720(.A(new_n847), .B1(new_n916), .B2(new_n920), .ZN(new_n921));
  INV_X1    g0721(.A(new_n744), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n922), .A2(new_n742), .ZN(new_n923));
  OAI211_X1 g0723(.A(KEYINPUT31), .B(new_n696), .C1(new_n923), .C2(new_n748), .ZN(new_n924));
  NAND3_X1  g0724(.A1(new_n732), .A2(new_n750), .A3(new_n924), .ZN(new_n925));
  AND2_X1   g0725(.A1(new_n921), .A2(new_n925), .ZN(new_n926));
  AND3_X1   g0726(.A1(new_n915), .A2(new_n926), .A3(KEYINPUT40), .ZN(new_n927));
  INV_X1    g0727(.A(KEYINPUT38), .ZN(new_n928));
  NAND3_X1  g0728(.A1(new_n909), .A2(new_n413), .A3(new_n910), .ZN(new_n929));
  NAND3_X1  g0729(.A1(new_n911), .A2(new_n929), .A3(new_n454), .ZN(new_n930));
  AOI21_X1  g0730(.A(new_n913), .B1(new_n930), .B2(KEYINPUT37), .ZN(new_n931));
  NOR2_X1   g0731(.A1(new_n458), .A2(new_n911), .ZN(new_n932));
  OAI21_X1  g0732(.A(new_n928), .B1(new_n931), .B2(new_n932), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n914), .A2(new_n933), .ZN(new_n934));
  AOI21_X1  g0734(.A(KEYINPUT40), .B1(new_n926), .B2(new_n934), .ZN(new_n935));
  NOR2_X1   g0735(.A1(new_n927), .A2(new_n935), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n528), .A2(new_n925), .ZN(new_n937));
  XNOR2_X1  g0737(.A(new_n936), .B(new_n937), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n938), .A2(G330), .ZN(new_n939));
  INV_X1    g0739(.A(KEYINPUT39), .ZN(new_n940));
  NOR3_X1   g0740(.A1(new_n931), .A2(new_n932), .A3(new_n928), .ZN(new_n941));
  NAND2_X1  g0741(.A1(new_n885), .A2(new_n890), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n942), .A2(KEYINPUT103), .ZN(new_n943));
  NAND3_X1  g0743(.A1(new_n885), .A2(new_n886), .A3(new_n890), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n943), .A2(new_n944), .ZN(new_n945));
  OAI21_X1  g0745(.A(new_n940), .B1(new_n941), .B2(new_n945), .ZN(new_n946));
  NAND3_X1  g0746(.A1(new_n510), .A2(new_n518), .A3(new_n697), .ZN(new_n947));
  INV_X1    g0747(.A(new_n947), .ZN(new_n948));
  NAND3_X1  g0748(.A1(new_n914), .A2(new_n933), .A3(KEYINPUT39), .ZN(new_n949));
  NAND3_X1  g0749(.A1(new_n946), .A2(new_n948), .A3(new_n949), .ZN(new_n950));
  AND2_X1   g0750(.A1(new_n916), .A2(new_n920), .ZN(new_n951));
  NAND3_X1  g0751(.A1(new_n840), .A2(new_n697), .A3(new_n841), .ZN(new_n952));
  AOI21_X1  g0752(.A(new_n951), .B1(new_n843), .B2(new_n952), .ZN(new_n953));
  AOI22_X1  g0753(.A1(new_n953), .A2(new_n934), .B1(new_n653), .B2(new_n694), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n950), .A2(new_n954), .ZN(new_n955));
  XNOR2_X1  g0755(.A(new_n939), .B(new_n955), .ZN(new_n956));
  OR2_X1    g0756(.A1(new_n480), .A2(new_n527), .ZN(new_n957));
  AOI21_X1  g0757(.A(new_n957), .B1(new_n728), .B2(new_n730), .ZN(new_n958));
  NOR2_X1   g0758(.A1(new_n958), .A2(new_n664), .ZN(new_n959));
  XNOR2_X1  g0759(.A(new_n956), .B(new_n959), .ZN(new_n960));
  OAI21_X1  g0760(.A(new_n960), .B1(new_n208), .B2(new_n763), .ZN(new_n961));
  AOI21_X1  g0761(.A(new_n251), .B1(new_n587), .B2(KEYINPUT35), .ZN(new_n962));
  OAI211_X1 g0762(.A(new_n962), .B(new_n235), .C1(KEYINPUT35), .C2(new_n587), .ZN(new_n963));
  XNOR2_X1  g0763(.A(new_n963), .B(KEYINPUT36), .ZN(new_n964));
  OAI21_X1  g0764(.A(G77), .B1(new_n228), .B2(new_n415), .ZN(new_n965));
  OAI22_X1  g0765(.A1(new_n965), .A2(new_n236), .B1(G50), .B2(new_n415), .ZN(new_n966));
  NAND3_X1  g0766(.A1(new_n966), .A2(G1), .A3(new_n271), .ZN(new_n967));
  NAND3_X1  g0767(.A1(new_n961), .A2(new_n964), .A3(new_n967), .ZN(new_n968));
  XOR2_X1   g0768(.A(new_n968), .B(KEYINPUT104), .Z(G367));
  NOR2_X1   g0769(.A1(new_n677), .A2(new_n697), .ZN(new_n970));
  NAND3_X1  g0770(.A1(new_n601), .A2(new_n603), .A3(new_n696), .ZN(new_n971));
  AOI21_X1  g0771(.A(new_n970), .B1(new_n722), .B2(new_n971), .ZN(new_n972));
  XOR2_X1   g0772(.A(KEYINPUT105), .B(KEYINPUT42), .Z(new_n973));
  INV_X1    g0773(.A(new_n973), .ZN(new_n974));
  OR3_X1    g0774(.A1(new_n708), .A2(new_n972), .A3(new_n974), .ZN(new_n975));
  OAI21_X1  g0775(.A(new_n974), .B1(new_n708), .B2(new_n972), .ZN(new_n976));
  INV_X1    g0776(.A(new_n972), .ZN(new_n977));
  AOI21_X1  g0777(.A(new_n592), .B1(new_n977), .B2(new_n702), .ZN(new_n978));
  OAI211_X1 g0778(.A(new_n975), .B(new_n976), .C1(new_n696), .C2(new_n978), .ZN(new_n979));
  INV_X1    g0779(.A(KEYINPUT106), .ZN(new_n980));
  NAND2_X1  g0780(.A1(new_n639), .A2(new_n641), .ZN(new_n981));
  NAND2_X1  g0781(.A1(new_n981), .A2(new_n696), .ZN(new_n982));
  NAND2_X1  g0782(.A1(new_n643), .A2(new_n982), .ZN(new_n983));
  OAI21_X1  g0783(.A(new_n983), .B1(new_n637), .B2(new_n982), .ZN(new_n984));
  NAND2_X1  g0784(.A1(new_n984), .A2(KEYINPUT43), .ZN(new_n985));
  NAND3_X1  g0785(.A1(new_n979), .A2(new_n980), .A3(new_n985), .ZN(new_n986));
  INV_X1    g0786(.A(new_n986), .ZN(new_n987));
  AOI21_X1  g0787(.A(new_n980), .B1(new_n979), .B2(new_n985), .ZN(new_n988));
  OAI22_X1  g0788(.A1(new_n987), .A2(new_n988), .B1(KEYINPUT43), .B2(new_n984), .ZN(new_n989));
  INV_X1    g0789(.A(new_n988), .ZN(new_n990));
  NOR2_X1   g0790(.A1(new_n984), .A2(KEYINPUT43), .ZN(new_n991));
  NAND3_X1  g0791(.A1(new_n990), .A2(new_n991), .A3(new_n986), .ZN(new_n992));
  NOR2_X1   g0792(.A1(new_n707), .A2(new_n972), .ZN(new_n993));
  AND3_X1   g0793(.A1(new_n989), .A2(new_n992), .A3(new_n993), .ZN(new_n994));
  AOI21_X1  g0794(.A(new_n993), .B1(new_n989), .B2(new_n992), .ZN(new_n995));
  NOR2_X1   g0795(.A1(new_n994), .A2(new_n995), .ZN(new_n996));
  XNOR2_X1  g0796(.A(new_n715), .B(KEYINPUT41), .ZN(new_n997));
  INV_X1    g0797(.A(new_n997), .ZN(new_n998));
  OAI21_X1  g0798(.A(new_n977), .B1(new_n711), .B2(new_n712), .ZN(new_n999));
  XNOR2_X1  g0799(.A(new_n999), .B(KEYINPUT45), .ZN(new_n1000));
  INV_X1    g0800(.A(new_n712), .ZN(new_n1001));
  NAND3_X1  g0801(.A1(new_n1001), .A2(new_n710), .A3(new_n972), .ZN(new_n1002));
  XNOR2_X1  g0802(.A(new_n1002), .B(KEYINPUT44), .ZN(new_n1003));
  OAI21_X1  g0803(.A(new_n706), .B1(new_n1000), .B2(new_n1003), .ZN(new_n1004));
  NAND2_X1  g0804(.A1(new_n685), .A2(new_n697), .ZN(new_n1005));
  NAND2_X1  g0805(.A1(new_n705), .A2(new_n1005), .ZN(new_n1006));
  AND3_X1   g0806(.A1(new_n701), .A2(new_n708), .A3(new_n1006), .ZN(new_n1007));
  AOI21_X1  g0807(.A(new_n701), .B1(new_n708), .B2(new_n1006), .ZN(new_n1008));
  NOR2_X1   g0808(.A1(new_n1007), .A2(new_n1008), .ZN(new_n1009));
  AOI21_X1  g0809(.A(new_n1009), .B1(new_n756), .B2(new_n758), .ZN(new_n1010));
  INV_X1    g0810(.A(KEYINPUT45), .ZN(new_n1011));
  XNOR2_X1  g0811(.A(new_n999), .B(new_n1011), .ZN(new_n1012));
  INV_X1    g0812(.A(KEYINPUT44), .ZN(new_n1013));
  XNOR2_X1  g0813(.A(new_n1002), .B(new_n1013), .ZN(new_n1014));
  NAND3_X1  g0814(.A1(new_n1012), .A2(new_n1014), .A3(new_n707), .ZN(new_n1015));
  NAND3_X1  g0815(.A1(new_n1004), .A2(new_n1010), .A3(new_n1015), .ZN(new_n1016));
  AOI21_X1  g0816(.A(new_n998), .B1(new_n1016), .B2(new_n759), .ZN(new_n1017));
  NAND2_X1  g0817(.A1(new_n764), .A2(G1), .ZN(new_n1018));
  OAI21_X1  g0818(.A(new_n996), .B1(new_n1017), .B2(new_n1018), .ZN(new_n1019));
  NAND2_X1  g0819(.A1(new_n1019), .A2(KEYINPUT107), .ZN(new_n1020));
  INV_X1    g0820(.A(KEYINPUT107), .ZN(new_n1021));
  OAI211_X1 g0821(.A(new_n996), .B(new_n1021), .C1(new_n1017), .C2(new_n1018), .ZN(new_n1022));
  NAND2_X1  g0822(.A1(new_n1020), .A2(new_n1022), .ZN(new_n1023));
  NOR2_X1   g0823(.A1(new_n808), .A2(new_n218), .ZN(new_n1024));
  NAND2_X1  g0824(.A1(new_n795), .A2(G116), .ZN(new_n1025));
  INV_X1    g0825(.A(KEYINPUT46), .ZN(new_n1026));
  AOI22_X1  g0826(.A1(new_n1025), .A2(new_n1026), .B1(G311), .B2(new_n790), .ZN(new_n1027));
  OAI211_X1 g0827(.A(new_n1027), .B(new_n419), .C1(new_n249), .C2(new_n803), .ZN(new_n1028));
  AOI21_X1  g0828(.A(new_n1028), .B1(G303), .B2(new_n786), .ZN(new_n1029));
  OAI21_X1  g0829(.A(new_n1029), .B1(new_n1026), .B2(new_n1025), .ZN(new_n1030));
  AOI211_X1 g0830(.A(new_n1024), .B(new_n1030), .C1(G294), .C2(new_n798), .ZN(new_n1031));
  XNOR2_X1  g0831(.A(KEYINPUT108), .B(G317), .ZN(new_n1032));
  INV_X1    g0832(.A(new_n1032), .ZN(new_n1033));
  OAI221_X1 g0833(.A(new_n1031), .B1(new_n806), .B2(new_n824), .C1(new_n873), .C2(new_n1033), .ZN(new_n1034));
  NOR2_X1   g0834(.A1(new_n824), .A2(new_n202), .ZN(new_n1035));
  INV_X1    g0835(.A(G159), .ZN(new_n1036));
  OAI22_X1  g0836(.A1(new_n808), .A2(new_n225), .B1(new_n1036), .B2(new_n799), .ZN(new_n1037));
  NOR2_X1   g0837(.A1(new_n821), .A2(new_n415), .ZN(new_n1038));
  OAI21_X1  g0838(.A(new_n341), .B1(new_n796), .B2(new_n228), .ZN(new_n1039));
  NOR3_X1   g0839(.A1(new_n1037), .A2(new_n1038), .A3(new_n1039), .ZN(new_n1040));
  NAND2_X1  g0840(.A1(new_n784), .A2(G137), .ZN(new_n1041));
  AOI22_X1  g0841(.A1(new_n790), .A2(G143), .B1(G150), .B2(new_n786), .ZN(new_n1042));
  NAND3_X1  g0842(.A1(new_n1040), .A2(new_n1041), .A3(new_n1042), .ZN(new_n1043));
  OAI21_X1  g0843(.A(new_n1034), .B1(new_n1035), .B2(new_n1043), .ZN(new_n1044));
  XNOR2_X1  g0844(.A(new_n1044), .B(KEYINPUT47), .ZN(new_n1045));
  NAND2_X1  g0845(.A1(new_n1045), .A2(new_n769), .ZN(new_n1046));
  OR2_X1    g0846(.A1(new_n984), .A2(new_n835), .ZN(new_n1047));
  OAI221_X1 g0847(.A(new_n771), .B1(new_n212), .B2(new_n471), .C1(new_n241), .C2(new_n774), .ZN(new_n1048));
  NAND4_X1  g0848(.A1(new_n1046), .A2(new_n766), .A3(new_n1047), .A4(new_n1048), .ZN(new_n1049));
  NAND2_X1  g0849(.A1(new_n1023), .A2(new_n1049), .ZN(G387));
  INV_X1    g0850(.A(new_n1009), .ZN(new_n1051));
  NAND2_X1  g0851(.A1(new_n759), .A2(new_n1051), .ZN(new_n1052));
  NAND3_X1  g0852(.A1(new_n756), .A2(new_n758), .A3(new_n1009), .ZN(new_n1053));
  NAND3_X1  g0853(.A1(new_n1052), .A2(new_n1053), .A3(new_n715), .ZN(new_n1054));
  NOR2_X1   g0854(.A1(new_n362), .A2(G50), .ZN(new_n1055));
  XNOR2_X1  g0855(.A(new_n1055), .B(KEYINPUT50), .ZN(new_n1056));
  NAND2_X1  g0856(.A1(G68), .A2(G77), .ZN(new_n1057));
  NAND4_X1  g0857(.A1(new_n1056), .A2(new_n718), .A3(new_n297), .A4(new_n1057), .ZN(new_n1058));
  AOI21_X1  g0858(.A(new_n774), .B1(new_n246), .B2(G45), .ZN(new_n1059));
  NOR3_X1   g0859(.A1(new_n718), .A2(new_n714), .A3(new_n419), .ZN(new_n1060));
  OAI21_X1  g0860(.A(new_n1058), .B1(new_n1059), .B2(new_n1060), .ZN(new_n1061));
  NAND2_X1  g0861(.A1(new_n714), .A2(new_n249), .ZN(new_n1062));
  AOI21_X1  g0862(.A(new_n772), .B1(new_n1061), .B2(new_n1062), .ZN(new_n1063));
  NOR2_X1   g0863(.A1(new_n821), .A2(new_n471), .ZN(new_n1064));
  AOI21_X1  g0864(.A(new_n1064), .B1(new_n378), .B2(new_n798), .ZN(new_n1065));
  OAI21_X1  g0865(.A(new_n1065), .B1(new_n415), .B2(new_n824), .ZN(new_n1066));
  AOI22_X1  g0866(.A1(new_n784), .A2(G150), .B1(G159), .B2(new_n790), .ZN(new_n1067));
  OAI221_X1 g0867(.A(new_n1067), .B1(new_n202), .B2(new_n825), .C1(new_n225), .C2(new_n796), .ZN(new_n1068));
  OR4_X1    g0868(.A1(new_n419), .A2(new_n1066), .A3(new_n1024), .A4(new_n1068), .ZN(new_n1069));
  AOI22_X1  g0869(.A1(G303), .A2(new_n810), .B1(new_n798), .B2(G311), .ZN(new_n1070));
  OAI21_X1  g0870(.A(new_n1070), .B1(new_n825), .B2(new_n1033), .ZN(new_n1071));
  AOI21_X1  g0871(.A(new_n1071), .B1(G322), .B2(new_n790), .ZN(new_n1072));
  XOR2_X1   g0872(.A(new_n1072), .B(KEYINPUT48), .Z(new_n1073));
  OAI221_X1 g0873(.A(new_n1073), .B1(new_n806), .B2(new_n803), .C1(new_n550), .C2(new_n796), .ZN(new_n1074));
  XOR2_X1   g0874(.A(new_n1074), .B(KEYINPUT49), .Z(new_n1075));
  AOI21_X1  g0875(.A(new_n341), .B1(new_n784), .B2(G326), .ZN(new_n1076));
  OAI21_X1  g0876(.A(new_n1076), .B1(new_n251), .B2(new_n808), .ZN(new_n1077));
  OAI21_X1  g0877(.A(new_n1069), .B1(new_n1075), .B2(new_n1077), .ZN(new_n1078));
  AOI21_X1  g0878(.A(new_n1063), .B1(new_n1078), .B2(new_n769), .ZN(new_n1079));
  INV_X1    g0879(.A(new_n705), .ZN(new_n1080));
  OAI211_X1 g0880(.A(new_n1079), .B(new_n766), .C1(new_n1080), .C2(new_n835), .ZN(new_n1081));
  XNOR2_X1  g0881(.A(new_n1081), .B(KEYINPUT109), .ZN(new_n1082));
  NAND2_X1  g0882(.A1(new_n1051), .A2(new_n1018), .ZN(new_n1083));
  NAND3_X1  g0883(.A1(new_n1054), .A2(new_n1082), .A3(new_n1083), .ZN(new_n1084));
  XNOR2_X1  g0884(.A(new_n1084), .B(KEYINPUT110), .ZN(G393));
  NAND2_X1  g0885(.A1(new_n1004), .A2(new_n1015), .ZN(new_n1086));
  NAND2_X1  g0886(.A1(new_n1086), .A2(new_n1052), .ZN(new_n1087));
  NAND3_X1  g0887(.A1(new_n1087), .A2(new_n715), .A3(new_n1016), .ZN(new_n1088));
  NAND3_X1  g0888(.A1(new_n1004), .A2(new_n1018), .A3(new_n1015), .ZN(new_n1089));
  AOI22_X1  g0889(.A1(new_n790), .A2(G150), .B1(G159), .B2(new_n786), .ZN(new_n1090));
  XNOR2_X1  g0890(.A(new_n1090), .B(KEYINPUT51), .ZN(new_n1091));
  OAI21_X1  g0891(.A(new_n341), .B1(new_n796), .B2(new_n415), .ZN(new_n1092));
  NOR2_X1   g0892(.A1(new_n1091), .A2(new_n1092), .ZN(new_n1093));
  OAI21_X1  g0893(.A(new_n1093), .B1(new_n216), .B2(new_n808), .ZN(new_n1094));
  NOR2_X1   g0894(.A1(new_n821), .A2(new_n225), .ZN(new_n1095));
  AOI21_X1  g0895(.A(new_n1095), .B1(G50), .B2(new_n798), .ZN(new_n1096));
  OAI21_X1  g0896(.A(new_n1096), .B1(new_n362), .B2(new_n824), .ZN(new_n1097));
  XOR2_X1   g0897(.A(new_n1097), .B(KEYINPUT111), .Z(new_n1098));
  AOI211_X1 g0898(.A(new_n1094), .B(new_n1098), .C1(G143), .C2(new_n784), .ZN(new_n1099));
  AOI22_X1  g0899(.A1(new_n790), .A2(G317), .B1(G311), .B2(new_n786), .ZN(new_n1100));
  XNOR2_X1  g0900(.A(new_n1100), .B(KEYINPUT52), .ZN(new_n1101));
  AOI211_X1 g0901(.A(new_n341), .B(new_n1101), .C1(G322), .C2(new_n784), .ZN(new_n1102));
  OAI22_X1  g0902(.A1(new_n824), .A2(new_n550), .B1(new_n799), .B2(new_n293), .ZN(new_n1103));
  AOI211_X1 g0903(.A(new_n1103), .B(new_n830), .C1(G283), .C2(new_n795), .ZN(new_n1104));
  OAI211_X1 g0904(.A(new_n1102), .B(new_n1104), .C1(new_n251), .C2(new_n803), .ZN(new_n1105));
  XOR2_X1   g0905(.A(new_n1105), .B(KEYINPUT112), .Z(new_n1106));
  OAI21_X1  g0906(.A(new_n769), .B1(new_n1099), .B2(new_n1106), .ZN(new_n1107));
  INV_X1    g0907(.A(new_n252), .ZN(new_n1108));
  OAI221_X1 g0908(.A(new_n771), .B1(new_n218), .B2(new_n212), .C1(new_n1108), .C2(new_n774), .ZN(new_n1109));
  AOI21_X1  g0909(.A(new_n765), .B1(new_n972), .B2(new_n770), .ZN(new_n1110));
  NAND3_X1  g0910(.A1(new_n1107), .A2(new_n1109), .A3(new_n1110), .ZN(new_n1111));
  NAND3_X1  g0911(.A1(new_n1088), .A2(new_n1089), .A3(new_n1111), .ZN(G390));
  NAND2_X1  g0912(.A1(new_n843), .A2(new_n952), .ZN(new_n1113));
  NAND2_X1  g0913(.A1(new_n916), .A2(new_n920), .ZN(new_n1114));
  NAND2_X1  g0914(.A1(new_n1113), .A2(new_n1114), .ZN(new_n1115));
  AOI22_X1  g0915(.A1(new_n946), .A2(new_n949), .B1(new_n1115), .B2(new_n947), .ZN(new_n1116));
  INV_X1    g0916(.A(new_n952), .ZN(new_n1117));
  AOI21_X1  g0917(.A(new_n696), .B1(new_n723), .B2(new_n726), .ZN(new_n1118));
  AOI21_X1  g0918(.A(new_n1117), .B1(new_n1118), .B2(new_n842), .ZN(new_n1119));
  OAI21_X1  g0919(.A(new_n947), .B1(new_n1119), .B2(new_n951), .ZN(new_n1120));
  NOR2_X1   g0920(.A1(new_n941), .A2(new_n945), .ZN(new_n1121));
  NOR2_X1   g0921(.A1(new_n1120), .A2(new_n1121), .ZN(new_n1122));
  NAND4_X1  g0922(.A1(new_n753), .A2(G330), .A3(new_n848), .A4(new_n1114), .ZN(new_n1123));
  NOR3_X1   g0923(.A1(new_n1116), .A2(new_n1122), .A3(new_n1123), .ZN(new_n1124));
  NAND4_X1  g0924(.A1(new_n925), .A2(G330), .A3(new_n848), .A4(new_n1114), .ZN(new_n1125));
  INV_X1    g0925(.A(new_n1125), .ZN(new_n1126));
  AND3_X1   g0926(.A1(new_n914), .A2(new_n933), .A3(KEYINPUT39), .ZN(new_n1127));
  AOI21_X1  g0927(.A(KEYINPUT39), .B1(new_n893), .B2(new_n914), .ZN(new_n1128));
  OAI22_X1  g0928(.A1(new_n1127), .A2(new_n1128), .B1(new_n948), .B2(new_n953), .ZN(new_n1129));
  OAI211_X1 g0929(.A(new_n915), .B(new_n947), .C1(new_n951), .C2(new_n1119), .ZN(new_n1130));
  AOI21_X1  g0930(.A(new_n1126), .B1(new_n1129), .B2(new_n1130), .ZN(new_n1131));
  OAI21_X1  g0931(.A(new_n1018), .B1(new_n1124), .B2(new_n1131), .ZN(new_n1132));
  NAND2_X1  g0932(.A1(new_n946), .A2(new_n949), .ZN(new_n1133));
  OAI21_X1  g0933(.A(new_n341), .B1(new_n808), .B2(new_n202), .ZN(new_n1134));
  NAND2_X1  g0934(.A1(new_n795), .A2(G150), .ZN(new_n1135));
  XNOR2_X1  g0935(.A(new_n1135), .B(KEYINPUT53), .ZN(new_n1136));
  AOI211_X1 g0936(.A(new_n1134), .B(new_n1136), .C1(G159), .C2(new_n822), .ZN(new_n1137));
  NAND2_X1  g0937(.A1(new_n798), .A2(G137), .ZN(new_n1138));
  NAND2_X1  g0938(.A1(new_n786), .A2(G132), .ZN(new_n1139));
  XNOR2_X1  g0939(.A(KEYINPUT54), .B(G143), .ZN(new_n1140));
  INV_X1    g0940(.A(G128), .ZN(new_n1141));
  OAI22_X1  g0941(.A1(new_n824), .A2(new_n1140), .B1(new_n789), .B2(new_n1141), .ZN(new_n1142));
  AOI21_X1  g0942(.A(new_n1142), .B1(new_n784), .B2(G125), .ZN(new_n1143));
  NAND4_X1  g0943(.A1(new_n1137), .A2(new_n1138), .A3(new_n1139), .A4(new_n1143), .ZN(new_n1144));
  OAI21_X1  g0944(.A(new_n871), .B1(new_n873), .B2(new_n550), .ZN(new_n1145));
  OAI21_X1  g0945(.A(new_n817), .B1(new_n1145), .B2(KEYINPUT115), .ZN(new_n1146));
  AOI211_X1 g0946(.A(new_n1095), .B(new_n1146), .C1(KEYINPUT115), .C2(new_n1145), .ZN(new_n1147));
  NAND2_X1  g0947(.A1(new_n786), .A2(G116), .ZN(new_n1148));
  AOI22_X1  g0948(.A1(new_n790), .A2(G283), .B1(G97), .B2(new_n810), .ZN(new_n1149));
  NAND4_X1  g0949(.A1(new_n1147), .A2(new_n419), .A3(new_n1148), .A4(new_n1149), .ZN(new_n1150));
  NOR2_X1   g0950(.A1(new_n799), .A2(new_n249), .ZN(new_n1151));
  OAI21_X1  g0951(.A(new_n1144), .B1(new_n1150), .B2(new_n1151), .ZN(new_n1152));
  AOI22_X1  g0952(.A1(new_n1133), .A2(new_n852), .B1(new_n769), .B2(new_n1152), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n855), .A2(new_n362), .ZN(new_n1154));
  NAND3_X1  g0954(.A1(new_n1153), .A2(new_n766), .A3(new_n1154), .ZN(new_n1155));
  INV_X1    g0955(.A(KEYINPUT116), .ZN(new_n1156));
  NAND2_X1  g0956(.A1(new_n1155), .A2(new_n1156), .ZN(new_n1157));
  NAND4_X1  g0957(.A1(new_n1153), .A2(KEYINPUT116), .A3(new_n766), .A4(new_n1154), .ZN(new_n1158));
  NAND3_X1  g0958(.A1(new_n1132), .A2(new_n1157), .A3(new_n1158), .ZN(new_n1159));
  XNOR2_X1  g0959(.A(new_n1159), .B(KEYINPUT117), .ZN(new_n1160));
  OAI21_X1  g0960(.A(new_n1125), .B1(new_n1116), .B2(new_n1122), .ZN(new_n1161));
  AND3_X1   g0961(.A1(new_n528), .A2(G330), .A3(new_n925), .ZN(new_n1162));
  NOR3_X1   g0962(.A1(new_n958), .A2(new_n1162), .A3(new_n664), .ZN(new_n1163));
  NAND3_X1  g0963(.A1(new_n925), .A2(G330), .A3(new_n848), .ZN(new_n1164));
  NAND2_X1  g0964(.A1(new_n1164), .A2(new_n951), .ZN(new_n1165));
  AND3_X1   g0965(.A1(new_n1165), .A2(new_n1119), .A3(new_n1123), .ZN(new_n1166));
  INV_X1    g0966(.A(new_n1113), .ZN(new_n1167));
  NAND3_X1  g0967(.A1(new_n753), .A2(G330), .A3(new_n848), .ZN(new_n1168));
  NAND2_X1  g0968(.A1(new_n1168), .A2(new_n951), .ZN(new_n1169));
  AOI21_X1  g0969(.A(new_n1167), .B1(new_n1169), .B2(new_n1125), .ZN(new_n1170));
  OAI21_X1  g0970(.A(new_n1163), .B1(new_n1166), .B2(new_n1170), .ZN(new_n1171));
  INV_X1    g0971(.A(new_n1123), .ZN(new_n1172));
  NAND3_X1  g0972(.A1(new_n1129), .A2(new_n1130), .A3(new_n1172), .ZN(new_n1173));
  NAND3_X1  g0973(.A1(new_n1161), .A2(new_n1171), .A3(new_n1173), .ZN(new_n1174));
  NAND2_X1  g0974(.A1(new_n1174), .A2(KEYINPUT113), .ZN(new_n1175));
  INV_X1    g0975(.A(KEYINPUT113), .ZN(new_n1176));
  NAND4_X1  g0976(.A1(new_n1161), .A2(new_n1171), .A3(new_n1176), .A4(new_n1173), .ZN(new_n1177));
  NAND2_X1  g0977(.A1(new_n731), .A2(new_n528), .ZN(new_n1178));
  NAND3_X1  g0978(.A1(new_n528), .A2(new_n925), .A3(G330), .ZN(new_n1179));
  NAND3_X1  g0979(.A1(new_n1178), .A2(new_n665), .A3(new_n1179), .ZN(new_n1180));
  INV_X1    g0980(.A(new_n1170), .ZN(new_n1181));
  NAND3_X1  g0981(.A1(new_n1165), .A2(new_n1119), .A3(new_n1123), .ZN(new_n1182));
  AOI21_X1  g0982(.A(new_n1180), .B1(new_n1181), .B2(new_n1182), .ZN(new_n1183));
  OAI21_X1  g0983(.A(new_n1183), .B1(new_n1124), .B2(new_n1131), .ZN(new_n1184));
  NAND4_X1  g0984(.A1(new_n1175), .A2(new_n715), .A3(new_n1177), .A4(new_n1184), .ZN(new_n1185));
  INV_X1    g0985(.A(KEYINPUT114), .ZN(new_n1186));
  AND2_X1   g0986(.A1(new_n1185), .A2(new_n1186), .ZN(new_n1187));
  NOR2_X1   g0987(.A1(new_n1185), .A2(new_n1186), .ZN(new_n1188));
  OAI21_X1  g0988(.A(new_n1160), .B1(new_n1187), .B2(new_n1188), .ZN(G378));
  INV_X1    g0989(.A(new_n1018), .ZN(new_n1190));
  INV_X1    g0990(.A(KEYINPUT119), .ZN(new_n1191));
  XOR2_X1   g0991(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1192));
  OAI21_X1  g0992(.A(new_n1192), .B1(new_n663), .B2(new_n375), .ZN(new_n1193));
  INV_X1    g0993(.A(new_n1192), .ZN(new_n1194));
  NAND2_X1  g0994(.A1(new_n398), .A2(new_n1194), .ZN(new_n1195));
  NAND2_X1  g0995(.A1(new_n1193), .A2(new_n1195), .ZN(new_n1196));
  NOR2_X1   g0996(.A1(new_n394), .A2(new_n694), .ZN(new_n1197));
  INV_X1    g0997(.A(new_n1197), .ZN(new_n1198));
  NAND2_X1  g0998(.A1(new_n1196), .A2(new_n1198), .ZN(new_n1199));
  NAND3_X1  g0999(.A1(new_n1193), .A2(new_n1197), .A3(new_n1195), .ZN(new_n1200));
  NAND2_X1  g1000(.A1(new_n1199), .A2(new_n1200), .ZN(new_n1201));
  INV_X1    g1001(.A(KEYINPUT118), .ZN(new_n1202));
  NAND2_X1  g1002(.A1(new_n1201), .A2(new_n1202), .ZN(new_n1203));
  AND3_X1   g1003(.A1(new_n950), .A2(new_n1203), .A3(new_n954), .ZN(new_n1204));
  AOI21_X1  g1004(.A(new_n1203), .B1(new_n950), .B2(new_n954), .ZN(new_n1205));
  NAND3_X1  g1005(.A1(new_n915), .A2(new_n926), .A3(KEYINPUT40), .ZN(new_n1206));
  AND2_X1   g1006(.A1(new_n926), .A2(new_n934), .ZN(new_n1207));
  OAI211_X1 g1007(.A(new_n1206), .B(G330), .C1(new_n1207), .C2(KEYINPUT40), .ZN(new_n1208));
  NOR3_X1   g1008(.A1(new_n1204), .A2(new_n1205), .A3(new_n1208), .ZN(new_n1209));
  INV_X1    g1009(.A(G330), .ZN(new_n1210));
  NOR3_X1   g1010(.A1(new_n927), .A2(new_n935), .A3(new_n1210), .ZN(new_n1211));
  INV_X1    g1011(.A(new_n1203), .ZN(new_n1212));
  NAND2_X1  g1012(.A1(new_n955), .A2(new_n1212), .ZN(new_n1213));
  NAND3_X1  g1013(.A1(new_n950), .A2(new_n1203), .A3(new_n954), .ZN(new_n1214));
  AOI21_X1  g1014(.A(new_n1211), .B1(new_n1213), .B2(new_n1214), .ZN(new_n1215));
  OAI21_X1  g1015(.A(new_n1191), .B1(new_n1209), .B2(new_n1215), .ZN(new_n1216));
  OAI21_X1  g1016(.A(new_n1208), .B1(new_n1204), .B2(new_n1205), .ZN(new_n1217));
  NAND3_X1  g1017(.A1(new_n1213), .A2(new_n1211), .A3(new_n1214), .ZN(new_n1218));
  NAND3_X1  g1018(.A1(new_n1217), .A2(new_n1218), .A3(KEYINPUT119), .ZN(new_n1219));
  AOI21_X1  g1019(.A(new_n1190), .B1(new_n1216), .B2(new_n1219), .ZN(new_n1220));
  NAND2_X1  g1020(.A1(new_n1201), .A2(new_n852), .ZN(new_n1221));
  AOI22_X1  g1021(.A1(new_n784), .A2(G283), .B1(new_n807), .B2(G58), .ZN(new_n1222));
  OAI21_X1  g1022(.A(new_n1222), .B1(new_n249), .B2(new_n825), .ZN(new_n1223));
  AOI211_X1 g1023(.A(new_n1038), .B(new_n1223), .C1(new_n470), .C2(new_n810), .ZN(new_n1224));
  OAI21_X1  g1024(.A(new_n419), .B1(new_n789), .B2(new_n251), .ZN(new_n1225));
  AOI211_X1 g1025(.A(G41), .B(new_n1225), .C1(G77), .C2(new_n795), .ZN(new_n1226));
  OAI211_X1 g1026(.A(new_n1224), .B(new_n1226), .C1(new_n218), .C2(new_n799), .ZN(new_n1227));
  XOR2_X1   g1027(.A(new_n1227), .B(KEYINPUT58), .Z(new_n1228));
  OAI21_X1  g1028(.A(new_n202), .B1(new_n286), .B2(G41), .ZN(new_n1229));
  AOI22_X1  g1029(.A1(new_n822), .A2(G150), .B1(G128), .B2(new_n786), .ZN(new_n1230));
  AOI22_X1  g1030(.A1(new_n790), .A2(G125), .B1(G132), .B2(new_n798), .ZN(new_n1231));
  OAI211_X1 g1031(.A(new_n1230), .B(new_n1231), .C1(new_n796), .C2(new_n1140), .ZN(new_n1232));
  AOI21_X1  g1032(.A(new_n1232), .B1(G137), .B2(new_n810), .ZN(new_n1233));
  INV_X1    g1033(.A(KEYINPUT59), .ZN(new_n1234));
  AOI21_X1  g1034(.A(G33), .B1(new_n1233), .B2(new_n1234), .ZN(new_n1235));
  AOI21_X1  g1035(.A(G41), .B1(new_n784), .B2(G124), .ZN(new_n1236));
  OAI211_X1 g1036(.A(new_n1235), .B(new_n1236), .C1(new_n1036), .C2(new_n808), .ZN(new_n1237));
  NOR2_X1   g1037(.A1(new_n1233), .A2(new_n1234), .ZN(new_n1238));
  OAI21_X1  g1038(.A(new_n1229), .B1(new_n1237), .B2(new_n1238), .ZN(new_n1239));
  OAI21_X1  g1039(.A(new_n769), .B1(new_n1228), .B2(new_n1239), .ZN(new_n1240));
  NAND2_X1  g1040(.A1(new_n855), .A2(new_n202), .ZN(new_n1241));
  NAND4_X1  g1041(.A1(new_n1221), .A2(new_n766), .A3(new_n1240), .A4(new_n1241), .ZN(new_n1242));
  INV_X1    g1042(.A(new_n1242), .ZN(new_n1243));
  OAI21_X1  g1043(.A(KEYINPUT120), .B1(new_n1220), .B2(new_n1243), .ZN(new_n1244));
  AND3_X1   g1044(.A1(new_n1217), .A2(new_n1218), .A3(KEYINPUT119), .ZN(new_n1245));
  AOI21_X1  g1045(.A(KEYINPUT119), .B1(new_n1217), .B2(new_n1218), .ZN(new_n1246));
  OAI21_X1  g1046(.A(new_n1018), .B1(new_n1245), .B2(new_n1246), .ZN(new_n1247));
  INV_X1    g1047(.A(KEYINPUT120), .ZN(new_n1248));
  NAND3_X1  g1048(.A1(new_n1247), .A2(new_n1248), .A3(new_n1242), .ZN(new_n1249));
  NAND2_X1  g1049(.A1(new_n1244), .A2(new_n1249), .ZN(new_n1250));
  NAND2_X1  g1050(.A1(new_n1217), .A2(new_n1218), .ZN(new_n1251));
  AOI21_X1  g1051(.A(new_n1171), .B1(new_n1161), .B2(new_n1173), .ZN(new_n1252));
  INV_X1    g1052(.A(KEYINPUT121), .ZN(new_n1253));
  NOR3_X1   g1053(.A1(new_n1252), .A2(new_n1253), .A3(new_n1180), .ZN(new_n1254));
  AOI21_X1  g1054(.A(KEYINPUT121), .B1(new_n1184), .B2(new_n1163), .ZN(new_n1255));
  OAI211_X1 g1055(.A(KEYINPUT57), .B(new_n1251), .C1(new_n1254), .C2(new_n1255), .ZN(new_n1256));
  OAI21_X1  g1056(.A(new_n1253), .B1(new_n1252), .B2(new_n1180), .ZN(new_n1257));
  NAND3_X1  g1057(.A1(new_n1184), .A2(KEYINPUT121), .A3(new_n1163), .ZN(new_n1258));
  AOI22_X1  g1058(.A1(new_n1219), .A2(new_n1216), .B1(new_n1257), .B2(new_n1258), .ZN(new_n1259));
  OAI211_X1 g1059(.A(new_n715), .B(new_n1256), .C1(new_n1259), .C2(KEYINPUT57), .ZN(new_n1260));
  NAND2_X1  g1060(.A1(new_n1250), .A2(new_n1260), .ZN(new_n1261));
  INV_X1    g1061(.A(KEYINPUT122), .ZN(new_n1262));
  NOR2_X1   g1062(.A1(new_n1261), .A2(new_n1262), .ZN(new_n1263));
  INV_X1    g1063(.A(new_n1263), .ZN(new_n1264));
  AOI21_X1  g1064(.A(KEYINPUT122), .B1(new_n1250), .B2(new_n1260), .ZN(new_n1265));
  INV_X1    g1065(.A(new_n1265), .ZN(new_n1266));
  NAND2_X1  g1066(.A1(new_n1264), .A2(new_n1266), .ZN(G375));
  NOR2_X1   g1067(.A1(new_n1166), .A2(new_n1170), .ZN(new_n1268));
  NAND2_X1  g1068(.A1(new_n1268), .A2(new_n1180), .ZN(new_n1269));
  NAND3_X1  g1069(.A1(new_n1269), .A2(new_n997), .A3(new_n1171), .ZN(new_n1270));
  NAND2_X1  g1070(.A1(new_n951), .A2(new_n852), .ZN(new_n1271));
  NOR2_X1   g1071(.A1(new_n799), .A2(new_n1140), .ZN(new_n1272));
  OAI22_X1  g1072(.A1(new_n796), .A2(new_n1036), .B1(new_n789), .B2(new_n874), .ZN(new_n1273));
  AOI21_X1  g1073(.A(new_n1273), .B1(G58), .B2(new_n807), .ZN(new_n1274));
  NAND2_X1  g1074(.A1(new_n784), .A2(G128), .ZN(new_n1275));
  NAND2_X1  g1075(.A1(new_n822), .A2(G50), .ZN(new_n1276));
  AOI21_X1  g1076(.A(new_n419), .B1(G150), .B2(new_n810), .ZN(new_n1277));
  NAND4_X1  g1077(.A1(new_n1274), .A2(new_n1275), .A3(new_n1276), .A4(new_n1277), .ZN(new_n1278));
  AOI211_X1 g1078(.A(new_n1272), .B(new_n1278), .C1(G137), .C2(new_n786), .ZN(new_n1279));
  AOI21_X1  g1079(.A(new_n1064), .B1(G283), .B2(new_n786), .ZN(new_n1280));
  AOI22_X1  g1080(.A1(new_n807), .A2(G77), .B1(G97), .B2(new_n795), .ZN(new_n1281));
  OAI211_X1 g1081(.A(new_n1280), .B(new_n1281), .C1(new_n293), .C2(new_n873), .ZN(new_n1282));
  NOR2_X1   g1082(.A1(new_n799), .A2(new_n251), .ZN(new_n1283));
  NOR2_X1   g1083(.A1(new_n824), .A2(new_n249), .ZN(new_n1284));
  OAI21_X1  g1084(.A(new_n419), .B1(new_n789), .B2(new_n550), .ZN(new_n1285));
  NOR4_X1   g1085(.A1(new_n1282), .A2(new_n1283), .A3(new_n1284), .A4(new_n1285), .ZN(new_n1286));
  OAI21_X1  g1086(.A(new_n769), .B1(new_n1279), .B2(new_n1286), .ZN(new_n1287));
  AOI21_X1  g1087(.A(new_n765), .B1(new_n855), .B2(new_n415), .ZN(new_n1288));
  XOR2_X1   g1088(.A(new_n1288), .B(KEYINPUT124), .Z(new_n1289));
  AND3_X1   g1089(.A1(new_n1271), .A2(new_n1287), .A3(new_n1289), .ZN(new_n1290));
  INV_X1    g1090(.A(new_n1268), .ZN(new_n1291));
  XOR2_X1   g1091(.A(new_n1018), .B(KEYINPUT123), .Z(new_n1292));
  AOI21_X1  g1092(.A(new_n1290), .B1(new_n1291), .B2(new_n1292), .ZN(new_n1293));
  NAND2_X1  g1093(.A1(new_n1270), .A2(new_n1293), .ZN(G381));
  AND2_X1   g1094(.A1(new_n1160), .A2(new_n1185), .ZN(new_n1295));
  NAND3_X1  g1095(.A1(new_n1264), .A2(new_n1266), .A3(new_n1295), .ZN(new_n1296));
  INV_X1    g1096(.A(G390), .ZN(new_n1297));
  AND3_X1   g1097(.A1(new_n1023), .A2(new_n1049), .A3(new_n1297), .ZN(new_n1298));
  NOR2_X1   g1098(.A1(G381), .A2(G384), .ZN(new_n1299));
  NOR2_X1   g1099(.A1(G393), .A2(G396), .ZN(new_n1300));
  NAND3_X1  g1100(.A1(new_n1298), .A2(new_n1299), .A3(new_n1300), .ZN(new_n1301));
  OR2_X1    g1101(.A1(new_n1296), .A2(new_n1301), .ZN(G407));
  AND2_X1   g1102(.A1(new_n1301), .A2(G343), .ZN(new_n1303));
  OAI21_X1  g1103(.A(G213), .B1(new_n1296), .B2(new_n1303), .ZN(G409));
  NOR2_X1   g1104(.A1(new_n691), .A2(G343), .ZN(new_n1305));
  NAND3_X1  g1105(.A1(new_n1250), .A2(G378), .A3(new_n1260), .ZN(new_n1306));
  NAND2_X1  g1106(.A1(new_n1257), .A2(new_n1258), .ZN(new_n1307));
  OAI211_X1 g1107(.A(new_n1307), .B(new_n997), .C1(new_n1245), .C2(new_n1246), .ZN(new_n1308));
  NAND2_X1  g1108(.A1(new_n1251), .A2(new_n1292), .ZN(new_n1309));
  NAND3_X1  g1109(.A1(new_n1308), .A2(new_n1242), .A3(new_n1309), .ZN(new_n1310));
  NAND2_X1  g1110(.A1(new_n1295), .A2(new_n1310), .ZN(new_n1311));
  AOI21_X1  g1111(.A(new_n1305), .B1(new_n1306), .B2(new_n1311), .ZN(new_n1312));
  INV_X1    g1112(.A(KEYINPUT60), .ZN(new_n1313));
  OAI211_X1 g1113(.A(new_n715), .B(new_n1171), .C1(new_n1269), .C2(new_n1313), .ZN(new_n1314));
  AOI21_X1  g1114(.A(KEYINPUT60), .B1(new_n1268), .B2(new_n1180), .ZN(new_n1315));
  OAI21_X1  g1115(.A(new_n1293), .B1(new_n1314), .B2(new_n1315), .ZN(new_n1316));
  NAND3_X1  g1116(.A1(new_n1316), .A2(new_n851), .A3(new_n878), .ZN(new_n1317));
  OAI211_X1 g1117(.A(G384), .B(new_n1293), .C1(new_n1314), .C2(new_n1315), .ZN(new_n1318));
  NAND2_X1  g1118(.A1(new_n1317), .A2(new_n1318), .ZN(new_n1319));
  INV_X1    g1119(.A(KEYINPUT63), .ZN(new_n1320));
  NOR2_X1   g1120(.A1(new_n1319), .A2(new_n1320), .ZN(new_n1321));
  AOI21_X1  g1121(.A(KEYINPUT61), .B1(new_n1312), .B2(new_n1321), .ZN(new_n1322));
  AOI21_X1  g1122(.A(new_n1297), .B1(new_n1023), .B2(new_n1049), .ZN(new_n1323));
  AND2_X1   g1123(.A1(G393), .A2(G396), .ZN(new_n1324));
  OAI22_X1  g1124(.A1(new_n1298), .A2(new_n1323), .B1(new_n1300), .B2(new_n1324), .ZN(new_n1325));
  NAND2_X1  g1125(.A1(G387), .A2(G390), .ZN(new_n1326));
  NAND3_X1  g1126(.A1(new_n1023), .A2(new_n1049), .A3(new_n1297), .ZN(new_n1327));
  XNOR2_X1  g1127(.A(G393), .B(new_n837), .ZN(new_n1328));
  NAND3_X1  g1128(.A1(new_n1326), .A2(new_n1327), .A3(new_n1328), .ZN(new_n1329));
  NAND2_X1  g1129(.A1(new_n1325), .A2(new_n1329), .ZN(new_n1330));
  NAND2_X1  g1130(.A1(new_n1306), .A2(new_n1311), .ZN(new_n1331));
  INV_X1    g1131(.A(KEYINPUT125), .ZN(new_n1332));
  NAND2_X1  g1132(.A1(new_n1331), .A2(new_n1332), .ZN(new_n1333));
  INV_X1    g1133(.A(new_n1305), .ZN(new_n1334));
  NAND3_X1  g1134(.A1(new_n1306), .A2(new_n1311), .A3(KEYINPUT125), .ZN(new_n1335));
  NAND3_X1  g1135(.A1(new_n1333), .A2(new_n1334), .A3(new_n1335), .ZN(new_n1336));
  NAND2_X1  g1136(.A1(new_n1305), .A2(G2897), .ZN(new_n1337));
  XOR2_X1   g1137(.A(new_n1319), .B(new_n1337), .Z(new_n1338));
  INV_X1    g1138(.A(new_n1338), .ZN(new_n1339));
  AOI21_X1  g1139(.A(new_n1320), .B1(new_n1336), .B2(new_n1339), .ZN(new_n1340));
  INV_X1    g1140(.A(new_n1319), .ZN(new_n1341));
  NAND4_X1  g1141(.A1(new_n1333), .A2(new_n1334), .A3(new_n1341), .A4(new_n1335), .ZN(new_n1342));
  INV_X1    g1142(.A(new_n1342), .ZN(new_n1343));
  OAI211_X1 g1143(.A(new_n1322), .B(new_n1330), .C1(new_n1340), .C2(new_n1343), .ZN(new_n1344));
  NOR2_X1   g1144(.A1(new_n1330), .A2(KEYINPUT126), .ZN(new_n1345));
  INV_X1    g1145(.A(KEYINPUT126), .ZN(new_n1346));
  AOI21_X1  g1146(.A(new_n1346), .B1(new_n1325), .B2(new_n1329), .ZN(new_n1347));
  NOR2_X1   g1147(.A1(new_n1345), .A2(new_n1347), .ZN(new_n1348));
  INV_X1    g1148(.A(KEYINPUT62), .ZN(new_n1349));
  NOR2_X1   g1149(.A1(new_n1319), .A2(new_n1349), .ZN(new_n1350));
  AND2_X1   g1150(.A1(new_n1312), .A2(new_n1350), .ZN(new_n1351));
  AOI21_X1  g1151(.A(new_n1351), .B1(new_n1342), .B2(new_n1349), .ZN(new_n1352));
  INV_X1    g1152(.A(KEYINPUT61), .ZN(new_n1353));
  OAI21_X1  g1153(.A(new_n1353), .B1(new_n1312), .B2(new_n1338), .ZN(new_n1354));
  OAI21_X1  g1154(.A(new_n1348), .B1(new_n1352), .B2(new_n1354), .ZN(new_n1355));
  NAND2_X1  g1155(.A1(new_n1344), .A2(new_n1355), .ZN(G405));
  OAI21_X1  g1156(.A(new_n1295), .B1(new_n1263), .B2(new_n1265), .ZN(new_n1357));
  INV_X1    g1157(.A(KEYINPUT127), .ZN(new_n1358));
  NAND2_X1  g1158(.A1(new_n1357), .A2(new_n1358), .ZN(new_n1359));
  OAI211_X1 g1159(.A(KEYINPUT127), .B(new_n1295), .C1(new_n1263), .C2(new_n1265), .ZN(new_n1360));
  NAND3_X1  g1160(.A1(new_n1359), .A2(new_n1306), .A3(new_n1360), .ZN(new_n1361));
  AND3_X1   g1161(.A1(new_n1325), .A2(new_n1329), .A3(new_n1319), .ZN(new_n1362));
  AOI21_X1  g1162(.A(new_n1319), .B1(new_n1325), .B2(new_n1329), .ZN(new_n1363));
  NOR2_X1   g1163(.A1(new_n1362), .A2(new_n1363), .ZN(new_n1364));
  XNOR2_X1  g1164(.A(new_n1361), .B(new_n1364), .ZN(G402));
endmodule


