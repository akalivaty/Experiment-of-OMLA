

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n510, n511, n512, n513,
         n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
         n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
         n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590,
         n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601,
         n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612,
         n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623,
         n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634,
         n635, n636, n637, n638, n639, n640, n641, n642, n643, n644, n645,
         n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, n656,
         n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n667,
         n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678,
         n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689,
         n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700,
         n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711,
         n712, n713, n714, n715, n716, n717, n718, n719, n720, n721, n722,
         n723, n724, n725, n726, n727, n728, n729, n730, n731, n732, n733,
         n734, n735, n736, n737, n738, n739, n740, n741, n742, n743, n744,
         n745, n746, n747, n748, n749, n750, n751, n752, n753, n754, n755,
         n756, n757, n758, n759, n760, n761, n762, n763, n764, n765, n766,
         n767, n768, n769, n770, n771, n772, n773, n774, n775, n776, n777,
         n778, n779, n780, n781, n782, n783, n784, n785, n786, n787, n788,
         n789, n790, n791, n792, n793, n794, n795, n796, n797, n798, n799,
         n800, n801, n802, n803, n804, n805, n806, n807, n808, n809, n810,
         n811, n812, n813, n814, n815, n816, n817, n818, n819, n820, n821,
         n822, n823, n824, n825, n826, n827, n828, n829, n830, n831, n832,
         n833, n834, n835, n836, n837, n838, n839, n840, n841, n842, n843,
         n844, n845, n846, n847, n848, n849, n850, n851, n852, n853, n854,
         n855, n856, n857, n858, n859, n860, n861, n862, n863, n864, n865,
         n866, n867, n868, n869, n870, n871, n872, n873, n874, n875, n876,
         n877, n878, n879, n880, n881, n882, n883, n884, n885, n886, n887,
         n888, n889, n890, n891, n892, n893, n894, n895, n896, n897, n898,
         n899, n900, n901, n902, n903, n904, n905, n906, n907, n908, n909,
         n910, n911, n912, n913, n914, n915, n916, n917, n918, n919, n920,
         n921, n922, n923, n924, n925, n926, n927, n928, n929, n930, n931,
         n932, n933, n934, n935, n936, n937, n938, n939, n940, n941, n942,
         n943, n944, n945, n946, n947, n948, n949, n950, n951, n952, n953,
         n954, n955, n956, n957, n958, n959, n960, n961, n962, n963, n964,
         n965, n966, n967, n968, n969, n970, n971, n972, n973, n974, n975,
         n976, n977, n978, n979, n980, n981, n982, n983, n984, n985, n986,
         n987, n988, n989, n990, n991, n992, n993, n994, n995, n996, n997,
         n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007,
         n1008, n1009;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NOR2_X1 U547 ( .A1(n721), .A2(n720), .ZN(n728) );
  INV_X1 U548 ( .A(n738), .ZN(n759) );
  XNOR2_X1 U549 ( .A(n767), .B(n766), .ZN(n768) );
  NOR2_X2 U550 ( .A1(n536), .A2(n535), .ZN(G160) );
  INV_X1 U551 ( .A(KEYINPUT97), .ZN(n710) );
  XNOR2_X1 U552 ( .A(n711), .B(n710), .ZN(n737) );
  NOR2_X1 U553 ( .A1(G651), .A2(n642), .ZN(n637) );
  INV_X1 U554 ( .A(G651), .ZN(n518) );
  NOR2_X1 U555 ( .A1(G543), .A2(n518), .ZN(n511) );
  XNOR2_X1 U556 ( .A(KEYINPUT1), .B(KEYINPUT67), .ZN(n510) );
  XNOR2_X1 U557 ( .A(n511), .B(n510), .ZN(n641) );
  NAND2_X1 U558 ( .A1(G63), .A2(n641), .ZN(n513) );
  XOR2_X1 U559 ( .A(KEYINPUT0), .B(G543), .Z(n642) );
  NAND2_X1 U560 ( .A1(G51), .A2(n637), .ZN(n512) );
  NAND2_X1 U561 ( .A1(n513), .A2(n512), .ZN(n514) );
  XNOR2_X1 U562 ( .A(KEYINPUT6), .B(n514), .ZN(n523) );
  NOR2_X1 U563 ( .A1(G543), .A2(G651), .ZN(n515) );
  XNOR2_X1 U564 ( .A(n515), .B(KEYINPUT64), .ZN(n628) );
  NAND2_X1 U565 ( .A1(n628), .A2(G89), .ZN(n516) );
  XOR2_X1 U566 ( .A(KEYINPUT73), .B(n516), .Z(n517) );
  XNOR2_X1 U567 ( .A(n517), .B(KEYINPUT4), .ZN(n520) );
  NOR2_X1 U568 ( .A1(n642), .A2(n518), .ZN(n631) );
  NAND2_X1 U569 ( .A1(G76), .A2(n631), .ZN(n519) );
  NAND2_X1 U570 ( .A1(n520), .A2(n519), .ZN(n521) );
  XOR2_X1 U571 ( .A(n521), .B(KEYINPUT5), .Z(n522) );
  NOR2_X1 U572 ( .A1(n523), .A2(n522), .ZN(n524) );
  XOR2_X1 U573 ( .A(KEYINPUT7), .B(n524), .Z(n525) );
  XNOR2_X1 U574 ( .A(KEYINPUT74), .B(n525), .ZN(G168) );
  XOR2_X1 U575 ( .A(KEYINPUT8), .B(G168), .Z(G286) );
  AND2_X1 U576 ( .A1(G2104), .A2(G2105), .ZN(n871) );
  NAND2_X1 U577 ( .A1(G113), .A2(n871), .ZN(n528) );
  NOR2_X1 U578 ( .A1(G2104), .A2(G2105), .ZN(n526) );
  XOR2_X2 U579 ( .A(KEYINPUT17), .B(n526), .Z(n867) );
  NAND2_X1 U580 ( .A1(G137), .A2(n867), .ZN(n527) );
  NAND2_X1 U581 ( .A1(n528), .A2(n527), .ZN(n536) );
  INV_X1 U582 ( .A(KEYINPUT23), .ZN(n530) );
  XNOR2_X1 U583 ( .A(G2104), .B(KEYINPUT65), .ZN(n531) );
  NOR2_X4 U584 ( .A1(G2105), .A2(n531), .ZN(n866) );
  NAND2_X1 U585 ( .A1(G101), .A2(n866), .ZN(n529) );
  XNOR2_X1 U586 ( .A(n530), .B(n529), .ZN(n534) );
  AND2_X1 U587 ( .A1(n531), .A2(G2105), .ZN(n549) );
  INV_X1 U588 ( .A(n549), .ZN(n532) );
  INV_X1 U589 ( .A(n532), .ZN(n870) );
  NAND2_X1 U590 ( .A1(n870), .A2(G125), .ZN(n533) );
  NAND2_X1 U591 ( .A1(n534), .A2(n533), .ZN(n535) );
  AND2_X1 U592 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U593 ( .A(G108), .ZN(G238) );
  INV_X1 U594 ( .A(G132), .ZN(G219) );
  INV_X1 U595 ( .A(G82), .ZN(G220) );
  NAND2_X1 U596 ( .A1(n631), .A2(G77), .ZN(n538) );
  NAND2_X1 U597 ( .A1(G90), .A2(n628), .ZN(n537) );
  NAND2_X1 U598 ( .A1(n538), .A2(n537), .ZN(n539) );
  XNOR2_X1 U599 ( .A(n539), .B(KEYINPUT9), .ZN(n541) );
  NAND2_X1 U600 ( .A1(G52), .A2(n637), .ZN(n540) );
  NAND2_X1 U601 ( .A1(n541), .A2(n540), .ZN(n544) );
  NAND2_X1 U602 ( .A1(n641), .A2(G64), .ZN(n542) );
  XOR2_X1 U603 ( .A(KEYINPUT68), .B(n542), .Z(n543) );
  NOR2_X1 U604 ( .A1(n544), .A2(n543), .ZN(G171) );
  NAND2_X1 U605 ( .A1(G102), .A2(n866), .ZN(n545) );
  XNOR2_X1 U606 ( .A(n545), .B(KEYINPUT90), .ZN(n548) );
  NAND2_X1 U607 ( .A1(G114), .A2(n871), .ZN(n546) );
  XOR2_X1 U608 ( .A(KEYINPUT89), .B(n546), .Z(n547) );
  NAND2_X1 U609 ( .A1(n548), .A2(n547), .ZN(n554) );
  NAND2_X1 U610 ( .A1(n549), .A2(G126), .ZN(n550) );
  XNOR2_X1 U611 ( .A(n550), .B(KEYINPUT88), .ZN(n552) );
  NAND2_X1 U612 ( .A1(G138), .A2(n867), .ZN(n551) );
  NAND2_X1 U613 ( .A1(n552), .A2(n551), .ZN(n553) );
  NOR2_X1 U614 ( .A1(n554), .A2(n553), .ZN(G164) );
  NAND2_X1 U615 ( .A1(G7), .A2(G661), .ZN(n555) );
  XNOR2_X1 U616 ( .A(n555), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U617 ( .A(G223), .ZN(n810) );
  NAND2_X1 U618 ( .A1(n810), .A2(G567), .ZN(n556) );
  XOR2_X1 U619 ( .A(KEYINPUT11), .B(n556), .Z(G234) );
  NAND2_X1 U620 ( .A1(G56), .A2(n641), .ZN(n557) );
  XOR2_X1 U621 ( .A(KEYINPUT14), .B(n557), .Z(n563) );
  NAND2_X1 U622 ( .A1(G81), .A2(n628), .ZN(n558) );
  XNOR2_X1 U623 ( .A(n558), .B(KEYINPUT12), .ZN(n560) );
  NAND2_X1 U624 ( .A1(G68), .A2(n631), .ZN(n559) );
  NAND2_X1 U625 ( .A1(n560), .A2(n559), .ZN(n561) );
  XOR2_X1 U626 ( .A(KEYINPUT13), .B(n561), .Z(n562) );
  NOR2_X1 U627 ( .A1(n563), .A2(n562), .ZN(n565) );
  NAND2_X1 U628 ( .A1(n637), .A2(G43), .ZN(n564) );
  NAND2_X1 U629 ( .A1(n565), .A2(n564), .ZN(n973) );
  XNOR2_X1 U630 ( .A(G860), .B(KEYINPUT71), .ZN(n586) );
  OR2_X1 U631 ( .A1(n973), .A2(n586), .ZN(G153) );
  INV_X1 U632 ( .A(G171), .ZN(G301) );
  NAND2_X1 U633 ( .A1(n641), .A2(G66), .ZN(n567) );
  NAND2_X1 U634 ( .A1(G92), .A2(n628), .ZN(n566) );
  NAND2_X1 U635 ( .A1(n567), .A2(n566), .ZN(n571) );
  NAND2_X1 U636 ( .A1(G79), .A2(n631), .ZN(n569) );
  NAND2_X1 U637 ( .A1(G54), .A2(n637), .ZN(n568) );
  NAND2_X1 U638 ( .A1(n569), .A2(n568), .ZN(n570) );
  NOR2_X1 U639 ( .A1(n571), .A2(n570), .ZN(n573) );
  XNOR2_X1 U640 ( .A(KEYINPUT72), .B(KEYINPUT15), .ZN(n572) );
  XNOR2_X1 U641 ( .A(n573), .B(n572), .ZN(n889) );
  NOR2_X1 U642 ( .A1(n889), .A2(G868), .ZN(n575) );
  INV_X1 U643 ( .A(G868), .ZN(n583) );
  NOR2_X1 U644 ( .A1(n583), .A2(G301), .ZN(n574) );
  NOR2_X1 U645 ( .A1(n575), .A2(n574), .ZN(G284) );
  NAND2_X1 U646 ( .A1(n631), .A2(G78), .ZN(n577) );
  NAND2_X1 U647 ( .A1(G91), .A2(n628), .ZN(n576) );
  NAND2_X1 U648 ( .A1(n577), .A2(n576), .ZN(n582) );
  NAND2_X1 U649 ( .A1(G65), .A2(n641), .ZN(n579) );
  NAND2_X1 U650 ( .A1(G53), .A2(n637), .ZN(n578) );
  NAND2_X1 U651 ( .A1(n579), .A2(n578), .ZN(n580) );
  XOR2_X1 U652 ( .A(KEYINPUT69), .B(n580), .Z(n581) );
  NOR2_X1 U653 ( .A1(n582), .A2(n581), .ZN(n964) );
  XOR2_X1 U654 ( .A(n964), .B(KEYINPUT70), .Z(G299) );
  NAND2_X1 U655 ( .A1(G868), .A2(G286), .ZN(n585) );
  NAND2_X1 U656 ( .A1(G299), .A2(n583), .ZN(n584) );
  NAND2_X1 U657 ( .A1(n585), .A2(n584), .ZN(G297) );
  NAND2_X1 U658 ( .A1(n586), .A2(G559), .ZN(n587) );
  INV_X1 U659 ( .A(n889), .ZN(n952) );
  NAND2_X1 U660 ( .A1(n587), .A2(n952), .ZN(n588) );
  XNOR2_X1 U661 ( .A(n588), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U662 ( .A1(G868), .A2(n973), .ZN(n589) );
  XOR2_X1 U663 ( .A(KEYINPUT75), .B(n589), .Z(n593) );
  NAND2_X1 U664 ( .A1(G868), .A2(n952), .ZN(n590) );
  NOR2_X1 U665 ( .A1(G559), .A2(n590), .ZN(n591) );
  XNOR2_X1 U666 ( .A(KEYINPUT76), .B(n591), .ZN(n592) );
  NOR2_X1 U667 ( .A1(n593), .A2(n592), .ZN(G282) );
  NAND2_X1 U668 ( .A1(G99), .A2(n866), .ZN(n595) );
  NAND2_X1 U669 ( .A1(G111), .A2(n871), .ZN(n594) );
  NAND2_X1 U670 ( .A1(n595), .A2(n594), .ZN(n596) );
  XNOR2_X1 U671 ( .A(KEYINPUT78), .B(n596), .ZN(n602) );
  NAND2_X1 U672 ( .A1(n870), .A2(G123), .ZN(n597) );
  XNOR2_X1 U673 ( .A(n597), .B(KEYINPUT18), .ZN(n599) );
  NAND2_X1 U674 ( .A1(G135), .A2(n867), .ZN(n598) );
  NAND2_X1 U675 ( .A1(n599), .A2(n598), .ZN(n600) );
  XOR2_X1 U676 ( .A(KEYINPUT77), .B(n600), .Z(n601) );
  NOR2_X1 U677 ( .A1(n602), .A2(n601), .ZN(n908) );
  XNOR2_X1 U678 ( .A(G2096), .B(n908), .ZN(n604) );
  INV_X1 U679 ( .A(G2100), .ZN(n603) );
  NAND2_X1 U680 ( .A1(n604), .A2(n603), .ZN(G156) );
  NAND2_X1 U681 ( .A1(n952), .A2(G559), .ZN(n605) );
  XNOR2_X1 U682 ( .A(n973), .B(n605), .ZN(n654) );
  NOR2_X1 U683 ( .A1(n654), .A2(G860), .ZN(n613) );
  NAND2_X1 U684 ( .A1(n641), .A2(G67), .ZN(n608) );
  NAND2_X1 U685 ( .A1(n628), .A2(G93), .ZN(n606) );
  XOR2_X1 U686 ( .A(KEYINPUT79), .B(n606), .Z(n607) );
  NAND2_X1 U687 ( .A1(n608), .A2(n607), .ZN(n612) );
  NAND2_X1 U688 ( .A1(G80), .A2(n631), .ZN(n610) );
  NAND2_X1 U689 ( .A1(G55), .A2(n637), .ZN(n609) );
  NAND2_X1 U690 ( .A1(n610), .A2(n609), .ZN(n611) );
  NOR2_X1 U691 ( .A1(n612), .A2(n611), .ZN(n646) );
  XNOR2_X1 U692 ( .A(n613), .B(n646), .ZN(G145) );
  NAND2_X1 U693 ( .A1(G62), .A2(n641), .ZN(n615) );
  NAND2_X1 U694 ( .A1(G50), .A2(n637), .ZN(n614) );
  NAND2_X1 U695 ( .A1(n615), .A2(n614), .ZN(n616) );
  XOR2_X1 U696 ( .A(KEYINPUT80), .B(n616), .Z(n620) );
  NAND2_X1 U697 ( .A1(n628), .A2(G88), .ZN(n618) );
  NAND2_X1 U698 ( .A1(n631), .A2(G75), .ZN(n617) );
  AND2_X1 U699 ( .A1(n618), .A2(n617), .ZN(n619) );
  NAND2_X1 U700 ( .A1(n620), .A2(n619), .ZN(G303) );
  INV_X1 U701 ( .A(G303), .ZN(G166) );
  NAND2_X1 U702 ( .A1(G72), .A2(n631), .ZN(n622) );
  NAND2_X1 U703 ( .A1(G47), .A2(n637), .ZN(n621) );
  NAND2_X1 U704 ( .A1(n622), .A2(n621), .ZN(n625) );
  NAND2_X1 U705 ( .A1(n628), .A2(G85), .ZN(n623) );
  XOR2_X1 U706 ( .A(KEYINPUT66), .B(n623), .Z(n624) );
  NOR2_X1 U707 ( .A1(n625), .A2(n624), .ZN(n627) );
  NAND2_X1 U708 ( .A1(n641), .A2(G60), .ZN(n626) );
  NAND2_X1 U709 ( .A1(n627), .A2(n626), .ZN(G290) );
  NAND2_X1 U710 ( .A1(n641), .A2(G61), .ZN(n630) );
  NAND2_X1 U711 ( .A1(G86), .A2(n628), .ZN(n629) );
  NAND2_X1 U712 ( .A1(n630), .A2(n629), .ZN(n634) );
  NAND2_X1 U713 ( .A1(n631), .A2(G73), .ZN(n632) );
  XOR2_X1 U714 ( .A(KEYINPUT2), .B(n632), .Z(n633) );
  NOR2_X1 U715 ( .A1(n634), .A2(n633), .ZN(n636) );
  NAND2_X1 U716 ( .A1(n637), .A2(G48), .ZN(n635) );
  NAND2_X1 U717 ( .A1(n636), .A2(n635), .ZN(G305) );
  NAND2_X1 U718 ( .A1(G49), .A2(n637), .ZN(n639) );
  NAND2_X1 U719 ( .A1(G74), .A2(G651), .ZN(n638) );
  NAND2_X1 U720 ( .A1(n639), .A2(n638), .ZN(n640) );
  NOR2_X1 U721 ( .A1(n641), .A2(n640), .ZN(n644) );
  NAND2_X1 U722 ( .A1(n642), .A2(G87), .ZN(n643) );
  NAND2_X1 U723 ( .A1(n644), .A2(n643), .ZN(G288) );
  NOR2_X1 U724 ( .A1(G868), .A2(n646), .ZN(n645) );
  XNOR2_X1 U725 ( .A(n645), .B(KEYINPUT83), .ZN(n657) );
  XOR2_X1 U726 ( .A(KEYINPUT82), .B(KEYINPUT81), .Z(n648) );
  XNOR2_X1 U727 ( .A(KEYINPUT19), .B(n646), .ZN(n647) );
  XNOR2_X1 U728 ( .A(n648), .B(n647), .ZN(n651) );
  XNOR2_X1 U729 ( .A(G166), .B(G290), .ZN(n649) );
  XNOR2_X1 U730 ( .A(n649), .B(G305), .ZN(n650) );
  XNOR2_X1 U731 ( .A(n651), .B(n650), .ZN(n653) );
  XNOR2_X1 U732 ( .A(G288), .B(G299), .ZN(n652) );
  XNOR2_X1 U733 ( .A(n653), .B(n652), .ZN(n892) );
  XOR2_X1 U734 ( .A(n892), .B(n654), .Z(n655) );
  NAND2_X1 U735 ( .A1(G868), .A2(n655), .ZN(n656) );
  NAND2_X1 U736 ( .A1(n657), .A2(n656), .ZN(G295) );
  NAND2_X1 U737 ( .A1(G2084), .A2(G2078), .ZN(n658) );
  XOR2_X1 U738 ( .A(KEYINPUT20), .B(n658), .Z(n659) );
  NAND2_X1 U739 ( .A1(G2090), .A2(n659), .ZN(n660) );
  XNOR2_X1 U740 ( .A(KEYINPUT21), .B(n660), .ZN(n661) );
  NAND2_X1 U741 ( .A1(n661), .A2(G2072), .ZN(n662) );
  XNOR2_X1 U742 ( .A(KEYINPUT84), .B(n662), .ZN(G158) );
  XNOR2_X1 U743 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U744 ( .A1(G220), .A2(G219), .ZN(n663) );
  XOR2_X1 U745 ( .A(KEYINPUT22), .B(n663), .Z(n664) );
  NOR2_X1 U746 ( .A1(G218), .A2(n664), .ZN(n665) );
  XOR2_X1 U747 ( .A(KEYINPUT85), .B(n665), .Z(n666) );
  NAND2_X1 U748 ( .A1(G96), .A2(n666), .ZN(n814) );
  NAND2_X1 U749 ( .A1(G2106), .A2(n814), .ZN(n667) );
  XNOR2_X1 U750 ( .A(n667), .B(KEYINPUT86), .ZN(n671) );
  NAND2_X1 U751 ( .A1(G120), .A2(G69), .ZN(n668) );
  NOR2_X1 U752 ( .A1(G238), .A2(n668), .ZN(n669) );
  NAND2_X1 U753 ( .A1(G57), .A2(n669), .ZN(n815) );
  NAND2_X1 U754 ( .A1(G567), .A2(n815), .ZN(n670) );
  NAND2_X1 U755 ( .A1(n671), .A2(n670), .ZN(n672) );
  XOR2_X1 U756 ( .A(KEYINPUT87), .B(n672), .Z(n816) );
  NAND2_X1 U757 ( .A1(G661), .A2(G483), .ZN(n673) );
  NOR2_X1 U758 ( .A1(n816), .A2(n673), .ZN(n813) );
  NAND2_X1 U759 ( .A1(n813), .A2(G36), .ZN(G176) );
  NAND2_X1 U760 ( .A1(G117), .A2(n871), .ZN(n675) );
  NAND2_X1 U761 ( .A1(G141), .A2(n867), .ZN(n674) );
  NAND2_X1 U762 ( .A1(n675), .A2(n674), .ZN(n678) );
  NAND2_X1 U763 ( .A1(n866), .A2(G105), .ZN(n676) );
  XOR2_X1 U764 ( .A(KEYINPUT38), .B(n676), .Z(n677) );
  NOR2_X1 U765 ( .A1(n678), .A2(n677), .ZN(n680) );
  NAND2_X1 U766 ( .A1(n870), .A2(G129), .ZN(n679) );
  NAND2_X1 U767 ( .A1(n680), .A2(n679), .ZN(n881) );
  NAND2_X1 U768 ( .A1(n881), .A2(G1996), .ZN(n689) );
  NAND2_X1 U769 ( .A1(G95), .A2(n866), .ZN(n682) );
  NAND2_X1 U770 ( .A1(G107), .A2(n871), .ZN(n681) );
  NAND2_X1 U771 ( .A1(n682), .A2(n681), .ZN(n685) );
  NAND2_X1 U772 ( .A1(n867), .A2(G131), .ZN(n683) );
  XOR2_X1 U773 ( .A(KEYINPUT94), .B(n683), .Z(n684) );
  NOR2_X1 U774 ( .A1(n685), .A2(n684), .ZN(n687) );
  NAND2_X1 U775 ( .A1(n870), .A2(G119), .ZN(n686) );
  NAND2_X1 U776 ( .A1(n687), .A2(n686), .ZN(n878) );
  NAND2_X1 U777 ( .A1(G1991), .A2(n878), .ZN(n688) );
  NAND2_X1 U778 ( .A1(n689), .A2(n688), .ZN(n690) );
  XNOR2_X1 U779 ( .A(n690), .B(KEYINPUT95), .ZN(n907) );
  NOR2_X1 U780 ( .A1(G164), .A2(G1384), .ZN(n707) );
  NAND2_X1 U781 ( .A1(G160), .A2(G40), .ZN(n705) );
  NOR2_X1 U782 ( .A1(n707), .A2(n705), .ZN(n691) );
  XOR2_X1 U783 ( .A(KEYINPUT91), .B(n691), .Z(n804) );
  INV_X1 U784 ( .A(n804), .ZN(n692) );
  NOR2_X1 U785 ( .A1(n907), .A2(n692), .ZN(n795) );
  XOR2_X1 U786 ( .A(KEYINPUT96), .B(n795), .Z(n704) );
  XNOR2_X1 U787 ( .A(KEYINPUT93), .B(KEYINPUT35), .ZN(n696) );
  NAND2_X1 U788 ( .A1(G128), .A2(n870), .ZN(n694) );
  NAND2_X1 U789 ( .A1(G116), .A2(n871), .ZN(n693) );
  NAND2_X1 U790 ( .A1(n694), .A2(n693), .ZN(n695) );
  XNOR2_X1 U791 ( .A(n696), .B(n695), .ZN(n702) );
  NAND2_X1 U792 ( .A1(n866), .A2(G104), .ZN(n697) );
  XNOR2_X1 U793 ( .A(n697), .B(KEYINPUT92), .ZN(n699) );
  NAND2_X1 U794 ( .A1(G140), .A2(n867), .ZN(n698) );
  NAND2_X1 U795 ( .A1(n699), .A2(n698), .ZN(n700) );
  XNOR2_X1 U796 ( .A(KEYINPUT34), .B(n700), .ZN(n701) );
  NOR2_X1 U797 ( .A1(n702), .A2(n701), .ZN(n703) );
  XNOR2_X1 U798 ( .A(KEYINPUT36), .B(n703), .ZN(n885) );
  XNOR2_X1 U799 ( .A(G2067), .B(KEYINPUT37), .ZN(n801) );
  NOR2_X1 U800 ( .A1(n885), .A2(n801), .ZN(n913) );
  NAND2_X1 U801 ( .A1(n804), .A2(n913), .ZN(n799) );
  NAND2_X1 U802 ( .A1(n704), .A2(n799), .ZN(n790) );
  INV_X1 U803 ( .A(n705), .ZN(n706) );
  NAND2_X1 U804 ( .A1(n707), .A2(n706), .ZN(n711) );
  INV_X1 U805 ( .A(n711), .ZN(n738) );
  NAND2_X1 U806 ( .A1(G8), .A2(n759), .ZN(n783) );
  NOR2_X1 U807 ( .A1(G1981), .A2(G305), .ZN(n708) );
  XOR2_X1 U808 ( .A(n708), .B(KEYINPUT24), .Z(n709) );
  NOR2_X1 U809 ( .A1(n783), .A2(n709), .ZN(n788) );
  NOR2_X1 U810 ( .A1(G2084), .A2(n759), .ZN(n743) );
  NAND2_X1 U811 ( .A1(G8), .A2(n743), .ZN(n757) );
  NOR2_X1 U812 ( .A1(G1966), .A2(n783), .ZN(n755) );
  INV_X1 U813 ( .A(n737), .ZN(n712) );
  NAND2_X1 U814 ( .A1(n712), .A2(G2072), .ZN(n713) );
  XNOR2_X1 U815 ( .A(n713), .B(KEYINPUT27), .ZN(n715) );
  AND2_X1 U816 ( .A1(G1956), .A2(n737), .ZN(n714) );
  NOR2_X1 U817 ( .A1(n715), .A2(n714), .ZN(n731) );
  NOR2_X1 U818 ( .A1(n731), .A2(n964), .ZN(n718) );
  XNOR2_X1 U819 ( .A(KEYINPUT28), .B(KEYINPUT99), .ZN(n716) );
  XNOR2_X1 U820 ( .A(n716), .B(KEYINPUT98), .ZN(n717) );
  XNOR2_X1 U821 ( .A(n718), .B(n717), .ZN(n735) );
  NAND2_X1 U822 ( .A1(G1348), .A2(n759), .ZN(n719) );
  XOR2_X1 U823 ( .A(KEYINPUT100), .B(n719), .Z(n721) );
  INV_X1 U824 ( .A(G2067), .ZN(n929) );
  NOR2_X1 U825 ( .A1(n929), .A2(n737), .ZN(n720) );
  NAND2_X1 U826 ( .A1(n952), .A2(n728), .ZN(n727) );
  AND2_X1 U827 ( .A1(n738), .A2(G1996), .ZN(n722) );
  XOR2_X1 U828 ( .A(n722), .B(KEYINPUT26), .Z(n724) );
  NAND2_X1 U829 ( .A1(n759), .A2(G1341), .ZN(n723) );
  NAND2_X1 U830 ( .A1(n724), .A2(n723), .ZN(n725) );
  OR2_X1 U831 ( .A1(n973), .A2(n725), .ZN(n726) );
  NAND2_X1 U832 ( .A1(n727), .A2(n726), .ZN(n730) );
  OR2_X1 U833 ( .A1(n728), .A2(n952), .ZN(n729) );
  NAND2_X1 U834 ( .A1(n730), .A2(n729), .ZN(n733) );
  NAND2_X1 U835 ( .A1(n731), .A2(n964), .ZN(n732) );
  NAND2_X1 U836 ( .A1(n733), .A2(n732), .ZN(n734) );
  NAND2_X1 U837 ( .A1(n735), .A2(n734), .ZN(n736) );
  XNOR2_X1 U838 ( .A(n736), .B(KEYINPUT29), .ZN(n742) );
  XOR2_X1 U839 ( .A(KEYINPUT25), .B(G2078), .Z(n935) );
  NOR2_X1 U840 ( .A1(n935), .A2(n737), .ZN(n740) );
  NOR2_X1 U841 ( .A1(n738), .A2(G1961), .ZN(n739) );
  NOR2_X1 U842 ( .A1(n740), .A2(n739), .ZN(n747) );
  NOR2_X1 U843 ( .A1(G301), .A2(n747), .ZN(n741) );
  NOR2_X1 U844 ( .A1(n742), .A2(n741), .ZN(n752) );
  NOR2_X1 U845 ( .A1(n755), .A2(n743), .ZN(n744) );
  NAND2_X1 U846 ( .A1(G8), .A2(n744), .ZN(n745) );
  XNOR2_X1 U847 ( .A(KEYINPUT30), .B(n745), .ZN(n746) );
  NOR2_X1 U848 ( .A1(G168), .A2(n746), .ZN(n749) );
  AND2_X1 U849 ( .A1(G301), .A2(n747), .ZN(n748) );
  NOR2_X1 U850 ( .A1(n749), .A2(n748), .ZN(n750) );
  XNOR2_X1 U851 ( .A(n750), .B(KEYINPUT31), .ZN(n751) );
  NOR2_X1 U852 ( .A1(n752), .A2(n751), .ZN(n753) );
  XNOR2_X1 U853 ( .A(n753), .B(KEYINPUT101), .ZN(n758) );
  XOR2_X1 U854 ( .A(n758), .B(KEYINPUT102), .Z(n754) );
  NOR2_X1 U855 ( .A1(n755), .A2(n754), .ZN(n756) );
  NAND2_X1 U856 ( .A1(n757), .A2(n756), .ZN(n769) );
  NAND2_X1 U857 ( .A1(n758), .A2(G286), .ZN(n764) );
  NOR2_X1 U858 ( .A1(G1971), .A2(n783), .ZN(n761) );
  NOR2_X1 U859 ( .A1(G2090), .A2(n759), .ZN(n760) );
  NOR2_X1 U860 ( .A1(n761), .A2(n760), .ZN(n762) );
  NAND2_X1 U861 ( .A1(n762), .A2(G303), .ZN(n763) );
  NAND2_X1 U862 ( .A1(n764), .A2(n763), .ZN(n765) );
  NAND2_X1 U863 ( .A1(G8), .A2(n765), .ZN(n767) );
  XOR2_X1 U864 ( .A(KEYINPUT32), .B(KEYINPUT103), .Z(n766) );
  NAND2_X1 U865 ( .A1(n769), .A2(n768), .ZN(n781) );
  NOR2_X1 U866 ( .A1(G1976), .A2(G288), .ZN(n961) );
  NOR2_X1 U867 ( .A1(G1971), .A2(G303), .ZN(n770) );
  NOR2_X1 U868 ( .A1(n961), .A2(n770), .ZN(n771) );
  NAND2_X1 U869 ( .A1(n781), .A2(n771), .ZN(n772) );
  NAND2_X1 U870 ( .A1(G1976), .A2(G288), .ZN(n962) );
  NAND2_X1 U871 ( .A1(n772), .A2(n962), .ZN(n773) );
  NOR2_X1 U872 ( .A1(n783), .A2(n773), .ZN(n774) );
  NOR2_X1 U873 ( .A1(KEYINPUT33), .A2(n774), .ZN(n777) );
  NAND2_X1 U874 ( .A1(n961), .A2(KEYINPUT33), .ZN(n775) );
  NOR2_X1 U875 ( .A1(n775), .A2(n783), .ZN(n776) );
  NOR2_X1 U876 ( .A1(n777), .A2(n776), .ZN(n778) );
  XOR2_X1 U877 ( .A(G1981), .B(G305), .Z(n957) );
  NAND2_X1 U878 ( .A1(n778), .A2(n957), .ZN(n786) );
  NOR2_X1 U879 ( .A1(G2090), .A2(G303), .ZN(n779) );
  XNOR2_X1 U880 ( .A(n779), .B(KEYINPUT104), .ZN(n780) );
  NAND2_X1 U881 ( .A1(n780), .A2(G8), .ZN(n782) );
  NAND2_X1 U882 ( .A1(n782), .A2(n781), .ZN(n784) );
  NAND2_X1 U883 ( .A1(n784), .A2(n783), .ZN(n785) );
  NAND2_X1 U884 ( .A1(n786), .A2(n785), .ZN(n787) );
  NOR2_X1 U885 ( .A1(n788), .A2(n787), .ZN(n789) );
  NOR2_X1 U886 ( .A1(n790), .A2(n789), .ZN(n792) );
  XNOR2_X1 U887 ( .A(G1986), .B(G290), .ZN(n970) );
  NAND2_X1 U888 ( .A1(n970), .A2(n804), .ZN(n791) );
  NAND2_X1 U889 ( .A1(n792), .A2(n791), .ZN(n807) );
  XOR2_X1 U890 ( .A(KEYINPUT105), .B(KEYINPUT39), .Z(n798) );
  NOR2_X1 U891 ( .A1(G1996), .A2(n881), .ZN(n904) );
  NOR2_X1 U892 ( .A1(G1986), .A2(G290), .ZN(n793) );
  NOR2_X1 U893 ( .A1(G1991), .A2(n878), .ZN(n909) );
  NOR2_X1 U894 ( .A1(n793), .A2(n909), .ZN(n794) );
  NOR2_X1 U895 ( .A1(n795), .A2(n794), .ZN(n796) );
  NOR2_X1 U896 ( .A1(n904), .A2(n796), .ZN(n797) );
  XNOR2_X1 U897 ( .A(n798), .B(n797), .ZN(n800) );
  NAND2_X1 U898 ( .A1(n800), .A2(n799), .ZN(n803) );
  NAND2_X1 U899 ( .A1(n885), .A2(n801), .ZN(n802) );
  XNOR2_X1 U900 ( .A(KEYINPUT106), .B(n802), .ZN(n919) );
  NAND2_X1 U901 ( .A1(n803), .A2(n919), .ZN(n805) );
  NAND2_X1 U902 ( .A1(n805), .A2(n804), .ZN(n806) );
  NAND2_X1 U903 ( .A1(n807), .A2(n806), .ZN(n809) );
  XOR2_X1 U904 ( .A(KEYINPUT107), .B(KEYINPUT40), .Z(n808) );
  XNOR2_X1 U905 ( .A(n809), .B(n808), .ZN(G329) );
  NAND2_X1 U906 ( .A1(G2106), .A2(n810), .ZN(G217) );
  AND2_X1 U907 ( .A1(G15), .A2(G2), .ZN(n811) );
  NAND2_X1 U908 ( .A1(G661), .A2(n811), .ZN(G259) );
  NAND2_X1 U909 ( .A1(G3), .A2(G1), .ZN(n812) );
  NAND2_X1 U910 ( .A1(n813), .A2(n812), .ZN(G188) );
  XNOR2_X1 U911 ( .A(G120), .B(KEYINPUT111), .ZN(G236) );
  XOR2_X1 U912 ( .A(G69), .B(KEYINPUT112), .Z(G235) );
  INV_X1 U914 ( .A(G96), .ZN(G221) );
  NOR2_X1 U915 ( .A1(n815), .A2(n814), .ZN(G325) );
  INV_X1 U916 ( .A(G325), .ZN(G261) );
  XNOR2_X1 U917 ( .A(KEYINPUT113), .B(n816), .ZN(G319) );
  XOR2_X1 U918 ( .A(G2096), .B(KEYINPUT43), .Z(n818) );
  XNOR2_X1 U919 ( .A(G2090), .B(KEYINPUT42), .ZN(n817) );
  XNOR2_X1 U920 ( .A(n818), .B(n817), .ZN(n819) );
  XOR2_X1 U921 ( .A(n819), .B(G2678), .Z(n821) );
  XNOR2_X1 U922 ( .A(G2067), .B(G2072), .ZN(n820) );
  XNOR2_X1 U923 ( .A(n821), .B(n820), .ZN(n825) );
  XOR2_X1 U924 ( .A(KEYINPUT114), .B(G2100), .Z(n823) );
  XNOR2_X1 U925 ( .A(G2084), .B(G2078), .ZN(n822) );
  XNOR2_X1 U926 ( .A(n823), .B(n822), .ZN(n824) );
  XNOR2_X1 U927 ( .A(n825), .B(n824), .ZN(G227) );
  XOR2_X1 U928 ( .A(G1981), .B(G1971), .Z(n827) );
  XNOR2_X1 U929 ( .A(G1986), .B(G1966), .ZN(n826) );
  XNOR2_X1 U930 ( .A(n827), .B(n826), .ZN(n828) );
  XOR2_X1 U931 ( .A(n828), .B(KEYINPUT41), .Z(n830) );
  XNOR2_X1 U932 ( .A(G1996), .B(G1991), .ZN(n829) );
  XNOR2_X1 U933 ( .A(n830), .B(n829), .ZN(n834) );
  XOR2_X1 U934 ( .A(G2474), .B(G1976), .Z(n832) );
  XNOR2_X1 U935 ( .A(G1961), .B(G1956), .ZN(n831) );
  XNOR2_X1 U936 ( .A(n832), .B(n831), .ZN(n833) );
  XNOR2_X1 U937 ( .A(n834), .B(n833), .ZN(G229) );
  XNOR2_X1 U938 ( .A(KEYINPUT109), .B(G2427), .ZN(n844) );
  XOR2_X1 U939 ( .A(G2443), .B(G2438), .Z(n836) );
  XNOR2_X1 U940 ( .A(G2430), .B(G2454), .ZN(n835) );
  XNOR2_X1 U941 ( .A(n836), .B(n835), .ZN(n840) );
  XOR2_X1 U942 ( .A(KEYINPUT108), .B(G2435), .Z(n838) );
  XNOR2_X1 U943 ( .A(G1348), .B(G1341), .ZN(n837) );
  XNOR2_X1 U944 ( .A(n838), .B(n837), .ZN(n839) );
  XOR2_X1 U945 ( .A(n840), .B(n839), .Z(n842) );
  XNOR2_X1 U946 ( .A(G2446), .B(G2451), .ZN(n841) );
  XNOR2_X1 U947 ( .A(n842), .B(n841), .ZN(n843) );
  XNOR2_X1 U948 ( .A(n844), .B(n843), .ZN(n845) );
  NAND2_X1 U949 ( .A1(n845), .A2(G14), .ZN(n846) );
  XOR2_X1 U950 ( .A(KEYINPUT110), .B(n846), .Z(G401) );
  NAND2_X1 U951 ( .A1(n870), .A2(G124), .ZN(n847) );
  XNOR2_X1 U952 ( .A(n847), .B(KEYINPUT44), .ZN(n849) );
  NAND2_X1 U953 ( .A1(G112), .A2(n871), .ZN(n848) );
  NAND2_X1 U954 ( .A1(n849), .A2(n848), .ZN(n853) );
  NAND2_X1 U955 ( .A1(G100), .A2(n866), .ZN(n851) );
  NAND2_X1 U956 ( .A1(G136), .A2(n867), .ZN(n850) );
  NAND2_X1 U957 ( .A1(n851), .A2(n850), .ZN(n852) );
  NOR2_X1 U958 ( .A1(n853), .A2(n852), .ZN(G162) );
  XOR2_X1 U959 ( .A(KEYINPUT117), .B(KEYINPUT46), .Z(n864) );
  NAND2_X1 U960 ( .A1(G106), .A2(n866), .ZN(n855) );
  NAND2_X1 U961 ( .A1(G142), .A2(n867), .ZN(n854) );
  NAND2_X1 U962 ( .A1(n855), .A2(n854), .ZN(n856) );
  XNOR2_X1 U963 ( .A(n856), .B(KEYINPUT45), .ZN(n858) );
  NAND2_X1 U964 ( .A1(G130), .A2(n870), .ZN(n857) );
  NAND2_X1 U965 ( .A1(n858), .A2(n857), .ZN(n861) );
  NAND2_X1 U966 ( .A1(G118), .A2(n871), .ZN(n859) );
  XNOR2_X1 U967 ( .A(KEYINPUT115), .B(n859), .ZN(n860) );
  NOR2_X1 U968 ( .A1(n861), .A2(n860), .ZN(n862) );
  XNOR2_X1 U969 ( .A(KEYINPUT48), .B(n862), .ZN(n863) );
  XNOR2_X1 U970 ( .A(n864), .B(n863), .ZN(n865) );
  XNOR2_X1 U971 ( .A(n908), .B(n865), .ZN(n880) );
  NAND2_X1 U972 ( .A1(G103), .A2(n866), .ZN(n869) );
  NAND2_X1 U973 ( .A1(G139), .A2(n867), .ZN(n868) );
  NAND2_X1 U974 ( .A1(n869), .A2(n868), .ZN(n876) );
  NAND2_X1 U975 ( .A1(G127), .A2(n870), .ZN(n873) );
  NAND2_X1 U976 ( .A1(G115), .A2(n871), .ZN(n872) );
  NAND2_X1 U977 ( .A1(n873), .A2(n872), .ZN(n874) );
  XOR2_X1 U978 ( .A(KEYINPUT47), .B(n874), .Z(n875) );
  NOR2_X1 U979 ( .A1(n876), .A2(n875), .ZN(n877) );
  XOR2_X1 U980 ( .A(KEYINPUT116), .B(n877), .Z(n920) );
  XNOR2_X1 U981 ( .A(n878), .B(n920), .ZN(n879) );
  XNOR2_X1 U982 ( .A(n880), .B(n879), .ZN(n887) );
  XNOR2_X1 U983 ( .A(n881), .B(G162), .ZN(n883) );
  XNOR2_X1 U984 ( .A(G164), .B(G160), .ZN(n882) );
  XNOR2_X1 U985 ( .A(n883), .B(n882), .ZN(n884) );
  XOR2_X1 U986 ( .A(n885), .B(n884), .Z(n886) );
  XNOR2_X1 U987 ( .A(n887), .B(n886), .ZN(n888) );
  NOR2_X1 U988 ( .A1(G37), .A2(n888), .ZN(G395) );
  XNOR2_X1 U989 ( .A(n973), .B(KEYINPUT118), .ZN(n891) );
  XNOR2_X1 U990 ( .A(G171), .B(n889), .ZN(n890) );
  XNOR2_X1 U991 ( .A(n891), .B(n890), .ZN(n894) );
  XOR2_X1 U992 ( .A(G286), .B(n892), .Z(n893) );
  XNOR2_X1 U993 ( .A(n894), .B(n893), .ZN(n895) );
  NOR2_X1 U994 ( .A1(G37), .A2(n895), .ZN(n896) );
  XOR2_X1 U995 ( .A(KEYINPUT119), .B(n896), .Z(G397) );
  NOR2_X1 U996 ( .A1(G227), .A2(G229), .ZN(n898) );
  XNOR2_X1 U997 ( .A(KEYINPUT49), .B(KEYINPUT120), .ZN(n897) );
  XNOR2_X1 U998 ( .A(n898), .B(n897), .ZN(n899) );
  NOR2_X1 U999 ( .A1(n899), .A2(G401), .ZN(n901) );
  NOR2_X1 U1000 ( .A1(G395), .A2(G397), .ZN(n900) );
  AND2_X1 U1001 ( .A1(n901), .A2(n900), .ZN(n902) );
  NAND2_X1 U1002 ( .A1(G319), .A2(n902), .ZN(G225) );
  INV_X1 U1003 ( .A(G225), .ZN(G308) );
  INV_X1 U1004 ( .A(G57), .ZN(G237) );
  XOR2_X1 U1005 ( .A(G2090), .B(G162), .Z(n903) );
  NOR2_X1 U1006 ( .A1(n904), .A2(n903), .ZN(n905) );
  XOR2_X1 U1007 ( .A(KEYINPUT51), .B(n905), .Z(n906) );
  NAND2_X1 U1008 ( .A1(n907), .A2(n906), .ZN(n917) );
  NOR2_X1 U1009 ( .A1(n909), .A2(n908), .ZN(n910) );
  XOR2_X1 U1010 ( .A(KEYINPUT121), .B(n910), .Z(n912) );
  XNOR2_X1 U1011 ( .A(G160), .B(G2084), .ZN(n911) );
  NAND2_X1 U1012 ( .A1(n912), .A2(n911), .ZN(n914) );
  NOR2_X1 U1013 ( .A1(n914), .A2(n913), .ZN(n915) );
  XOR2_X1 U1014 ( .A(KEYINPUT122), .B(n915), .Z(n916) );
  NOR2_X1 U1015 ( .A1(n917), .A2(n916), .ZN(n918) );
  NAND2_X1 U1016 ( .A1(n919), .A2(n918), .ZN(n925) );
  XOR2_X1 U1017 ( .A(G164), .B(G2078), .Z(n922) );
  XNOR2_X1 U1018 ( .A(G2072), .B(n920), .ZN(n921) );
  NOR2_X1 U1019 ( .A1(n922), .A2(n921), .ZN(n923) );
  XOR2_X1 U1020 ( .A(KEYINPUT50), .B(n923), .Z(n924) );
  NOR2_X1 U1021 ( .A1(n925), .A2(n924), .ZN(n926) );
  XNOR2_X1 U1022 ( .A(KEYINPUT52), .B(n926), .ZN(n927) );
  INV_X1 U1023 ( .A(KEYINPUT55), .ZN(n948) );
  NAND2_X1 U1024 ( .A1(n927), .A2(n948), .ZN(n928) );
  NAND2_X1 U1025 ( .A1(n928), .A2(G29), .ZN(n1008) );
  XNOR2_X1 U1026 ( .A(G2090), .B(G35), .ZN(n943) );
  XNOR2_X1 U1027 ( .A(G26), .B(n929), .ZN(n934) );
  XOR2_X1 U1028 ( .A(G2072), .B(G33), .Z(n930) );
  NAND2_X1 U1029 ( .A1(n930), .A2(G28), .ZN(n932) );
  XNOR2_X1 U1030 ( .A(G25), .B(G1991), .ZN(n931) );
  NOR2_X1 U1031 ( .A1(n932), .A2(n931), .ZN(n933) );
  NAND2_X1 U1032 ( .A1(n934), .A2(n933), .ZN(n940) );
  XNOR2_X1 U1033 ( .A(G1996), .B(G32), .ZN(n937) );
  XNOR2_X1 U1034 ( .A(n935), .B(G27), .ZN(n936) );
  NOR2_X1 U1035 ( .A1(n937), .A2(n936), .ZN(n938) );
  XNOR2_X1 U1036 ( .A(n938), .B(KEYINPUT123), .ZN(n939) );
  NOR2_X1 U1037 ( .A1(n940), .A2(n939), .ZN(n941) );
  XNOR2_X1 U1038 ( .A(KEYINPUT53), .B(n941), .ZN(n942) );
  NOR2_X1 U1039 ( .A1(n943), .A2(n942), .ZN(n946) );
  XOR2_X1 U1040 ( .A(G2084), .B(G34), .Z(n944) );
  XNOR2_X1 U1041 ( .A(KEYINPUT54), .B(n944), .ZN(n945) );
  NAND2_X1 U1042 ( .A1(n946), .A2(n945), .ZN(n947) );
  XNOR2_X1 U1043 ( .A(n948), .B(n947), .ZN(n950) );
  INV_X1 U1044 ( .A(G29), .ZN(n949) );
  NAND2_X1 U1045 ( .A1(n950), .A2(n949), .ZN(n951) );
  NAND2_X1 U1046 ( .A1(G11), .A2(n951), .ZN(n1006) );
  XNOR2_X1 U1047 ( .A(G16), .B(KEYINPUT56), .ZN(n979) );
  XNOR2_X1 U1048 ( .A(G171), .B(G1961), .ZN(n955) );
  XNOR2_X1 U1049 ( .A(G1348), .B(KEYINPUT124), .ZN(n953) );
  XNOR2_X1 U1050 ( .A(n953), .B(n952), .ZN(n954) );
  NAND2_X1 U1051 ( .A1(n955), .A2(n954), .ZN(n956) );
  XNOR2_X1 U1052 ( .A(n956), .B(KEYINPUT125), .ZN(n977) );
  XNOR2_X1 U1053 ( .A(G1966), .B(G168), .ZN(n958) );
  NAND2_X1 U1054 ( .A1(n958), .A2(n957), .ZN(n959) );
  XNOR2_X1 U1055 ( .A(KEYINPUT57), .B(n959), .ZN(n972) );
  XNOR2_X1 U1056 ( .A(G1971), .B(G166), .ZN(n960) );
  XNOR2_X1 U1057 ( .A(n960), .B(KEYINPUT126), .ZN(n968) );
  INV_X1 U1058 ( .A(n961), .ZN(n963) );
  NAND2_X1 U1059 ( .A1(n963), .A2(n962), .ZN(n966) );
  XOR2_X1 U1060 ( .A(n964), .B(G1956), .Z(n965) );
  NOR2_X1 U1061 ( .A1(n966), .A2(n965), .ZN(n967) );
  NAND2_X1 U1062 ( .A1(n968), .A2(n967), .ZN(n969) );
  NOR2_X1 U1063 ( .A1(n970), .A2(n969), .ZN(n971) );
  NAND2_X1 U1064 ( .A1(n972), .A2(n971), .ZN(n975) );
  XNOR2_X1 U1065 ( .A(G1341), .B(n973), .ZN(n974) );
  NOR2_X1 U1066 ( .A1(n975), .A2(n974), .ZN(n976) );
  NAND2_X1 U1067 ( .A1(n977), .A2(n976), .ZN(n978) );
  NAND2_X1 U1068 ( .A1(n979), .A2(n978), .ZN(n1004) );
  INV_X1 U1069 ( .A(G16), .ZN(n1002) );
  XNOR2_X1 U1070 ( .A(G1348), .B(KEYINPUT59), .ZN(n980) );
  XNOR2_X1 U1071 ( .A(n980), .B(G4), .ZN(n984) );
  XNOR2_X1 U1072 ( .A(G1956), .B(G20), .ZN(n982) );
  XNOR2_X1 U1073 ( .A(G1981), .B(G6), .ZN(n981) );
  NOR2_X1 U1074 ( .A1(n982), .A2(n981), .ZN(n983) );
  NAND2_X1 U1075 ( .A1(n984), .A2(n983), .ZN(n987) );
  XOR2_X1 U1076 ( .A(KEYINPUT127), .B(G1341), .Z(n985) );
  XNOR2_X1 U1077 ( .A(G19), .B(n985), .ZN(n986) );
  NOR2_X1 U1078 ( .A1(n987), .A2(n986), .ZN(n988) );
  XNOR2_X1 U1079 ( .A(KEYINPUT60), .B(n988), .ZN(n992) );
  XNOR2_X1 U1080 ( .A(G1966), .B(G21), .ZN(n990) );
  XNOR2_X1 U1081 ( .A(G5), .B(G1961), .ZN(n989) );
  NOR2_X1 U1082 ( .A1(n990), .A2(n989), .ZN(n991) );
  NAND2_X1 U1083 ( .A1(n992), .A2(n991), .ZN(n999) );
  XNOR2_X1 U1084 ( .A(G1971), .B(G22), .ZN(n994) );
  XNOR2_X1 U1085 ( .A(G23), .B(G1976), .ZN(n993) );
  NOR2_X1 U1086 ( .A1(n994), .A2(n993), .ZN(n996) );
  XOR2_X1 U1087 ( .A(G1986), .B(G24), .Z(n995) );
  NAND2_X1 U1088 ( .A1(n996), .A2(n995), .ZN(n997) );
  XNOR2_X1 U1089 ( .A(KEYINPUT58), .B(n997), .ZN(n998) );
  NOR2_X1 U1090 ( .A1(n999), .A2(n998), .ZN(n1000) );
  XNOR2_X1 U1091 ( .A(KEYINPUT61), .B(n1000), .ZN(n1001) );
  NAND2_X1 U1092 ( .A1(n1002), .A2(n1001), .ZN(n1003) );
  NAND2_X1 U1093 ( .A1(n1004), .A2(n1003), .ZN(n1005) );
  NOR2_X1 U1094 ( .A1(n1006), .A2(n1005), .ZN(n1007) );
  NAND2_X1 U1095 ( .A1(n1008), .A2(n1007), .ZN(n1009) );
  XOR2_X1 U1096 ( .A(KEYINPUT62), .B(n1009), .Z(G311) );
  INV_X1 U1097 ( .A(G311), .ZN(G150) );
endmodule

