

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
         n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598,
         n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609,
         n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620,
         n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631,
         n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642,
         n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653,
         n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664,
         n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675,
         n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686,
         n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697,
         n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708,
         n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719,
         n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, n730,
         n731, n732, n733, n734, n735, n736, n737, n738, n739, n740, n741,
         n742, n743, n744, n745, n746, n747, n748, n749, n750, n751, n752,
         n753, n754;

  XNOR2_X1 U367 ( .A(n502), .B(n501), .ZN(n572) );
  XNOR2_X1 U368 ( .A(n470), .B(n469), .ZN(n739) );
  BUF_X1 U369 ( .A(G146), .Z(n346) );
  XNOR2_X1 U370 ( .A(n471), .B(G125), .ZN(n434) );
  NAND2_X2 U371 ( .A1(n620), .A2(n619), .ZN(n625) );
  AND2_X2 U372 ( .A1(n533), .A2(n686), .ZN(n530) );
  NOR2_X1 U373 ( .A1(G953), .A2(G237), .ZN(n438) );
  XNOR2_X1 U374 ( .A(n739), .B(n473), .ZN(n489) );
  NAND2_X2 U375 ( .A1(n357), .A2(n356), .ZN(n578) );
  AND2_X2 U376 ( .A1(n358), .A2(n400), .ZN(n356) );
  AND2_X4 U377 ( .A1(n625), .A2(n624), .ZN(n719) );
  XNOR2_X2 U378 ( .A(n733), .B(n353), .ZN(n645) );
  XNOR2_X2 U379 ( .A(n453), .B(n414), .ZN(n470) );
  XNOR2_X2 U380 ( .A(n408), .B(n485), .ZN(n733) );
  XOR2_X2 U381 ( .A(G131), .B(KEYINPUT70), .Z(n468) );
  XNOR2_X2 U382 ( .A(n684), .B(n504), .ZN(n590) );
  INV_X1 U383 ( .A(KEYINPUT48), .ZN(n384) );
  INV_X4 U384 ( .A(G953), .ZN(n742) );
  NOR2_X1 U385 ( .A1(n383), .A2(n378), .ZN(n387) );
  XNOR2_X1 U386 ( .A(n588), .B(KEYINPUT74), .ZN(n386) );
  XNOR2_X1 U387 ( .A(n601), .B(n367), .ZN(n389) );
  NOR2_X1 U388 ( .A1(n610), .A2(n594), .ZN(n595) );
  XNOR2_X1 U389 ( .A(n517), .B(n516), .ZN(n533) );
  XNOR2_X1 U390 ( .A(n392), .B(n391), .ZN(n724) );
  INV_X2 U391 ( .A(G128), .ZN(n355) );
  XNOR2_X1 U392 ( .A(G119), .B(G116), .ZN(n405) );
  INV_X2 U393 ( .A(n520), .ZN(n531) );
  XNOR2_X2 U394 ( .A(n430), .B(n429), .ZN(n520) );
  XNOR2_X2 U395 ( .A(n531), .B(KEYINPUT91), .ZN(n534) );
  NAND2_X1 U396 ( .A1(n750), .A2(KEYINPUT46), .ZN(n380) );
  XNOR2_X1 U397 ( .A(n369), .B(n407), .ZN(n485) );
  XNOR2_X1 U398 ( .A(n405), .B(KEYINPUT3), .ZN(n369) );
  INV_X1 U399 ( .A(KEYINPUT71), .ZN(n406) );
  XNOR2_X1 U400 ( .A(KEYINPUT87), .B(G110), .ZN(n403) );
  NAND2_X1 U401 ( .A1(n645), .A2(n618), .ZN(n352) );
  INV_X1 U402 ( .A(KEYINPUT30), .ZN(n375) );
  NAND2_X1 U403 ( .A1(n558), .A2(n375), .ZN(n374) );
  NAND2_X1 U404 ( .A1(n695), .A2(n375), .ZN(n373) );
  NOR2_X1 U405 ( .A1(n389), .A2(n608), .ZN(n383) );
  XNOR2_X1 U406 ( .A(n456), .B(n455), .ZN(n495) );
  XOR2_X1 U407 ( .A(KEYINPUT8), .B(KEYINPUT69), .Z(n455) );
  XNOR2_X1 U408 ( .A(n454), .B(KEYINPUT81), .ZN(n456) );
  XNOR2_X1 U409 ( .A(n434), .B(n433), .ZN(n494) );
  XOR2_X1 U410 ( .A(G137), .B(G140), .Z(n492) );
  AND2_X1 U411 ( .A1(n377), .A2(n564), .ZN(n376) );
  INV_X1 U412 ( .A(KEYINPUT19), .ZN(n398) );
  NAND2_X1 U413 ( .A1(n695), .A2(KEYINPUT19), .ZN(n400) );
  NOR2_X1 U414 ( .A1(n572), .A2(n515), .ZN(n517) );
  XNOR2_X1 U415 ( .A(n496), .B(n395), .ZN(n394) );
  XNOR2_X1 U416 ( .A(G119), .B(KEYINPUT24), .ZN(n395) );
  XNOR2_X1 U417 ( .A(KEYINPUT88), .B(KEYINPUT17), .ZN(n409) );
  XNOR2_X1 U418 ( .A(KEYINPUT18), .B(KEYINPUT79), .ZN(n411) );
  XOR2_X1 U419 ( .A(KEYINPUT66), .B(G101), .Z(n472) );
  AND2_X1 U420 ( .A1(n388), .A2(n608), .ZN(n382) );
  NAND2_X1 U421 ( .A1(n636), .A2(n751), .ZN(n549) );
  NOR2_X1 U422 ( .A1(n754), .A2(n587), .ZN(n588) );
  NOR2_X1 U423 ( .A1(n695), .A2(n375), .ZN(n372) );
  XNOR2_X1 U424 ( .A(n446), .B(n445), .ZN(n536) );
  XNOR2_X1 U425 ( .A(n370), .B(n368), .ZN(n488) );
  XNOR2_X1 U426 ( .A(n487), .B(n486), .ZN(n370) );
  INV_X1 U427 ( .A(n485), .ZN(n368) );
  XNOR2_X1 U428 ( .A(G134), .B(G116), .ZN(n447) );
  XNOR2_X1 U429 ( .A(G143), .B(G140), .ZN(n431) );
  XNOR2_X1 U430 ( .A(G113), .B(KEYINPUT11), .ZN(n435) );
  XNOR2_X1 U431 ( .A(n475), .B(n474), .ZN(n476) );
  NAND2_X1 U432 ( .A1(n399), .A2(n350), .ZN(n357) );
  NOR2_X1 U433 ( .A1(n558), .A2(n397), .ZN(n364) );
  INV_X1 U434 ( .A(n572), .ZN(n363) );
  XNOR2_X1 U435 ( .A(n390), .B(KEYINPUT95), .ZN(n565) );
  XNOR2_X1 U436 ( .A(n396), .B(n393), .ZN(n392) );
  INV_X1 U437 ( .A(n738), .ZN(n391) );
  XNOR2_X1 U438 ( .A(n394), .B(n497), .ZN(n393) );
  XNOR2_X1 U439 ( .A(n415), .B(n416), .ZN(n353) );
  XNOR2_X1 U440 ( .A(n470), .B(n472), .ZN(n415) );
  INV_X1 U441 ( .A(KEYINPUT40), .ZN(n367) );
  XNOR2_X1 U442 ( .A(n597), .B(KEYINPUT112), .ZN(n752) );
  NAND2_X2 U443 ( .A1(n361), .A2(n359), .ZN(n636) );
  AND2_X1 U444 ( .A1(n365), .A2(n362), .ZN(n361) );
  NAND2_X1 U445 ( .A1(n360), .A2(KEYINPUT64), .ZN(n359) );
  NOR2_X1 U446 ( .A1(n364), .A2(n363), .ZN(n362) );
  XNOR2_X1 U447 ( .A(n389), .B(G131), .ZN(G33) );
  INV_X1 U448 ( .A(G122), .ZN(n637) );
  INV_X1 U449 ( .A(n750), .ZN(n388) );
  INV_X1 U450 ( .A(G146), .ZN(n471) );
  OR2_X1 U451 ( .A1(G902), .A2(n720), .ZN(n347) );
  OR2_X1 U452 ( .A1(n590), .A2(n542), .ZN(n348) );
  INV_X1 U453 ( .A(n684), .ZN(n558) );
  AND2_X1 U454 ( .A1(n374), .A2(n373), .ZN(n349) );
  AND2_X1 U455 ( .A1(n611), .A2(n398), .ZN(n350) );
  AND2_X1 U456 ( .A1(n558), .A2(n397), .ZN(n351) );
  XNOR2_X1 U457 ( .A(n494), .B(n493), .ZN(n738) );
  INV_X1 U458 ( .A(KEYINPUT64), .ZN(n397) );
  XNOR2_X2 U459 ( .A(n352), .B(n419), .ZN(n567) );
  NOR2_X1 U460 ( .A1(n354), .A2(n348), .ZN(n658) );
  XNOR2_X2 U461 ( .A(n354), .B(KEYINPUT103), .ZN(n366) );
  NAND2_X2 U462 ( .A1(n503), .A2(n482), .ZN(n354) );
  XNOR2_X2 U463 ( .A(n355), .B(G143), .ZN(n453) );
  INV_X1 U464 ( .A(n567), .ZN(n399) );
  NAND2_X1 U465 ( .A1(n567), .A2(KEYINPUT19), .ZN(n358) );
  INV_X1 U466 ( .A(n366), .ZN(n360) );
  NAND2_X1 U467 ( .A1(n366), .A2(n351), .ZN(n365) );
  NAND2_X1 U468 ( .A1(n349), .A2(n371), .ZN(n377) );
  NAND2_X1 U469 ( .A1(n684), .A2(n372), .ZN(n371) );
  NAND2_X1 U470 ( .A1(n565), .A2(n376), .ZN(n566) );
  AND2_X2 U471 ( .A1(n623), .A2(n621), .ZN(n741) );
  NAND2_X1 U472 ( .A1(n381), .A2(n379), .ZN(n378) );
  AND2_X1 U473 ( .A1(n752), .A2(n380), .ZN(n379) );
  NAND2_X1 U474 ( .A1(n389), .A2(n382), .ZN(n381) );
  XNOR2_X2 U475 ( .A(n385), .B(n384), .ZN(n623) );
  NAND2_X1 U476 ( .A1(n387), .A2(n386), .ZN(n385) );
  NAND2_X1 U477 ( .A1(n533), .A2(n576), .ZN(n390) );
  NAND2_X1 U478 ( .A1(n495), .A2(G221), .ZN(n396) );
  XNOR2_X2 U479 ( .A(n474), .B(G122), .ZN(n432) );
  NAND2_X1 U480 ( .A1(n399), .A2(n611), .ZN(n594) );
  BUF_X1 U481 ( .A(n567), .Z(n614) );
  XNOR2_X1 U482 ( .A(n629), .B(n628), .ZN(n401) );
  AND2_X1 U483 ( .A1(n549), .A2(KEYINPUT44), .ZN(n402) );
  INV_X2 U484 ( .A(G104), .ZN(n474) );
  INV_X1 U485 ( .A(KEYINPUT46), .ZN(n608) );
  XNOR2_X1 U486 ( .A(n477), .B(n476), .ZN(n478) );
  INV_X1 U487 ( .A(KEYINPUT67), .ZN(n516) );
  XNOR2_X1 U488 ( .A(n472), .B(n346), .ZN(n473) );
  XNOR2_X1 U489 ( .A(n468), .B(G134), .ZN(n469) );
  INV_X1 U490 ( .A(KEYINPUT10), .ZN(n433) );
  NOR2_X1 U491 ( .A1(n550), .A2(n402), .ZN(n551) );
  XNOR2_X1 U492 ( .A(n489), .B(n479), .ZN(n629) );
  XNOR2_X1 U493 ( .A(n444), .B(n443), .ZN(n445) );
  NAND2_X1 U494 ( .A1(n552), .A2(n551), .ZN(n553) );
  NOR2_X1 U495 ( .A1(n724), .A2(G902), .ZN(n502) );
  INV_X1 U496 ( .A(n726), .ZN(n632) );
  XNOR2_X1 U497 ( .A(n403), .B(G107), .ZN(n477) );
  XNOR2_X1 U498 ( .A(n432), .B(KEYINPUT16), .ZN(n404) );
  XNOR2_X1 U499 ( .A(n477), .B(n404), .ZN(n408) );
  XNOR2_X1 U500 ( .A(n406), .B(G113), .ZN(n407) );
  XNOR2_X1 U501 ( .A(n434), .B(n409), .ZN(n413) );
  NAND2_X1 U502 ( .A1(n742), .A2(G224), .ZN(n410) );
  XNOR2_X1 U503 ( .A(n411), .B(n410), .ZN(n412) );
  XNOR2_X1 U504 ( .A(n413), .B(n412), .ZN(n416) );
  INV_X1 U505 ( .A(KEYINPUT4), .ZN(n414) );
  XNOR2_X1 U506 ( .A(KEYINPUT15), .B(G902), .ZN(n618) );
  INV_X1 U507 ( .A(G902), .ZN(n418) );
  INV_X1 U508 ( .A(G237), .ZN(n417) );
  NAND2_X1 U509 ( .A1(n418), .A2(n417), .ZN(n420) );
  NAND2_X1 U510 ( .A1(n420), .A2(G210), .ZN(n419) );
  NAND2_X1 U511 ( .A1(n420), .A2(G214), .ZN(n422) );
  INV_X1 U512 ( .A(KEYINPUT89), .ZN(n421) );
  XNOR2_X1 U513 ( .A(n422), .B(n421), .ZN(n611) );
  INV_X1 U514 ( .A(n611), .ZN(n695) );
  NAND2_X1 U515 ( .A1(G234), .A2(G237), .ZN(n423) );
  XNOR2_X1 U516 ( .A(n423), .B(KEYINPUT90), .ZN(n424) );
  XNOR2_X1 U517 ( .A(KEYINPUT14), .B(n424), .ZN(n426) );
  NAND2_X1 U518 ( .A1(G952), .A2(n426), .ZN(n708) );
  NOR2_X1 U519 ( .A1(n708), .A2(G953), .ZN(n563) );
  AND2_X1 U520 ( .A1(G953), .A2(G902), .ZN(n425) );
  NAND2_X1 U521 ( .A1(n426), .A2(n425), .ZN(n559) );
  NOR2_X1 U522 ( .A1(n559), .A2(G898), .ZN(n427) );
  OR2_X1 U523 ( .A1(n563), .A2(n427), .ZN(n428) );
  NAND2_X1 U524 ( .A1(n578), .A2(n428), .ZN(n430) );
  INV_X1 U525 ( .A(KEYINPUT0), .ZN(n429) );
  XNOR2_X1 U526 ( .A(n432), .B(n431), .ZN(n437) );
  XNOR2_X1 U527 ( .A(n494), .B(n435), .ZN(n436) );
  XOR2_X1 U528 ( .A(n437), .B(n436), .Z(n442) );
  XOR2_X1 U529 ( .A(KEYINPUT77), .B(n438), .Z(n483) );
  NAND2_X1 U530 ( .A1(G214), .A2(n483), .ZN(n439) );
  XNOR2_X1 U531 ( .A(n439), .B(KEYINPUT12), .ZN(n440) );
  XNOR2_X1 U532 ( .A(n468), .B(n440), .ZN(n441) );
  XNOR2_X1 U533 ( .A(n442), .B(n441), .ZN(n639) );
  NOR2_X1 U534 ( .A1(G902), .A2(n639), .ZN(n446) );
  XNOR2_X1 U535 ( .A(KEYINPUT97), .B(KEYINPUT13), .ZN(n444) );
  INV_X1 U536 ( .A(G475), .ZN(n443) );
  XOR2_X1 U537 ( .A(G122), .B(G107), .Z(n448) );
  XNOR2_X1 U538 ( .A(n448), .B(n447), .ZN(n452) );
  XOR2_X1 U539 ( .A(KEYINPUT7), .B(KEYINPUT101), .Z(n450) );
  XNOR2_X1 U540 ( .A(KEYINPUT100), .B(KEYINPUT99), .ZN(n449) );
  XNOR2_X1 U541 ( .A(n450), .B(n449), .ZN(n451) );
  XNOR2_X1 U542 ( .A(n452), .B(n451), .ZN(n460) );
  XOR2_X1 U543 ( .A(n453), .B(KEYINPUT9), .Z(n458) );
  NAND2_X1 U544 ( .A1(G234), .A2(n742), .ZN(n454) );
  NAND2_X1 U545 ( .A1(G217), .A2(n495), .ZN(n457) );
  XNOR2_X1 U546 ( .A(n458), .B(n457), .ZN(n459) );
  XNOR2_X1 U547 ( .A(n460), .B(n459), .ZN(n720) );
  XNOR2_X1 U548 ( .A(G478), .B(n347), .ZN(n538) );
  OR2_X1 U549 ( .A1(n536), .A2(n538), .ZN(n602) );
  NAND2_X1 U550 ( .A1(n618), .A2(G234), .ZN(n461) );
  XNOR2_X1 U551 ( .A(n461), .B(KEYINPUT20), .ZN(n498) );
  NAND2_X1 U552 ( .A1(n498), .A2(G221), .ZN(n463) );
  INV_X1 U553 ( .A(KEYINPUT21), .ZN(n462) );
  XNOR2_X1 U554 ( .A(n463), .B(n462), .ZN(n680) );
  INV_X1 U555 ( .A(KEYINPUT94), .ZN(n464) );
  XNOR2_X1 U556 ( .A(n680), .B(n464), .ZN(n515) );
  NOR2_X1 U557 ( .A1(n602), .A2(n515), .ZN(n465) );
  NAND2_X1 U558 ( .A1(n520), .A2(n465), .ZN(n467) );
  INV_X1 U559 ( .A(KEYINPUT22), .ZN(n466) );
  XNOR2_X2 U560 ( .A(n467), .B(n466), .ZN(n503) );
  NAND2_X1 U561 ( .A1(G227), .A2(n742), .ZN(n475) );
  XNOR2_X1 U562 ( .A(n478), .B(n492), .ZN(n479) );
  NOR2_X1 U563 ( .A1(n629), .A2(G902), .ZN(n481) );
  INV_X1 U564 ( .A(G469), .ZN(n480) );
  XNOR2_X2 U565 ( .A(n481), .B(n480), .ZN(n576) );
  XNOR2_X2 U566 ( .A(n576), .B(KEYINPUT1), .ZN(n686) );
  INV_X1 U567 ( .A(n686), .ZN(n482) );
  NAND2_X1 U568 ( .A1(G210), .A2(n483), .ZN(n487) );
  XOR2_X1 U569 ( .A(KEYINPUT96), .B(KEYINPUT5), .Z(n484) );
  XNOR2_X1 U570 ( .A(n484), .B(G137), .ZN(n486) );
  XNOR2_X1 U571 ( .A(n489), .B(n488), .ZN(n650) );
  NOR2_X1 U572 ( .A1(n650), .A2(G902), .ZN(n491) );
  INV_X1 U573 ( .A(G472), .ZN(n490) );
  XNOR2_X2 U574 ( .A(n491), .B(n490), .ZN(n684) );
  INV_X1 U575 ( .A(n492), .ZN(n493) );
  XOR2_X1 U576 ( .A(KEYINPUT92), .B(KEYINPUT23), .Z(n497) );
  XNOR2_X1 U577 ( .A(G128), .B(G110), .ZN(n496) );
  NAND2_X1 U578 ( .A1(G217), .A2(n498), .ZN(n500) );
  XNOR2_X1 U579 ( .A(KEYINPUT93), .B(KEYINPUT25), .ZN(n499) );
  XNOR2_X1 U580 ( .A(n500), .B(n499), .ZN(n501) );
  INV_X1 U581 ( .A(KEYINPUT6), .ZN(n504) );
  INV_X1 U582 ( .A(KEYINPUT102), .ZN(n505) );
  XNOR2_X1 U583 ( .A(n572), .B(n505), .ZN(n681) );
  INV_X1 U584 ( .A(n681), .ZN(n542) );
  NAND2_X1 U585 ( .A1(n542), .A2(n686), .ZN(n506) );
  NOR2_X1 U586 ( .A1(n590), .A2(n506), .ZN(n507) );
  NAND2_X1 U587 ( .A1(n503), .A2(n507), .ZN(n508) );
  XNOR2_X1 U588 ( .A(n508), .B(KEYINPUT32), .ZN(n751) );
  INV_X1 U589 ( .A(n549), .ZN(n511) );
  INV_X1 U590 ( .A(KEYINPUT44), .ZN(n509) );
  AND2_X1 U591 ( .A1(n509), .A2(KEYINPUT84), .ZN(n510) );
  NAND2_X1 U592 ( .A1(n511), .A2(n510), .ZN(n514) );
  INV_X1 U593 ( .A(KEYINPUT84), .ZN(n512) );
  NAND2_X1 U594 ( .A1(n549), .A2(n512), .ZN(n513) );
  NAND2_X1 U595 ( .A1(n514), .A2(n513), .ZN(n528) );
  NAND2_X1 U596 ( .A1(n530), .A2(n590), .ZN(n519) );
  XNOR2_X1 U597 ( .A(KEYINPUT72), .B(KEYINPUT33), .ZN(n518) );
  XNOR2_X2 U598 ( .A(n519), .B(n518), .ZN(n710) );
  NAND2_X1 U599 ( .A1(n710), .A2(n534), .ZN(n522) );
  XNOR2_X1 U600 ( .A(KEYINPUT73), .B(KEYINPUT34), .ZN(n521) );
  XNOR2_X1 U601 ( .A(n522), .B(n521), .ZN(n525) );
  NAND2_X1 U602 ( .A1(n536), .A2(n538), .ZN(n524) );
  INV_X1 U603 ( .A(KEYINPUT104), .ZN(n523) );
  XNOR2_X1 U604 ( .A(n524), .B(n523), .ZN(n557) );
  NAND2_X1 U605 ( .A1(n525), .A2(n557), .ZN(n526) );
  XNOR2_X2 U606 ( .A(n526), .B(KEYINPUT35), .ZN(n529) );
  INV_X1 U607 ( .A(n529), .ZN(n527) );
  NAND2_X1 U608 ( .A1(n528), .A2(n527), .ZN(n552) );
  NAND2_X1 U609 ( .A1(n529), .A2(KEYINPUT44), .ZN(n546) );
  NAND2_X1 U610 ( .A1(n530), .A2(n684), .ZN(n691) );
  NOR2_X1 U611 ( .A1(n691), .A2(n531), .ZN(n532) );
  XNOR2_X1 U612 ( .A(n532), .B(KEYINPUT31), .ZN(n676) );
  AND2_X1 U613 ( .A1(n565), .A2(n558), .ZN(n535) );
  NAND2_X1 U614 ( .A1(n535), .A2(n534), .ZN(n661) );
  NAND2_X1 U615 ( .A1(n676), .A2(n661), .ZN(n541) );
  XOR2_X1 U616 ( .A(KEYINPUT98), .B(n536), .Z(n537) );
  NAND2_X1 U617 ( .A1(n537), .A2(n538), .ZN(n677) );
  INV_X1 U618 ( .A(n537), .ZN(n540) );
  INV_X1 U619 ( .A(n538), .ZN(n539) );
  NAND2_X1 U620 ( .A1(n540), .A2(n539), .ZN(n673) );
  NAND2_X1 U621 ( .A1(n677), .A2(n673), .ZN(n699) );
  XNOR2_X1 U622 ( .A(KEYINPUT80), .B(n699), .ZN(n582) );
  NAND2_X1 U623 ( .A1(n541), .A2(n582), .ZN(n544) );
  INV_X1 U624 ( .A(n658), .ZN(n543) );
  AND2_X1 U625 ( .A1(n544), .A2(n543), .ZN(n545) );
  NAND2_X1 U626 ( .A1(n546), .A2(n545), .ZN(n548) );
  INV_X1 U627 ( .A(KEYINPUT83), .ZN(n547) );
  XNOR2_X1 U628 ( .A(n548), .B(n547), .ZN(n550) );
  XNOR2_X2 U629 ( .A(n553), .B(KEYINPUT45), .ZN(n727) );
  INV_X1 U630 ( .A(n618), .ZN(n554) );
  NAND2_X1 U631 ( .A1(n727), .A2(n554), .ZN(n556) );
  INV_X1 U632 ( .A(KEYINPUT82), .ZN(n555) );
  XNOR2_X1 U633 ( .A(n556), .B(n555), .ZN(n616) );
  INV_X1 U634 ( .A(n557), .ZN(n570) );
  XOR2_X1 U635 ( .A(n559), .B(KEYINPUT105), .Z(n560) );
  NOR2_X1 U636 ( .A1(G900), .A2(n560), .ZN(n561) );
  XNOR2_X1 U637 ( .A(n561), .B(KEYINPUT106), .ZN(n562) );
  NOR2_X1 U638 ( .A1(n563), .A2(n562), .ZN(n574) );
  INV_X1 U639 ( .A(n574), .ZN(n564) );
  XNOR2_X1 U640 ( .A(n566), .B(KEYINPUT78), .ZN(n599) );
  NOR2_X1 U641 ( .A1(n599), .A2(n614), .ZN(n568) );
  XNOR2_X1 U642 ( .A(n568), .B(KEYINPUT109), .ZN(n569) );
  NOR2_X1 U643 ( .A1(n570), .A2(n569), .ZN(n571) );
  XNOR2_X1 U644 ( .A(KEYINPUT110), .B(n571), .ZN(n754) );
  NAND2_X1 U645 ( .A1(n572), .A2(n680), .ZN(n573) );
  NOR2_X1 U646 ( .A1(n574), .A2(n573), .ZN(n589) );
  AND2_X1 U647 ( .A1(n684), .A2(n589), .ZN(n575) );
  XNOR2_X1 U648 ( .A(KEYINPUT28), .B(n575), .ZN(n577) );
  NAND2_X1 U649 ( .A1(n577), .A2(n576), .ZN(n605) );
  INV_X1 U650 ( .A(n578), .ZN(n579) );
  NOR2_X1 U651 ( .A1(n605), .A2(n579), .ZN(n670) );
  NAND2_X1 U652 ( .A1(n670), .A2(n699), .ZN(n580) );
  NAND2_X1 U653 ( .A1(n580), .A2(KEYINPUT47), .ZN(n586) );
  XOR2_X1 U654 ( .A(KEYINPUT68), .B(KEYINPUT47), .Z(n581) );
  NAND2_X1 U655 ( .A1(n582), .A2(n581), .ZN(n583) );
  XNOR2_X1 U656 ( .A(KEYINPUT75), .B(n583), .ZN(n584) );
  NAND2_X1 U657 ( .A1(n584), .A2(n670), .ZN(n585) );
  NAND2_X1 U658 ( .A1(n586), .A2(n585), .ZN(n587) );
  NAND2_X1 U659 ( .A1(n590), .A2(n589), .ZN(n591) );
  XNOR2_X1 U660 ( .A(KEYINPUT107), .B(n591), .ZN(n592) );
  INV_X1 U661 ( .A(n673), .ZN(n671) );
  NAND2_X1 U662 ( .A1(n592), .A2(n671), .ZN(n593) );
  XNOR2_X1 U663 ( .A(KEYINPUT108), .B(n593), .ZN(n610) );
  XNOR2_X1 U664 ( .A(n595), .B(KEYINPUT36), .ZN(n596) );
  NAND2_X1 U665 ( .A1(n596), .A2(n686), .ZN(n597) );
  XOR2_X1 U666 ( .A(KEYINPUT76), .B(KEYINPUT38), .Z(n598) );
  XNOR2_X1 U667 ( .A(n614), .B(n598), .ZN(n696) );
  NOR2_X1 U668 ( .A1(n599), .A2(n696), .ZN(n600) );
  XNOR2_X1 U669 ( .A(n600), .B(KEYINPUT39), .ZN(n609) );
  NOR2_X1 U670 ( .A1(n609), .A2(n673), .ZN(n601) );
  XOR2_X1 U671 ( .A(KEYINPUT111), .B(KEYINPUT41), .Z(n604) );
  NOR2_X1 U672 ( .A1(n695), .A2(n696), .ZN(n700) );
  INV_X1 U673 ( .A(n602), .ZN(n697) );
  NAND2_X1 U674 ( .A1(n700), .A2(n697), .ZN(n603) );
  XNOR2_X1 U675 ( .A(n604), .B(n603), .ZN(n711) );
  INV_X1 U676 ( .A(n605), .ZN(n606) );
  NAND2_X1 U677 ( .A1(n711), .A2(n606), .ZN(n607) );
  XOR2_X1 U678 ( .A(KEYINPUT42), .B(n607), .Z(n750) );
  NOR2_X1 U679 ( .A1(n609), .A2(n677), .ZN(n679) );
  NOR2_X1 U680 ( .A1(n610), .A2(n686), .ZN(n612) );
  NAND2_X1 U681 ( .A1(n612), .A2(n611), .ZN(n613) );
  XNOR2_X1 U682 ( .A(n613), .B(KEYINPUT43), .ZN(n615) );
  AND2_X1 U683 ( .A1(n615), .A2(n614), .ZN(n635) );
  NOR2_X1 U684 ( .A1(n679), .A2(n635), .ZN(n621) );
  NAND2_X1 U685 ( .A1(n616), .A2(n741), .ZN(n620) );
  INV_X1 U686 ( .A(KEYINPUT2), .ZN(n617) );
  OR2_X1 U687 ( .A1(n618), .A2(n617), .ZN(n619) );
  AND2_X1 U688 ( .A1(n621), .A2(n727), .ZN(n622) );
  AND2_X1 U689 ( .A1(n623), .A2(n622), .ZN(n709) );
  NAND2_X1 U690 ( .A1(n709), .A2(KEYINPUT2), .ZN(n624) );
  NAND2_X1 U691 ( .A1(n719), .A2(G469), .ZN(n630) );
  XOR2_X1 U692 ( .A(KEYINPUT122), .B(KEYINPUT121), .Z(n627) );
  XNOR2_X1 U693 ( .A(KEYINPUT57), .B(KEYINPUT58), .ZN(n626) );
  XNOR2_X1 U694 ( .A(n627), .B(n626), .ZN(n628) );
  XNOR2_X1 U695 ( .A(n630), .B(n401), .ZN(n633) );
  INV_X1 U696 ( .A(G952), .ZN(n631) );
  AND2_X1 U697 ( .A1(n631), .A2(G953), .ZN(n726) );
  NAND2_X1 U698 ( .A1(n633), .A2(n632), .ZN(n634) );
  XNOR2_X1 U699 ( .A(n634), .B(KEYINPUT123), .ZN(G54) );
  XOR2_X1 U700 ( .A(n635), .B(G140), .Z(G42) );
  XNOR2_X1 U701 ( .A(n636), .B(G110), .ZN(G12) );
  XNOR2_X1 U702 ( .A(n529), .B(n637), .ZN(G24) );
  NAND2_X1 U703 ( .A1(n719), .A2(G475), .ZN(n641) );
  XNOR2_X1 U704 ( .A(KEYINPUT65), .B(KEYINPUT59), .ZN(n638) );
  XNOR2_X1 U705 ( .A(n639), .B(n638), .ZN(n640) );
  XNOR2_X1 U706 ( .A(n641), .B(n640), .ZN(n642) );
  NOR2_X2 U707 ( .A1(n642), .A2(n726), .ZN(n643) );
  XNOR2_X1 U708 ( .A(n643), .B(KEYINPUT60), .ZN(G60) );
  NAND2_X1 U709 ( .A1(n719), .A2(G210), .ZN(n647) );
  XNOR2_X1 U710 ( .A(KEYINPUT54), .B(KEYINPUT55), .ZN(n644) );
  XNOR2_X1 U711 ( .A(n645), .B(n644), .ZN(n646) );
  XNOR2_X1 U712 ( .A(n647), .B(n646), .ZN(n648) );
  NOR2_X2 U713 ( .A1(n648), .A2(n726), .ZN(n649) );
  XNOR2_X1 U714 ( .A(n649), .B(KEYINPUT56), .ZN(G51) );
  NAND2_X1 U715 ( .A1(n719), .A2(G472), .ZN(n652) );
  XNOR2_X1 U716 ( .A(n650), .B(KEYINPUT62), .ZN(n651) );
  XNOR2_X1 U717 ( .A(n652), .B(n651), .ZN(n653) );
  NOR2_X2 U718 ( .A1(n653), .A2(n726), .ZN(n657) );
  XOR2_X1 U719 ( .A(KEYINPUT85), .B(KEYINPUT113), .Z(n655) );
  XNOR2_X1 U720 ( .A(KEYINPUT86), .B(KEYINPUT63), .ZN(n654) );
  XNOR2_X1 U721 ( .A(n655), .B(n654), .ZN(n656) );
  XNOR2_X1 U722 ( .A(n657), .B(n656), .ZN(G57) );
  XOR2_X1 U723 ( .A(G101), .B(n658), .Z(n659) );
  XNOR2_X1 U724 ( .A(KEYINPUT114), .B(n659), .ZN(G3) );
  NOR2_X1 U725 ( .A1(n673), .A2(n661), .ZN(n660) );
  XOR2_X1 U726 ( .A(G104), .B(n660), .Z(G6) );
  NOR2_X1 U727 ( .A1(n661), .A2(n677), .ZN(n665) );
  XOR2_X1 U728 ( .A(KEYINPUT115), .B(KEYINPUT26), .Z(n663) );
  XNOR2_X1 U729 ( .A(G107), .B(KEYINPUT27), .ZN(n662) );
  XNOR2_X1 U730 ( .A(n663), .B(n662), .ZN(n664) );
  XNOR2_X1 U731 ( .A(n665), .B(n664), .ZN(G9) );
  XOR2_X1 U732 ( .A(KEYINPUT116), .B(KEYINPUT29), .Z(n668) );
  INV_X1 U733 ( .A(n677), .ZN(n666) );
  NAND2_X1 U734 ( .A1(n666), .A2(n670), .ZN(n667) );
  XNOR2_X1 U735 ( .A(n668), .B(n667), .ZN(n669) );
  XNOR2_X1 U736 ( .A(G128), .B(n669), .ZN(G30) );
  NAND2_X1 U737 ( .A1(n671), .A2(n670), .ZN(n672) );
  XNOR2_X1 U738 ( .A(n672), .B(n346), .ZN(G48) );
  NOR2_X1 U739 ( .A1(n673), .A2(n676), .ZN(n675) );
  XNOR2_X1 U740 ( .A(G113), .B(KEYINPUT117), .ZN(n674) );
  XNOR2_X1 U741 ( .A(n675), .B(n674), .ZN(G15) );
  NOR2_X1 U742 ( .A1(n677), .A2(n676), .ZN(n678) );
  XOR2_X1 U743 ( .A(G116), .B(n678), .Z(G18) );
  XOR2_X1 U744 ( .A(G134), .B(n679), .Z(G36) );
  XOR2_X1 U745 ( .A(KEYINPUT120), .B(KEYINPUT53), .Z(n718) );
  NOR2_X1 U746 ( .A1(n681), .A2(n680), .ZN(n682) );
  XOR2_X1 U747 ( .A(KEYINPUT49), .B(n682), .Z(n683) );
  NOR2_X1 U748 ( .A1(n684), .A2(n683), .ZN(n685) );
  XOR2_X1 U749 ( .A(KEYINPUT118), .B(n685), .Z(n689) );
  NOR2_X1 U750 ( .A1(n533), .A2(n686), .ZN(n687) );
  XNOR2_X1 U751 ( .A(KEYINPUT50), .B(n687), .ZN(n688) );
  NOR2_X1 U752 ( .A1(n689), .A2(n688), .ZN(n690) );
  XNOR2_X1 U753 ( .A(n690), .B(KEYINPUT119), .ZN(n692) );
  NAND2_X1 U754 ( .A1(n692), .A2(n691), .ZN(n693) );
  XOR2_X1 U755 ( .A(KEYINPUT51), .B(n693), .Z(n694) );
  NAND2_X1 U756 ( .A1(n711), .A2(n694), .ZN(n705) );
  NAND2_X1 U757 ( .A1(n696), .A2(n695), .ZN(n698) );
  NAND2_X1 U758 ( .A1(n698), .A2(n697), .ZN(n702) );
  NAND2_X1 U759 ( .A1(n700), .A2(n699), .ZN(n701) );
  NAND2_X1 U760 ( .A1(n702), .A2(n701), .ZN(n703) );
  NAND2_X1 U761 ( .A1(n703), .A2(n710), .ZN(n704) );
  NAND2_X1 U762 ( .A1(n705), .A2(n704), .ZN(n706) );
  XOR2_X1 U763 ( .A(KEYINPUT52), .B(n706), .Z(n707) );
  NOR2_X1 U764 ( .A1(n708), .A2(n707), .ZN(n715) );
  XNOR2_X1 U765 ( .A(n709), .B(KEYINPUT2), .ZN(n713) );
  NAND2_X1 U766 ( .A1(n711), .A2(n710), .ZN(n712) );
  NAND2_X1 U767 ( .A1(n713), .A2(n712), .ZN(n714) );
  NOR2_X1 U768 ( .A1(n715), .A2(n714), .ZN(n716) );
  NAND2_X1 U769 ( .A1(n716), .A2(n742), .ZN(n717) );
  XNOR2_X1 U770 ( .A(n718), .B(n717), .ZN(G75) );
  NAND2_X1 U771 ( .A1(n719), .A2(G478), .ZN(n721) );
  XNOR2_X1 U772 ( .A(n721), .B(n720), .ZN(n722) );
  NOR2_X1 U773 ( .A1(n726), .A2(n722), .ZN(G63) );
  NAND2_X1 U774 ( .A1(n719), .A2(G217), .ZN(n723) );
  XNOR2_X1 U775 ( .A(n724), .B(n723), .ZN(n725) );
  NOR2_X1 U776 ( .A1(n726), .A2(n725), .ZN(G66) );
  NAND2_X1 U777 ( .A1(n727), .A2(n742), .ZN(n731) );
  NAND2_X1 U778 ( .A1(G953), .A2(G224), .ZN(n728) );
  XNOR2_X1 U779 ( .A(KEYINPUT61), .B(n728), .ZN(n729) );
  NAND2_X1 U780 ( .A1(n729), .A2(G898), .ZN(n730) );
  NAND2_X1 U781 ( .A1(n731), .A2(n730), .ZN(n737) );
  XNOR2_X1 U782 ( .A(G101), .B(KEYINPUT124), .ZN(n732) );
  XNOR2_X1 U783 ( .A(n733), .B(n732), .ZN(n735) );
  NOR2_X1 U784 ( .A1(G898), .A2(n742), .ZN(n734) );
  NOR2_X1 U785 ( .A1(n735), .A2(n734), .ZN(n736) );
  XNOR2_X1 U786 ( .A(n737), .B(n736), .ZN(G69) );
  XOR2_X1 U787 ( .A(n738), .B(n739), .Z(n740) );
  XNOR2_X1 U788 ( .A(KEYINPUT125), .B(n740), .ZN(n744) );
  XOR2_X1 U789 ( .A(n744), .B(n741), .Z(n743) );
  NAND2_X1 U790 ( .A1(n743), .A2(n742), .ZN(n748) );
  XNOR2_X1 U791 ( .A(G227), .B(n744), .ZN(n745) );
  NAND2_X1 U792 ( .A1(n745), .A2(G900), .ZN(n746) );
  NAND2_X1 U793 ( .A1(G953), .A2(n746), .ZN(n747) );
  NAND2_X1 U794 ( .A1(n748), .A2(n747), .ZN(G72) );
  XOR2_X1 U795 ( .A(G137), .B(KEYINPUT126), .Z(n749) );
  XNOR2_X1 U796 ( .A(n750), .B(n749), .ZN(G39) );
  XNOR2_X1 U797 ( .A(G119), .B(n751), .ZN(G21) );
  XOR2_X1 U798 ( .A(G125), .B(n752), .Z(n753) );
  XNOR2_X1 U799 ( .A(KEYINPUT37), .B(n753), .ZN(G27) );
  XOR2_X1 U800 ( .A(G143), .B(n754), .Z(G45) );
endmodule

