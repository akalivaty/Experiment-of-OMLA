//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 0 0 1 0 1 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 1 0 0 0 0 0 1 0 0 0 0 1 1 1 0 0 0 1 1 1 1 1 0 0 1 1 0 1 1 1 1 0 0 1 1 1 1 1 0 0 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:27:31 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n710,
    new_n711, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n721, new_n722, new_n724, new_n725, new_n726, new_n728,
    new_n729, new_n730, new_n731, new_n732, new_n733, new_n734, new_n735,
    new_n736, new_n737, new_n739, new_n740, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n750, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n774, new_n775,
    new_n776, new_n777, new_n778, new_n779, new_n780, new_n781, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n906, new_n907, new_n908, new_n909, new_n910,
    new_n911, new_n912, new_n913, new_n914, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n934,
    new_n935, new_n936, new_n937, new_n938, new_n939, new_n940, new_n941,
    new_n943, new_n944, new_n945, new_n946, new_n947, new_n948, new_n949,
    new_n950, new_n951, new_n952, new_n953, new_n954, new_n955, new_n956,
    new_n957, new_n959, new_n960, new_n961, new_n962, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012;
  OAI21_X1  g000(.A(G214), .B1(G237), .B2(G902), .ZN(new_n187));
  OAI21_X1  g001(.A(G210), .B1(G237), .B2(G902), .ZN(new_n188));
  INV_X1    g002(.A(KEYINPUT3), .ZN(new_n189));
  NAND2_X1  g003(.A1(new_n189), .A2(G104), .ZN(new_n190));
  AND2_X1   g004(.A1(KEYINPUT79), .A2(G107), .ZN(new_n191));
  NOR2_X1   g005(.A1(KEYINPUT79), .A2(G107), .ZN(new_n192));
  NOR3_X1   g006(.A1(new_n190), .A2(new_n191), .A3(new_n192), .ZN(new_n193));
  INV_X1    g007(.A(G104), .ZN(new_n194));
  AOI21_X1  g008(.A(G107), .B1(new_n194), .B2(KEYINPUT3), .ZN(new_n195));
  NOR2_X1   g009(.A1(new_n194), .A2(KEYINPUT3), .ZN(new_n196));
  NOR2_X1   g010(.A1(new_n195), .A2(new_n196), .ZN(new_n197));
  OAI21_X1  g011(.A(G101), .B1(new_n193), .B2(new_n197), .ZN(new_n198));
  OR2_X1    g012(.A1(KEYINPUT79), .A2(G107), .ZN(new_n199));
  NAND2_X1  g013(.A1(KEYINPUT79), .A2(G107), .ZN(new_n200));
  NAND3_X1  g014(.A1(new_n196), .A2(new_n199), .A3(new_n200), .ZN(new_n201));
  INV_X1    g015(.A(G107), .ZN(new_n202));
  OAI21_X1  g016(.A(new_n202), .B1(new_n189), .B2(G104), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n203), .A2(new_n190), .ZN(new_n204));
  INV_X1    g018(.A(G101), .ZN(new_n205));
  NAND3_X1  g019(.A1(new_n201), .A2(new_n204), .A3(new_n205), .ZN(new_n206));
  NAND3_X1  g020(.A1(new_n198), .A2(KEYINPUT4), .A3(new_n206), .ZN(new_n207));
  XNOR2_X1  g021(.A(G116), .B(G119), .ZN(new_n208));
  INV_X1    g022(.A(new_n208), .ZN(new_n209));
  XNOR2_X1  g023(.A(KEYINPUT2), .B(G113), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  INV_X1    g025(.A(new_n210), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n212), .A2(new_n208), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n211), .A2(new_n213), .ZN(new_n214));
  INV_X1    g028(.A(KEYINPUT4), .ZN(new_n215));
  OAI211_X1 g029(.A(new_n215), .B(G101), .C1(new_n193), .C2(new_n197), .ZN(new_n216));
  NAND3_X1  g030(.A1(new_n207), .A2(new_n214), .A3(new_n216), .ZN(new_n217));
  AOI21_X1  g031(.A(new_n205), .B1(G104), .B2(G107), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n199), .A2(new_n200), .ZN(new_n219));
  OAI21_X1  g033(.A(new_n218), .B1(new_n219), .B2(G104), .ZN(new_n220));
  AND2_X1   g034(.A1(new_n206), .A2(new_n220), .ZN(new_n221));
  INV_X1    g035(.A(KEYINPUT5), .ZN(new_n222));
  INV_X1    g036(.A(G119), .ZN(new_n223));
  NAND3_X1  g037(.A1(new_n222), .A2(new_n223), .A3(G116), .ZN(new_n224));
  OAI211_X1 g038(.A(G113), .B(new_n224), .C1(new_n209), .C2(new_n222), .ZN(new_n225));
  NAND3_X1  g039(.A1(new_n221), .A2(new_n213), .A3(new_n225), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n217), .A2(new_n226), .ZN(new_n227));
  XNOR2_X1  g041(.A(G110), .B(G122), .ZN(new_n228));
  INV_X1    g042(.A(new_n228), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n227), .A2(new_n229), .ZN(new_n230));
  NAND3_X1  g044(.A1(new_n217), .A2(new_n226), .A3(new_n228), .ZN(new_n231));
  NAND3_X1  g045(.A1(new_n230), .A2(KEYINPUT6), .A3(new_n231), .ZN(new_n232));
  XNOR2_X1  g046(.A(KEYINPUT83), .B(G224), .ZN(new_n233));
  INV_X1    g047(.A(G953), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n233), .A2(new_n234), .ZN(new_n235));
  XOR2_X1   g049(.A(new_n235), .B(KEYINPUT82), .Z(new_n236));
  INV_X1    g050(.A(new_n236), .ZN(new_n237));
  INV_X1    g051(.A(G125), .ZN(new_n238));
  AND2_X1   g052(.A1(KEYINPUT0), .A2(G128), .ZN(new_n239));
  NOR2_X1   g053(.A1(KEYINPUT0), .A2(G128), .ZN(new_n240));
  NOR2_X1   g054(.A1(new_n239), .A2(new_n240), .ZN(new_n241));
  INV_X1    g055(.A(G146), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n242), .A2(KEYINPUT64), .ZN(new_n243));
  INV_X1    g057(.A(KEYINPUT64), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n244), .A2(G146), .ZN(new_n245));
  AOI21_X1  g059(.A(G143), .B1(new_n243), .B2(new_n245), .ZN(new_n246));
  INV_X1    g060(.A(G143), .ZN(new_n247));
  NOR2_X1   g061(.A1(new_n247), .A2(G146), .ZN(new_n248));
  OAI21_X1  g062(.A(new_n241), .B1(new_n246), .B2(new_n248), .ZN(new_n249));
  INV_X1    g063(.A(KEYINPUT65), .ZN(new_n250));
  NOR2_X1   g064(.A1(new_n242), .A2(G143), .ZN(new_n251));
  XNOR2_X1  g065(.A(KEYINPUT64), .B(G146), .ZN(new_n252));
  AOI21_X1  g066(.A(new_n251), .B1(new_n252), .B2(G143), .ZN(new_n253));
  AOI22_X1  g067(.A1(new_n249), .A2(new_n250), .B1(new_n239), .B2(new_n253), .ZN(new_n254));
  OAI211_X1 g068(.A(KEYINPUT65), .B(new_n241), .C1(new_n246), .C2(new_n248), .ZN(new_n255));
  AOI21_X1  g069(.A(new_n238), .B1(new_n254), .B2(new_n255), .ZN(new_n256));
  NAND3_X1  g070(.A1(new_n243), .A2(new_n245), .A3(G143), .ZN(new_n257));
  INV_X1    g071(.A(new_n251), .ZN(new_n258));
  INV_X1    g072(.A(G128), .ZN(new_n259));
  NOR2_X1   g073(.A1(new_n259), .A2(KEYINPUT1), .ZN(new_n260));
  NAND3_X1  g074(.A1(new_n257), .A2(new_n258), .A3(new_n260), .ZN(new_n261));
  AOI21_X1  g075(.A(new_n259), .B1(new_n257), .B2(KEYINPUT1), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n243), .A2(new_n245), .ZN(new_n263));
  AOI21_X1  g077(.A(new_n248), .B1(new_n263), .B2(new_n247), .ZN(new_n264));
  OAI211_X1 g078(.A(new_n238), .B(new_n261), .C1(new_n262), .C2(new_n264), .ZN(new_n265));
  INV_X1    g079(.A(new_n265), .ZN(new_n266));
  OAI21_X1  g080(.A(new_n237), .B1(new_n256), .B2(new_n266), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n249), .A2(new_n250), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n253), .A2(new_n239), .ZN(new_n269));
  NAND3_X1  g083(.A1(new_n268), .A2(new_n255), .A3(new_n269), .ZN(new_n270));
  NAND2_X1  g084(.A1(new_n270), .A2(G125), .ZN(new_n271));
  NAND3_X1  g085(.A1(new_n271), .A2(new_n265), .A3(new_n236), .ZN(new_n272));
  NAND2_X1  g086(.A1(new_n267), .A2(new_n272), .ZN(new_n273));
  INV_X1    g087(.A(KEYINPUT6), .ZN(new_n274));
  NAND3_X1  g088(.A1(new_n227), .A2(new_n274), .A3(new_n229), .ZN(new_n275));
  NAND3_X1  g089(.A1(new_n232), .A2(new_n273), .A3(new_n275), .ZN(new_n276));
  INV_X1    g090(.A(KEYINPUT84), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n276), .A2(new_n277), .ZN(new_n278));
  NAND4_X1  g092(.A1(new_n232), .A2(KEYINPUT84), .A3(new_n273), .A4(new_n275), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n278), .A2(new_n279), .ZN(new_n280));
  INV_X1    g094(.A(G902), .ZN(new_n281));
  NAND4_X1  g095(.A1(new_n271), .A2(KEYINPUT7), .A3(new_n265), .A4(new_n235), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n235), .A2(KEYINPUT7), .ZN(new_n283));
  OAI21_X1  g097(.A(new_n283), .B1(new_n256), .B2(new_n266), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n282), .A2(new_n284), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n225), .A2(new_n213), .ZN(new_n286));
  NAND2_X1  g100(.A1(new_n206), .A2(new_n220), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n286), .A2(new_n287), .ZN(new_n288));
  AND2_X1   g102(.A1(new_n226), .A2(new_n288), .ZN(new_n289));
  XOR2_X1   g103(.A(new_n228), .B(KEYINPUT8), .Z(new_n290));
  OAI21_X1  g104(.A(new_n231), .B1(new_n289), .B2(new_n290), .ZN(new_n291));
  OAI21_X1  g105(.A(new_n281), .B1(new_n285), .B2(new_n291), .ZN(new_n292));
  INV_X1    g106(.A(new_n292), .ZN(new_n293));
  AOI21_X1  g107(.A(new_n188), .B1(new_n280), .B2(new_n293), .ZN(new_n294));
  INV_X1    g108(.A(new_n188), .ZN(new_n295));
  AOI211_X1 g109(.A(new_n295), .B(new_n292), .C1(new_n278), .C2(new_n279), .ZN(new_n296));
  OAI21_X1  g110(.A(new_n187), .B1(new_n294), .B2(new_n296), .ZN(new_n297));
  XNOR2_X1  g111(.A(KEYINPUT9), .B(G234), .ZN(new_n298));
  OAI21_X1  g112(.A(G221), .B1(new_n298), .B2(G902), .ZN(new_n299));
  XNOR2_X1  g113(.A(new_n299), .B(KEYINPUT78), .ZN(new_n300));
  INV_X1    g114(.A(new_n300), .ZN(new_n301));
  INV_X1    g115(.A(G469), .ZN(new_n302));
  XOR2_X1   g116(.A(KEYINPUT70), .B(G902), .Z(new_n303));
  XNOR2_X1  g117(.A(G110), .B(G140), .ZN(new_n304));
  INV_X1    g118(.A(G227), .ZN(new_n305));
  NOR2_X1   g119(.A1(new_n305), .A2(G953), .ZN(new_n306));
  XNOR2_X1  g120(.A(new_n304), .B(new_n306), .ZN(new_n307));
  AND3_X1   g121(.A1(new_n257), .A2(new_n258), .A3(new_n260), .ZN(new_n308));
  OAI21_X1  g122(.A(KEYINPUT1), .B1(new_n247), .B2(G146), .ZN(new_n309));
  AOI22_X1  g123(.A1(new_n257), .A2(new_n258), .B1(G128), .B2(new_n309), .ZN(new_n310));
  OAI211_X1 g124(.A(new_n206), .B(new_n220), .C1(new_n308), .C2(new_n310), .ZN(new_n311));
  INV_X1    g125(.A(KEYINPUT10), .ZN(new_n312));
  AND3_X1   g126(.A1(new_n206), .A2(KEYINPUT10), .A3(new_n220), .ZN(new_n313));
  OAI21_X1  g127(.A(new_n261), .B1(new_n262), .B2(new_n264), .ZN(new_n314));
  AOI22_X1  g128(.A1(new_n311), .A2(new_n312), .B1(new_n313), .B2(new_n314), .ZN(new_n315));
  INV_X1    g129(.A(G134), .ZN(new_n316));
  OAI21_X1  g130(.A(KEYINPUT11), .B1(new_n316), .B2(G137), .ZN(new_n317));
  INV_X1    g131(.A(KEYINPUT11), .ZN(new_n318));
  INV_X1    g132(.A(G137), .ZN(new_n319));
  NAND3_X1  g133(.A1(new_n318), .A2(new_n319), .A3(G134), .ZN(new_n320));
  AND2_X1   g134(.A1(new_n317), .A2(new_n320), .ZN(new_n321));
  OAI21_X1  g135(.A(KEYINPUT66), .B1(new_n319), .B2(G134), .ZN(new_n322));
  INV_X1    g136(.A(KEYINPUT66), .ZN(new_n323));
  NAND3_X1  g137(.A1(new_n323), .A2(new_n316), .A3(G137), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n322), .A2(new_n324), .ZN(new_n325));
  OAI21_X1  g139(.A(G131), .B1(new_n321), .B2(new_n325), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n317), .A2(new_n320), .ZN(new_n327));
  INV_X1    g141(.A(G131), .ZN(new_n328));
  NAND4_X1  g142(.A1(new_n327), .A2(new_n328), .A3(new_n322), .A4(new_n324), .ZN(new_n329));
  AND2_X1   g143(.A1(new_n326), .A2(new_n329), .ZN(new_n330));
  NAND4_X1  g144(.A1(new_n254), .A2(new_n207), .A3(new_n255), .A4(new_n216), .ZN(new_n331));
  AND3_X1   g145(.A1(new_n315), .A2(new_n330), .A3(new_n331), .ZN(new_n332));
  AOI21_X1  g146(.A(new_n330), .B1(new_n315), .B2(new_n331), .ZN(new_n333));
  OAI211_X1 g147(.A(KEYINPUT81), .B(new_n307), .C1(new_n332), .C2(new_n333), .ZN(new_n334));
  INV_X1    g148(.A(new_n307), .ZN(new_n335));
  NAND3_X1  g149(.A1(new_n315), .A2(new_n330), .A3(new_n331), .ZN(new_n336));
  OAI21_X1  g150(.A(new_n311), .B1(new_n314), .B2(new_n221), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n326), .A2(new_n329), .ZN(new_n338));
  AND3_X1   g152(.A1(new_n337), .A2(KEYINPUT12), .A3(new_n338), .ZN(new_n339));
  AOI21_X1  g153(.A(KEYINPUT12), .B1(new_n337), .B2(new_n338), .ZN(new_n340));
  OAI211_X1 g154(.A(new_n335), .B(new_n336), .C1(new_n339), .C2(new_n340), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n334), .A2(new_n341), .ZN(new_n342));
  NOR2_X1   g156(.A1(new_n308), .A2(new_n310), .ZN(new_n343));
  OAI21_X1  g157(.A(new_n312), .B1(new_n343), .B2(new_n287), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n313), .A2(new_n314), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n207), .A2(new_n216), .ZN(new_n346));
  OAI211_X1 g160(.A(new_n344), .B(new_n345), .C1(new_n346), .C2(new_n270), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n347), .A2(new_n338), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n348), .A2(new_n336), .ZN(new_n349));
  AOI21_X1  g163(.A(KEYINPUT81), .B1(new_n349), .B2(new_n307), .ZN(new_n350));
  OAI211_X1 g164(.A(new_n302), .B(new_n303), .C1(new_n342), .C2(new_n350), .ZN(new_n351));
  INV_X1    g165(.A(new_n351), .ZN(new_n352));
  OAI21_X1  g166(.A(new_n336), .B1(new_n339), .B2(new_n340), .ZN(new_n353));
  NAND2_X1  g167(.A1(new_n353), .A2(new_n307), .ZN(new_n354));
  INV_X1    g168(.A(KEYINPUT80), .ZN(new_n355));
  AOI21_X1  g169(.A(new_n355), .B1(new_n336), .B2(new_n335), .ZN(new_n356));
  NAND3_X1  g170(.A1(new_n336), .A2(new_n355), .A3(new_n335), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n357), .A2(new_n348), .ZN(new_n358));
  OAI211_X1 g172(.A(new_n354), .B(G469), .C1(new_n356), .C2(new_n358), .ZN(new_n359));
  NOR2_X1   g173(.A1(new_n302), .A2(new_n281), .ZN(new_n360));
  INV_X1    g174(.A(new_n360), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n359), .A2(new_n361), .ZN(new_n362));
  OAI21_X1  g176(.A(new_n301), .B1(new_n352), .B2(new_n362), .ZN(new_n363));
  INV_X1    g177(.A(G475), .ZN(new_n364));
  XNOR2_X1  g178(.A(G113), .B(G122), .ZN(new_n365));
  XNOR2_X1  g179(.A(new_n365), .B(new_n194), .ZN(new_n366));
  NAND2_X1  g180(.A1(KEYINPUT18), .A2(G131), .ZN(new_n367));
  INV_X1    g181(.A(G237), .ZN(new_n368));
  NAND3_X1  g182(.A1(new_n368), .A2(new_n234), .A3(G214), .ZN(new_n369));
  INV_X1    g183(.A(KEYINPUT85), .ZN(new_n370));
  AOI21_X1  g184(.A(G143), .B1(new_n369), .B2(new_n370), .ZN(new_n371));
  INV_X1    g185(.A(KEYINPUT86), .ZN(new_n372));
  NAND4_X1  g186(.A1(new_n368), .A2(new_n234), .A3(KEYINPUT85), .A4(G214), .ZN(new_n373));
  AND3_X1   g187(.A1(new_n371), .A2(new_n372), .A3(new_n373), .ZN(new_n374));
  NAND4_X1  g188(.A1(new_n368), .A2(new_n234), .A3(G143), .A4(G214), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n375), .A2(KEYINPUT86), .ZN(new_n376));
  AOI21_X1  g190(.A(new_n376), .B1(new_n371), .B2(new_n373), .ZN(new_n377));
  OAI21_X1  g191(.A(new_n367), .B1(new_n374), .B2(new_n377), .ZN(new_n378));
  INV_X1    g192(.A(G140), .ZN(new_n379));
  AND3_X1   g193(.A1(new_n379), .A2(KEYINPUT72), .A3(G125), .ZN(new_n380));
  XNOR2_X1  g194(.A(G125), .B(G140), .ZN(new_n381));
  INV_X1    g195(.A(KEYINPUT72), .ZN(new_n382));
  AOI21_X1  g196(.A(new_n380), .B1(new_n381), .B2(new_n382), .ZN(new_n383));
  NAND2_X1  g197(.A1(new_n383), .A2(G146), .ZN(new_n384));
  INV_X1    g198(.A(new_n381), .ZN(new_n385));
  OAI21_X1  g199(.A(new_n384), .B1(new_n263), .B2(new_n385), .ZN(new_n386));
  NAND2_X1  g200(.A1(new_n369), .A2(new_n370), .ZN(new_n387));
  NAND3_X1  g201(.A1(new_n387), .A2(new_n247), .A3(new_n373), .ZN(new_n388));
  INV_X1    g202(.A(new_n376), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n388), .A2(new_n389), .ZN(new_n390));
  NAND3_X1  g204(.A1(new_n371), .A2(new_n372), .A3(new_n373), .ZN(new_n391));
  NAND3_X1  g205(.A1(new_n390), .A2(G131), .A3(new_n391), .ZN(new_n392));
  INV_X1    g206(.A(KEYINPUT18), .ZN(new_n393));
  OAI211_X1 g207(.A(new_n378), .B(new_n386), .C1(new_n392), .C2(new_n393), .ZN(new_n394));
  OAI21_X1  g208(.A(new_n328), .B1(new_n374), .B2(new_n377), .ZN(new_n395));
  INV_X1    g209(.A(KEYINPUT17), .ZN(new_n396));
  AND3_X1   g210(.A1(new_n395), .A2(new_n396), .A3(new_n392), .ZN(new_n397));
  NAND4_X1  g211(.A1(new_n390), .A2(KEYINPUT17), .A3(G131), .A4(new_n391), .ZN(new_n398));
  AOI21_X1  g212(.A(KEYINPUT16), .B1(new_n379), .B2(G125), .ZN(new_n399));
  AOI21_X1  g213(.A(new_n399), .B1(new_n383), .B2(KEYINPUT16), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n400), .A2(new_n242), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n379), .A2(G125), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n238), .A2(G140), .ZN(new_n403));
  NAND3_X1  g217(.A1(new_n402), .A2(new_n403), .A3(new_n382), .ZN(new_n404));
  NAND3_X1  g218(.A1(new_n379), .A2(KEYINPUT72), .A3(G125), .ZN(new_n405));
  NAND3_X1  g219(.A1(new_n404), .A2(KEYINPUT16), .A3(new_n405), .ZN(new_n406));
  INV_X1    g220(.A(new_n399), .ZN(new_n407));
  AOI21_X1  g221(.A(new_n242), .B1(new_n406), .B2(new_n407), .ZN(new_n408));
  INV_X1    g222(.A(new_n408), .ZN(new_n409));
  NAND3_X1  g223(.A1(new_n398), .A2(new_n401), .A3(new_n409), .ZN(new_n410));
  OAI211_X1 g224(.A(new_n366), .B(new_n394), .C1(new_n397), .C2(new_n410), .ZN(new_n411));
  INV_X1    g225(.A(new_n411), .ZN(new_n412));
  NAND3_X1  g226(.A1(new_n395), .A2(new_n396), .A3(new_n392), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n406), .A2(new_n407), .ZN(new_n414));
  NOR2_X1   g228(.A1(new_n414), .A2(G146), .ZN(new_n415));
  NOR2_X1   g229(.A1(new_n415), .A2(new_n408), .ZN(new_n416));
  NAND3_X1  g230(.A1(new_n413), .A2(new_n416), .A3(new_n398), .ZN(new_n417));
  AOI21_X1  g231(.A(new_n366), .B1(new_n417), .B2(new_n394), .ZN(new_n418));
  OAI21_X1  g232(.A(new_n281), .B1(new_n412), .B2(new_n418), .ZN(new_n419));
  AOI21_X1  g233(.A(new_n364), .B1(new_n419), .B2(KEYINPUT89), .ZN(new_n420));
  INV_X1    g234(.A(KEYINPUT89), .ZN(new_n421));
  OAI211_X1 g235(.A(new_n421), .B(new_n281), .C1(new_n412), .C2(new_n418), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n420), .A2(new_n422), .ZN(new_n423));
  NOR2_X1   g237(.A1(G475), .A2(G902), .ZN(new_n424));
  NOR3_X1   g238(.A1(new_n374), .A2(new_n377), .A3(new_n328), .ZN(new_n425));
  AOI21_X1  g239(.A(G131), .B1(new_n390), .B2(new_n391), .ZN(new_n426));
  OAI21_X1  g240(.A(KEYINPUT87), .B1(new_n425), .B2(new_n426), .ZN(new_n427));
  INV_X1    g241(.A(KEYINPUT73), .ZN(new_n428));
  AOI21_X1  g242(.A(new_n428), .B1(new_n414), .B2(G146), .ZN(new_n429));
  AOI211_X1 g243(.A(KEYINPUT73), .B(new_n242), .C1(new_n406), .C2(new_n407), .ZN(new_n430));
  NOR2_X1   g244(.A1(new_n429), .A2(new_n430), .ZN(new_n431));
  NAND3_X1  g245(.A1(new_n383), .A2(KEYINPUT88), .A3(KEYINPUT19), .ZN(new_n432));
  AND2_X1   g246(.A1(new_n383), .A2(KEYINPUT19), .ZN(new_n433));
  INV_X1    g247(.A(KEYINPUT88), .ZN(new_n434));
  OAI21_X1  g248(.A(new_n434), .B1(new_n385), .B2(KEYINPUT19), .ZN(new_n435));
  OAI21_X1  g249(.A(new_n432), .B1(new_n433), .B2(new_n435), .ZN(new_n436));
  NAND2_X1  g250(.A1(new_n436), .A2(new_n252), .ZN(new_n437));
  INV_X1    g251(.A(KEYINPUT87), .ZN(new_n438));
  NAND3_X1  g252(.A1(new_n395), .A2(new_n438), .A3(new_n392), .ZN(new_n439));
  NAND4_X1  g253(.A1(new_n427), .A2(new_n431), .A3(new_n437), .A4(new_n439), .ZN(new_n440));
  AOI21_X1  g254(.A(new_n366), .B1(new_n440), .B2(new_n394), .ZN(new_n441));
  OAI21_X1  g255(.A(new_n424), .B1(new_n441), .B2(new_n412), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n442), .A2(KEYINPUT20), .ZN(new_n443));
  INV_X1    g257(.A(KEYINPUT20), .ZN(new_n444));
  OAI211_X1 g258(.A(new_n444), .B(new_n424), .C1(new_n441), .C2(new_n412), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n443), .A2(new_n445), .ZN(new_n446));
  XNOR2_X1  g260(.A(G116), .B(G122), .ZN(new_n447));
  INV_X1    g261(.A(KEYINPUT14), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n447), .A2(new_n448), .ZN(new_n449));
  INV_X1    g263(.A(G122), .ZN(new_n450));
  NOR2_X1   g264(.A1(new_n450), .A2(G116), .ZN(new_n451));
  AOI21_X1  g265(.A(new_n202), .B1(new_n451), .B2(KEYINPUT14), .ZN(new_n452));
  NOR2_X1   g266(.A1(new_n191), .A2(new_n192), .ZN(new_n453));
  AOI22_X1  g267(.A1(new_n449), .A2(new_n452), .B1(new_n453), .B2(new_n447), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n247), .A2(G128), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n259), .A2(G143), .ZN(new_n456));
  AND3_X1   g270(.A1(new_n455), .A2(new_n456), .A3(new_n316), .ZN(new_n457));
  AOI21_X1  g271(.A(new_n316), .B1(new_n455), .B2(new_n456), .ZN(new_n458));
  INV_X1    g272(.A(KEYINPUT90), .ZN(new_n459));
  NOR3_X1   g273(.A1(new_n457), .A2(new_n458), .A3(new_n459), .ZN(new_n460));
  NOR2_X1   g274(.A1(new_n259), .A2(G143), .ZN(new_n461));
  NOR2_X1   g275(.A1(new_n247), .A2(G128), .ZN(new_n462));
  OAI21_X1  g276(.A(G134), .B1(new_n461), .B2(new_n462), .ZN(new_n463));
  NAND3_X1  g277(.A1(new_n455), .A2(new_n456), .A3(new_n316), .ZN(new_n464));
  AOI21_X1  g278(.A(KEYINPUT90), .B1(new_n463), .B2(new_n464), .ZN(new_n465));
  OAI21_X1  g279(.A(new_n454), .B1(new_n460), .B2(new_n465), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n450), .A2(G116), .ZN(new_n467));
  INV_X1    g281(.A(G116), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n468), .A2(G122), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n467), .A2(new_n469), .ZN(new_n470));
  NAND2_X1  g284(.A1(new_n219), .A2(new_n470), .ZN(new_n471));
  NAND2_X1  g285(.A1(new_n453), .A2(new_n447), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n471), .A2(new_n472), .ZN(new_n473));
  INV_X1    g287(.A(KEYINPUT13), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n455), .A2(new_n474), .ZN(new_n475));
  NAND3_X1  g289(.A1(new_n247), .A2(KEYINPUT13), .A3(G128), .ZN(new_n476));
  NAND3_X1  g290(.A1(new_n475), .A2(new_n476), .A3(new_n456), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n477), .A2(G134), .ZN(new_n478));
  NAND3_X1  g292(.A1(new_n473), .A2(new_n478), .A3(new_n464), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n234), .A2(G217), .ZN(new_n480));
  NOR2_X1   g294(.A1(new_n298), .A2(new_n480), .ZN(new_n481));
  AND3_X1   g295(.A1(new_n466), .A2(new_n479), .A3(new_n481), .ZN(new_n482));
  AOI21_X1  g296(.A(new_n481), .B1(new_n466), .B2(new_n479), .ZN(new_n483));
  OAI21_X1  g297(.A(new_n303), .B1(new_n482), .B2(new_n483), .ZN(new_n484));
  NAND2_X1  g298(.A1(new_n484), .A2(KEYINPUT91), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n466), .A2(new_n479), .ZN(new_n486));
  OR2_X1    g300(.A1(new_n298), .A2(new_n480), .ZN(new_n487));
  NAND2_X1  g301(.A1(new_n486), .A2(new_n487), .ZN(new_n488));
  NAND3_X1  g302(.A1(new_n466), .A2(new_n479), .A3(new_n481), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  INV_X1    g304(.A(KEYINPUT91), .ZN(new_n491));
  NAND3_X1  g305(.A1(new_n490), .A2(new_n491), .A3(new_n303), .ZN(new_n492));
  INV_X1    g306(.A(G478), .ZN(new_n493));
  NOR2_X1   g307(.A1(new_n493), .A2(KEYINPUT15), .ZN(new_n494));
  NAND3_X1  g308(.A1(new_n485), .A2(new_n492), .A3(new_n494), .ZN(new_n495));
  INV_X1    g309(.A(KEYINPUT92), .ZN(new_n496));
  OR3_X1    g310(.A1(new_n484), .A2(new_n496), .A3(new_n494), .ZN(new_n497));
  OAI21_X1  g311(.A(new_n496), .B1(new_n484), .B2(new_n494), .ZN(new_n498));
  AND3_X1   g312(.A1(new_n495), .A2(new_n497), .A3(new_n498), .ZN(new_n499));
  INV_X1    g313(.A(G952), .ZN(new_n500));
  AND2_X1   g314(.A1(new_n500), .A2(KEYINPUT93), .ZN(new_n501));
  NOR2_X1   g315(.A1(new_n500), .A2(KEYINPUT93), .ZN(new_n502));
  OAI21_X1  g316(.A(new_n234), .B1(new_n501), .B2(new_n502), .ZN(new_n503));
  AOI21_X1  g317(.A(new_n503), .B1(G234), .B2(G237), .ZN(new_n504));
  INV_X1    g318(.A(new_n504), .ZN(new_n505));
  AOI211_X1 g319(.A(new_n234), .B(new_n303), .C1(G234), .C2(G237), .ZN(new_n506));
  INV_X1    g320(.A(new_n506), .ZN(new_n507));
  XNOR2_X1  g321(.A(KEYINPUT21), .B(G898), .ZN(new_n508));
  XNOR2_X1  g322(.A(new_n508), .B(KEYINPUT94), .ZN(new_n509));
  OAI21_X1  g323(.A(new_n505), .B1(new_n507), .B2(new_n509), .ZN(new_n510));
  NAND4_X1  g324(.A1(new_n423), .A2(new_n446), .A3(new_n499), .A4(new_n510), .ZN(new_n511));
  NOR3_X1   g325(.A1(new_n297), .A2(new_n363), .A3(new_n511), .ZN(new_n512));
  INV_X1    g326(.A(KEYINPUT77), .ZN(new_n513));
  INV_X1    g327(.A(G217), .ZN(new_n514));
  AOI21_X1  g328(.A(new_n514), .B1(new_n303), .B2(G234), .ZN(new_n515));
  INV_X1    g329(.A(KEYINPUT75), .ZN(new_n516));
  NOR2_X1   g330(.A1(new_n516), .A2(KEYINPUT25), .ZN(new_n517));
  INV_X1    g331(.A(new_n517), .ZN(new_n518));
  XNOR2_X1  g332(.A(KEYINPUT22), .B(G137), .ZN(new_n519));
  NAND3_X1  g333(.A1(new_n234), .A2(G221), .A3(G234), .ZN(new_n520));
  XNOR2_X1  g334(.A(new_n519), .B(new_n520), .ZN(new_n521));
  OAI21_X1  g335(.A(KEYINPUT73), .B1(new_n400), .B2(new_n242), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n223), .A2(G128), .ZN(new_n523));
  NAND3_X1  g337(.A1(new_n259), .A2(KEYINPUT23), .A3(G119), .ZN(new_n524));
  NOR2_X1   g338(.A1(new_n223), .A2(G128), .ZN(new_n525));
  OAI211_X1 g339(.A(new_n523), .B(new_n524), .C1(new_n525), .C2(KEYINPUT23), .ZN(new_n526));
  OR2_X1    g340(.A1(new_n526), .A2(G110), .ZN(new_n527));
  XNOR2_X1  g341(.A(KEYINPUT24), .B(G110), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n259), .A2(G119), .ZN(new_n529));
  INV_X1    g343(.A(KEYINPUT71), .ZN(new_n530));
  AND3_X1   g344(.A1(new_n523), .A2(new_n529), .A3(new_n530), .ZN(new_n531));
  AOI21_X1  g345(.A(new_n530), .B1(new_n523), .B2(new_n529), .ZN(new_n532));
  OAI21_X1  g346(.A(new_n528), .B1(new_n531), .B2(new_n532), .ZN(new_n533));
  AOI22_X1  g347(.A1(new_n527), .A2(new_n533), .B1(new_n252), .B2(new_n381), .ZN(new_n534));
  NAND2_X1  g348(.A1(new_n408), .A2(new_n428), .ZN(new_n535));
  NAND3_X1  g349(.A1(new_n522), .A2(new_n534), .A3(new_n535), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n536), .A2(KEYINPUT74), .ZN(new_n537));
  INV_X1    g351(.A(KEYINPUT74), .ZN(new_n538));
  NAND4_X1  g352(.A1(new_n522), .A2(new_n534), .A3(new_n538), .A4(new_n535), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n537), .A2(new_n539), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n526), .A2(G110), .ZN(new_n541));
  OR2_X1    g355(.A1(new_n531), .A2(new_n532), .ZN(new_n542));
  OAI21_X1  g356(.A(new_n541), .B1(new_n542), .B2(new_n528), .ZN(new_n543));
  AOI21_X1  g357(.A(new_n543), .B1(new_n409), .B2(new_n401), .ZN(new_n544));
  INV_X1    g358(.A(new_n544), .ZN(new_n545));
  AOI21_X1  g359(.A(new_n521), .B1(new_n540), .B2(new_n545), .ZN(new_n546));
  INV_X1    g360(.A(new_n521), .ZN(new_n547));
  AOI211_X1 g361(.A(new_n544), .B(new_n547), .C1(new_n537), .C2(new_n539), .ZN(new_n548));
  NOR2_X1   g362(.A1(new_n546), .A2(new_n548), .ZN(new_n549));
  AOI21_X1  g363(.A(new_n518), .B1(new_n549), .B2(new_n303), .ZN(new_n550));
  AOI21_X1  g364(.A(new_n538), .B1(new_n431), .B2(new_n534), .ZN(new_n551));
  INV_X1    g365(.A(new_n539), .ZN(new_n552));
  OAI21_X1  g366(.A(new_n545), .B1(new_n551), .B2(new_n552), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n553), .A2(new_n547), .ZN(new_n554));
  NAND3_X1  g368(.A1(new_n540), .A2(new_n545), .A3(new_n521), .ZN(new_n555));
  NAND4_X1  g369(.A1(new_n554), .A2(new_n555), .A3(new_n303), .A4(new_n518), .ZN(new_n556));
  INV_X1    g370(.A(new_n556), .ZN(new_n557));
  OAI21_X1  g371(.A(new_n515), .B1(new_n550), .B2(new_n557), .ZN(new_n558));
  INV_X1    g372(.A(new_n515), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n559), .A2(new_n281), .ZN(new_n560));
  XNOR2_X1  g374(.A(new_n560), .B(KEYINPUT76), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n549), .A2(new_n561), .ZN(new_n562));
  AOI21_X1  g376(.A(new_n513), .B1(new_n558), .B2(new_n562), .ZN(new_n563));
  NAND3_X1  g377(.A1(new_n554), .A2(new_n555), .A3(new_n303), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n564), .A2(new_n517), .ZN(new_n565));
  AOI21_X1  g379(.A(new_n559), .B1(new_n565), .B2(new_n556), .ZN(new_n566));
  INV_X1    g380(.A(new_n562), .ZN(new_n567));
  NOR3_X1   g381(.A1(new_n566), .A2(KEYINPUT77), .A3(new_n567), .ZN(new_n568));
  NOR2_X1   g382(.A1(new_n563), .A2(new_n568), .ZN(new_n569));
  NAND3_X1  g383(.A1(new_n368), .A2(new_n234), .A3(G210), .ZN(new_n570));
  XOR2_X1   g384(.A(new_n570), .B(KEYINPUT27), .Z(new_n571));
  XNOR2_X1  g385(.A(KEYINPUT26), .B(G101), .ZN(new_n572));
  XNOR2_X1  g386(.A(new_n571), .B(new_n572), .ZN(new_n573));
  INV_X1    g387(.A(new_n573), .ZN(new_n574));
  XOR2_X1   g388(.A(KEYINPUT67), .B(KEYINPUT28), .Z(new_n575));
  NAND3_X1  g389(.A1(new_n254), .A2(new_n338), .A3(new_n255), .ZN(new_n576));
  INV_X1    g390(.A(new_n214), .ZN(new_n577));
  NOR2_X1   g391(.A1(new_n316), .A2(G137), .ZN(new_n578));
  NOR2_X1   g392(.A1(new_n319), .A2(G134), .ZN(new_n579));
  OAI21_X1  g393(.A(G131), .B1(new_n578), .B2(new_n579), .ZN(new_n580));
  AND2_X1   g394(.A1(new_n329), .A2(new_n580), .ZN(new_n581));
  NAND2_X1  g395(.A1(new_n581), .A2(new_n314), .ZN(new_n582));
  AND3_X1   g396(.A1(new_n576), .A2(new_n577), .A3(new_n582), .ZN(new_n583));
  AOI21_X1  g397(.A(new_n577), .B1(new_n576), .B2(new_n582), .ZN(new_n584));
  OAI21_X1  g398(.A(new_n575), .B1(new_n583), .B2(new_n584), .ZN(new_n585));
  NAND3_X1  g399(.A1(new_n576), .A2(new_n577), .A3(new_n582), .ZN(new_n586));
  INV_X1    g400(.A(KEYINPUT28), .ZN(new_n587));
  NAND2_X1  g401(.A1(new_n586), .A2(new_n587), .ZN(new_n588));
  AOI21_X1  g402(.A(new_n574), .B1(new_n585), .B2(new_n588), .ZN(new_n589));
  INV_X1    g403(.A(new_n589), .ZN(new_n590));
  OAI21_X1  g404(.A(new_n582), .B1(new_n270), .B2(new_n330), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n591), .A2(KEYINPUT30), .ZN(new_n592));
  INV_X1    g406(.A(KEYINPUT30), .ZN(new_n593));
  NAND3_X1  g407(.A1(new_n576), .A2(new_n593), .A3(new_n582), .ZN(new_n594));
  NAND2_X1  g408(.A1(new_n592), .A2(new_n594), .ZN(new_n595));
  AOI21_X1  g409(.A(new_n583), .B1(new_n595), .B2(new_n214), .ZN(new_n596));
  AOI21_X1  g410(.A(KEYINPUT31), .B1(new_n596), .B2(new_n574), .ZN(new_n597));
  AND3_X1   g411(.A1(new_n576), .A2(new_n593), .A3(new_n582), .ZN(new_n598));
  AOI21_X1  g412(.A(new_n593), .B1(new_n576), .B2(new_n582), .ZN(new_n599));
  OAI21_X1  g413(.A(new_n214), .B1(new_n598), .B2(new_n599), .ZN(new_n600));
  NAND4_X1  g414(.A1(new_n600), .A2(KEYINPUT31), .A3(new_n574), .A4(new_n586), .ZN(new_n601));
  INV_X1    g415(.A(new_n601), .ZN(new_n602));
  OAI21_X1  g416(.A(new_n590), .B1(new_n597), .B2(new_n602), .ZN(new_n603));
  INV_X1    g417(.A(KEYINPUT32), .ZN(new_n604));
  NOR2_X1   g418(.A1(G472), .A2(G902), .ZN(new_n605));
  NAND3_X1  g419(.A1(new_n603), .A2(new_n604), .A3(new_n605), .ZN(new_n606));
  NAND3_X1  g420(.A1(new_n600), .A2(new_n574), .A3(new_n586), .ZN(new_n607));
  INV_X1    g421(.A(KEYINPUT31), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  AOI21_X1  g423(.A(new_n589), .B1(new_n609), .B2(new_n601), .ZN(new_n610));
  INV_X1    g424(.A(new_n605), .ZN(new_n611));
  OAI21_X1  g425(.A(KEYINPUT32), .B1(new_n610), .B2(new_n611), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n606), .A2(new_n612), .ZN(new_n613));
  INV_X1    g427(.A(new_n303), .ZN(new_n614));
  INV_X1    g428(.A(KEYINPUT69), .ZN(new_n615));
  OAI211_X1 g429(.A(new_n615), .B(KEYINPUT28), .C1(new_n583), .C2(new_n584), .ZN(new_n616));
  NAND2_X1  g430(.A1(new_n616), .A2(new_n588), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n591), .A2(new_n214), .ZN(new_n618));
  NAND2_X1  g432(.A1(new_n618), .A2(new_n586), .ZN(new_n619));
  AOI21_X1  g433(.A(new_n615), .B1(new_n619), .B2(KEYINPUT28), .ZN(new_n620));
  NOR2_X1   g434(.A1(new_n617), .A2(new_n620), .ZN(new_n621));
  INV_X1    g435(.A(KEYINPUT29), .ZN(new_n622));
  NOR2_X1   g436(.A1(new_n573), .A2(new_n622), .ZN(new_n623));
  AOI21_X1  g437(.A(new_n614), .B1(new_n621), .B2(new_n623), .ZN(new_n624));
  AOI21_X1  g438(.A(new_n577), .B1(new_n592), .B2(new_n594), .ZN(new_n625));
  OAI21_X1  g439(.A(new_n573), .B1(new_n625), .B2(new_n583), .ZN(new_n626));
  NAND3_X1  g440(.A1(new_n585), .A2(new_n574), .A3(new_n588), .ZN(new_n627));
  NAND3_X1  g441(.A1(new_n626), .A2(new_n622), .A3(new_n627), .ZN(new_n628));
  INV_X1    g442(.A(KEYINPUT68), .ZN(new_n629));
  NAND2_X1  g443(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  NAND4_X1  g444(.A1(new_n626), .A2(KEYINPUT68), .A3(new_n627), .A4(new_n622), .ZN(new_n631));
  NAND3_X1  g445(.A1(new_n624), .A2(new_n630), .A3(new_n631), .ZN(new_n632));
  NAND2_X1  g446(.A1(new_n632), .A2(G472), .ZN(new_n633));
  NAND2_X1  g447(.A1(new_n613), .A2(new_n633), .ZN(new_n634));
  NAND3_X1  g448(.A1(new_n512), .A2(new_n569), .A3(new_n634), .ZN(new_n635));
  XNOR2_X1  g449(.A(new_n635), .B(G101), .ZN(G3));
  OAI21_X1  g450(.A(G472), .B1(new_n610), .B2(new_n614), .ZN(new_n637));
  NAND2_X1  g451(.A1(new_n603), .A2(new_n605), .ZN(new_n638));
  NAND2_X1  g452(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  NOR2_X1   g453(.A1(new_n639), .A2(new_n363), .ZN(new_n640));
  OAI211_X1 g454(.A(new_n187), .B(new_n510), .C1(new_n294), .C2(new_n296), .ZN(new_n641));
  NAND2_X1  g455(.A1(new_n423), .A2(new_n446), .ZN(new_n642));
  NAND3_X1  g456(.A1(new_n485), .A2(new_n492), .A3(new_n493), .ZN(new_n643));
  INV_X1    g457(.A(KEYINPUT95), .ZN(new_n644));
  OR2_X1    g458(.A1(new_n644), .A2(KEYINPUT33), .ZN(new_n645));
  NAND2_X1  g459(.A1(new_n644), .A2(KEYINPUT33), .ZN(new_n646));
  NAND2_X1  g460(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  MUX2_X1   g461(.A(new_n647), .B(new_n646), .S(new_n490), .Z(new_n648));
  NAND2_X1  g462(.A1(new_n303), .A2(G478), .ZN(new_n649));
  OAI21_X1  g463(.A(new_n643), .B1(new_n648), .B2(new_n649), .ZN(new_n650));
  NAND2_X1  g464(.A1(new_n642), .A2(new_n650), .ZN(new_n651));
  NOR2_X1   g465(.A1(new_n641), .A2(new_n651), .ZN(new_n652));
  NAND3_X1  g466(.A1(new_n569), .A2(new_n640), .A3(new_n652), .ZN(new_n653));
  XOR2_X1   g467(.A(KEYINPUT34), .B(G104), .Z(new_n654));
  XNOR2_X1  g468(.A(new_n653), .B(new_n654), .ZN(G6));
  INV_X1    g469(.A(new_n641), .ZN(new_n656));
  AOI21_X1  g470(.A(new_n499), .B1(new_n422), .B2(new_n420), .ZN(new_n657));
  NAND3_X1  g471(.A1(new_n442), .A2(KEYINPUT96), .A3(KEYINPUT20), .ZN(new_n658));
  INV_X1    g472(.A(KEYINPUT96), .ZN(new_n659));
  NAND3_X1  g473(.A1(new_n443), .A2(new_n659), .A3(new_n445), .ZN(new_n660));
  AND3_X1   g474(.A1(new_n657), .A2(new_n658), .A3(new_n660), .ZN(new_n661));
  NAND4_X1  g475(.A1(new_n569), .A2(new_n640), .A3(new_n656), .A4(new_n661), .ZN(new_n662));
  XOR2_X1   g476(.A(KEYINPUT35), .B(G107), .Z(new_n663));
  XNOR2_X1  g477(.A(new_n662), .B(new_n663), .ZN(new_n664));
  XNOR2_X1  g478(.A(KEYINPUT97), .B(KEYINPUT98), .ZN(new_n665));
  XNOR2_X1  g479(.A(new_n664), .B(new_n665), .ZN(G9));
  NOR2_X1   g480(.A1(new_n547), .A2(KEYINPUT36), .ZN(new_n667));
  XNOR2_X1  g481(.A(new_n553), .B(new_n667), .ZN(new_n668));
  AND2_X1   g482(.A1(new_n668), .A2(new_n561), .ZN(new_n669));
  NOR2_X1   g483(.A1(new_n566), .A2(new_n669), .ZN(new_n670));
  NOR2_X1   g484(.A1(new_n639), .A2(new_n670), .ZN(new_n671));
  NAND2_X1  g485(.A1(new_n512), .A2(new_n671), .ZN(new_n672));
  XOR2_X1   g486(.A(KEYINPUT37), .B(G110), .Z(new_n673));
  XNOR2_X1  g487(.A(new_n672), .B(new_n673), .ZN(G12));
  NOR2_X1   g488(.A1(new_n297), .A2(new_n363), .ZN(new_n675));
  INV_X1    g489(.A(G900), .ZN(new_n676));
  AOI21_X1  g490(.A(new_n504), .B1(new_n506), .B2(new_n676), .ZN(new_n677));
  INV_X1    g491(.A(new_n677), .ZN(new_n678));
  AND4_X1   g492(.A1(new_n658), .A2(new_n657), .A3(new_n660), .A4(new_n678), .ZN(new_n679));
  NAND2_X1  g493(.A1(new_n668), .A2(new_n561), .ZN(new_n680));
  NAND2_X1  g494(.A1(new_n558), .A2(new_n680), .ZN(new_n681));
  NAND4_X1  g495(.A1(new_n675), .A2(new_n634), .A3(new_n679), .A4(new_n681), .ZN(new_n682));
  XNOR2_X1  g496(.A(new_n682), .B(G128), .ZN(G30));
  NAND2_X1  g497(.A1(new_n280), .A2(new_n293), .ZN(new_n684));
  NAND2_X1  g498(.A1(new_n684), .A2(new_n295), .ZN(new_n685));
  NAND3_X1  g499(.A1(new_n280), .A2(new_n293), .A3(new_n188), .ZN(new_n686));
  NAND2_X1  g500(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  XNOR2_X1  g501(.A(new_n687), .B(KEYINPUT38), .ZN(new_n688));
  INV_X1    g502(.A(new_n499), .ZN(new_n689));
  NAND2_X1  g503(.A1(new_n642), .A2(new_n689), .ZN(new_n690));
  INV_X1    g504(.A(new_n690), .ZN(new_n691));
  NAND4_X1  g505(.A1(new_n688), .A2(new_n187), .A3(new_n670), .A4(new_n691), .ZN(new_n692));
  NOR2_X1   g506(.A1(new_n619), .A2(new_n574), .ZN(new_n693));
  INV_X1    g507(.A(new_n693), .ZN(new_n694));
  INV_X1    g508(.A(KEYINPUT99), .ZN(new_n695));
  OAI211_X1 g509(.A(new_n694), .B(new_n695), .C1(new_n596), .C2(new_n573), .ZN(new_n696));
  AOI21_X1  g510(.A(new_n573), .B1(new_n600), .B2(new_n586), .ZN(new_n697));
  OAI21_X1  g511(.A(KEYINPUT99), .B1(new_n697), .B2(new_n693), .ZN(new_n698));
  NAND3_X1  g512(.A1(new_n696), .A2(new_n281), .A3(new_n698), .ZN(new_n699));
  AOI22_X1  g513(.A1(new_n606), .A2(new_n612), .B1(G472), .B2(new_n699), .ZN(new_n700));
  AND2_X1   g514(.A1(new_n359), .A2(new_n361), .ZN(new_n701));
  AOI21_X1  g515(.A(new_n300), .B1(new_n701), .B2(new_n351), .ZN(new_n702));
  XOR2_X1   g516(.A(new_n677), .B(KEYINPUT39), .Z(new_n703));
  NAND2_X1  g517(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  AOI21_X1  g518(.A(new_n700), .B1(KEYINPUT40), .B2(new_n704), .ZN(new_n705));
  OAI21_X1  g519(.A(new_n705), .B1(KEYINPUT40), .B2(new_n704), .ZN(new_n706));
  NOR2_X1   g520(.A1(new_n692), .A2(new_n706), .ZN(new_n707));
  XNOR2_X1  g521(.A(new_n707), .B(KEYINPUT100), .ZN(new_n708));
  XNOR2_X1  g522(.A(new_n708), .B(G143), .ZN(G45));
  AND3_X1   g523(.A1(new_n642), .A2(new_n650), .A3(new_n678), .ZN(new_n710));
  NAND4_X1  g524(.A1(new_n675), .A2(new_n634), .A3(new_n681), .A4(new_n710), .ZN(new_n711));
  XNOR2_X1  g525(.A(new_n711), .B(G146), .ZN(G48));
  OAI21_X1  g526(.A(new_n303), .B1(new_n342), .B2(new_n350), .ZN(new_n713));
  NAND2_X1  g527(.A1(new_n713), .A2(G469), .ZN(new_n714));
  NAND3_X1  g528(.A1(new_n714), .A2(new_n301), .A3(new_n351), .ZN(new_n715));
  INV_X1    g529(.A(new_n715), .ZN(new_n716));
  NAND4_X1  g530(.A1(new_n569), .A2(new_n652), .A3(new_n634), .A4(new_n716), .ZN(new_n717));
  XOR2_X1   g531(.A(KEYINPUT41), .B(G113), .Z(new_n718));
  XNOR2_X1  g532(.A(new_n718), .B(KEYINPUT101), .ZN(new_n719));
  XNOR2_X1  g533(.A(new_n717), .B(new_n719), .ZN(G15));
  AOI21_X1  g534(.A(new_n715), .B1(new_n613), .B2(new_n633), .ZN(new_n721));
  NAND4_X1  g535(.A1(new_n569), .A2(new_n721), .A3(new_n656), .A4(new_n661), .ZN(new_n722));
  XNOR2_X1  g536(.A(new_n722), .B(G116), .ZN(G18));
  NOR3_X1   g537(.A1(new_n297), .A2(new_n715), .A3(new_n511), .ZN(new_n724));
  AOI21_X1  g538(.A(new_n670), .B1(new_n613), .B2(new_n633), .ZN(new_n725));
  NAND2_X1  g539(.A1(new_n724), .A2(new_n725), .ZN(new_n726));
  XNOR2_X1  g540(.A(new_n726), .B(G119), .ZN(G21));
  NOR3_X1   g541(.A1(new_n641), .A2(new_n690), .A3(new_n715), .ZN(new_n728));
  NOR2_X1   g542(.A1(new_n566), .A2(new_n567), .ZN(new_n729));
  NAND2_X1  g543(.A1(new_n609), .A2(new_n601), .ZN(new_n730));
  OAI21_X1  g544(.A(new_n573), .B1(new_n617), .B2(new_n620), .ZN(new_n731));
  AOI21_X1  g545(.A(new_n611), .B1(new_n730), .B2(new_n731), .ZN(new_n732));
  INV_X1    g546(.A(KEYINPUT102), .ZN(new_n733));
  NAND2_X1  g547(.A1(new_n637), .A2(new_n733), .ZN(new_n734));
  OAI211_X1 g548(.A(KEYINPUT102), .B(G472), .C1(new_n610), .C2(new_n614), .ZN(new_n735));
  AOI21_X1  g549(.A(new_n732), .B1(new_n734), .B2(new_n735), .ZN(new_n736));
  NAND3_X1  g550(.A1(new_n728), .A2(new_n729), .A3(new_n736), .ZN(new_n737));
  XNOR2_X1  g551(.A(new_n737), .B(G122), .ZN(G24));
  NOR2_X1   g552(.A1(new_n297), .A2(new_n715), .ZN(new_n739));
  NAND4_X1  g553(.A1(new_n736), .A2(new_n739), .A3(new_n681), .A4(new_n710), .ZN(new_n740));
  XNOR2_X1  g554(.A(new_n740), .B(G125), .ZN(G27));
  NAND3_X1  g555(.A1(new_n685), .A2(new_n187), .A3(new_n686), .ZN(new_n742));
  NOR2_X1   g556(.A1(new_n742), .A2(new_n363), .ZN(new_n743));
  NAND4_X1  g557(.A1(new_n569), .A2(new_n634), .A3(new_n743), .A4(new_n710), .ZN(new_n744));
  XOR2_X1   g558(.A(KEYINPUT103), .B(KEYINPUT42), .Z(new_n745));
  AND3_X1   g559(.A1(new_n743), .A2(KEYINPUT42), .A3(new_n710), .ZN(new_n746));
  AND2_X1   g560(.A1(new_n634), .A2(new_n729), .ZN(new_n747));
  AOI22_X1  g561(.A1(new_n744), .A2(new_n745), .B1(new_n746), .B2(new_n747), .ZN(new_n748));
  XNOR2_X1  g562(.A(new_n748), .B(new_n328), .ZN(G33));
  NAND4_X1  g563(.A1(new_n569), .A2(new_n634), .A3(new_n743), .A4(new_n679), .ZN(new_n750));
  XNOR2_X1  g564(.A(new_n750), .B(G134), .ZN(G36));
  NAND3_X1  g565(.A1(new_n423), .A2(new_n446), .A3(new_n650), .ZN(new_n752));
  XOR2_X1   g566(.A(new_n752), .B(KEYINPUT43), .Z(new_n753));
  AND2_X1   g567(.A1(new_n639), .A2(new_n681), .ZN(new_n754));
  NAND2_X1  g568(.A1(new_n753), .A2(new_n754), .ZN(new_n755));
  INV_X1    g569(.A(new_n755), .ZN(new_n756));
  NOR2_X1   g570(.A1(new_n756), .A2(KEYINPUT44), .ZN(new_n757));
  INV_X1    g571(.A(new_n187), .ZN(new_n758));
  NOR3_X1   g572(.A1(new_n294), .A2(new_n296), .A3(new_n758), .ZN(new_n759));
  INV_X1    g573(.A(KEYINPUT44), .ZN(new_n760));
  OAI21_X1  g574(.A(new_n759), .B1(new_n755), .B2(new_n760), .ZN(new_n761));
  OAI21_X1  g575(.A(new_n354), .B1(new_n356), .B2(new_n358), .ZN(new_n762));
  INV_X1    g576(.A(KEYINPUT45), .ZN(new_n763));
  OR2_X1    g577(.A1(new_n762), .A2(new_n763), .ZN(new_n764));
  AOI21_X1  g578(.A(new_n302), .B1(new_n762), .B2(new_n763), .ZN(new_n765));
  NAND2_X1  g579(.A1(new_n764), .A2(new_n765), .ZN(new_n766));
  NAND2_X1  g580(.A1(new_n766), .A2(new_n361), .ZN(new_n767));
  INV_X1    g581(.A(new_n767), .ZN(new_n768));
  AND2_X1   g582(.A1(new_n768), .A2(KEYINPUT46), .ZN(new_n769));
  OAI21_X1  g583(.A(new_n351), .B1(new_n768), .B2(KEYINPUT46), .ZN(new_n770));
  OAI211_X1 g584(.A(new_n301), .B(new_n703), .C1(new_n769), .C2(new_n770), .ZN(new_n771));
  NOR3_X1   g585(.A1(new_n757), .A2(new_n761), .A3(new_n771), .ZN(new_n772));
  XNOR2_X1  g586(.A(new_n772), .B(new_n319), .ZN(G39));
  OAI21_X1  g587(.A(new_n301), .B1(new_n769), .B2(new_n770), .ZN(new_n774));
  INV_X1    g588(.A(KEYINPUT104), .ZN(new_n775));
  OAI21_X1  g589(.A(new_n774), .B1(new_n775), .B2(KEYINPUT47), .ZN(new_n776));
  INV_X1    g590(.A(new_n569), .ZN(new_n777));
  XOR2_X1   g591(.A(KEYINPUT104), .B(KEYINPUT47), .Z(new_n778));
  OAI211_X1 g592(.A(new_n301), .B(new_n778), .C1(new_n769), .C2(new_n770), .ZN(new_n779));
  NOR4_X1   g593(.A1(new_n634), .A2(new_n651), .A3(new_n677), .A4(new_n742), .ZN(new_n780));
  NAND4_X1  g594(.A1(new_n776), .A2(new_n777), .A3(new_n779), .A4(new_n780), .ZN(new_n781));
  XNOR2_X1  g595(.A(new_n781), .B(G140), .ZN(G42));
  NAND3_X1  g596(.A1(new_n729), .A2(new_n187), .A3(new_n301), .ZN(new_n783));
  OR2_X1    g597(.A1(new_n783), .A2(new_n752), .ZN(new_n784));
  AND2_X1   g598(.A1(new_n714), .A2(new_n351), .ZN(new_n785));
  INV_X1    g599(.A(new_n785), .ZN(new_n786));
  AOI22_X1  g600(.A1(new_n784), .A2(KEYINPUT105), .B1(KEYINPUT49), .B2(new_n786), .ZN(new_n787));
  OAI21_X1  g601(.A(new_n787), .B1(KEYINPUT105), .B2(new_n784), .ZN(new_n788));
  XNOR2_X1  g602(.A(new_n788), .B(KEYINPUT106), .ZN(new_n789));
  NAND2_X1  g603(.A1(new_n699), .A2(G472), .ZN(new_n790));
  AOI21_X1  g604(.A(new_n604), .B1(new_n603), .B2(new_n605), .ZN(new_n791));
  NOR3_X1   g605(.A1(new_n610), .A2(KEYINPUT32), .A3(new_n611), .ZN(new_n792));
  OAI21_X1  g606(.A(new_n790), .B1(new_n791), .B2(new_n792), .ZN(new_n793));
  NOR2_X1   g607(.A1(new_n786), .A2(KEYINPUT49), .ZN(new_n794));
  OR4_X1    g608(.A1(new_n688), .A2(new_n789), .A3(new_n793), .A4(new_n794), .ZN(new_n795));
  INV_X1    g609(.A(KEYINPUT53), .ZN(new_n796));
  NAND4_X1  g610(.A1(new_n495), .A2(new_n497), .A3(new_n498), .A4(new_n678), .ZN(new_n797));
  AOI21_X1  g611(.A(new_n797), .B1(new_n420), .B2(new_n422), .ZN(new_n798));
  AND3_X1   g612(.A1(new_n798), .A2(new_n658), .A3(new_n660), .ZN(new_n799));
  NAND3_X1  g613(.A1(new_n799), .A2(new_n759), .A3(KEYINPUT108), .ZN(new_n800));
  INV_X1    g614(.A(KEYINPUT108), .ZN(new_n801));
  NAND3_X1  g615(.A1(new_n798), .A2(new_n658), .A3(new_n660), .ZN(new_n802));
  OAI21_X1  g616(.A(new_n801), .B1(new_n742), .B2(new_n802), .ZN(new_n803));
  NAND4_X1  g617(.A1(new_n725), .A2(new_n800), .A3(new_n803), .A4(new_n702), .ZN(new_n804));
  NAND4_X1  g618(.A1(new_n736), .A2(new_n743), .A3(new_n681), .A4(new_n710), .ZN(new_n805));
  NAND3_X1  g619(.A1(new_n804), .A2(new_n750), .A3(new_n805), .ZN(new_n806));
  NAND2_X1  g620(.A1(new_n806), .A2(KEYINPUT109), .ZN(new_n807));
  INV_X1    g621(.A(KEYINPUT109), .ZN(new_n808));
  NAND4_X1  g622(.A1(new_n804), .A2(new_n750), .A3(new_n805), .A4(new_n808), .ZN(new_n809));
  NAND2_X1  g623(.A1(new_n807), .A2(new_n809), .ZN(new_n810));
  AOI22_X1  g624(.A1(new_n725), .A2(new_n724), .B1(new_n512), .B2(new_n671), .ZN(new_n811));
  AOI21_X1  g625(.A(new_n758), .B1(new_n685), .B2(new_n686), .ZN(new_n812));
  NAND3_X1  g626(.A1(new_n423), .A2(new_n689), .A3(new_n446), .ZN(new_n813));
  INV_X1    g627(.A(new_n813), .ZN(new_n814));
  INV_X1    g628(.A(KEYINPUT107), .ZN(new_n815));
  NAND4_X1  g629(.A1(new_n812), .A2(new_n814), .A3(new_n815), .A4(new_n510), .ZN(new_n816));
  OAI21_X1  g630(.A(KEYINPUT107), .B1(new_n641), .B2(new_n813), .ZN(new_n817));
  NAND4_X1  g631(.A1(new_n816), .A2(new_n569), .A3(new_n817), .A4(new_n640), .ZN(new_n818));
  NAND4_X1  g632(.A1(new_n811), .A2(new_n635), .A3(new_n818), .A4(new_n653), .ZN(new_n819));
  NAND3_X1  g633(.A1(new_n722), .A2(new_n717), .A3(new_n737), .ZN(new_n820));
  NOR2_X1   g634(.A1(new_n819), .A2(new_n820), .ZN(new_n821));
  INV_X1    g635(.A(new_n748), .ZN(new_n822));
  NAND3_X1  g636(.A1(new_n810), .A2(new_n821), .A3(new_n822), .ZN(new_n823));
  INV_X1    g637(.A(KEYINPUT110), .ZN(new_n824));
  OAI211_X1 g638(.A(new_n301), .B(new_n678), .C1(new_n352), .C2(new_n362), .ZN(new_n825));
  NOR3_X1   g639(.A1(new_n700), .A2(new_n681), .A3(new_n825), .ZN(new_n826));
  NOR2_X1   g640(.A1(new_n297), .A2(new_n690), .ZN(new_n827));
  AOI21_X1  g641(.A(new_n824), .B1(new_n826), .B2(new_n827), .ZN(new_n828));
  NOR2_X1   g642(.A1(new_n825), .A2(new_n681), .ZN(new_n829));
  AND4_X1   g643(.A1(new_n824), .A2(new_n829), .A3(new_n827), .A4(new_n793), .ZN(new_n830));
  NOR2_X1   g644(.A1(new_n828), .A2(new_n830), .ZN(new_n831));
  NAND3_X1  g645(.A1(new_n740), .A2(new_n682), .A3(new_n711), .ZN(new_n832));
  OAI21_X1  g646(.A(KEYINPUT52), .B1(new_n831), .B2(new_n832), .ZN(new_n833));
  AND3_X1   g647(.A1(new_n740), .A2(new_n682), .A3(new_n711), .ZN(new_n834));
  AOI211_X1 g648(.A(new_n300), .B(new_n677), .C1(new_n701), .C2(new_n351), .ZN(new_n835));
  NAND3_X1  g649(.A1(new_n793), .A2(new_n670), .A3(new_n835), .ZN(new_n836));
  NAND2_X1  g650(.A1(new_n691), .A2(new_n812), .ZN(new_n837));
  OAI21_X1  g651(.A(KEYINPUT110), .B1(new_n836), .B2(new_n837), .ZN(new_n838));
  NAND4_X1  g652(.A1(new_n829), .A2(new_n827), .A3(new_n824), .A4(new_n793), .ZN(new_n839));
  NAND2_X1  g653(.A1(new_n838), .A2(new_n839), .ZN(new_n840));
  INV_X1    g654(.A(KEYINPUT52), .ZN(new_n841));
  NAND3_X1  g655(.A1(new_n834), .A2(new_n840), .A3(new_n841), .ZN(new_n842));
  NAND2_X1  g656(.A1(new_n833), .A2(new_n842), .ZN(new_n843));
  OAI21_X1  g657(.A(new_n796), .B1(new_n823), .B2(new_n843), .ZN(new_n844));
  AND3_X1   g658(.A1(new_n834), .A2(new_n840), .A3(new_n841), .ZN(new_n845));
  AOI21_X1  g659(.A(new_n841), .B1(new_n834), .B2(new_n840), .ZN(new_n846));
  NOR2_X1   g660(.A1(new_n845), .A2(new_n846), .ZN(new_n847));
  NOR3_X1   g661(.A1(new_n819), .A2(new_n748), .A3(new_n820), .ZN(new_n848));
  NAND4_X1  g662(.A1(new_n847), .A2(KEYINPUT53), .A3(new_n810), .A4(new_n848), .ZN(new_n849));
  INV_X1    g663(.A(KEYINPUT54), .ZN(new_n850));
  NAND3_X1  g664(.A1(new_n844), .A2(new_n849), .A3(new_n850), .ZN(new_n851));
  INV_X1    g665(.A(KEYINPUT112), .ZN(new_n852));
  NAND2_X1  g666(.A1(new_n851), .A2(new_n852), .ZN(new_n853));
  NAND4_X1  g667(.A1(new_n844), .A2(new_n849), .A3(KEYINPUT112), .A4(new_n850), .ZN(new_n854));
  NAND2_X1  g668(.A1(new_n853), .A2(new_n854), .ZN(new_n855));
  NAND2_X1  g669(.A1(new_n844), .A2(new_n849), .ZN(new_n856));
  NAND2_X1  g670(.A1(new_n856), .A2(KEYINPUT54), .ZN(new_n857));
  INV_X1    g671(.A(KEYINPUT111), .ZN(new_n858));
  NAND2_X1  g672(.A1(new_n857), .A2(new_n858), .ZN(new_n859));
  AND4_X1   g673(.A1(new_n504), .A2(new_n753), .A3(new_n716), .A4(new_n759), .ZN(new_n860));
  NAND2_X1  g674(.A1(new_n860), .A2(new_n747), .ZN(new_n861));
  XNOR2_X1  g675(.A(new_n861), .B(KEYINPUT48), .ZN(new_n862));
  NAND3_X1  g676(.A1(new_n700), .A2(new_n716), .A3(new_n759), .ZN(new_n863));
  NOR3_X1   g677(.A1(new_n777), .A2(new_n505), .A3(new_n863), .ZN(new_n864));
  INV_X1    g678(.A(new_n651), .ZN(new_n865));
  AOI21_X1  g679(.A(new_n503), .B1(new_n864), .B2(new_n865), .ZN(new_n866));
  AND2_X1   g680(.A1(new_n753), .A2(new_n504), .ZN(new_n867));
  NAND2_X1  g681(.A1(new_n736), .A2(new_n729), .ZN(new_n868));
  INV_X1    g682(.A(new_n868), .ZN(new_n869));
  NAND3_X1  g683(.A1(new_n867), .A2(new_n739), .A3(new_n869), .ZN(new_n870));
  AOI21_X1  g684(.A(KEYINPUT114), .B1(new_n866), .B2(new_n870), .ZN(new_n871));
  AND3_X1   g685(.A1(new_n866), .A2(KEYINPUT114), .A3(new_n870), .ZN(new_n872));
  OAI21_X1  g686(.A(new_n862), .B1(new_n871), .B2(new_n872), .ZN(new_n873));
  INV_X1    g687(.A(KEYINPUT115), .ZN(new_n874));
  NAND2_X1  g688(.A1(new_n873), .A2(new_n874), .ZN(new_n875));
  OAI211_X1 g689(.A(new_n862), .B(KEYINPUT115), .C1(new_n871), .C2(new_n872), .ZN(new_n876));
  AND2_X1   g690(.A1(new_n786), .A2(KEYINPUT113), .ZN(new_n877));
  NOR2_X1   g691(.A1(new_n786), .A2(KEYINPUT113), .ZN(new_n878));
  NOR3_X1   g692(.A1(new_n877), .A2(new_n878), .A3(new_n301), .ZN(new_n879));
  AOI21_X1  g693(.A(new_n879), .B1(new_n776), .B2(new_n779), .ZN(new_n880));
  NAND3_X1  g694(.A1(new_n867), .A2(new_n869), .A3(new_n759), .ZN(new_n881));
  OR2_X1    g695(.A1(new_n880), .A2(new_n881), .ZN(new_n882));
  NOR3_X1   g696(.A1(new_n688), .A2(new_n187), .A3(new_n715), .ZN(new_n883));
  NAND3_X1  g697(.A1(new_n883), .A2(new_n867), .A3(new_n869), .ZN(new_n884));
  XNOR2_X1  g698(.A(new_n884), .B(KEYINPUT50), .ZN(new_n885));
  INV_X1    g699(.A(new_n885), .ZN(new_n886));
  INV_X1    g700(.A(KEYINPUT51), .ZN(new_n887));
  NAND2_X1  g701(.A1(new_n736), .A2(new_n681), .ZN(new_n888));
  INV_X1    g702(.A(new_n888), .ZN(new_n889));
  NOR2_X1   g703(.A1(new_n642), .A2(new_n650), .ZN(new_n890));
  AOI22_X1  g704(.A1(new_n860), .A2(new_n889), .B1(new_n864), .B2(new_n890), .ZN(new_n891));
  NAND4_X1  g705(.A1(new_n882), .A2(new_n886), .A3(new_n887), .A4(new_n891), .ZN(new_n892));
  OAI21_X1  g706(.A(new_n891), .B1(new_n880), .B2(new_n881), .ZN(new_n893));
  OAI21_X1  g707(.A(KEYINPUT51), .B1(new_n893), .B2(new_n885), .ZN(new_n894));
  AOI22_X1  g708(.A1(new_n875), .A2(new_n876), .B1(new_n892), .B2(new_n894), .ZN(new_n895));
  AOI21_X1  g709(.A(new_n850), .B1(new_n844), .B2(new_n849), .ZN(new_n896));
  NAND2_X1  g710(.A1(new_n896), .A2(KEYINPUT111), .ZN(new_n897));
  AND4_X1   g711(.A1(new_n855), .A2(new_n859), .A3(new_n895), .A4(new_n897), .ZN(new_n898));
  NOR2_X1   g712(.A1(G952), .A2(G953), .ZN(new_n899));
  OAI21_X1  g713(.A(new_n795), .B1(new_n898), .B2(new_n899), .ZN(G75));
  NOR2_X1   g714(.A1(new_n234), .A2(G952), .ZN(new_n901));
  XNOR2_X1  g715(.A(new_n901), .B(KEYINPUT118), .ZN(new_n902));
  NAND3_X1  g716(.A1(new_n856), .A2(new_n614), .A3(new_n295), .ZN(new_n903));
  INV_X1    g717(.A(KEYINPUT56), .ZN(new_n904));
  NAND2_X1  g718(.A1(new_n903), .A2(new_n904), .ZN(new_n905));
  NAND2_X1  g719(.A1(new_n232), .A2(new_n275), .ZN(new_n906));
  XNOR2_X1  g720(.A(new_n906), .B(new_n273), .ZN(new_n907));
  XNOR2_X1  g721(.A(KEYINPUT116), .B(KEYINPUT55), .ZN(new_n908));
  XOR2_X1   g722(.A(new_n907), .B(new_n908), .Z(new_n909));
  OAI21_X1  g723(.A(new_n902), .B1(new_n905), .B2(new_n909), .ZN(new_n910));
  NAND2_X1  g724(.A1(new_n905), .A2(new_n909), .ZN(new_n911));
  INV_X1    g725(.A(KEYINPUT117), .ZN(new_n912));
  NAND2_X1  g726(.A1(new_n911), .A2(new_n912), .ZN(new_n913));
  NAND3_X1  g727(.A1(new_n905), .A2(KEYINPUT117), .A3(new_n909), .ZN(new_n914));
  AOI21_X1  g728(.A(new_n910), .B1(new_n913), .B2(new_n914), .ZN(G51));
  XNOR2_X1  g729(.A(KEYINPUT119), .B(KEYINPUT57), .ZN(new_n916));
  XNOR2_X1  g730(.A(new_n916), .B(new_n360), .ZN(new_n917));
  INV_X1    g731(.A(new_n851), .ZN(new_n918));
  OAI21_X1  g732(.A(new_n917), .B1(new_n918), .B2(new_n896), .ZN(new_n919));
  OAI21_X1  g733(.A(new_n919), .B1(new_n350), .B2(new_n342), .ZN(new_n920));
  NAND4_X1  g734(.A1(new_n856), .A2(new_n614), .A3(new_n764), .A4(new_n765), .ZN(new_n921));
  AOI21_X1  g735(.A(new_n901), .B1(new_n920), .B2(new_n921), .ZN(G54));
  INV_X1    g736(.A(KEYINPUT120), .ZN(new_n923));
  NAND4_X1  g737(.A1(new_n856), .A2(KEYINPUT58), .A3(G475), .A4(new_n614), .ZN(new_n924));
  NOR2_X1   g738(.A1(new_n441), .A2(new_n412), .ZN(new_n925));
  NAND2_X1  g739(.A1(new_n924), .A2(new_n925), .ZN(new_n926));
  INV_X1    g740(.A(new_n901), .ZN(new_n927));
  NAND2_X1  g741(.A1(new_n926), .A2(new_n927), .ZN(new_n928));
  NOR2_X1   g742(.A1(new_n924), .A2(new_n925), .ZN(new_n929));
  OAI21_X1  g743(.A(new_n923), .B1(new_n928), .B2(new_n929), .ZN(new_n930));
  AOI21_X1  g744(.A(new_n901), .B1(new_n924), .B2(new_n925), .ZN(new_n931));
  OAI211_X1 g745(.A(new_n931), .B(KEYINPUT120), .C1(new_n925), .C2(new_n924), .ZN(new_n932));
  NAND2_X1  g746(.A1(new_n930), .A2(new_n932), .ZN(G60));
  NAND2_X1  g747(.A1(G478), .A2(G902), .ZN(new_n934));
  XOR2_X1   g748(.A(new_n934), .B(KEYINPUT59), .Z(new_n935));
  NOR2_X1   g749(.A1(new_n648), .A2(new_n935), .ZN(new_n936));
  OAI21_X1  g750(.A(new_n936), .B1(new_n918), .B2(new_n896), .ZN(new_n937));
  NAND2_X1  g751(.A1(new_n937), .A2(new_n902), .ZN(new_n938));
  NAND3_X1  g752(.A1(new_n855), .A2(new_n859), .A3(new_n897), .ZN(new_n939));
  INV_X1    g753(.A(new_n935), .ZN(new_n940));
  NAND2_X1  g754(.A1(new_n939), .A2(new_n940), .ZN(new_n941));
  AOI21_X1  g755(.A(new_n938), .B1(new_n941), .B2(new_n648), .ZN(G63));
  NAND2_X1  g756(.A1(G217), .A2(G902), .ZN(new_n943));
  XNOR2_X1  g757(.A(new_n943), .B(KEYINPUT60), .ZN(new_n944));
  AOI21_X1  g758(.A(new_n944), .B1(new_n844), .B2(new_n849), .ZN(new_n945));
  XNOR2_X1  g759(.A(new_n668), .B(KEYINPUT121), .ZN(new_n946));
  AND2_X1   g760(.A1(new_n945), .A2(new_n946), .ZN(new_n947));
  INV_X1    g761(.A(new_n902), .ZN(new_n948));
  INV_X1    g762(.A(KEYINPUT122), .ZN(new_n949));
  INV_X1    g763(.A(KEYINPUT61), .ZN(new_n950));
  AOI21_X1  g764(.A(new_n948), .B1(new_n949), .B2(new_n950), .ZN(new_n951));
  OAI21_X1  g765(.A(new_n951), .B1(new_n945), .B2(new_n549), .ZN(new_n952));
  NOR2_X1   g766(.A1(new_n947), .A2(new_n952), .ZN(new_n953));
  NOR2_X1   g767(.A1(new_n949), .A2(new_n950), .ZN(new_n954));
  INV_X1    g768(.A(new_n954), .ZN(new_n955));
  NOR2_X1   g769(.A1(new_n953), .A2(new_n955), .ZN(new_n956));
  NOR3_X1   g770(.A1(new_n947), .A2(new_n952), .A3(new_n954), .ZN(new_n957));
  NOR2_X1   g771(.A1(new_n956), .A2(new_n957), .ZN(G66));
  NAND2_X1  g772(.A1(new_n509), .A2(new_n233), .ZN(new_n959));
  NAND2_X1  g773(.A1(new_n959), .A2(G953), .ZN(new_n960));
  OAI21_X1  g774(.A(new_n960), .B1(new_n821), .B2(G953), .ZN(new_n961));
  OAI21_X1  g775(.A(new_n906), .B1(G898), .B2(new_n234), .ZN(new_n962));
  XNOR2_X1  g776(.A(new_n961), .B(new_n962), .ZN(G69));
  OAI21_X1  g777(.A(G953), .B1(new_n305), .B2(new_n676), .ZN(new_n964));
  NAND2_X1  g778(.A1(new_n964), .A2(KEYINPUT126), .ZN(new_n965));
  OR2_X1    g779(.A1(new_n964), .A2(KEYINPUT126), .ZN(new_n966));
  INV_X1    g780(.A(new_n772), .ZN(new_n967));
  AND3_X1   g781(.A1(new_n569), .A2(new_n634), .A3(new_n743), .ZN(new_n968));
  INV_X1    g782(.A(new_n703), .ZN(new_n969));
  AOI21_X1  g783(.A(new_n969), .B1(new_n651), .B2(new_n813), .ZN(new_n970));
  NAND3_X1  g784(.A1(new_n968), .A2(KEYINPUT123), .A3(new_n970), .ZN(new_n971));
  AND2_X1   g785(.A1(new_n968), .A2(new_n970), .ZN(new_n972));
  OR2_X1    g786(.A1(new_n972), .A2(KEYINPUT123), .ZN(new_n973));
  AND3_X1   g787(.A1(new_n967), .A2(new_n971), .A3(new_n973), .ZN(new_n974));
  INV_X1    g788(.A(KEYINPUT100), .ZN(new_n975));
  XNOR2_X1  g789(.A(new_n707), .B(new_n975), .ZN(new_n976));
  OAI21_X1  g790(.A(KEYINPUT62), .B1(new_n976), .B2(new_n832), .ZN(new_n977));
  INV_X1    g791(.A(KEYINPUT62), .ZN(new_n978));
  NAND3_X1  g792(.A1(new_n708), .A2(new_n978), .A3(new_n834), .ZN(new_n979));
  NAND4_X1  g793(.A1(new_n974), .A2(new_n977), .A3(new_n781), .A4(new_n979), .ZN(new_n980));
  XOR2_X1   g794(.A(new_n595), .B(new_n436), .Z(new_n981));
  AND2_X1   g795(.A1(new_n981), .A2(new_n234), .ZN(new_n982));
  NAND2_X1  g796(.A1(new_n980), .A2(new_n982), .ZN(new_n983));
  INV_X1    g797(.A(new_n983), .ZN(new_n984));
  AOI21_X1  g798(.A(new_n981), .B1(new_n676), .B2(G953), .ZN(new_n985));
  INV_X1    g799(.A(new_n985), .ZN(new_n986));
  NAND3_X1  g800(.A1(new_n967), .A2(KEYINPUT124), .A3(new_n834), .ZN(new_n987));
  AND3_X1   g801(.A1(new_n781), .A2(new_n822), .A3(new_n750), .ZN(new_n988));
  NAND2_X1  g802(.A1(new_n747), .A2(new_n827), .ZN(new_n989));
  NOR2_X1   g803(.A1(new_n771), .A2(new_n989), .ZN(new_n990));
  XNOR2_X1  g804(.A(new_n990), .B(KEYINPUT125), .ZN(new_n991));
  INV_X1    g805(.A(KEYINPUT124), .ZN(new_n992));
  OAI21_X1  g806(.A(new_n992), .B1(new_n772), .B2(new_n832), .ZN(new_n993));
  NAND4_X1  g807(.A1(new_n987), .A2(new_n988), .A3(new_n991), .A4(new_n993), .ZN(new_n994));
  AOI21_X1  g808(.A(new_n986), .B1(new_n994), .B2(new_n234), .ZN(new_n995));
  OAI211_X1 g809(.A(new_n965), .B(new_n966), .C1(new_n984), .C2(new_n995), .ZN(new_n996));
  INV_X1    g810(.A(new_n995), .ZN(new_n997));
  NAND4_X1  g811(.A1(new_n997), .A2(KEYINPUT126), .A3(new_n983), .A4(new_n964), .ZN(new_n998));
  AND2_X1   g812(.A1(new_n996), .A2(new_n998), .ZN(G72));
  NAND2_X1  g813(.A1(new_n596), .A2(new_n573), .ZN(new_n1000));
  NAND2_X1  g814(.A1(G472), .A2(G902), .ZN(new_n1001));
  XOR2_X1   g815(.A(new_n1001), .B(KEYINPUT63), .Z(new_n1002));
  INV_X1    g816(.A(new_n821), .ZN(new_n1003));
  OAI21_X1  g817(.A(new_n1002), .B1(new_n994), .B2(new_n1003), .ZN(new_n1004));
  AOI21_X1  g818(.A(new_n1000), .B1(new_n1004), .B2(KEYINPUT127), .ZN(new_n1005));
  INV_X1    g819(.A(KEYINPUT127), .ZN(new_n1006));
  OAI211_X1 g820(.A(new_n1006), .B(new_n1002), .C1(new_n994), .C2(new_n1003), .ZN(new_n1007));
  NAND2_X1  g821(.A1(new_n1005), .A2(new_n1007), .ZN(new_n1008));
  OAI21_X1  g822(.A(new_n1002), .B1(new_n980), .B2(new_n1003), .ZN(new_n1009));
  AOI21_X1  g823(.A(new_n901), .B1(new_n1009), .B2(new_n697), .ZN(new_n1010));
  INV_X1    g824(.A(new_n697), .ZN(new_n1011));
  NAND4_X1  g825(.A1(new_n856), .A2(new_n1011), .A3(new_n1002), .A4(new_n1000), .ZN(new_n1012));
  AND3_X1   g826(.A1(new_n1008), .A2(new_n1010), .A3(new_n1012), .ZN(G57));
endmodule


